netcdf SN99880 {
dimensions:
	time = UNLIMITED ; // (59360 currently)
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Time of measurement" ;
		time:calendar = "standard" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:axis = "T" ;
	double latitude ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:units = "degree_north" ;
	double longitude ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:units = "degree_east" ;
	float air_temperature_2m(time) ;
		air_temperature_2m:long_name = "Air temperature" ;
		air_temperature_2m:coverage_content_type = "coordinate" ;
		air_temperature_2m:standard_name = "air_temperature" ;
		air_temperature_2m:units = "K" ;
	float air_pressure_at_sea_level(time) ;
		air_pressure_at_sea_level:long_name = "Air pressure at sea level" ;
		air_pressure_at_sea_level:coverage_content_type = "coordinate" ;
		air_pressure_at_sea_level:standard_name = "air_pressure_at_sea_level" ;
		air_pressure_at_sea_level:units = "Pa" ;
	float air_pressure_at_sea_level_qnh(time) ;
		air_pressure_at_sea_level_qnh:long_name = "Air pressure (QNH)" ;
		air_pressure_at_sea_level_qnh:coverage_content_type = "coordinate" ;
		air_pressure_at_sea_level_qnh:standard_name = "air_pressure_at_sea_level_qnh" ;
		air_pressure_at_sea_level_qnh:units = "hPa" ;
	float wind_speed_10m(time) ;
		wind_speed_10m:long_name = "Mean wind speed" ;
		wind_speed_10m:coverage_content_type = "coordinate" ;
		wind_speed_10m:standard_name = "wind_speed" ;
		wind_speed_10m:units = "m s-1" ;
	float relative_humidity(time) ;
		relative_humidity:long_name = "Relative air humidity" ;
		relative_humidity:coverage_content_type = "coordinate" ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:units = "1" ;
	float surface_air_pressure_2m(time) ;
		surface_air_pressure_2m:long_name = "Air pressure at station level" ;
		surface_air_pressure_2m:coverage_content_type = "coordinate" ;
		surface_air_pressure_2m:standard_name = "surface_air_pressure" ;
		surface_air_pressure_2m:units = "Pa" ;
	float wind_from_direction_10m(time) ;
		wind_from_direction_10m:long_name = "Wind direction" ;
		wind_from_direction_10m:coverage_content_type = "coordinate" ;
		wind_from_direction_10m:standard_name = "wind_from_direction" ;
		wind_from_direction_10m:units = "degree" ;

// global attributes:
		:station_name = "PYRAMIDEN" ;
		:wigos_identifier = "0-20000-0-01024" ;
		:wmo_identifier = "01024" ;
		:date_created = "2019-09-03T09:58:12.415858+00:00" ;
		:Conventions = "ACDD-1.3 CF-1.6" ;
		:title = "Observations from station PYRAMIDEN SN99880" ;
		:institution = "Norwegian Meteorological Institute" ;
		:source = "Meterological surface observation via frost.met.no" ;
		:history = "https://github.com/ferrighi/netcdf-ld-prototype/blob/master/files/data-provenance-sios.ttl" ;
		:references = "" ;
		:acknowledgment = "frost.met.no" ;
		:comment = "Observations based on data from frost.met.no" ;
		:creator_email = "observasjon@met.no" ;
		:creator_name = "Norwegian Meteorological Institute" ;
		:creator_url = "https://met.no" ;
		:geospatial_bounds = "POINT(16.360300 78.655700)" ;
		:geospatial_bounds_crs = "latlon" ;
		:geospatial_lat_max = "78.655700" ;
		:geospatial_lat_min = "78.655700" ;
		:geospatial_lon_max = "16.360300" ;
		:geospatial_lon_min = "16.360300" ;
		:id = "metno_obs_SN99880" ;
		:keywords = "observations" ;
		:metadata_link = "https://oaipmh.met.no/oai/?verb=GetRecord&metadataPrefix=iso&identifier=SN99880" ;
		:summary = "Surface meteorological observations from the observation network operated by the Norwegian Meteorological Institute. Data are received and quality controlled using the local KVALOBS system. Observation stations are normally operated according to WMO requirements, although specifications are not followed on some remote stations for practical matters. Stations may have more parameters than reported in this dataset." ;
		:time_coverage_start = "2012-11-16T10:00:00" ;
		:time_coverage_end = "2019-09-03T10:00:00" ;
		:featureType = "timeSeries" ;
}
