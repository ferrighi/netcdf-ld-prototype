netcdf SN99938 {
dimensions:
	time = UNLIMITED ; // (65718 currently)
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Time of measurement" ;
		time:calendar = "standard" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:axis = "T" ;
	double latitude ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:units = "degree_north" ;
	double longitude ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:units = "degree_east" ;
	float air_pressure_at_sea_level(time) ;
		air_pressure_at_sea_level:long_name = "Air pressure at sea level" ;
		air_pressure_at_sea_level:standard_name = "air_pressure_at_sea_level" ;
		air_pressure_at_sea_level:unit = "Pa" ;
	float surface_air_pressure_2m(time) ;
		surface_air_pressure_2m:long_name = "Air pressure at station level" ;
		surface_air_pressure_2m:standard_name = "surface_air_pressure" ;
		surface_air_pressure_2m:unit = "Pa" ;
	float air_temperature_2m(time) ;
		air_temperature_2m:long_name = "Air temperature" ;
		air_temperature_2m:standard_name = "air_temperature" ;
		air_temperature_2m:unit = "K" ;
	float air_pressure_at_sea_level_qnh(time) ;
		air_pressure_at_sea_level_qnh:long_name = "Air pressure (QNH)" ;
		air_pressure_at_sea_level_qnh:standard_name = "air_pressure_at_sea_level" ;
		air_pressure_at_sea_level_qnh:unit = "Pa" ;
	float wind_speed_10m(time) ;
		wind_speed_10m:long_name = "Mean wind speed" ;
		wind_speed_10m:standard_name = "wind_speed" ;
		wind_speed_10m:unit = "m s-1" ;
	float wind_from_direction_10m(time) ;
		wind_from_direction_10m:long_name = "Wind direction" ;
		wind_from_direction_10m:standard_name = "wind_from_direction" ;
		wind_from_direction_10m:unit = "degree" ;
	float relative_humidity(time) ;
		relative_humidity:long_name = "Relative air humidity" ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:unit = "1" ;

// global attributes:
		:wigos = "unknown" ;
		string :station_name = "KVITØYA" ;
		:wmo_identifier = "01011" ;
		:date_created = "2019-03-02T07:01:38.400294+00:00" ;
		:time_coverage_end = "2019-03-02T07:00:00" ;
		string :title = "Observations from station KVITØYA SN99938" ;
		:metadata_link = "https://oaipmh.met.no/oai/?verb=GetRecord&metadataPrefix=iso&identifier=SN99938" ;
		:acknowledgment = "frost.met.no" ;
		:comment = "Observations based on data from frost.met.no" ;
		:institution = "Norwegian Meteorological Institute" ;
		:featureType = "timeSeries" ;
		:id = "metno_obs_SN99938" ;
		:references = "" ;
		:geospatial_lat_min = "80.105800" ;
		:Conventions = "ACDD-1.3,CF-1.6" ;
		:creator_name = "Norwegian Meteorological Institute" ;
		:keywords = "observations" ;
		:history = "data-provenance-sios.ttl" ;
		:creator_url = "https://met.no" ;
		:geospatial_lon_max = "31.464300" ;
		:summary = "Surface meteorological observations from the observation network operated by the Norwegian Meteorological Institute. Data are received and quality controlled using the local KVALOBS system. Observation stations are normally operated according to WMO requirements, although specifications are not followed on some remote stations for practical matters. Stations may have more parameters than reported in this dataset." ;
		:geospatial_lon_min = "31.464300" ;
		:geospatial_bounds = "POINT(31.464300 80.105800)" ;
		:geospatial_lat_max = "80.105800" ;
		:creator_email = "observasjon@met.no" ;
		:geospatial_bounds_crs = "latlon" ;
		:source = "Meterological surface observation via frost.met.no" ;
		:time_coverage_start = "1996-01-01T03:00:00" ;
		:wigos_identifier = "unknown" ;
data:

 time = 820465200, 820486800, 820508400, 820551600, 820573200, 820594800, 
    820638000, 820659600, 820681200, 820724400, 820767600, 820810800, 
    820832400, 820854000, 820897200, 820918800, 820940400, 820983600, 
    821005200, 821026800, 821048400, 821091600, 821113200, 821156400, 
    821178000, 821199600, 821242800, 821264400, 821286000, 821329200, 
    821350800, 821372400, 821415600, 821437200, 821458800, 821523600, 
    821545200, 821588400, 821610000, 821631600, 821653200, 821696400, 
    821782800, 821804400, 821847600, 821869200, 821890800, 821934000, 
    821955600, 821977200, 822020400, 822042000, 822063600, 822128400, 
    822150000, 822214800, 822236400, 822279600, 822301200, 822366000, 
    822452400, 822474000, 822495600, 822517200, 822538800, 822560400, 
    822603600, 822625200, 822646800, 822668400, 822690000, 822711600, 
    822733200, 822754800, 822798000, 822819600, 822841200, 822884400, 
    822906000, 822927600, 822970800, 823014000, 823057200, 823078800, 
    823100400, 823143600, 823165200, 823186800, 823251600, 823273200, 
    823316400, 823338000, 823359600, 823381200, 823402800, 823424400, 
    823446000, 823467600, 823489200, 823510800, 823532400, 823575600, 
    823597200, 823662000, 823683600, 823705200, 823748400, 823770000, 
    823791600, 823834800, 823856400, 823878000, 823921200, 823964400, 
    824007600, 824029200, 824050800, 824072400, 824094000, 824115600, 
    824137200, 824158800, 824180400, 824223600, 824245200, 824266800, 
    824288400, 824310000, 824374800, 824396400, 824439600, 824461200, 
    824526000, 824547600, 824569200, 824634000, 824655600, 824720400, 
    824742000, 824806800, 824828400, 824850000, 824871600, 824979600, 
    825044400, 825066000, 991353600, 991364400, 991375200, 991386000, 
    991450800, 991461600, 991483200, 991494000, 991526400, 991537200, 
    991548000, 991569600, 991580400, 991623600, 991634400, 991656000, 
    991666800, 991710000, 991720800, 991742400, 991753200, 991796400, 
    991807200, 1009789200, 1096592400, 1096596000, 1096603200, 1096963200, 
    1099270800, 1099274400, 1099278000, 1101862800, 1101866400, 1104541200, 
    1107068400, 1107219600, 1107223200, 1109638800, 1109642400, 1109646000, 
    1109732400, 1112317200, 1112320800, 1112324400, 1112367600, 1114909200, 
    1114912800, 1114916400, 1114923600, 1114981200, 1115521200, 1313571600, 
    1313575200, 1313578800, 1313582400, 1313586000, 1313589600, 1313593200, 
    1313596800, 1313600400, 1313604000, 1313607600, 1313611200, 1313614800, 
    1313618400, 1313622000, 1313625600, 1313629200, 1313632800, 1313636400, 
    1313640000, 1313643600, 1313647200, 1313650800, 1313654400, 1313658000, 
    1313661600, 1313665200, 1313668800, 1313672400, 1313676000, 1313679600, 
    1313683200, 1313686800, 1313690400, 1313694000, 1313697600, 1313701200, 
    1313704800, 1313708400, 1313712000, 1313715600, 1313719200, 1313722800, 
    1313726400, 1313730000, 1313733600, 1313737200, 1313740800, 1313744400, 
    1313748000, 1313751600, 1313755200, 1313758800, 1313762400, 1313766000, 
    1313769600, 1313773200, 1313776800, 1313780400, 1313784000, 1313787600, 
    1313791200, 1313794800, 1313798400, 1313802000, 1313805600, 1313809200, 
    1313812800, 1313816400, 1313820000, 1313823600, 1313827200, 1313830800, 
    1313834400, 1313838000, 1313841600, 1313845200, 1313848800, 1313852400, 
    1313856000, 1313859600, 1313863200, 1313866800, 1313870400, 1313874000, 
    1313877600, 1313881200, 1313884800, 1313888400, 1313892000, 1313895600, 
    1313899200, 1313902800, 1313906400, 1313910000, 1313913600, 1313917200, 
    1313920800, 1313924400, 1313928000, 1313931600, 1313935200, 1313938800, 
    1313942400, 1313946000, 1313949600, 1313953200, 1313956800, 1313960400, 
    1313964000, 1313967600, 1313971200, 1313974800, 1313978400, 1313982000, 
    1313985600, 1313989200, 1313992800, 1313996400, 1314000000, 1314003600, 
    1314007200, 1314010800, 1314014400, 1314018000, 1314021600, 1314025200, 
    1314028800, 1314032400, 1314036000, 1314039600, 1314043200, 1314046800, 
    1314050400, 1314054000, 1314057600, 1314061200, 1314064800, 1314068400, 
    1314072000, 1314075600, 1314079200, 1314082800, 1314086400, 1314090000, 
    1314093600, 1314097200, 1314100800, 1314104400, 1314108000, 1314111600, 
    1314115200, 1314118800, 1314122400, 1314126000, 1314129600, 1314133200, 
    1314136800, 1314140400, 1314144000, 1314147600, 1314151200, 1314154800, 
    1314158400, 1314162000, 1314165600, 1314169200, 1314172800, 1314176400, 
    1314180000, 1314183600, 1314187200, 1314190800, 1314194400, 1314198000, 
    1314201600, 1314205200, 1314208800, 1314212400, 1314216000, 1314219600, 
    1314223200, 1314226800, 1314230400, 1314234000, 1314237600, 1314241200, 
    1314244800, 1314248400, 1314252000, 1314255600, 1314259200, 1314262800, 
    1314266400, 1314270000, 1314273600, 1314277200, 1314280800, 1314284400, 
    1314288000, 1314291600, 1314295200, 1314298800, 1314302400, 1314306000, 
    1314309600, 1314313200, 1314316800, 1314320400, 1314324000, 1314327600, 
    1314331200, 1314334800, 1314338400, 1314342000, 1314345600, 1314349200, 
    1314352800, 1314356400, 1314360000, 1314363600, 1314367200, 1314370800, 
    1314374400, 1314378000, 1314381600, 1314385200, 1314388800, 1314392400, 
    1314396000, 1314399600, 1314403200, 1314406800, 1314410400, 1314414000, 
    1314417600, 1314421200, 1314424800, 1314428400, 1314432000, 1314435600, 
    1314439200, 1314442800, 1314446400, 1314450000, 1314453600, 1314457200, 
    1314460800, 1314464400, 1314468000, 1314471600, 1314475200, 1314478800, 
    1314482400, 1314486000, 1314489600, 1314493200, 1314496800, 1314500400, 
    1314504000, 1314507600, 1314511200, 1314514800, 1314518400, 1314522000, 
    1314525600, 1314529200, 1314532800, 1314536400, 1314540000, 1314543600, 
    1314547200, 1314550800, 1314554400, 1314558000, 1314561600, 1314565200, 
    1314568800, 1314572400, 1314576000, 1314579600, 1314583200, 1314586800, 
    1314590400, 1314594000, 1314597600, 1314601200, 1314604800, 1314608400, 
    1314612000, 1314615600, 1314619200, 1314622800, 1314626400, 1314630000, 
    1314633600, 1314637200, 1314640800, 1314644400, 1314648000, 1314651600, 
    1314655200, 1314658800, 1314662400, 1314666000, 1314669600, 1314673200, 
    1314676800, 1314680400, 1314684000, 1314687600, 1314691200, 1314694800, 
    1314698400, 1314702000, 1314705600, 1314709200, 1314712800, 1314716400, 
    1314720000, 1314723600, 1314727200, 1314730800, 1314734400, 1314738000, 
    1314741600, 1314745200, 1314748800, 1314752400, 1314756000, 1314759600, 
    1314763200, 1314766800, 1314770400, 1314774000, 1314777600, 1314781200, 
    1314784800, 1314788400, 1314792000, 1314795600, 1314799200, 1314802800, 
    1314806400, 1314810000, 1314813600, 1314817200, 1314820800, 1314824400, 
    1314828000, 1314831600, 1314835200, 1314838800, 1314842400, 1314846000, 
    1314849600, 1314853200, 1314856800, 1314860400, 1314864000, 1314867600, 
    1314871200, 1314874800, 1314878400, 1314882000, 1314885600, 1314889200, 
    1314892800, 1314896400, 1314900000, 1314903600, 1314907200, 1314910800, 
    1314914400, 1314918000, 1314921600, 1314925200, 1314928800, 1314932400, 
    1314936000, 1314939600, 1314943200, 1314946800, 1314950400, 1314954000, 
    1314957600, 1314961200, 1314964800, 1314968400, 1314972000, 1314975600, 
    1314979200, 1314982800, 1314986400, 1314990000, 1314993600, 1314997200, 
    1315000800, 1315004400, 1315008000, 1315011600, 1315015200, 1315018800, 
    1315022400, 1315026000, 1315029600, 1315033200, 1315036800, 1315040400, 
    1315044000, 1315047600, 1315051200, 1315054800, 1315058400, 1315062000, 
    1315065600, 1315069200, 1315072800, 1315076400, 1315080000, 1315083600, 
    1315087200, 1315090800, 1315094400, 1315098000, 1315101600, 1315105200, 
    1315108800, 1315112400, 1315116000, 1315119600, 1315123200, 1315126800, 
    1315130400, 1315134000, 1315137600, 1315141200, 1315144800, 1315148400, 
    1315152000, 1315155600, 1315159200, 1315162800, 1315166400, 1315170000, 
    1315173600, 1315177200, 1315180800, 1315184400, 1315188000, 1315191600, 
    1315195200, 1315198800, 1315202400, 1315206000, 1315209600, 1315213200, 
    1315216800, 1315220400, 1315224000, 1315227600, 1315231200, 1315234800, 
    1315238400, 1315242000, 1315245600, 1315249200, 1315252800, 1315256400, 
    1315260000, 1315263600, 1315267200, 1315270800, 1315274400, 1315278000, 
    1315281600, 1315285200, 1315288800, 1315292400, 1315296000, 1315299600, 
    1315303200, 1315306800, 1315310400, 1315314000, 1315317600, 1315321200, 
    1315324800, 1315328400, 1315332000, 1315335600, 1315339200, 1315342800, 
    1315346400, 1315350000, 1315353600, 1315357200, 1315360800, 1315364400, 
    1315368000, 1315371600, 1315375200, 1315378800, 1315382400, 1315386000, 
    1315389600, 1315393200, 1315396800, 1315400400, 1315404000, 1315407600, 
    1315411200, 1315414800, 1315418400, 1315422000, 1315425600, 1315429200, 
    1315432800, 1315436400, 1315440000, 1315443600, 1315447200, 1315450800, 
    1315454400, 1315458000, 1315461600, 1315465200, 1315468800, 1315472400, 
    1315476000, 1315479600, 1315483200, 1315486800, 1315490400, 1315494000, 
    1315497600, 1315501200, 1315504800, 1315508400, 1315512000, 1315515600, 
    1315519200, 1315522800, 1315526400, 1315530000, 1315533600, 1315537200, 
    1315540800, 1315544400, 1315548000, 1315551600, 1315555200, 1315558800, 
    1315562400, 1315566000, 1315569600, 1315573200, 1315576800, 1315580400, 
    1315584000, 1315587600, 1315591200, 1315594800, 1315598400, 1315602000, 
    1315605600, 1315609200, 1315612800, 1315616400, 1315620000, 1315623600, 
    1315627200, 1315630800, 1315634400, 1315638000, 1315641600, 1315645200, 
    1315648800, 1315652400, 1315656000, 1315659600, 1315663200, 1315666800, 
    1315670400, 1315674000, 1315677600, 1315681200, 1315684800, 1315688400, 
    1315692000, 1315695600, 1315699200, 1315702800, 1315706400, 1315710000, 
    1315713600, 1315717200, 1315720800, 1315724400, 1315728000, 1315731600, 
    1315735200, 1315738800, 1315742400, 1315746000, 1315749600, 1315753200, 
    1315756800, 1315760400, 1315764000, 1315767600, 1315771200, 1315774800, 
    1315778400, 1315782000, 1315785600, 1315789200, 1315792800, 1315796400, 
    1315800000, 1315803600, 1315807200, 1315810800, 1315814400, 1315818000, 
    1315821600, 1315825200, 1315828800, 1315832400, 1315836000, 1315839600, 
    1315843200, 1315846800, 1315850400, 1315854000, 1315857600, 1315861200, 
    1315864800, 1315868400, 1315872000, 1315875600, 1315879200, 1315882800, 
    1315886400, 1315890000, 1315893600, 1315897200, 1315900800, 1315904400, 
    1315908000, 1315911600, 1315915200, 1315918800, 1315922400, 1315926000, 
    1315929600, 1315933200, 1315936800, 1315940400, 1315944000, 1315947600, 
    1315951200, 1315954800, 1315958400, 1315962000, 1315965600, 1315969200, 
    1315972800, 1315976400, 1315980000, 1315983600, 1315987200, 1315990800, 
    1315994400, 1315998000, 1316001600, 1316005200, 1316008800, 1316012400, 
    1316016000, 1316019600, 1316023200, 1316026800, 1316030400, 1316034000, 
    1316037600, 1316041200, 1316044800, 1316048400, 1316052000, 1316055600, 
    1316059200, 1316062800, 1316066400, 1316070000, 1316073600, 1316077200, 
    1316080800, 1316084400, 1316088000, 1316091600, 1316095200, 1316098800, 
    1316102400, 1316106000, 1316109600, 1316113200, 1316116800, 1316120400, 
    1316124000, 1316127600, 1316131200, 1316134800, 1316138400, 1316142000, 
    1316145600, 1316149200, 1316152800, 1316156400, 1316160000, 1316163600, 
    1316167200, 1316170800, 1316174400, 1316178000, 1316181600, 1316185200, 
    1316188800, 1316192400, 1316196000, 1316199600, 1316203200, 1316206800, 
    1316210400, 1316214000, 1316217600, 1316221200, 1316224800, 1316228400, 
    1316232000, 1316235600, 1316239200, 1316242800, 1316246400, 1316250000, 
    1316253600, 1316257200, 1316260800, 1316264400, 1316268000, 1316271600, 
    1316275200, 1316278800, 1316282400, 1316286000, 1316289600, 1316293200, 
    1316296800, 1316300400, 1316304000, 1316307600, 1316311200, 1316314800, 
    1316318400, 1316322000, 1316325600, 1316329200, 1316332800, 1316336400, 
    1316340000, 1316343600, 1316347200, 1316350800, 1316354400, 1316358000, 
    1316361600, 1316365200, 1316368800, 1316372400, 1316376000, 1316379600, 
    1316383200, 1316386800, 1316390400, 1316394000, 1316397600, 1316401200, 
    1316404800, 1316408400, 1316412000, 1316415600, 1316419200, 1316422800, 
    1316426400, 1316430000, 1316433600, 1316437200, 1316440800, 1316444400, 
    1316448000, 1316451600, 1316455200, 1316458800, 1316462400, 1316466000, 
    1316469600, 1316473200, 1316476800, 1316480400, 1316484000, 1316487600, 
    1316491200, 1316494800, 1316498400, 1316502000, 1316505600, 1316509200, 
    1316512800, 1316516400, 1316520000, 1316523600, 1316527200, 1316530800, 
    1316534400, 1316538000, 1316541600, 1316545200, 1316548800, 1316552400, 
    1316556000, 1316559600, 1316563200, 1316566800, 1316570400, 1316574000, 
    1316577600, 1316581200, 1316584800, 1316588400, 1316592000, 1316595600, 
    1316599200, 1316602800, 1316606400, 1316610000, 1316613600, 1316617200, 
    1316620800, 1316624400, 1316628000, 1316631600, 1316635200, 1316638800, 
    1316642400, 1316646000, 1316649600, 1316653200, 1316656800, 1316660400, 
    1316664000, 1316667600, 1316671200, 1316674800, 1316678400, 1316682000, 
    1316685600, 1316689200, 1316692800, 1316696400, 1316700000, 1316703600, 
    1316707200, 1316710800, 1316714400, 1316718000, 1316721600, 1316725200, 
    1316728800, 1316732400, 1316736000, 1316739600, 1316743200, 1316746800, 
    1316750400, 1316754000, 1316757600, 1316761200, 1316764800, 1316768400, 
    1316772000, 1316775600, 1316779200, 1316782800, 1316786400, 1316790000, 
    1316793600, 1316797200, 1316800800, 1316804400, 1316808000, 1316811600, 
    1316815200, 1316818800, 1316822400, 1316826000, 1316829600, 1316833200, 
    1316836800, 1316840400, 1316844000, 1316847600, 1316851200, 1316854800, 
    1316858400, 1316862000, 1316865600, 1316869200, 1316872800, 1316876400, 
    1316880000, 1316883600, 1316887200, 1316890800, 1316894400, 1316898000, 
    1316901600, 1316905200, 1316908800, 1316912400, 1316916000, 1316919600, 
    1316923200, 1316926800, 1316930400, 1316934000, 1316937600, 1316941200, 
    1316944800, 1316948400, 1316952000, 1316955600, 1316959200, 1316962800, 
    1316966400, 1316970000, 1316973600, 1316977200, 1316980800, 1316984400, 
    1316988000, 1316991600, 1316995200, 1316998800, 1317002400, 1317006000, 
    1317009600, 1317013200, 1317016800, 1317020400, 1317024000, 1317027600, 
    1317031200, 1317034800, 1317038400, 1317042000, 1317045600, 1317049200, 
    1317052800, 1317056400, 1317060000, 1317063600, 1317067200, 1317070800, 
    1317074400, 1317078000, 1317081600, 1317085200, 1317088800, 1317092400, 
    1317096000, 1317099600, 1317103200, 1317106800, 1317110400, 1317114000, 
    1317117600, 1317121200, 1317124800, 1317128400, 1317132000, 1317135600, 
    1317139200, 1317142800, 1317146400, 1317150000, 1317153600, 1317157200, 
    1317160800, 1317164400, 1317168000, 1317171600, 1317175200, 1317178800, 
    1317182400, 1317186000, 1317189600, 1317193200, 1317196800, 1317200400, 
    1317204000, 1317207600, 1317211200, 1317214800, 1317218400, 1317222000, 
    1317225600, 1317229200, 1317232800, 1317236400, 1317240000, 1317243600, 
    1317247200, 1317250800, 1317254400, 1317258000, 1317261600, 1317265200, 
    1317268800, 1317272400, 1317276000, 1317279600, 1317283200, 1317286800, 
    1317290400, 1317294000, 1317297600, 1317301200, 1317304800, 1317308400, 
    1317312000, 1317315600, 1317319200, 1317322800, 1317326400, 1317330000, 
    1317333600, 1317337200, 1317340800, 1317344400, 1317348000, 1317351600, 
    1317355200, 1317358800, 1317362400, 1317366000, 1317369600, 1317373200, 
    1317376800, 1317380400, 1317384000, 1317387600, 1317391200, 1317394800, 
    1317398400, 1317402000, 1317405600, 1317409200, 1317412800, 1317416400, 
    1317420000, 1317423600, 1317427200, 1317430800, 1317434400, 1317438000, 
    1317441600, 1317445200, 1317448800, 1317452400, 1317456000, 1317459600, 
    1317463200, 1317466800, 1317470400, 1317474000, 1317477600, 1317481200, 
    1317484800, 1317488400, 1317492000, 1317495600, 1317499200, 1317502800, 
    1317506400, 1317510000, 1317513600, 1317517200, 1317520800, 1317524400, 
    1317528000, 1317531600, 1317535200, 1317538800, 1317542400, 1317546000, 
    1317549600, 1317553200, 1317556800, 1317560400, 1317564000, 1317567600, 
    1317571200, 1317574800, 1317578400, 1317582000, 1317585600, 1317589200, 
    1317592800, 1317596400, 1317600000, 1317603600, 1317607200, 1317610800, 
    1317614400, 1317618000, 1317621600, 1317625200, 1317628800, 1317632400, 
    1317636000, 1317639600, 1317643200, 1317646800, 1317650400, 1317654000, 
    1317657600, 1317661200, 1317664800, 1317668400, 1317672000, 1317675600, 
    1317679200, 1317682800, 1317686400, 1317690000, 1317693600, 1317697200, 
    1317700800, 1317704400, 1317708000, 1317711600, 1317715200, 1317718800, 
    1317722400, 1317726000, 1317729600, 1317733200, 1317736800, 1317740400, 
    1317744000, 1317747600, 1317751200, 1317754800, 1317758400, 1317762000, 
    1317765600, 1317769200, 1317772800, 1317776400, 1317780000, 1317783600, 
    1317787200, 1317790800, 1317794400, 1317798000, 1317801600, 1317805200, 
    1317808800, 1317812400, 1317816000, 1317819600, 1317823200, 1317826800, 
    1317830400, 1317834000, 1317837600, 1317841200, 1317844800, 1317848400, 
    1317852000, 1317855600, 1317859200, 1317862800, 1317866400, 1317870000, 
    1317873600, 1317877200, 1317880800, 1317884400, 1317888000, 1317891600, 
    1317895200, 1317898800, 1317902400, 1317906000, 1317909600, 1317913200, 
    1317916800, 1317920400, 1317924000, 1317927600, 1317931200, 1317934800, 
    1317938400, 1317942000, 1317945600, 1317949200, 1317952800, 1317956400, 
    1317960000, 1317963600, 1317967200, 1317970800, 1317974400, 1317978000, 
    1317981600, 1317985200, 1317988800, 1317992400, 1317996000, 1317999600, 
    1318003200, 1318006800, 1318010400, 1318014000, 1318017600, 1318021200, 
    1318024800, 1318028400, 1318032000, 1318035600, 1318039200, 1318042800, 
    1318046400, 1318050000, 1318053600, 1318057200, 1318060800, 1318064400, 
    1318068000, 1318071600, 1318075200, 1318078800, 1318082400, 1318086000, 
    1318089600, 1318093200, 1318096800, 1318100400, 1318104000, 1318107600, 
    1318111200, 1318114800, 1318118400, 1318122000, 1318125600, 1318129200, 
    1318132800, 1318136400, 1318140000, 1318143600, 1318147200, 1318150800, 
    1318154400, 1318158000, 1318161600, 1318165200, 1318168800, 1318172400, 
    1318176000, 1318179600, 1318183200, 1318186800, 1318190400, 1318194000, 
    1318197600, 1318201200, 1318204800, 1318208400, 1318212000, 1318215600, 
    1318219200, 1318222800, 1318226400, 1318230000, 1318233600, 1318237200, 
    1318240800, 1318244400, 1318248000, 1318251600, 1318255200, 1318258800, 
    1318262400, 1318266000, 1318269600, 1318273200, 1318276800, 1318280400, 
    1318284000, 1318287600, 1318291200, 1318294800, 1318298400, 1318302000, 
    1318305600, 1318309200, 1318312800, 1318316400, 1318320000, 1318323600, 
    1318327200, 1318330800, 1318334400, 1318338000, 1318341600, 1318345200, 
    1318348800, 1318352400, 1318356000, 1318359600, 1318363200, 1318366800, 
    1318370400, 1318374000, 1318377600, 1318381200, 1318384800, 1318388400, 
    1318392000, 1318395600, 1318399200, 1318402800, 1318406400, 1318410000, 
    1318413600, 1318417200, 1318420800, 1318424400, 1318428000, 1318431600, 
    1318435200, 1318438800, 1318442400, 1318446000, 1318449600, 1318453200, 
    1318456800, 1318460400, 1318464000, 1318467600, 1318471200, 1318474800, 
    1318478400, 1318482000, 1318485600, 1318489200, 1318492800, 1318496400, 
    1318500000, 1318503600, 1318507200, 1318510800, 1318514400, 1318518000, 
    1318521600, 1318525200, 1318528800, 1318532400, 1318536000, 1318539600, 
    1318543200, 1318546800, 1318550400, 1318554000, 1318557600, 1318561200, 
    1318564800, 1318568400, 1318572000, 1318575600, 1318579200, 1318582800, 
    1318586400, 1318590000, 1318593600, 1318597200, 1318600800, 1318604400, 
    1318608000, 1318611600, 1318615200, 1318618800, 1318622400, 1318626000, 
    1318629600, 1318633200, 1318636800, 1318640400, 1318644000, 1318647600, 
    1318651200, 1318654800, 1318658400, 1318662000, 1318665600, 1318669200, 
    1318672800, 1318676400, 1318680000, 1318683600, 1318687200, 1318690800, 
    1318694400, 1318698000, 1318701600, 1318705200, 1318708800, 1318712400, 
    1318716000, 1318719600, 1318723200, 1318726800, 1318730400, 1318734000, 
    1318737600, 1318741200, 1318744800, 1318748400, 1318752000, 1318755600, 
    1318759200, 1318762800, 1318766400, 1318770000, 1318773600, 1318777200, 
    1318780800, 1318784400, 1318788000, 1318791600, 1318795200, 1318798800, 
    1318802400, 1318806000, 1318809600, 1318813200, 1318816800, 1318820400, 
    1318824000, 1318827600, 1318831200, 1318834800, 1318838400, 1318842000, 
    1318845600, 1318849200, 1318852800, 1318856400, 1318860000, 1318863600, 
    1318867200, 1318870800, 1318874400, 1318878000, 1318881600, 1318885200, 
    1318888800, 1318892400, 1318896000, 1318899600, 1318903200, 1318906800, 
    1318910400, 1318914000, 1318917600, 1318921200, 1318924800, 1318928400, 
    1318932000, 1318935600, 1318939200, 1318942800, 1318946400, 1318950000, 
    1318953600, 1318957200, 1318960800, 1318964400, 1318968000, 1318971600, 
    1318975200, 1318978800, 1318982400, 1318986000, 1318989600, 1318993200, 
    1318996800, 1319000400, 1319004000, 1319007600, 1319011200, 1319014800, 
    1319018400, 1319022000, 1319025600, 1319029200, 1319032800, 1319036400, 
    1319040000, 1319043600, 1319047200, 1319050800, 1319054400, 1319058000, 
    1319061600, 1319065200, 1319068800, 1319072400, 1319076000, 1319079600, 
    1319083200, 1319086800, 1319090400, 1319094000, 1319097600, 1319101200, 
    1319104800, 1319108400, 1319112000, 1319115600, 1319119200, 1319122800, 
    1319126400, 1319130000, 1319133600, 1319137200, 1319140800, 1319144400, 
    1319148000, 1319151600, 1319155200, 1319158800, 1319162400, 1319166000, 
    1319169600, 1319173200, 1319176800, 1319180400, 1319184000, 1319187600, 
    1319191200, 1319194800, 1319198400, 1319202000, 1319205600, 1319209200, 
    1319212800, 1319216400, 1319220000, 1319223600, 1319227200, 1319230800, 
    1319234400, 1319238000, 1319241600, 1319245200, 1319248800, 1319252400, 
    1319256000, 1319259600, 1319263200, 1319266800, 1319270400, 1319274000, 
    1319277600, 1319281200, 1319284800, 1319288400, 1319292000, 1319295600, 
    1319299200, 1319302800, 1319306400, 1319310000, 1319313600, 1319317200, 
    1319320800, 1319324400, 1319328000, 1319331600, 1319335200, 1319338800, 
    1319342400, 1319346000, 1319349600, 1319353200, 1319356800, 1319360400, 
    1319364000, 1319367600, 1319371200, 1319374800, 1319378400, 1319382000, 
    1319385600, 1319389200, 1319392800, 1319396400, 1319400000, 1319403600, 
    1319407200, 1319410800, 1319414400, 1319418000, 1319421600, 1319425200, 
    1319428800, 1319432400, 1319436000, 1319439600, 1319443200, 1319446800, 
    1319450400, 1319454000, 1319457600, 1319461200, 1319464800, 1319468400, 
    1319472000, 1319475600, 1319479200, 1319482800, 1319486400, 1319490000, 
    1319493600, 1319497200, 1319500800, 1319504400, 1319508000, 1319511600, 
    1319515200, 1319518800, 1319522400, 1319526000, 1319529600, 1319533200, 
    1319536800, 1319540400, 1319544000, 1319547600, 1319551200, 1319554800, 
    1319558400, 1319562000, 1319565600, 1319569200, 1319572800, 1319576400, 
    1319580000, 1319583600, 1319587200, 1319590800, 1319594400, 1319598000, 
    1319601600, 1319605200, 1319608800, 1319612400, 1319616000, 1319619600, 
    1319623200, 1319626800, 1319630400, 1319634000, 1319637600, 1319641200, 
    1319644800, 1319648400, 1319652000, 1319655600, 1319659200, 1319662800, 
    1319666400, 1319670000, 1319673600, 1319677200, 1319680800, 1319684400, 
    1319688000, 1319691600, 1319695200, 1319698800, 1319702400, 1319706000, 
    1319709600, 1319713200, 1319716800, 1319720400, 1319724000, 1319727600, 
    1319731200, 1319734800, 1319738400, 1319742000, 1319745600, 1319749200, 
    1319752800, 1319756400, 1319760000, 1319763600, 1319767200, 1319770800, 
    1319774400, 1319778000, 1319781600, 1319785200, 1319788800, 1319792400, 
    1319796000, 1319799600, 1319803200, 1319806800, 1319810400, 1319814000, 
    1319817600, 1319821200, 1319824800, 1319828400, 1319832000, 1319835600, 
    1319839200, 1319842800, 1319846400, 1319850000, 1319853600, 1319857200, 
    1319860800, 1319864400, 1319868000, 1319871600, 1319875200, 1319878800, 
    1319882400, 1319886000, 1319889600, 1319893200, 1319896800, 1319900400, 
    1319904000, 1319907600, 1319911200, 1319914800, 1319918400, 1319922000, 
    1319925600, 1319929200, 1319932800, 1319936400, 1319940000, 1319943600, 
    1319947200, 1319950800, 1319954400, 1319958000, 1319961600, 1319965200, 
    1319968800, 1319972400, 1319976000, 1319979600, 1319983200, 1319986800, 
    1319990400, 1319994000, 1319997600, 1320001200, 1320004800, 1320008400, 
    1320012000, 1320015600, 1320019200, 1320022800, 1320026400, 1320030000, 
    1320033600, 1320037200, 1320040800, 1320044400, 1320048000, 1320051600, 
    1320055200, 1320058800, 1320062400, 1320066000, 1320069600, 1320073200, 
    1320076800, 1320080400, 1320084000, 1320087600, 1320091200, 1320094800, 
    1320098400, 1320102000, 1320105600, 1320109200, 1320112800, 1320116400, 
    1320120000, 1320123600, 1320127200, 1320130800, 1320134400, 1320138000, 
    1320141600, 1320145200, 1320148800, 1320152400, 1320156000, 1320159600, 
    1320163200, 1320166800, 1320170400, 1320174000, 1320177600, 1320181200, 
    1320184800, 1320188400, 1320192000, 1320195600, 1320199200, 1320202800, 
    1320206400, 1320210000, 1320213600, 1320217200, 1320220800, 1320224400, 
    1320228000, 1320231600, 1320235200, 1320238800, 1320242400, 1320246000, 
    1320249600, 1320253200, 1320256800, 1320260400, 1320264000, 1320267600, 
    1320271200, 1320274800, 1320278400, 1320282000, 1320285600, 1320289200, 
    1320292800, 1320296400, 1320300000, 1320303600, 1320307200, 1320310800, 
    1320314400, 1320318000, 1320321600, 1320325200, 1320328800, 1320332400, 
    1320336000, 1320339600, 1320343200, 1320346800, 1320350400, 1320354000, 
    1320357600, 1320361200, 1320364800, 1320368400, 1320372000, 1320375600, 
    1320379200, 1320382800, 1320386400, 1320390000, 1320393600, 1320397200, 
    1320400800, 1320404400, 1320408000, 1320411600, 1320415200, 1320418800, 
    1320422400, 1320426000, 1320429600, 1320433200, 1320436800, 1320440400, 
    1320444000, 1320447600, 1320451200, 1320454800, 1320458400, 1320462000, 
    1320465600, 1320469200, 1320472800, 1320476400, 1320480000, 1320483600, 
    1320487200, 1320490800, 1320494400, 1320498000, 1320501600, 1320505200, 
    1320508800, 1320512400, 1320516000, 1320519600, 1320523200, 1320526800, 
    1320530400, 1320534000, 1320537600, 1320541200, 1320544800, 1320548400, 
    1320552000, 1320555600, 1320559200, 1320562800, 1320566400, 1320570000, 
    1320573600, 1320577200, 1320580800, 1320584400, 1320588000, 1320591600, 
    1320595200, 1320598800, 1320602400, 1320606000, 1320609600, 1320613200, 
    1320616800, 1320620400, 1320624000, 1320627600, 1320631200, 1320634800, 
    1320638400, 1320642000, 1320645600, 1320649200, 1320652800, 1320656400, 
    1320660000, 1320663600, 1320667200, 1320670800, 1320674400, 1320678000, 
    1320681600, 1320685200, 1320688800, 1320692400, 1320696000, 1320699600, 
    1320703200, 1320706800, 1320710400, 1320714000, 1320717600, 1320721200, 
    1320724800, 1320728400, 1320732000, 1320735600, 1320739200, 1320742800, 
    1320746400, 1320750000, 1320753600, 1320757200, 1320760800, 1320764400, 
    1320768000, 1320771600, 1320775200, 1320778800, 1320782400, 1320786000, 
    1320789600, 1320793200, 1320796800, 1320800400, 1320804000, 1320807600, 
    1320811200, 1320814800, 1320818400, 1320822000, 1320825600, 1320829200, 
    1320832800, 1320836400, 1320840000, 1320843600, 1320847200, 1320850800, 
    1320854400, 1320858000, 1320861600, 1320865200, 1320868800, 1320872400, 
    1320876000, 1320879600, 1320883200, 1320886800, 1320890400, 1320894000, 
    1320897600, 1320901200, 1320904800, 1320908400, 1320912000, 1320915600, 
    1320919200, 1320922800, 1320926400, 1320930000, 1320933600, 1320937200, 
    1321362000, 1321365600, 1321369200, 1321372800, 1321376400, 1321380000, 
    1321383600, 1321387200, 1321390800, 1321394400, 1321398000, 1321401600, 
    1321405200, 1321408800, 1321412400, 1321416000, 1321419600, 1321423200, 
    1321426800, 1321430400, 1321434000, 1321437600, 1321441200, 1321444800, 
    1321448400, 1321452000, 1321455600, 1321459200, 1321462800, 1321466400, 
    1321470000, 1321473600, 1321477200, 1321480800, 1321484400, 1321488000, 
    1321491600, 1321495200, 1321498800, 1321502400, 1321506000, 1321509600, 
    1321513200, 1321516800, 1321520400, 1321524000, 1321527600, 1321531200, 
    1321534800, 1321538400, 1321542000, 1321545600, 1321549200, 1321552800, 
    1321556400, 1321560000, 1321563600, 1321567200, 1321570800, 1321574400, 
    1321578000, 1321581600, 1321585200, 1321588800, 1321592400, 1321596000, 
    1321599600, 1321603200, 1321606800, 1321610400, 1321614000, 1321617600, 
    1321621200, 1321624800, 1321628400, 1321632000, 1321635600, 1321639200, 
    1321642800, 1321646400, 1321650000, 1321653600, 1321657200, 1321660800, 
    1321664400, 1321668000, 1321671600, 1321675200, 1321678800, 1321682400, 
    1321686000, 1321689600, 1321693200, 1321696800, 1321700400, 1321704000, 
    1321707600, 1321711200, 1321714800, 1321718400, 1321722000, 1321725600, 
    1321729200, 1321732800, 1321736400, 1321740000, 1321743600, 1321747200, 
    1321750800, 1321754400, 1321758000, 1321761600, 1321765200, 1321768800, 
    1321772400, 1321776000, 1321779600, 1321783200, 1321786800, 1321790400, 
    1321794000, 1321797600, 1321801200, 1321804800, 1321808400, 1321812000, 
    1321815600, 1321819200, 1321822800, 1321826400, 1321830000, 1321833600, 
    1321837200, 1321840800, 1321844400, 1321848000, 1321851600, 1321855200, 
    1321858800, 1321862400, 1321866000, 1321869600, 1321873200, 1321876800, 
    1321880400, 1321884000, 1321887600, 1321891200, 1321894800, 1321898400, 
    1321902000, 1321905600, 1321909200, 1321912800, 1321916400, 1321920000, 
    1321923600, 1321927200, 1321930800, 1321934400, 1321938000, 1321941600, 
    1321945200, 1321948800, 1321952400, 1321956000, 1321959600, 1321963200, 
    1321966800, 1321970400, 1321974000, 1321977600, 1321981200, 1321984800, 
    1321988400, 1321992000, 1321995600, 1321999200, 1322002800, 1322053200, 
    1322056800, 1322060400, 1322064000, 1322067600, 1322071200, 1322074800, 
    1322078400, 1322082000, 1322085600, 1322089200, 1322092800, 1322096400, 
    1322100000, 1322103600, 1322107200, 1322110800, 1322114400, 1322118000, 
    1322121600, 1322125200, 1322128800, 1322132400, 1322136000, 1322139600, 
    1322143200, 1322146800, 1322150400, 1322154000, 1322157600, 1322161200, 
    1322164800, 1322168400, 1322172000, 1322175600, 1322179200, 1322182800, 
    1322186400, 1322190000, 1322193600, 1322197200, 1322200800, 1322204400, 
    1322208000, 1322211600, 1322215200, 1322218800, 1322222400, 1322226000, 
    1322229600, 1322233200, 1322236800, 1322240400, 1322244000, 1322247600, 
    1322251200, 1322254800, 1322258400, 1322262000, 1322265600, 1322269200, 
    1322272800, 1322276400, 1322280000, 1322283600, 1322287200, 1322290800, 
    1322294400, 1322298000, 1322301600, 1322305200, 1322308800, 1322312400, 
    1322316000, 1322319600, 1322323200, 1322326800, 1322330400, 1322334000, 
    1322337600, 1322341200, 1322344800, 1322348400, 1322352000, 1322355600, 
    1322359200, 1322362800, 1322366400, 1322370000, 1322373600, 1322377200, 
    1322380800, 1322384400, 1322388000, 1322391600, 1322395200, 1322398800, 
    1322402400, 1322406000, 1322409600, 1322413200, 1322416800, 1322420400, 
    1322424000, 1322427600, 1322431200, 1322434800, 1322438400, 1322442000, 
    1322445600, 1322449200, 1322452800, 1322456400, 1322460000, 1322463600, 
    1322467200, 1322470800, 1322474400, 1322478000, 1322481600, 1322485200, 
    1322488800, 1322492400, 1322496000, 1322499600, 1322503200, 1322506800, 
    1322510400, 1322514000, 1322517600, 1322521200, 1322524800, 1322528400, 
    1322532000, 1322535600, 1322539200, 1322542800, 1322546400, 1322550000, 
    1322553600, 1322557200, 1322560800, 1322564400, 1322568000, 1322571600, 
    1322575200, 1322578800, 1322582400, 1322586000, 1322589600, 1322593200, 
    1322596800, 1322600400, 1322604000, 1322607600, 1322611200, 1322614800, 
    1322618400, 1322622000, 1322625600, 1322629200, 1322632800, 1322636400, 
    1322640000, 1322643600, 1322647200, 1322650800, 1322654400, 1322658000, 
    1322661600, 1322665200, 1322668800, 1322672400, 1322676000, 1322679600, 
    1322683200, 1322686800, 1322690400, 1322694000, 1322697600, 1322701200, 
    1322704800, 1322708400, 1322712000, 1322715600, 1322719200, 1322722800, 
    1322726400, 1322730000, 1322733600, 1322737200, 1322740800, 1322744400, 
    1322748000, 1322751600, 1322755200, 1322758800, 1322762400, 1322766000, 
    1322769600, 1322773200, 1322776800, 1322780400, 1322784000, 1322787600, 
    1322791200, 1322794800, 1322798400, 1322802000, 1322805600, 1322809200, 
    1322812800, 1322816400, 1322820000, 1322823600, 1322827200, 1322830800, 
    1322834400, 1322838000, 1322841600, 1322845200, 1322848800, 1322852400, 
    1322856000, 1322859600, 1322863200, 1322866800, 1322870400, 1322874000, 
    1322877600, 1322881200, 1322884800, 1322888400, 1322892000, 1322895600, 
    1322899200, 1322902800, 1322906400, 1322910000, 1322913600, 1322917200, 
    1322920800, 1322924400, 1322928000, 1322931600, 1322935200, 1322938800, 
    1322942400, 1322946000, 1322949600, 1322953200, 1322956800, 1322960400, 
    1322964000, 1322967600, 1322971200, 1322974800, 1322978400, 1322982000, 
    1322985600, 1322989200, 1322992800, 1322996400, 1323000000, 1323003600, 
    1323007200, 1323010800, 1323014400, 1323018000, 1323021600, 1323025200, 
    1323028800, 1323032400, 1323036000, 1323039600, 1323043200, 1323046800, 
    1323050400, 1323054000, 1323057600, 1323061200, 1323064800, 1323068400, 
    1323072000, 1323075600, 1323079200, 1323082800, 1323086400, 1323090000, 
    1323093600, 1323097200, 1323100800, 1323104400, 1323108000, 1323111600, 
    1323115200, 1323118800, 1323122400, 1323126000, 1323129600, 1323133200, 
    1323136800, 1323140400, 1323144000, 1323147600, 1323151200, 1323154800, 
    1323158400, 1323162000, 1323165600, 1323169200, 1323172800, 1323176400, 
    1323180000, 1323183600, 1323187200, 1323190800, 1323194400, 1323198000, 
    1323201600, 1323205200, 1323208800, 1323212400, 1323435600, 1323439200, 
    1323442800, 1323446400, 1323450000, 1323453600, 1323457200, 1323460800, 
    1323464400, 1323468000, 1323471600, 1323475200, 1323478800, 1323482400, 
    1323486000, 1323489600, 1323493200, 1323496800, 1323500400, 1323504000, 
    1323507600, 1323511200, 1323514800, 1323518400, 1323522000, 1323525600, 
    1323529200, 1323532800, 1323536400, 1323540000, 1323543600, 1323547200, 
    1323550800, 1323554400, 1323558000, 1323561600, 1323565200, 1323568800, 
    1323572400, 1323576000, 1323579600, 1323583200, 1323586800, 1323590400, 
    1323594000, 1323597600, 1323601200, 1323604800, 1323608400, 1323612000, 
    1323615600, 1323619200, 1323622800, 1323626400, 1323630000, 1323633600, 
    1323637200, 1323640800, 1323644400, 1323648000, 1323651600, 1323655200, 
    1323658800, 1323662400, 1323666000, 1323669600, 1323673200, 1323676800, 
    1323680400, 1323687600, 1323691200, 1323694800, 1323698400, 1323702000, 
    1323705600, 1323709200, 1323712800, 1323716400, 1323720000, 1323723600, 
    1323727200, 1323730800, 1323734400, 1323738000, 1323741600, 1323745200, 
    1323748800, 1323752400, 1323756000, 1323759600, 1323763200, 1323766800, 
    1323770400, 1323774000, 1323777600, 1323781200, 1323784800, 1323788400, 
    1323792000, 1323795600, 1323799200, 1323802800, 1323806400, 1323810000, 
    1323813600, 1323817200, 1323820800, 1323824400, 1323828000, 1323831600, 
    1323835200, 1323838800, 1323842400, 1323846000, 1323849600, 1323853200, 
    1323856800, 1323860400, 1323864000, 1323867600, 1323871200, 1323874800, 
    1323878400, 1323882000, 1323885600, 1323889200, 1323892800, 1323896400, 
    1323900000, 1323903600, 1323907200, 1323910800, 1323914400, 1323918000, 
    1323921600, 1323925200, 1323928800, 1323932400, 1323936000, 1323939600, 
    1323943200, 1323946800, 1323950400, 1323954000, 1323957600, 1323961200, 
    1323964800, 1323968400, 1324303200, 1324306800, 1324310400, 1324314000, 
    1324404000, 1324407600, 1324411200, 1324414800, 1324418400, 1324422000, 
    1324425600, 1324429200, 1324432800, 1324436400, 1324440000, 1324443600, 
    1324447200, 1324450800, 1324454400, 1324458000, 1324461600, 1324465200, 
    1324468800, 1324472400, 1324476000, 1324479600, 1324483200, 1324486800, 
    1324490400, 1324494000, 1324497600, 1324501200, 1324504800, 1324508400, 
    1324512000, 1324515600, 1324519200, 1324522800, 1324526400, 1324530000, 
    1324533600, 1324537200, 1324540800, 1324544400, 1324548000, 1324551600, 
    1324555200, 1324558800, 1324562400, 1324566000, 1324569600, 1324573200, 
    1324576800, 1324580400, 1324584000, 1324587600, 1324591200, 1324594800, 
    1324598400, 1324602000, 1324605600, 1324609200, 1324612800, 1324616400, 
    1324620000, 1324623600, 1324627200, 1324630800, 1324634400, 1324638000, 
    1324641600, 1324645200, 1324648800, 1324652400, 1324656000, 1324659600, 
    1324663200, 1324666800, 1324670400, 1324674000, 1324677600, 1324681200, 
    1324684800, 1324688400, 1324692000, 1324695600, 1324699200, 1324702800, 
    1324706400, 1324710000, 1324713600, 1324717200, 1324720800, 1324724400, 
    1324728000, 1324731600, 1324735200, 1324738800, 1324742400, 1324746000, 
    1324749600, 1324753200, 1324756800, 1324760400, 1324764000, 1324767600, 
    1324771200, 1324774800, 1324778400, 1324782000, 1324785600, 1324789200, 
    1324792800, 1324796400, 1324800000, 1324803600, 1324807200, 1324810800, 
    1324814400, 1324818000, 1324821600, 1324825200, 1324828800, 1324832400, 
    1324836000, 1324839600, 1324843200, 1324846800, 1324850400, 1324854000, 
    1324857600, 1324861200, 1324864800, 1324868400, 1324872000, 1324875600, 
    1324879200, 1324882800, 1324886400, 1324890000, 1324893600, 1324897200, 
    1324900800, 1324904400, 1324908000, 1324911600, 1324915200, 1324918800, 
    1324922400, 1324926000, 1324929600, 1324933200, 1324936800, 1324940400, 
    1324944000, 1324947600, 1324951200, 1324954800, 1324958400, 1324962000, 
    1324965600, 1324969200, 1324972800, 1324976400, 1324980000, 1324983600, 
    1324987200, 1324990800, 1324994400, 1324998000, 1325001600, 1325005200, 
    1325008800, 1325012400, 1325016000, 1325019600, 1325023200, 1325026800, 
    1325030400, 1325034000, 1325037600, 1325041200, 1325044800, 1325048400, 
    1325052000, 1325055600, 1325059200, 1325062800, 1325066400, 1325070000, 
    1325073600, 1325077200, 1325080800, 1325084400, 1325088000, 1325091600, 
    1325095200, 1325098800, 1325102400, 1325106000, 1325109600, 1325113200, 
    1325116800, 1325120400, 1325124000, 1325127600, 1325131200, 1325134800, 
    1325138400, 1325142000, 1325145600, 1325149200, 1325152800, 1325156400, 
    1325160000, 1325163600, 1325167200, 1325170800, 1325174400, 1325178000, 
    1325181600, 1325185200, 1325188800, 1325192400, 1325196000, 1325199600, 
    1325203200, 1325206800, 1325210400, 1325214000, 1325217600, 1325221200, 
    1325224800, 1325228400, 1325232000, 1325235600, 1325239200, 1325242800, 
    1325246400, 1325250000, 1325253600, 1325257200, 1325260800, 1325264400, 
    1325268000, 1325271600, 1325275200, 1325278800, 1325282400, 1325286000, 
    1325289600, 1325293200, 1325296800, 1325300400, 1325304000, 1325307600, 
    1325311200, 1325314800, 1325318400, 1325322000, 1325325600, 1325329200, 
    1325332800, 1325336400, 1325340000, 1325343600, 1325347200, 1325350800, 
    1325354400, 1325358000, 1325361600, 1325365200, 1325368800, 1325372400, 
    1325376000, 1325379600, 1325383200, 1325386800, 1325390400, 1325394000, 
    1325397600, 1325401200, 1325404800, 1325408400, 1325412000, 1325415600, 
    1325419200, 1325422800, 1325426400, 1325430000, 1325433600, 1325437200, 
    1325440800, 1325444400, 1325448000, 1325451600, 1325455200, 1325458800, 
    1325462400, 1325466000, 1325469600, 1325473200, 1325476800, 1325480400, 
    1325484000, 1325487600, 1325491200, 1325494800, 1325502000, 1325505600, 
    1325509200, 1325512800, 1325516400, 1325520000, 1325523600, 1325527200, 
    1325530800, 1325534400, 1325538000, 1325541600, 1325545200, 1325548800, 
    1325552400, 1325556000, 1325559600, 1325563200, 1325566800, 1325570400, 
    1325574000, 1325577600, 1325581200, 1325584800, 1325588400, 1325592000, 
    1325595600, 1325599200, 1325602800, 1325606400, 1325610000, 1325613600, 
    1325617200, 1325620800, 1325624400, 1325628000, 1325631600, 1325635200, 
    1325638800, 1325642400, 1325646000, 1325649600, 1325653200, 1325656800, 
    1325660400, 1325664000, 1325667600, 1325671200, 1325674800, 1325678400, 
    1325682000, 1325685600, 1325689200, 1325692800, 1325696400, 1325700000, 
    1325703600, 1325707200, 1325710800, 1325714400, 1325718000, 1325721600, 
    1325725200, 1325728800, 1325732400, 1325736000, 1325739600, 1325743200, 
    1325746800, 1325750400, 1325754000, 1325757600, 1325761200, 1325764800, 
    1325768400, 1325772000, 1325775600, 1325779200, 1325782800, 1325786400, 
    1325790000, 1325793600, 1325797200, 1325800800, 1325804400, 1325808000, 
    1325811600, 1325815200, 1325818800, 1325822400, 1325826000, 1325829600, 
    1325833200, 1325836800, 1325840400, 1325844000, 1325847600, 1325851200, 
    1325854800, 1325858400, 1325862000, 1325865600, 1325869200, 1325872800, 
    1325876400, 1325880000, 1325883600, 1325887200, 1325890800, 1325894400, 
    1325898000, 1325901600, 1325905200, 1325908800, 1325912400, 1325916000, 
    1325919600, 1325923200, 1325926800, 1325930400, 1325934000, 1325937600, 
    1325941200, 1325944800, 1325948400, 1325952000, 1325955600, 1325959200, 
    1325962800, 1325966400, 1325970000, 1325973600, 1325977200, 1325980800, 
    1325984400, 1325988000, 1325991600, 1325995200, 1325998800, 1326002400, 
    1326006000, 1326009600, 1326013200, 1326016800, 1326020400, 1326024000, 
    1326027600, 1326031200, 1326034800, 1326038400, 1326042000, 1326045600, 
    1326049200, 1326052800, 1326056400, 1326060000, 1326063600, 1326067200, 
    1326070800, 1326074400, 1326078000, 1326081600, 1326085200, 1326088800, 
    1326092400, 1326096000, 1326099600, 1326103200, 1326106800, 1326110400, 
    1326114000, 1326117600, 1326121200, 1326124800, 1326128400, 1326132000, 
    1326135600, 1326139200, 1326142800, 1326146400, 1326150000, 1326189600, 
    1326193200, 1326196800, 1326200400, 1326204000, 1326207600, 1326211200, 
    1326214800, 1326456000, 1326459600, 1326463200, 1326466800, 1326470400, 
    1326474000, 1326477600, 1326481200, 1326484800, 1326488400, 1326492000, 
    1326495600, 1326499200, 1326502800, 1326506400, 1326510000, 1326513600, 
    1326517200, 1326520800, 1326524400, 1326528000, 1326531600, 1326535200, 
    1326538800, 1326542400, 1326546000, 1326549600, 1326553200, 1326556800, 
    1326560400, 1326564000, 1326567600, 1326571200, 1326574800, 1326578400, 
    1326582000, 1326585600, 1326589200, 1326592800, 1326596400, 1326600000, 
    1326603600, 1326607200, 1326610800, 1326614400, 1326618000, 1326621600, 
    1326625200, 1326628800, 1326632400, 1326636000, 1326639600, 1326643200, 
    1326646800, 1326650400, 1326654000, 1326657600, 1326661200, 1326664800, 
    1326668400, 1326672000, 1326675600, 1326679200, 1326682800, 1326686400, 
    1326690000, 1326693600, 1326697200, 1326700800, 1326704400, 1326708000, 
    1326711600, 1326715200, 1326718800, 1326722400, 1326726000, 1326729600, 
    1326733200, 1326736800, 1326740400, 1326744000, 1326747600, 1326751200, 
    1326754800, 1326758400, 1326762000, 1326765600, 1326769200, 1326772800, 
    1326776400, 1326780000, 1326783600, 1326787200, 1326790800, 1326794400, 
    1326798000, 1326801600, 1326805200, 1326808800, 1326812400, 1326816000, 
    1326819600, 1326823200, 1326826800, 1326830400, 1326834000, 1326837600, 
    1326841200, 1326844800, 1326848400, 1326852000, 1326855600, 1326859200, 
    1326862800, 1326866400, 1326870000, 1326873600, 1326877200, 1326880800, 
    1326884400, 1326888000, 1326891600, 1326895200, 1326898800, 1326902400, 
    1326906000, 1326909600, 1326913200, 1326916800, 1326920400, 1326924000, 
    1326927600, 1326931200, 1326934800, 1326938400, 1326942000, 1326945600, 
    1326949200, 1326952800, 1326956400, 1326960000, 1326963600, 1326967200, 
    1326970800, 1326974400, 1326978000, 1326981600, 1326985200, 1326988800, 
    1326992400, 1326996000, 1326999600, 1327003200, 1327006800, 1327010400, 
    1327014000, 1327017600, 1327021200, 1327024800, 1327028400, 1327032000, 
    1327035600, 1327039200, 1327042800, 1327046400, 1327050000, 1327053600, 
    1327057200, 1327060800, 1327064400, 1327068000, 1327071600, 1327075200, 
    1327078800, 1327082400, 1327086000, 1327089600, 1327093200, 1327096800, 
    1327100400, 1327104000, 1327107600, 1327111200, 1327114800, 1327118400, 
    1327122000, 1327125600, 1327129200, 1327132800, 1327136400, 1327140000, 
    1327143600, 1327147200, 1327150800, 1327154400, 1327158000, 1327161600, 
    1327165200, 1327168800, 1327172400, 1327176000, 1327179600, 1327183200, 
    1327186800, 1327190400, 1327194000, 1327197600, 1327201200, 1327204800, 
    1327208400, 1327212000, 1327215600, 1327219200, 1327222800, 1327226400, 
    1327230000, 1327233600, 1327237200, 1327240800, 1327244400, 1327248000, 
    1327251600, 1327255200, 1327258800, 1327262400, 1327266000, 1327269600, 
    1327273200, 1327276800, 1327280400, 1327284000, 1327287600, 1327291200, 
    1327294800, 1327298400, 1327302000, 1327305600, 1327309200, 1327312800, 
    1327316400, 1327320000, 1327323600, 1327327200, 1327330800, 1327334400, 
    1327338000, 1327341600, 1327345200, 1327348800, 1327352400, 1327356000, 
    1327359600, 1327363200, 1327366800, 1327370400, 1327374000, 1327377600, 
    1327381200, 1327384800, 1327388400, 1327392000, 1327395600, 1327399200, 
    1327402800, 1327406400, 1327410000, 1327413600, 1327417200, 1327420800, 
    1327424400, 1327428000, 1327431600, 1327435200, 1327438800, 1327442400, 
    1327446000, 1327449600, 1327453200, 1327456800, 1327460400, 1327464000, 
    1327467600, 1327471200, 1327474800, 1327478400, 1327482000, 1327485600, 
    1327489200, 1327492800, 1327496400, 1327500000, 1327503600, 1327507200, 
    1327510800, 1327514400, 1327518000, 1327521600, 1327525200, 1327528800, 
    1327532400, 1327536000, 1327539600, 1327543200, 1327546800, 1327550400, 
    1327554000, 1327557600, 1327561200, 1327564800, 1327568400, 1327572000, 
    1327575600, 1327579200, 1327582800, 1327586400, 1327590000, 1327593600, 
    1327597200, 1327600800, 1327604400, 1327608000, 1327611600, 1327615200, 
    1327618800, 1327622400, 1327626000, 1327629600, 1327633200, 1327636800, 
    1327640400, 1327644000, 1327647600, 1327651200, 1327654800, 1327658400, 
    1327662000, 1327665600, 1327669200, 1327672800, 1327676400, 1327680000, 
    1327683600, 1327687200, 1327690800, 1327694400, 1327698000, 1327701600, 
    1327705200, 1327708800, 1327712400, 1327716000, 1327719600, 1327723200, 
    1327726800, 1327730400, 1327734000, 1327737600, 1327741200, 1327744800, 
    1327748400, 1327752000, 1327755600, 1327759200, 1327762800, 1327766400, 
    1327770000, 1327773600, 1327777200, 1327780800, 1327784400, 1327788000, 
    1327791600, 1327795200, 1327798800, 1327802400, 1327806000, 1327809600, 
    1327813200, 1327816800, 1327820400, 1327824000, 1327827600, 1327831200, 
    1327834800, 1327838400, 1327842000, 1327845600, 1327849200, 1327852800, 
    1327856400, 1327860000, 1327863600, 1327867200, 1327870800, 1327874400, 
    1327878000, 1327881600, 1327885200, 1327888800, 1327892400, 1327896000, 
    1327899600, 1327903200, 1327906800, 1327910400, 1327914000, 1327917600, 
    1327921200, 1327924800, 1327928400, 1327932000, 1327935600, 1327939200, 
    1327942800, 1327946400, 1327950000, 1327953600, 1327957200, 1327960800, 
    1327964400, 1327968000, 1327971600, 1327975200, 1327978800, 1327982400, 
    1327986000, 1327989600, 1327993200, 1327996800, 1328000400, 1328004000, 
    1328007600, 1328011200, 1328014800, 1328018400, 1328022000, 1328025600, 
    1328029200, 1328032800, 1328036400, 1328040000, 1328043600, 1328047200, 
    1328050800, 1328054400, 1328058000, 1328061600, 1328065200, 1328068800, 
    1328072400, 1328076000, 1328079600, 1328083200, 1328086800, 1328090400, 
    1328094000, 1328097600, 1328101200, 1328104800, 1328108400, 1328112000, 
    1328115600, 1328119200, 1328122800, 1328126400, 1328130000, 1328133600, 
    1328137200, 1328140800, 1328144400, 1328148000, 1328151600, 1328155200, 
    1328158800, 1328162400, 1328166000, 1328169600, 1328173200, 1328176800, 
    1328180400, 1328184000, 1328187600, 1328191200, 1328194800, 1328198400, 
    1328202000, 1328205600, 1328209200, 1328212800, 1328216400, 1328220000, 
    1328223600, 1328227200, 1328230800, 1328234400, 1328238000, 1328241600, 
    1328245200, 1328248800, 1328252400, 1328256000, 1328259600, 1328266800, 
    1328270400, 1328274000, 1328277600, 1328281200, 1328284800, 1328288400, 
    1328292000, 1328295600, 1328299200, 1328302800, 1328306400, 1328310000, 
    1328313600, 1328317200, 1328320800, 1328324400, 1328328000, 1328331600, 
    1328335200, 1328338800, 1328342400, 1328346000, 1328349600, 1328353200, 
    1328356800, 1328360400, 1328364000, 1328367600, 1328371200, 1328374800, 
    1328378400, 1328382000, 1328385600, 1328389200, 1328392800, 1328396400, 
    1328400000, 1328403600, 1328407200, 1328410800, 1328414400, 1328418000, 
    1328421600, 1328425200, 1328428800, 1328432400, 1328436000, 1328439600, 
    1328443200, 1328446800, 1328450400, 1328454000, 1328457600, 1328461200, 
    1328464800, 1328468400, 1328472000, 1328475600, 1328479200, 1328482800, 
    1328486400, 1328490000, 1328493600, 1328497200, 1328500800, 1328504400, 
    1328508000, 1328511600, 1328515200, 1328518800, 1328522400, 1328526000, 
    1328529600, 1328533200, 1328536800, 1328540400, 1328544000, 1328547600, 
    1328551200, 1328554800, 1328558400, 1328562000, 1328565600, 1328569200, 
    1328572800, 1328576400, 1328580000, 1328583600, 1328587200, 1328590800, 
    1328594400, 1328598000, 1328601600, 1328605200, 1328608800, 1328612400, 
    1328616000, 1328619600, 1328623200, 1328626800, 1328630400, 1328634000, 
    1328637600, 1328641200, 1328644800, 1328648400, 1328652000, 1328655600, 
    1328659200, 1328662800, 1328666400, 1328670000, 1328673600, 1328677200, 
    1328680800, 1328684400, 1328688000, 1328691600, 1328695200, 1328698800, 
    1328702400, 1328706000, 1328709600, 1328713200, 1328716800, 1328720400, 
    1328724000, 1328727600, 1328731200, 1328734800, 1328738400, 1328742000, 
    1328745600, 1328749200, 1328752800, 1328756400, 1328760000, 1328763600, 
    1328767200, 1328770800, 1328774400, 1328778000, 1328781600, 1328788800, 
    1328792400, 1328796000, 1328799600, 1328803200, 1328806800, 1328810400, 
    1328814000, 1328817600, 1328821200, 1328824800, 1328828400, 1328832000, 
    1328835600, 1328839200, 1328842800, 1328846400, 1328850000, 1328853600, 
    1328857200, 1328860800, 1328864400, 1328868000, 1328871600, 1328875200, 
    1328878800, 1328882400, 1328886000, 1328889600, 1328893200, 1328896800, 
    1328900400, 1328904000, 1328907600, 1328911200, 1328914800, 1328918400, 
    1328922000, 1328925600, 1328929200, 1328932800, 1328936400, 1328940000, 
    1328943600, 1328947200, 1328950800, 1328954400, 1328958000, 1328961600, 
    1328965200, 1328968800, 1328972400, 1328976000, 1328979600, 1328983200, 
    1328986800, 1328990400, 1328994000, 1328997600, 1329001200, 1329004800, 
    1329008400, 1329012000, 1329015600, 1329019200, 1329022800, 1329026400, 
    1329030000, 1329033600, 1329037200, 1329040800, 1329044400, 1329048000, 
    1329051600, 1329055200, 1329058800, 1329062400, 1329066000, 1329069600, 
    1329073200, 1329076800, 1329080400, 1329084000, 1329087600, 1329091200, 
    1329094800, 1329098400, 1329102000, 1329105600, 1329109200, 1329112800, 
    1329116400, 1329120000, 1329123600, 1329127200, 1329130800, 1329134400, 
    1329138000, 1329141600, 1329145200, 1329148800, 1329152400, 1329156000, 
    1329159600, 1329163200, 1329166800, 1329170400, 1329174000, 1329177600, 
    1329181200, 1329184800, 1329188400, 1329192000, 1329195600, 1329199200, 
    1329202800, 1329206400, 1329210000, 1329213600, 1329217200, 1329220800, 
    1329224400, 1329228000, 1329231600, 1329235200, 1329238800, 1329242400, 
    1329246000, 1329249600, 1329253200, 1329256800, 1329260400, 1329264000, 
    1329267600, 1329271200, 1329274800, 1329278400, 1329282000, 1329285600, 
    1329289200, 1329292800, 1329296400, 1329300000, 1329303600, 1329307200, 
    1329310800, 1329314400, 1329318000, 1329321600, 1329325200, 1329328800, 
    1329332400, 1329336000, 1329339600, 1329343200, 1329346800, 1329350400, 
    1329354000, 1329357600, 1329361200, 1329364800, 1329368400, 1329372000, 
    1329375600, 1329379200, 1329382800, 1329386400, 1329390000, 1329393600, 
    1329397200, 1329400800, 1329404400, 1329408000, 1329411600, 1329415200, 
    1329418800, 1329422400, 1329426000, 1329429600, 1329433200, 1329436800, 
    1329440400, 1329444000, 1329447600, 1329451200, 1329454800, 1329458400, 
    1329462000, 1329465600, 1329469200, 1329472800, 1329476400, 1329480000, 
    1329483600, 1329487200, 1329490800, 1329494400, 1329498000, 1329501600, 
    1329505200, 1329508800, 1329512400, 1329516000, 1329519600, 1329523200, 
    1329526800, 1329530400, 1329534000, 1329537600, 1329541200, 1329544800, 
    1329548400, 1329552000, 1329555600, 1329559200, 1329562800, 1329566400, 
    1329570000, 1329573600, 1329577200, 1329580800, 1329584400, 1329588000, 
    1329591600, 1329595200, 1329598800, 1329602400, 1329606000, 1329609600, 
    1329613200, 1329616800, 1329620400, 1329624000, 1329627600, 1329631200, 
    1329634800, 1329638400, 1329642000, 1329645600, 1329649200, 1329652800, 
    1329656400, 1329660000, 1329663600, 1329667200, 1329670800, 1329674400, 
    1329678000, 1329681600, 1329685200, 1329688800, 1329692400, 1329696000, 
    1329699600, 1329703200, 1329706800, 1329710400, 1329714000, 1329717600, 
    1329721200, 1329724800, 1329728400, 1329732000, 1329735600, 1329739200, 
    1329742800, 1329746400, 1329750000, 1329753600, 1329757200, 1329760800, 
    1329764400, 1329768000, 1329771600, 1329775200, 1329778800, 1329782400, 
    1329786000, 1329789600, 1329793200, 1329796800, 1329800400, 1329804000, 
    1329807600, 1329811200, 1329814800, 1329818400, 1329822000, 1329825600, 
    1329829200, 1329832800, 1329836400, 1329840000, 1329843600, 1329847200, 
    1329850800, 1329854400, 1329858000, 1329861600, 1329865200, 1329868800, 
    1329872400, 1329876000, 1329879600, 1329883200, 1329886800, 1329890400, 
    1329894000, 1329897600, 1329901200, 1329904800, 1329908400, 1329912000, 
    1329915600, 1329919200, 1329922800, 1329926400, 1329930000, 1329933600, 
    1329937200, 1329940800, 1329944400, 1329948000, 1329951600, 1329955200, 
    1329958800, 1329962400, 1329966000, 1329969600, 1329973200, 1329976800, 
    1329980400, 1329984000, 1329987600, 1329991200, 1329994800, 1329998400, 
    1330002000, 1330005600, 1330009200, 1330012800, 1330016400, 1330020000, 
    1330023600, 1330027200, 1330030800, 1330034400, 1330038000, 1330084800, 
    1330088400, 1330092000, 1330095600, 1330099200, 1330102800, 1330106400, 
    1330110000, 1330113600, 1330117200, 1330120800, 1330124400, 1330128000, 
    1330131600, 1330135200, 1330138800, 1330142400, 1330146000, 1330149600, 
    1330153200, 1330156800, 1330160400, 1330164000, 1330167600, 1330171200, 
    1330174800, 1330178400, 1330182000, 1330185600, 1330189200, 1330192800, 
    1330196400, 1330200000, 1330203600, 1330207200, 1330210800, 1330214400, 
    1330218000, 1330221600, 1330225200, 1330228800, 1330232400, 1330236000, 
    1330239600, 1330243200, 1330246800, 1330250400, 1330254000, 1330257600, 
    1330261200, 1330264800, 1330268400, 1330272000, 1330275600, 1330279200, 
    1330282800, 1330286400, 1330290000, 1330293600, 1330297200, 1330300800, 
    1330304400, 1330308000, 1330311600, 1330315200, 1330318800, 1330322400, 
    1330326000, 1330329600, 1330333200, 1330336800, 1330340400, 1330344000, 
    1330347600, 1330351200, 1330354800, 1330358400, 1330362000, 1330365600, 
    1330369200, 1330372800, 1330376400, 1330380000, 1330383600, 1330387200, 
    1330390800, 1330394400, 1330398000, 1330401600, 1330405200, 1330408800, 
    1330412400, 1330416000, 1330419600, 1330423200, 1330426800, 1330430400, 
    1330434000, 1330437600, 1330441200, 1330444800, 1330448400, 1330452000, 
    1330455600, 1330459200, 1330462800, 1330466400, 1330470000, 1330473600, 
    1330477200, 1330480800, 1330484400, 1330488000, 1330491600, 1330495200, 
    1330498800, 1330502400, 1330506000, 1330509600, 1330513200, 1330516800, 
    1330520400, 1330524000, 1330527600, 1330531200, 1330534800, 1330538400, 
    1330542000, 1330545600, 1330549200, 1330552800, 1330556400, 1330560000, 
    1330563600, 1330567200, 1330570800, 1330574400, 1330578000, 1330581600, 
    1330585200, 1330588800, 1330592400, 1330596000, 1330599600, 1330603200, 
    1330606800, 1330610400, 1330614000, 1330617600, 1330621200, 1330624800, 
    1330628400, 1330632000, 1330635600, 1330639200, 1330642800, 1330646400, 
    1330650000, 1330653600, 1330657200, 1330660800, 1330664400, 1330668000, 
    1330671600, 1330675200, 1330678800, 1330682400, 1330686000, 1330689600, 
    1330693200, 1330696800, 1330700400, 1330704000, 1330707600, 1330711200, 
    1330714800, 1330718400, 1330722000, 1330725600, 1330729200, 1330732800, 
    1330736400, 1330740000, 1330743600, 1330747200, 1330750800, 1330754400, 
    1330758000, 1330761600, 1330765200, 1330768800, 1330772400, 1330776000, 
    1330779600, 1330783200, 1330786800, 1330790400, 1330794000, 1330797600, 
    1330801200, 1330804800, 1330808400, 1330812000, 1330815600, 1330819200, 
    1330822800, 1330826400, 1330830000, 1330833600, 1330837200, 1330840800, 
    1330844400, 1330848000, 1330851600, 1330855200, 1330858800, 1330862400, 
    1330866000, 1330869600, 1330873200, 1330876800, 1330880400, 1330884000, 
    1330887600, 1330891200, 1330894800, 1330898400, 1330902000, 1330905600, 
    1330909200, 1330912800, 1330916400, 1330920000, 1330923600, 1330927200, 
    1330930800, 1330934400, 1330938000, 1330941600, 1330945200, 1330948800, 
    1330952400, 1330956000, 1330959600, 1330963200, 1330966800, 1330970400, 
    1330974000, 1330977600, 1330981200, 1330984800, 1330988400, 1330992000, 
    1330995600, 1330999200, 1331002800, 1331006400, 1331010000, 1331013600, 
    1331017200, 1331020800, 1331024400, 1331028000, 1331031600, 1331035200, 
    1331038800, 1331042400, 1331046000, 1331049600, 1331053200, 1331056800, 
    1331060400, 1331064000, 1331067600, 1331071200, 1331074800, 1331078400, 
    1331082000, 1331085600, 1331089200, 1331092800, 1331096400, 1331100000, 
    1331103600, 1331107200, 1331110800, 1331114400, 1331118000, 1331121600, 
    1331125200, 1331128800, 1331132400, 1331136000, 1331139600, 1331143200, 
    1331146800, 1331150400, 1331154000, 1331157600, 1331161200, 1331164800, 
    1331168400, 1331172000, 1331175600, 1331179200, 1331182800, 1331186400, 
    1331190000, 1331193600, 1331197200, 1331200800, 1331204400, 1331208000, 
    1331211600, 1331215200, 1331218800, 1331222400, 1331226000, 1331229600, 
    1331233200, 1331236800, 1331240400, 1331244000, 1331247600, 1331251200, 
    1331254800, 1331258400, 1331262000, 1331265600, 1331269200, 1331272800, 
    1331276400, 1331280000, 1331283600, 1331287200, 1331290800, 1331294400, 
    1331298000, 1331301600, 1331305200, 1331308800, 1331312400, 1331316000, 
    1331319600, 1331323200, 1331326800, 1331330400, 1331334000, 1331337600, 
    1331341200, 1331344800, 1331348400, 1331352000, 1331355600, 1331359200, 
    1331362800, 1331366400, 1331370000, 1331373600, 1331377200, 1331380800, 
    1331384400, 1331388000, 1331391600, 1331395200, 1331398800, 1331402400, 
    1331406000, 1331409600, 1331413200, 1331416800, 1331420400, 1331424000, 
    1331427600, 1331431200, 1331434800, 1331438400, 1331442000, 1331445600, 
    1331449200, 1331452800, 1331456400, 1331460000, 1331463600, 1331467200, 
    1331470800, 1331474400, 1331478000, 1331481600, 1331485200, 1331488800, 
    1331492400, 1331496000, 1331499600, 1331503200, 1331506800, 1331510400, 
    1331514000, 1331517600, 1331521200, 1331524800, 1331528400, 1331532000, 
    1331535600, 1331539200, 1331542800, 1331546400, 1331550000, 1331553600, 
    1331557200, 1331560800, 1331564400, 1331568000, 1331571600, 1331575200, 
    1331578800, 1331582400, 1331586000, 1331589600, 1331593200, 1331596800, 
    1331600400, 1331604000, 1331607600, 1331611200, 1331614800, 1331618400, 
    1331622000, 1331625600, 1331629200, 1331632800, 1331636400, 1331640000, 
    1331643600, 1331647200, 1331650800, 1331654400, 1331658000, 1331661600, 
    1331665200, 1331668800, 1331672400, 1331676000, 1331679600, 1331683200, 
    1331686800, 1331690400, 1331694000, 1331697600, 1331701200, 1331704800, 
    1331708400, 1331712000, 1331715600, 1331719200, 1331722800, 1331726400, 
    1331730000, 1331733600, 1331737200, 1331740800, 1331744400, 1331748000, 
    1331751600, 1331755200, 1331758800, 1331762400, 1331766000, 1331769600, 
    1331773200, 1331776800, 1331780400, 1331784000, 1331787600, 1331791200, 
    1331794800, 1331798400, 1331802000, 1331805600, 1331809200, 1331812800, 
    1331816400, 1331820000, 1331823600, 1331827200, 1331830800, 1331834400, 
    1331838000, 1331841600, 1331845200, 1331848800, 1331852400, 1331856000, 
    1331859600, 1331863200, 1331866800, 1331870400, 1331874000, 1331877600, 
    1331881200, 1331884800, 1331888400, 1331892000, 1331895600, 1331899200, 
    1331902800, 1331906400, 1331910000, 1331913600, 1331917200, 1331920800, 
    1331924400, 1331928000, 1331931600, 1331935200, 1331938800, 1331942400, 
    1331946000, 1331949600, 1331953200, 1331956800, 1331960400, 1331964000, 
    1331967600, 1331971200, 1331974800, 1331978400, 1331982000, 1331985600, 
    1331989200, 1331992800, 1331996400, 1332000000, 1332003600, 1332007200, 
    1332010800, 1332014400, 1332018000, 1332021600, 1332025200, 1332028800, 
    1332032400, 1332036000, 1332039600, 1332043200, 1332046800, 1332050400, 
    1332054000, 1332057600, 1332061200, 1332064800, 1332068400, 1332072000, 
    1332075600, 1332079200, 1332082800, 1332086400, 1332090000, 1332093600, 
    1332097200, 1332100800, 1332104400, 1332108000, 1332111600, 1332115200, 
    1332118800, 1332122400, 1332126000, 1332129600, 1332133200, 1332136800, 
    1332140400, 1332144000, 1332147600, 1332151200, 1332154800, 1332158400, 
    1332162000, 1332165600, 1332169200, 1332172800, 1332176400, 1332180000, 
    1332183600, 1332187200, 1332190800, 1332194400, 1332198000, 1332201600, 
    1332205200, 1332208800, 1332212400, 1332216000, 1332219600, 1332223200, 
    1332226800, 1332230400, 1332234000, 1332237600, 1332241200, 1332244800, 
    1332248400, 1332252000, 1332255600, 1332259200, 1332262800, 1332266400, 
    1332270000, 1332273600, 1332277200, 1332280800, 1332284400, 1332288000, 
    1332291600, 1332295200, 1332298800, 1332302400, 1332306000, 1332309600, 
    1332313200, 1332316800, 1332320400, 1332324000, 1332327600, 1332331200, 
    1332334800, 1332338400, 1332342000, 1332345600, 1332349200, 1332352800, 
    1332356400, 1332360000, 1332363600, 1332367200, 1332370800, 1332374400, 
    1332378000, 1332381600, 1332385200, 1332388800, 1332392400, 1332396000, 
    1332399600, 1332403200, 1332406800, 1332410400, 1332414000, 1332417600, 
    1332421200, 1332424800, 1332428400, 1332432000, 1332435600, 1332439200, 
    1332442800, 1332446400, 1332450000, 1332453600, 1332457200, 1332460800, 
    1332464400, 1332468000, 1332471600, 1332475200, 1332478800, 1332482400, 
    1332486000, 1332489600, 1332493200, 1332496800, 1332500400, 1332504000, 
    1332507600, 1332511200, 1332514800, 1332518400, 1332522000, 1332525600, 
    1332529200, 1332532800, 1332536400, 1332540000, 1332543600, 1332547200, 
    1332550800, 1332554400, 1332558000, 1332561600, 1332565200, 1332568800, 
    1332572400, 1332576000, 1332579600, 1332583200, 1332586800, 1332590400, 
    1332594000, 1332597600, 1332601200, 1332604800, 1332608400, 1332612000, 
    1332615600, 1332619200, 1332622800, 1332626400, 1332630000, 1332633600, 
    1332637200, 1332640800, 1332644400, 1332648000, 1332651600, 1332655200, 
    1332658800, 1332662400, 1332666000, 1332669600, 1332673200, 1332676800, 
    1332680400, 1332684000, 1332687600, 1332691200, 1332694800, 1332698400, 
    1332702000, 1332705600, 1332709200, 1332712800, 1332716400, 1332720000, 
    1332723600, 1332727200, 1332730800, 1332734400, 1332738000, 1332741600, 
    1332745200, 1332748800, 1332752400, 1332756000, 1332759600, 1332763200, 
    1332766800, 1332770400, 1332774000, 1332777600, 1332781200, 1332784800, 
    1332788400, 1332792000, 1332795600, 1332799200, 1332802800, 1332806400, 
    1332810000, 1332813600, 1332817200, 1332820800, 1332824400, 1332828000, 
    1332831600, 1332835200, 1332838800, 1332842400, 1332846000, 1332849600, 
    1332853200, 1332856800, 1332860400, 1332864000, 1332867600, 1332871200, 
    1332874800, 1332878400, 1332882000, 1332885600, 1332889200, 1332892800, 
    1332896400, 1332900000, 1332903600, 1332907200, 1332910800, 1332914400, 
    1332918000, 1332921600, 1332925200, 1332928800, 1332932400, 1332936000, 
    1332939600, 1332943200, 1332946800, 1332950400, 1332954000, 1332957600, 
    1332961200, 1332964800, 1332968400, 1332972000, 1332975600, 1332979200, 
    1332982800, 1332986400, 1332990000, 1332993600, 1332997200, 1333000800, 
    1333004400, 1333008000, 1333011600, 1333015200, 1333018800, 1333022400, 
    1333026000, 1333029600, 1333033200, 1333036800, 1333040400, 1333044000, 
    1333047600, 1333051200, 1333054800, 1333058400, 1333062000, 1333065600, 
    1333069200, 1333072800, 1333076400, 1333080000, 1333083600, 1333087200, 
    1333090800, 1333094400, 1333098000, 1333101600, 1333105200, 1333108800, 
    1333112400, 1333116000, 1333119600, 1333123200, 1333126800, 1333130400, 
    1333134000, 1333137600, 1333141200, 1333144800, 1333148400, 1333152000, 
    1333155600, 1333159200, 1333162800, 1333166400, 1333170000, 1333173600, 
    1333177200, 1333180800, 1333184400, 1333188000, 1333191600, 1333195200, 
    1333198800, 1333202400, 1333206000, 1333209600, 1333213200, 1333216800, 
    1333220400, 1333224000, 1333227600, 1333231200, 1333234800, 1333238400, 
    1333242000, 1333245600, 1333249200, 1333252800, 1333256400, 1333260000, 
    1333263600, 1333267200, 1333270800, 1333274400, 1333278000, 1333281600, 
    1333285200, 1333288800, 1333292400, 1333296000, 1333299600, 1333303200, 
    1333306800, 1333310400, 1333314000, 1333317600, 1333321200, 1333324800, 
    1333328400, 1333332000, 1333335600, 1333339200, 1333342800, 1333346400, 
    1333350000, 1333353600, 1333357200, 1333360800, 1333364400, 1333368000, 
    1333371600, 1333375200, 1333378800, 1333382400, 1333386000, 1333389600, 
    1333393200, 1333396800, 1333400400, 1333404000, 1333407600, 1333411200, 
    1333414800, 1333418400, 1333422000, 1333425600, 1333429200, 1333432800, 
    1333436400, 1333440000, 1333443600, 1333447200, 1333450800, 1333454400, 
    1333458000, 1333461600, 1333465200, 1333468800, 1333472400, 1333476000, 
    1333479600, 1333483200, 1333486800, 1333490400, 1333494000, 1333497600, 
    1333501200, 1333504800, 1333508400, 1333512000, 1333515600, 1333519200, 
    1333522800, 1333526400, 1333530000, 1333533600, 1333537200, 1333540800, 
    1333544400, 1333548000, 1333551600, 1333555200, 1333558800, 1333562400, 
    1333566000, 1333569600, 1333573200, 1333576800, 1333580400, 1333584000, 
    1333587600, 1333591200, 1333594800, 1333598400, 1333602000, 1333605600, 
    1333609200, 1333612800, 1333616400, 1333620000, 1333623600, 1333627200, 
    1333630800, 1333634400, 1333638000, 1333641600, 1333645200, 1333648800, 
    1333652400, 1333656000, 1333659600, 1333663200, 1333666800, 1333670400, 
    1333674000, 1333677600, 1333681200, 1333684800, 1333688400, 1333692000, 
    1333695600, 1333699200, 1333702800, 1333706400, 1333710000, 1333713600, 
    1333717200, 1333720800, 1333724400, 1333728000, 1333731600, 1333735200, 
    1333738800, 1333742400, 1333746000, 1333749600, 1333753200, 1333756800, 
    1333760400, 1333764000, 1333767600, 1333771200, 1333774800, 1333778400, 
    1333782000, 1333785600, 1333789200, 1333792800, 1333796400, 1333800000, 
    1333803600, 1333807200, 1333810800, 1333814400, 1333818000, 1333821600, 
    1333825200, 1333828800, 1333832400, 1333836000, 1333839600, 1333843200, 
    1333846800, 1333850400, 1333854000, 1333857600, 1333861200, 1333864800, 
    1333868400, 1333872000, 1333875600, 1333879200, 1333882800, 1333886400, 
    1333890000, 1333893600, 1333897200, 1333900800, 1333904400, 1333908000, 
    1333911600, 1333915200, 1333918800, 1333922400, 1333926000, 1333929600, 
    1333933200, 1333936800, 1333940400, 1333944000, 1333947600, 1333951200, 
    1333954800, 1333958400, 1333962000, 1333965600, 1333969200, 1333972800, 
    1333976400, 1333980000, 1333983600, 1333987200, 1333990800, 1333994400, 
    1333998000, 1334001600, 1334005200, 1334008800, 1334012400, 1334016000, 
    1334019600, 1334023200, 1334026800, 1334030400, 1334034000, 1334037600, 
    1334041200, 1334044800, 1334048400, 1334052000, 1334055600, 1334059200, 
    1334062800, 1334066400, 1334070000, 1334073600, 1334077200, 1334080800, 
    1334084400, 1334088000, 1334091600, 1334095200, 1334098800, 1334102400, 
    1334106000, 1334109600, 1334113200, 1334116800, 1334120400, 1334124000, 
    1334127600, 1334131200, 1334134800, 1334138400, 1334142000, 1334145600, 
    1334149200, 1334152800, 1334156400, 1334160000, 1334163600, 1334167200, 
    1334170800, 1334174400, 1334178000, 1334181600, 1334185200, 1334188800, 
    1334192400, 1334196000, 1334199600, 1334203200, 1334206800, 1334210400, 
    1334214000, 1334217600, 1334221200, 1334224800, 1334228400, 1334232000, 
    1334235600, 1334239200, 1334242800, 1334246400, 1334250000, 1334253600, 
    1334257200, 1334260800, 1334264400, 1334268000, 1334271600, 1334275200, 
    1334278800, 1334282400, 1334286000, 1334289600, 1334293200, 1334296800, 
    1334300400, 1334304000, 1334307600, 1334311200, 1334314800, 1334318400, 
    1334322000, 1334325600, 1334329200, 1334332800, 1334336400, 1334340000, 
    1334343600, 1334347200, 1334350800, 1334354400, 1334358000, 1334361600, 
    1334365200, 1334368800, 1334372400, 1334376000, 1334379600, 1334383200, 
    1334386800, 1334390400, 1334394000, 1334397600, 1334401200, 1334404800, 
    1334408400, 1334412000, 1334415600, 1334419200, 1334422800, 1334426400, 
    1334430000, 1334433600, 1334437200, 1334440800, 1334444400, 1334448000, 
    1334451600, 1334455200, 1334458800, 1334462400, 1334466000, 1334469600, 
    1334473200, 1334476800, 1334480400, 1334484000, 1334487600, 1334491200, 
    1334494800, 1334498400, 1334502000, 1334505600, 1334509200, 1334512800, 
    1334516400, 1334520000, 1334523600, 1334527200, 1334530800, 1334534400, 
    1334538000, 1334541600, 1334545200, 1334548800, 1334552400, 1334556000, 
    1334559600, 1334563200, 1334566800, 1334570400, 1334574000, 1334577600, 
    1334581200, 1334584800, 1334588400, 1334592000, 1334595600, 1334599200, 
    1334602800, 1334606400, 1334610000, 1334613600, 1334617200, 1334620800, 
    1334624400, 1334628000, 1334631600, 1334635200, 1334638800, 1334642400, 
    1334646000, 1334649600, 1334653200, 1334656800, 1334660400, 1334664000, 
    1334667600, 1334671200, 1334674800, 1334678400, 1334682000, 1334685600, 
    1334689200, 1334692800, 1334696400, 1334700000, 1334703600, 1334707200, 
    1334710800, 1334714400, 1334718000, 1334721600, 1334725200, 1334728800, 
    1334732400, 1334736000, 1334739600, 1334743200, 1334746800, 1334750400, 
    1334754000, 1334757600, 1334761200, 1334764800, 1334768400, 1334772000, 
    1334775600, 1334779200, 1334782800, 1334786400, 1334790000, 1334793600, 
    1334797200, 1334800800, 1334804400, 1334808000, 1334811600, 1334815200, 
    1334818800, 1334822400, 1334826000, 1334829600, 1334833200, 1334836800, 
    1334840400, 1334844000, 1334847600, 1334851200, 1334854800, 1334858400, 
    1334862000, 1334865600, 1334869200, 1334872800, 1334876400, 1334880000, 
    1334883600, 1334887200, 1334890800, 1334894400, 1334898000, 1334901600, 
    1334905200, 1334908800, 1334912400, 1334916000, 1334919600, 1334923200, 
    1334926800, 1334930400, 1334934000, 1334937600, 1334941200, 1334944800, 
    1334948400, 1334952000, 1334955600, 1334959200, 1334962800, 1334966400, 
    1334970000, 1334973600, 1334977200, 1334980800, 1334984400, 1334988000, 
    1334991600, 1334995200, 1334998800, 1335002400, 1335006000, 1335009600, 
    1335013200, 1335016800, 1335020400, 1335024000, 1335027600, 1335031200, 
    1335034800, 1335038400, 1335042000, 1335045600, 1335049200, 1335052800, 
    1335056400, 1335060000, 1335063600, 1335067200, 1335070800, 1335074400, 
    1335078000, 1335081600, 1335085200, 1335088800, 1335092400, 1335096000, 
    1335099600, 1335103200, 1335106800, 1335110400, 1335114000, 1335117600, 
    1335121200, 1335124800, 1335128400, 1335132000, 1335135600, 1335139200, 
    1335142800, 1335146400, 1335150000, 1335153600, 1335157200, 1335160800, 
    1335164400, 1335168000, 1335171600, 1335175200, 1335178800, 1335182400, 
    1335186000, 1335189600, 1335193200, 1335196800, 1335200400, 1335204000, 
    1335207600, 1335211200, 1335214800, 1335218400, 1335222000, 1335225600, 
    1335229200, 1335232800, 1335236400, 1335240000, 1335243600, 1335247200, 
    1335250800, 1335254400, 1335258000, 1335261600, 1335265200, 1335268800, 
    1335272400, 1335276000, 1335279600, 1335283200, 1335286800, 1335290400, 
    1335294000, 1335297600, 1335301200, 1335304800, 1335308400, 1335312000, 
    1335315600, 1335319200, 1335322800, 1335326400, 1335330000, 1335333600, 
    1335337200, 1335340800, 1335344400, 1335348000, 1335351600, 1335355200, 
    1335358800, 1335362400, 1335366000, 1335369600, 1335373200, 1335376800, 
    1335380400, 1335384000, 1335387600, 1335391200, 1335394800, 1335398400, 
    1335402000, 1335405600, 1335409200, 1335412800, 1335416400, 1335420000, 
    1335423600, 1335427200, 1335430800, 1335434400, 1335438000, 1335441600, 
    1335445200, 1335448800, 1335452400, 1335456000, 1335459600, 1335463200, 
    1335466800, 1335470400, 1335474000, 1335477600, 1335481200, 1335484800, 
    1335488400, 1335492000, 1335495600, 1335499200, 1335502800, 1335506400, 
    1335510000, 1335513600, 1335517200, 1335520800, 1335524400, 1335528000, 
    1335531600, 1335535200, 1335538800, 1335542400, 1335546000, 1335549600, 
    1335553200, 1335556800, 1335560400, 1335564000, 1335567600, 1335571200, 
    1335574800, 1335578400, 1335582000, 1335585600, 1335589200, 1335592800, 
    1335596400, 1335600000, 1335603600, 1335607200, 1335610800, 1335614400, 
    1335618000, 1335621600, 1335625200, 1335628800, 1335632400, 1335636000, 
    1335639600, 1335643200, 1335646800, 1335650400, 1335654000, 1335657600, 
    1335661200, 1335664800, 1335668400, 1335672000, 1335675600, 1335679200, 
    1335682800, 1335686400, 1335690000, 1335693600, 1335697200, 1335700800, 
    1335704400, 1335708000, 1335711600, 1335715200, 1335718800, 1335722400, 
    1335726000, 1335729600, 1335733200, 1335736800, 1335740400, 1335744000, 
    1335747600, 1335751200, 1335754800, 1335758400, 1335762000, 1335765600, 
    1335769200, 1335772800, 1335776400, 1335780000, 1335783600, 1335787200, 
    1335790800, 1335794400, 1335798000, 1335801600, 1335805200, 1335808800, 
    1335812400, 1335816000, 1335819600, 1335823200, 1335826800, 1335830400, 
    1335834000, 1335837600, 1335841200, 1335844800, 1335848400, 1335852000, 
    1335855600, 1335859200, 1335862800, 1335866400, 1335870000, 1335873600, 
    1335877200, 1335880800, 1335884400, 1335888000, 1335891600, 1335895200, 
    1335898800, 1335902400, 1335906000, 1335909600, 1335913200, 1335916800, 
    1335920400, 1335924000, 1335927600, 1335931200, 1335934800, 1335938400, 
    1335942000, 1335945600, 1335949200, 1335952800, 1335956400, 1335960000, 
    1335963600, 1335967200, 1335970800, 1335974400, 1335978000, 1335981600, 
    1335985200, 1335988800, 1335992400, 1335996000, 1335999600, 1336003200, 
    1336006800, 1336010400, 1336014000, 1336017600, 1336021200, 1336024800, 
    1336028400, 1336032000, 1336035600, 1336039200, 1336042800, 1336046400, 
    1336050000, 1336053600, 1336057200, 1336060800, 1336064400, 1336068000, 
    1336071600, 1336075200, 1336078800, 1336082400, 1336086000, 1336089600, 
    1336093200, 1336096800, 1336100400, 1336104000, 1336107600, 1336111200, 
    1336114800, 1336118400, 1336122000, 1336125600, 1336129200, 1336132800, 
    1336136400, 1336140000, 1336143600, 1336147200, 1336150800, 1336154400, 
    1336158000, 1336161600, 1336165200, 1336168800, 1336172400, 1336176000, 
    1336179600, 1336183200, 1336186800, 1336190400, 1336194000, 1336197600, 
    1336201200, 1336204800, 1336208400, 1336212000, 1336215600, 1336219200, 
    1336222800, 1336226400, 1336230000, 1336233600, 1336237200, 1336240800, 
    1336244400, 1336248000, 1336251600, 1336255200, 1336258800, 1336262400, 
    1336266000, 1336269600, 1336273200, 1336276800, 1336280400, 1336284000, 
    1336287600, 1336291200, 1336294800, 1336298400, 1336302000, 1336305600, 
    1336309200, 1336312800, 1336316400, 1336320000, 1336323600, 1336327200, 
    1336330800, 1336334400, 1336338000, 1336341600, 1336345200, 1336348800, 
    1336352400, 1336356000, 1336359600, 1336363200, 1336366800, 1336370400, 
    1336374000, 1336377600, 1336381200, 1336384800, 1336388400, 1336392000, 
    1336395600, 1336399200, 1336402800, 1336406400, 1336410000, 1336413600, 
    1336417200, 1336420800, 1336424400, 1336428000, 1336431600, 1336435200, 
    1336438800, 1336442400, 1336446000, 1336449600, 1336453200, 1336456800, 
    1336460400, 1336464000, 1336467600, 1336471200, 1336474800, 1336478400, 
    1336482000, 1336485600, 1336489200, 1336492800, 1336496400, 1336500000, 
    1336503600, 1336507200, 1336510800, 1336514400, 1336518000, 1336521600, 
    1336525200, 1336528800, 1336532400, 1336536000, 1336539600, 1336543200, 
    1336546800, 1336550400, 1336554000, 1336557600, 1336561200, 1336564800, 
    1336568400, 1336572000, 1336575600, 1336579200, 1336582800, 1336586400, 
    1336590000, 1336593600, 1336597200, 1336600800, 1336604400, 1336608000, 
    1336611600, 1336615200, 1336618800, 1336622400, 1336626000, 1336629600, 
    1336633200, 1336636800, 1336640400, 1336644000, 1336647600, 1336651200, 
    1336654800, 1336658400, 1336662000, 1336665600, 1336669200, 1336672800, 
    1336676400, 1336680000, 1336683600, 1336687200, 1336690800, 1336694400, 
    1336698000, 1336701600, 1336705200, 1336708800, 1336712400, 1336716000, 
    1336719600, 1336723200, 1336726800, 1336730400, 1336734000, 1336737600, 
    1336741200, 1336744800, 1336748400, 1336752000, 1336755600, 1336759200, 
    1336762800, 1336766400, 1336770000, 1336773600, 1336777200, 1336780800, 
    1336784400, 1336788000, 1336791600, 1336795200, 1336798800, 1336802400, 
    1336806000, 1336809600, 1336813200, 1336816800, 1336820400, 1336824000, 
    1336827600, 1336831200, 1336834800, 1336838400, 1336842000, 1336845600, 
    1336849200, 1336852800, 1336856400, 1336860000, 1336863600, 1336867200, 
    1336870800, 1336874400, 1336878000, 1336881600, 1336885200, 1336888800, 
    1336892400, 1336896000, 1336899600, 1336903200, 1336906800, 1336910400, 
    1336914000, 1336917600, 1336921200, 1336924800, 1336928400, 1336932000, 
    1336935600, 1336939200, 1336942800, 1336946400, 1336950000, 1336953600, 
    1336957200, 1336960800, 1336964400, 1336968000, 1336971600, 1336975200, 
    1336978800, 1336982400, 1336986000, 1336989600, 1336993200, 1336996800, 
    1337000400, 1337004000, 1337007600, 1337011200, 1337014800, 1337018400, 
    1337022000, 1337025600, 1337029200, 1337032800, 1337036400, 1337040000, 
    1337043600, 1337047200, 1337050800, 1337054400, 1337058000, 1337061600, 
    1337065200, 1337068800, 1337072400, 1337076000, 1337079600, 1337083200, 
    1337086800, 1337090400, 1337094000, 1337097600, 1337101200, 1337104800, 
    1337108400, 1337112000, 1337115600, 1337119200, 1337122800, 1337126400, 
    1337130000, 1337133600, 1337137200, 1337140800, 1337144400, 1337148000, 
    1337151600, 1337155200, 1337158800, 1337162400, 1337166000, 1337169600, 
    1337173200, 1337176800, 1337180400, 1337184000, 1337187600, 1337191200, 
    1337194800, 1337198400, 1337202000, 1337205600, 1337209200, 1337212800, 
    1337216400, 1337220000, 1337223600, 1337227200, 1337230800, 1337234400, 
    1337238000, 1337241600, 1337245200, 1337248800, 1337252400, 1337256000, 
    1337259600, 1337263200, 1337266800, 1337270400, 1337274000, 1337277600, 
    1337281200, 1337284800, 1337288400, 1337292000, 1337295600, 1337299200, 
    1337302800, 1337306400, 1337310000, 1337313600, 1337317200, 1337320800, 
    1337324400, 1337328000, 1337331600, 1337335200, 1337338800, 1337342400, 
    1337346000, 1337349600, 1337353200, 1337356800, 1337360400, 1337364000, 
    1337367600, 1337371200, 1337374800, 1337378400, 1337382000, 1337385600, 
    1337389200, 1337392800, 1337396400, 1337400000, 1337403600, 1337407200, 
    1337410800, 1337414400, 1337418000, 1337421600, 1337425200, 1337428800, 
    1337432400, 1337436000, 1337439600, 1337443200, 1337446800, 1337450400, 
    1337454000, 1337457600, 1337461200, 1337464800, 1337468400, 1337472000, 
    1337475600, 1337479200, 1337482800, 1337486400, 1337490000, 1337493600, 
    1337497200, 1337500800, 1337504400, 1337508000, 1337511600, 1337515200, 
    1337518800, 1337522400, 1337526000, 1337529600, 1337533200, 1337536800, 
    1337540400, 1337544000, 1337547600, 1337551200, 1337554800, 1337558400, 
    1337562000, 1337565600, 1337569200, 1337572800, 1337576400, 1337580000, 
    1337583600, 1337587200, 1337590800, 1337594400, 1337598000, 1337601600, 
    1337605200, 1337608800, 1337612400, 1337616000, 1337619600, 1337623200, 
    1337626800, 1337630400, 1337634000, 1337637600, 1337641200, 1337644800, 
    1337648400, 1337652000, 1337655600, 1337659200, 1337662800, 1337666400, 
    1337670000, 1337673600, 1337677200, 1337680800, 1337684400, 1337688000, 
    1337691600, 1337695200, 1337698800, 1337702400, 1337706000, 1337709600, 
    1337713200, 1337716800, 1337720400, 1337724000, 1337727600, 1337731200, 
    1337734800, 1337738400, 1337742000, 1337745600, 1337749200, 1337752800, 
    1337756400, 1337760000, 1337763600, 1337767200, 1337770800, 1337774400, 
    1337778000, 1337781600, 1337785200, 1337788800, 1337792400, 1337796000, 
    1337799600, 1337803200, 1337806800, 1337810400, 1337814000, 1337817600, 
    1337821200, 1337824800, 1337828400, 1337832000, 1337835600, 1337839200, 
    1337842800, 1337846400, 1337850000, 1337853600, 1337857200, 1337860800, 
    1337864400, 1337868000, 1337871600, 1337875200, 1337878800, 1337882400, 
    1337886000, 1337889600, 1337893200, 1337896800, 1337900400, 1337904000, 
    1337907600, 1337911200, 1337914800, 1337918400, 1337922000, 1337925600, 
    1337929200, 1337932800, 1337936400, 1337940000, 1337943600, 1337947200, 
    1337950800, 1337954400, 1337958000, 1337961600, 1337965200, 1337968800, 
    1337972400, 1337976000, 1337979600, 1337983200, 1337986800, 1337990400, 
    1337994000, 1337997600, 1338001200, 1338004800, 1338008400, 1338012000, 
    1338015600, 1338019200, 1338022800, 1338026400, 1338030000, 1338033600, 
    1338037200, 1338040800, 1338044400, 1338048000, 1338051600, 1338055200, 
    1338058800, 1338062400, 1338066000, 1338069600, 1338073200, 1338076800, 
    1338080400, 1338084000, 1338087600, 1338091200, 1338094800, 1338098400, 
    1338102000, 1338105600, 1338109200, 1338112800, 1338116400, 1338120000, 
    1338123600, 1338127200, 1338130800, 1338134400, 1338138000, 1338141600, 
    1338145200, 1338148800, 1338152400, 1338156000, 1338159600, 1338163200, 
    1338166800, 1338170400, 1338174000, 1338177600, 1338181200, 1338184800, 
    1338188400, 1338192000, 1338195600, 1338199200, 1338202800, 1338206400, 
    1338210000, 1338213600, 1338217200, 1338220800, 1338224400, 1338228000, 
    1338231600, 1338235200, 1338238800, 1338242400, 1338246000, 1338249600, 
    1338253200, 1338256800, 1338260400, 1338264000, 1338267600, 1338271200, 
    1338274800, 1338278400, 1338282000, 1338285600, 1338289200, 1338292800, 
    1338296400, 1338300000, 1338303600, 1338307200, 1338310800, 1338314400, 
    1338318000, 1338321600, 1338325200, 1338328800, 1338332400, 1338336000, 
    1338339600, 1338343200, 1338346800, 1338350400, 1338354000, 1338357600, 
    1338361200, 1338364800, 1338368400, 1338372000, 1338375600, 1338379200, 
    1338382800, 1338386400, 1338390000, 1338393600, 1338397200, 1338400800, 
    1338404400, 1338408000, 1338411600, 1338415200, 1338418800, 1338422400, 
    1338426000, 1338429600, 1338433200, 1338436800, 1338440400, 1338444000, 
    1338447600, 1338451200, 1338454800, 1338458400, 1338462000, 1338465600, 
    1338469200, 1338472800, 1338476400, 1338480000, 1338483600, 1338487200, 
    1338490800, 1338494400, 1338498000, 1338501600, 1338505200, 1338508800, 
    1338512400, 1338516000, 1338519600, 1338523200, 1338526800, 1338530400, 
    1338534000, 1338537600, 1338541200, 1338544800, 1338548400, 1338552000, 
    1338555600, 1338559200, 1338562800, 1338566400, 1338570000, 1338573600, 
    1338577200, 1338580800, 1338584400, 1338588000, 1338591600, 1338595200, 
    1338598800, 1338602400, 1338606000, 1338609600, 1338613200, 1338616800, 
    1338620400, 1338624000, 1338627600, 1338631200, 1338634800, 1338638400, 
    1338642000, 1338645600, 1338649200, 1338652800, 1338656400, 1338660000, 
    1338663600, 1338667200, 1338670800, 1338674400, 1338678000, 1338681600, 
    1338685200, 1338688800, 1338692400, 1338696000, 1338699600, 1338703200, 
    1338706800, 1338710400, 1338714000, 1338717600, 1338721200, 1338724800, 
    1338728400, 1338732000, 1338735600, 1338739200, 1338742800, 1338746400, 
    1338750000, 1338753600, 1338757200, 1338760800, 1338764400, 1338768000, 
    1338771600, 1338775200, 1338778800, 1338782400, 1338786000, 1338789600, 
    1338793200, 1338796800, 1338800400, 1338804000, 1338807600, 1338811200, 
    1338814800, 1338818400, 1338822000, 1338825600, 1338829200, 1338832800, 
    1338836400, 1338840000, 1338843600, 1338847200, 1338850800, 1338854400, 
    1338858000, 1338861600, 1338865200, 1338868800, 1338872400, 1338876000, 
    1338879600, 1338883200, 1338886800, 1338890400, 1338894000, 1338897600, 
    1338901200, 1338904800, 1338908400, 1338912000, 1338915600, 1338919200, 
    1338922800, 1338926400, 1338930000, 1338933600, 1338937200, 1338940800, 
    1338944400, 1338948000, 1338951600, 1338955200, 1338958800, 1338962400, 
    1338966000, 1338969600, 1338973200, 1338976800, 1338980400, 1338984000, 
    1338987600, 1338991200, 1338994800, 1338998400, 1339002000, 1339005600, 
    1339009200, 1339012800, 1339016400, 1339020000, 1339023600, 1339027200, 
    1339030800, 1339034400, 1339038000, 1339041600, 1339045200, 1339048800, 
    1339052400, 1339056000, 1339059600, 1339063200, 1339066800, 1339070400, 
    1339074000, 1339077600, 1339081200, 1339084800, 1339088400, 1339092000, 
    1339095600, 1339099200, 1339102800, 1339106400, 1339110000, 1339113600, 
    1339117200, 1339120800, 1339124400, 1339128000, 1339131600, 1339135200, 
    1339138800, 1339142400, 1339146000, 1339149600, 1339153200, 1339156800, 
    1339160400, 1339164000, 1339167600, 1339171200, 1339174800, 1339178400, 
    1339182000, 1339185600, 1339189200, 1339192800, 1339196400, 1339200000, 
    1339203600, 1339207200, 1339210800, 1339214400, 1339218000, 1339221600, 
    1339225200, 1339228800, 1339232400, 1339236000, 1339239600, 1339243200, 
    1339246800, 1339250400, 1339254000, 1339257600, 1339261200, 1339264800, 
    1339268400, 1339272000, 1339275600, 1339279200, 1339282800, 1339286400, 
    1339290000, 1339293600, 1339297200, 1339300800, 1339304400, 1339308000, 
    1339311600, 1339315200, 1339318800, 1339322400, 1339326000, 1339329600, 
    1339333200, 1339336800, 1339340400, 1339344000, 1339347600, 1339351200, 
    1339354800, 1339358400, 1339362000, 1339365600, 1339369200, 1339372800, 
    1339376400, 1339380000, 1339383600, 1339387200, 1339390800, 1339394400, 
    1339398000, 1339401600, 1339405200, 1339408800, 1339412400, 1339416000, 
    1339419600, 1339423200, 1339426800, 1339430400, 1339434000, 1339437600, 
    1339441200, 1339444800, 1339448400, 1339452000, 1339455600, 1339459200, 
    1339462800, 1339466400, 1339470000, 1339473600, 1339477200, 1339480800, 
    1339484400, 1339488000, 1339491600, 1339495200, 1339498800, 1339502400, 
    1339506000, 1339509600, 1339513200, 1339516800, 1339520400, 1339524000, 
    1339527600, 1339531200, 1339534800, 1339538400, 1339542000, 1339545600, 
    1339549200, 1339552800, 1339556400, 1339560000, 1339563600, 1339567200, 
    1339570800, 1339574400, 1339578000, 1339581600, 1339585200, 1339588800, 
    1339592400, 1339596000, 1339599600, 1339603200, 1339606800, 1339610400, 
    1339614000, 1339617600, 1339621200, 1339624800, 1339628400, 1339632000, 
    1339635600, 1339639200, 1339642800, 1339646400, 1339650000, 1339653600, 
    1339657200, 1339660800, 1339664400, 1339668000, 1339671600, 1339675200, 
    1339678800, 1339682400, 1339686000, 1339689600, 1339693200, 1339696800, 
    1339700400, 1339704000, 1339707600, 1339711200, 1339714800, 1339718400, 
    1339722000, 1339725600, 1339729200, 1339732800, 1339736400, 1339740000, 
    1339743600, 1339747200, 1339750800, 1339754400, 1339758000, 1339761600, 
    1339765200, 1339768800, 1339772400, 1339776000, 1339779600, 1339783200, 
    1339786800, 1339790400, 1339794000, 1339797600, 1339801200, 1339804800, 
    1339808400, 1339812000, 1339815600, 1339819200, 1339822800, 1339826400, 
    1339830000, 1339833600, 1339837200, 1339840800, 1339844400, 1339848000, 
    1339851600, 1339855200, 1339858800, 1339862400, 1339866000, 1339869600, 
    1339873200, 1339876800, 1339880400, 1339884000, 1339887600, 1339891200, 
    1339894800, 1339898400, 1339902000, 1339905600, 1339909200, 1339912800, 
    1339916400, 1339920000, 1339923600, 1339927200, 1339930800, 1339934400, 
    1339938000, 1339941600, 1339945200, 1339948800, 1339952400, 1339956000, 
    1339959600, 1339963200, 1339966800, 1339970400, 1339974000, 1339977600, 
    1339981200, 1339984800, 1339988400, 1339992000, 1339995600, 1339999200, 
    1340002800, 1340006400, 1340010000, 1340013600, 1340017200, 1340020800, 
    1340024400, 1340028000, 1340031600, 1340035200, 1340038800, 1340042400, 
    1340046000, 1340049600, 1340053200, 1340056800, 1340060400, 1340064000, 
    1340067600, 1340071200, 1340074800, 1340078400, 1340082000, 1340085600, 
    1340089200, 1340092800, 1340096400, 1340100000, 1340103600, 1340107200, 
    1340110800, 1340114400, 1340118000, 1340121600, 1340125200, 1340128800, 
    1340132400, 1340136000, 1340139600, 1340143200, 1340146800, 1340150400, 
    1340154000, 1340157600, 1340161200, 1340164800, 1340168400, 1340172000, 
    1340175600, 1340179200, 1340186400, 1340190000, 1340193600, 1340197200, 
    1340200800, 1340204400, 1340208000, 1340211600, 1340215200, 1340218800, 
    1340222400, 1340226000, 1340229600, 1340233200, 1340236800, 1340240400, 
    1340244000, 1340247600, 1340251200, 1340254800, 1340258400, 1340262000, 
    1340265600, 1340269200, 1340272800, 1340276400, 1340280000, 1340283600, 
    1340287200, 1340290800, 1340294400, 1340298000, 1340301600, 1340305200, 
    1340308800, 1340312400, 1340316000, 1340319600, 1340323200, 1340326800, 
    1340330400, 1340334000, 1340337600, 1340341200, 1340344800, 1340348400, 
    1340352000, 1340355600, 1340359200, 1340362800, 1340366400, 1340370000, 
    1340373600, 1340377200, 1340380800, 1340384400, 1340388000, 1340391600, 
    1340395200, 1340398800, 1340402400, 1340406000, 1340409600, 1340413200, 
    1340416800, 1340420400, 1340424000, 1340427600, 1340431200, 1340434800, 
    1340438400, 1340442000, 1340445600, 1340449200, 1340452800, 1340456400, 
    1340460000, 1340463600, 1340467200, 1340470800, 1340474400, 1340478000, 
    1340481600, 1340485200, 1340488800, 1340492400, 1340496000, 1340499600, 
    1340503200, 1340506800, 1340510400, 1340514000, 1340517600, 1340521200, 
    1340524800, 1340528400, 1340532000, 1340535600, 1340539200, 1340542800, 
    1340546400, 1340550000, 1340553600, 1340557200, 1340560800, 1340564400, 
    1340568000, 1340571600, 1340575200, 1340578800, 1340582400, 1340586000, 
    1340589600, 1340593200, 1340596800, 1340600400, 1340604000, 1340607600, 
    1340611200, 1340614800, 1340618400, 1340622000, 1340625600, 1340629200, 
    1340632800, 1340636400, 1340640000, 1340643600, 1340647200, 1340650800, 
    1340654400, 1340658000, 1340661600, 1340665200, 1340668800, 1340672400, 
    1340676000, 1340679600, 1340683200, 1340686800, 1340690400, 1340694000, 
    1340697600, 1340701200, 1340704800, 1340708400, 1340712000, 1340715600, 
    1340719200, 1340722800, 1340726400, 1340730000, 1340733600, 1340737200, 
    1340740800, 1340744400, 1340748000, 1340751600, 1340755200, 1340758800, 
    1340762400, 1340766000, 1340769600, 1340773200, 1340776800, 1340780400, 
    1340784000, 1340787600, 1340791200, 1340794800, 1340798400, 1340802000, 
    1340805600, 1340809200, 1340812800, 1340816400, 1340820000, 1340823600, 
    1340827200, 1340830800, 1340834400, 1340838000, 1340841600, 1340845200, 
    1340848800, 1340852400, 1340856000, 1340859600, 1340863200, 1340866800, 
    1340870400, 1340874000, 1340877600, 1340881200, 1340884800, 1340888400, 
    1340892000, 1340895600, 1340899200, 1340902800, 1340906400, 1340910000, 
    1340913600, 1340917200, 1340920800, 1340924400, 1340928000, 1340931600, 
    1340935200, 1340938800, 1340942400, 1340946000, 1340949600, 1340953200, 
    1340956800, 1340960400, 1340964000, 1340967600, 1340971200, 1340974800, 
    1340978400, 1340982000, 1340985600, 1340989200, 1340992800, 1340996400, 
    1341000000, 1341003600, 1341007200, 1341010800, 1341014400, 1341018000, 
    1341021600, 1341025200, 1341028800, 1341032400, 1341036000, 1341039600, 
    1341043200, 1341046800, 1341050400, 1341054000, 1341057600, 1341061200, 
    1341064800, 1341068400, 1341072000, 1341075600, 1341079200, 1341082800, 
    1341086400, 1341090000, 1341093600, 1341097200, 1341100800, 1341104400, 
    1341108000, 1341111600, 1341115200, 1341118800, 1341122400, 1341126000, 
    1341129600, 1341133200, 1341136800, 1341140400, 1341144000, 1341147600, 
    1341151200, 1341154800, 1341158400, 1341162000, 1341165600, 1341169200, 
    1341172800, 1341176400, 1341180000, 1341183600, 1341187200, 1341190800, 
    1341194400, 1341198000, 1341201600, 1341205200, 1341208800, 1341212400, 
    1341216000, 1341219600, 1341223200, 1341226800, 1341230400, 1341234000, 
    1341237600, 1341241200, 1341244800, 1341248400, 1341252000, 1341255600, 
    1341259200, 1341262800, 1341266400, 1341270000, 1341273600, 1341277200, 
    1341280800, 1341284400, 1341288000, 1341291600, 1341295200, 1341298800, 
    1341302400, 1341306000, 1341309600, 1341313200, 1341316800, 1341320400, 
    1341324000, 1341327600, 1341331200, 1341334800, 1341338400, 1341342000, 
    1341345600, 1341349200, 1341352800, 1341356400, 1341360000, 1341363600, 
    1341367200, 1341370800, 1341374400, 1341378000, 1341381600, 1341385200, 
    1341388800, 1341392400, 1341396000, 1341399600, 1341403200, 1341406800, 
    1341410400, 1341414000, 1341417600, 1341421200, 1341424800, 1341428400, 
    1341432000, 1341435600, 1341439200, 1341442800, 1341446400, 1341450000, 
    1341453600, 1341457200, 1341460800, 1341464400, 1341468000, 1341471600, 
    1341475200, 1341478800, 1341482400, 1341486000, 1341489600, 1341493200, 
    1341496800, 1341500400, 1341504000, 1341507600, 1341511200, 1341514800, 
    1341518400, 1341522000, 1341525600, 1341529200, 1341532800, 1341536400, 
    1341540000, 1341543600, 1341547200, 1341550800, 1341554400, 1341558000, 
    1341561600, 1341565200, 1341568800, 1341572400, 1341576000, 1341579600, 
    1341583200, 1341586800, 1341590400, 1341594000, 1341597600, 1341601200, 
    1341604800, 1341608400, 1341612000, 1341615600, 1341619200, 1341622800, 
    1341626400, 1341630000, 1341633600, 1341637200, 1341640800, 1341644400, 
    1341648000, 1341651600, 1341655200, 1341658800, 1341662400, 1341666000, 
    1341669600, 1341673200, 1341676800, 1341680400, 1341684000, 1341687600, 
    1341691200, 1341694800, 1341698400, 1341702000, 1341705600, 1341709200, 
    1341712800, 1341716400, 1341720000, 1341723600, 1341727200, 1341730800, 
    1341734400, 1341738000, 1341741600, 1341745200, 1341748800, 1341752400, 
    1341756000, 1341759600, 1341763200, 1341766800, 1341770400, 1341774000, 
    1341777600, 1341781200, 1341784800, 1341788400, 1341792000, 1341795600, 
    1341799200, 1341802800, 1341806400, 1341810000, 1341813600, 1341817200, 
    1341820800, 1341824400, 1341828000, 1341831600, 1341835200, 1341838800, 
    1341842400, 1341846000, 1341849600, 1341853200, 1341856800, 1341860400, 
    1341864000, 1341867600, 1341871200, 1341874800, 1341878400, 1341882000, 
    1341885600, 1341889200, 1341892800, 1341896400, 1341900000, 1341903600, 
    1341907200, 1341910800, 1341914400, 1341918000, 1341921600, 1341925200, 
    1341928800, 1341932400, 1341936000, 1341939600, 1341943200, 1341946800, 
    1341950400, 1341954000, 1341957600, 1341961200, 1341964800, 1341968400, 
    1341972000, 1341975600, 1341979200, 1341982800, 1341986400, 1341990000, 
    1341993600, 1341997200, 1342000800, 1342004400, 1342008000, 1342011600, 
    1342015200, 1342018800, 1342022400, 1342026000, 1342029600, 1342033200, 
    1342036800, 1342040400, 1342044000, 1342047600, 1342051200, 1342054800, 
    1342058400, 1342062000, 1342065600, 1342069200, 1342072800, 1342076400, 
    1342080000, 1342083600, 1342087200, 1342090800, 1342094400, 1342098000, 
    1342101600, 1342105200, 1342108800, 1342112400, 1342116000, 1342119600, 
    1342123200, 1342126800, 1342130400, 1342134000, 1342137600, 1342141200, 
    1342144800, 1342148400, 1342152000, 1342155600, 1342159200, 1342162800, 
    1342166400, 1342170000, 1342173600, 1342177200, 1342180800, 1342184400, 
    1342188000, 1342191600, 1342195200, 1342198800, 1342202400, 1342206000, 
    1342209600, 1342213200, 1342216800, 1342220400, 1342224000, 1342227600, 
    1342231200, 1342234800, 1342238400, 1342242000, 1342245600, 1342249200, 
    1342252800, 1342256400, 1342260000, 1342263600, 1342267200, 1342270800, 
    1342274400, 1342278000, 1342281600, 1342285200, 1342288800, 1342292400, 
    1342296000, 1342299600, 1342303200, 1342306800, 1342310400, 1342314000, 
    1342317600, 1342321200, 1342324800, 1342328400, 1342332000, 1342335600, 
    1342339200, 1342342800, 1342346400, 1342350000, 1342353600, 1342357200, 
    1342360800, 1342364400, 1342368000, 1342371600, 1342375200, 1342378800, 
    1342382400, 1342386000, 1342389600, 1342393200, 1342396800, 1342400400, 
    1342404000, 1342407600, 1342411200, 1342414800, 1342418400, 1342422000, 
    1342425600, 1342429200, 1342432800, 1342436400, 1342440000, 1342443600, 
    1342447200, 1342450800, 1342454400, 1342458000, 1342461600, 1342465200, 
    1342468800, 1342472400, 1342476000, 1342479600, 1342483200, 1342486800, 
    1342490400, 1342494000, 1342497600, 1342501200, 1342504800, 1342508400, 
    1342512000, 1342515600, 1342519200, 1342522800, 1342526400, 1342530000, 
    1342533600, 1342537200, 1342540800, 1342544400, 1342548000, 1342551600, 
    1342555200, 1342558800, 1342562400, 1342566000, 1342569600, 1342573200, 
    1342576800, 1342580400, 1342584000, 1342587600, 1342591200, 1342594800, 
    1342598400, 1342602000, 1342605600, 1342609200, 1342612800, 1342616400, 
    1342620000, 1342623600, 1342627200, 1342630800, 1342634400, 1342638000, 
    1342641600, 1342645200, 1342648800, 1342652400, 1342656000, 1342659600, 
    1342663200, 1342666800, 1342670400, 1342674000, 1342677600, 1342681200, 
    1342684800, 1342688400, 1342692000, 1342695600, 1342699200, 1342702800, 
    1342706400, 1342710000, 1342713600, 1342717200, 1342720800, 1342724400, 
    1342728000, 1342731600, 1342735200, 1342738800, 1342742400, 1342746000, 
    1342749600, 1342753200, 1342756800, 1342760400, 1342764000, 1342767600, 
    1342771200, 1342774800, 1342778400, 1342782000, 1342785600, 1342789200, 
    1342792800, 1342796400, 1342800000, 1342803600, 1342807200, 1342810800, 
    1342814400, 1342818000, 1342821600, 1342825200, 1342828800, 1342832400, 
    1342836000, 1342839600, 1342843200, 1342846800, 1342850400, 1342854000, 
    1342857600, 1342861200, 1342864800, 1342868400, 1342872000, 1342875600, 
    1342879200, 1342882800, 1342886400, 1342890000, 1342893600, 1342897200, 
    1342900800, 1342904400, 1342908000, 1342911600, 1342915200, 1342918800, 
    1342922400, 1342926000, 1342929600, 1342933200, 1342936800, 1342940400, 
    1342944000, 1342947600, 1342951200, 1342954800, 1342958400, 1342962000, 
    1342965600, 1342969200, 1342972800, 1342976400, 1342980000, 1342983600, 
    1342987200, 1342990800, 1342994400, 1342998000, 1343001600, 1343005200, 
    1343008800, 1343012400, 1343016000, 1343019600, 1343023200, 1343026800, 
    1343030400, 1343034000, 1343037600, 1343041200, 1343044800, 1343048400, 
    1343052000, 1343055600, 1343059200, 1343062800, 1343066400, 1343070000, 
    1343073600, 1343077200, 1343080800, 1343084400, 1343088000, 1343091600, 
    1343095200, 1343098800, 1343102400, 1343106000, 1343109600, 1343113200, 
    1343116800, 1343120400, 1343124000, 1343127600, 1343131200, 1343134800, 
    1343138400, 1343142000, 1343145600, 1343149200, 1343152800, 1343156400, 
    1343160000, 1343163600, 1343167200, 1343170800, 1343174400, 1343178000, 
    1343181600, 1343185200, 1343188800, 1343192400, 1343196000, 1343199600, 
    1343203200, 1343206800, 1343210400, 1343214000, 1343217600, 1343221200, 
    1343224800, 1343228400, 1343232000, 1343235600, 1343239200, 1343242800, 
    1343246400, 1343250000, 1343253600, 1343257200, 1343260800, 1343264400, 
    1343268000, 1343271600, 1343275200, 1343278800, 1343282400, 1343286000, 
    1343289600, 1343293200, 1343296800, 1343300400, 1343304000, 1343307600, 
    1343311200, 1343314800, 1343318400, 1343322000, 1343325600, 1343329200, 
    1343332800, 1343336400, 1343340000, 1343343600, 1343347200, 1343350800, 
    1343354400, 1343358000, 1343361600, 1343365200, 1343368800, 1343372400, 
    1343376000, 1343379600, 1343383200, 1343386800, 1343390400, 1343394000, 
    1343397600, 1343401200, 1343404800, 1343408400, 1343412000, 1343415600, 
    1343419200, 1343422800, 1343426400, 1343430000, 1343433600, 1343437200, 
    1343440800, 1343444400, 1343448000, 1343451600, 1343455200, 1343458800, 
    1343462400, 1343466000, 1343469600, 1343473200, 1343476800, 1343480400, 
    1343484000, 1343487600, 1343491200, 1343494800, 1343498400, 1343502000, 
    1343505600, 1343509200, 1343512800, 1343516400, 1343520000, 1343523600, 
    1343527200, 1343530800, 1343534400, 1343538000, 1343541600, 1343545200, 
    1343548800, 1343552400, 1343556000, 1343559600, 1343563200, 1343566800, 
    1343570400, 1343574000, 1343577600, 1343581200, 1343584800, 1343588400, 
    1343592000, 1343595600, 1343599200, 1343602800, 1343606400, 1343610000, 
    1343613600, 1343617200, 1343620800, 1343624400, 1343628000, 1343631600, 
    1343635200, 1343638800, 1343642400, 1343646000, 1343649600, 1343653200, 
    1343656800, 1343660400, 1343664000, 1343667600, 1343671200, 1343674800, 
    1343678400, 1343682000, 1343685600, 1343689200, 1343692800, 1343696400, 
    1343700000, 1343703600, 1343707200, 1343710800, 1343714400, 1343718000, 
    1343721600, 1343725200, 1343728800, 1343732400, 1343736000, 1343739600, 
    1343743200, 1343746800, 1343750400, 1343754000, 1343757600, 1343761200, 
    1343764800, 1343768400, 1343772000, 1343775600, 1343779200, 1343782800, 
    1343786400, 1343790000, 1343793600, 1343797200, 1343800800, 1343804400, 
    1343808000, 1343811600, 1343815200, 1343818800, 1343822400, 1343826000, 
    1343829600, 1343833200, 1343836800, 1343840400, 1343844000, 1343847600, 
    1343851200, 1343854800, 1343858400, 1343862000, 1343865600, 1343869200, 
    1343872800, 1343876400, 1343880000, 1343883600, 1343887200, 1343890800, 
    1343894400, 1343898000, 1343901600, 1343905200, 1343908800, 1343912400, 
    1343916000, 1343919600, 1343923200, 1343926800, 1343930400, 1343934000, 
    1343937600, 1343941200, 1343944800, 1343948400, 1343952000, 1343955600, 
    1343959200, 1343962800, 1343966400, 1343970000, 1343973600, 1343977200, 
    1343980800, 1343984400, 1343988000, 1343991600, 1343995200, 1343998800, 
    1344002400, 1344006000, 1344009600, 1344013200, 1344016800, 1344020400, 
    1344024000, 1344027600, 1344031200, 1344034800, 1344038400, 1344042000, 
    1344045600, 1344049200, 1344052800, 1344056400, 1344060000, 1344063600, 
    1344067200, 1344070800, 1344074400, 1344078000, 1344081600, 1344085200, 
    1344088800, 1344092400, 1344096000, 1344099600, 1344103200, 1344106800, 
    1344110400, 1344114000, 1344117600, 1344121200, 1344124800, 1344128400, 
    1344132000, 1344135600, 1344139200, 1344142800, 1344146400, 1344150000, 
    1344153600, 1344157200, 1344160800, 1344164400, 1344168000, 1344171600, 
    1344175200, 1344178800, 1344182400, 1344186000, 1344189600, 1344193200, 
    1344196800, 1344200400, 1344204000, 1344207600, 1344211200, 1344214800, 
    1344218400, 1344222000, 1344225600, 1344229200, 1344232800, 1344236400, 
    1344240000, 1344243600, 1344247200, 1344250800, 1344254400, 1344258000, 
    1344261600, 1344265200, 1344268800, 1344272400, 1344276000, 1344279600, 
    1344283200, 1344286800, 1344290400, 1344294000, 1344297600, 1344301200, 
    1344304800, 1344308400, 1344312000, 1344315600, 1344319200, 1344322800, 
    1344326400, 1344330000, 1344333600, 1344337200, 1344340800, 1344344400, 
    1344348000, 1344351600, 1344355200, 1344358800, 1344362400, 1344366000, 
    1344369600, 1344373200, 1344376800, 1344380400, 1344384000, 1344387600, 
    1344391200, 1344394800, 1344398400, 1344402000, 1344405600, 1344409200, 
    1344412800, 1344416400, 1344420000, 1344423600, 1344427200, 1344430800, 
    1344434400, 1344438000, 1344441600, 1344445200, 1344448800, 1344452400, 
    1344456000, 1344459600, 1344463200, 1344466800, 1344470400, 1344474000, 
    1344477600, 1344481200, 1344484800, 1344488400, 1344492000, 1344495600, 
    1344499200, 1344502800, 1344506400, 1344510000, 1344513600, 1344517200, 
    1344520800, 1344524400, 1344528000, 1344531600, 1344535200, 1344538800, 
    1344542400, 1344546000, 1344549600, 1344553200, 1344556800, 1344560400, 
    1344564000, 1344567600, 1344571200, 1344574800, 1344578400, 1344582000, 
    1344585600, 1344589200, 1344592800, 1344596400, 1344600000, 1344603600, 
    1344607200, 1344610800, 1344614400, 1344618000, 1344621600, 1344625200, 
    1344628800, 1344632400, 1344636000, 1344639600, 1344643200, 1344646800, 
    1344650400, 1344654000, 1344657600, 1344661200, 1344664800, 1344668400, 
    1344672000, 1344675600, 1344679200, 1344682800, 1344686400, 1344690000, 
    1344693600, 1344697200, 1344700800, 1344704400, 1344708000, 1344711600, 
    1344715200, 1344718800, 1344722400, 1344726000, 1344729600, 1344733200, 
    1344736800, 1344740400, 1344744000, 1344747600, 1344751200, 1344754800, 
    1344758400, 1344762000, 1344765600, 1344769200, 1344772800, 1344776400, 
    1344780000, 1344783600, 1344787200, 1344790800, 1344794400, 1344798000, 
    1344801600, 1344805200, 1344808800, 1344812400, 1344816000, 1344819600, 
    1344823200, 1344826800, 1344830400, 1344834000, 1344837600, 1344841200, 
    1344844800, 1344848400, 1344852000, 1344855600, 1344859200, 1344862800, 
    1344866400, 1344870000, 1344873600, 1344877200, 1344880800, 1344884400, 
    1344888000, 1344891600, 1344895200, 1344898800, 1344902400, 1344906000, 
    1344909600, 1344913200, 1344916800, 1344920400, 1344924000, 1344927600, 
    1344931200, 1344934800, 1344938400, 1344942000, 1344945600, 1344949200, 
    1344952800, 1344956400, 1344960000, 1344963600, 1344967200, 1344970800, 
    1344974400, 1344978000, 1344981600, 1344985200, 1344988800, 1344992400, 
    1344996000, 1344999600, 1345003200, 1345006800, 1345010400, 1345014000, 
    1345017600, 1345021200, 1345024800, 1345028400, 1345032000, 1345035600, 
    1345039200, 1345042800, 1345046400, 1345050000, 1345053600, 1345057200, 
    1345060800, 1345064400, 1345068000, 1345071600, 1345075200, 1345078800, 
    1345082400, 1345086000, 1345089600, 1345093200, 1345096800, 1345100400, 
    1345104000, 1345107600, 1345111200, 1345114800, 1345118400, 1345122000, 
    1345125600, 1345129200, 1345132800, 1345136400, 1345140000, 1345143600, 
    1345147200, 1345150800, 1345154400, 1345158000, 1345161600, 1345165200, 
    1345168800, 1345172400, 1345176000, 1345179600, 1345183200, 1345186800, 
    1345190400, 1345194000, 1345197600, 1345201200, 1345204800, 1345208400, 
    1345212000, 1345215600, 1345219200, 1345222800, 1345226400, 1345230000, 
    1345233600, 1345237200, 1345240800, 1345244400, 1345248000, 1345251600, 
    1345255200, 1345258800, 1345262400, 1345266000, 1345269600, 1345273200, 
    1345276800, 1345280400, 1345284000, 1345287600, 1345291200, 1345294800, 
    1345298400, 1345302000, 1345305600, 1345309200, 1345312800, 1345316400, 
    1345320000, 1345323600, 1345327200, 1345330800, 1345334400, 1345338000, 
    1345341600, 1345345200, 1345348800, 1345352400, 1345356000, 1345359600, 
    1345363200, 1345366800, 1345370400, 1345374000, 1345377600, 1345381200, 
    1345384800, 1345388400, 1345392000, 1345395600, 1345399200, 1345402800, 
    1345406400, 1345410000, 1345413600, 1345417200, 1345420800, 1345424400, 
    1345428000, 1345431600, 1345435200, 1345438800, 1345442400, 1345446000, 
    1345449600, 1345453200, 1345456800, 1345460400, 1345464000, 1345467600, 
    1345471200, 1345474800, 1345478400, 1345482000, 1345485600, 1345489200, 
    1345492800, 1345496400, 1345500000, 1345503600, 1345507200, 1345510800, 
    1345514400, 1345518000, 1345521600, 1345525200, 1345528800, 1345532400, 
    1345536000, 1345539600, 1345543200, 1345546800, 1345550400, 1345554000, 
    1345557600, 1345561200, 1345564800, 1345568400, 1345572000, 1345575600, 
    1345579200, 1345582800, 1345586400, 1345590000, 1345593600, 1345597200, 
    1345600800, 1345604400, 1345608000, 1345611600, 1345615200, 1345618800, 
    1345622400, 1345626000, 1345629600, 1345633200, 1345636800, 1345640400, 
    1345644000, 1345647600, 1345651200, 1345654800, 1345658400, 1345662000, 
    1345665600, 1345669200, 1345672800, 1345676400, 1345680000, 1345683600, 
    1345687200, 1345690800, 1345694400, 1345698000, 1345701600, 1345705200, 
    1345708800, 1345712400, 1345716000, 1345719600, 1345723200, 1345726800, 
    1345730400, 1345734000, 1345737600, 1345741200, 1345744800, 1345748400, 
    1345752000, 1345755600, 1345759200, 1345762800, 1345766400, 1345770000, 
    1345773600, 1345777200, 1345780800, 1345784400, 1345788000, 1345791600, 
    1345795200, 1345798800, 1345802400, 1345806000, 1345809600, 1345813200, 
    1345816800, 1345820400, 1345824000, 1345827600, 1345831200, 1345834800, 
    1345838400, 1345842000, 1345845600, 1345849200, 1345852800, 1345856400, 
    1345860000, 1345863600, 1345867200, 1345870800, 1345874400, 1345878000, 
    1345881600, 1345885200, 1345888800, 1345892400, 1345896000, 1345899600, 
    1345903200, 1345906800, 1345910400, 1345914000, 1345917600, 1345921200, 
    1345924800, 1345928400, 1345932000, 1345935600, 1345939200, 1345942800, 
    1345946400, 1345950000, 1345953600, 1345957200, 1345960800, 1345964400, 
    1345968000, 1345971600, 1345975200, 1345978800, 1345982400, 1345986000, 
    1345989600, 1345993200, 1345996800, 1346000400, 1346004000, 1346007600, 
    1346011200, 1346014800, 1346018400, 1346022000, 1346025600, 1346029200, 
    1346032800, 1346036400, 1346040000, 1346043600, 1346047200, 1346050800, 
    1346054400, 1346058000, 1346061600, 1346065200, 1346068800, 1346072400, 
    1346076000, 1346079600, 1346083200, 1346086800, 1346090400, 1346094000, 
    1346097600, 1346101200, 1346104800, 1346108400, 1346112000, 1346115600, 
    1346119200, 1346122800, 1346126400, 1346130000, 1346133600, 1346137200, 
    1346140800, 1346144400, 1346148000, 1346151600, 1346155200, 1346158800, 
    1346162400, 1346166000, 1346169600, 1346173200, 1346176800, 1346180400, 
    1346184000, 1346187600, 1346191200, 1346194800, 1346198400, 1346202000, 
    1346205600, 1346209200, 1346212800, 1346216400, 1346220000, 1346223600, 
    1346227200, 1346230800, 1346234400, 1346238000, 1346241600, 1346245200, 
    1346248800, 1346252400, 1346256000, 1346259600, 1346263200, 1346266800, 
    1346270400, 1346274000, 1346277600, 1346281200, 1346284800, 1346288400, 
    1346292000, 1346295600, 1346299200, 1346302800, 1346306400, 1346310000, 
    1346313600, 1346317200, 1346320800, 1346324400, 1346328000, 1346331600, 
    1346335200, 1346338800, 1346342400, 1346346000, 1346349600, 1346353200, 
    1346356800, 1346360400, 1346364000, 1346367600, 1346371200, 1346374800, 
    1346378400, 1346382000, 1346385600, 1346389200, 1346392800, 1346396400, 
    1346400000, 1346403600, 1346407200, 1346410800, 1346414400, 1346418000, 
    1346421600, 1346425200, 1346428800, 1346432400, 1346436000, 1346439600, 
    1346443200, 1346446800, 1346450400, 1346454000, 1346457600, 1346461200, 
    1346464800, 1346468400, 1346472000, 1346475600, 1346479200, 1346482800, 
    1346486400, 1346490000, 1346493600, 1346497200, 1346500800, 1346504400, 
    1346508000, 1346511600, 1346515200, 1346518800, 1346522400, 1346526000, 
    1346529600, 1346533200, 1346536800, 1346540400, 1346544000, 1346547600, 
    1346551200, 1346554800, 1346558400, 1346562000, 1346565600, 1346569200, 
    1346572800, 1346576400, 1346580000, 1346583600, 1346587200, 1346590800, 
    1346594400, 1346598000, 1346601600, 1346605200, 1346608800, 1346612400, 
    1346616000, 1346619600, 1346623200, 1346626800, 1346630400, 1346634000, 
    1346637600, 1346641200, 1346644800, 1346648400, 1346652000, 1346655600, 
    1346659200, 1346662800, 1346666400, 1346670000, 1346673600, 1346677200, 
    1346680800, 1346684400, 1346688000, 1346691600, 1346695200, 1346698800, 
    1346702400, 1346706000, 1346709600, 1346713200, 1346716800, 1346720400, 
    1346724000, 1346727600, 1346731200, 1346734800, 1346738400, 1346742000, 
    1346745600, 1346749200, 1346752800, 1346756400, 1346760000, 1346763600, 
    1346767200, 1346770800, 1346774400, 1346778000, 1346781600, 1346785200, 
    1346788800, 1346792400, 1346796000, 1346799600, 1346803200, 1346806800, 
    1346810400, 1346814000, 1346817600, 1346821200, 1346824800, 1346828400, 
    1346832000, 1346835600, 1346839200, 1346842800, 1346846400, 1346850000, 
    1346853600, 1346857200, 1346860800, 1346864400, 1346868000, 1346871600, 
    1346875200, 1346878800, 1346882400, 1346886000, 1346889600, 1346893200, 
    1346896800, 1346900400, 1346904000, 1346907600, 1346911200, 1346914800, 
    1346918400, 1346922000, 1346925600, 1346929200, 1346932800, 1346936400, 
    1346940000, 1346943600, 1346947200, 1346950800, 1346954400, 1346958000, 
    1346961600, 1346965200, 1346968800, 1346972400, 1346976000, 1346979600, 
    1346983200, 1346986800, 1346990400, 1346994000, 1346997600, 1347001200, 
    1347004800, 1347008400, 1347012000, 1347015600, 1347019200, 1347022800, 
    1347026400, 1347030000, 1347033600, 1347037200, 1347040800, 1347044400, 
    1347048000, 1347051600, 1347055200, 1347058800, 1347062400, 1347066000, 
    1347069600, 1347073200, 1347076800, 1347080400, 1347084000, 1347087600, 
    1347091200, 1347094800, 1347098400, 1347102000, 1347105600, 1347109200, 
    1347112800, 1347116400, 1347120000, 1347123600, 1347127200, 1347130800, 
    1347134400, 1347138000, 1347141600, 1347145200, 1347148800, 1347152400, 
    1347156000, 1347159600, 1347163200, 1347166800, 1347170400, 1347174000, 
    1347177600, 1347181200, 1347184800, 1347188400, 1347192000, 1347195600, 
    1347199200, 1347202800, 1347206400, 1347210000, 1347213600, 1347217200, 
    1347220800, 1347224400, 1347228000, 1347231600, 1347235200, 1347238800, 
    1347242400, 1347246000, 1347249600, 1347253200, 1347256800, 1347260400, 
    1347264000, 1347267600, 1347271200, 1347274800, 1347278400, 1347282000, 
    1347285600, 1347289200, 1347292800, 1347296400, 1347300000, 1347303600, 
    1347307200, 1347310800, 1347314400, 1347318000, 1347321600, 1347325200, 
    1347328800, 1347332400, 1347336000, 1347339600, 1347343200, 1347346800, 
    1347350400, 1347354000, 1347357600, 1347361200, 1347364800, 1347368400, 
    1347372000, 1347375600, 1347379200, 1347382800, 1347386400, 1347390000, 
    1347393600, 1347397200, 1347400800, 1347404400, 1347408000, 1347411600, 
    1347415200, 1347418800, 1347422400, 1347426000, 1347429600, 1347433200, 
    1347436800, 1347440400, 1347444000, 1347447600, 1347451200, 1347454800, 
    1347458400, 1347462000, 1347465600, 1347469200, 1347472800, 1347476400, 
    1347480000, 1347483600, 1347487200, 1347490800, 1347494400, 1347498000, 
    1347501600, 1347505200, 1347508800, 1347512400, 1347516000, 1347519600, 
    1347523200, 1347526800, 1347530400, 1347534000, 1347537600, 1347541200, 
    1347544800, 1347548400, 1347552000, 1347555600, 1347559200, 1347562800, 
    1347566400, 1347570000, 1347573600, 1347577200, 1347580800, 1347584400, 
    1347588000, 1347591600, 1347595200, 1347598800, 1347602400, 1347606000, 
    1347609600, 1347613200, 1347616800, 1347620400, 1347624000, 1347627600, 
    1347631200, 1347634800, 1347638400, 1347642000, 1347645600, 1347649200, 
    1347652800, 1347656400, 1347660000, 1347663600, 1347667200, 1347670800, 
    1347674400, 1347678000, 1347681600, 1347685200, 1347688800, 1347692400, 
    1347696000, 1347699600, 1347703200, 1347706800, 1347710400, 1347714000, 
    1347717600, 1347721200, 1347724800, 1347728400, 1347732000, 1347735600, 
    1347739200, 1347742800, 1347746400, 1347750000, 1347753600, 1347757200, 
    1347760800, 1347764400, 1347768000, 1347771600, 1347775200, 1347778800, 
    1347782400, 1347786000, 1347789600, 1347793200, 1347796800, 1347800400, 
    1347804000, 1347807600, 1347811200, 1347814800, 1347818400, 1347822000, 
    1347825600, 1347829200, 1347832800, 1347836400, 1347840000, 1347843600, 
    1347847200, 1347850800, 1347854400, 1347858000, 1347861600, 1347865200, 
    1347868800, 1347872400, 1347876000, 1347879600, 1347883200, 1347886800, 
    1347890400, 1347894000, 1347897600, 1347901200, 1347904800, 1347908400, 
    1347912000, 1347915600, 1347919200, 1347922800, 1347926400, 1347930000, 
    1347933600, 1347937200, 1347940800, 1347944400, 1347948000, 1347951600, 
    1347955200, 1347958800, 1347962400, 1347966000, 1347969600, 1347973200, 
    1347976800, 1347980400, 1347984000, 1347987600, 1347991200, 1347994800, 
    1347998400, 1348002000, 1348005600, 1348009200, 1348012800, 1348016400, 
    1348020000, 1348023600, 1348027200, 1348030800, 1348034400, 1348038000, 
    1348041600, 1348045200, 1348048800, 1348052400, 1348056000, 1348059600, 
    1348063200, 1348066800, 1348070400, 1348074000, 1348077600, 1348081200, 
    1348084800, 1348088400, 1348092000, 1348095600, 1348099200, 1348102800, 
    1348106400, 1348110000, 1348113600, 1348117200, 1348120800, 1348124400, 
    1348128000, 1348131600, 1348135200, 1348138800, 1348142400, 1348146000, 
    1348149600, 1348153200, 1348156800, 1348160400, 1348164000, 1348167600, 
    1348171200, 1348174800, 1348178400, 1348182000, 1348185600, 1348189200, 
    1348192800, 1348196400, 1348200000, 1348203600, 1348207200, 1348210800, 
    1348214400, 1348218000, 1348221600, 1348225200, 1348228800, 1348232400, 
    1348236000, 1348239600, 1348243200, 1348246800, 1348250400, 1348254000, 
    1348257600, 1348261200, 1348264800, 1348268400, 1348272000, 1348275600, 
    1348279200, 1348282800, 1348286400, 1348290000, 1348293600, 1348297200, 
    1348300800, 1348304400, 1348308000, 1348311600, 1348315200, 1348318800, 
    1348322400, 1348326000, 1348329600, 1348333200, 1348336800, 1348340400, 
    1348344000, 1348347600, 1348351200, 1348354800, 1348358400, 1348362000, 
    1348365600, 1348369200, 1348372800, 1348376400, 1348380000, 1348383600, 
    1348387200, 1348390800, 1348394400, 1348398000, 1348401600, 1348405200, 
    1348408800, 1348412400, 1348416000, 1348419600, 1348423200, 1348426800, 
    1348430400, 1348434000, 1348437600, 1348441200, 1348444800, 1348448400, 
    1348452000, 1348455600, 1348459200, 1348462800, 1348466400, 1348470000, 
    1348473600, 1348477200, 1348480800, 1348484400, 1348488000, 1348491600, 
    1348495200, 1348498800, 1348502400, 1348506000, 1348509600, 1348513200, 
    1348516800, 1348520400, 1348524000, 1348527600, 1348531200, 1348534800, 
    1348538400, 1348542000, 1348545600, 1348549200, 1348552800, 1348556400, 
    1348560000, 1348563600, 1348567200, 1348570800, 1348574400, 1348578000, 
    1348581600, 1348585200, 1348588800, 1348592400, 1348596000, 1348599600, 
    1348603200, 1348606800, 1348610400, 1348614000, 1348617600, 1348621200, 
    1348624800, 1348628400, 1348632000, 1348635600, 1348639200, 1348642800, 
    1348646400, 1348650000, 1348653600, 1348657200, 1348660800, 1348664400, 
    1348668000, 1348671600, 1348675200, 1348678800, 1348682400, 1348686000, 
    1348689600, 1348693200, 1348696800, 1348700400, 1348704000, 1348707600, 
    1348711200, 1348714800, 1348718400, 1348722000, 1348725600, 1348729200, 
    1348732800, 1348736400, 1348740000, 1348743600, 1348747200, 1348750800, 
    1348754400, 1348758000, 1348761600, 1348765200, 1348768800, 1348772400, 
    1348776000, 1348779600, 1348783200, 1348786800, 1348790400, 1348794000, 
    1348797600, 1348801200, 1348804800, 1348808400, 1348812000, 1348815600, 
    1348819200, 1348822800, 1348826400, 1348830000, 1348833600, 1348837200, 
    1348840800, 1348844400, 1348848000, 1348851600, 1348855200, 1348858800, 
    1348862400, 1348866000, 1348869600, 1348873200, 1348876800, 1348880400, 
    1348884000, 1348887600, 1348891200, 1348894800, 1348898400, 1348902000, 
    1348905600, 1348909200, 1348912800, 1348916400, 1348920000, 1348923600, 
    1348927200, 1348930800, 1348934400, 1348938000, 1348941600, 1348945200, 
    1348948800, 1348952400, 1348956000, 1348959600, 1348963200, 1348966800, 
    1348970400, 1348974000, 1348977600, 1348981200, 1348984800, 1348988400, 
    1348992000, 1348995600, 1348999200, 1349002800, 1349006400, 1349010000, 
    1349013600, 1349017200, 1349020800, 1349024400, 1349028000, 1349031600, 
    1349035200, 1349038800, 1349042400, 1349046000, 1349049600, 1349053200, 
    1349056800, 1349060400, 1349064000, 1349067600, 1349071200, 1349074800, 
    1349078400, 1349082000, 1349085600, 1349089200, 1349092800, 1349096400, 
    1349100000, 1349103600, 1349107200, 1349110800, 1349114400, 1349118000, 
    1349121600, 1349125200, 1349128800, 1349132400, 1349136000, 1349139600, 
    1349143200, 1349146800, 1349150400, 1349154000, 1349157600, 1349161200, 
    1349164800, 1349168400, 1349172000, 1349175600, 1349179200, 1349182800, 
    1349186400, 1349190000, 1349193600, 1349197200, 1349200800, 1349204400, 
    1349208000, 1349211600, 1349215200, 1349218800, 1349222400, 1349226000, 
    1349229600, 1349233200, 1349236800, 1349240400, 1349244000, 1349247600, 
    1349251200, 1349254800, 1349258400, 1349262000, 1349265600, 1349269200, 
    1349272800, 1349276400, 1349280000, 1349283600, 1349287200, 1349290800, 
    1349294400, 1349298000, 1349301600, 1349305200, 1349308800, 1349312400, 
    1349316000, 1349319600, 1349323200, 1349326800, 1349330400, 1349334000, 
    1349337600, 1349341200, 1349344800, 1349348400, 1349352000, 1349355600, 
    1349359200, 1349362800, 1349366400, 1349370000, 1349373600, 1349377200, 
    1349380800, 1349384400, 1349388000, 1349391600, 1349395200, 1349398800, 
    1349402400, 1349406000, 1349409600, 1349413200, 1349416800, 1349420400, 
    1349424000, 1349427600, 1349431200, 1349434800, 1349438400, 1349442000, 
    1349445600, 1349449200, 1349452800, 1349456400, 1349460000, 1349463600, 
    1349467200, 1349470800, 1349474400, 1349478000, 1349481600, 1349485200, 
    1349488800, 1349492400, 1349496000, 1349499600, 1349503200, 1349506800, 
    1349510400, 1349514000, 1349517600, 1349521200, 1349524800, 1349528400, 
    1349532000, 1349535600, 1349539200, 1349542800, 1349546400, 1349550000, 
    1349553600, 1349557200, 1349560800, 1349564400, 1349568000, 1349571600, 
    1349575200, 1349578800, 1349582400, 1349586000, 1349589600, 1349593200, 
    1349596800, 1349600400, 1349604000, 1349607600, 1349611200, 1349614800, 
    1349618400, 1349622000, 1349625600, 1349629200, 1349632800, 1349636400, 
    1349640000, 1349643600, 1349647200, 1349650800, 1349654400, 1349658000, 
    1349661600, 1349665200, 1349668800, 1349672400, 1349676000, 1349679600, 
    1349683200, 1349686800, 1349690400, 1349694000, 1349697600, 1349701200, 
    1349704800, 1349708400, 1349712000, 1349715600, 1349719200, 1349722800, 
    1349726400, 1349730000, 1349733600, 1349737200, 1349740800, 1349744400, 
    1349748000, 1349751600, 1349755200, 1349758800, 1349762400, 1349766000, 
    1349769600, 1349773200, 1349776800, 1349780400, 1349784000, 1349787600, 
    1349791200, 1349794800, 1349798400, 1349802000, 1349805600, 1349809200, 
    1349812800, 1349816400, 1349820000, 1349823600, 1349827200, 1349830800, 
    1349834400, 1349838000, 1349841600, 1349845200, 1349848800, 1349852400, 
    1349856000, 1349859600, 1349863200, 1349866800, 1349870400, 1349874000, 
    1349877600, 1349881200, 1349884800, 1349888400, 1349892000, 1349895600, 
    1349899200, 1349902800, 1349906400, 1349910000, 1349913600, 1349917200, 
    1349920800, 1349924400, 1349928000, 1349931600, 1349935200, 1349938800, 
    1349942400, 1349946000, 1349949600, 1349953200, 1349956800, 1349960400, 
    1349964000, 1349967600, 1349971200, 1349974800, 1349978400, 1349982000, 
    1349985600, 1349989200, 1349992800, 1349996400, 1350000000, 1350003600, 
    1350007200, 1350010800, 1350014400, 1350018000, 1350021600, 1350025200, 
    1350028800, 1350032400, 1350036000, 1350039600, 1350043200, 1350046800, 
    1350050400, 1350054000, 1350057600, 1350061200, 1350064800, 1350068400, 
    1350072000, 1350075600, 1350079200, 1350082800, 1350086400, 1350090000, 
    1350093600, 1350097200, 1350100800, 1350104400, 1350108000, 1350111600, 
    1350115200, 1350118800, 1350122400, 1350126000, 1350129600, 1350133200, 
    1350136800, 1350140400, 1350144000, 1350147600, 1350151200, 1350154800, 
    1350158400, 1350162000, 1350165600, 1350169200, 1350172800, 1350176400, 
    1350180000, 1350183600, 1350187200, 1350190800, 1350194400, 1350198000, 
    1350201600, 1350205200, 1350208800, 1350212400, 1350216000, 1350219600, 
    1350223200, 1350226800, 1350230400, 1350234000, 1350237600, 1350241200, 
    1350244800, 1350248400, 1350252000, 1350255600, 1350259200, 1350262800, 
    1350266400, 1350270000, 1350273600, 1350277200, 1350280800, 1350284400, 
    1350288000, 1350291600, 1350295200, 1350298800, 1350302400, 1350306000, 
    1350309600, 1350313200, 1350316800, 1350320400, 1350324000, 1350327600, 
    1350331200, 1350334800, 1350338400, 1350342000, 1350345600, 1350349200, 
    1350352800, 1350356400, 1350360000, 1350363600, 1350367200, 1350370800, 
    1350374400, 1350378000, 1350381600, 1350385200, 1350388800, 1350392400, 
    1350396000, 1350399600, 1350403200, 1350406800, 1350410400, 1350414000, 
    1350417600, 1350421200, 1350424800, 1350428400, 1350432000, 1350435600, 
    1350439200, 1350442800, 1350446400, 1350450000, 1350453600, 1350457200, 
    1350460800, 1350464400, 1350468000, 1350471600, 1350475200, 1350478800, 
    1350482400, 1350486000, 1350489600, 1350493200, 1350496800, 1350500400, 
    1350504000, 1350507600, 1350511200, 1350514800, 1350518400, 1350522000, 
    1350525600, 1350529200, 1350532800, 1350536400, 1350540000, 1350543600, 
    1350547200, 1350550800, 1350554400, 1350558000, 1350561600, 1350565200, 
    1350568800, 1350572400, 1350576000, 1350579600, 1350583200, 1350586800, 
    1350590400, 1350594000, 1350597600, 1350601200, 1350604800, 1350608400, 
    1350612000, 1350615600, 1350619200, 1350622800, 1350626400, 1350630000, 
    1350633600, 1350637200, 1350640800, 1350644400, 1350648000, 1350651600, 
    1350655200, 1350658800, 1350662400, 1350666000, 1350669600, 1350673200, 
    1350676800, 1350680400, 1350684000, 1350687600, 1350691200, 1350694800, 
    1350698400, 1350702000, 1350705600, 1350709200, 1350712800, 1350716400, 
    1350720000, 1350723600, 1350727200, 1350730800, 1350734400, 1350738000, 
    1350741600, 1350745200, 1350748800, 1350752400, 1350756000, 1350759600, 
    1350763200, 1350766800, 1350770400, 1350774000, 1350777600, 1350781200, 
    1350784800, 1350788400, 1350792000, 1350795600, 1350799200, 1350802800, 
    1350806400, 1350810000, 1350813600, 1350817200, 1350820800, 1350824400, 
    1350828000, 1350831600, 1350835200, 1350838800, 1350842400, 1350846000, 
    1350849600, 1350853200, 1350856800, 1350860400, 1350864000, 1350867600, 
    1350871200, 1350874800, 1350878400, 1350882000, 1350885600, 1350889200, 
    1350892800, 1350896400, 1350900000, 1350903600, 1350907200, 1350910800, 
    1350914400, 1350918000, 1350921600, 1350925200, 1350928800, 1350932400, 
    1350936000, 1350939600, 1350943200, 1350946800, 1350950400, 1350954000, 
    1350957600, 1350961200, 1350964800, 1350968400, 1350972000, 1350975600, 
    1350979200, 1350982800, 1350986400, 1350990000, 1350993600, 1350997200, 
    1351000800, 1351004400, 1351008000, 1351011600, 1351015200, 1351018800, 
    1351022400, 1351026000, 1351029600, 1351033200, 1351036800, 1351040400, 
    1351044000, 1351047600, 1351051200, 1351054800, 1351058400, 1351062000, 
    1351065600, 1351069200, 1351072800, 1351076400, 1351080000, 1351083600, 
    1351087200, 1351090800, 1351094400, 1351098000, 1351101600, 1351105200, 
    1351108800, 1351112400, 1351116000, 1351119600, 1351123200, 1351126800, 
    1351130400, 1351134000, 1351137600, 1351141200, 1351144800, 1351148400, 
    1351152000, 1351155600, 1351159200, 1351162800, 1351166400, 1351170000, 
    1351173600, 1351177200, 1351180800, 1351184400, 1351188000, 1351191600, 
    1351195200, 1351198800, 1351202400, 1351206000, 1351209600, 1351213200, 
    1351216800, 1351220400, 1351224000, 1351227600, 1351231200, 1351234800, 
    1351238400, 1351242000, 1351245600, 1351249200, 1351252800, 1351256400, 
    1351260000, 1351263600, 1351267200, 1351270800, 1351274400, 1351278000, 
    1351281600, 1351285200, 1351288800, 1351292400, 1351296000, 1351299600, 
    1351303200, 1351306800, 1351310400, 1351314000, 1351317600, 1351321200, 
    1351324800, 1351328400, 1351332000, 1351335600, 1351339200, 1351342800, 
    1351346400, 1351350000, 1351353600, 1351357200, 1351360800, 1351364400, 
    1351368000, 1351371600, 1351375200, 1351378800, 1351382400, 1351386000, 
    1351389600, 1351393200, 1351396800, 1351400400, 1351404000, 1351407600, 
    1351411200, 1351414800, 1351418400, 1351422000, 1351425600, 1351429200, 
    1351432800, 1351436400, 1351440000, 1351443600, 1351447200, 1351450800, 
    1351454400, 1351458000, 1351461600, 1351465200, 1351468800, 1351472400, 
    1351476000, 1351479600, 1351483200, 1351486800, 1351490400, 1351494000, 
    1351497600, 1351501200, 1351504800, 1351508400, 1351512000, 1351515600, 
    1351519200, 1351522800, 1351526400, 1351530000, 1351533600, 1351537200, 
    1351540800, 1351544400, 1351591200, 1351594800, 1351598400, 1351602000, 
    1351605600, 1351609200, 1351612800, 1351616400, 1351620000, 1351623600, 
    1351627200, 1351630800, 1351634400, 1351638000, 1351641600, 1351645200, 
    1351648800, 1351652400, 1351656000, 1351659600, 1351663200, 1351666800, 
    1351670400, 1351674000, 1351677600, 1351681200, 1351684800, 1351688400, 
    1351692000, 1351695600, 1351699200, 1351702800, 1351706400, 1351710000, 
    1351713600, 1351717200, 1351720800, 1351724400, 1351728000, 1351731600, 
    1351735200, 1351738800, 1351742400, 1351746000, 1351749600, 1351753200, 
    1351756800, 1351760400, 1351764000, 1351767600, 1351771200, 1351774800, 
    1351778400, 1351782000, 1351785600, 1351789200, 1351792800, 1351796400, 
    1351800000, 1351803600, 1351807200, 1351810800, 1351814400, 1351818000, 
    1351821600, 1351825200, 1351828800, 1351832400, 1351836000, 1351839600, 
    1351843200, 1351846800, 1351850400, 1351854000, 1351857600, 1351861200, 
    1351864800, 1351868400, 1351872000, 1351875600, 1351879200, 1351882800, 
    1351886400, 1351890000, 1351893600, 1351897200, 1351900800, 1351904400, 
    1351908000, 1351911600, 1351915200, 1351918800, 1351922400, 1351926000, 
    1351929600, 1351933200, 1351936800, 1351940400, 1351944000, 1351947600, 
    1351951200, 1351954800, 1351958400, 1351962000, 1351965600, 1351969200, 
    1351972800, 1351976400, 1351980000, 1351983600, 1351987200, 1351990800, 
    1351994400, 1351998000, 1352001600, 1352005200, 1352008800, 1352012400, 
    1352016000, 1352019600, 1352023200, 1352026800, 1352030400, 1352034000, 
    1352037600, 1352041200, 1352044800, 1352048400, 1352052000, 1352055600, 
    1352059200, 1352062800, 1352066400, 1352070000, 1352073600, 1352077200, 
    1352080800, 1352084400, 1352088000, 1352091600, 1352095200, 1352098800, 
    1352102400, 1352106000, 1352109600, 1352113200, 1352116800, 1352120400, 
    1352124000, 1352127600, 1352131200, 1352134800, 1352138400, 1352142000, 
    1352145600, 1352149200, 1352152800, 1352156400, 1352160000, 1352163600, 
    1352167200, 1352170800, 1352174400, 1352178000, 1352181600, 1352185200, 
    1352188800, 1352192400, 1352196000, 1352199600, 1352203200, 1352206800, 
    1352210400, 1352214000, 1352217600, 1352221200, 1352224800, 1352228400, 
    1352232000, 1352235600, 1352239200, 1352242800, 1352246400, 1352250000, 
    1352253600, 1352257200, 1352260800, 1352264400, 1352268000, 1352271600, 
    1352275200, 1352278800, 1352282400, 1352286000, 1352289600, 1352293200, 
    1352296800, 1352300400, 1352304000, 1352307600, 1352311200, 1352314800, 
    1352318400, 1352322000, 1352325600, 1352329200, 1352332800, 1352336400, 
    1352340000, 1352343600, 1352347200, 1352350800, 1352354400, 1352358000, 
    1352361600, 1352365200, 1352368800, 1352372400, 1352376000, 1352379600, 
    1352383200, 1352386800, 1352390400, 1352394000, 1352397600, 1352401200, 
    1352404800, 1352408400, 1352412000, 1352415600, 1352419200, 1352422800, 
    1352426400, 1352430000, 1352433600, 1352437200, 1352440800, 1352444400, 
    1352448000, 1352451600, 1352455200, 1352458800, 1352462400, 1352466000, 
    1352469600, 1352473200, 1352476800, 1352480400, 1352484000, 1352487600, 
    1352491200, 1352494800, 1352498400, 1352502000, 1352505600, 1352509200, 
    1352512800, 1352516400, 1352520000, 1352523600, 1352527200, 1352530800, 
    1352534400, 1352538000, 1352541600, 1352545200, 1352548800, 1352552400, 
    1352556000, 1352559600, 1352563200, 1352566800, 1352570400, 1352574000, 
    1352577600, 1352581200, 1352584800, 1352588400, 1352592000, 1352595600, 
    1352599200, 1352602800, 1352606400, 1352610000, 1352613600, 1352617200, 
    1352620800, 1352624400, 1352628000, 1352631600, 1352635200, 1352638800, 
    1352642400, 1352646000, 1352649600, 1352653200, 1352656800, 1352660400, 
    1352664000, 1352667600, 1352671200, 1352674800, 1352678400, 1352682000, 
    1352685600, 1352689200, 1352692800, 1352696400, 1352700000, 1352703600, 
    1352707200, 1352710800, 1352714400, 1352718000, 1352721600, 1352725200, 
    1352728800, 1352732400, 1352736000, 1352739600, 1352743200, 1352746800, 
    1352750400, 1352754000, 1352757600, 1352761200, 1352764800, 1352768400, 
    1352772000, 1352775600, 1352779200, 1352782800, 1352786400, 1352790000, 
    1352793600, 1352797200, 1352800800, 1352804400, 1352808000, 1352811600, 
    1352815200, 1352818800, 1352822400, 1352826000, 1352829600, 1352833200, 
    1352836800, 1352840400, 1352844000, 1352847600, 1352851200, 1352854800, 
    1352858400, 1352862000, 1352865600, 1352869200, 1352872800, 1352876400, 
    1352880000, 1352883600, 1352887200, 1352890800, 1352894400, 1352898000, 
    1352901600, 1352905200, 1352908800, 1352912400, 1352916000, 1352919600, 
    1352923200, 1352926800, 1352930400, 1352934000, 1352937600, 1352941200, 
    1352944800, 1352948400, 1352952000, 1352955600, 1352959200, 1352962800, 
    1352966400, 1352970000, 1352973600, 1352977200, 1352980800, 1352984400, 
    1352988000, 1352991600, 1352995200, 1352998800, 1353002400, 1353006000, 
    1353009600, 1353013200, 1353016800, 1353020400, 1353024000, 1353027600, 
    1353031200, 1353034800, 1353038400, 1353042000, 1353045600, 1353049200, 
    1353052800, 1353056400, 1353060000, 1353063600, 1353067200, 1353070800, 
    1353074400, 1353078000, 1353081600, 1353085200, 1353088800, 1353092400, 
    1353096000, 1353099600, 1353103200, 1353106800, 1353110400, 1353114000, 
    1353117600, 1353121200, 1353124800, 1353128400, 1353132000, 1353135600, 
    1353139200, 1353142800, 1353146400, 1353150000, 1353153600, 1353157200, 
    1353160800, 1353164400, 1353168000, 1353171600, 1353175200, 1353178800, 
    1353182400, 1353186000, 1353189600, 1353193200, 1353196800, 1353200400, 
    1353204000, 1353207600, 1353211200, 1353214800, 1353218400, 1353222000, 
    1353225600, 1353229200, 1353232800, 1353236400, 1353240000, 1353243600, 
    1353247200, 1353250800, 1353254400, 1353258000, 1353261600, 1353265200, 
    1353268800, 1353272400, 1353276000, 1353279600, 1353283200, 1353286800, 
    1353290400, 1353294000, 1353297600, 1353301200, 1353304800, 1353308400, 
    1353312000, 1353315600, 1353319200, 1353322800, 1353326400, 1353330000, 
    1353333600, 1353337200, 1353340800, 1353344400, 1353348000, 1353351600, 
    1353355200, 1353358800, 1353362400, 1353366000, 1353369600, 1353373200, 
    1353376800, 1353380400, 1353384000, 1353387600, 1353391200, 1353394800, 
    1353398400, 1353402000, 1353405600, 1353409200, 1353412800, 1353416400, 
    1353420000, 1353423600, 1353427200, 1353430800, 1353434400, 1353438000, 
    1353441600, 1353445200, 1353448800, 1353452400, 1353456000, 1353459600, 
    1353463200, 1353466800, 1353470400, 1353474000, 1353477600, 1353481200, 
    1353484800, 1353488400, 1353492000, 1353495600, 1353499200, 1353502800, 
    1353506400, 1353510000, 1353513600, 1353517200, 1353520800, 1353524400, 
    1353528000, 1353531600, 1353535200, 1353538800, 1353542400, 1353546000, 
    1353549600, 1353553200, 1353556800, 1353560400, 1353564000, 1353567600, 
    1353571200, 1353574800, 1353578400, 1353582000, 1353585600, 1353589200, 
    1353592800, 1353596400, 1353600000, 1353603600, 1353607200, 1353610800, 
    1353614400, 1353618000, 1353621600, 1353625200, 1353628800, 1353632400, 
    1353636000, 1353639600, 1353643200, 1353646800, 1353650400, 1353654000, 
    1353657600, 1353661200, 1353664800, 1353668400, 1353672000, 1353675600, 
    1353679200, 1353682800, 1353686400, 1353690000, 1353693600, 1353697200, 
    1353700800, 1353704400, 1353708000, 1353711600, 1353715200, 1353718800, 
    1353722400, 1353726000, 1353729600, 1353733200, 1353736800, 1353740400, 
    1353744000, 1353747600, 1353751200, 1353754800, 1353758400, 1353762000, 
    1353765600, 1353769200, 1353772800, 1353776400, 1353780000, 1353783600, 
    1353787200, 1353790800, 1353794400, 1353798000, 1353801600, 1353805200, 
    1353808800, 1353812400, 1353816000, 1353819600, 1353823200, 1353826800, 
    1353830400, 1353834000, 1353837600, 1353841200, 1353844800, 1353848400, 
    1353852000, 1353855600, 1353859200, 1353862800, 1353866400, 1353870000, 
    1353873600, 1353877200, 1353880800, 1353884400, 1353888000, 1353891600, 
    1353895200, 1353898800, 1353902400, 1353906000, 1353909600, 1353913200, 
    1353916800, 1353920400, 1353924000, 1353927600, 1353931200, 1353934800, 
    1353938400, 1353942000, 1353945600, 1353949200, 1353952800, 1353956400, 
    1353960000, 1353963600, 1353967200, 1353970800, 1353974400, 1353978000, 
    1353981600, 1353985200, 1353988800, 1353992400, 1353996000, 1353999600, 
    1354003200, 1354006800, 1354010400, 1354014000, 1354017600, 1354021200, 
    1354024800, 1354028400, 1354032000, 1354035600, 1354039200, 1354042800, 
    1354046400, 1354050000, 1354053600, 1354057200, 1354060800, 1354064400, 
    1354068000, 1354071600, 1354075200, 1354078800, 1354082400, 1354086000, 
    1354089600, 1354093200, 1354096800, 1354100400, 1354104000, 1354107600, 
    1354111200, 1354114800, 1354118400, 1354122000, 1354125600, 1354129200, 
    1354132800, 1354136400, 1354140000, 1354143600, 1354147200, 1354150800, 
    1354154400, 1354158000, 1354161600, 1354165200, 1354168800, 1354172400, 
    1354176000, 1354179600, 1354183200, 1354186800, 1354190400, 1354194000, 
    1354197600, 1354201200, 1354204800, 1354208400, 1354212000, 1354215600, 
    1354219200, 1354222800, 1354226400, 1354230000, 1354233600, 1354237200, 
    1354240800, 1354244400, 1354248000, 1354251600, 1354255200, 1354258800, 
    1354262400, 1354266000, 1354269600, 1354273200, 1354276800, 1354280400, 
    1354284000, 1354287600, 1354291200, 1354294800, 1354298400, 1354302000, 
    1354305600, 1354309200, 1354312800, 1354316400, 1354320000, 1354323600, 
    1354327200, 1354330800, 1354334400, 1354338000, 1354341600, 1354345200, 
    1354348800, 1354352400, 1354356000, 1354359600, 1354363200, 1354366800, 
    1354370400, 1354374000, 1354377600, 1354381200, 1354384800, 1354388400, 
    1354392000, 1354395600, 1354399200, 1354402800, 1354406400, 1354410000, 
    1354413600, 1354417200, 1354420800, 1354424400, 1354428000, 1354431600, 
    1354435200, 1354438800, 1354442400, 1354446000, 1354449600, 1354453200, 
    1354456800, 1354460400, 1354464000, 1354467600, 1354471200, 1354474800, 
    1354478400, 1354482000, 1354485600, 1354489200, 1354492800, 1354496400, 
    1354500000, 1354503600, 1354507200, 1354510800, 1354514400, 1354518000, 
    1354521600, 1354525200, 1354528800, 1354532400, 1354536000, 1354539600, 
    1354543200, 1354546800, 1354550400, 1354554000, 1354557600, 1354561200, 
    1354564800, 1354568400, 1354572000, 1354575600, 1354579200, 1354582800, 
    1354586400, 1354590000, 1354593600, 1354597200, 1354600800, 1354604400, 
    1354608000, 1354611600, 1354615200, 1354618800, 1354622400, 1354626000, 
    1354629600, 1354633200, 1354636800, 1354640400, 1354644000, 1354647600, 
    1354651200, 1354654800, 1354658400, 1354662000, 1354665600, 1354669200, 
    1354672800, 1354676400, 1354680000, 1354683600, 1354687200, 1354690800, 
    1354694400, 1354698000, 1354701600, 1354705200, 1354708800, 1354712400, 
    1354716000, 1354719600, 1354723200, 1354726800, 1354730400, 1354734000, 
    1354737600, 1354741200, 1354744800, 1354748400, 1354752000, 1354755600, 
    1354759200, 1354762800, 1354766400, 1354770000, 1354773600, 1354777200, 
    1354780800, 1354784400, 1354788000, 1354791600, 1354795200, 1354798800, 
    1354802400, 1354806000, 1354809600, 1354813200, 1354816800, 1354820400, 
    1354824000, 1354827600, 1354831200, 1354834800, 1354838400, 1354842000, 
    1354845600, 1354849200, 1354852800, 1354856400, 1354860000, 1354863600, 
    1354867200, 1354870800, 1354874400, 1354878000, 1354881600, 1354885200, 
    1354888800, 1354892400, 1354896000, 1354899600, 1354903200, 1354906800, 
    1354910400, 1354914000, 1354917600, 1354921200, 1354924800, 1354928400, 
    1354932000, 1354935600, 1354939200, 1354942800, 1354946400, 1354950000, 
    1354953600, 1354957200, 1354960800, 1354964400, 1354968000, 1354971600, 
    1354975200, 1354978800, 1354982400, 1354986000, 1354989600, 1354993200, 
    1354996800, 1355000400, 1355004000, 1355007600, 1355011200, 1355014800, 
    1355018400, 1355022000, 1355025600, 1355029200, 1355032800, 1355036400, 
    1355040000, 1355043600, 1355047200, 1355050800, 1355054400, 1355058000, 
    1355061600, 1355065200, 1355068800, 1355072400, 1355076000, 1355079600, 
    1355083200, 1355086800, 1355090400, 1355094000, 1355097600, 1355101200, 
    1355104800, 1355108400, 1355112000, 1355115600, 1355119200, 1355122800, 
    1355126400, 1355130000, 1355133600, 1355137200, 1355140800, 1355144400, 
    1355148000, 1355151600, 1355155200, 1355158800, 1355162400, 1355166000, 
    1355169600, 1355173200, 1355176800, 1355180400, 1355184000, 1355187600, 
    1355191200, 1355194800, 1355198400, 1355202000, 1355205600, 1355209200, 
    1355212800, 1355216400, 1355220000, 1355223600, 1355227200, 1355230800, 
    1355234400, 1355238000, 1355241600, 1355245200, 1355248800, 1355252400, 
    1355256000, 1355259600, 1355263200, 1355266800, 1355270400, 1355274000, 
    1355277600, 1355281200, 1355284800, 1355288400, 1355292000, 1355295600, 
    1355299200, 1355302800, 1355306400, 1355310000, 1355313600, 1355317200, 
    1355320800, 1355324400, 1355328000, 1355331600, 1355335200, 1355338800, 
    1355342400, 1355346000, 1355349600, 1355353200, 1355356800, 1355360400, 
    1355364000, 1355367600, 1355371200, 1355374800, 1355378400, 1355382000, 
    1355385600, 1355389200, 1355392800, 1355396400, 1355400000, 1355403600, 
    1355407200, 1355410800, 1355414400, 1355418000, 1355421600, 1355425200, 
    1355428800, 1355432400, 1355436000, 1355439600, 1355443200, 1355446800, 
    1355450400, 1355454000, 1355457600, 1355461200, 1355464800, 1355468400, 
    1355472000, 1355475600, 1355479200, 1355482800, 1355486400, 1355490000, 
    1355493600, 1355497200, 1355500800, 1355504400, 1355508000, 1355511600, 
    1355515200, 1355518800, 1355522400, 1355526000, 1355529600, 1355533200, 
    1355536800, 1355540400, 1355544000, 1355547600, 1355551200, 1355554800, 
    1355558400, 1355562000, 1355565600, 1355569200, 1355572800, 1355576400, 
    1355580000, 1355583600, 1355587200, 1355590800, 1355594400, 1355598000, 
    1355601600, 1355605200, 1355608800, 1355612400, 1355616000, 1355619600, 
    1355623200, 1355626800, 1355630400, 1355634000, 1355637600, 1355641200, 
    1355644800, 1355648400, 1355652000, 1355655600, 1355659200, 1355662800, 
    1355666400, 1355670000, 1355673600, 1355677200, 1355680800, 1355684400, 
    1355688000, 1355691600, 1355695200, 1355698800, 1355702400, 1355706000, 
    1355709600, 1355713200, 1355716800, 1355720400, 1355724000, 1355727600, 
    1355731200, 1355734800, 1355738400, 1355742000, 1355745600, 1355749200, 
    1355752800, 1355756400, 1355760000, 1355763600, 1355767200, 1355770800, 
    1355774400, 1355778000, 1355781600, 1355785200, 1355788800, 1355792400, 
    1355796000, 1355799600, 1355803200, 1355806800, 1355810400, 1355814000, 
    1355817600, 1355821200, 1355824800, 1355828400, 1355832000, 1355835600, 
    1355839200, 1355842800, 1355846400, 1355850000, 1355853600, 1355857200, 
    1355860800, 1355864400, 1355868000, 1355871600, 1355875200, 1355878800, 
    1355882400, 1355886000, 1355889600, 1355893200, 1355896800, 1355900400, 
    1355904000, 1355907600, 1355911200, 1355914800, 1355918400, 1355922000, 
    1355925600, 1355929200, 1355932800, 1355936400, 1355940000, 1355943600, 
    1355947200, 1355950800, 1355954400, 1355958000, 1355961600, 1355965200, 
    1355968800, 1355972400, 1355976000, 1355979600, 1355983200, 1355986800, 
    1355990400, 1355994000, 1355997600, 1356001200, 1356004800, 1356008400, 
    1356012000, 1356015600, 1356019200, 1356022800, 1356026400, 1356030000, 
    1356033600, 1356037200, 1356040800, 1356044400, 1356048000, 1356051600, 
    1356055200, 1356058800, 1356062400, 1356066000, 1356069600, 1356073200, 
    1356076800, 1356080400, 1356084000, 1356087600, 1356091200, 1356094800, 
    1356098400, 1356102000, 1356105600, 1356109200, 1356112800, 1356116400, 
    1356120000, 1356123600, 1356127200, 1356130800, 1356134400, 1356138000, 
    1356141600, 1356145200, 1356148800, 1356152400, 1356156000, 1356159600, 
    1356163200, 1356166800, 1356170400, 1356174000, 1356177600, 1356181200, 
    1356184800, 1356188400, 1356192000, 1356195600, 1356199200, 1356202800, 
    1356206400, 1356210000, 1356213600, 1356217200, 1356220800, 1356224400, 
    1356228000, 1356231600, 1356235200, 1356238800, 1356242400, 1356246000, 
    1356249600, 1356253200, 1356256800, 1356260400, 1356264000, 1356267600, 
    1356271200, 1356274800, 1356278400, 1356282000, 1356285600, 1356289200, 
    1356292800, 1356296400, 1356300000, 1356303600, 1356307200, 1356310800, 
    1356314400, 1356318000, 1356321600, 1356325200, 1356328800, 1356332400, 
    1356336000, 1356339600, 1356343200, 1356346800, 1356350400, 1356354000, 
    1356357600, 1356361200, 1356364800, 1356368400, 1356372000, 1356375600, 
    1356379200, 1356382800, 1356386400, 1356390000, 1356393600, 1356397200, 
    1356400800, 1356404400, 1356408000, 1356411600, 1356415200, 1356418800, 
    1356422400, 1356426000, 1356429600, 1356433200, 1356436800, 1356440400, 
    1356444000, 1356447600, 1356451200, 1356454800, 1356458400, 1356462000, 
    1356465600, 1356469200, 1356472800, 1356476400, 1356480000, 1356483600, 
    1356487200, 1356490800, 1356494400, 1356498000, 1356501600, 1356505200, 
    1356508800, 1356512400, 1356516000, 1356519600, 1356523200, 1356526800, 
    1356530400, 1356534000, 1356537600, 1356541200, 1356544800, 1356548400, 
    1356552000, 1356555600, 1356559200, 1356562800, 1356566400, 1356570000, 
    1356573600, 1356577200, 1356580800, 1356584400, 1356588000, 1356591600, 
    1356595200, 1356598800, 1356602400, 1356606000, 1356609600, 1356613200, 
    1356616800, 1356620400, 1356624000, 1356627600, 1356631200, 1356634800, 
    1356638400, 1356642000, 1356645600, 1356649200, 1356652800, 1356656400, 
    1356660000, 1356663600, 1356667200, 1356670800, 1356674400, 1356678000, 
    1356681600, 1356685200, 1356688800, 1356692400, 1356696000, 1356699600, 
    1356703200, 1356706800, 1356710400, 1356714000, 1356717600, 1356721200, 
    1356724800, 1356728400, 1356732000, 1356735600, 1356739200, 1356742800, 
    1356746400, 1356750000, 1356753600, 1356757200, 1356760800, 1356764400, 
    1356768000, 1356771600, 1356775200, 1356778800, 1356782400, 1356786000, 
    1356789600, 1356793200, 1356796800, 1356800400, 1356804000, 1356807600, 
    1356811200, 1356814800, 1356818400, 1356822000, 1356825600, 1356829200, 
    1356832800, 1356836400, 1356840000, 1356843600, 1356847200, 1356850800, 
    1356854400, 1356858000, 1356861600, 1356865200, 1356868800, 1356872400, 
    1356876000, 1356879600, 1356883200, 1356886800, 1356890400, 1356894000, 
    1356897600, 1356901200, 1356904800, 1356908400, 1356912000, 1356915600, 
    1356919200, 1356922800, 1356926400, 1356930000, 1356933600, 1356937200, 
    1356940800, 1356944400, 1356948000, 1356951600, 1356955200, 1356958800, 
    1356962400, 1356966000, 1356969600, 1356973200, 1356976800, 1356980400, 
    1356984000, 1356987600, 1356991200, 1356994800, 1356998400, 1357002000, 
    1357005600, 1357009200, 1357012800, 1357016400, 1357020000, 1357023600, 
    1357027200, 1357030800, 1357034400, 1357038000, 1357041600, 1357045200, 
    1357048800, 1357052400, 1357056000, 1357059600, 1357063200, 1357066800, 
    1357070400, 1357074000, 1357077600, 1357081200, 1357084800, 1357088400, 
    1357092000, 1357095600, 1357099200, 1357102800, 1357106400, 1357110000, 
    1357113600, 1357117200, 1357120800, 1357124400, 1357128000, 1357131600, 
    1357135200, 1357138800, 1357142400, 1357146000, 1357149600, 1357153200, 
    1357156800, 1357160400, 1357164000, 1357167600, 1357171200, 1357174800, 
    1357178400, 1357182000, 1357185600, 1357189200, 1357192800, 1357196400, 
    1357200000, 1357203600, 1357207200, 1357210800, 1357214400, 1357218000, 
    1357221600, 1357225200, 1357228800, 1357232400, 1357236000, 1357239600, 
    1357243200, 1357246800, 1357250400, 1357254000, 1357257600, 1357261200, 
    1357264800, 1357268400, 1357272000, 1357275600, 1357279200, 1357282800, 
    1357286400, 1357290000, 1357293600, 1357297200, 1357300800, 1357304400, 
    1357308000, 1357311600, 1357315200, 1357318800, 1357322400, 1357326000, 
    1357329600, 1357333200, 1357336800, 1357340400, 1357344000, 1357347600, 
    1357351200, 1357354800, 1357358400, 1357362000, 1357365600, 1357369200, 
    1357372800, 1357376400, 1357380000, 1357383600, 1357387200, 1357390800, 
    1357394400, 1357398000, 1357401600, 1357405200, 1357408800, 1357412400, 
    1357416000, 1357419600, 1357423200, 1357426800, 1357430400, 1357434000, 
    1357437600, 1357441200, 1357444800, 1357448400, 1357452000, 1357455600, 
    1357459200, 1357462800, 1357466400, 1357470000, 1357473600, 1357477200, 
    1357480800, 1357484400, 1357488000, 1357491600, 1357495200, 1357498800, 
    1357502400, 1357506000, 1357509600, 1357513200, 1357516800, 1357520400, 
    1357524000, 1357527600, 1357531200, 1357534800, 1357538400, 1357542000, 
    1357545600, 1357549200, 1357552800, 1357556400, 1357560000, 1357563600, 
    1357567200, 1357570800, 1357574400, 1357578000, 1357581600, 1357585200, 
    1357588800, 1357592400, 1357596000, 1357599600, 1357603200, 1357606800, 
    1357610400, 1357614000, 1357617600, 1357621200, 1357624800, 1357628400, 
    1357632000, 1357635600, 1357639200, 1357642800, 1357646400, 1357650000, 
    1357653600, 1357657200, 1357660800, 1357664400, 1357668000, 1357671600, 
    1357675200, 1357678800, 1357682400, 1357686000, 1357689600, 1357693200, 
    1357696800, 1357700400, 1357704000, 1357707600, 1357711200, 1357714800, 
    1357718400, 1357722000, 1357725600, 1357729200, 1357732800, 1357736400, 
    1357740000, 1357743600, 1357747200, 1357750800, 1357754400, 1357758000, 
    1357761600, 1357765200, 1357768800, 1357772400, 1357776000, 1357779600, 
    1357783200, 1357786800, 1357790400, 1357794000, 1357797600, 1357801200, 
    1357804800, 1357808400, 1357812000, 1357815600, 1357819200, 1357822800, 
    1357826400, 1357830000, 1357833600, 1357837200, 1357840800, 1357844400, 
    1357848000, 1357851600, 1357855200, 1357858800, 1357862400, 1357866000, 
    1357869600, 1357873200, 1357876800, 1357880400, 1357884000, 1357887600, 
    1357891200, 1357894800, 1357898400, 1357902000, 1357905600, 1357909200, 
    1357912800, 1357916400, 1357920000, 1357923600, 1357927200, 1357930800, 
    1357934400, 1357938000, 1357941600, 1357945200, 1357948800, 1357952400, 
    1357956000, 1357959600, 1357963200, 1357966800, 1357970400, 1357974000, 
    1357977600, 1357981200, 1357984800, 1357988400, 1357992000, 1357995600, 
    1357999200, 1358002800, 1358006400, 1358010000, 1358013600, 1358017200, 
    1358020800, 1358024400, 1358028000, 1358031600, 1358035200, 1358038800, 
    1358042400, 1358046000, 1358049600, 1358053200, 1358056800, 1358060400, 
    1358064000, 1358067600, 1358071200, 1358074800, 1358078400, 1358082000, 
    1358085600, 1358089200, 1358092800, 1358096400, 1358100000, 1358103600, 
    1358107200, 1358110800, 1358114400, 1358118000, 1358121600, 1358125200, 
    1358128800, 1358132400, 1358136000, 1358139600, 1358143200, 1358146800, 
    1358150400, 1358154000, 1358157600, 1358161200, 1358164800, 1358168400, 
    1358172000, 1358175600, 1358179200, 1358182800, 1358186400, 1358190000, 
    1358193600, 1358197200, 1358200800, 1358204400, 1358208000, 1358211600, 
    1358215200, 1358218800, 1358222400, 1358226000, 1358229600, 1358233200, 
    1358236800, 1358240400, 1358244000, 1358247600, 1358251200, 1358254800, 
    1358258400, 1358262000, 1358265600, 1358269200, 1358272800, 1358276400, 
    1358280000, 1358283600, 1358287200, 1358290800, 1358294400, 1358298000, 
    1358301600, 1358305200, 1358308800, 1358312400, 1358316000, 1358319600, 
    1358323200, 1358326800, 1358330400, 1358334000, 1358337600, 1358341200, 
    1358344800, 1358348400, 1358352000, 1358355600, 1358359200, 1358362800, 
    1358366400, 1358370000, 1358373600, 1358377200, 1358380800, 1358384400, 
    1358388000, 1358391600, 1358395200, 1358398800, 1358402400, 1358406000, 
    1358409600, 1358413200, 1358416800, 1358420400, 1358424000, 1358427600, 
    1358431200, 1358434800, 1358438400, 1358442000, 1358445600, 1358449200, 
    1358452800, 1358456400, 1358460000, 1358463600, 1358467200, 1358470800, 
    1358474400, 1358478000, 1358481600, 1358485200, 1358488800, 1358492400, 
    1358496000, 1358499600, 1358503200, 1358506800, 1358510400, 1358514000, 
    1358517600, 1358521200, 1358524800, 1358528400, 1358532000, 1358535600, 
    1358539200, 1358542800, 1358546400, 1358550000, 1358553600, 1358557200, 
    1358560800, 1358564400, 1358568000, 1358571600, 1358575200, 1358578800, 
    1358582400, 1358586000, 1358589600, 1358593200, 1358596800, 1358600400, 
    1358604000, 1358607600, 1358611200, 1358614800, 1358618400, 1358622000, 
    1358625600, 1358629200, 1358632800, 1358636400, 1358640000, 1358643600, 
    1358647200, 1358650800, 1358654400, 1358658000, 1358661600, 1358665200, 
    1358668800, 1358672400, 1358676000, 1358679600, 1358683200, 1358686800, 
    1358690400, 1358694000, 1358697600, 1358701200, 1358704800, 1358708400, 
    1358712000, 1358715600, 1358719200, 1358722800, 1358726400, 1358730000, 
    1358733600, 1358737200, 1358740800, 1358744400, 1358748000, 1358751600, 
    1358755200, 1358758800, 1358762400, 1358766000, 1358769600, 1358773200, 
    1358776800, 1358780400, 1358784000, 1358787600, 1358791200, 1358794800, 
    1358798400, 1358802000, 1358805600, 1358809200, 1358812800, 1358816400, 
    1358820000, 1358823600, 1358827200, 1358830800, 1358834400, 1358838000, 
    1358841600, 1358845200, 1358848800, 1358852400, 1358856000, 1358859600, 
    1358863200, 1358866800, 1358870400, 1358874000, 1358877600, 1358881200, 
    1358884800, 1358888400, 1358892000, 1358895600, 1358899200, 1358902800, 
    1358906400, 1358910000, 1358913600, 1358917200, 1358920800, 1358924400, 
    1358928000, 1358931600, 1358935200, 1358938800, 1358942400, 1358946000, 
    1358949600, 1358953200, 1358956800, 1358960400, 1358964000, 1358967600, 
    1358971200, 1358974800, 1358978400, 1358982000, 1358985600, 1358989200, 
    1358992800, 1358996400, 1359000000, 1359003600, 1359007200, 1359010800, 
    1359014400, 1359018000, 1359021600, 1359025200, 1359028800, 1359032400, 
    1359036000, 1359039600, 1359043200, 1359046800, 1359050400, 1359054000, 
    1359057600, 1359061200, 1359064800, 1359068400, 1359072000, 1359075600, 
    1359079200, 1359082800, 1359086400, 1359090000, 1359093600, 1359097200, 
    1359100800, 1359104400, 1359108000, 1359111600, 1359115200, 1359118800, 
    1359122400, 1359126000, 1359129600, 1359133200, 1359136800, 1359140400, 
    1359144000, 1359147600, 1359151200, 1359154800, 1359158400, 1359162000, 
    1359165600, 1359169200, 1359172800, 1359176400, 1359180000, 1359183600, 
    1359187200, 1359190800, 1359194400, 1359198000, 1359201600, 1359205200, 
    1359208800, 1359212400, 1359216000, 1359219600, 1359223200, 1359226800, 
    1359230400, 1359234000, 1359237600, 1359241200, 1359244800, 1359248400, 
    1359252000, 1359255600, 1359259200, 1359262800, 1359266400, 1359270000, 
    1359273600, 1359277200, 1359280800, 1359284400, 1359288000, 1359291600, 
    1359295200, 1359298800, 1359302400, 1359306000, 1359309600, 1359313200, 
    1359316800, 1359320400, 1359324000, 1359327600, 1359331200, 1359334800, 
    1359338400, 1359342000, 1359345600, 1359349200, 1359352800, 1359356400, 
    1359360000, 1359363600, 1359367200, 1359370800, 1359374400, 1359378000, 
    1359381600, 1359385200, 1359388800, 1359392400, 1359396000, 1359399600, 
    1359403200, 1359406800, 1359410400, 1359414000, 1359417600, 1359421200, 
    1359424800, 1359428400, 1359432000, 1359435600, 1359439200, 1359442800, 
    1359446400, 1359450000, 1359453600, 1359457200, 1359460800, 1359464400, 
    1359468000, 1359471600, 1359475200, 1359478800, 1359482400, 1359486000, 
    1359489600, 1359493200, 1359496800, 1359500400, 1359504000, 1359507600, 
    1359511200, 1359514800, 1359518400, 1359522000, 1359525600, 1359529200, 
    1359532800, 1359536400, 1359540000, 1359543600, 1359547200, 1359550800, 
    1359554400, 1359558000, 1359561600, 1359565200, 1359568800, 1359572400, 
    1359576000, 1359579600, 1359583200, 1359586800, 1359590400, 1359594000, 
    1359597600, 1359601200, 1359604800, 1359608400, 1359612000, 1359615600, 
    1359619200, 1359622800, 1359626400, 1359630000, 1359633600, 1359637200, 
    1359640800, 1359644400, 1359648000, 1359651600, 1359655200, 1359658800, 
    1359662400, 1359666000, 1359669600, 1359673200, 1359676800, 1359680400, 
    1359684000, 1359687600, 1359691200, 1359694800, 1359698400, 1359702000, 
    1359705600, 1359709200, 1359712800, 1359716400, 1359720000, 1359723600, 
    1359727200, 1359730800, 1359734400, 1359738000, 1359741600, 1359745200, 
    1359748800, 1359752400, 1359756000, 1359759600, 1359763200, 1359766800, 
    1359770400, 1359774000, 1359777600, 1359781200, 1359784800, 1359788400, 
    1359792000, 1359795600, 1359799200, 1359802800, 1359806400, 1359810000, 
    1359813600, 1359817200, 1359820800, 1359824400, 1359828000, 1359831600, 
    1359835200, 1359838800, 1359842400, 1359846000, 1359849600, 1359853200, 
    1359856800, 1359860400, 1359864000, 1359867600, 1359871200, 1359874800, 
    1359878400, 1359882000, 1359885600, 1359889200, 1359892800, 1359896400, 
    1359900000, 1359903600, 1359907200, 1359910800, 1359914400, 1359918000, 
    1359921600, 1359925200, 1359928800, 1359932400, 1359936000, 1359939600, 
    1359943200, 1359946800, 1359950400, 1359954000, 1359957600, 1359961200, 
    1359964800, 1359968400, 1359972000, 1359975600, 1359979200, 1359982800, 
    1359986400, 1359990000, 1359993600, 1359997200, 1360000800, 1360004400, 
    1360008000, 1360011600, 1360015200, 1360018800, 1360022400, 1360026000, 
    1360029600, 1360033200, 1360036800, 1360040400, 1360044000, 1360047600, 
    1360051200, 1360054800, 1360058400, 1360062000, 1360065600, 1360069200, 
    1360072800, 1360076400, 1360080000, 1360083600, 1360087200, 1360090800, 
    1360094400, 1360098000, 1360101600, 1360105200, 1360108800, 1360112400, 
    1360116000, 1360119600, 1360123200, 1360126800, 1360130400, 1360134000, 
    1360137600, 1360141200, 1360144800, 1360148400, 1360152000, 1360155600, 
    1360159200, 1360162800, 1360166400, 1360170000, 1360173600, 1360177200, 
    1360180800, 1360184400, 1360188000, 1360191600, 1360195200, 1360198800, 
    1360202400, 1360206000, 1360209600, 1360213200, 1360216800, 1360220400, 
    1360224000, 1360227600, 1360231200, 1360234800, 1360238400, 1360242000, 
    1360245600, 1360249200, 1360252800, 1360256400, 1360260000, 1360263600, 
    1360267200, 1360270800, 1360274400, 1360278000, 1360281600, 1360285200, 
    1360288800, 1360292400, 1360296000, 1360299600, 1360303200, 1360306800, 
    1360310400, 1360314000, 1360317600, 1360321200, 1360324800, 1360328400, 
    1360332000, 1360335600, 1360339200, 1360342800, 1360346400, 1360350000, 
    1360353600, 1360357200, 1360360800, 1360364400, 1360368000, 1360371600, 
    1360375200, 1360378800, 1360382400, 1360386000, 1360389600, 1360393200, 
    1360396800, 1360400400, 1360404000, 1360407600, 1360411200, 1360414800, 
    1360418400, 1360422000, 1360425600, 1360429200, 1360432800, 1360436400, 
    1360440000, 1360443600, 1360447200, 1360450800, 1360454400, 1360458000, 
    1360461600, 1360465200, 1360468800, 1360472400, 1360476000, 1360479600, 
    1360483200, 1360486800, 1360490400, 1360494000, 1360497600, 1360501200, 
    1360504800, 1360508400, 1360512000, 1360515600, 1360519200, 1360522800, 
    1360526400, 1360530000, 1360533600, 1360537200, 1360540800, 1360544400, 
    1360548000, 1360551600, 1360555200, 1360558800, 1360562400, 1360566000, 
    1360569600, 1360573200, 1360576800, 1360580400, 1360584000, 1360587600, 
    1360591200, 1360594800, 1360598400, 1360602000, 1360605600, 1360609200, 
    1360612800, 1360616400, 1360620000, 1360623600, 1360627200, 1360630800, 
    1360634400, 1360638000, 1360641600, 1360645200, 1360648800, 1360652400, 
    1360656000, 1360659600, 1360663200, 1360666800, 1360670400, 1360674000, 
    1360677600, 1360681200, 1360684800, 1360688400, 1360692000, 1360695600, 
    1360699200, 1360702800, 1360706400, 1360710000, 1360713600, 1360717200, 
    1360720800, 1360724400, 1360728000, 1360731600, 1360735200, 1360738800, 
    1360742400, 1360746000, 1360749600, 1360753200, 1360756800, 1360760400, 
    1360764000, 1360767600, 1360771200, 1360774800, 1360778400, 1360782000, 
    1360785600, 1360789200, 1360792800, 1360796400, 1360800000, 1360803600, 
    1360807200, 1360810800, 1360814400, 1360818000, 1360821600, 1360825200, 
    1360828800, 1360832400, 1360836000, 1360839600, 1360843200, 1360846800, 
    1360850400, 1360854000, 1360857600, 1360861200, 1360864800, 1360868400, 
    1360872000, 1360875600, 1360879200, 1360882800, 1360886400, 1360890000, 
    1360893600, 1360897200, 1360900800, 1360904400, 1360908000, 1360911600, 
    1360915200, 1360918800, 1360922400, 1360926000, 1360929600, 1360933200, 
    1360936800, 1360940400, 1360944000, 1360947600, 1360951200, 1360954800, 
    1360958400, 1360962000, 1360965600, 1360969200, 1360972800, 1360976400, 
    1360980000, 1360983600, 1360987200, 1360990800, 1360994400, 1360998000, 
    1361001600, 1361005200, 1361008800, 1361012400, 1361016000, 1361019600, 
    1361023200, 1361026800, 1361030400, 1361034000, 1361037600, 1361041200, 
    1361044800, 1361048400, 1361052000, 1361055600, 1361059200, 1361062800, 
    1361066400, 1361070000, 1361073600, 1361077200, 1361080800, 1361084400, 
    1361088000, 1361091600, 1361095200, 1361098800, 1361102400, 1361106000, 
    1361109600, 1361113200, 1361116800, 1361120400, 1361124000, 1361127600, 
    1361131200, 1361134800, 1361138400, 1361142000, 1361145600, 1361149200, 
    1361152800, 1361156400, 1361160000, 1361163600, 1361167200, 1361170800, 
    1361174400, 1361178000, 1361181600, 1361185200, 1361188800, 1361192400, 
    1361196000, 1361199600, 1361203200, 1361206800, 1361210400, 1361214000, 
    1361217600, 1361221200, 1361224800, 1361228400, 1361232000, 1361235600, 
    1361239200, 1361242800, 1361246400, 1361250000, 1361253600, 1361257200, 
    1361260800, 1361264400, 1361268000, 1361271600, 1361275200, 1361278800, 
    1361282400, 1361286000, 1361289600, 1361293200, 1361296800, 1361300400, 
    1361304000, 1361307600, 1361311200, 1361314800, 1361318400, 1361322000, 
    1361325600, 1361329200, 1361332800, 1361336400, 1361340000, 1361343600, 
    1361347200, 1361350800, 1361354400, 1361358000, 1361361600, 1361365200, 
    1361368800, 1361372400, 1361376000, 1361379600, 1361383200, 1361386800, 
    1361390400, 1361394000, 1361397600, 1361401200, 1361404800, 1361408400, 
    1361412000, 1361415600, 1361419200, 1361422800, 1361426400, 1361430000, 
    1361433600, 1361437200, 1361440800, 1361444400, 1361448000, 1361451600, 
    1361455200, 1361458800, 1361462400, 1361466000, 1361469600, 1361473200, 
    1361476800, 1361480400, 1361484000, 1361487600, 1361491200, 1361494800, 
    1361498400, 1361502000, 1361505600, 1361509200, 1361512800, 1361516400, 
    1361520000, 1361523600, 1361527200, 1361530800, 1361534400, 1361538000, 
    1361541600, 1361545200, 1361548800, 1361552400, 1361556000, 1361559600, 
    1361563200, 1361566800, 1361570400, 1361574000, 1361577600, 1361581200, 
    1361584800, 1361588400, 1361592000, 1361595600, 1361599200, 1361602800, 
    1361606400, 1361610000, 1361613600, 1361617200, 1361620800, 1361624400, 
    1361628000, 1361631600, 1361635200, 1361638800, 1361642400, 1361646000, 
    1361649600, 1361653200, 1361656800, 1361660400, 1361664000, 1361667600, 
    1361671200, 1361674800, 1361678400, 1361682000, 1361685600, 1361689200, 
    1361692800, 1361696400, 1361700000, 1361703600, 1361707200, 1361710800, 
    1361714400, 1361718000, 1361721600, 1361725200, 1361728800, 1361732400, 
    1361736000, 1361739600, 1361743200, 1361746800, 1361750400, 1361754000, 
    1361757600, 1361761200, 1361764800, 1361768400, 1361772000, 1361775600, 
    1361779200, 1361782800, 1361786400, 1361790000, 1361793600, 1361797200, 
    1361800800, 1361804400, 1361808000, 1361811600, 1361815200, 1361818800, 
    1361822400, 1361826000, 1361829600, 1361833200, 1361836800, 1361840400, 
    1361844000, 1361847600, 1361851200, 1361854800, 1361858400, 1361862000, 
    1361865600, 1361869200, 1361872800, 1361876400, 1361880000, 1361883600, 
    1361887200, 1361890800, 1361894400, 1361898000, 1361901600, 1361905200, 
    1361908800, 1361912400, 1361916000, 1361919600, 1361923200, 1361926800, 
    1361930400, 1361934000, 1361937600, 1361941200, 1361944800, 1361948400, 
    1361952000, 1361955600, 1361959200, 1361962800, 1361966400, 1361970000, 
    1361973600, 1361977200, 1361980800, 1361984400, 1361988000, 1361991600, 
    1361995200, 1361998800, 1362002400, 1362006000, 1362009600, 1362013200, 
    1362016800, 1362020400, 1362024000, 1362027600, 1362031200, 1362034800, 
    1362038400, 1362042000, 1362045600, 1362049200, 1362052800, 1362056400, 
    1362060000, 1362063600, 1362067200, 1362070800, 1362074400, 1362078000, 
    1362081600, 1362085200, 1362088800, 1362092400, 1362096000, 1362099600, 
    1362103200, 1362106800, 1362110400, 1362114000, 1362117600, 1362121200, 
    1362124800, 1362128400, 1362132000, 1362135600, 1362139200, 1362142800, 
    1362146400, 1362150000, 1362153600, 1362157200, 1362160800, 1362164400, 
    1362168000, 1362171600, 1362175200, 1362178800, 1362182400, 1362186000, 
    1362189600, 1362193200, 1362196800, 1362200400, 1362204000, 1362207600, 
    1362211200, 1362214800, 1362218400, 1362222000, 1362225600, 1362229200, 
    1362232800, 1362236400, 1362240000, 1362243600, 1362247200, 1362250800, 
    1362254400, 1362258000, 1362261600, 1362265200, 1362268800, 1362272400, 
    1362276000, 1362279600, 1362283200, 1362286800, 1362290400, 1362294000, 
    1362297600, 1362301200, 1362304800, 1362308400, 1362312000, 1362315600, 
    1362319200, 1362322800, 1362326400, 1362330000, 1362333600, 1362337200, 
    1362340800, 1362344400, 1362348000, 1362351600, 1362355200, 1362358800, 
    1362362400, 1362366000, 1362369600, 1362373200, 1362376800, 1362380400, 
    1362384000, 1362387600, 1362391200, 1362394800, 1362398400, 1362402000, 
    1362405600, 1362409200, 1362412800, 1362416400, 1362420000, 1362423600, 
    1362427200, 1362430800, 1362434400, 1362438000, 1362441600, 1362445200, 
    1362448800, 1362452400, 1362456000, 1362459600, 1362463200, 1362466800, 
    1362470400, 1362474000, 1362477600, 1362481200, 1362484800, 1362488400, 
    1362492000, 1362495600, 1362499200, 1362502800, 1362506400, 1362510000, 
    1362513600, 1362517200, 1362520800, 1362524400, 1362528000, 1362531600, 
    1362535200, 1362538800, 1362542400, 1362546000, 1362549600, 1362553200, 
    1362556800, 1362560400, 1362564000, 1362567600, 1362571200, 1362574800, 
    1362578400, 1362582000, 1362585600, 1362589200, 1362592800, 1362596400, 
    1362600000, 1362603600, 1362607200, 1362610800, 1362614400, 1362618000, 
    1362621600, 1362625200, 1362628800, 1362632400, 1362636000, 1362639600, 
    1362643200, 1362646800, 1362650400, 1362654000, 1362657600, 1362661200, 
    1362664800, 1362668400, 1362672000, 1362675600, 1362679200, 1362682800, 
    1362686400, 1362690000, 1362693600, 1362697200, 1362700800, 1362704400, 
    1362708000, 1362711600, 1362715200, 1362718800, 1362722400, 1362726000, 
    1362729600, 1362733200, 1362736800, 1362740400, 1362744000, 1362747600, 
    1362751200, 1362754800, 1362758400, 1362762000, 1362765600, 1362769200, 
    1362772800, 1362776400, 1362780000, 1362783600, 1362787200, 1362790800, 
    1362794400, 1362798000, 1362801600, 1362805200, 1362808800, 1362812400, 
    1362816000, 1362819600, 1362823200, 1362826800, 1362830400, 1362834000, 
    1362837600, 1362841200, 1362844800, 1362848400, 1362852000, 1362855600, 
    1362859200, 1362862800, 1362866400, 1362870000, 1362873600, 1362877200, 
    1362880800, 1362884400, 1362888000, 1362891600, 1362895200, 1362898800, 
    1362902400, 1362906000, 1362909600, 1362913200, 1362916800, 1362920400, 
    1362924000, 1362927600, 1362931200, 1362934800, 1362938400, 1362942000, 
    1362945600, 1362949200, 1362952800, 1362956400, 1362960000, 1362963600, 
    1362967200, 1362970800, 1362974400, 1362978000, 1362981600, 1362985200, 
    1362988800, 1362992400, 1362996000, 1362999600, 1363003200, 1363006800, 
    1363010400, 1363014000, 1363017600, 1363021200, 1363024800, 1363028400, 
    1363032000, 1363035600, 1363039200, 1363042800, 1363046400, 1363050000, 
    1363053600, 1363057200, 1363060800, 1363064400, 1363068000, 1363071600, 
    1363075200, 1363078800, 1363082400, 1363086000, 1363089600, 1363093200, 
    1363096800, 1363100400, 1363104000, 1363107600, 1363111200, 1363114800, 
    1363118400, 1363122000, 1363125600, 1363129200, 1363132800, 1363136400, 
    1363140000, 1363143600, 1363147200, 1363150800, 1363154400, 1363158000, 
    1363161600, 1363165200, 1363168800, 1363172400, 1363176000, 1363179600, 
    1363183200, 1363186800, 1363190400, 1363194000, 1363197600, 1363201200, 
    1363204800, 1363208400, 1363212000, 1363215600, 1363219200, 1363222800, 
    1363226400, 1363230000, 1363233600, 1363237200, 1363240800, 1363244400, 
    1363248000, 1363251600, 1363255200, 1363258800, 1363262400, 1363266000, 
    1363269600, 1363273200, 1363276800, 1363280400, 1363284000, 1363287600, 
    1363291200, 1363294800, 1363298400, 1363302000, 1363305600, 1363309200, 
    1363312800, 1363316400, 1363320000, 1363323600, 1363327200, 1363330800, 
    1363334400, 1363338000, 1363341600, 1363345200, 1363348800, 1363352400, 
    1363356000, 1363359600, 1363363200, 1363366800, 1363370400, 1363374000, 
    1363377600, 1363381200, 1363384800, 1363388400, 1363392000, 1363395600, 
    1363399200, 1363402800, 1363406400, 1363410000, 1363413600, 1363417200, 
    1363420800, 1363424400, 1363428000, 1363431600, 1363435200, 1363438800, 
    1363442400, 1363446000, 1363449600, 1363453200, 1363456800, 1363460400, 
    1363464000, 1363467600, 1363471200, 1363474800, 1363478400, 1363482000, 
    1363485600, 1363489200, 1363492800, 1363496400, 1363500000, 1363503600, 
    1363507200, 1363510800, 1363514400, 1363518000, 1363521600, 1363525200, 
    1363528800, 1363532400, 1363536000, 1363539600, 1363543200, 1363546800, 
    1363550400, 1363554000, 1363557600, 1363561200, 1363564800, 1363568400, 
    1363572000, 1363575600, 1363579200, 1363582800, 1363586400, 1363590000, 
    1363593600, 1363597200, 1363600800, 1363604400, 1363608000, 1363611600, 
    1363615200, 1363618800, 1363622400, 1363626000, 1363629600, 1363633200, 
    1363636800, 1363640400, 1363644000, 1363647600, 1363651200, 1363654800, 
    1363658400, 1363662000, 1363665600, 1363669200, 1363672800, 1363676400, 
    1363680000, 1363683600, 1363687200, 1363690800, 1363694400, 1363698000, 
    1363701600, 1363705200, 1363708800, 1363712400, 1363716000, 1363719600, 
    1363723200, 1363726800, 1363730400, 1363734000, 1363737600, 1363741200, 
    1363744800, 1363748400, 1363752000, 1363755600, 1363759200, 1363762800, 
    1363766400, 1363770000, 1363773600, 1363777200, 1363780800, 1363784400, 
    1363788000, 1363791600, 1363795200, 1363798800, 1363802400, 1363806000, 
    1363809600, 1363813200, 1363816800, 1363820400, 1363824000, 1363827600, 
    1363831200, 1363834800, 1363838400, 1363842000, 1363845600, 1363849200, 
    1363852800, 1363856400, 1363860000, 1363863600, 1363867200, 1363870800, 
    1363874400, 1363878000, 1363881600, 1363885200, 1363888800, 1363892400, 
    1363896000, 1363899600, 1363903200, 1363906800, 1363910400, 1363914000, 
    1363917600, 1363921200, 1363924800, 1363928400, 1363932000, 1363935600, 
    1363939200, 1363942800, 1363946400, 1363950000, 1363953600, 1363957200, 
    1363960800, 1363964400, 1363968000, 1363971600, 1363975200, 1363978800, 
    1363982400, 1363986000, 1363989600, 1363993200, 1363996800, 1364000400, 
    1364004000, 1364007600, 1364011200, 1364014800, 1364018400, 1364022000, 
    1364025600, 1364029200, 1364032800, 1364036400, 1364040000, 1364043600, 
    1364047200, 1364050800, 1364054400, 1364058000, 1364061600, 1364065200, 
    1364068800, 1364072400, 1364076000, 1364079600, 1364083200, 1364086800, 
    1364090400, 1364094000, 1364097600, 1364101200, 1364104800, 1364108400, 
    1364112000, 1364115600, 1364119200, 1364122800, 1364126400, 1364130000, 
    1364133600, 1364137200, 1364140800, 1364144400, 1364148000, 1364151600, 
    1364155200, 1364158800, 1364162400, 1364166000, 1364169600, 1364173200, 
    1364176800, 1364180400, 1364184000, 1364187600, 1364191200, 1364194800, 
    1364198400, 1364202000, 1364205600, 1364209200, 1364212800, 1364216400, 
    1364220000, 1364223600, 1364227200, 1364230800, 1364234400, 1364238000, 
    1364241600, 1364245200, 1364248800, 1364252400, 1364256000, 1364259600, 
    1364263200, 1364266800, 1364270400, 1364274000, 1364277600, 1364281200, 
    1364284800, 1364288400, 1364292000, 1364295600, 1364299200, 1364302800, 
    1364306400, 1364310000, 1364313600, 1364317200, 1364320800, 1364324400, 
    1364328000, 1364331600, 1364335200, 1364338800, 1364342400, 1364346000, 
    1364349600, 1364353200, 1364356800, 1364360400, 1364364000, 1364367600, 
    1364371200, 1364374800, 1364378400, 1364382000, 1364385600, 1364389200, 
    1364392800, 1364396400, 1364400000, 1364403600, 1364407200, 1364410800, 
    1364414400, 1364418000, 1364421600, 1364425200, 1364428800, 1364432400, 
    1364436000, 1364439600, 1364443200, 1364446800, 1364450400, 1364454000, 
    1364457600, 1364461200, 1364464800, 1364468400, 1364472000, 1364475600, 
    1364479200, 1364482800, 1364486400, 1364490000, 1364493600, 1364497200, 
    1364500800, 1364504400, 1364508000, 1364511600, 1364515200, 1364518800, 
    1364522400, 1364526000, 1364529600, 1364533200, 1364536800, 1364540400, 
    1364544000, 1364547600, 1364551200, 1364554800, 1364558400, 1364562000, 
    1364565600, 1364569200, 1364572800, 1364576400, 1364580000, 1364583600, 
    1364587200, 1364590800, 1364594400, 1364598000, 1364601600, 1364605200, 
    1364608800, 1364612400, 1364616000, 1364619600, 1364623200, 1364626800, 
    1364630400, 1364634000, 1364637600, 1364641200, 1364644800, 1364648400, 
    1364652000, 1364655600, 1364659200, 1364662800, 1364666400, 1364670000, 
    1364673600, 1364677200, 1364680800, 1364684400, 1364688000, 1364691600, 
    1364695200, 1364698800, 1364702400, 1364706000, 1364709600, 1364713200, 
    1364716800, 1364720400, 1364724000, 1364727600, 1364731200, 1364734800, 
    1364738400, 1364742000, 1364745600, 1364749200, 1364752800, 1364756400, 
    1364760000, 1364763600, 1364767200, 1364770800, 1364774400, 1364778000, 
    1364781600, 1364785200, 1364788800, 1364792400, 1364796000, 1364799600, 
    1364803200, 1364806800, 1364810400, 1364814000, 1364817600, 1364821200, 
    1364824800, 1364828400, 1364832000, 1364835600, 1364839200, 1364842800, 
    1364846400, 1364850000, 1364853600, 1364857200, 1364860800, 1364864400, 
    1364868000, 1364871600, 1364875200, 1364878800, 1364882400, 1364886000, 
    1364889600, 1364893200, 1364896800, 1364900400, 1364904000, 1364907600, 
    1364911200, 1364914800, 1364918400, 1364922000, 1364925600, 1364929200, 
    1364932800, 1364936400, 1364940000, 1364943600, 1364947200, 1364950800, 
    1364954400, 1364958000, 1364961600, 1364965200, 1364968800, 1364972400, 
    1364976000, 1364979600, 1364983200, 1364986800, 1364990400, 1364994000, 
    1364997600, 1365001200, 1365004800, 1365008400, 1365012000, 1365015600, 
    1365019200, 1365022800, 1365026400, 1365030000, 1365033600, 1365037200, 
    1365040800, 1365044400, 1365048000, 1365051600, 1365055200, 1365058800, 
    1365062400, 1365066000, 1365069600, 1365073200, 1365076800, 1365080400, 
    1365084000, 1365087600, 1365091200, 1365094800, 1365098400, 1365102000, 
    1365105600, 1365109200, 1365112800, 1365116400, 1365120000, 1365123600, 
    1365127200, 1365130800, 1365134400, 1365138000, 1365141600, 1365145200, 
    1365148800, 1365152400, 1365156000, 1365159600, 1365163200, 1365166800, 
    1365170400, 1365174000, 1365177600, 1365181200, 1365184800, 1365188400, 
    1365192000, 1365195600, 1365199200, 1365202800, 1365206400, 1365210000, 
    1365213600, 1365217200, 1365220800, 1365224400, 1365228000, 1365231600, 
    1365235200, 1365238800, 1365242400, 1365246000, 1365249600, 1365253200, 
    1365256800, 1365260400, 1365264000, 1365267600, 1365271200, 1365274800, 
    1365278400, 1365282000, 1365285600, 1365289200, 1365292800, 1365296400, 
    1365300000, 1365303600, 1365307200, 1365310800, 1365314400, 1365318000, 
    1365321600, 1365325200, 1365328800, 1365332400, 1365336000, 1365339600, 
    1365343200, 1365346800, 1365350400, 1365354000, 1365357600, 1365361200, 
    1365364800, 1365368400, 1365372000, 1365375600, 1365379200, 1365382800, 
    1365386400, 1365390000, 1365393600, 1365397200, 1365400800, 1365404400, 
    1365408000, 1365411600, 1365415200, 1365418800, 1365422400, 1365426000, 
    1365429600, 1365433200, 1365436800, 1365440400, 1365444000, 1365447600, 
    1365451200, 1365454800, 1365458400, 1365462000, 1365465600, 1365469200, 
    1365472800, 1365476400, 1365480000, 1365483600, 1365487200, 1365490800, 
    1365494400, 1365498000, 1365501600, 1365505200, 1365508800, 1365512400, 
    1365516000, 1365519600, 1365523200, 1365526800, 1365530400, 1365534000, 
    1365537600, 1365541200, 1365544800, 1365548400, 1365552000, 1365555600, 
    1365559200, 1365562800, 1365566400, 1365570000, 1365573600, 1365577200, 
    1365580800, 1365584400, 1365588000, 1365591600, 1365595200, 1365598800, 
    1365602400, 1365606000, 1365609600, 1365613200, 1365616800, 1365620400, 
    1365624000, 1365627600, 1365631200, 1365634800, 1365638400, 1365642000, 
    1365645600, 1365649200, 1365652800, 1365656400, 1365660000, 1365663600, 
    1365667200, 1365670800, 1365674400, 1365678000, 1365681600, 1365685200, 
    1365688800, 1365692400, 1365696000, 1365699600, 1365703200, 1365706800, 
    1365710400, 1365714000, 1365717600, 1365721200, 1365724800, 1365728400, 
    1365732000, 1365735600, 1365739200, 1365742800, 1365746400, 1365750000, 
    1365753600, 1365757200, 1365760800, 1365764400, 1365768000, 1365771600, 
    1365775200, 1365778800, 1365782400, 1365786000, 1365789600, 1365793200, 
    1365796800, 1365800400, 1365804000, 1365807600, 1365811200, 1365814800, 
    1365818400, 1365822000, 1365825600, 1365829200, 1365832800, 1365836400, 
    1365840000, 1365843600, 1365847200, 1365850800, 1365854400, 1365858000, 
    1365861600, 1365865200, 1365868800, 1365872400, 1365876000, 1365879600, 
    1365883200, 1365886800, 1365890400, 1365894000, 1365897600, 1365901200, 
    1365904800, 1365908400, 1365912000, 1365915600, 1365919200, 1365922800, 
    1365926400, 1365930000, 1365933600, 1365937200, 1365940800, 1365944400, 
    1365948000, 1365951600, 1365955200, 1365958800, 1365962400, 1365966000, 
    1365969600, 1365973200, 1365976800, 1365980400, 1365984000, 1365987600, 
    1365991200, 1365994800, 1365998400, 1366002000, 1366005600, 1366009200, 
    1366012800, 1366016400, 1366020000, 1366023600, 1366027200, 1366030800, 
    1366034400, 1366038000, 1366041600, 1366045200, 1366048800, 1366052400, 
    1366056000, 1366059600, 1366063200, 1366066800, 1366070400, 1366074000, 
    1366077600, 1366081200, 1366084800, 1366088400, 1366092000, 1366095600, 
    1366099200, 1366102800, 1366106400, 1366110000, 1366113600, 1366117200, 
    1366120800, 1366124400, 1366128000, 1366131600, 1366135200, 1366138800, 
    1366142400, 1366146000, 1366149600, 1366153200, 1366156800, 1366160400, 
    1366164000, 1366167600, 1366171200, 1366174800, 1366178400, 1366182000, 
    1366185600, 1366189200, 1366192800, 1366196400, 1366200000, 1366203600, 
    1366207200, 1366210800, 1366214400, 1366218000, 1366221600, 1366225200, 
    1366228800, 1366232400, 1366236000, 1366239600, 1366243200, 1366246800, 
    1366250400, 1366254000, 1366257600, 1366261200, 1366264800, 1366268400, 
    1366272000, 1366275600, 1366279200, 1366282800, 1366286400, 1366290000, 
    1366293600, 1366297200, 1366300800, 1366304400, 1366308000, 1366311600, 
    1366315200, 1366318800, 1366322400, 1366326000, 1366329600, 1366333200, 
    1366336800, 1366340400, 1366344000, 1366347600, 1366351200, 1366354800, 
    1366358400, 1366362000, 1366365600, 1366369200, 1366372800, 1366376400, 
    1366380000, 1366383600, 1366387200, 1366390800, 1366394400, 1366398000, 
    1366401600, 1366405200, 1366408800, 1366412400, 1366416000, 1366419600, 
    1366423200, 1366426800, 1366430400, 1366434000, 1366437600, 1366441200, 
    1366444800, 1366448400, 1366452000, 1366455600, 1366459200, 1366462800, 
    1366466400, 1366470000, 1366473600, 1366477200, 1366480800, 1366484400, 
    1366488000, 1366491600, 1366495200, 1366498800, 1366502400, 1366506000, 
    1366509600, 1366513200, 1366516800, 1366520400, 1366524000, 1366527600, 
    1366531200, 1366534800, 1366538400, 1366542000, 1366545600, 1366549200, 
    1366552800, 1366556400, 1366560000, 1366563600, 1366567200, 1366570800, 
    1366574400, 1366578000, 1366581600, 1366585200, 1366588800, 1366592400, 
    1366596000, 1366599600, 1366603200, 1366606800, 1366610400, 1366614000, 
    1366617600, 1366621200, 1366624800, 1366628400, 1366632000, 1366635600, 
    1366639200, 1366642800, 1366646400, 1366650000, 1366653600, 1366657200, 
    1366660800, 1366664400, 1366668000, 1366671600, 1366675200, 1366678800, 
    1366682400, 1366686000, 1366689600, 1366693200, 1366696800, 1366700400, 
    1366704000, 1366707600, 1366711200, 1366714800, 1366718400, 1366722000, 
    1366725600, 1366729200, 1366732800, 1366736400, 1366740000, 1366743600, 
    1366747200, 1366750800, 1366754400, 1366758000, 1366761600, 1366765200, 
    1366768800, 1366772400, 1366776000, 1366779600, 1366783200, 1366786800, 
    1366790400, 1366794000, 1366797600, 1366801200, 1366804800, 1366808400, 
    1366812000, 1366815600, 1366819200, 1366822800, 1366826400, 1366830000, 
    1366833600, 1366837200, 1366840800, 1366844400, 1366848000, 1366851600, 
    1366855200, 1366858800, 1366862400, 1366866000, 1366869600, 1366873200, 
    1366876800, 1366880400, 1366884000, 1366887600, 1366891200, 1366894800, 
    1366898400, 1366902000, 1366905600, 1366909200, 1366912800, 1366916400, 
    1366920000, 1366923600, 1366927200, 1366930800, 1366934400, 1366938000, 
    1366941600, 1366945200, 1366948800, 1366952400, 1366956000, 1366959600, 
    1366963200, 1366966800, 1366970400, 1366974000, 1366977600, 1366981200, 
    1366984800, 1366988400, 1366992000, 1366995600, 1366999200, 1367002800, 
    1367006400, 1367010000, 1367013600, 1367017200, 1367020800, 1367024400, 
    1367028000, 1367031600, 1367035200, 1367038800, 1367042400, 1367046000, 
    1367049600, 1367053200, 1367056800, 1367060400, 1367064000, 1367067600, 
    1367071200, 1367074800, 1367078400, 1367082000, 1367085600, 1367089200, 
    1367092800, 1367096400, 1367100000, 1367103600, 1367107200, 1367110800, 
    1367114400, 1367118000, 1367121600, 1367125200, 1367128800, 1367132400, 
    1367136000, 1367139600, 1367143200, 1367146800, 1367150400, 1367154000, 
    1367157600, 1367161200, 1367164800, 1367168400, 1367172000, 1367175600, 
    1367179200, 1367182800, 1367186400, 1367190000, 1367193600, 1367197200, 
    1367200800, 1367204400, 1367208000, 1367211600, 1367215200, 1367218800, 
    1367222400, 1367226000, 1367229600, 1367233200, 1367236800, 1367240400, 
    1367244000, 1367247600, 1367251200, 1367254800, 1367258400, 1367262000, 
    1367265600, 1367269200, 1367272800, 1367276400, 1367280000, 1367283600, 
    1367287200, 1367290800, 1367294400, 1367298000, 1367301600, 1367305200, 
    1367308800, 1367312400, 1367316000, 1367319600, 1367323200, 1367326800, 
    1367330400, 1367334000, 1367337600, 1367341200, 1367344800, 1367348400, 
    1367352000, 1367355600, 1367359200, 1367362800, 1367366400, 1367370000, 
    1367373600, 1367377200, 1367380800, 1367384400, 1367388000, 1367391600, 
    1367395200, 1367398800, 1367402400, 1367406000, 1367409600, 1367413200, 
    1367416800, 1367420400, 1367424000, 1367427600, 1367431200, 1367434800, 
    1367438400, 1367442000, 1367445600, 1367449200, 1367452800, 1367456400, 
    1367460000, 1367463600, 1367467200, 1367470800, 1367474400, 1367478000, 
    1367481600, 1367485200, 1367488800, 1367492400, 1367496000, 1367499600, 
    1367503200, 1367506800, 1367510400, 1367514000, 1367517600, 1367521200, 
    1367524800, 1367528400, 1367532000, 1367535600, 1367539200, 1367542800, 
    1367546400, 1367550000, 1367553600, 1367557200, 1367560800, 1367564400, 
    1367568000, 1367571600, 1367575200, 1367578800, 1367582400, 1367586000, 
    1367589600, 1367593200, 1367596800, 1367600400, 1367604000, 1367607600, 
    1367611200, 1367614800, 1367618400, 1367622000, 1367625600, 1367629200, 
    1367632800, 1367636400, 1367640000, 1367643600, 1367647200, 1367650800, 
    1367654400, 1367658000, 1367661600, 1367665200, 1367668800, 1367672400, 
    1367676000, 1367679600, 1367683200, 1367686800, 1367690400, 1367694000, 
    1367697600, 1367701200, 1367704800, 1367708400, 1367712000, 1367715600, 
    1367719200, 1367722800, 1367726400, 1367730000, 1367733600, 1367737200, 
    1367740800, 1367744400, 1367748000, 1367751600, 1367755200, 1367758800, 
    1367762400, 1367766000, 1367769600, 1367773200, 1367776800, 1367780400, 
    1367784000, 1367787600, 1367791200, 1367794800, 1367798400, 1367802000, 
    1367805600, 1367809200, 1367812800, 1367816400, 1367820000, 1367823600, 
    1367827200, 1367830800, 1367834400, 1367838000, 1367841600, 1367845200, 
    1367848800, 1367852400, 1367856000, 1367859600, 1367863200, 1367866800, 
    1367870400, 1367874000, 1367877600, 1367881200, 1367884800, 1367888400, 
    1367892000, 1367895600, 1367899200, 1367902800, 1367906400, 1367910000, 
    1367913600, 1367917200, 1367920800, 1367924400, 1367928000, 1367931600, 
    1367935200, 1367938800, 1367942400, 1367946000, 1367949600, 1367953200, 
    1367956800, 1367960400, 1367964000, 1367967600, 1367971200, 1367974800, 
    1367978400, 1367982000, 1367985600, 1367989200, 1367992800, 1367996400, 
    1368000000, 1368003600, 1368007200, 1368010800, 1368014400, 1368018000, 
    1368021600, 1368025200, 1368028800, 1368032400, 1368036000, 1368039600, 
    1368043200, 1368046800, 1368050400, 1368054000, 1368057600, 1368061200, 
    1368064800, 1368068400, 1368072000, 1368075600, 1368079200, 1368082800, 
    1368086400, 1368090000, 1368093600, 1368097200, 1368100800, 1368104400, 
    1368108000, 1368111600, 1368115200, 1368118800, 1368122400, 1368126000, 
    1368129600, 1368133200, 1368136800, 1368140400, 1368144000, 1368147600, 
    1368151200, 1368154800, 1368158400, 1368162000, 1368165600, 1368169200, 
    1368172800, 1368176400, 1368180000, 1368183600, 1368187200, 1368190800, 
    1368194400, 1368198000, 1368201600, 1368205200, 1368208800, 1368212400, 
    1368216000, 1368219600, 1368223200, 1368226800, 1368230400, 1368234000, 
    1368237600, 1368241200, 1368244800, 1368248400, 1368252000, 1368255600, 
    1368259200, 1368262800, 1368266400, 1368270000, 1368273600, 1368277200, 
    1368280800, 1368284400, 1368288000, 1368291600, 1368295200, 1368298800, 
    1368302400, 1368306000, 1368309600, 1368313200, 1368316800, 1368320400, 
    1368324000, 1368327600, 1368331200, 1368334800, 1368338400, 1368342000, 
    1368345600, 1368349200, 1368352800, 1368356400, 1368360000, 1368363600, 
    1368367200, 1368370800, 1368374400, 1368378000, 1368381600, 1368385200, 
    1368388800, 1368392400, 1368396000, 1368399600, 1368403200, 1368406800, 
    1368410400, 1368414000, 1368417600, 1368421200, 1368424800, 1368428400, 
    1368432000, 1368435600, 1368439200, 1368442800, 1368446400, 1368450000, 
    1368453600, 1368457200, 1368460800, 1368464400, 1368468000, 1368471600, 
    1368475200, 1368478800, 1368482400, 1368486000, 1368489600, 1368493200, 
    1368496800, 1368500400, 1368504000, 1368507600, 1368511200, 1368514800, 
    1368518400, 1368522000, 1368525600, 1368529200, 1368532800, 1368536400, 
    1368540000, 1368543600, 1368547200, 1368550800, 1368554400, 1368558000, 
    1368561600, 1368565200, 1368568800, 1368572400, 1368576000, 1368579600, 
    1368583200, 1368586800, 1368590400, 1368594000, 1368597600, 1368601200, 
    1368604800, 1368608400, 1368612000, 1368615600, 1368619200, 1368622800, 
    1368626400, 1368630000, 1368633600, 1368637200, 1368640800, 1368644400, 
    1368648000, 1368651600, 1368655200, 1368658800, 1368662400, 1368666000, 
    1368669600, 1368673200, 1368676800, 1368680400, 1368684000, 1368687600, 
    1368691200, 1368694800, 1368698400, 1368702000, 1368705600, 1368709200, 
    1368712800, 1368716400, 1368720000, 1368723600, 1368727200, 1368730800, 
    1368734400, 1368738000, 1368741600, 1368745200, 1368748800, 1368752400, 
    1368756000, 1368759600, 1368763200, 1368766800, 1368770400, 1368774000, 
    1368777600, 1368781200, 1368784800, 1368788400, 1368792000, 1368795600, 
    1368799200, 1368802800, 1368806400, 1368810000, 1368813600, 1368817200, 
    1368820800, 1368824400, 1368828000, 1368831600, 1368835200, 1368838800, 
    1368842400, 1368846000, 1368849600, 1368853200, 1368856800, 1368860400, 
    1368864000, 1368867600, 1368871200, 1368874800, 1368878400, 1368882000, 
    1368885600, 1368889200, 1368892800, 1368896400, 1368900000, 1368903600, 
    1368907200, 1368910800, 1368914400, 1368918000, 1368921600, 1368925200, 
    1368928800, 1368932400, 1368936000, 1368939600, 1368943200, 1368946800, 
    1368950400, 1368954000, 1368957600, 1368961200, 1368964800, 1368968400, 
    1368972000, 1368975600, 1368979200, 1368982800, 1368986400, 1368990000, 
    1368993600, 1368997200, 1369000800, 1369004400, 1369008000, 1369011600, 
    1369015200, 1369018800, 1369022400, 1369026000, 1369029600, 1369033200, 
    1369036800, 1369040400, 1369044000, 1369047600, 1369051200, 1369054800, 
    1369058400, 1369062000, 1369065600, 1369069200, 1369072800, 1369076400, 
    1369080000, 1369083600, 1369087200, 1369090800, 1369094400, 1369098000, 
    1369101600, 1369105200, 1369108800, 1369112400, 1369116000, 1369119600, 
    1369123200, 1369126800, 1369130400, 1369134000, 1369137600, 1369141200, 
    1369144800, 1369148400, 1369152000, 1369155600, 1369159200, 1369162800, 
    1369166400, 1369170000, 1369173600, 1369177200, 1369180800, 1369184400, 
    1369188000, 1369191600, 1369195200, 1369198800, 1369202400, 1369206000, 
    1369209600, 1369213200, 1369216800, 1369220400, 1369224000, 1369227600, 
    1369231200, 1369234800, 1369238400, 1369242000, 1369245600, 1369249200, 
    1369252800, 1369256400, 1369260000, 1369263600, 1369267200, 1369270800, 
    1369274400, 1369278000, 1369281600, 1369285200, 1369288800, 1369292400, 
    1369296000, 1369299600, 1369303200, 1369306800, 1369310400, 1369314000, 
    1369317600, 1369321200, 1369324800, 1369328400, 1369332000, 1369335600, 
    1369339200, 1369342800, 1369346400, 1369350000, 1369353600, 1369357200, 
    1369360800, 1369364400, 1369368000, 1369371600, 1369375200, 1369378800, 
    1369382400, 1369386000, 1369389600, 1369393200, 1369396800, 1369400400, 
    1369404000, 1369407600, 1369411200, 1369414800, 1369418400, 1369422000, 
    1369425600, 1369429200, 1369432800, 1369436400, 1369440000, 1369443600, 
    1369447200, 1369450800, 1369454400, 1369458000, 1369461600, 1369465200, 
    1369468800, 1369472400, 1369476000, 1369479600, 1369483200, 1369486800, 
    1369490400, 1369494000, 1369497600, 1369501200, 1369504800, 1369508400, 
    1369512000, 1369515600, 1369519200, 1369522800, 1369526400, 1369530000, 
    1369533600, 1369537200, 1369540800, 1369544400, 1369548000, 1369551600, 
    1369555200, 1369558800, 1369562400, 1369566000, 1369569600, 1369573200, 
    1369576800, 1369580400, 1369584000, 1369587600, 1369591200, 1369594800, 
    1369598400, 1369602000, 1369605600, 1369609200, 1369612800, 1369616400, 
    1369620000, 1369623600, 1369627200, 1369630800, 1369634400, 1369638000, 
    1369641600, 1369645200, 1369648800, 1369652400, 1369656000, 1369659600, 
    1369663200, 1369666800, 1369670400, 1369674000, 1369677600, 1369681200, 
    1369684800, 1369688400, 1369692000, 1369695600, 1369699200, 1369702800, 
    1369706400, 1369710000, 1369713600, 1369717200, 1369720800, 1369724400, 
    1369728000, 1369731600, 1369735200, 1369738800, 1369742400, 1369746000, 
    1369749600, 1369753200, 1369756800, 1369760400, 1369764000, 1369767600, 
    1369771200, 1369774800, 1369778400, 1369782000, 1369785600, 1369789200, 
    1369792800, 1369796400, 1369800000, 1369803600, 1369807200, 1369810800, 
    1369814400, 1369818000, 1369821600, 1369825200, 1369828800, 1369832400, 
    1369836000, 1369839600, 1369843200, 1369846800, 1369850400, 1369854000, 
    1369857600, 1369861200, 1369864800, 1369868400, 1369872000, 1369875600, 
    1369879200, 1369882800, 1369886400, 1369890000, 1369893600, 1369897200, 
    1369900800, 1369904400, 1369908000, 1369911600, 1369915200, 1369918800, 
    1369922400, 1369926000, 1369929600, 1369933200, 1369936800, 1369940400, 
    1369944000, 1369947600, 1369951200, 1369954800, 1369958400, 1369962000, 
    1369965600, 1369969200, 1369972800, 1369976400, 1369980000, 1369983600, 
    1369987200, 1369990800, 1369994400, 1369998000, 1370001600, 1370005200, 
    1370008800, 1370012400, 1370016000, 1370019600, 1370023200, 1370026800, 
    1370030400, 1370034000, 1370037600, 1370041200, 1370044800, 1370048400, 
    1370052000, 1370055600, 1370059200, 1370062800, 1370066400, 1370070000, 
    1370073600, 1370077200, 1370080800, 1370084400, 1370088000, 1370091600, 
    1370095200, 1370098800, 1370102400, 1370106000, 1370109600, 1370113200, 
    1370116800, 1370120400, 1370124000, 1370127600, 1370131200, 1370134800, 
    1370138400, 1370142000, 1370145600, 1370149200, 1370152800, 1370156400, 
    1370160000, 1370163600, 1370167200, 1370170800, 1370174400, 1370178000, 
    1370181600, 1370185200, 1370188800, 1370192400, 1370196000, 1370199600, 
    1370203200, 1370206800, 1370210400, 1370214000, 1370217600, 1370221200, 
    1370224800, 1370228400, 1370232000, 1370235600, 1370239200, 1370242800, 
    1370246400, 1370250000, 1370253600, 1370257200, 1370260800, 1370264400, 
    1370268000, 1370271600, 1370275200, 1370278800, 1370282400, 1370286000, 
    1370289600, 1370293200, 1370296800, 1370300400, 1370304000, 1370307600, 
    1370311200, 1370314800, 1370318400, 1370322000, 1370325600, 1370329200, 
    1370332800, 1370336400, 1370340000, 1370343600, 1370347200, 1370350800, 
    1370354400, 1370358000, 1370361600, 1370365200, 1370368800, 1370372400, 
    1370376000, 1370379600, 1370383200, 1370386800, 1370390400, 1370394000, 
    1370397600, 1370401200, 1370404800, 1370408400, 1370412000, 1370415600, 
    1370419200, 1370422800, 1370426400, 1370430000, 1370433600, 1370437200, 
    1370440800, 1370444400, 1370448000, 1370451600, 1370455200, 1370458800, 
    1370462400, 1370466000, 1370469600, 1370473200, 1370476800, 1370480400, 
    1370484000, 1370487600, 1370491200, 1370494800, 1370498400, 1370502000, 
    1370505600, 1370509200, 1370512800, 1370516400, 1370520000, 1370523600, 
    1370527200, 1370530800, 1370534400, 1370538000, 1370541600, 1370545200, 
    1370548800, 1370552400, 1370556000, 1370559600, 1370563200, 1370566800, 
    1370570400, 1370574000, 1370577600, 1370581200, 1370584800, 1370588400, 
    1370592000, 1370595600, 1370599200, 1370602800, 1370606400, 1370610000, 
    1370613600, 1370617200, 1370620800, 1370624400, 1370628000, 1370631600, 
    1370635200, 1370638800, 1370642400, 1370646000, 1370649600, 1370653200, 
    1370656800, 1370660400, 1370664000, 1370667600, 1370671200, 1370674800, 
    1370678400, 1370682000, 1370685600, 1370689200, 1370692800, 1370696400, 
    1370700000, 1370703600, 1370707200, 1370710800, 1370714400, 1370718000, 
    1370721600, 1370725200, 1370728800, 1370732400, 1370736000, 1370739600, 
    1370743200, 1370746800, 1370750400, 1370754000, 1370757600, 1370761200, 
    1370764800, 1370768400, 1370772000, 1370775600, 1370779200, 1370782800, 
    1370786400, 1370790000, 1370793600, 1370797200, 1370800800, 1370804400, 
    1370808000, 1370811600, 1370815200, 1370818800, 1370822400, 1370826000, 
    1370829600, 1370833200, 1370836800, 1370840400, 1370844000, 1370847600, 
    1370851200, 1370854800, 1370858400, 1370862000, 1370865600, 1370869200, 
    1370872800, 1370876400, 1370880000, 1370883600, 1370887200, 1370890800, 
    1370894400, 1370898000, 1370901600, 1370905200, 1370908800, 1370912400, 
    1370916000, 1370919600, 1370923200, 1370926800, 1370930400, 1370934000, 
    1370937600, 1370941200, 1370944800, 1370948400, 1370952000, 1370955600, 
    1370959200, 1370962800, 1370966400, 1370970000, 1370973600, 1370977200, 
    1370980800, 1370984400, 1370988000, 1370991600, 1370995200, 1370998800, 
    1371002400, 1371006000, 1371009600, 1371013200, 1371016800, 1371020400, 
    1371024000, 1371027600, 1371031200, 1371034800, 1371038400, 1371042000, 
    1371045600, 1371049200, 1371052800, 1371056400, 1371060000, 1371063600, 
    1371067200, 1371070800, 1371074400, 1371078000, 1371081600, 1371085200, 
    1371088800, 1371092400, 1371096000, 1371099600, 1371103200, 1371106800, 
    1371110400, 1371114000, 1371117600, 1371121200, 1371124800, 1371128400, 
    1371132000, 1371135600, 1371139200, 1371142800, 1371146400, 1371150000, 
    1371153600, 1371157200, 1371160800, 1371164400, 1371168000, 1371171600, 
    1371175200, 1371178800, 1371182400, 1371186000, 1371189600, 1371193200, 
    1371196800, 1371200400, 1371204000, 1371207600, 1371211200, 1371214800, 
    1371218400, 1371222000, 1371225600, 1371229200, 1371232800, 1371236400, 
    1371240000, 1371243600, 1371247200, 1371250800, 1371254400, 1371258000, 
    1371261600, 1371265200, 1371268800, 1371272400, 1371276000, 1371279600, 
    1371283200, 1371286800, 1371290400, 1371294000, 1371297600, 1371301200, 
    1371304800, 1371308400, 1371312000, 1371315600, 1371319200, 1371322800, 
    1371326400, 1371330000, 1371333600, 1371337200, 1371340800, 1371344400, 
    1371348000, 1371351600, 1371355200, 1371358800, 1371362400, 1371366000, 
    1371369600, 1371373200, 1371376800, 1371380400, 1371384000, 1371387600, 
    1371391200, 1371394800, 1371398400, 1371402000, 1371405600, 1371409200, 
    1371412800, 1371416400, 1371420000, 1371423600, 1371427200, 1371430800, 
    1371434400, 1371438000, 1371441600, 1371445200, 1371448800, 1371452400, 
    1371456000, 1371459600, 1371463200, 1371466800, 1371470400, 1371474000, 
    1371477600, 1371481200, 1371484800, 1371488400, 1371492000, 1371495600, 
    1371499200, 1371502800, 1371506400, 1371510000, 1371513600, 1371517200, 
    1371520800, 1371524400, 1371528000, 1371531600, 1371535200, 1371538800, 
    1371542400, 1371546000, 1371549600, 1371553200, 1371556800, 1371560400, 
    1371564000, 1371567600, 1371571200, 1371574800, 1371578400, 1371582000, 
    1371585600, 1371589200, 1371592800, 1371596400, 1371600000, 1371603600, 
    1371607200, 1371610800, 1371614400, 1371618000, 1371621600, 1371625200, 
    1371628800, 1371632400, 1371636000, 1371639600, 1371643200, 1371646800, 
    1371650400, 1371654000, 1371657600, 1371661200, 1371664800, 1371668400, 
    1371672000, 1371675600, 1371679200, 1371682800, 1371686400, 1371690000, 
    1371693600, 1371697200, 1371700800, 1371704400, 1371708000, 1371711600, 
    1371715200, 1371718800, 1371722400, 1371726000, 1371729600, 1371733200, 
    1371736800, 1371740400, 1371744000, 1371747600, 1371751200, 1371754800, 
    1371758400, 1371762000, 1371765600, 1371769200, 1371772800, 1371776400, 
    1371780000, 1371783600, 1371787200, 1371790800, 1371794400, 1371798000, 
    1371801600, 1371805200, 1371808800, 1371812400, 1371816000, 1371819600, 
    1371823200, 1371826800, 1371830400, 1371834000, 1371837600, 1371841200, 
    1371844800, 1371848400, 1371852000, 1371855600, 1371859200, 1371862800, 
    1371866400, 1371870000, 1371873600, 1371877200, 1371880800, 1371884400, 
    1371888000, 1371891600, 1371895200, 1371898800, 1371902400, 1371906000, 
    1371909600, 1371913200, 1371916800, 1371920400, 1371924000, 1371927600, 
    1371931200, 1371934800, 1371938400, 1371942000, 1371945600, 1371949200, 
    1371952800, 1371956400, 1371960000, 1371963600, 1371967200, 1371970800, 
    1371974400, 1371978000, 1371981600, 1371985200, 1371988800, 1371992400, 
    1371996000, 1371999600, 1372003200, 1372006800, 1372010400, 1372014000, 
    1372017600, 1372021200, 1372024800, 1372028400, 1372032000, 1372035600, 
    1372039200, 1372042800, 1372046400, 1372050000, 1372053600, 1372057200, 
    1372060800, 1372064400, 1372068000, 1372071600, 1372075200, 1372078800, 
    1372082400, 1372086000, 1372089600, 1372093200, 1372096800, 1372100400, 
    1372104000, 1372107600, 1372111200, 1372114800, 1372118400, 1372122000, 
    1372125600, 1372129200, 1372132800, 1372136400, 1372140000, 1372143600, 
    1372147200, 1372150800, 1372154400, 1372158000, 1372161600, 1372165200, 
    1372168800, 1372172400, 1372176000, 1372179600, 1372183200, 1372186800, 
    1372190400, 1372194000, 1372197600, 1372201200, 1372204800, 1372208400, 
    1372212000, 1372215600, 1372219200, 1372222800, 1372226400, 1372230000, 
    1372233600, 1372237200, 1372240800, 1372244400, 1372248000, 1372251600, 
    1372255200, 1372258800, 1372262400, 1372266000, 1372269600, 1372273200, 
    1372276800, 1372280400, 1372284000, 1372287600, 1372291200, 1372294800, 
    1372298400, 1372302000, 1372305600, 1372309200, 1372312800, 1372316400, 
    1372320000, 1372323600, 1372327200, 1372330800, 1372334400, 1372338000, 
    1372341600, 1372345200, 1372348800, 1372352400, 1372356000, 1372359600, 
    1372363200, 1372366800, 1372370400, 1372374000, 1372377600, 1372381200, 
    1372384800, 1372388400, 1372392000, 1372395600, 1372399200, 1372402800, 
    1372406400, 1372410000, 1372413600, 1372417200, 1372420800, 1372424400, 
    1372428000, 1372431600, 1372435200, 1372438800, 1372442400, 1372446000, 
    1372449600, 1372453200, 1372456800, 1372460400, 1372464000, 1372467600, 
    1372471200, 1372474800, 1372478400, 1372482000, 1372485600, 1372489200, 
    1372492800, 1372496400, 1372500000, 1372503600, 1372507200, 1372510800, 
    1372514400, 1372518000, 1372521600, 1372525200, 1372528800, 1372532400, 
    1372536000, 1372539600, 1372543200, 1372546800, 1372550400, 1372554000, 
    1372557600, 1372561200, 1372564800, 1372568400, 1372572000, 1372575600, 
    1372579200, 1372582800, 1372586400, 1372590000, 1372593600, 1372597200, 
    1372600800, 1372604400, 1372608000, 1372611600, 1372615200, 1372618800, 
    1372622400, 1372626000, 1372629600, 1372633200, 1372636800, 1372640400, 
    1372644000, 1372647600, 1372651200, 1372654800, 1372658400, 1372662000, 
    1372665600, 1372669200, 1372672800, 1372676400, 1372680000, 1372683600, 
    1372687200, 1372690800, 1372694400, 1372698000, 1372701600, 1372705200, 
    1372708800, 1372712400, 1372716000, 1372719600, 1372723200, 1372726800, 
    1372730400, 1372734000, 1372737600, 1372741200, 1372744800, 1372748400, 
    1372752000, 1372755600, 1372759200, 1372762800, 1372766400, 1372770000, 
    1372773600, 1372777200, 1372780800, 1372784400, 1372788000, 1372791600, 
    1372795200, 1372798800, 1372802400, 1372806000, 1372809600, 1372813200, 
    1372816800, 1372820400, 1372824000, 1372827600, 1372831200, 1372834800, 
    1372838400, 1372842000, 1372845600, 1372849200, 1372852800, 1372856400, 
    1372860000, 1372863600, 1372867200, 1372870800, 1372874400, 1372878000, 
    1372881600, 1372885200, 1372888800, 1372892400, 1372896000, 1372899600, 
    1372903200, 1372906800, 1372910400, 1372914000, 1372917600, 1372921200, 
    1372924800, 1372928400, 1372932000, 1372935600, 1372939200, 1372942800, 
    1372946400, 1372950000, 1372953600, 1372957200, 1372960800, 1372964400, 
    1372968000, 1372971600, 1372975200, 1372978800, 1372982400, 1372986000, 
    1372989600, 1372993200, 1372996800, 1373000400, 1373004000, 1373007600, 
    1373011200, 1373014800, 1373018400, 1373022000, 1373025600, 1373029200, 
    1373032800, 1373036400, 1373040000, 1373043600, 1373047200, 1373050800, 
    1373054400, 1373058000, 1373061600, 1373065200, 1373068800, 1373072400, 
    1373076000, 1373079600, 1373083200, 1373086800, 1373090400, 1373094000, 
    1373097600, 1373101200, 1373104800, 1373108400, 1373112000, 1373115600, 
    1373119200, 1373122800, 1373126400, 1373130000, 1373133600, 1373137200, 
    1373140800, 1373144400, 1373148000, 1373151600, 1373155200, 1373158800, 
    1373162400, 1373166000, 1373169600, 1373173200, 1373176800, 1373180400, 
    1373184000, 1373187600, 1373191200, 1373194800, 1373198400, 1373202000, 
    1373205600, 1373209200, 1373212800, 1373216400, 1373220000, 1373223600, 
    1373227200, 1373230800, 1373234400, 1373238000, 1373241600, 1373245200, 
    1373248800, 1373252400, 1373256000, 1373259600, 1373263200, 1373266800, 
    1373270400, 1373274000, 1373277600, 1373281200, 1373284800, 1373288400, 
    1373292000, 1373295600, 1373299200, 1373302800, 1373306400, 1373310000, 
    1373313600, 1373317200, 1373320800, 1373324400, 1373328000, 1373331600, 
    1373335200, 1373338800, 1373342400, 1373346000, 1373349600, 1373353200, 
    1373356800, 1373360400, 1373364000, 1373367600, 1373371200, 1373374800, 
    1373378400, 1373382000, 1373385600, 1373389200, 1373392800, 1373396400, 
    1373400000, 1373403600, 1373407200, 1373410800, 1373414400, 1373418000, 
    1373421600, 1373425200, 1373428800, 1373432400, 1373436000, 1373439600, 
    1373443200, 1373446800, 1373450400, 1373454000, 1373457600, 1373461200, 
    1373464800, 1373468400, 1373472000, 1373475600, 1373479200, 1373482800, 
    1373486400, 1373490000, 1373493600, 1373497200, 1373500800, 1373504400, 
    1373508000, 1373511600, 1373515200, 1373518800, 1373522400, 1373526000, 
    1373529600, 1373533200, 1373536800, 1373540400, 1373544000, 1373547600, 
    1373551200, 1373554800, 1373558400, 1373562000, 1373565600, 1373569200, 
    1373572800, 1373576400, 1373580000, 1373583600, 1373587200, 1373590800, 
    1373594400, 1373598000, 1373601600, 1373605200, 1373608800, 1373612400, 
    1373616000, 1373619600, 1373623200, 1373626800, 1373630400, 1373634000, 
    1373637600, 1373641200, 1373644800, 1373648400, 1373652000, 1373655600, 
    1373659200, 1373662800, 1373666400, 1373670000, 1373673600, 1373677200, 
    1373680800, 1373684400, 1373688000, 1373691600, 1373695200, 1373698800, 
    1373702400, 1373706000, 1373709600, 1373713200, 1373716800, 1373720400, 
    1373724000, 1373727600, 1373731200, 1373734800, 1373738400, 1373742000, 
    1373745600, 1373749200, 1373752800, 1373756400, 1373760000, 1373763600, 
    1373767200, 1373770800, 1373774400, 1373778000, 1373781600, 1373785200, 
    1373788800, 1373792400, 1373796000, 1373799600, 1373803200, 1373806800, 
    1373810400, 1373814000, 1373817600, 1373821200, 1373824800, 1373828400, 
    1373832000, 1373835600, 1373839200, 1373842800, 1373846400, 1373850000, 
    1373853600, 1373857200, 1373860800, 1373864400, 1373868000, 1373871600, 
    1373875200, 1373878800, 1373882400, 1373886000, 1373889600, 1373893200, 
    1373896800, 1373900400, 1373904000, 1373907600, 1373911200, 1373914800, 
    1373918400, 1373922000, 1373925600, 1373929200, 1373932800, 1373936400, 
    1373940000, 1373943600, 1373947200, 1373950800, 1373954400, 1373958000, 
    1373961600, 1373965200, 1373968800, 1373972400, 1373976000, 1373979600, 
    1373983200, 1373986800, 1373990400, 1373994000, 1373997600, 1374001200, 
    1374004800, 1374008400, 1374012000, 1374015600, 1374019200, 1374022800, 
    1374026400, 1374030000, 1374033600, 1374037200, 1374040800, 1374044400, 
    1374048000, 1374051600, 1374055200, 1374058800, 1374062400, 1374066000, 
    1374069600, 1374073200, 1374076800, 1374080400, 1374084000, 1374087600, 
    1374091200, 1374094800, 1374098400, 1374102000, 1374105600, 1374109200, 
    1374112800, 1374116400, 1374120000, 1374123600, 1374127200, 1374130800, 
    1374134400, 1374138000, 1374141600, 1374145200, 1374148800, 1374152400, 
    1374156000, 1374159600, 1374163200, 1374166800, 1374170400, 1374174000, 
    1374177600, 1374181200, 1374184800, 1374188400, 1374192000, 1374195600, 
    1374199200, 1374202800, 1374206400, 1374210000, 1374213600, 1374217200, 
    1374220800, 1374224400, 1374228000, 1374231600, 1374235200, 1374238800, 
    1374242400, 1374246000, 1374249600, 1374253200, 1374256800, 1374260400, 
    1374264000, 1374267600, 1374271200, 1374274800, 1374278400, 1374282000, 
    1374285600, 1374289200, 1374292800, 1374296400, 1374300000, 1374303600, 
    1374307200, 1374310800, 1374314400, 1374318000, 1374321600, 1374325200, 
    1374328800, 1374332400, 1374336000, 1374339600, 1374343200, 1374346800, 
    1374350400, 1374354000, 1374357600, 1374361200, 1374364800, 1374368400, 
    1374372000, 1374375600, 1374379200, 1374382800, 1374386400, 1374390000, 
    1374393600, 1374397200, 1374400800, 1374404400, 1374408000, 1374411600, 
    1374415200, 1374418800, 1374422400, 1374426000, 1374429600, 1374433200, 
    1374436800, 1374440400, 1374444000, 1374447600, 1374451200, 1374454800, 
    1374458400, 1374462000, 1374465600, 1374469200, 1374472800, 1374476400, 
    1374480000, 1374483600, 1374487200, 1374490800, 1374494400, 1374498000, 
    1374501600, 1374505200, 1374508800, 1374512400, 1374516000, 1374519600, 
    1374523200, 1374526800, 1374530400, 1374534000, 1374537600, 1374541200, 
    1374544800, 1374548400, 1374552000, 1374555600, 1374559200, 1374562800, 
    1374566400, 1374570000, 1374573600, 1374577200, 1374580800, 1374584400, 
    1374588000, 1374591600, 1374595200, 1374598800, 1374602400, 1374606000, 
    1374609600, 1374613200, 1374616800, 1374620400, 1374624000, 1374627600, 
    1374631200, 1374634800, 1374638400, 1374642000, 1374645600, 1374649200, 
    1374652800, 1374656400, 1374660000, 1374663600, 1374667200, 1374670800, 
    1374674400, 1374678000, 1374681600, 1374685200, 1374688800, 1374692400, 
    1374696000, 1374699600, 1374703200, 1374706800, 1374710400, 1374714000, 
    1374717600, 1374721200, 1374724800, 1374728400, 1374732000, 1374735600, 
    1374739200, 1374742800, 1374746400, 1374750000, 1374753600, 1374757200, 
    1374760800, 1374764400, 1374768000, 1374771600, 1374775200, 1374778800, 
    1374782400, 1374786000, 1374789600, 1374793200, 1374796800, 1374800400, 
    1374804000, 1374807600, 1374811200, 1374814800, 1374818400, 1374822000, 
    1374825600, 1374829200, 1374832800, 1374836400, 1374840000, 1374843600, 
    1374847200, 1374850800, 1374854400, 1374858000, 1374861600, 1374865200, 
    1374868800, 1374872400, 1374876000, 1374879600, 1374883200, 1374886800, 
    1374890400, 1374894000, 1374897600, 1374901200, 1374904800, 1374908400, 
    1374912000, 1374915600, 1374919200, 1374922800, 1374926400, 1374930000, 
    1374933600, 1374937200, 1374940800, 1374944400, 1374948000, 1374951600, 
    1374955200, 1374958800, 1374962400, 1374966000, 1374969600, 1374973200, 
    1374976800, 1374980400, 1374984000, 1374987600, 1374991200, 1374994800, 
    1374998400, 1375002000, 1375005600, 1375009200, 1375012800, 1375016400, 
    1375020000, 1375023600, 1375027200, 1375030800, 1375034400, 1375038000, 
    1375041600, 1375045200, 1375048800, 1375052400, 1375056000, 1375059600, 
    1375063200, 1375066800, 1375070400, 1375074000, 1375077600, 1375081200, 
    1375084800, 1375088400, 1375092000, 1375095600, 1375099200, 1375102800, 
    1375106400, 1375110000, 1375113600, 1375117200, 1375120800, 1375124400, 
    1375128000, 1375131600, 1375135200, 1375138800, 1375142400, 1375146000, 
    1375149600, 1375153200, 1375156800, 1375160400, 1375164000, 1375167600, 
    1375171200, 1375174800, 1375178400, 1375182000, 1375185600, 1375189200, 
    1375192800, 1375196400, 1375200000, 1375203600, 1375207200, 1375210800, 
    1375214400, 1375218000, 1375221600, 1375225200, 1375228800, 1375232400, 
    1375236000, 1375239600, 1375243200, 1375246800, 1375250400, 1375254000, 
    1375257600, 1375261200, 1375264800, 1375268400, 1375272000, 1375275600, 
    1375279200, 1375282800, 1375286400, 1375290000, 1375293600, 1375297200, 
    1375300800, 1375304400, 1375308000, 1375311600, 1375315200, 1375318800, 
    1375322400, 1375326000, 1375329600, 1375333200, 1375336800, 1375340400, 
    1375344000, 1375347600, 1375351200, 1375354800, 1375358400, 1375362000, 
    1375365600, 1375369200, 1375372800, 1375376400, 1375380000, 1375383600, 
    1375387200, 1375390800, 1375394400, 1375398000, 1375401600, 1375405200, 
    1375408800, 1375412400, 1375416000, 1375419600, 1375423200, 1375426800, 
    1375430400, 1375434000, 1375437600, 1375441200, 1375444800, 1375448400, 
    1375452000, 1375455600, 1375459200, 1375462800, 1375466400, 1375470000, 
    1375473600, 1375477200, 1375480800, 1375484400, 1375488000, 1375491600, 
    1375495200, 1375498800, 1375502400, 1375506000, 1375509600, 1375513200, 
    1375516800, 1375520400, 1375524000, 1375527600, 1375531200, 1375534800, 
    1375538400, 1375542000, 1375545600, 1375549200, 1375552800, 1375556400, 
    1375560000, 1375563600, 1375567200, 1375570800, 1375574400, 1375578000, 
    1375581600, 1375585200, 1375588800, 1375592400, 1375596000, 1375599600, 
    1375603200, 1375606800, 1375610400, 1375614000, 1375617600, 1375621200, 
    1375624800, 1375628400, 1375632000, 1375635600, 1375639200, 1375642800, 
    1375646400, 1375650000, 1375653600, 1375657200, 1375660800, 1375664400, 
    1375668000, 1375671600, 1375675200, 1375678800, 1375682400, 1375686000, 
    1375689600, 1375693200, 1375696800, 1375700400, 1375704000, 1375707600, 
    1375711200, 1375714800, 1375718400, 1375722000, 1375725600, 1375729200, 
    1375732800, 1375736400, 1375740000, 1375743600, 1375747200, 1375750800, 
    1375754400, 1375758000, 1375761600, 1375765200, 1375768800, 1375772400, 
    1375776000, 1375779600, 1375783200, 1375786800, 1375790400, 1375794000, 
    1375797600, 1375801200, 1375804800, 1375808400, 1375812000, 1375815600, 
    1375819200, 1375822800, 1375826400, 1375830000, 1375833600, 1375837200, 
    1375840800, 1375844400, 1375848000, 1375851600, 1375855200, 1375858800, 
    1375862400, 1375866000, 1375869600, 1375873200, 1375876800, 1375880400, 
    1375884000, 1375887600, 1375891200, 1375894800, 1375898400, 1375902000, 
    1375905600, 1375909200, 1375912800, 1375916400, 1375920000, 1375923600, 
    1375927200, 1375930800, 1375934400, 1375938000, 1375941600, 1375945200, 
    1375948800, 1375952400, 1375956000, 1375959600, 1375963200, 1375966800, 
    1375970400, 1375974000, 1375977600, 1375981200, 1375984800, 1375988400, 
    1375992000, 1375995600, 1375999200, 1376002800, 1376006400, 1376010000, 
    1376013600, 1376017200, 1376020800, 1376024400, 1376028000, 1376031600, 
    1376035200, 1376038800, 1376042400, 1376046000, 1376049600, 1376053200, 
    1376056800, 1376060400, 1376064000, 1376067600, 1376071200, 1376074800, 
    1376078400, 1376082000, 1376085600, 1376089200, 1376092800, 1376096400, 
    1376100000, 1376103600, 1376107200, 1376110800, 1376114400, 1376118000, 
    1376121600, 1376125200, 1376128800, 1376132400, 1376136000, 1376139600, 
    1376143200, 1376146800, 1376150400, 1376154000, 1376157600, 1376161200, 
    1376164800, 1376168400, 1376172000, 1376175600, 1376179200, 1376182800, 
    1376186400, 1376190000, 1376193600, 1376197200, 1376200800, 1376204400, 
    1376208000, 1376211600, 1376215200, 1376218800, 1376222400, 1376226000, 
    1376229600, 1376233200, 1376236800, 1376240400, 1376244000, 1376247600, 
    1376251200, 1376254800, 1376258400, 1376262000, 1376265600, 1376269200, 
    1376272800, 1376276400, 1376280000, 1376283600, 1376287200, 1376290800, 
    1376294400, 1376298000, 1376301600, 1376305200, 1376308800, 1376312400, 
    1376316000, 1376319600, 1376323200, 1376326800, 1376330400, 1376334000, 
    1376337600, 1376341200, 1376344800, 1376348400, 1376352000, 1376355600, 
    1376359200, 1376362800, 1376366400, 1376370000, 1376373600, 1376377200, 
    1376380800, 1376384400, 1376388000, 1376391600, 1376395200, 1376398800, 
    1376402400, 1376406000, 1376409600, 1376413200, 1376416800, 1376420400, 
    1376424000, 1376427600, 1376431200, 1376434800, 1376438400, 1376442000, 
    1376445600, 1376449200, 1376452800, 1376456400, 1376460000, 1376463600, 
    1376467200, 1376470800, 1376474400, 1376478000, 1376481600, 1376485200, 
    1376488800, 1376492400, 1376496000, 1376499600, 1376503200, 1376506800, 
    1376510400, 1376514000, 1376517600, 1376521200, 1376524800, 1376528400, 
    1376532000, 1376535600, 1376539200, 1376542800, 1376546400, 1376550000, 
    1376553600, 1376557200, 1376560800, 1376564400, 1376568000, 1376571600, 
    1376575200, 1376578800, 1376582400, 1376586000, 1376589600, 1376593200, 
    1376596800, 1376600400, 1376604000, 1376607600, 1376611200, 1376614800, 
    1376618400, 1376622000, 1376625600, 1376629200, 1376632800, 1376636400, 
    1376640000, 1376643600, 1376647200, 1376650800, 1376654400, 1376658000, 
    1376661600, 1376665200, 1376668800, 1376672400, 1376676000, 1376679600, 
    1376683200, 1376686800, 1376690400, 1376694000, 1376697600, 1376701200, 
    1376704800, 1376708400, 1376712000, 1376715600, 1376719200, 1376722800, 
    1376726400, 1376730000, 1376733600, 1376737200, 1376740800, 1376744400, 
    1376748000, 1376751600, 1376755200, 1376758800, 1376762400, 1376766000, 
    1376769600, 1376773200, 1376776800, 1376780400, 1376784000, 1376787600, 
    1376791200, 1376794800, 1376798400, 1376802000, 1376805600, 1376809200, 
    1376812800, 1376816400, 1376820000, 1376823600, 1376827200, 1376830800, 
    1376834400, 1376838000, 1376841600, 1376845200, 1376848800, 1376852400, 
    1376856000, 1376859600, 1376863200, 1376866800, 1376870400, 1376874000, 
    1376877600, 1376881200, 1376884800, 1376888400, 1376892000, 1376895600, 
    1376899200, 1376902800, 1376906400, 1376910000, 1376913600, 1376917200, 
    1376920800, 1376924400, 1376928000, 1376931600, 1376935200, 1376938800, 
    1376942400, 1376946000, 1376949600, 1376953200, 1376956800, 1376960400, 
    1376964000, 1376967600, 1376971200, 1376974800, 1376978400, 1376982000, 
    1376985600, 1376989200, 1376992800, 1376996400, 1377000000, 1377003600, 
    1377007200, 1377010800, 1377014400, 1377018000, 1377021600, 1377025200, 
    1377028800, 1377032400, 1377036000, 1377039600, 1377043200, 1377046800, 
    1377050400, 1377054000, 1377057600, 1377061200, 1377064800, 1377068400, 
    1377072000, 1377075600, 1377079200, 1377082800, 1377086400, 1377090000, 
    1377093600, 1377097200, 1377100800, 1377104400, 1377108000, 1377111600, 
    1377115200, 1377118800, 1377122400, 1377126000, 1377129600, 1377133200, 
    1377136800, 1377140400, 1377144000, 1377147600, 1377151200, 1377154800, 
    1377158400, 1377162000, 1377165600, 1377169200, 1377172800, 1377176400, 
    1377180000, 1377183600, 1377187200, 1377190800, 1377194400, 1377198000, 
    1377201600, 1377205200, 1377208800, 1377212400, 1377216000, 1377219600, 
    1377223200, 1377226800, 1377230400, 1377234000, 1377237600, 1377241200, 
    1377244800, 1377248400, 1377252000, 1377255600, 1377259200, 1377262800, 
    1377266400, 1377270000, 1377273600, 1377277200, 1377280800, 1377284400, 
    1377288000, 1377291600, 1377295200, 1377298800, 1377302400, 1377306000, 
    1377309600, 1377313200, 1377316800, 1377320400, 1377324000, 1377327600, 
    1377331200, 1377334800, 1377338400, 1377342000, 1377345600, 1377349200, 
    1377352800, 1377356400, 1377360000, 1377363600, 1377367200, 1377370800, 
    1377374400, 1377378000, 1377381600, 1377385200, 1377388800, 1377392400, 
    1377396000, 1377399600, 1377403200, 1377406800, 1377410400, 1377414000, 
    1377417600, 1377421200, 1377424800, 1377428400, 1377432000, 1377435600, 
    1377439200, 1377442800, 1377446400, 1377450000, 1377453600, 1377457200, 
    1377460800, 1377464400, 1377468000, 1377471600, 1377475200, 1377478800, 
    1377482400, 1377486000, 1377489600, 1377493200, 1377496800, 1377500400, 
    1377504000, 1377507600, 1377511200, 1377514800, 1377518400, 1377522000, 
    1377525600, 1377529200, 1377532800, 1377536400, 1377540000, 1377543600, 
    1377547200, 1377550800, 1377554400, 1377558000, 1377561600, 1377565200, 
    1377568800, 1377572400, 1377576000, 1377579600, 1377583200, 1377586800, 
    1377590400, 1377594000, 1377597600, 1377601200, 1377604800, 1377608400, 
    1377612000, 1377615600, 1377619200, 1377622800, 1377626400, 1377630000, 
    1377633600, 1377637200, 1377640800, 1377644400, 1377648000, 1377651600, 
    1377655200, 1377658800, 1377662400, 1377666000, 1377669600, 1377673200, 
    1377676800, 1377680400, 1377684000, 1377687600, 1377691200, 1377694800, 
    1377698400, 1377702000, 1377705600, 1377709200, 1377712800, 1377716400, 
    1377720000, 1377723600, 1377727200, 1377730800, 1377734400, 1377738000, 
    1377741600, 1377745200, 1377748800, 1377752400, 1377756000, 1377759600, 
    1377763200, 1377766800, 1377770400, 1377774000, 1377777600, 1377781200, 
    1377784800, 1377788400, 1377792000, 1377795600, 1377799200, 1377802800, 
    1377806400, 1377810000, 1377813600, 1377817200, 1377820800, 1377824400, 
    1377828000, 1377831600, 1377835200, 1377838800, 1377842400, 1377846000, 
    1377849600, 1377853200, 1377856800, 1377860400, 1377864000, 1377867600, 
    1377871200, 1377874800, 1377878400, 1377882000, 1377885600, 1377889200, 
    1377892800, 1377896400, 1377900000, 1377903600, 1377907200, 1377910800, 
    1377914400, 1377918000, 1377921600, 1377925200, 1377928800, 1377932400, 
    1377936000, 1377939600, 1377943200, 1377946800, 1377950400, 1377954000, 
    1377957600, 1377961200, 1377964800, 1377968400, 1377972000, 1377975600, 
    1377979200, 1377982800, 1377986400, 1377990000, 1377993600, 1377997200, 
    1378000800, 1378004400, 1378008000, 1378011600, 1378015200, 1378018800, 
    1378022400, 1378026000, 1378029600, 1378033200, 1378036800, 1378040400, 
    1378044000, 1378047600, 1378051200, 1378054800, 1378058400, 1378062000, 
    1378065600, 1378069200, 1378072800, 1378076400, 1378080000, 1378083600, 
    1378087200, 1378090800, 1378094400, 1378098000, 1378101600, 1378105200, 
    1378108800, 1378112400, 1378116000, 1378119600, 1378123200, 1378126800, 
    1378130400, 1378134000, 1378137600, 1378141200, 1378144800, 1378148400, 
    1378152000, 1378155600, 1378159200, 1378162800, 1378166400, 1378170000, 
    1378173600, 1378177200, 1378180800, 1378184400, 1378188000, 1378191600, 
    1378195200, 1378198800, 1378202400, 1378206000, 1378209600, 1378213200, 
    1378216800, 1378220400, 1378224000, 1378227600, 1378231200, 1378234800, 
    1378238400, 1378242000, 1378245600, 1378249200, 1378252800, 1378256400, 
    1378260000, 1378263600, 1378267200, 1378270800, 1378274400, 1378278000, 
    1378281600, 1378285200, 1378288800, 1378292400, 1378296000, 1378299600, 
    1378303200, 1378306800, 1378310400, 1378314000, 1378317600, 1378321200, 
    1378324800, 1378328400, 1378332000, 1378335600, 1378339200, 1378342800, 
    1378346400, 1378350000, 1378353600, 1378357200, 1378360800, 1378364400, 
    1378368000, 1378371600, 1378375200, 1378378800, 1378382400, 1378386000, 
    1378389600, 1378393200, 1378396800, 1378400400, 1378404000, 1378407600, 
    1378411200, 1378414800, 1378418400, 1378422000, 1378425600, 1378429200, 
    1378432800, 1378436400, 1378440000, 1378443600, 1378447200, 1378450800, 
    1378454400, 1378458000, 1378461600, 1378465200, 1378468800, 1378472400, 
    1378476000, 1378479600, 1378483200, 1378486800, 1378490400, 1378494000, 
    1378497600, 1378501200, 1378504800, 1378508400, 1378512000, 1378515600, 
    1378519200, 1378522800, 1378526400, 1378530000, 1378533600, 1378537200, 
    1378540800, 1378544400, 1378548000, 1378551600, 1378555200, 1378558800, 
    1378562400, 1378566000, 1378569600, 1378573200, 1378576800, 1378580400, 
    1378584000, 1378587600, 1378591200, 1378594800, 1378598400, 1378602000, 
    1378605600, 1378609200, 1378612800, 1378616400, 1378620000, 1378623600, 
    1378627200, 1378630800, 1378634400, 1378638000, 1378641600, 1378645200, 
    1378648800, 1378652400, 1378656000, 1378659600, 1378663200, 1378666800, 
    1378670400, 1378674000, 1378677600, 1378681200, 1378684800, 1378688400, 
    1378692000, 1378695600, 1378699200, 1378702800, 1378706400, 1378710000, 
    1378713600, 1378717200, 1378720800, 1378724400, 1378728000, 1378731600, 
    1378735200, 1378738800, 1378742400, 1378746000, 1378749600, 1378753200, 
    1378756800, 1378760400, 1378764000, 1378767600, 1378771200, 1378774800, 
    1378778400, 1378782000, 1378785600, 1378789200, 1378792800, 1378796400, 
    1378800000, 1378803600, 1378807200, 1378810800, 1378814400, 1378818000, 
    1378821600, 1378825200, 1378828800, 1378832400, 1378836000, 1378839600, 
    1378843200, 1378846800, 1378850400, 1378854000, 1378857600, 1378861200, 
    1378864800, 1378868400, 1378872000, 1378875600, 1378879200, 1378882800, 
    1378886400, 1378890000, 1378893600, 1378897200, 1378900800, 1378904400, 
    1378908000, 1378911600, 1378915200, 1378918800, 1378922400, 1378926000, 
    1378929600, 1378933200, 1378936800, 1378940400, 1378944000, 1378947600, 
    1378951200, 1378954800, 1378958400, 1378962000, 1378965600, 1378969200, 
    1378972800, 1378976400, 1378980000, 1378983600, 1378987200, 1378990800, 
    1378994400, 1378998000, 1379001600, 1379005200, 1379008800, 1379012400, 
    1379016000, 1379019600, 1379023200, 1379026800, 1379030400, 1379034000, 
    1379037600, 1379041200, 1379044800, 1379048400, 1379052000, 1379055600, 
    1379059200, 1379062800, 1379066400, 1379070000, 1379073600, 1379077200, 
    1379080800, 1379084400, 1379088000, 1379091600, 1379095200, 1379098800, 
    1379102400, 1379106000, 1379109600, 1379113200, 1379116800, 1379120400, 
    1379124000, 1379127600, 1379131200, 1379134800, 1379138400, 1379142000, 
    1379145600, 1379149200, 1379152800, 1379156400, 1379160000, 1379163600, 
    1379167200, 1379170800, 1379174400, 1379178000, 1379181600, 1379185200, 
    1379188800, 1379192400, 1379196000, 1379199600, 1379203200, 1379206800, 
    1379210400, 1379214000, 1379217600, 1379221200, 1379224800, 1379228400, 
    1379232000, 1379235600, 1379239200, 1379242800, 1379246400, 1379250000, 
    1379253600, 1379257200, 1379260800, 1379264400, 1379268000, 1379271600, 
    1379275200, 1379278800, 1379282400, 1379286000, 1379289600, 1379293200, 
    1379296800, 1379300400, 1379304000, 1379307600, 1379311200, 1379314800, 
    1379318400, 1379322000, 1379325600, 1379329200, 1379332800, 1379336400, 
    1379340000, 1379343600, 1379347200, 1379350800, 1379354400, 1379358000, 
    1379361600, 1379365200, 1379368800, 1379372400, 1379376000, 1379379600, 
    1379383200, 1379386800, 1379390400, 1379394000, 1379397600, 1379401200, 
    1379404800, 1379408400, 1379412000, 1379415600, 1379419200, 1379422800, 
    1379426400, 1379430000, 1379433600, 1379437200, 1379440800, 1379444400, 
    1379448000, 1379451600, 1379455200, 1379458800, 1379462400, 1379466000, 
    1379469600, 1379473200, 1379476800, 1379480400, 1379484000, 1379487600, 
    1379491200, 1379494800, 1379498400, 1379502000, 1379505600, 1379509200, 
    1379512800, 1379516400, 1379520000, 1379523600, 1379527200, 1379530800, 
    1379534400, 1379538000, 1379541600, 1379545200, 1379548800, 1379552400, 
    1379556000, 1379559600, 1379563200, 1379566800, 1379570400, 1379574000, 
    1379577600, 1379581200, 1379584800, 1379588400, 1379592000, 1379595600, 
    1379599200, 1379602800, 1379606400, 1379610000, 1379613600, 1379617200, 
    1379620800, 1379624400, 1379628000, 1379631600, 1379635200, 1379638800, 
    1379642400, 1379646000, 1379649600, 1379653200, 1379656800, 1379660400, 
    1379664000, 1379667600, 1379671200, 1379674800, 1379678400, 1379682000, 
    1379685600, 1379689200, 1379692800, 1379696400, 1379700000, 1379703600, 
    1379707200, 1379710800, 1379714400, 1379718000, 1379721600, 1379725200, 
    1379728800, 1379732400, 1379736000, 1379739600, 1379743200, 1379746800, 
    1379750400, 1379754000, 1379757600, 1379761200, 1379764800, 1379768400, 
    1379772000, 1379775600, 1379779200, 1379782800, 1379786400, 1379790000, 
    1379793600, 1379797200, 1379800800, 1379804400, 1379808000, 1379811600, 
    1379815200, 1379818800, 1379822400, 1379826000, 1379829600, 1379833200, 
    1379836800, 1379840400, 1379844000, 1379847600, 1379851200, 1379854800, 
    1379858400, 1379862000, 1379865600, 1379869200, 1379872800, 1379876400, 
    1379880000, 1379883600, 1379887200, 1379890800, 1379894400, 1379898000, 
    1379901600, 1379905200, 1379908800, 1379912400, 1379916000, 1379919600, 
    1379923200, 1379926800, 1379930400, 1379934000, 1379937600, 1379941200, 
    1379944800, 1379948400, 1379952000, 1379955600, 1379959200, 1379962800, 
    1379966400, 1379970000, 1379973600, 1379977200, 1379980800, 1379984400, 
    1379988000, 1379991600, 1379995200, 1379998800, 1380002400, 1380006000, 
    1380009600, 1380013200, 1380016800, 1380020400, 1380024000, 1380027600, 
    1380031200, 1380034800, 1380038400, 1380042000, 1380045600, 1380049200, 
    1380052800, 1380056400, 1380060000, 1380063600, 1380067200, 1380070800, 
    1380074400, 1380078000, 1380081600, 1380085200, 1380088800, 1380092400, 
    1380096000, 1380099600, 1380103200, 1380106800, 1380110400, 1380114000, 
    1380117600, 1380121200, 1380124800, 1380128400, 1380132000, 1380135600, 
    1380139200, 1380142800, 1380146400, 1380150000, 1380153600, 1380157200, 
    1380160800, 1380164400, 1380168000, 1380171600, 1380175200, 1380178800, 
    1380182400, 1380186000, 1380189600, 1380193200, 1380196800, 1380200400, 
    1380204000, 1380207600, 1380211200, 1380214800, 1380218400, 1380222000, 
    1380225600, 1380229200, 1380232800, 1380236400, 1380240000, 1380243600, 
    1380247200, 1380250800, 1380254400, 1380258000, 1380261600, 1380265200, 
    1380268800, 1380272400, 1380276000, 1380279600, 1380283200, 1380286800, 
    1380290400, 1380294000, 1380297600, 1380301200, 1380304800, 1380308400, 
    1380312000, 1380315600, 1380319200, 1380322800, 1380326400, 1380330000, 
    1380333600, 1380337200, 1380340800, 1380344400, 1380348000, 1380351600, 
    1380355200, 1380358800, 1380362400, 1380366000, 1380369600, 1380373200, 
    1380376800, 1380380400, 1380384000, 1380387600, 1380391200, 1380394800, 
    1380398400, 1380402000, 1380405600, 1380409200, 1380412800, 1380416400, 
    1380420000, 1380423600, 1380427200, 1380430800, 1380434400, 1380438000, 
    1380441600, 1380445200, 1380448800, 1380452400, 1380456000, 1380459600, 
    1380463200, 1380466800, 1380470400, 1380474000, 1380477600, 1380481200, 
    1380484800, 1380488400, 1380492000, 1380495600, 1380499200, 1380502800, 
    1380506400, 1380510000, 1380513600, 1380517200, 1380520800, 1380524400, 
    1380528000, 1380531600, 1380535200, 1380538800, 1380542400, 1380546000, 
    1380549600, 1380553200, 1380556800, 1380560400, 1380564000, 1380567600, 
    1380571200, 1380574800, 1380578400, 1380582000, 1380585600, 1380589200, 
    1380592800, 1380596400, 1380600000, 1380603600, 1380607200, 1380610800, 
    1380614400, 1380618000, 1380621600, 1380625200, 1380628800, 1380632400, 
    1380636000, 1380639600, 1380643200, 1380646800, 1380650400, 1380654000, 
    1380657600, 1380661200, 1380664800, 1380668400, 1380672000, 1380675600, 
    1380679200, 1380682800, 1380686400, 1380690000, 1380693600, 1380697200, 
    1380700800, 1380704400, 1380708000, 1380711600, 1380715200, 1380718800, 
    1380722400, 1380726000, 1380729600, 1380733200, 1380736800, 1380740400, 
    1380744000, 1380747600, 1380751200, 1380754800, 1380758400, 1380762000, 
    1380765600, 1380769200, 1380772800, 1380776400, 1380780000, 1380783600, 
    1380787200, 1380790800, 1380794400, 1380798000, 1380801600, 1380805200, 
    1380808800, 1380812400, 1380816000, 1380819600, 1380823200, 1380826800, 
    1380830400, 1380834000, 1380837600, 1380841200, 1380844800, 1380848400, 
    1380852000, 1380855600, 1380859200, 1380862800, 1380866400, 1380870000, 
    1380873600, 1380877200, 1380880800, 1380884400, 1380888000, 1380891600, 
    1380895200, 1380898800, 1380902400, 1380906000, 1380909600, 1380913200, 
    1380916800, 1380920400, 1380924000, 1380927600, 1380931200, 1380934800, 
    1380938400, 1380942000, 1380945600, 1380949200, 1380952800, 1380956400, 
    1380960000, 1380963600, 1380967200, 1380970800, 1380974400, 1380978000, 
    1380981600, 1380985200, 1380988800, 1380992400, 1380996000, 1380999600, 
    1381003200, 1381006800, 1381010400, 1381014000, 1381017600, 1381021200, 
    1381024800, 1381028400, 1381032000, 1381035600, 1381039200, 1381042800, 
    1381046400, 1381050000, 1381053600, 1381057200, 1381060800, 1381064400, 
    1381068000, 1381071600, 1381075200, 1381078800, 1381082400, 1381086000, 
    1381089600, 1381093200, 1381096800, 1381100400, 1381104000, 1381107600, 
    1381111200, 1381114800, 1381118400, 1381122000, 1381125600, 1381129200, 
    1381132800, 1381136400, 1381140000, 1381143600, 1381147200, 1381150800, 
    1381154400, 1381158000, 1381161600, 1381165200, 1381168800, 1381172400, 
    1381176000, 1381179600, 1381183200, 1381186800, 1381190400, 1381194000, 
    1381197600, 1381201200, 1381204800, 1381208400, 1381212000, 1381215600, 
    1381219200, 1381222800, 1381226400, 1381230000, 1381233600, 1381237200, 
    1381240800, 1381244400, 1381248000, 1381251600, 1381255200, 1381258800, 
    1381262400, 1381266000, 1381269600, 1381273200, 1381276800, 1381280400, 
    1381284000, 1381287600, 1381291200, 1381294800, 1381298400, 1381302000, 
    1381305600, 1381309200, 1381312800, 1381316400, 1381320000, 1381323600, 
    1381327200, 1381330800, 1381334400, 1381338000, 1381341600, 1381345200, 
    1381348800, 1381352400, 1381356000, 1381359600, 1381363200, 1381366800, 
    1381370400, 1381374000, 1381377600, 1381381200, 1381384800, 1381388400, 
    1381392000, 1381395600, 1381399200, 1381402800, 1381406400, 1381410000, 
    1381413600, 1381417200, 1381420800, 1381424400, 1381428000, 1381431600, 
    1381435200, 1381438800, 1381442400, 1381446000, 1381449600, 1381453200, 
    1381456800, 1381460400, 1381464000, 1381467600, 1381471200, 1381474800, 
    1381478400, 1381482000, 1381485600, 1381489200, 1381492800, 1381496400, 
    1381500000, 1381503600, 1381507200, 1381510800, 1381514400, 1381518000, 
    1381521600, 1381525200, 1381528800, 1381532400, 1381536000, 1381539600, 
    1381543200, 1381546800, 1381550400, 1381554000, 1381557600, 1381561200, 
    1381564800, 1381568400, 1381572000, 1381575600, 1381579200, 1381582800, 
    1381586400, 1381590000, 1381593600, 1381597200, 1381600800, 1381604400, 
    1381608000, 1381611600, 1381615200, 1381618800, 1381622400, 1381626000, 
    1381629600, 1381633200, 1381636800, 1381640400, 1381644000, 1381647600, 
    1381651200, 1381654800, 1381658400, 1381662000, 1381665600, 1381669200, 
    1381672800, 1381676400, 1381680000, 1381683600, 1381687200, 1381690800, 
    1381694400, 1381698000, 1381701600, 1381705200, 1381708800, 1381712400, 
    1381716000, 1381719600, 1381723200, 1381726800, 1381730400, 1381734000, 
    1381737600, 1381741200, 1381744800, 1381748400, 1381752000, 1381755600, 
    1381759200, 1381762800, 1381766400, 1381770000, 1381773600, 1381777200, 
    1381780800, 1381784400, 1381788000, 1381791600, 1381795200, 1381798800, 
    1381802400, 1381806000, 1381809600, 1381813200, 1381816800, 1381820400, 
    1381824000, 1381827600, 1381831200, 1381834800, 1381838400, 1381842000, 
    1381845600, 1381849200, 1381852800, 1381856400, 1381860000, 1381863600, 
    1381867200, 1381870800, 1381874400, 1381878000, 1381881600, 1381885200, 
    1381888800, 1381892400, 1381896000, 1381899600, 1381903200, 1381906800, 
    1381910400, 1381914000, 1381917600, 1381921200, 1381924800, 1381928400, 
    1381932000, 1381935600, 1381939200, 1381942800, 1381946400, 1381950000, 
    1381953600, 1381957200, 1381960800, 1381964400, 1381968000, 1381971600, 
    1381975200, 1381978800, 1381982400, 1381986000, 1381989600, 1381993200, 
    1381996800, 1382000400, 1382004000, 1382007600, 1382011200, 1382014800, 
    1382018400, 1382022000, 1382025600, 1382029200, 1382032800, 1382036400, 
    1382040000, 1382043600, 1382047200, 1382050800, 1382054400, 1382058000, 
    1382061600, 1382065200, 1382068800, 1382072400, 1382076000, 1382079600, 
    1382083200, 1382086800, 1382090400, 1382094000, 1382097600, 1382101200, 
    1382104800, 1382108400, 1382112000, 1382115600, 1382119200, 1382122800, 
    1382126400, 1382130000, 1382133600, 1382137200, 1382140800, 1382144400, 
    1382148000, 1382151600, 1382155200, 1382158800, 1382162400, 1382166000, 
    1382169600, 1382173200, 1382176800, 1382180400, 1382184000, 1382187600, 
    1382191200, 1382194800, 1382198400, 1382202000, 1382205600, 1382209200, 
    1382212800, 1382216400, 1382220000, 1382223600, 1382227200, 1382230800, 
    1382234400, 1382238000, 1382241600, 1382245200, 1382248800, 1382252400, 
    1382256000, 1382259600, 1382263200, 1382266800, 1382270400, 1382274000, 
    1382277600, 1382281200, 1382284800, 1382288400, 1382292000, 1382295600, 
    1382299200, 1382302800, 1382306400, 1382310000, 1382313600, 1382317200, 
    1382320800, 1382324400, 1382328000, 1382331600, 1382335200, 1382338800, 
    1382342400, 1382346000, 1382349600, 1382353200, 1382356800, 1382360400, 
    1382364000, 1382367600, 1382371200, 1382374800, 1382378400, 1382382000, 
    1382385600, 1382389200, 1382392800, 1382396400, 1382400000, 1382403600, 
    1382407200, 1382410800, 1382414400, 1382418000, 1382421600, 1382425200, 
    1382428800, 1382432400, 1382436000, 1382439600, 1382443200, 1382446800, 
    1382450400, 1382454000, 1382457600, 1382461200, 1382464800, 1382468400, 
    1382472000, 1382475600, 1382479200, 1382482800, 1382486400, 1382490000, 
    1382493600, 1382497200, 1382500800, 1382504400, 1382508000, 1382511600, 
    1382515200, 1382518800, 1382522400, 1382526000, 1382529600, 1382533200, 
    1382536800, 1382540400, 1382544000, 1382547600, 1382551200, 1382554800, 
    1382558400, 1382562000, 1382565600, 1382569200, 1382572800, 1382576400, 
    1382580000, 1382583600, 1382587200, 1382590800, 1382594400, 1382598000, 
    1382601600, 1382605200, 1382608800, 1382612400, 1382616000, 1382619600, 
    1382623200, 1382626800, 1382630400, 1382634000, 1382637600, 1382641200, 
    1382644800, 1382648400, 1382652000, 1382655600, 1382659200, 1382662800, 
    1382666400, 1382670000, 1382673600, 1382677200, 1382680800, 1382684400, 
    1382688000, 1382691600, 1382695200, 1382698800, 1382702400, 1382706000, 
    1382709600, 1382713200, 1382716800, 1382720400, 1382724000, 1382727600, 
    1382731200, 1382734800, 1382738400, 1382742000, 1382745600, 1382749200, 
    1382752800, 1382756400, 1382760000, 1382763600, 1382767200, 1382770800, 
    1382774400, 1382778000, 1382781600, 1382785200, 1382788800, 1382792400, 
    1382796000, 1382799600, 1382803200, 1382806800, 1382810400, 1382814000, 
    1382817600, 1382821200, 1382824800, 1382828400, 1382832000, 1382835600, 
    1382839200, 1382842800, 1382846400, 1382850000, 1382853600, 1382857200, 
    1382860800, 1382864400, 1382868000, 1382871600, 1382875200, 1382878800, 
    1382882400, 1382886000, 1382889600, 1382893200, 1382896800, 1382900400, 
    1382904000, 1382907600, 1382911200, 1382914800, 1382918400, 1382922000, 
    1382925600, 1382929200, 1382932800, 1382936400, 1382940000, 1382943600, 
    1382947200, 1382950800, 1382954400, 1382958000, 1382961600, 1382965200, 
    1382968800, 1382972400, 1382976000, 1382979600, 1382983200, 1382986800, 
    1382990400, 1382994000, 1382997600, 1383001200, 1383004800, 1383008400, 
    1383012000, 1383015600, 1383019200, 1383022800, 1383026400, 1383030000, 
    1383033600, 1383037200, 1383040800, 1383044400, 1383048000, 1383051600, 
    1383055200, 1383058800, 1383062400, 1383066000, 1383069600, 1383073200, 
    1383076800, 1383080400, 1383084000, 1383087600, 1383091200, 1383094800, 
    1383098400, 1383102000, 1383105600, 1383109200, 1383112800, 1383116400, 
    1383120000, 1383123600, 1383127200, 1383130800, 1383134400, 1383138000, 
    1383141600, 1383145200, 1383148800, 1383152400, 1383156000, 1383159600, 
    1383163200, 1383166800, 1383170400, 1383174000, 1383177600, 1383181200, 
    1383184800, 1383188400, 1383192000, 1383195600, 1383199200, 1383202800, 
    1383206400, 1383210000, 1383213600, 1383217200, 1383220800, 1383224400, 
    1383228000, 1383231600, 1383235200, 1383238800, 1383242400, 1383246000, 
    1383249600, 1383253200, 1383256800, 1383260400, 1383264000, 1383267600, 
    1383271200, 1383274800, 1383278400, 1383282000, 1383285600, 1383289200, 
    1383292800, 1383296400, 1383300000, 1383303600, 1383307200, 1383310800, 
    1383314400, 1383318000, 1383321600, 1383325200, 1383328800, 1383332400, 
    1383336000, 1383339600, 1383343200, 1383346800, 1383350400, 1383354000, 
    1383357600, 1383361200, 1383364800, 1383368400, 1383372000, 1383375600, 
    1383379200, 1383382800, 1383386400, 1383390000, 1383393600, 1383397200, 
    1383400800, 1383404400, 1383408000, 1383411600, 1383415200, 1383418800, 
    1383422400, 1383426000, 1383429600, 1383433200, 1383436800, 1383440400, 
    1383444000, 1383447600, 1383451200, 1383454800, 1383458400, 1383462000, 
    1383465600, 1383469200, 1383472800, 1383476400, 1383480000, 1383483600, 
    1383487200, 1383490800, 1383494400, 1383498000, 1383501600, 1383505200, 
    1383508800, 1383512400, 1383516000, 1383519600, 1383523200, 1383526800, 
    1383530400, 1383534000, 1383537600, 1383541200, 1383544800, 1383548400, 
    1383552000, 1383555600, 1383559200, 1383562800, 1383566400, 1383570000, 
    1383573600, 1383577200, 1383580800, 1383584400, 1383588000, 1383591600, 
    1383595200, 1383598800, 1383602400, 1383606000, 1383609600, 1383613200, 
    1383616800, 1383620400, 1383624000, 1383627600, 1383631200, 1383634800, 
    1383638400, 1383642000, 1383645600, 1383649200, 1383652800, 1383656400, 
    1383660000, 1383663600, 1383667200, 1383670800, 1383674400, 1383678000, 
    1383681600, 1383685200, 1383688800, 1383692400, 1383696000, 1383699600, 
    1383703200, 1383706800, 1383710400, 1383714000, 1383717600, 1383721200, 
    1383724800, 1383728400, 1383732000, 1383735600, 1383739200, 1383742800, 
    1383746400, 1383750000, 1383753600, 1383757200, 1383760800, 1383764400, 
    1383768000, 1383771600, 1383775200, 1383778800, 1383782400, 1383786000, 
    1383789600, 1383793200, 1383796800, 1383800400, 1383804000, 1383807600, 
    1383811200, 1383814800, 1383818400, 1383822000, 1383825600, 1383829200, 
    1383832800, 1383836400, 1383840000, 1383843600, 1383847200, 1383850800, 
    1383854400, 1383858000, 1383861600, 1383865200, 1383868800, 1383872400, 
    1383876000, 1383879600, 1383883200, 1383886800, 1383890400, 1383894000, 
    1383897600, 1383901200, 1383904800, 1383908400, 1383912000, 1383915600, 
    1383919200, 1383922800, 1383926400, 1383930000, 1383933600, 1383937200, 
    1383940800, 1383944400, 1383948000, 1383951600, 1383955200, 1383958800, 
    1383962400, 1383966000, 1383969600, 1383973200, 1383976800, 1383980400, 
    1383984000, 1383987600, 1383991200, 1383994800, 1383998400, 1384002000, 
    1384005600, 1384009200, 1384012800, 1384016400, 1384020000, 1384023600, 
    1384027200, 1384030800, 1384034400, 1384038000, 1384041600, 1384045200, 
    1384048800, 1384052400, 1384056000, 1384059600, 1384063200, 1384066800, 
    1384070400, 1384074000, 1384077600, 1384081200, 1384084800, 1384088400, 
    1384092000, 1384095600, 1384099200, 1384102800, 1384106400, 1384110000, 
    1384113600, 1384117200, 1384120800, 1384124400, 1384128000, 1384131600, 
    1384135200, 1384138800, 1384142400, 1384146000, 1384149600, 1384153200, 
    1384156800, 1384160400, 1384164000, 1384167600, 1384171200, 1384174800, 
    1384178400, 1384182000, 1384185600, 1384189200, 1384192800, 1384196400, 
    1384200000, 1384203600, 1384207200, 1384210800, 1384214400, 1384218000, 
    1384221600, 1384225200, 1384228800, 1384232400, 1384236000, 1384239600, 
    1384243200, 1384246800, 1384250400, 1384254000, 1384257600, 1384261200, 
    1384264800, 1384268400, 1384272000, 1384275600, 1384279200, 1384282800, 
    1384286400, 1384290000, 1384293600, 1384297200, 1384300800, 1384304400, 
    1384308000, 1384311600, 1384315200, 1384318800, 1384322400, 1384326000, 
    1384329600, 1384333200, 1384336800, 1384340400, 1384344000, 1384347600, 
    1384351200, 1384354800, 1384358400, 1384362000, 1384365600, 1384369200, 
    1384372800, 1384376400, 1384380000, 1384383600, 1384387200, 1384390800, 
    1384394400, 1384398000, 1384401600, 1384405200, 1384408800, 1384412400, 
    1384416000, 1384419600, 1384423200, 1384426800, 1384430400, 1384434000, 
    1384437600, 1384441200, 1384444800, 1384448400, 1384452000, 1384455600, 
    1384459200, 1384462800, 1384466400, 1384470000, 1384473600, 1384477200, 
    1384480800, 1384484400, 1384488000, 1384491600, 1384495200, 1384498800, 
    1384502400, 1384506000, 1384509600, 1384513200, 1384516800, 1384520400, 
    1384524000, 1384527600, 1384531200, 1384534800, 1384538400, 1384542000, 
    1384545600, 1384549200, 1384552800, 1384556400, 1384560000, 1384563600, 
    1384567200, 1384570800, 1384574400, 1384578000, 1384581600, 1384585200, 
    1384588800, 1384592400, 1384596000, 1384599600, 1384603200, 1384606800, 
    1384610400, 1384614000, 1384617600, 1384621200, 1384624800, 1384628400, 
    1384632000, 1384635600, 1384639200, 1384642800, 1384646400, 1384650000, 
    1384653600, 1384657200, 1384660800, 1384664400, 1384668000, 1384671600, 
    1384675200, 1384678800, 1384682400, 1384686000, 1384689600, 1384693200, 
    1384696800, 1384700400, 1384704000, 1384707600, 1384711200, 1384714800, 
    1384718400, 1384722000, 1384725600, 1384729200, 1384732800, 1384736400, 
    1384740000, 1384743600, 1384747200, 1384750800, 1384754400, 1384758000, 
    1384761600, 1384765200, 1384768800, 1384772400, 1384776000, 1384779600, 
    1384783200, 1384786800, 1384790400, 1384794000, 1384797600, 1384801200, 
    1384804800, 1384808400, 1384812000, 1384815600, 1384819200, 1384822800, 
    1384826400, 1384830000, 1384833600, 1384837200, 1384840800, 1384844400, 
    1384848000, 1384851600, 1384855200, 1384858800, 1384862400, 1384866000, 
    1384869600, 1384873200, 1384876800, 1384880400, 1384884000, 1384887600, 
    1384891200, 1384894800, 1384898400, 1384902000, 1384905600, 1384909200, 
    1384912800, 1384916400, 1384920000, 1384923600, 1384927200, 1384930800, 
    1384934400, 1384938000, 1384941600, 1384945200, 1384948800, 1384952400, 
    1384956000, 1384959600, 1384963200, 1384966800, 1384970400, 1384974000, 
    1384977600, 1384981200, 1384984800, 1384988400, 1384992000, 1384995600, 
    1384999200, 1385002800, 1385006400, 1385010000, 1385013600, 1385017200, 
    1385020800, 1385024400, 1385028000, 1385031600, 1385035200, 1385038800, 
    1385042400, 1385046000, 1385049600, 1385053200, 1385056800, 1385060400, 
    1385064000, 1385067600, 1385071200, 1385074800, 1385078400, 1385082000, 
    1385085600, 1385089200, 1385092800, 1385096400, 1385100000, 1385103600, 
    1385107200, 1385110800, 1385114400, 1385118000, 1385121600, 1385125200, 
    1385128800, 1385132400, 1385136000, 1385139600, 1385143200, 1385146800, 
    1385150400, 1385154000, 1385157600, 1385161200, 1385164800, 1385168400, 
    1385172000, 1385175600, 1385179200, 1385182800, 1385186400, 1385190000, 
    1385193600, 1385197200, 1385200800, 1385204400, 1385208000, 1385211600, 
    1385215200, 1385218800, 1385222400, 1385226000, 1385229600, 1385233200, 
    1385236800, 1385240400, 1385244000, 1385247600, 1385251200, 1385254800, 
    1385258400, 1385262000, 1385265600, 1385269200, 1385272800, 1385276400, 
    1385280000, 1385283600, 1385287200, 1385290800, 1385294400, 1385298000, 
    1385301600, 1385305200, 1385308800, 1385312400, 1385316000, 1385319600, 
    1385323200, 1385326800, 1385330400, 1385334000, 1385337600, 1385341200, 
    1385344800, 1385348400, 1385352000, 1385355600, 1385359200, 1385362800, 
    1385366400, 1385370000, 1385373600, 1385377200, 1385380800, 1385384400, 
    1385388000, 1385391600, 1385395200, 1385398800, 1385402400, 1385406000, 
    1385409600, 1385413200, 1385416800, 1385420400, 1385424000, 1385427600, 
    1385431200, 1385434800, 1385438400, 1385442000, 1385445600, 1385449200, 
    1385452800, 1385456400, 1385460000, 1385463600, 1385467200, 1385470800, 
    1385474400, 1385478000, 1385481600, 1385485200, 1385488800, 1385492400, 
    1385496000, 1385499600, 1385503200, 1385506800, 1385510400, 1385514000, 
    1385517600, 1385521200, 1385524800, 1385528400, 1385532000, 1385535600, 
    1385539200, 1385542800, 1385546400, 1385550000, 1385553600, 1385557200, 
    1385560800, 1385564400, 1385568000, 1385571600, 1385575200, 1385578800, 
    1385582400, 1385586000, 1385589600, 1385593200, 1385596800, 1385600400, 
    1385604000, 1385607600, 1385611200, 1385614800, 1385618400, 1385622000, 
    1385625600, 1385629200, 1385632800, 1385636400, 1385640000, 1385643600, 
    1385647200, 1385650800, 1385654400, 1385658000, 1385661600, 1385665200, 
    1385668800, 1385672400, 1385676000, 1385679600, 1385683200, 1385686800, 
    1385690400, 1385694000, 1385697600, 1385701200, 1385704800, 1385708400, 
    1385712000, 1385715600, 1385719200, 1385722800, 1385726400, 1385730000, 
    1385733600, 1385737200, 1385740800, 1385744400, 1385748000, 1385751600, 
    1385755200, 1385758800, 1385762400, 1385766000, 1385769600, 1385773200, 
    1385776800, 1385780400, 1385784000, 1385787600, 1385791200, 1385794800, 
    1385798400, 1385802000, 1385805600, 1385809200, 1385812800, 1385816400, 
    1385820000, 1385823600, 1385827200, 1385830800, 1385834400, 1385838000, 
    1385841600, 1385845200, 1385848800, 1385852400, 1385856000, 1385859600, 
    1385863200, 1385866800, 1385870400, 1385874000, 1385877600, 1385881200, 
    1385884800, 1385888400, 1385892000, 1385895600, 1385899200, 1385902800, 
    1385906400, 1385910000, 1385913600, 1385917200, 1385920800, 1385924400, 
    1385928000, 1385931600, 1385935200, 1385938800, 1385942400, 1385946000, 
    1385949600, 1385953200, 1385956800, 1385960400, 1385964000, 1385967600, 
    1385971200, 1385974800, 1385978400, 1385982000, 1385985600, 1385989200, 
    1385992800, 1385996400, 1386000000, 1386003600, 1386007200, 1386010800, 
    1386014400, 1386018000, 1386021600, 1386025200, 1386028800, 1386032400, 
    1386036000, 1386039600, 1386043200, 1386046800, 1386050400, 1386054000, 
    1386057600, 1386061200, 1386064800, 1386068400, 1386072000, 1386075600, 
    1386079200, 1386082800, 1386086400, 1386090000, 1386093600, 1386097200, 
    1386100800, 1386104400, 1386108000, 1386111600, 1386115200, 1386118800, 
    1386122400, 1386126000, 1386129600, 1386133200, 1386136800, 1386140400, 
    1386144000, 1386147600, 1386151200, 1386154800, 1386158400, 1386162000, 
    1386165600, 1386169200, 1386172800, 1386176400, 1386180000, 1386183600, 
    1386187200, 1386190800, 1386194400, 1386198000, 1386201600, 1386205200, 
    1386208800, 1386212400, 1386216000, 1386219600, 1386223200, 1386226800, 
    1386230400, 1386234000, 1386237600, 1386241200, 1386244800, 1386248400, 
    1386252000, 1386255600, 1386259200, 1386262800, 1386266400, 1386270000, 
    1386273600, 1386277200, 1386280800, 1386284400, 1386288000, 1386291600, 
    1386295200, 1386298800, 1386302400, 1386306000, 1386309600, 1386313200, 
    1386316800, 1386320400, 1386324000, 1386327600, 1386331200, 1386334800, 
    1386338400, 1386342000, 1386345600, 1386349200, 1386352800, 1386356400, 
    1386360000, 1386363600, 1386367200, 1386370800, 1386374400, 1386378000, 
    1386381600, 1386385200, 1386388800, 1386392400, 1386396000, 1386399600, 
    1386403200, 1386406800, 1386410400, 1386414000, 1386417600, 1386421200, 
    1386424800, 1386428400, 1386432000, 1386435600, 1386439200, 1386442800, 
    1386446400, 1386450000, 1386453600, 1386457200, 1386460800, 1386464400, 
    1386468000, 1386471600, 1386475200, 1386478800, 1386482400, 1386486000, 
    1386489600, 1386493200, 1386496800, 1386500400, 1386504000, 1386507600, 
    1386511200, 1386514800, 1386518400, 1386522000, 1386525600, 1386529200, 
    1386532800, 1386536400, 1386540000, 1386543600, 1386547200, 1386550800, 
    1386554400, 1386558000, 1386561600, 1386565200, 1386568800, 1386572400, 
    1386576000, 1386579600, 1386583200, 1386586800, 1386590400, 1386594000, 
    1386597600, 1386601200, 1386604800, 1386608400, 1386612000, 1386615600, 
    1386619200, 1386622800, 1386626400, 1386630000, 1386633600, 1386637200, 
    1386640800, 1386644400, 1386648000, 1386651600, 1386655200, 1386658800, 
    1386662400, 1386666000, 1386669600, 1386673200, 1386676800, 1386680400, 
    1386684000, 1386687600, 1386691200, 1386694800, 1386698400, 1386702000, 
    1386705600, 1386709200, 1386712800, 1386716400, 1386720000, 1386723600, 
    1386727200, 1386730800, 1386734400, 1386738000, 1386741600, 1386745200, 
    1386748800, 1386752400, 1386756000, 1386759600, 1386763200, 1386766800, 
    1386770400, 1386774000, 1386777600, 1386781200, 1386784800, 1386788400, 
    1386792000, 1386795600, 1386799200, 1386802800, 1386806400, 1386810000, 
    1386813600, 1386817200, 1386820800, 1386824400, 1386828000, 1386831600, 
    1386835200, 1386838800, 1386842400, 1386846000, 1386849600, 1386853200, 
    1386856800, 1386860400, 1386864000, 1386867600, 1386871200, 1386874800, 
    1386878400, 1386882000, 1386885600, 1386889200, 1386892800, 1386896400, 
    1386900000, 1386903600, 1386907200, 1386910800, 1386914400, 1386918000, 
    1386921600, 1386925200, 1386928800, 1386932400, 1386936000, 1386939600, 
    1386943200, 1386946800, 1386950400, 1386954000, 1386957600, 1386961200, 
    1386964800, 1386968400, 1386972000, 1386975600, 1386979200, 1386982800, 
    1386986400, 1386990000, 1386993600, 1386997200, 1387000800, 1387004400, 
    1387008000, 1387011600, 1387015200, 1387018800, 1387022400, 1387026000, 
    1387029600, 1387033200, 1387036800, 1387040400, 1387044000, 1387047600, 
    1387051200, 1387054800, 1387058400, 1387062000, 1387065600, 1387069200, 
    1387072800, 1387076400, 1387080000, 1387083600, 1387087200, 1387090800, 
    1387094400, 1387098000, 1387101600, 1387105200, 1387108800, 1387112400, 
    1387116000, 1387119600, 1387123200, 1387126800, 1387130400, 1387134000, 
    1387137600, 1387141200, 1387144800, 1387148400, 1387152000, 1387155600, 
    1387159200, 1387162800, 1387166400, 1387170000, 1387173600, 1387177200, 
    1387180800, 1387184400, 1387188000, 1387191600, 1387195200, 1387198800, 
    1387202400, 1387206000, 1387209600, 1387213200, 1387216800, 1387220400, 
    1387224000, 1387227600, 1387231200, 1387234800, 1387238400, 1387242000, 
    1387245600, 1387249200, 1387252800, 1387256400, 1387260000, 1387263600, 
    1387267200, 1387270800, 1387274400, 1387278000, 1387281600, 1387285200, 
    1387288800, 1387292400, 1387296000, 1387299600, 1387303200, 1387306800, 
    1387310400, 1387314000, 1387317600, 1387321200, 1387324800, 1387328400, 
    1387332000, 1387335600, 1387339200, 1387342800, 1387346400, 1387350000, 
    1387353600, 1387357200, 1387360800, 1387364400, 1387368000, 1387371600, 
    1387375200, 1387378800, 1387382400, 1387386000, 1387389600, 1387393200, 
    1387396800, 1387400400, 1387404000, 1387407600, 1387411200, 1387414800, 
    1387418400, 1387422000, 1387425600, 1387429200, 1387432800, 1387436400, 
    1387440000, 1387443600, 1387447200, 1387450800, 1387454400, 1387458000, 
    1387461600, 1387465200, 1387468800, 1387472400, 1387476000, 1387479600, 
    1387483200, 1387486800, 1387490400, 1387494000, 1387497600, 1387501200, 
    1387504800, 1387508400, 1387512000, 1387515600, 1387519200, 1387522800, 
    1387526400, 1387530000, 1387533600, 1387537200, 1387540800, 1387544400, 
    1387548000, 1387551600, 1387555200, 1387558800, 1387562400, 1387566000, 
    1387569600, 1387573200, 1387576800, 1387580400, 1387584000, 1387587600, 
    1387591200, 1387594800, 1387598400, 1387602000, 1387605600, 1387609200, 
    1387612800, 1387616400, 1387620000, 1387623600, 1387627200, 1387630800, 
    1387634400, 1387638000, 1387641600, 1387645200, 1387648800, 1387652400, 
    1387656000, 1387659600, 1387663200, 1387666800, 1387670400, 1387674000, 
    1387677600, 1387681200, 1387684800, 1387688400, 1387692000, 1387695600, 
    1387699200, 1387702800, 1387706400, 1387710000, 1387713600, 1387717200, 
    1387720800, 1387724400, 1387728000, 1387731600, 1387735200, 1387738800, 
    1387742400, 1387746000, 1387749600, 1387753200, 1387756800, 1387760400, 
    1387764000, 1387767600, 1387771200, 1387774800, 1387778400, 1387782000, 
    1387785600, 1387789200, 1387792800, 1387796400, 1387800000, 1387803600, 
    1387807200, 1387810800, 1387814400, 1387818000, 1387821600, 1387825200, 
    1387828800, 1387832400, 1387836000, 1387839600, 1387843200, 1387846800, 
    1387850400, 1387854000, 1387857600, 1387861200, 1387864800, 1387868400, 
    1387872000, 1387875600, 1387879200, 1387882800, 1387886400, 1387890000, 
    1387893600, 1387897200, 1387900800, 1387904400, 1387908000, 1387911600, 
    1387915200, 1387918800, 1387922400, 1387926000, 1387929600, 1387933200, 
    1387936800, 1387940400, 1387944000, 1387947600, 1387951200, 1387954800, 
    1387958400, 1387962000, 1387965600, 1387969200, 1387972800, 1387976400, 
    1387980000, 1387983600, 1387987200, 1387990800, 1387994400, 1387998000, 
    1388001600, 1388005200, 1388008800, 1388012400, 1388016000, 1388019600, 
    1388023200, 1388026800, 1388030400, 1388034000, 1388037600, 1388041200, 
    1388044800, 1388048400, 1388052000, 1388055600, 1388059200, 1388062800, 
    1388066400, 1388070000, 1388073600, 1388077200, 1388080800, 1388084400, 
    1388088000, 1388091600, 1388095200, 1388098800, 1388102400, 1388106000, 
    1388109600, 1388113200, 1388116800, 1388120400, 1388124000, 1388127600, 
    1388131200, 1388134800, 1388138400, 1388142000, 1388145600, 1388149200, 
    1388152800, 1388156400, 1388160000, 1388163600, 1388167200, 1388170800, 
    1388174400, 1388178000, 1388181600, 1388185200, 1388188800, 1388192400, 
    1388196000, 1388199600, 1388203200, 1388206800, 1388210400, 1388214000, 
    1388217600, 1388221200, 1388224800, 1388228400, 1388232000, 1388235600, 
    1388239200, 1388242800, 1388246400, 1388250000, 1388253600, 1388257200, 
    1388260800, 1388264400, 1388268000, 1388271600, 1388275200, 1388278800, 
    1388282400, 1388286000, 1388289600, 1388293200, 1388296800, 1388300400, 
    1388304000, 1388307600, 1388311200, 1388314800, 1388318400, 1388322000, 
    1388325600, 1388329200, 1388332800, 1388336400, 1388340000, 1388343600, 
    1388347200, 1388350800, 1388354400, 1388358000, 1388361600, 1388365200, 
    1388368800, 1388372400, 1388376000, 1388379600, 1388383200, 1388386800, 
    1388390400, 1388394000, 1388397600, 1388401200, 1388404800, 1388408400, 
    1388412000, 1388415600, 1388419200, 1388422800, 1388426400, 1388430000, 
    1388433600, 1388437200, 1388440800, 1388444400, 1388448000, 1388451600, 
    1388455200, 1388458800, 1388462400, 1388466000, 1388469600, 1388473200, 
    1388476800, 1388480400, 1388484000, 1388487600, 1388491200, 1388494800, 
    1388498400, 1388502000, 1388505600, 1388509200, 1388512800, 1388516400, 
    1388520000, 1388523600, 1388527200, 1388530800, 1388534400, 1388538000, 
    1388541600, 1388545200, 1388548800, 1388552400, 1388556000, 1388559600, 
    1388563200, 1388566800, 1388570400, 1388574000, 1388577600, 1388581200, 
    1388584800, 1388588400, 1388592000, 1388595600, 1388599200, 1388602800, 
    1388606400, 1388610000, 1388613600, 1388617200, 1388620800, 1388624400, 
    1388628000, 1388631600, 1388635200, 1388638800, 1388642400, 1388646000, 
    1388649600, 1388653200, 1388656800, 1388660400, 1388664000, 1388667600, 
    1388671200, 1388674800, 1388678400, 1388682000, 1388685600, 1388689200, 
    1388692800, 1388696400, 1388700000, 1388703600, 1388707200, 1388710800, 
    1388714400, 1388718000, 1388721600, 1388725200, 1388728800, 1388732400, 
    1388736000, 1388739600, 1388743200, 1388746800, 1388750400, 1388754000, 
    1388757600, 1388761200, 1388764800, 1388768400, 1388772000, 1388775600, 
    1388779200, 1388782800, 1388786400, 1388790000, 1388793600, 1388797200, 
    1388800800, 1388804400, 1388808000, 1388811600, 1388815200, 1388818800, 
    1388822400, 1388826000, 1388829600, 1388833200, 1388836800, 1388840400, 
    1388844000, 1388847600, 1388851200, 1388854800, 1388858400, 1388862000, 
    1388865600, 1388869200, 1388872800, 1388876400, 1388880000, 1388883600, 
    1388887200, 1388890800, 1388894400, 1388898000, 1388901600, 1388905200, 
    1388908800, 1388912400, 1388916000, 1388919600, 1388923200, 1388926800, 
    1388930400, 1388934000, 1388937600, 1388941200, 1388944800, 1388948400, 
    1388952000, 1388955600, 1388959200, 1388962800, 1388966400, 1388970000, 
    1388973600, 1388977200, 1388980800, 1388984400, 1388988000, 1388991600, 
    1388995200, 1388998800, 1389002400, 1389006000, 1389009600, 1389013200, 
    1389016800, 1389020400, 1389024000, 1389027600, 1389031200, 1389034800, 
    1389038400, 1389042000, 1389045600, 1389049200, 1389052800, 1389056400, 
    1389060000, 1389063600, 1389067200, 1389070800, 1389074400, 1389078000, 
    1389081600, 1389085200, 1389088800, 1389092400, 1389096000, 1389099600, 
    1389103200, 1389106800, 1389110400, 1389114000, 1389117600, 1389121200, 
    1389124800, 1389128400, 1389132000, 1389135600, 1389139200, 1389142800, 
    1389146400, 1389150000, 1389153600, 1389157200, 1389160800, 1389164400, 
    1389168000, 1389171600, 1389175200, 1389178800, 1389182400, 1389186000, 
    1389189600, 1389193200, 1389196800, 1389200400, 1389204000, 1389207600, 
    1389211200, 1389214800, 1389218400, 1389222000, 1389225600, 1389229200, 
    1389232800, 1389236400, 1389240000, 1389243600, 1389247200, 1389250800, 
    1389254400, 1389258000, 1389261600, 1389265200, 1389268800, 1389272400, 
    1389276000, 1389279600, 1389283200, 1389286800, 1389290400, 1389294000, 
    1389297600, 1389301200, 1389304800, 1389308400, 1389312000, 1389315600, 
    1389319200, 1389322800, 1389326400, 1389330000, 1389333600, 1389337200, 
    1389340800, 1389344400, 1389348000, 1389351600, 1389355200, 1389358800, 
    1389362400, 1389366000, 1389369600, 1389373200, 1389376800, 1389380400, 
    1389384000, 1389387600, 1389391200, 1389394800, 1389398400, 1389402000, 
    1389405600, 1389409200, 1389412800, 1389416400, 1389420000, 1389423600, 
    1389427200, 1389430800, 1389434400, 1389438000, 1389441600, 1389445200, 
    1389448800, 1389452400, 1389456000, 1389459600, 1389463200, 1389466800, 
    1389470400, 1389474000, 1389477600, 1389481200, 1389484800, 1389488400, 
    1389492000, 1389495600, 1389499200, 1389502800, 1389506400, 1389510000, 
    1389513600, 1389517200, 1389520800, 1389524400, 1389528000, 1389531600, 
    1389535200, 1389538800, 1389542400, 1389546000, 1389549600, 1389553200, 
    1389556800, 1389560400, 1389564000, 1389567600, 1389571200, 1389574800, 
    1389578400, 1389582000, 1389585600, 1389589200, 1389592800, 1389596400, 
    1389600000, 1389603600, 1389607200, 1389610800, 1389614400, 1389618000, 
    1389621600, 1389625200, 1389628800, 1389632400, 1389636000, 1389639600, 
    1389643200, 1389646800, 1389650400, 1389654000, 1389657600, 1389661200, 
    1389664800, 1389668400, 1389672000, 1389675600, 1389679200, 1389682800, 
    1389686400, 1389690000, 1389693600, 1389697200, 1389700800, 1389704400, 
    1389708000, 1389711600, 1389715200, 1389718800, 1389722400, 1389726000, 
    1389729600, 1389733200, 1389736800, 1389740400, 1389744000, 1389747600, 
    1389751200, 1389754800, 1389758400, 1389762000, 1389765600, 1389769200, 
    1389772800, 1389776400, 1389780000, 1389783600, 1389787200, 1389790800, 
    1389794400, 1389798000, 1389801600, 1389805200, 1389808800, 1389812400, 
    1389816000, 1389819600, 1389823200, 1389826800, 1389830400, 1389834000, 
    1389837600, 1389841200, 1389844800, 1389848400, 1389852000, 1389855600, 
    1389859200, 1389862800, 1389866400, 1389870000, 1389873600, 1389877200, 
    1389880800, 1389884400, 1389888000, 1389891600, 1389895200, 1389898800, 
    1389902400, 1389906000, 1389909600, 1389913200, 1389916800, 1389920400, 
    1389924000, 1389927600, 1389931200, 1389934800, 1389938400, 1389942000, 
    1389945600, 1389949200, 1389952800, 1389956400, 1389960000, 1389963600, 
    1389967200, 1389970800, 1389974400, 1389978000, 1389981600, 1389985200, 
    1389988800, 1389992400, 1389996000, 1389999600, 1390003200, 1390006800, 
    1390010400, 1390014000, 1390017600, 1390021200, 1390024800, 1390028400, 
    1390032000, 1390035600, 1390039200, 1390042800, 1390046400, 1390050000, 
    1390053600, 1390057200, 1390060800, 1390064400, 1390068000, 1390071600, 
    1390075200, 1390078800, 1390082400, 1390086000, 1390089600, 1390093200, 
    1390096800, 1390100400, 1390104000, 1390107600, 1390111200, 1390114800, 
    1390118400, 1390122000, 1390125600, 1390129200, 1390132800, 1390136400, 
    1390140000, 1390143600, 1390147200, 1390150800, 1390154400, 1390158000, 
    1390161600, 1390165200, 1390168800, 1390172400, 1390176000, 1390179600, 
    1390183200, 1390186800, 1390190400, 1390194000, 1390197600, 1390201200, 
    1390204800, 1390208400, 1390212000, 1390215600, 1390219200, 1390222800, 
    1390226400, 1390230000, 1390233600, 1390237200, 1390240800, 1390244400, 
    1390248000, 1390251600, 1390255200, 1390258800, 1390262400, 1390266000, 
    1390269600, 1390273200, 1390276800, 1390280400, 1390284000, 1390287600, 
    1390291200, 1390294800, 1390298400, 1390302000, 1390305600, 1390309200, 
    1390312800, 1390316400, 1390320000, 1390323600, 1390327200, 1390330800, 
    1390334400, 1390338000, 1390341600, 1390345200, 1390348800, 1390352400, 
    1390356000, 1390359600, 1390363200, 1390366800, 1390370400, 1390374000, 
    1390377600, 1390381200, 1390384800, 1390388400, 1390392000, 1390395600, 
    1390399200, 1390402800, 1390406400, 1390410000, 1390413600, 1390417200, 
    1390420800, 1390424400, 1390428000, 1390431600, 1390435200, 1390438800, 
    1390442400, 1390446000, 1390449600, 1390453200, 1390456800, 1390460400, 
    1390464000, 1390467600, 1390471200, 1390474800, 1390478400, 1390482000, 
    1390485600, 1390489200, 1390492800, 1390496400, 1390500000, 1390503600, 
    1390507200, 1390510800, 1390514400, 1390518000, 1390521600, 1390525200, 
    1390528800, 1390532400, 1390536000, 1390539600, 1390543200, 1390546800, 
    1390550400, 1390554000, 1390557600, 1390561200, 1390564800, 1390568400, 
    1390572000, 1390575600, 1390579200, 1390582800, 1390586400, 1390590000, 
    1390593600, 1390597200, 1390600800, 1390604400, 1390608000, 1390611600, 
    1390615200, 1390618800, 1390622400, 1390626000, 1390629600, 1390633200, 
    1390636800, 1390640400, 1390644000, 1390647600, 1390651200, 1390654800, 
    1390658400, 1390662000, 1390665600, 1390669200, 1390672800, 1390676400, 
    1390680000, 1390683600, 1390687200, 1390690800, 1390694400, 1390698000, 
    1390701600, 1390705200, 1390708800, 1390712400, 1390716000, 1390719600, 
    1390723200, 1390726800, 1390730400, 1390734000, 1390737600, 1390741200, 
    1390744800, 1390748400, 1390752000, 1390755600, 1390759200, 1390762800, 
    1390766400, 1390770000, 1390773600, 1390777200, 1390780800, 1390784400, 
    1390788000, 1390791600, 1390795200, 1390798800, 1390802400, 1390806000, 
    1390809600, 1390813200, 1390816800, 1390820400, 1390824000, 1390827600, 
    1390831200, 1390834800, 1390838400, 1390842000, 1390845600, 1390849200, 
    1390852800, 1390856400, 1390860000, 1390863600, 1390867200, 1390870800, 
    1390874400, 1390878000, 1390881600, 1390885200, 1390888800, 1390892400, 
    1390896000, 1390899600, 1390903200, 1390906800, 1390910400, 1390914000, 
    1390917600, 1390921200, 1390924800, 1390928400, 1390932000, 1390935600, 
    1390939200, 1390942800, 1390946400, 1390950000, 1390953600, 1390957200, 
    1390960800, 1390964400, 1390968000, 1390971600, 1390975200, 1390978800, 
    1390982400, 1390986000, 1390989600, 1390993200, 1390996800, 1391000400, 
    1391004000, 1391007600, 1391011200, 1391014800, 1391018400, 1391022000, 
    1391025600, 1391029200, 1391032800, 1391036400, 1391040000, 1391043600, 
    1391047200, 1391050800, 1391054400, 1391058000, 1391061600, 1391065200, 
    1391068800, 1391072400, 1391076000, 1391079600, 1391083200, 1391086800, 
    1391090400, 1391094000, 1391097600, 1391101200, 1391104800, 1391108400, 
    1391112000, 1391115600, 1391119200, 1391122800, 1391126400, 1391130000, 
    1391133600, 1391137200, 1391140800, 1391144400, 1391148000, 1391151600, 
    1391155200, 1391158800, 1391162400, 1391166000, 1391169600, 1391173200, 
    1391176800, 1391180400, 1391184000, 1391187600, 1391191200, 1391194800, 
    1391198400, 1391202000, 1391205600, 1391209200, 1391212800, 1391216400, 
    1391220000, 1391223600, 1391227200, 1391230800, 1391234400, 1391238000, 
    1391241600, 1391245200, 1391248800, 1391252400, 1391256000, 1391259600, 
    1391263200, 1391266800, 1391270400, 1391274000, 1391277600, 1391281200, 
    1391284800, 1391288400, 1391292000, 1391295600, 1391299200, 1391302800, 
    1391306400, 1391310000, 1391313600, 1391317200, 1391320800, 1391324400, 
    1391328000, 1391331600, 1391335200, 1391338800, 1391342400, 1391346000, 
    1391349600, 1391353200, 1391356800, 1391360400, 1391364000, 1391367600, 
    1391371200, 1391374800, 1391378400, 1391382000, 1391385600, 1391389200, 
    1391392800, 1391396400, 1391400000, 1391403600, 1391407200, 1391410800, 
    1391414400, 1391418000, 1391421600, 1391425200, 1391428800, 1391432400, 
    1391436000, 1391439600, 1391443200, 1391446800, 1391450400, 1391454000, 
    1391457600, 1391461200, 1391464800, 1391468400, 1391472000, 1391475600, 
    1391479200, 1391482800, 1391486400, 1391490000, 1391493600, 1391497200, 
    1391500800, 1391504400, 1391508000, 1391511600, 1391515200, 1391518800, 
    1391522400, 1391526000, 1391529600, 1391533200, 1391536800, 1391540400, 
    1391544000, 1391547600, 1391551200, 1391554800, 1391558400, 1391562000, 
    1391565600, 1391569200, 1391572800, 1391576400, 1391580000, 1391583600, 
    1391587200, 1391590800, 1391594400, 1391598000, 1391601600, 1391605200, 
    1391608800, 1391612400, 1391616000, 1391619600, 1391623200, 1391626800, 
    1391630400, 1391634000, 1391637600, 1391641200, 1391644800, 1391648400, 
    1391652000, 1391655600, 1391659200, 1391662800, 1391666400, 1391670000, 
    1391673600, 1391677200, 1391680800, 1391684400, 1391688000, 1391691600, 
    1391695200, 1391698800, 1391702400, 1391706000, 1391709600, 1391713200, 
    1391716800, 1391720400, 1391724000, 1391727600, 1391731200, 1391734800, 
    1391738400, 1391742000, 1391745600, 1391749200, 1391752800, 1391756400, 
    1391760000, 1391763600, 1391767200, 1391770800, 1391774400, 1391778000, 
    1391781600, 1391785200, 1391788800, 1391792400, 1391796000, 1391799600, 
    1391803200, 1391806800, 1391810400, 1391814000, 1391817600, 1391821200, 
    1391824800, 1391828400, 1391832000, 1391835600, 1391839200, 1391842800, 
    1391846400, 1391850000, 1391853600, 1391857200, 1391860800, 1391864400, 
    1391868000, 1391871600, 1391875200, 1391878800, 1391882400, 1391886000, 
    1391889600, 1391893200, 1391896800, 1391900400, 1391904000, 1391907600, 
    1391911200, 1391914800, 1391918400, 1391922000, 1391925600, 1391929200, 
    1391932800, 1391936400, 1391940000, 1391943600, 1391947200, 1391950800, 
    1391954400, 1391958000, 1391961600, 1391965200, 1391968800, 1391972400, 
    1391976000, 1391979600, 1391983200, 1391986800, 1391990400, 1391994000, 
    1391997600, 1392001200, 1392004800, 1392008400, 1392012000, 1392015600, 
    1392019200, 1392022800, 1392026400, 1392030000, 1392033600, 1392037200, 
    1392040800, 1392044400, 1392048000, 1392051600, 1392055200, 1392058800, 
    1392062400, 1392066000, 1392069600, 1392073200, 1392076800, 1392080400, 
    1392084000, 1392087600, 1392091200, 1392094800, 1392098400, 1392102000, 
    1392105600, 1392109200, 1392112800, 1392116400, 1392120000, 1392123600, 
    1392127200, 1392130800, 1392134400, 1392138000, 1392141600, 1392145200, 
    1392148800, 1392152400, 1392156000, 1392159600, 1392163200, 1392166800, 
    1392170400, 1392174000, 1392177600, 1392181200, 1392184800, 1392188400, 
    1392192000, 1392195600, 1392199200, 1392202800, 1392206400, 1392210000, 
    1392213600, 1392217200, 1392220800, 1392224400, 1392228000, 1392231600, 
    1392235200, 1392238800, 1392242400, 1392246000, 1392249600, 1392253200, 
    1392256800, 1392260400, 1392264000, 1392267600, 1392271200, 1392274800, 
    1392278400, 1392282000, 1392285600, 1392289200, 1392292800, 1392296400, 
    1392300000, 1392303600, 1392307200, 1392310800, 1392314400, 1392318000, 
    1392321600, 1392325200, 1392328800, 1392332400, 1392336000, 1392339600, 
    1392343200, 1392346800, 1392350400, 1392354000, 1392357600, 1392361200, 
    1392364800, 1392368400, 1392372000, 1392375600, 1392379200, 1392382800, 
    1392386400, 1392390000, 1392393600, 1392397200, 1392400800, 1392404400, 
    1392408000, 1392411600, 1392415200, 1392418800, 1392422400, 1392426000, 
    1392429600, 1392433200, 1392436800, 1392440400, 1392444000, 1392447600, 
    1392451200, 1392454800, 1392458400, 1392462000, 1392465600, 1392469200, 
    1392472800, 1392476400, 1392480000, 1392483600, 1392487200, 1392490800, 
    1392494400, 1392498000, 1392501600, 1392505200, 1392508800, 1392512400, 
    1392516000, 1392519600, 1392523200, 1392526800, 1392530400, 1392534000, 
    1392537600, 1392541200, 1392544800, 1392548400, 1392552000, 1392555600, 
    1392559200, 1392562800, 1392566400, 1392570000, 1392573600, 1392577200, 
    1392580800, 1392584400, 1392588000, 1392591600, 1392595200, 1392598800, 
    1392602400, 1392606000, 1392609600, 1392613200, 1392616800, 1392620400, 
    1392624000, 1392627600, 1392631200, 1392634800, 1392638400, 1392642000, 
    1392645600, 1392649200, 1392652800, 1392656400, 1392660000, 1392663600, 
    1392667200, 1392670800, 1392674400, 1392678000, 1392681600, 1392685200, 
    1392688800, 1392692400, 1392696000, 1392699600, 1392703200, 1392706800, 
    1392710400, 1392714000, 1392717600, 1392721200, 1392724800, 1392728400, 
    1392732000, 1392735600, 1392739200, 1392742800, 1392746400, 1392750000, 
    1392753600, 1392757200, 1392760800, 1392764400, 1392768000, 1392771600, 
    1392775200, 1392778800, 1392782400, 1392786000, 1392789600, 1392793200, 
    1392796800, 1392800400, 1392804000, 1392807600, 1392811200, 1392814800, 
    1392818400, 1392822000, 1392825600, 1392829200, 1392832800, 1392836400, 
    1392840000, 1392843600, 1392847200, 1392850800, 1392854400, 1392858000, 
    1392861600, 1392865200, 1392868800, 1392872400, 1392876000, 1392879600, 
    1392883200, 1392886800, 1392890400, 1392894000, 1392897600, 1392901200, 
    1392904800, 1392908400, 1392912000, 1392915600, 1392919200, 1392922800, 
    1392926400, 1392930000, 1392933600, 1392937200, 1392940800, 1392944400, 
    1392948000, 1392951600, 1392955200, 1392958800, 1392962400, 1392966000, 
    1392969600, 1392973200, 1392976800, 1392980400, 1392984000, 1392987600, 
    1392991200, 1392994800, 1392998400, 1393002000, 1393005600, 1393009200, 
    1393012800, 1393016400, 1393020000, 1393023600, 1393027200, 1393030800, 
    1393034400, 1393038000, 1393041600, 1393045200, 1393048800, 1393052400, 
    1393056000, 1393059600, 1393063200, 1393066800, 1393070400, 1393074000, 
    1393077600, 1393081200, 1393084800, 1393088400, 1393092000, 1393095600, 
    1393099200, 1393102800, 1393106400, 1393110000, 1393113600, 1393117200, 
    1393120800, 1393124400, 1393128000, 1393131600, 1393135200, 1393138800, 
    1393142400, 1393146000, 1393149600, 1393153200, 1393156800, 1393160400, 
    1393164000, 1393167600, 1393171200, 1393174800, 1393178400, 1393182000, 
    1393185600, 1393189200, 1393192800, 1393196400, 1393200000, 1393203600, 
    1393207200, 1393210800, 1393214400, 1393218000, 1393221600, 1393225200, 
    1393228800, 1393232400, 1393236000, 1393239600, 1393243200, 1393246800, 
    1393250400, 1393254000, 1393257600, 1393261200, 1393264800, 1393268400, 
    1393272000, 1393275600, 1393279200, 1393282800, 1393286400, 1393290000, 
    1393293600, 1393297200, 1393300800, 1393304400, 1393308000, 1393311600, 
    1393315200, 1393318800, 1393322400, 1393326000, 1393329600, 1393333200, 
    1393336800, 1393340400, 1393344000, 1393347600, 1393351200, 1393354800, 
    1393358400, 1393362000, 1393365600, 1393369200, 1393372800, 1393376400, 
    1393380000, 1393383600, 1393387200, 1393390800, 1393394400, 1393398000, 
    1393401600, 1393405200, 1393408800, 1393412400, 1393416000, 1393419600, 
    1393423200, 1393426800, 1393430400, 1393434000, 1393437600, 1393441200, 
    1393444800, 1393448400, 1393452000, 1393455600, 1393459200, 1393462800, 
    1393466400, 1393470000, 1393473600, 1393477200, 1393480800, 1393484400, 
    1393488000, 1393491600, 1393495200, 1393498800, 1393502400, 1393506000, 
    1393509600, 1393513200, 1393516800, 1393520400, 1393524000, 1393527600, 
    1393531200, 1393534800, 1393538400, 1393542000, 1393545600, 1393549200, 
    1393552800, 1393556400, 1393560000, 1393563600, 1393567200, 1393570800, 
    1393574400, 1393578000, 1393581600, 1393585200, 1393588800, 1393592400, 
    1393596000, 1393599600, 1393603200, 1393606800, 1393610400, 1393614000, 
    1393617600, 1393621200, 1393624800, 1393628400, 1393632000, 1393635600, 
    1393639200, 1393642800, 1393646400, 1393650000, 1393653600, 1393657200, 
    1393660800, 1393664400, 1393668000, 1393671600, 1393675200, 1393678800, 
    1393682400, 1393686000, 1393689600, 1393693200, 1393696800, 1393700400, 
    1393704000, 1393707600, 1393711200, 1393714800, 1393718400, 1393722000, 
    1393725600, 1393729200, 1393732800, 1393736400, 1393740000, 1393743600, 
    1393747200, 1393750800, 1393754400, 1393758000, 1393761600, 1393765200, 
    1393768800, 1393772400, 1393776000, 1393779600, 1393783200, 1393786800, 
    1393790400, 1393794000, 1393797600, 1393801200, 1393804800, 1393808400, 
    1393812000, 1393815600, 1393819200, 1393822800, 1393826400, 1393830000, 
    1393833600, 1393837200, 1393840800, 1393844400, 1393848000, 1393851600, 
    1393855200, 1393858800, 1393862400, 1393866000, 1393869600, 1393873200, 
    1393876800, 1393880400, 1393884000, 1393887600, 1393891200, 1393894800, 
    1393898400, 1393902000, 1393905600, 1393909200, 1393912800, 1393916400, 
    1393920000, 1393923600, 1393927200, 1393930800, 1393934400, 1393938000, 
    1393941600, 1393945200, 1393948800, 1393952400, 1393956000, 1393959600, 
    1393963200, 1393966800, 1393970400, 1393974000, 1393977600, 1393981200, 
    1393984800, 1393988400, 1393992000, 1393995600, 1393999200, 1394002800, 
    1394006400, 1394010000, 1394013600, 1394017200, 1394020800, 1394024400, 
    1394028000, 1394031600, 1394035200, 1394038800, 1394042400, 1394046000, 
    1394049600, 1394053200, 1394056800, 1394060400, 1394064000, 1394067600, 
    1394071200, 1394074800, 1394078400, 1394082000, 1394085600, 1394089200, 
    1394092800, 1394096400, 1394100000, 1394103600, 1394107200, 1394110800, 
    1394114400, 1394118000, 1394121600, 1394125200, 1394128800, 1394132400, 
    1394136000, 1394139600, 1394143200, 1394146800, 1394150400, 1394154000, 
    1394157600, 1394161200, 1394164800, 1394168400, 1394172000, 1394175600, 
    1394179200, 1394182800, 1394186400, 1394190000, 1394193600, 1394197200, 
    1394200800, 1394204400, 1394208000, 1394211600, 1394215200, 1394218800, 
    1394222400, 1394226000, 1394229600, 1394233200, 1394236800, 1394240400, 
    1394244000, 1394247600, 1394251200, 1394254800, 1394258400, 1394262000, 
    1394265600, 1394269200, 1394272800, 1394276400, 1394280000, 1394283600, 
    1394287200, 1394290800, 1394294400, 1394298000, 1394301600, 1394305200, 
    1394308800, 1394312400, 1394316000, 1394319600, 1394323200, 1394326800, 
    1394330400, 1394334000, 1394337600, 1394341200, 1394344800, 1394348400, 
    1394352000, 1394355600, 1394359200, 1394362800, 1394366400, 1394370000, 
    1394373600, 1394377200, 1394380800, 1394384400, 1394388000, 1394391600, 
    1394395200, 1394398800, 1394402400, 1394406000, 1394409600, 1394413200, 
    1394416800, 1394420400, 1394424000, 1394427600, 1394431200, 1394434800, 
    1394438400, 1394442000, 1394445600, 1394449200, 1394452800, 1394456400, 
    1394460000, 1394463600, 1394467200, 1394470800, 1394474400, 1394478000, 
    1394481600, 1394485200, 1394488800, 1394492400, 1394496000, 1394499600, 
    1394503200, 1394506800, 1394510400, 1394514000, 1394517600, 1394521200, 
    1394524800, 1394528400, 1394532000, 1394535600, 1394539200, 1394542800, 
    1394546400, 1394550000, 1394553600, 1394557200, 1394560800, 1394564400, 
    1394568000, 1394571600, 1394575200, 1394578800, 1394582400, 1394586000, 
    1394589600, 1394593200, 1394596800, 1394600400, 1394604000, 1394607600, 
    1394611200, 1394614800, 1394618400, 1394622000, 1394625600, 1394629200, 
    1394632800, 1394636400, 1394640000, 1394643600, 1394647200, 1394650800, 
    1394654400, 1394658000, 1394661600, 1394665200, 1394668800, 1394672400, 
    1394676000, 1394679600, 1394683200, 1394686800, 1394690400, 1394694000, 
    1394697600, 1394701200, 1394704800, 1394708400, 1394712000, 1394715600, 
    1394719200, 1394722800, 1394726400, 1394730000, 1394733600, 1394737200, 
    1394740800, 1394744400, 1394748000, 1394751600, 1394755200, 1394758800, 
    1394762400, 1394766000, 1394769600, 1394773200, 1394776800, 1394780400, 
    1394784000, 1394787600, 1394791200, 1394794800, 1394798400, 1394802000, 
    1394805600, 1394809200, 1394812800, 1394816400, 1394820000, 1394823600, 
    1394827200, 1394830800, 1394834400, 1394838000, 1394841600, 1394845200, 
    1394848800, 1394852400, 1394856000, 1394859600, 1394863200, 1394866800, 
    1394870400, 1394874000, 1394877600, 1394881200, 1394884800, 1394888400, 
    1394892000, 1394895600, 1394899200, 1394902800, 1394906400, 1394910000, 
    1394913600, 1394917200, 1394920800, 1394924400, 1394928000, 1394931600, 
    1394935200, 1394938800, 1394942400, 1394946000, 1394949600, 1394953200, 
    1394956800, 1394960400, 1394964000, 1394967600, 1394971200, 1394974800, 
    1394978400, 1394982000, 1394985600, 1394989200, 1394992800, 1394996400, 
    1395000000, 1395003600, 1395007200, 1395010800, 1395014400, 1395018000, 
    1395021600, 1395025200, 1395028800, 1395032400, 1395036000, 1395039600, 
    1395043200, 1395046800, 1395050400, 1395054000, 1395057600, 1395061200, 
    1395064800, 1395068400, 1395072000, 1395075600, 1395079200, 1395082800, 
    1395086400, 1395090000, 1395093600, 1395097200, 1395100800, 1395104400, 
    1395108000, 1395111600, 1395115200, 1395118800, 1395122400, 1395126000, 
    1395129600, 1395133200, 1395136800, 1395140400, 1395144000, 1395147600, 
    1395151200, 1395154800, 1395158400, 1395162000, 1395165600, 1395169200, 
    1395172800, 1395176400, 1395180000, 1395183600, 1395187200, 1395190800, 
    1395194400, 1395198000, 1395201600, 1395205200, 1395208800, 1395212400, 
    1395216000, 1395219600, 1395223200, 1395226800, 1395230400, 1395234000, 
    1395237600, 1395241200, 1395244800, 1395248400, 1395252000, 1395255600, 
    1395259200, 1395262800, 1395266400, 1395270000, 1395273600, 1395277200, 
    1395280800, 1395284400, 1395288000, 1395291600, 1395295200, 1395298800, 
    1395302400, 1395306000, 1395309600, 1395313200, 1395316800, 1395320400, 
    1395324000, 1395327600, 1395331200, 1395334800, 1395338400, 1395342000, 
    1395345600, 1395349200, 1395352800, 1395356400, 1395360000, 1395363600, 
    1395367200, 1395370800, 1395374400, 1395378000, 1395381600, 1395385200, 
    1395388800, 1395392400, 1395396000, 1395399600, 1395403200, 1395406800, 
    1395410400, 1395414000, 1395417600, 1395421200, 1395424800, 1395428400, 
    1395432000, 1395435600, 1395439200, 1395442800, 1395446400, 1395450000, 
    1395453600, 1395457200, 1395460800, 1395464400, 1395468000, 1395471600, 
    1395475200, 1395478800, 1395482400, 1395486000, 1395489600, 1395493200, 
    1395496800, 1395500400, 1395504000, 1395507600, 1395511200, 1395514800, 
    1395518400, 1395522000, 1395525600, 1395529200, 1395532800, 1395536400, 
    1395540000, 1395543600, 1395547200, 1395550800, 1395554400, 1395558000, 
    1395561600, 1395565200, 1395568800, 1395572400, 1395576000, 1395579600, 
    1395583200, 1395586800, 1395590400, 1395594000, 1395597600, 1395601200, 
    1395604800, 1395608400, 1395612000, 1395615600, 1395619200, 1395622800, 
    1395626400, 1395630000, 1395633600, 1395637200, 1395640800, 1395644400, 
    1395648000, 1395651600, 1395655200, 1395658800, 1395662400, 1395666000, 
    1395669600, 1395673200, 1395676800, 1395680400, 1395684000, 1395687600, 
    1395691200, 1395694800, 1395698400, 1395702000, 1395705600, 1395709200, 
    1395712800, 1395716400, 1395720000, 1395723600, 1395727200, 1395730800, 
    1395734400, 1395738000, 1395741600, 1395745200, 1395748800, 1395752400, 
    1395756000, 1395759600, 1395763200, 1395766800, 1395770400, 1395774000, 
    1395777600, 1395781200, 1395784800, 1395788400, 1395792000, 1395795600, 
    1395799200, 1395802800, 1395806400, 1395810000, 1395813600, 1395817200, 
    1395820800, 1395824400, 1395828000, 1395831600, 1395835200, 1395838800, 
    1395842400, 1395846000, 1395849600, 1395853200, 1395856800, 1395860400, 
    1395864000, 1395867600, 1395871200, 1395874800, 1395878400, 1395882000, 
    1395885600, 1395889200, 1395892800, 1395896400, 1395900000, 1395903600, 
    1395907200, 1395910800, 1395914400, 1395918000, 1395921600, 1395925200, 
    1395928800, 1395932400, 1395936000, 1395939600, 1395943200, 1395946800, 
    1395950400, 1395954000, 1395957600, 1395961200, 1395964800, 1395968400, 
    1395972000, 1395975600, 1395979200, 1395982800, 1395986400, 1395990000, 
    1395993600, 1395997200, 1396000800, 1396004400, 1396008000, 1396011600, 
    1396015200, 1396018800, 1396022400, 1396026000, 1396029600, 1396033200, 
    1396036800, 1396040400, 1396044000, 1396047600, 1396051200, 1396054800, 
    1396058400, 1396062000, 1396065600, 1396069200, 1396072800, 1396076400, 
    1396080000, 1396083600, 1396087200, 1396090800, 1396094400, 1396098000, 
    1396101600, 1396105200, 1396108800, 1396112400, 1396116000, 1396119600, 
    1396123200, 1396126800, 1396130400, 1396134000, 1396137600, 1396141200, 
    1396144800, 1396148400, 1396152000, 1396155600, 1396159200, 1396162800, 
    1396166400, 1396170000, 1396173600, 1396177200, 1396180800, 1396184400, 
    1396188000, 1396191600, 1396195200, 1396198800, 1396202400, 1396206000, 
    1396209600, 1396213200, 1396216800, 1396220400, 1396224000, 1396227600, 
    1396231200, 1396234800, 1396238400, 1396242000, 1396245600, 1396249200, 
    1396252800, 1396256400, 1396260000, 1396263600, 1396267200, 1396270800, 
    1396274400, 1396278000, 1396281600, 1396285200, 1396288800, 1396292400, 
    1396296000, 1396299600, 1396303200, 1396306800, 1396310400, 1396314000, 
    1396317600, 1396321200, 1396324800, 1396328400, 1396332000, 1396335600, 
    1396339200, 1396342800, 1396346400, 1396350000, 1396353600, 1396357200, 
    1396360800, 1396364400, 1396368000, 1396371600, 1396375200, 1396378800, 
    1396382400, 1396386000, 1396389600, 1396393200, 1396396800, 1396400400, 
    1396404000, 1396407600, 1396411200, 1396414800, 1396418400, 1396422000, 
    1396425600, 1396429200, 1396432800, 1396436400, 1396440000, 1396443600, 
    1396447200, 1396450800, 1396454400, 1396458000, 1396461600, 1396465200, 
    1396468800, 1396472400, 1396476000, 1396479600, 1396483200, 1396486800, 
    1396490400, 1396494000, 1396497600, 1396501200, 1396504800, 1396508400, 
    1396512000, 1396515600, 1396519200, 1396522800, 1396526400, 1396530000, 
    1396533600, 1396537200, 1396540800, 1396544400, 1396548000, 1396551600, 
    1396555200, 1396558800, 1396562400, 1396566000, 1396569600, 1396573200, 
    1396576800, 1396580400, 1396584000, 1396587600, 1396591200, 1396594800, 
    1396598400, 1396602000, 1396605600, 1396609200, 1396612800, 1396616400, 
    1396620000, 1396623600, 1396627200, 1396630800, 1396634400, 1396638000, 
    1396641600, 1396645200, 1396648800, 1396652400, 1396656000, 1396659600, 
    1396663200, 1396666800, 1396670400, 1396674000, 1396677600, 1396681200, 
    1396684800, 1396688400, 1396692000, 1396695600, 1396699200, 1396702800, 
    1396706400, 1396710000, 1396713600, 1396717200, 1396720800, 1396724400, 
    1396728000, 1396731600, 1396735200, 1396738800, 1396742400, 1396746000, 
    1396749600, 1396753200, 1396756800, 1396760400, 1396764000, 1396767600, 
    1396771200, 1396774800, 1396778400, 1396782000, 1396785600, 1396789200, 
    1396792800, 1396796400, 1396800000, 1396803600, 1396807200, 1396810800, 
    1396814400, 1396818000, 1396821600, 1396825200, 1396828800, 1396832400, 
    1396836000, 1396839600, 1396843200, 1396846800, 1396850400, 1396854000, 
    1396857600, 1396861200, 1396864800, 1396868400, 1396872000, 1396875600, 
    1396879200, 1396882800, 1396886400, 1396890000, 1396893600, 1396897200, 
    1396900800, 1396904400, 1396908000, 1396911600, 1396915200, 1396918800, 
    1396922400, 1396926000, 1396929600, 1396933200, 1396936800, 1396940400, 
    1396944000, 1396947600, 1396951200, 1396954800, 1396958400, 1396962000, 
    1396965600, 1396969200, 1396972800, 1396976400, 1396980000, 1396983600, 
    1396987200, 1396990800, 1396994400, 1396998000, 1397001600, 1397005200, 
    1397008800, 1397012400, 1397016000, 1397019600, 1397023200, 1397026800, 
    1397030400, 1397034000, 1397037600, 1397041200, 1397044800, 1397048400, 
    1397052000, 1397055600, 1397059200, 1397062800, 1397066400, 1397070000, 
    1397073600, 1397077200, 1397080800, 1397084400, 1397088000, 1397091600, 
    1397095200, 1397098800, 1397102400, 1397106000, 1397109600, 1397113200, 
    1397116800, 1397120400, 1397124000, 1397127600, 1397131200, 1397134800, 
    1397138400, 1397142000, 1397145600, 1397149200, 1397152800, 1397156400, 
    1397160000, 1397163600, 1397167200, 1397170800, 1397174400, 1397178000, 
    1397181600, 1397185200, 1397188800, 1397192400, 1397196000, 1397199600, 
    1397203200, 1397206800, 1397210400, 1397214000, 1397217600, 1397221200, 
    1397224800, 1397228400, 1397232000, 1397235600, 1397239200, 1397242800, 
    1397246400, 1397250000, 1397253600, 1397257200, 1397260800, 1397264400, 
    1397268000, 1397271600, 1397275200, 1397278800, 1397282400, 1397286000, 
    1397289600, 1397293200, 1397296800, 1397300400, 1397304000, 1397307600, 
    1397311200, 1397314800, 1397318400, 1397322000, 1397325600, 1397329200, 
    1397332800, 1397336400, 1397340000, 1397343600, 1397347200, 1397350800, 
    1397354400, 1397358000, 1397361600, 1397365200, 1397368800, 1397372400, 
    1397376000, 1397379600, 1397383200, 1397386800, 1397390400, 1397394000, 
    1397397600, 1397401200, 1397404800, 1397408400, 1397412000, 1397415600, 
    1397419200, 1397422800, 1397426400, 1397430000, 1397433600, 1397437200, 
    1397440800, 1397444400, 1397448000, 1397451600, 1397455200, 1397458800, 
    1397462400, 1397466000, 1397469600, 1397473200, 1397476800, 1397480400, 
    1397484000, 1397487600, 1397491200, 1397494800, 1397498400, 1397502000, 
    1397505600, 1397509200, 1397512800, 1397516400, 1397520000, 1397523600, 
    1397527200, 1397530800, 1397534400, 1397538000, 1397541600, 1397545200, 
    1397548800, 1397552400, 1397556000, 1397559600, 1397563200, 1397566800, 
    1397570400, 1397574000, 1397577600, 1397581200, 1397584800, 1397588400, 
    1397592000, 1397595600, 1397599200, 1397602800, 1397606400, 1397610000, 
    1397613600, 1397617200, 1397620800, 1397624400, 1397628000, 1397631600, 
    1397635200, 1397638800, 1397642400, 1397646000, 1397649600, 1397653200, 
    1397656800, 1397660400, 1397664000, 1397667600, 1397671200, 1397674800, 
    1397678400, 1397682000, 1397685600, 1397689200, 1397692800, 1397696400, 
    1397700000, 1397703600, 1397707200, 1397710800, 1397714400, 1397718000, 
    1397721600, 1397725200, 1397728800, 1397732400, 1397736000, 1397739600, 
    1397743200, 1397746800, 1397750400, 1397754000, 1397757600, 1397761200, 
    1397764800, 1397768400, 1397772000, 1397775600, 1397779200, 1397782800, 
    1397786400, 1397790000, 1397793600, 1397797200, 1397800800, 1397804400, 
    1397808000, 1397811600, 1397815200, 1397818800, 1397822400, 1397826000, 
    1397829600, 1397833200, 1397836800, 1397840400, 1397844000, 1397847600, 
    1397851200, 1397854800, 1397858400, 1397862000, 1397865600, 1397869200, 
    1397872800, 1397876400, 1397880000, 1397883600, 1397887200, 1397890800, 
    1397894400, 1397898000, 1397901600, 1397905200, 1397908800, 1397912400, 
    1397916000, 1397919600, 1397923200, 1397926800, 1397930400, 1397934000, 
    1397937600, 1397941200, 1397944800, 1397948400, 1397952000, 1397955600, 
    1397959200, 1397962800, 1397966400, 1397970000, 1397973600, 1397977200, 
    1397980800, 1397984400, 1397988000, 1397991600, 1397995200, 1397998800, 
    1398002400, 1398006000, 1398009600, 1398013200, 1398016800, 1398020400, 
    1398024000, 1398027600, 1398031200, 1398034800, 1398038400, 1398042000, 
    1398045600, 1398049200, 1398052800, 1398056400, 1398060000, 1398063600, 
    1398067200, 1398070800, 1398074400, 1398078000, 1398081600, 1398085200, 
    1398088800, 1398092400, 1398096000, 1398099600, 1398103200, 1398106800, 
    1398110400, 1398114000, 1398117600, 1398121200, 1398124800, 1398128400, 
    1398132000, 1398135600, 1398139200, 1398142800, 1398146400, 1398150000, 
    1398153600, 1398157200, 1398160800, 1398164400, 1398168000, 1398171600, 
    1398175200, 1398178800, 1398182400, 1398186000, 1398189600, 1398193200, 
    1398196800, 1398200400, 1398204000, 1398207600, 1398211200, 1398214800, 
    1398218400, 1398222000, 1398225600, 1398229200, 1398232800, 1398236400, 
    1398240000, 1398243600, 1398247200, 1398250800, 1398254400, 1398258000, 
    1398261600, 1398265200, 1398268800, 1398272400, 1398276000, 1398279600, 
    1398283200, 1398286800, 1398290400, 1398294000, 1398297600, 1398301200, 
    1398304800, 1398308400, 1398312000, 1398315600, 1398319200, 1398322800, 
    1398326400, 1398330000, 1398333600, 1398337200, 1398340800, 1398344400, 
    1398348000, 1398351600, 1398355200, 1398358800, 1398362400, 1398366000, 
    1398369600, 1398373200, 1398376800, 1398380400, 1398384000, 1398387600, 
    1398391200, 1398394800, 1398398400, 1398402000, 1398405600, 1398409200, 
    1398412800, 1398416400, 1398420000, 1398423600, 1398427200, 1398430800, 
    1398434400, 1398438000, 1398441600, 1398445200, 1398448800, 1398452400, 
    1398456000, 1398459600, 1398463200, 1398466800, 1398470400, 1398474000, 
    1398477600, 1398481200, 1398484800, 1398488400, 1398492000, 1398495600, 
    1398499200, 1398502800, 1398506400, 1398510000, 1398513600, 1398517200, 
    1398520800, 1398524400, 1398528000, 1398531600, 1398535200, 1398538800, 
    1398542400, 1398546000, 1398549600, 1398553200, 1398556800, 1398560400, 
    1398564000, 1398567600, 1398571200, 1398574800, 1398578400, 1398582000, 
    1398585600, 1398589200, 1398592800, 1398596400, 1398600000, 1398603600, 
    1398607200, 1398610800, 1398614400, 1398618000, 1398621600, 1398625200, 
    1398628800, 1398632400, 1398636000, 1398639600, 1398643200, 1398646800, 
    1398650400, 1398654000, 1398657600, 1398661200, 1398664800, 1398668400, 
    1398672000, 1398675600, 1398679200, 1398682800, 1398686400, 1398690000, 
    1398693600, 1398697200, 1398700800, 1398704400, 1398708000, 1398711600, 
    1398715200, 1398718800, 1398722400, 1398726000, 1398729600, 1398733200, 
    1398736800, 1398740400, 1398744000, 1398747600, 1398751200, 1398754800, 
    1398758400, 1398762000, 1398765600, 1398769200, 1398772800, 1398776400, 
    1398780000, 1398783600, 1398787200, 1398790800, 1398794400, 1398798000, 
    1398801600, 1398805200, 1398808800, 1398812400, 1398816000, 1398819600, 
    1398823200, 1398826800, 1398830400, 1398834000, 1398837600, 1398841200, 
    1398844800, 1398848400, 1398852000, 1398855600, 1398859200, 1398862800, 
    1398866400, 1398870000, 1398873600, 1398877200, 1398880800, 1398884400, 
    1398888000, 1398891600, 1398895200, 1398898800, 1398902400, 1398906000, 
    1398909600, 1398913200, 1398916800, 1398920400, 1398924000, 1398927600, 
    1398931200, 1398934800, 1398938400, 1398942000, 1398945600, 1398949200, 
    1398952800, 1398956400, 1398960000, 1398963600, 1398967200, 1398970800, 
    1398974400, 1398978000, 1398981600, 1398985200, 1398988800, 1398992400, 
    1398996000, 1398999600, 1399003200, 1399006800, 1399010400, 1399014000, 
    1399017600, 1399021200, 1399024800, 1399028400, 1399032000, 1399035600, 
    1399039200, 1399042800, 1399046400, 1399050000, 1399053600, 1399057200, 
    1399060800, 1399064400, 1399068000, 1399071600, 1399075200, 1399078800, 
    1399082400, 1399086000, 1399089600, 1399093200, 1399096800, 1399100400, 
    1399104000, 1399107600, 1399111200, 1399114800, 1399118400, 1399122000, 
    1399125600, 1399129200, 1399132800, 1399136400, 1399140000, 1399143600, 
    1399147200, 1399150800, 1399154400, 1399158000, 1399161600, 1399165200, 
    1399168800, 1399172400, 1399176000, 1399179600, 1399183200, 1399186800, 
    1399190400, 1399194000, 1399197600, 1399201200, 1399204800, 1399208400, 
    1399212000, 1399215600, 1399219200, 1399222800, 1399226400, 1399230000, 
    1399233600, 1399237200, 1399240800, 1399244400, 1399248000, 1399251600, 
    1399255200, 1399258800, 1399262400, 1399266000, 1399269600, 1399273200, 
    1399276800, 1399280400, 1399284000, 1399287600, 1399291200, 1399294800, 
    1399298400, 1399302000, 1399305600, 1399309200, 1399312800, 1399316400, 
    1399320000, 1399323600, 1399327200, 1399330800, 1399334400, 1399338000, 
    1399341600, 1399345200, 1399348800, 1399352400, 1399356000, 1399359600, 
    1399363200, 1399366800, 1399370400, 1399374000, 1399377600, 1399381200, 
    1399384800, 1399388400, 1399392000, 1399395600, 1399399200, 1399402800, 
    1399406400, 1399410000, 1399413600, 1399417200, 1399420800, 1399424400, 
    1399428000, 1399431600, 1399435200, 1399438800, 1399442400, 1399446000, 
    1399449600, 1399453200, 1399456800, 1399460400, 1399464000, 1399467600, 
    1399471200, 1399474800, 1399478400, 1399482000, 1399485600, 1399489200, 
    1399492800, 1399496400, 1399500000, 1399503600, 1399507200, 1399510800, 
    1399514400, 1399518000, 1399521600, 1399525200, 1399528800, 1399532400, 
    1399536000, 1399539600, 1399543200, 1399546800, 1399550400, 1399554000, 
    1399557600, 1399561200, 1399564800, 1399568400, 1399572000, 1399575600, 
    1399579200, 1399582800, 1399586400, 1399590000, 1399593600, 1399597200, 
    1399600800, 1399604400, 1399608000, 1399611600, 1399615200, 1399618800, 
    1399622400, 1399626000, 1399629600, 1399633200, 1399636800, 1399640400, 
    1399644000, 1399647600, 1399651200, 1399654800, 1399658400, 1399662000, 
    1399665600, 1399669200, 1399672800, 1399676400, 1399680000, 1399683600, 
    1399687200, 1399690800, 1399694400, 1399698000, 1399701600, 1399705200, 
    1399708800, 1399712400, 1399716000, 1399719600, 1399723200, 1399726800, 
    1399730400, 1399734000, 1399737600, 1399741200, 1399744800, 1399748400, 
    1399752000, 1399755600, 1399759200, 1399762800, 1399766400, 1399770000, 
    1399773600, 1399777200, 1399780800, 1399784400, 1399788000, 1399791600, 
    1399795200, 1399798800, 1399802400, 1399806000, 1399809600, 1399813200, 
    1399816800, 1399820400, 1399824000, 1399827600, 1399831200, 1399834800, 
    1399838400, 1399842000, 1399845600, 1399849200, 1399852800, 1399856400, 
    1399860000, 1399863600, 1399867200, 1399870800, 1399874400, 1399878000, 
    1399881600, 1399885200, 1399888800, 1399892400, 1399896000, 1399899600, 
    1399903200, 1399906800, 1399910400, 1399914000, 1399917600, 1399921200, 
    1399924800, 1399928400, 1399932000, 1399935600, 1399939200, 1399942800, 
    1399946400, 1399950000, 1399953600, 1399957200, 1399960800, 1399964400, 
    1399968000, 1399971600, 1399975200, 1399978800, 1399982400, 1399986000, 
    1399989600, 1399993200, 1399996800, 1400000400, 1400004000, 1400007600, 
    1400011200, 1400014800, 1400018400, 1400022000, 1400025600, 1400029200, 
    1400032800, 1400036400, 1400040000, 1400043600, 1400047200, 1400050800, 
    1400054400, 1400058000, 1400061600, 1400065200, 1400068800, 1400072400, 
    1400076000, 1400079600, 1400083200, 1400086800, 1400090400, 1400094000, 
    1400097600, 1400101200, 1400104800, 1400108400, 1400112000, 1400115600, 
    1400119200, 1400122800, 1400126400, 1400130000, 1400133600, 1400137200, 
    1400140800, 1400144400, 1400148000, 1400151600, 1400155200, 1400158800, 
    1400162400, 1400166000, 1400169600, 1400173200, 1400176800, 1400180400, 
    1400184000, 1400187600, 1400191200, 1400194800, 1400198400, 1400202000, 
    1400205600, 1400209200, 1400212800, 1400216400, 1400220000, 1400223600, 
    1400227200, 1400230800, 1400234400, 1400238000, 1400241600, 1400245200, 
    1400248800, 1400252400, 1400256000, 1400259600, 1400263200, 1400266800, 
    1400270400, 1400274000, 1400277600, 1400281200, 1400284800, 1400288400, 
    1400292000, 1400295600, 1400299200, 1400302800, 1400306400, 1400310000, 
    1400313600, 1400317200, 1400320800, 1400324400, 1400328000, 1400331600, 
    1400335200, 1400338800, 1400342400, 1400346000, 1400349600, 1400353200, 
    1400356800, 1400360400, 1400364000, 1400367600, 1400371200, 1400374800, 
    1400378400, 1400382000, 1400385600, 1400389200, 1400392800, 1400396400, 
    1400400000, 1400403600, 1400407200, 1400410800, 1400414400, 1400418000, 
    1400421600, 1400425200, 1400428800, 1400432400, 1400436000, 1400439600, 
    1400443200, 1400446800, 1400450400, 1400454000, 1400457600, 1400461200, 
    1400464800, 1400468400, 1400472000, 1400475600, 1400479200, 1400482800, 
    1400486400, 1400490000, 1400493600, 1400497200, 1400500800, 1400504400, 
    1400508000, 1400511600, 1400515200, 1400518800, 1400522400, 1400526000, 
    1400529600, 1400533200, 1400536800, 1400540400, 1400544000, 1400547600, 
    1400551200, 1400554800, 1400558400, 1400562000, 1400565600, 1400569200, 
    1400572800, 1400576400, 1400580000, 1400583600, 1400587200, 1400590800, 
    1400594400, 1400598000, 1400601600, 1400605200, 1400608800, 1400612400, 
    1400616000, 1400619600, 1400623200, 1400626800, 1400630400, 1400634000, 
    1400637600, 1400641200, 1400644800, 1400648400, 1400652000, 1400655600, 
    1400659200, 1400662800, 1400666400, 1400670000, 1400673600, 1400677200, 
    1400680800, 1400684400, 1400688000, 1400691600, 1400695200, 1400698800, 
    1400702400, 1400706000, 1400709600, 1400713200, 1400716800, 1400720400, 
    1400724000, 1400727600, 1400731200, 1400734800, 1400738400, 1400742000, 
    1400745600, 1400749200, 1400752800, 1400756400, 1400760000, 1400763600, 
    1400767200, 1400770800, 1400774400, 1400778000, 1400781600, 1400785200, 
    1400788800, 1400792400, 1400796000, 1400799600, 1400803200, 1400806800, 
    1400810400, 1400814000, 1400817600, 1400821200, 1400824800, 1400828400, 
    1400832000, 1400835600, 1400839200, 1400842800, 1400846400, 1400850000, 
    1400853600, 1400857200, 1400860800, 1400864400, 1400868000, 1400871600, 
    1400875200, 1400878800, 1400882400, 1400886000, 1400889600, 1400893200, 
    1400896800, 1400900400, 1400904000, 1400907600, 1400911200, 1400914800, 
    1400918400, 1400922000, 1400925600, 1400929200, 1400932800, 1400936400, 
    1400940000, 1400943600, 1400947200, 1400950800, 1400954400, 1400958000, 
    1400961600, 1400965200, 1400968800, 1400972400, 1400976000, 1400979600, 
    1400983200, 1400986800, 1400990400, 1400994000, 1400997600, 1401001200, 
    1401004800, 1401008400, 1401012000, 1401015600, 1401019200, 1401022800, 
    1401026400, 1401030000, 1401033600, 1401037200, 1401040800, 1401044400, 
    1401048000, 1401051600, 1401055200, 1401058800, 1401062400, 1401066000, 
    1401069600, 1401073200, 1401076800, 1401080400, 1401084000, 1401087600, 
    1401091200, 1401094800, 1401098400, 1401102000, 1401105600, 1401109200, 
    1401112800, 1401116400, 1401120000, 1401123600, 1401127200, 1401130800, 
    1401134400, 1401138000, 1401141600, 1401145200, 1401148800, 1401152400, 
    1401156000, 1401159600, 1401163200, 1401166800, 1401170400, 1401174000, 
    1401177600, 1401181200, 1401184800, 1401188400, 1401192000, 1401195600, 
    1401199200, 1401202800, 1401206400, 1401210000, 1401213600, 1401217200, 
    1401220800, 1401224400, 1401228000, 1401231600, 1401235200, 1401238800, 
    1401242400, 1401246000, 1401249600, 1401253200, 1401256800, 1401260400, 
    1401264000, 1401267600, 1401271200, 1401274800, 1401278400, 1401282000, 
    1401285600, 1401289200, 1401292800, 1401296400, 1401300000, 1401303600, 
    1401307200, 1401310800, 1401314400, 1401318000, 1401321600, 1401325200, 
    1401328800, 1401332400, 1401336000, 1401339600, 1401343200, 1401346800, 
    1401350400, 1401354000, 1401357600, 1401361200, 1401364800, 1401368400, 
    1401372000, 1401375600, 1401379200, 1401382800, 1401386400, 1401390000, 
    1401393600, 1401397200, 1401400800, 1401404400, 1401408000, 1401411600, 
    1401415200, 1401418800, 1401422400, 1401426000, 1401429600, 1401433200, 
    1401436800, 1401440400, 1401444000, 1401447600, 1401451200, 1401454800, 
    1401458400, 1401462000, 1401465600, 1401469200, 1401472800, 1401476400, 
    1401480000, 1401483600, 1401487200, 1401490800, 1401494400, 1401498000, 
    1401501600, 1401505200, 1401508800, 1401512400, 1401516000, 1401519600, 
    1401523200, 1401526800, 1401530400, 1401534000, 1401537600, 1401541200, 
    1401544800, 1401548400, 1401552000, 1401555600, 1401559200, 1401562800, 
    1401566400, 1401570000, 1401573600, 1401577200, 1401580800, 1401584400, 
    1401588000, 1401591600, 1401595200, 1401598800, 1401602400, 1401606000, 
    1401609600, 1401613200, 1401616800, 1401620400, 1401624000, 1401627600, 
    1401631200, 1401634800, 1401638400, 1401642000, 1401645600, 1401649200, 
    1401652800, 1401656400, 1401660000, 1401663600, 1401667200, 1401670800, 
    1401674400, 1401678000, 1401681600, 1401685200, 1401688800, 1401692400, 
    1401696000, 1401699600, 1401703200, 1401706800, 1401710400, 1401714000, 
    1401717600, 1401721200, 1401724800, 1401728400, 1401732000, 1401735600, 
    1401739200, 1401742800, 1401746400, 1401750000, 1401753600, 1401757200, 
    1401760800, 1401764400, 1401768000, 1401771600, 1401775200, 1401778800, 
    1401782400, 1401786000, 1401789600, 1401793200, 1401796800, 1401800400, 
    1401804000, 1401807600, 1401811200, 1401814800, 1401818400, 1401822000, 
    1401825600, 1401829200, 1401832800, 1401836400, 1401840000, 1401843600, 
    1401847200, 1401850800, 1401854400, 1401858000, 1401861600, 1401865200, 
    1401868800, 1401872400, 1401876000, 1401879600, 1401883200, 1401886800, 
    1401890400, 1401894000, 1401897600, 1401901200, 1401904800, 1401908400, 
    1401912000, 1401915600, 1401919200, 1401922800, 1401926400, 1401930000, 
    1401933600, 1401937200, 1401940800, 1401944400, 1401948000, 1401951600, 
    1401955200, 1401958800, 1401962400, 1401966000, 1401969600, 1401973200, 
    1401976800, 1401980400, 1401984000, 1401987600, 1401991200, 1401994800, 
    1401998400, 1402002000, 1402005600, 1402009200, 1402012800, 1402016400, 
    1402020000, 1402023600, 1402027200, 1402030800, 1402034400, 1402038000, 
    1402041600, 1402045200, 1402048800, 1402052400, 1402056000, 1402059600, 
    1402063200, 1402066800, 1402070400, 1402074000, 1402077600, 1402081200, 
    1402084800, 1402088400, 1402092000, 1402095600, 1402099200, 1402102800, 
    1402106400, 1402110000, 1402113600, 1402117200, 1402120800, 1402124400, 
    1402128000, 1402131600, 1402135200, 1402138800, 1402142400, 1402146000, 
    1402149600, 1402153200, 1402156800, 1402160400, 1402164000, 1402167600, 
    1402171200, 1402174800, 1402178400, 1402182000, 1402185600, 1402189200, 
    1402192800, 1402196400, 1402200000, 1402203600, 1402207200, 1402210800, 
    1402214400, 1402218000, 1402221600, 1402225200, 1402228800, 1402232400, 
    1402236000, 1402239600, 1402243200, 1402246800, 1402250400, 1402254000, 
    1402257600, 1402261200, 1402264800, 1402268400, 1402272000, 1402275600, 
    1402279200, 1402282800, 1402286400, 1402290000, 1402293600, 1402297200, 
    1402300800, 1402304400, 1402308000, 1402311600, 1402315200, 1402318800, 
    1402322400, 1402326000, 1402329600, 1402333200, 1402336800, 1402340400, 
    1402344000, 1402347600, 1402351200, 1402354800, 1402358400, 1402362000, 
    1402365600, 1402369200, 1402372800, 1402376400, 1402380000, 1402383600, 
    1402387200, 1402390800, 1402394400, 1402398000, 1402401600, 1402405200, 
    1402408800, 1402412400, 1402416000, 1402419600, 1402423200, 1402426800, 
    1402430400, 1402434000, 1402437600, 1402441200, 1402444800, 1402448400, 
    1402452000, 1402455600, 1402459200, 1402462800, 1402466400, 1402470000, 
    1402473600, 1402477200, 1402480800, 1402484400, 1402488000, 1402491600, 
    1402495200, 1402498800, 1402502400, 1402506000, 1402509600, 1402513200, 
    1402516800, 1402520400, 1402524000, 1402527600, 1402531200, 1402534800, 
    1402538400, 1402542000, 1402545600, 1402549200, 1402552800, 1402556400, 
    1402560000, 1402563600, 1402567200, 1402570800, 1402574400, 1402578000, 
    1402581600, 1402585200, 1402588800, 1402592400, 1402596000, 1402599600, 
    1402603200, 1402606800, 1402610400, 1402614000, 1402617600, 1402621200, 
    1402624800, 1402628400, 1402632000, 1402635600, 1402639200, 1402642800, 
    1402646400, 1402650000, 1402653600, 1402657200, 1402660800, 1402664400, 
    1402668000, 1402671600, 1402675200, 1402678800, 1402682400, 1402686000, 
    1402689600, 1402693200, 1402696800, 1402700400, 1402704000, 1402707600, 
    1402711200, 1402714800, 1402718400, 1402722000, 1402725600, 1402729200, 
    1402732800, 1402736400, 1402740000, 1402743600, 1402747200, 1402750800, 
    1402754400, 1402758000, 1402761600, 1402765200, 1402768800, 1402772400, 
    1402776000, 1402779600, 1402783200, 1402786800, 1402790400, 1402794000, 
    1402797600, 1402801200, 1402804800, 1402808400, 1402812000, 1402815600, 
    1402819200, 1402822800, 1402826400, 1402830000, 1402833600, 1402837200, 
    1402840800, 1402844400, 1402848000, 1402851600, 1402855200, 1402858800, 
    1402862400, 1402866000, 1402869600, 1402873200, 1402876800, 1402880400, 
    1402884000, 1402887600, 1402891200, 1402894800, 1402898400, 1402902000, 
    1402905600, 1402909200, 1402912800, 1402916400, 1402920000, 1402923600, 
    1402927200, 1402930800, 1402934400, 1402938000, 1402941600, 1402945200, 
    1402948800, 1402952400, 1402956000, 1402959600, 1402963200, 1402966800, 
    1402970400, 1402974000, 1402977600, 1402981200, 1402984800, 1402988400, 
    1402992000, 1402995600, 1402999200, 1403002800, 1403006400, 1403010000, 
    1403013600, 1403017200, 1403020800, 1403024400, 1403028000, 1403031600, 
    1403035200, 1403038800, 1403042400, 1403046000, 1403049600, 1403053200, 
    1403056800, 1403060400, 1403064000, 1403067600, 1403071200, 1403074800, 
    1403078400, 1403082000, 1403085600, 1403089200, 1403092800, 1403096400, 
    1403100000, 1403103600, 1403107200, 1403110800, 1403114400, 1403118000, 
    1403121600, 1403125200, 1403128800, 1403132400, 1403136000, 1403139600, 
    1403143200, 1403146800, 1403150400, 1403154000, 1403157600, 1403161200, 
    1403164800, 1403168400, 1403172000, 1403175600, 1403179200, 1403182800, 
    1403186400, 1403190000, 1403193600, 1403197200, 1403200800, 1403204400, 
    1403208000, 1403211600, 1403215200, 1403218800, 1403222400, 1403226000, 
    1403229600, 1403233200, 1403236800, 1403240400, 1403244000, 1403247600, 
    1403251200, 1403254800, 1403258400, 1403262000, 1403265600, 1403269200, 
    1403272800, 1403276400, 1403280000, 1403283600, 1403287200, 1403290800, 
    1403294400, 1403298000, 1403301600, 1403305200, 1403308800, 1403312400, 
    1403316000, 1403319600, 1403323200, 1403326800, 1403330400, 1403334000, 
    1403337600, 1403341200, 1403344800, 1403348400, 1403352000, 1403355600, 
    1403359200, 1403362800, 1403366400, 1403370000, 1403373600, 1403377200, 
    1403380800, 1403384400, 1403388000, 1403391600, 1403395200, 1403398800, 
    1403402400, 1403406000, 1403409600, 1403413200, 1403416800, 1403420400, 
    1403424000, 1403427600, 1403431200, 1403434800, 1403438400, 1403442000, 
    1403445600, 1403449200, 1403452800, 1403456400, 1403460000, 1403463600, 
    1403467200, 1403470800, 1403474400, 1403478000, 1403481600, 1403485200, 
    1403488800, 1403492400, 1403496000, 1403499600, 1403503200, 1403506800, 
    1403510400, 1403514000, 1403517600, 1403521200, 1403524800, 1403528400, 
    1403532000, 1403535600, 1403539200, 1403542800, 1403546400, 1403550000, 
    1403553600, 1403557200, 1403560800, 1403564400, 1403568000, 1403571600, 
    1403575200, 1403578800, 1403582400, 1403586000, 1403589600, 1403593200, 
    1403596800, 1403600400, 1403604000, 1403607600, 1403611200, 1403614800, 
    1403618400, 1403622000, 1403625600, 1403629200, 1403632800, 1403636400, 
    1403640000, 1403643600, 1403647200, 1403650800, 1403654400, 1403658000, 
    1403661600, 1403665200, 1403668800, 1403672400, 1403676000, 1403679600, 
    1403683200, 1403686800, 1403690400, 1403694000, 1403697600, 1403701200, 
    1403704800, 1403708400, 1403712000, 1403715600, 1403719200, 1403722800, 
    1403726400, 1403730000, 1403733600, 1403737200, 1403740800, 1403744400, 
    1403748000, 1403751600, 1403755200, 1403758800, 1403762400, 1403766000, 
    1403769600, 1403773200, 1403776800, 1403780400, 1403784000, 1403787600, 
    1403791200, 1403794800, 1403798400, 1403802000, 1403805600, 1403809200, 
    1403812800, 1403816400, 1403820000, 1403823600, 1403827200, 1403830800, 
    1403834400, 1403838000, 1403841600, 1403845200, 1403848800, 1403852400, 
    1403856000, 1403859600, 1403863200, 1403866800, 1403870400, 1403874000, 
    1403877600, 1403881200, 1403884800, 1403888400, 1403892000, 1403895600, 
    1403899200, 1403902800, 1403906400, 1403910000, 1403913600, 1403917200, 
    1403920800, 1403924400, 1403928000, 1403931600, 1403935200, 1403938800, 
    1403942400, 1403946000, 1403949600, 1403953200, 1403956800, 1403960400, 
    1403964000, 1403967600, 1403971200, 1403974800, 1403978400, 1403982000, 
    1403985600, 1403989200, 1403992800, 1403996400, 1404000000, 1404003600, 
    1404007200, 1404010800, 1404014400, 1404018000, 1404021600, 1404025200, 
    1404028800, 1404032400, 1404036000, 1404039600, 1404043200, 1404046800, 
    1404050400, 1404054000, 1404057600, 1404061200, 1404064800, 1404068400, 
    1404072000, 1404075600, 1404079200, 1404082800, 1404086400, 1404090000, 
    1404093600, 1404097200, 1404100800, 1404104400, 1404108000, 1404111600, 
    1404115200, 1404118800, 1404122400, 1404126000, 1404129600, 1404133200, 
    1404136800, 1404140400, 1404144000, 1404147600, 1404151200, 1404154800, 
    1404158400, 1404162000, 1404165600, 1404169200, 1404172800, 1404176400, 
    1404180000, 1404183600, 1404187200, 1404190800, 1404194400, 1404198000, 
    1404201600, 1404205200, 1404208800, 1404212400, 1404216000, 1404219600, 
    1404223200, 1404226800, 1404230400, 1404234000, 1404237600, 1404241200, 
    1404244800, 1404248400, 1404252000, 1404255600, 1404259200, 1404262800, 
    1404266400, 1404270000, 1404273600, 1404277200, 1404280800, 1404284400, 
    1404288000, 1404291600, 1404295200, 1404298800, 1404302400, 1404306000, 
    1404309600, 1404313200, 1404316800, 1404320400, 1404324000, 1404327600, 
    1404331200, 1404334800, 1404338400, 1404342000, 1404345600, 1404349200, 
    1404352800, 1404356400, 1404360000, 1404363600, 1404367200, 1404370800, 
    1404374400, 1404378000, 1404381600, 1404385200, 1404388800, 1404392400, 
    1404396000, 1404399600, 1404403200, 1404406800, 1404410400, 1404414000, 
    1404417600, 1404421200, 1404424800, 1404428400, 1404432000, 1404435600, 
    1404439200, 1404442800, 1404446400, 1404450000, 1404453600, 1404457200, 
    1404460800, 1404464400, 1404468000, 1404471600, 1404475200, 1404478800, 
    1404482400, 1404486000, 1404489600, 1404493200, 1404496800, 1404500400, 
    1404504000, 1404507600, 1404511200, 1404514800, 1404518400, 1404522000, 
    1404525600, 1404529200, 1404532800, 1404536400, 1404540000, 1404543600, 
    1404547200, 1404550800, 1404554400, 1404558000, 1404561600, 1404565200, 
    1404568800, 1404572400, 1404576000, 1404579600, 1404583200, 1404586800, 
    1404590400, 1404594000, 1404597600, 1404601200, 1404604800, 1404608400, 
    1404612000, 1404615600, 1404619200, 1404622800, 1404626400, 1404630000, 
    1404633600, 1404637200, 1404640800, 1404644400, 1404648000, 1404651600, 
    1404655200, 1404658800, 1404662400, 1404666000, 1404669600, 1404673200, 
    1404676800, 1404680400, 1404684000, 1404687600, 1404691200, 1404694800, 
    1404698400, 1404702000, 1404705600, 1404709200, 1404712800, 1404716400, 
    1404720000, 1404723600, 1404727200, 1404730800, 1404734400, 1404738000, 
    1404741600, 1404745200, 1404748800, 1404752400, 1404756000, 1404759600, 
    1404763200, 1404766800, 1404770400, 1404774000, 1404777600, 1404781200, 
    1404784800, 1404788400, 1404792000, 1404795600, 1404799200, 1404802800, 
    1404806400, 1404810000, 1404813600, 1404817200, 1404820800, 1404824400, 
    1404828000, 1404831600, 1404835200, 1404838800, 1404842400, 1404846000, 
    1404849600, 1404853200, 1404856800, 1404860400, 1404864000, 1404867600, 
    1404871200, 1404874800, 1404878400, 1404882000, 1404885600, 1404889200, 
    1404892800, 1404896400, 1404900000, 1404903600, 1404907200, 1404910800, 
    1404914400, 1404918000, 1404921600, 1404925200, 1404928800, 1404932400, 
    1404936000, 1404939600, 1404943200, 1404946800, 1404950400, 1404954000, 
    1404957600, 1404961200, 1404964800, 1404968400, 1404972000, 1404975600, 
    1404979200, 1404982800, 1404986400, 1404990000, 1404993600, 1404997200, 
    1405000800, 1405004400, 1405008000, 1405011600, 1405015200, 1405018800, 
    1405022400, 1405026000, 1405029600, 1405033200, 1405036800, 1405040400, 
    1405044000, 1405047600, 1405051200, 1405054800, 1405058400, 1405062000, 
    1405065600, 1405069200, 1405072800, 1405076400, 1405080000, 1405083600, 
    1405087200, 1405090800, 1405094400, 1405098000, 1405101600, 1405105200, 
    1405108800, 1405112400, 1405116000, 1405119600, 1405123200, 1405126800, 
    1405130400, 1405134000, 1405137600, 1405141200, 1405144800, 1405148400, 
    1405152000, 1405155600, 1405159200, 1405162800, 1405166400, 1405170000, 
    1405173600, 1405177200, 1405180800, 1405184400, 1405188000, 1405191600, 
    1405195200, 1405198800, 1405202400, 1405206000, 1405209600, 1405213200, 
    1405216800, 1405220400, 1405224000, 1405227600, 1405231200, 1405234800, 
    1405238400, 1405242000, 1405245600, 1405249200, 1405252800, 1405256400, 
    1405260000, 1405263600, 1405267200, 1405270800, 1405274400, 1405278000, 
    1405281600, 1405285200, 1405288800, 1405292400, 1405296000, 1405299600, 
    1405303200, 1405306800, 1405310400, 1405314000, 1405317600, 1405321200, 
    1405324800, 1405328400, 1405332000, 1405335600, 1405339200, 1405342800, 
    1405346400, 1405350000, 1405353600, 1405357200, 1405360800, 1405364400, 
    1405368000, 1405371600, 1405375200, 1405378800, 1405382400, 1405386000, 
    1405389600, 1405393200, 1405396800, 1405400400, 1405404000, 1405407600, 
    1405411200, 1405414800, 1405418400, 1405422000, 1405425600, 1405429200, 
    1405432800, 1405436400, 1405440000, 1405443600, 1405447200, 1405450800, 
    1405454400, 1405458000, 1405461600, 1405465200, 1405468800, 1405472400, 
    1405476000, 1405479600, 1405483200, 1405486800, 1405490400, 1405494000, 
    1405497600, 1405501200, 1405504800, 1405508400, 1405512000, 1405515600, 
    1405519200, 1405522800, 1405526400, 1405530000, 1405533600, 1405537200, 
    1405540800, 1405544400, 1405548000, 1405551600, 1405555200, 1405558800, 
    1405562400, 1405566000, 1405569600, 1405573200, 1405576800, 1405580400, 
    1405584000, 1405587600, 1405591200, 1405594800, 1405598400, 1405602000, 
    1405605600, 1405609200, 1405612800, 1405616400, 1405620000, 1405623600, 
    1405627200, 1405630800, 1405634400, 1405638000, 1405641600, 1405645200, 
    1405648800, 1405652400, 1405656000, 1405659600, 1405663200, 1405666800, 
    1405670400, 1405674000, 1405677600, 1405681200, 1405684800, 1405688400, 
    1405692000, 1405695600, 1405699200, 1405702800, 1405706400, 1405710000, 
    1405713600, 1405717200, 1405720800, 1405724400, 1405728000, 1405731600, 
    1405735200, 1405738800, 1405742400, 1405746000, 1405749600, 1405753200, 
    1405756800, 1405760400, 1405764000, 1405767600, 1405771200, 1405774800, 
    1405778400, 1405782000, 1405785600, 1405789200, 1405792800, 1405796400, 
    1405800000, 1405803600, 1405807200, 1405810800, 1405814400, 1405818000, 
    1405821600, 1405825200, 1405828800, 1405832400, 1405836000, 1405839600, 
    1405843200, 1405846800, 1405850400, 1405854000, 1405857600, 1405861200, 
    1405864800, 1405868400, 1405872000, 1405875600, 1405879200, 1405882800, 
    1405886400, 1405890000, 1405893600, 1405897200, 1405900800, 1405904400, 
    1405908000, 1405911600, 1405915200, 1405918800, 1405922400, 1405926000, 
    1405929600, 1405933200, 1405936800, 1405940400, 1405944000, 1405947600, 
    1405951200, 1405954800, 1405958400, 1405962000, 1405965600, 1405969200, 
    1405972800, 1405976400, 1405980000, 1405983600, 1405987200, 1405990800, 
    1405994400, 1405998000, 1406001600, 1406005200, 1406008800, 1406012400, 
    1406016000, 1406019600, 1406023200, 1406026800, 1406030400, 1406034000, 
    1406037600, 1406041200, 1406044800, 1406048400, 1406052000, 1406055600, 
    1406059200, 1406062800, 1406066400, 1406070000, 1406073600, 1406077200, 
    1406080800, 1406084400, 1406088000, 1406091600, 1406095200, 1406098800, 
    1406102400, 1406106000, 1406109600, 1406113200, 1406116800, 1406120400, 
    1406124000, 1406127600, 1406131200, 1406134800, 1406138400, 1406142000, 
    1406145600, 1406149200, 1406152800, 1406156400, 1406160000, 1406163600, 
    1406167200, 1406170800, 1406174400, 1406178000, 1406181600, 1406185200, 
    1406188800, 1406192400, 1406196000, 1406199600, 1406203200, 1406206800, 
    1406210400, 1406214000, 1406217600, 1406221200, 1406224800, 1406228400, 
    1406232000, 1406235600, 1406239200, 1406242800, 1406246400, 1406250000, 
    1406253600, 1406257200, 1406260800, 1406264400, 1406268000, 1406271600, 
    1406275200, 1406278800, 1406282400, 1406286000, 1406289600, 1406293200, 
    1406296800, 1406300400, 1406304000, 1406307600, 1406311200, 1406314800, 
    1406318400, 1406322000, 1406325600, 1406329200, 1406332800, 1406336400, 
    1406340000, 1406343600, 1406347200, 1406350800, 1406354400, 1406358000, 
    1406361600, 1406365200, 1406368800, 1406372400, 1406376000, 1406379600, 
    1406383200, 1406386800, 1406390400, 1406394000, 1406397600, 1406401200, 
    1406404800, 1406408400, 1406412000, 1406415600, 1406419200, 1406422800, 
    1406426400, 1406430000, 1406433600, 1406437200, 1406440800, 1406444400, 
    1406448000, 1406451600, 1406455200, 1406458800, 1406462400, 1406466000, 
    1406469600, 1406473200, 1406476800, 1406480400, 1406484000, 1406487600, 
    1406491200, 1406494800, 1406498400, 1406502000, 1406505600, 1406509200, 
    1406512800, 1406516400, 1406520000, 1406523600, 1406527200, 1406530800, 
    1406534400, 1406538000, 1406541600, 1406545200, 1406548800, 1406552400, 
    1406556000, 1406559600, 1406563200, 1406566800, 1406570400, 1406574000, 
    1406577600, 1406581200, 1406584800, 1406588400, 1406592000, 1406595600, 
    1406599200, 1406602800, 1406606400, 1406610000, 1406613600, 1406617200, 
    1406620800, 1406624400, 1406628000, 1406631600, 1406635200, 1406638800, 
    1406642400, 1406646000, 1406649600, 1406653200, 1406656800, 1406660400, 
    1406664000, 1406667600, 1406671200, 1406674800, 1406678400, 1406682000, 
    1406685600, 1406689200, 1406692800, 1406696400, 1406700000, 1406703600, 
    1406707200, 1406710800, 1406714400, 1406718000, 1406721600, 1406725200, 
    1406728800, 1406732400, 1406736000, 1406739600, 1406743200, 1406746800, 
    1406750400, 1406754000, 1406757600, 1406761200, 1406764800, 1406768400, 
    1406772000, 1406775600, 1406779200, 1406782800, 1406786400, 1406790000, 
    1406793600, 1406797200, 1406800800, 1406804400, 1406808000, 1406811600, 
    1406815200, 1406818800, 1406822400, 1406826000, 1406829600, 1406833200, 
    1406836800, 1406840400, 1406844000, 1406847600, 1406851200, 1406854800, 
    1406858400, 1406862000, 1406865600, 1406869200, 1406872800, 1406876400, 
    1406880000, 1406883600, 1406887200, 1406890800, 1406894400, 1406898000, 
    1406901600, 1406905200, 1406908800, 1406912400, 1406916000, 1406919600, 
    1406923200, 1406926800, 1406930400, 1406934000, 1406937600, 1406941200, 
    1406944800, 1406948400, 1406952000, 1406955600, 1406959200, 1406962800, 
    1406966400, 1406970000, 1406973600, 1406977200, 1406980800, 1406984400, 
    1406988000, 1406991600, 1406995200, 1406998800, 1407002400, 1407006000, 
    1407009600, 1407013200, 1407016800, 1407020400, 1407024000, 1407027600, 
    1407031200, 1407034800, 1407038400, 1407042000, 1407045600, 1407049200, 
    1407052800, 1407056400, 1407060000, 1407063600, 1407067200, 1407070800, 
    1407074400, 1407078000, 1407081600, 1407085200, 1407088800, 1407092400, 
    1407096000, 1407099600, 1407103200, 1407106800, 1407110400, 1407114000, 
    1407117600, 1407121200, 1407124800, 1407128400, 1407132000, 1407135600, 
    1407139200, 1407142800, 1407146400, 1407150000, 1407153600, 1407157200, 
    1407160800, 1407164400, 1407168000, 1407171600, 1407175200, 1407178800, 
    1407182400, 1407186000, 1407189600, 1407193200, 1407196800, 1407200400, 
    1407204000, 1407207600, 1407211200, 1407214800, 1407218400, 1407222000, 
    1407225600, 1407229200, 1407232800, 1407236400, 1407240000, 1407243600, 
    1407247200, 1407250800, 1407254400, 1407258000, 1407261600, 1407265200, 
    1407268800, 1407272400, 1407276000, 1407279600, 1407283200, 1407286800, 
    1407290400, 1407294000, 1407297600, 1407301200, 1407304800, 1407308400, 
    1407312000, 1407315600, 1407319200, 1407322800, 1407326400, 1407330000, 
    1407333600, 1407337200, 1407340800, 1407344400, 1407348000, 1407351600, 
    1407355200, 1407358800, 1407362400, 1407366000, 1407369600, 1407373200, 
    1407376800, 1407380400, 1407384000, 1407387600, 1407391200, 1407394800, 
    1407398400, 1407402000, 1407405600, 1407409200, 1407412800, 1407416400, 
    1407420000, 1407423600, 1407427200, 1407430800, 1407434400, 1407438000, 
    1407441600, 1407445200, 1407448800, 1407452400, 1407456000, 1407459600, 
    1407463200, 1407466800, 1407470400, 1407474000, 1407477600, 1407481200, 
    1407484800, 1407488400, 1407492000, 1407495600, 1407499200, 1407502800, 
    1407506400, 1407510000, 1407513600, 1407517200, 1407520800, 1407524400, 
    1407528000, 1407531600, 1407535200, 1407538800, 1407542400, 1407546000, 
    1407549600, 1407553200, 1407556800, 1407560400, 1407564000, 1407567600, 
    1407571200, 1407574800, 1407578400, 1407582000, 1407585600, 1407589200, 
    1407592800, 1407596400, 1407600000, 1407603600, 1407607200, 1407610800, 
    1407614400, 1407618000, 1407621600, 1407625200, 1407628800, 1407632400, 
    1407636000, 1407639600, 1407643200, 1407646800, 1407650400, 1407654000, 
    1407657600, 1407661200, 1407664800, 1407668400, 1407672000, 1407675600, 
    1407679200, 1407682800, 1407686400, 1407690000, 1407693600, 1407697200, 
    1407700800, 1407704400, 1407708000, 1407711600, 1407715200, 1407718800, 
    1407722400, 1407726000, 1407729600, 1407733200, 1407736800, 1407740400, 
    1407744000, 1407747600, 1407751200, 1407754800, 1407758400, 1407762000, 
    1407765600, 1407769200, 1407772800, 1407776400, 1407780000, 1407783600, 
    1407787200, 1407790800, 1407794400, 1407798000, 1407801600, 1407805200, 
    1407808800, 1407812400, 1407816000, 1407819600, 1407823200, 1407826800, 
    1407830400, 1407834000, 1407837600, 1407841200, 1407844800, 1407848400, 
    1407852000, 1407855600, 1407859200, 1407862800, 1407866400, 1407870000, 
    1407873600, 1407877200, 1407880800, 1407884400, 1407888000, 1407891600, 
    1407895200, 1407898800, 1407902400, 1407906000, 1407909600, 1407913200, 
    1407916800, 1407920400, 1407924000, 1407927600, 1407931200, 1407934800, 
    1407938400, 1407942000, 1407945600, 1407949200, 1407952800, 1407956400, 
    1407960000, 1407963600, 1407967200, 1407970800, 1407974400, 1407978000, 
    1407981600, 1407985200, 1407988800, 1407992400, 1407996000, 1407999600, 
    1408003200, 1408006800, 1408010400, 1408014000, 1408017600, 1408021200, 
    1408024800, 1408028400, 1408032000, 1408035600, 1408039200, 1408042800, 
    1408046400, 1408050000, 1408053600, 1408057200, 1408060800, 1408064400, 
    1408068000, 1408071600, 1408075200, 1408078800, 1408082400, 1408086000, 
    1408089600, 1408093200, 1408096800, 1408100400, 1408104000, 1408107600, 
    1408111200, 1408114800, 1408118400, 1408122000, 1408125600, 1408129200, 
    1408132800, 1408136400, 1408140000, 1408143600, 1408147200, 1408150800, 
    1408154400, 1408158000, 1408161600, 1408165200, 1408168800, 1408172400, 
    1408176000, 1408179600, 1408183200, 1408186800, 1408190400, 1408194000, 
    1408197600, 1408201200, 1408204800, 1408208400, 1408212000, 1408215600, 
    1408219200, 1408222800, 1408226400, 1408230000, 1408233600, 1408237200, 
    1408240800, 1408244400, 1408248000, 1408251600, 1408255200, 1408258800, 
    1408262400, 1408266000, 1408269600, 1408273200, 1408276800, 1408280400, 
    1408284000, 1408287600, 1408291200, 1408294800, 1408298400, 1408302000, 
    1408305600, 1408309200, 1408312800, 1408316400, 1408320000, 1408323600, 
    1408327200, 1408330800, 1408334400, 1408338000, 1408341600, 1408345200, 
    1408348800, 1408352400, 1408356000, 1408359600, 1408363200, 1408366800, 
    1408370400, 1408374000, 1408377600, 1408381200, 1408384800, 1408388400, 
    1408392000, 1408395600, 1408399200, 1408402800, 1408406400, 1408410000, 
    1408413600, 1408417200, 1408420800, 1408424400, 1408428000, 1408431600, 
    1408435200, 1408438800, 1408442400, 1408446000, 1408449600, 1408453200, 
    1408456800, 1408460400, 1408464000, 1408467600, 1408471200, 1408474800, 
    1408478400, 1408482000, 1408485600, 1408489200, 1408492800, 1408496400, 
    1408500000, 1408503600, 1408507200, 1408510800, 1408514400, 1408518000, 
    1408521600, 1408525200, 1408528800, 1408532400, 1408536000, 1408539600, 
    1408543200, 1408546800, 1408550400, 1408554000, 1408557600, 1408561200, 
    1408564800, 1408568400, 1408572000, 1408575600, 1408579200, 1408582800, 
    1408586400, 1408590000, 1408593600, 1408597200, 1408600800, 1408604400, 
    1408608000, 1408611600, 1408615200, 1408618800, 1408622400, 1408626000, 
    1408629600, 1408633200, 1408636800, 1408640400, 1408644000, 1408647600, 
    1408651200, 1408654800, 1408658400, 1408662000, 1408665600, 1408669200, 
    1408672800, 1408676400, 1408680000, 1408683600, 1408687200, 1408690800, 
    1408694400, 1408698000, 1408701600, 1408705200, 1408708800, 1408712400, 
    1408716000, 1408719600, 1408723200, 1408726800, 1408730400, 1408734000, 
    1408737600, 1408741200, 1408744800, 1408748400, 1408752000, 1408755600, 
    1408759200, 1408762800, 1408766400, 1408770000, 1408773600, 1408777200, 
    1408780800, 1408784400, 1408788000, 1408791600, 1408795200, 1408798800, 
    1408802400, 1408806000, 1408809600, 1408813200, 1408816800, 1408820400, 
    1408824000, 1408827600, 1408831200, 1408834800, 1408838400, 1408842000, 
    1408845600, 1408849200, 1408852800, 1408856400, 1408860000, 1408863600, 
    1408867200, 1408870800, 1408874400, 1408878000, 1408881600, 1408885200, 
    1408888800, 1408892400, 1408896000, 1408899600, 1408903200, 1408906800, 
    1408910400, 1408914000, 1408917600, 1408921200, 1408924800, 1408928400, 
    1408932000, 1408935600, 1408939200, 1408942800, 1408946400, 1408950000, 
    1408953600, 1408957200, 1408960800, 1408964400, 1408968000, 1408971600, 
    1408975200, 1408978800, 1408982400, 1408986000, 1408989600, 1408993200, 
    1408996800, 1409000400, 1409004000, 1409007600, 1409011200, 1409014800, 
    1409018400, 1409022000, 1409025600, 1409029200, 1409032800, 1409036400, 
    1409040000, 1409043600, 1409047200, 1409050800, 1409054400, 1409058000, 
    1409061600, 1409065200, 1409068800, 1409072400, 1409076000, 1409079600, 
    1409083200, 1409086800, 1409090400, 1409094000, 1409097600, 1409101200, 
    1409104800, 1409108400, 1409112000, 1409115600, 1409119200, 1409122800, 
    1409126400, 1409130000, 1409133600, 1409137200, 1409140800, 1409144400, 
    1409148000, 1409151600, 1409155200, 1409158800, 1409162400, 1409166000, 
    1409169600, 1409173200, 1409176800, 1409180400, 1409184000, 1409187600, 
    1409191200, 1409194800, 1409198400, 1409202000, 1409205600, 1409209200, 
    1409212800, 1409216400, 1409220000, 1409223600, 1409227200, 1409230800, 
    1409234400, 1409238000, 1409241600, 1409245200, 1409248800, 1409252400, 
    1409256000, 1409259600, 1409263200, 1409266800, 1409270400, 1409274000, 
    1409277600, 1409281200, 1409284800, 1409288400, 1409292000, 1409295600, 
    1409299200, 1409302800, 1409306400, 1409310000, 1409313600, 1409317200, 
    1409320800, 1409324400, 1409328000, 1409331600, 1409335200, 1409338800, 
    1409342400, 1409346000, 1409349600, 1409353200, 1409356800, 1409360400, 
    1409364000, 1409367600, 1409371200, 1409374800, 1409378400, 1409382000, 
    1409385600, 1409389200, 1409392800, 1409396400, 1409400000, 1409403600, 
    1409407200, 1409410800, 1409414400, 1409418000, 1409421600, 1409425200, 
    1409428800, 1409432400, 1409436000, 1409439600, 1409443200, 1409446800, 
    1409450400, 1409454000, 1409457600, 1409461200, 1409464800, 1409468400, 
    1409472000, 1409475600, 1409479200, 1409482800, 1409486400, 1409490000, 
    1409493600, 1409497200, 1409500800, 1409504400, 1409508000, 1409511600, 
    1409515200, 1409518800, 1409522400, 1409526000, 1409529600, 1409533200, 
    1409536800, 1409540400, 1409544000, 1409547600, 1409551200, 1409554800, 
    1409558400, 1409562000, 1409565600, 1409569200, 1409572800, 1409576400, 
    1409580000, 1409583600, 1409587200, 1409590800, 1409594400, 1409598000, 
    1409601600, 1409605200, 1409608800, 1409612400, 1409616000, 1409619600, 
    1409623200, 1409626800, 1409630400, 1409634000, 1409637600, 1409641200, 
    1409644800, 1409648400, 1409652000, 1409655600, 1409659200, 1409662800, 
    1409666400, 1409670000, 1409673600, 1409677200, 1409680800, 1409684400, 
    1409688000, 1409691600, 1409695200, 1409698800, 1409702400, 1409706000, 
    1409709600, 1409713200, 1409716800, 1409720400, 1409724000, 1409727600, 
    1409731200, 1409734800, 1409738400, 1409742000, 1409745600, 1409749200, 
    1409752800, 1409756400, 1409760000, 1409763600, 1409767200, 1409770800, 
    1409774400, 1409778000, 1409781600, 1409785200, 1409788800, 1409792400, 
    1409796000, 1409799600, 1409803200, 1409806800, 1409810400, 1409814000, 
    1409817600, 1409821200, 1409824800, 1409828400, 1409832000, 1409835600, 
    1409839200, 1409842800, 1409846400, 1409850000, 1409853600, 1409857200, 
    1409860800, 1409864400, 1409868000, 1409871600, 1409875200, 1409878800, 
    1409882400, 1409886000, 1409889600, 1409893200, 1409896800, 1409900400, 
    1409904000, 1409907600, 1409911200, 1409914800, 1409918400, 1409922000, 
    1409925600, 1409929200, 1409932800, 1409936400, 1409940000, 1409943600, 
    1409947200, 1409950800, 1409954400, 1409958000, 1409961600, 1409965200, 
    1409968800, 1409972400, 1409976000, 1409979600, 1409983200, 1409986800, 
    1409990400, 1409994000, 1409997600, 1410001200, 1410004800, 1410008400, 
    1410012000, 1410015600, 1410019200, 1410022800, 1410026400, 1410030000, 
    1410033600, 1410037200, 1410040800, 1410044400, 1410048000, 1410051600, 
    1410055200, 1410058800, 1410062400, 1410066000, 1410069600, 1410073200, 
    1410076800, 1410080400, 1410084000, 1410087600, 1410091200, 1410094800, 
    1410098400, 1410102000, 1410105600, 1410109200, 1410112800, 1410116400, 
    1410120000, 1410123600, 1410127200, 1410130800, 1410134400, 1410138000, 
    1410141600, 1410145200, 1410148800, 1410152400, 1410156000, 1410159600, 
    1410163200, 1410166800, 1410170400, 1410174000, 1410177600, 1410181200, 
    1410184800, 1410188400, 1410192000, 1410195600, 1410199200, 1410202800, 
    1410206400, 1410210000, 1410213600, 1410217200, 1410220800, 1410224400, 
    1410228000, 1410231600, 1410235200, 1410238800, 1410242400, 1410246000, 
    1410249600, 1410253200, 1410256800, 1410260400, 1410264000, 1410267600, 
    1410271200, 1410274800, 1410278400, 1410282000, 1410285600, 1410289200, 
    1410292800, 1410296400, 1410300000, 1410303600, 1410307200, 1410310800, 
    1410314400, 1410318000, 1410321600, 1410325200, 1410328800, 1410332400, 
    1410336000, 1410339600, 1410343200, 1410346800, 1410350400, 1410354000, 
    1410357600, 1410361200, 1410364800, 1410368400, 1410372000, 1410375600, 
    1410379200, 1410382800, 1410386400, 1410390000, 1410393600, 1410397200, 
    1410400800, 1410404400, 1410408000, 1410411600, 1410415200, 1410418800, 
    1410422400, 1410426000, 1410429600, 1410433200, 1410436800, 1410440400, 
    1410444000, 1410447600, 1410451200, 1410454800, 1410458400, 1410462000, 
    1410465600, 1410469200, 1410472800, 1410476400, 1410480000, 1410483600, 
    1410487200, 1410490800, 1410494400, 1410498000, 1410501600, 1410505200, 
    1410508800, 1410512400, 1410516000, 1410519600, 1410523200, 1410526800, 
    1410530400, 1410534000, 1410537600, 1410541200, 1410544800, 1410548400, 
    1410552000, 1410555600, 1410559200, 1410562800, 1410566400, 1410570000, 
    1410573600, 1410577200, 1410580800, 1410584400, 1410588000, 1410591600, 
    1410595200, 1410598800, 1410602400, 1410606000, 1410609600, 1410613200, 
    1410616800, 1410620400, 1410624000, 1410627600, 1410631200, 1410634800, 
    1410638400, 1410642000, 1410645600, 1410649200, 1410652800, 1410656400, 
    1410660000, 1410663600, 1410667200, 1410670800, 1410674400, 1410678000, 
    1410681600, 1410685200, 1410688800, 1410692400, 1410696000, 1410699600, 
    1410703200, 1410706800, 1410710400, 1410714000, 1410717600, 1410721200, 
    1410724800, 1410728400, 1410732000, 1410735600, 1410739200, 1410742800, 
    1410746400, 1410750000, 1410753600, 1410757200, 1410760800, 1410764400, 
    1410768000, 1410771600, 1410775200, 1410778800, 1410782400, 1410786000, 
    1410789600, 1410793200, 1410796800, 1410800400, 1410804000, 1410807600, 
    1410811200, 1410814800, 1410818400, 1410822000, 1410825600, 1410829200, 
    1410832800, 1410836400, 1410840000, 1410843600, 1410847200, 1410850800, 
    1410854400, 1410858000, 1410861600, 1410865200, 1410868800, 1410872400, 
    1410876000, 1410879600, 1410883200, 1410886800, 1410890400, 1410894000, 
    1410897600, 1410901200, 1410904800, 1410908400, 1410912000, 1410915600, 
    1410919200, 1410922800, 1410926400, 1410930000, 1410933600, 1410937200, 
    1410940800, 1410944400, 1410948000, 1410951600, 1410955200, 1410958800, 
    1410962400, 1410966000, 1410969600, 1410973200, 1410976800, 1410980400, 
    1410984000, 1410987600, 1410991200, 1410994800, 1410998400, 1411002000, 
    1411005600, 1411009200, 1411012800, 1411016400, 1411020000, 1411023600, 
    1411027200, 1411030800, 1411034400, 1411038000, 1411041600, 1411045200, 
    1411048800, 1411052400, 1411056000, 1411059600, 1411063200, 1411066800, 
    1411070400, 1411074000, 1411077600, 1411081200, 1411084800, 1411088400, 
    1411092000, 1411095600, 1411099200, 1411102800, 1411106400, 1411110000, 
    1411113600, 1411117200, 1411120800, 1411124400, 1411128000, 1411131600, 
    1411135200, 1411138800, 1411142400, 1411146000, 1411149600, 1411153200, 
    1411156800, 1411160400, 1411164000, 1411167600, 1411171200, 1411174800, 
    1411178400, 1411182000, 1411185600, 1411189200, 1411192800, 1411196400, 
    1411200000, 1411203600, 1411207200, 1411210800, 1411214400, 1411218000, 
    1411221600, 1411225200, 1411228800, 1411232400, 1411236000, 1411239600, 
    1411243200, 1411246800, 1411250400, 1411254000, 1411257600, 1411261200, 
    1411264800, 1411268400, 1411272000, 1411275600, 1411279200, 1411282800, 
    1411286400, 1411290000, 1411293600, 1411297200, 1411300800, 1411304400, 
    1411308000, 1411311600, 1411315200, 1411318800, 1411322400, 1411326000, 
    1411329600, 1411333200, 1411336800, 1411340400, 1411344000, 1411347600, 
    1411351200, 1411354800, 1411358400, 1411362000, 1411365600, 1411369200, 
    1411372800, 1411376400, 1411380000, 1411383600, 1411387200, 1411390800, 
    1411394400, 1411398000, 1411401600, 1411405200, 1411408800, 1411412400, 
    1411416000, 1411419600, 1411423200, 1411426800, 1411430400, 1411434000, 
    1411437600, 1411441200, 1411444800, 1411448400, 1411452000, 1411455600, 
    1411459200, 1411462800, 1411466400, 1411470000, 1411473600, 1411477200, 
    1411480800, 1411484400, 1411488000, 1411491600, 1411495200, 1411498800, 
    1411502400, 1411506000, 1411509600, 1411513200, 1411516800, 1411520400, 
    1411524000, 1411527600, 1411531200, 1411534800, 1411538400, 1411542000, 
    1411545600, 1411549200, 1411552800, 1411556400, 1411560000, 1411563600, 
    1411567200, 1411570800, 1411574400, 1411578000, 1411581600, 1411585200, 
    1411588800, 1411592400, 1411596000, 1411599600, 1411603200, 1411606800, 
    1411610400, 1411614000, 1411617600, 1411621200, 1411624800, 1411628400, 
    1411632000, 1411635600, 1411639200, 1411642800, 1411646400, 1411650000, 
    1411653600, 1411657200, 1411660800, 1411664400, 1411668000, 1411671600, 
    1411675200, 1411678800, 1411682400, 1411686000, 1411689600, 1411693200, 
    1411696800, 1411700400, 1411704000, 1411707600, 1411711200, 1411714800, 
    1411718400, 1411722000, 1411725600, 1411729200, 1411732800, 1411736400, 
    1411740000, 1411743600, 1411747200, 1411750800, 1411754400, 1411758000, 
    1411761600, 1411765200, 1411768800, 1411772400, 1411776000, 1411779600, 
    1411783200, 1411786800, 1411790400, 1411794000, 1411797600, 1411801200, 
    1411804800, 1411808400, 1411812000, 1411815600, 1411819200, 1411822800, 
    1411826400, 1411830000, 1411833600, 1411837200, 1411840800, 1411844400, 
    1411848000, 1411851600, 1411855200, 1411858800, 1411862400, 1411866000, 
    1411869600, 1411873200, 1411876800, 1411880400, 1411884000, 1411887600, 
    1411891200, 1411894800, 1411898400, 1411902000, 1411905600, 1411909200, 
    1411912800, 1411916400, 1411920000, 1411923600, 1411927200, 1411930800, 
    1411934400, 1411938000, 1411941600, 1411945200, 1411948800, 1411952400, 
    1411956000, 1411959600, 1411963200, 1411966800, 1411970400, 1411974000, 
    1411977600, 1411981200, 1411984800, 1411988400, 1411992000, 1411995600, 
    1411999200, 1412002800, 1412006400, 1412010000, 1412013600, 1412017200, 
    1412020800, 1412024400, 1412028000, 1412031600, 1412035200, 1412038800, 
    1412042400, 1412046000, 1412049600, 1412053200, 1412056800, 1412060400, 
    1412064000, 1412067600, 1412071200, 1412074800, 1412078400, 1412082000, 
    1412085600, 1412089200, 1412092800, 1412096400, 1412100000, 1412103600, 
    1412107200, 1412110800, 1412114400, 1412118000, 1412121600, 1412125200, 
    1412128800, 1412132400, 1412136000, 1412139600, 1412143200, 1412146800, 
    1412150400, 1412154000, 1412157600, 1412161200, 1412164800, 1412168400, 
    1412172000, 1412175600, 1412179200, 1412182800, 1412186400, 1412190000, 
    1412193600, 1412197200, 1412200800, 1412204400, 1412208000, 1412211600, 
    1412215200, 1412218800, 1412222400, 1412226000, 1412229600, 1412233200, 
    1412236800, 1412240400, 1412244000, 1412247600, 1412251200, 1412254800, 
    1412258400, 1412262000, 1412265600, 1412269200, 1412272800, 1412276400, 
    1412280000, 1412283600, 1412287200, 1412290800, 1412294400, 1412298000, 
    1412301600, 1412305200, 1412308800, 1412312400, 1412316000, 1412319600, 
    1412323200, 1412326800, 1412330400, 1412334000, 1412337600, 1412341200, 
    1412344800, 1412348400, 1412352000, 1412355600, 1412359200, 1412362800, 
    1412366400, 1412370000, 1412373600, 1412377200, 1412380800, 1412384400, 
    1412388000, 1412391600, 1412395200, 1412398800, 1412402400, 1412406000, 
    1412409600, 1412413200, 1412416800, 1412420400, 1412424000, 1412427600, 
    1412431200, 1412434800, 1412438400, 1412442000, 1412445600, 1412449200, 
    1412452800, 1412456400, 1412460000, 1412463600, 1412467200, 1412470800, 
    1412474400, 1412478000, 1412481600, 1412485200, 1412488800, 1412492400, 
    1412496000, 1412499600, 1412503200, 1412506800, 1412510400, 1412514000, 
    1412517600, 1412521200, 1412524800, 1412528400, 1412532000, 1412535600, 
    1412539200, 1412542800, 1412546400, 1412550000, 1412553600, 1412557200, 
    1412560800, 1412564400, 1412568000, 1412571600, 1412575200, 1412578800, 
    1412582400, 1412586000, 1412589600, 1412593200, 1412596800, 1412600400, 
    1412604000, 1412607600, 1412611200, 1412614800, 1412618400, 1412622000, 
    1412625600, 1412629200, 1412632800, 1412636400, 1412640000, 1412643600, 
    1412647200, 1412650800, 1412654400, 1412658000, 1412661600, 1412665200, 
    1412668800, 1412672400, 1412676000, 1412679600, 1412683200, 1412686800, 
    1412690400, 1412694000, 1412697600, 1412701200, 1412704800, 1412708400, 
    1412712000, 1412715600, 1412719200, 1412722800, 1412726400, 1412730000, 
    1412733600, 1412737200, 1412740800, 1412744400, 1412748000, 1412751600, 
    1412755200, 1412758800, 1412762400, 1412766000, 1412769600, 1412773200, 
    1412776800, 1412780400, 1412784000, 1412787600, 1412791200, 1412794800, 
    1412798400, 1412802000, 1412805600, 1412809200, 1412812800, 1412816400, 
    1412820000, 1412823600, 1412827200, 1412830800, 1412834400, 1412838000, 
    1412841600, 1412845200, 1412848800, 1412852400, 1412856000, 1412859600, 
    1412863200, 1412866800, 1412870400, 1412874000, 1412877600, 1412881200, 
    1412884800, 1412888400, 1412892000, 1412895600, 1412899200, 1412902800, 
    1412906400, 1412910000, 1412913600, 1412917200, 1412920800, 1412924400, 
    1412928000, 1412931600, 1412935200, 1412938800, 1412942400, 1412946000, 
    1412949600, 1412953200, 1412956800, 1412960400, 1412964000, 1412967600, 
    1412971200, 1412974800, 1412978400, 1412982000, 1412985600, 1412989200, 
    1412992800, 1412996400, 1413000000, 1413003600, 1413007200, 1413010800, 
    1413014400, 1413018000, 1413021600, 1413025200, 1413028800, 1413032400, 
    1413036000, 1413039600, 1413043200, 1413046800, 1413050400, 1413054000, 
    1413057600, 1413061200, 1413064800, 1413068400, 1413072000, 1413075600, 
    1413079200, 1413082800, 1413086400, 1413090000, 1413093600, 1413097200, 
    1413100800, 1413104400, 1413108000, 1413111600, 1413115200, 1413118800, 
    1413122400, 1413126000, 1413129600, 1413133200, 1413136800, 1413140400, 
    1413144000, 1413147600, 1413151200, 1413154800, 1413158400, 1413162000, 
    1413165600, 1413169200, 1413172800, 1413176400, 1413180000, 1413183600, 
    1413187200, 1413190800, 1413194400, 1413198000, 1413201600, 1413205200, 
    1413208800, 1413212400, 1413216000, 1413219600, 1413223200, 1413226800, 
    1413230400, 1413234000, 1413237600, 1413241200, 1413244800, 1413248400, 
    1413252000, 1413255600, 1413259200, 1413262800, 1413266400, 1413270000, 
    1413273600, 1413277200, 1413280800, 1413284400, 1413288000, 1413291600, 
    1413295200, 1413298800, 1413302400, 1413306000, 1413309600, 1413313200, 
    1413316800, 1413320400, 1413324000, 1413327600, 1413331200, 1413334800, 
    1413338400, 1413342000, 1413345600, 1413349200, 1413352800, 1413356400, 
    1413360000, 1413363600, 1413367200, 1413370800, 1413374400, 1413378000, 
    1413381600, 1413385200, 1413388800, 1413392400, 1413396000, 1413399600, 
    1413403200, 1413406800, 1413410400, 1413414000, 1413417600, 1413421200, 
    1413424800, 1413428400, 1413432000, 1413435600, 1413439200, 1413442800, 
    1413446400, 1413450000, 1413453600, 1413457200, 1413460800, 1413464400, 
    1413468000, 1413471600, 1413475200, 1413478800, 1413482400, 1413486000, 
    1413489600, 1413493200, 1413496800, 1413500400, 1413504000, 1413507600, 
    1413511200, 1413514800, 1413518400, 1413522000, 1413525600, 1413529200, 
    1413532800, 1413536400, 1413540000, 1413543600, 1413547200, 1413550800, 
    1413554400, 1413558000, 1413561600, 1413565200, 1413568800, 1413572400, 
    1413576000, 1413579600, 1413583200, 1413586800, 1413590400, 1413594000, 
    1413597600, 1413601200, 1413604800, 1413608400, 1413612000, 1413615600, 
    1413619200, 1413622800, 1413626400, 1413630000, 1413633600, 1413637200, 
    1413640800, 1413644400, 1413648000, 1413651600, 1413655200, 1413658800, 
    1413662400, 1413666000, 1413669600, 1413673200, 1413676800, 1413680400, 
    1413684000, 1413687600, 1413691200, 1413694800, 1413698400, 1413702000, 
    1413705600, 1413709200, 1413712800, 1413716400, 1413720000, 1413723600, 
    1413727200, 1413730800, 1413734400, 1413738000, 1413741600, 1413745200, 
    1413748800, 1413752400, 1413756000, 1413759600, 1413763200, 1413766800, 
    1413770400, 1413774000, 1413777600, 1413781200, 1413784800, 1413788400, 
    1413792000, 1413795600, 1413799200, 1413802800, 1413806400, 1413810000, 
    1413813600, 1413817200, 1413820800, 1413824400, 1413828000, 1413831600, 
    1413835200, 1413838800, 1413842400, 1413846000, 1413849600, 1413853200, 
    1413856800, 1413860400, 1413864000, 1413867600, 1413871200, 1413874800, 
    1413878400, 1413882000, 1413885600, 1413889200, 1413892800, 1413896400, 
    1413900000, 1413903600, 1413907200, 1413910800, 1413914400, 1413918000, 
    1413921600, 1413925200, 1413928800, 1413932400, 1413936000, 1413939600, 
    1413943200, 1413946800, 1413950400, 1413954000, 1413957600, 1413961200, 
    1413964800, 1413968400, 1413972000, 1413975600, 1413979200, 1413982800, 
    1413986400, 1413990000, 1413993600, 1413997200, 1414000800, 1414004400, 
    1414008000, 1414011600, 1414015200, 1414018800, 1414022400, 1414026000, 
    1414029600, 1414033200, 1414036800, 1414040400, 1414044000, 1414047600, 
    1414051200, 1414054800, 1414058400, 1414062000, 1414065600, 1414069200, 
    1414072800, 1414076400, 1414080000, 1414083600, 1414087200, 1414090800, 
    1414094400, 1414098000, 1414101600, 1414105200, 1414108800, 1414112400, 
    1414116000, 1414119600, 1414123200, 1414126800, 1414130400, 1414134000, 
    1414137600, 1414141200, 1414144800, 1414148400, 1414152000, 1414155600, 
    1414159200, 1414162800, 1414166400, 1414170000, 1414173600, 1414177200, 
    1414180800, 1414184400, 1414188000, 1414191600, 1414195200, 1414198800, 
    1414202400, 1414206000, 1414209600, 1414213200, 1414216800, 1414220400, 
    1414224000, 1414227600, 1414231200, 1414234800, 1414238400, 1414242000, 
    1414245600, 1414249200, 1414252800, 1414256400, 1414260000, 1414263600, 
    1414267200, 1414270800, 1414274400, 1414278000, 1414281600, 1414285200, 
    1414288800, 1414292400, 1414296000, 1414299600, 1414303200, 1414306800, 
    1414310400, 1414314000, 1414317600, 1414321200, 1414324800, 1414328400, 
    1414332000, 1414335600, 1414339200, 1414342800, 1414346400, 1414350000, 
    1414353600, 1414357200, 1414360800, 1414364400, 1414368000, 1414371600, 
    1414375200, 1414378800, 1414382400, 1414386000, 1414389600, 1414393200, 
    1414396800, 1414400400, 1414404000, 1414407600, 1414411200, 1414414800, 
    1414418400, 1414422000, 1414425600, 1414429200, 1414432800, 1414436400, 
    1414440000, 1414443600, 1414447200, 1414450800, 1414454400, 1414458000, 
    1414461600, 1414465200, 1414468800, 1414472400, 1414476000, 1414479600, 
    1414483200, 1414486800, 1414490400, 1414494000, 1414497600, 1414501200, 
    1414504800, 1414508400, 1414512000, 1414515600, 1414519200, 1414522800, 
    1414526400, 1414530000, 1414533600, 1414537200, 1414540800, 1414544400, 
    1414548000, 1414551600, 1414555200, 1414558800, 1414562400, 1414566000, 
    1414569600, 1414573200, 1414576800, 1414580400, 1414584000, 1414587600, 
    1414591200, 1414594800, 1414598400, 1414602000, 1414605600, 1414609200, 
    1414612800, 1414616400, 1414620000, 1414623600, 1414627200, 1414630800, 
    1414634400, 1414638000, 1414641600, 1414645200, 1414648800, 1414652400, 
    1414656000, 1414659600, 1414663200, 1414666800, 1414670400, 1414674000, 
    1414677600, 1414681200, 1414684800, 1414688400, 1414692000, 1414695600, 
    1414699200, 1414702800, 1414706400, 1414710000, 1414713600, 1414717200, 
    1414720800, 1414724400, 1414728000, 1414731600, 1414735200, 1414738800, 
    1414742400, 1414746000, 1414749600, 1414753200, 1414756800, 1414760400, 
    1414764000, 1414767600, 1414771200, 1414774800, 1414778400, 1414782000, 
    1414785600, 1414789200, 1414792800, 1414796400, 1414800000, 1414803600, 
    1414807200, 1414810800, 1414814400, 1414818000, 1414821600, 1414825200, 
    1414828800, 1414832400, 1414836000, 1414839600, 1414843200, 1414846800, 
    1414850400, 1414854000, 1414857600, 1414861200, 1414864800, 1414868400, 
    1414872000, 1414875600, 1414879200, 1414882800, 1414886400, 1414890000, 
    1414893600, 1414897200, 1414900800, 1414904400, 1414908000, 1414911600, 
    1414915200, 1414918800, 1414922400, 1414926000, 1414929600, 1414933200, 
    1414936800, 1414940400, 1414944000, 1414947600, 1414951200, 1414954800, 
    1414958400, 1414962000, 1414965600, 1414969200, 1414972800, 1414976400, 
    1414980000, 1414983600, 1414987200, 1414990800, 1414994400, 1414998000, 
    1415001600, 1415005200, 1415008800, 1415012400, 1415016000, 1415019600, 
    1415023200, 1415026800, 1415030400, 1415034000, 1415037600, 1415041200, 
    1415044800, 1415048400, 1415052000, 1415055600, 1415059200, 1415062800, 
    1415066400, 1415070000, 1415073600, 1415077200, 1415080800, 1415084400, 
    1415088000, 1415091600, 1415095200, 1415098800, 1415102400, 1415106000, 
    1415109600, 1415113200, 1415116800, 1415120400, 1415124000, 1415127600, 
    1415131200, 1415134800, 1415138400, 1415142000, 1415145600, 1415149200, 
    1415152800, 1415156400, 1415160000, 1415163600, 1415167200, 1415170800, 
    1415174400, 1415178000, 1415181600, 1415185200, 1415188800, 1415192400, 
    1415196000, 1415199600, 1415203200, 1415206800, 1415210400, 1415214000, 
    1415217600, 1415221200, 1415224800, 1415228400, 1415232000, 1415235600, 
    1415239200, 1415242800, 1415246400, 1415250000, 1415253600, 1415257200, 
    1415260800, 1415264400, 1415268000, 1415271600, 1415275200, 1415278800, 
    1415282400, 1415286000, 1415289600, 1415293200, 1415296800, 1415300400, 
    1415304000, 1415307600, 1415311200, 1415314800, 1415318400, 1415322000, 
    1415325600, 1415329200, 1415332800, 1415336400, 1415340000, 1415343600, 
    1415347200, 1415350800, 1415354400, 1415358000, 1415361600, 1415365200, 
    1415368800, 1415372400, 1415376000, 1415379600, 1415383200, 1415386800, 
    1415390400, 1415394000, 1415397600, 1415401200, 1415404800, 1415408400, 
    1415412000, 1415415600, 1415419200, 1415422800, 1415426400, 1415430000, 
    1415433600, 1415437200, 1415440800, 1415444400, 1415448000, 1415451600, 
    1415455200, 1415458800, 1415462400, 1415466000, 1415469600, 1415473200, 
    1415476800, 1415480400, 1415484000, 1415487600, 1415491200, 1415494800, 
    1415498400, 1415502000, 1415505600, 1415509200, 1415512800, 1415516400, 
    1415520000, 1415523600, 1415527200, 1415530800, 1415534400, 1415538000, 
    1415541600, 1415545200, 1415548800, 1415552400, 1415556000, 1415559600, 
    1415563200, 1415566800, 1415570400, 1415574000, 1415577600, 1415581200, 
    1415584800, 1415588400, 1415592000, 1415595600, 1415599200, 1415602800, 
    1415606400, 1415610000, 1415613600, 1415617200, 1415620800, 1415624400, 
    1415628000, 1415631600, 1415635200, 1415638800, 1415642400, 1415646000, 
    1415649600, 1415653200, 1415656800, 1415660400, 1415664000, 1415667600, 
    1415671200, 1415674800, 1415678400, 1415682000, 1415685600, 1415689200, 
    1415692800, 1415696400, 1415700000, 1415703600, 1415707200, 1415710800, 
    1415714400, 1415718000, 1415721600, 1415725200, 1415728800, 1415732400, 
    1415736000, 1415739600, 1415743200, 1415746800, 1415750400, 1415754000, 
    1415757600, 1415761200, 1415764800, 1415768400, 1415772000, 1415775600, 
    1415779200, 1415782800, 1415786400, 1415790000, 1415793600, 1415797200, 
    1415800800, 1415804400, 1415808000, 1415811600, 1415815200, 1415818800, 
    1415822400, 1415826000, 1415829600, 1415833200, 1415836800, 1415840400, 
    1415844000, 1415847600, 1415851200, 1415854800, 1415858400, 1415862000, 
    1415865600, 1415869200, 1415872800, 1415876400, 1415880000, 1415883600, 
    1415887200, 1415890800, 1415894400, 1415898000, 1415901600, 1415905200, 
    1415908800, 1415912400, 1415916000, 1415919600, 1415923200, 1415926800, 
    1415930400, 1415934000, 1415937600, 1415941200, 1415944800, 1415948400, 
    1415952000, 1415955600, 1415959200, 1415962800, 1415966400, 1415970000, 
    1415973600, 1415977200, 1415980800, 1415984400, 1415988000, 1415991600, 
    1415995200, 1415998800, 1416002400, 1416006000, 1416009600, 1416013200, 
    1416016800, 1416020400, 1416024000, 1416027600, 1416031200, 1416034800, 
    1416038400, 1416042000, 1416045600, 1416049200, 1416052800, 1416056400, 
    1416060000, 1416063600, 1416067200, 1416070800, 1416074400, 1416078000, 
    1416081600, 1416085200, 1416088800, 1416092400, 1416096000, 1416099600, 
    1416103200, 1416106800, 1416110400, 1416114000, 1416117600, 1416121200, 
    1416124800, 1416128400, 1416132000, 1416135600, 1416139200, 1416142800, 
    1416146400, 1416150000, 1416153600, 1416157200, 1416160800, 1416164400, 
    1416168000, 1416171600, 1416175200, 1416178800, 1416182400, 1416186000, 
    1416189600, 1416193200, 1416196800, 1416200400, 1416204000, 1416207600, 
    1416211200, 1416214800, 1416218400, 1416222000, 1416225600, 1416229200, 
    1416232800, 1416236400, 1416240000, 1416243600, 1416247200, 1416250800, 
    1416254400, 1416258000, 1416261600, 1416265200, 1416268800, 1416272400, 
    1416276000, 1416279600, 1416283200, 1416286800, 1416290400, 1416294000, 
    1416297600, 1416301200, 1416304800, 1416308400, 1416312000, 1416315600, 
    1416319200, 1416322800, 1416326400, 1416330000, 1416333600, 1416337200, 
    1416340800, 1416344400, 1416348000, 1416351600, 1416355200, 1416358800, 
    1416362400, 1416366000, 1416369600, 1416373200, 1416376800, 1416380400, 
    1416384000, 1416387600, 1416391200, 1416394800, 1416398400, 1416402000, 
    1416405600, 1416409200, 1416412800, 1416416400, 1416420000, 1416423600, 
    1416427200, 1416430800, 1416434400, 1416438000, 1416441600, 1416445200, 
    1416448800, 1416452400, 1416456000, 1416459600, 1416463200, 1416466800, 
    1416470400, 1416474000, 1416477600, 1416481200, 1416484800, 1416488400, 
    1416492000, 1416495600, 1416499200, 1416502800, 1416506400, 1416510000, 
    1416513600, 1416517200, 1416520800, 1416524400, 1416528000, 1416531600, 
    1416535200, 1416538800, 1416542400, 1416546000, 1416549600, 1416553200, 
    1416556800, 1416560400, 1416564000, 1416567600, 1416571200, 1416574800, 
    1416578400, 1416582000, 1416585600, 1416589200, 1416592800, 1416596400, 
    1416600000, 1416603600, 1416607200, 1416610800, 1416614400, 1416618000, 
    1416621600, 1416625200, 1416628800, 1416632400, 1416636000, 1416639600, 
    1416643200, 1416646800, 1416650400, 1416654000, 1416657600, 1416661200, 
    1416664800, 1416668400, 1416672000, 1416675600, 1416679200, 1416682800, 
    1416686400, 1416690000, 1416693600, 1416697200, 1416700800, 1416704400, 
    1416708000, 1416711600, 1416715200, 1416718800, 1416722400, 1416726000, 
    1416729600, 1416733200, 1416736800, 1416740400, 1416744000, 1416747600, 
    1416751200, 1416754800, 1416758400, 1416762000, 1416765600, 1416769200, 
    1416772800, 1416776400, 1416780000, 1416783600, 1416787200, 1416790800, 
    1416794400, 1416798000, 1416801600, 1416805200, 1416808800, 1416812400, 
    1416816000, 1416819600, 1416823200, 1416826800, 1416830400, 1416834000, 
    1416837600, 1416841200, 1416844800, 1416848400, 1416852000, 1416855600, 
    1416859200, 1416862800, 1416866400, 1416870000, 1416873600, 1416877200, 
    1416880800, 1416884400, 1416888000, 1416891600, 1416895200, 1416898800, 
    1416902400, 1416906000, 1416909600, 1416913200, 1416916800, 1416920400, 
    1416924000, 1416927600, 1416931200, 1416934800, 1416938400, 1416942000, 
    1416945600, 1416949200, 1416952800, 1416956400, 1416960000, 1416963600, 
    1416967200, 1416970800, 1416974400, 1416978000, 1416981600, 1416985200, 
    1416988800, 1416992400, 1416996000, 1416999600, 1417003200, 1417006800, 
    1417010400, 1417014000, 1417017600, 1417021200, 1417024800, 1417028400, 
    1417032000, 1417035600, 1417039200, 1417042800, 1417046400, 1417050000, 
    1417053600, 1417057200, 1417060800, 1417064400, 1417068000, 1417071600, 
    1417075200, 1417078800, 1417082400, 1417086000, 1417089600, 1417093200, 
    1417096800, 1417100400, 1417104000, 1417107600, 1417111200, 1417114800, 
    1417118400, 1417122000, 1417125600, 1417129200, 1417132800, 1417136400, 
    1417140000, 1417143600, 1417147200, 1417150800, 1417154400, 1417158000, 
    1417161600, 1417165200, 1417168800, 1417172400, 1417176000, 1417179600, 
    1417183200, 1417186800, 1417190400, 1417194000, 1417197600, 1417201200, 
    1417204800, 1417208400, 1417212000, 1417215600, 1417219200, 1417222800, 
    1417226400, 1417230000, 1417233600, 1417237200, 1417240800, 1417244400, 
    1417248000, 1417251600, 1417255200, 1417258800, 1417262400, 1417266000, 
    1417269600, 1417273200, 1417276800, 1417280400, 1417284000, 1417287600, 
    1417291200, 1417294800, 1417298400, 1417302000, 1417305600, 1417309200, 
    1417312800, 1417316400, 1417320000, 1417323600, 1417327200, 1417330800, 
    1417334400, 1417338000, 1417341600, 1417345200, 1417348800, 1417352400, 
    1417356000, 1417359600, 1417363200, 1417366800, 1417370400, 1417374000, 
    1417377600, 1417381200, 1417384800, 1417388400, 1417392000, 1417395600, 
    1417399200, 1417402800, 1417406400, 1417410000, 1417413600, 1417417200, 
    1417420800, 1417424400, 1417428000, 1417431600, 1417435200, 1417438800, 
    1417442400, 1417446000, 1417449600, 1417453200, 1417456800, 1417460400, 
    1417464000, 1417467600, 1417471200, 1417474800, 1417478400, 1417482000, 
    1417485600, 1417489200, 1417492800, 1417496400, 1417500000, 1417503600, 
    1417507200, 1417510800, 1417514400, 1417518000, 1417521600, 1417525200, 
    1417528800, 1417532400, 1417536000, 1417539600, 1417543200, 1417546800, 
    1417550400, 1417554000, 1417557600, 1417561200, 1417564800, 1417568400, 
    1417572000, 1417575600, 1417579200, 1417582800, 1417586400, 1417590000, 
    1417593600, 1417597200, 1417600800, 1417604400, 1417608000, 1417611600, 
    1417615200, 1417618800, 1417622400, 1417626000, 1417629600, 1417633200, 
    1417636800, 1417640400, 1417644000, 1417647600, 1417651200, 1417654800, 
    1417658400, 1417662000, 1417665600, 1417669200, 1417672800, 1417676400, 
    1417680000, 1417683600, 1417687200, 1417690800, 1417694400, 1417698000, 
    1417701600, 1417705200, 1417708800, 1417712400, 1417716000, 1417719600, 
    1417723200, 1417726800, 1417730400, 1417734000, 1417737600, 1417741200, 
    1417744800, 1417748400, 1417752000, 1417755600, 1417759200, 1417762800, 
    1417766400, 1417770000, 1417773600, 1417777200, 1417780800, 1417784400, 
    1417788000, 1417791600, 1417795200, 1417798800, 1417802400, 1417806000, 
    1417809600, 1417813200, 1417816800, 1417820400, 1417824000, 1417827600, 
    1417831200, 1417834800, 1417838400, 1417842000, 1417845600, 1417849200, 
    1417852800, 1417856400, 1417860000, 1417863600, 1417867200, 1417870800, 
    1417874400, 1417878000, 1417881600, 1417885200, 1417888800, 1417892400, 
    1417896000, 1417899600, 1417903200, 1417906800, 1417910400, 1417914000, 
    1417917600, 1417921200, 1417924800, 1417928400, 1417932000, 1417935600, 
    1417939200, 1417942800, 1417946400, 1417950000, 1417953600, 1417957200, 
    1417960800, 1417964400, 1417968000, 1417971600, 1417975200, 1417978800, 
    1417982400, 1417986000, 1417989600, 1417993200, 1417996800, 1418000400, 
    1418004000, 1418007600, 1418011200, 1418014800, 1418018400, 1418022000, 
    1418025600, 1418029200, 1418032800, 1418036400, 1418040000, 1418043600, 
    1418047200, 1418050800, 1418054400, 1418058000, 1418061600, 1418065200, 
    1418068800, 1418072400, 1418076000, 1418079600, 1418083200, 1418086800, 
    1418090400, 1418094000, 1418097600, 1418101200, 1418104800, 1418108400, 
    1418112000, 1418115600, 1418119200, 1418122800, 1418126400, 1418130000, 
    1418133600, 1418137200, 1418140800, 1418144400, 1418148000, 1418151600, 
    1418155200, 1418158800, 1418162400, 1418166000, 1418169600, 1418173200, 
    1418176800, 1418180400, 1418184000, 1418187600, 1418191200, 1418194800, 
    1418198400, 1418202000, 1418205600, 1418209200, 1418212800, 1418216400, 
    1418220000, 1418223600, 1418227200, 1418230800, 1418234400, 1418238000, 
    1418241600, 1418245200, 1418248800, 1418252400, 1418256000, 1418259600, 
    1418263200, 1418266800, 1418270400, 1418274000, 1418277600, 1418281200, 
    1418284800, 1418288400, 1418292000, 1418295600, 1418299200, 1418302800, 
    1418306400, 1418310000, 1418313600, 1418317200, 1418320800, 1418324400, 
    1418328000, 1418331600, 1418335200, 1418338800, 1418342400, 1418346000, 
    1418349600, 1418353200, 1418356800, 1418360400, 1418364000, 1418367600, 
    1418371200, 1418374800, 1418378400, 1418382000, 1418385600, 1418389200, 
    1418392800, 1418396400, 1418400000, 1418403600, 1418407200, 1418410800, 
    1418414400, 1418418000, 1418421600, 1418425200, 1418428800, 1418432400, 
    1418436000, 1418439600, 1418443200, 1418446800, 1418450400, 1418454000, 
    1418457600, 1418461200, 1418464800, 1418468400, 1418472000, 1418475600, 
    1418479200, 1418482800, 1418486400, 1418490000, 1418493600, 1418497200, 
    1418500800, 1418504400, 1418508000, 1418511600, 1418515200, 1418518800, 
    1418522400, 1418526000, 1418529600, 1418533200, 1418536800, 1418540400, 
    1418544000, 1418547600, 1418551200, 1418554800, 1418558400, 1418562000, 
    1418565600, 1418569200, 1418572800, 1418576400, 1418580000, 1418583600, 
    1418587200, 1418590800, 1418594400, 1418598000, 1418601600, 1418605200, 
    1418608800, 1418612400, 1418616000, 1418619600, 1418623200, 1418626800, 
    1418630400, 1418634000, 1418637600, 1418641200, 1418644800, 1418648400, 
    1418652000, 1418655600, 1418659200, 1418662800, 1418666400, 1418670000, 
    1418673600, 1418677200, 1418680800, 1418684400, 1418688000, 1418691600, 
    1418695200, 1418698800, 1418702400, 1418706000, 1418709600, 1418713200, 
    1418716800, 1418720400, 1418724000, 1418727600, 1418731200, 1418734800, 
    1418738400, 1418742000, 1418745600, 1418749200, 1418752800, 1418756400, 
    1418760000, 1418763600, 1418767200, 1418770800, 1418774400, 1418778000, 
    1418781600, 1418785200, 1418788800, 1418792400, 1418796000, 1418799600, 
    1418803200, 1418806800, 1418810400, 1418814000, 1418817600, 1418821200, 
    1418824800, 1418828400, 1418832000, 1418835600, 1418839200, 1418842800, 
    1418846400, 1418850000, 1418853600, 1418857200, 1418860800, 1418864400, 
    1418868000, 1418871600, 1418875200, 1418878800, 1418882400, 1418886000, 
    1418889600, 1418893200, 1418896800, 1418900400, 1418904000, 1418907600, 
    1418911200, 1418914800, 1418918400, 1418922000, 1418925600, 1418929200, 
    1418932800, 1418936400, 1418940000, 1418943600, 1418947200, 1418950800, 
    1418954400, 1418958000, 1418961600, 1418965200, 1418968800, 1418972400, 
    1418976000, 1418979600, 1418983200, 1418986800, 1418990400, 1418994000, 
    1418997600, 1419001200, 1419004800, 1419008400, 1419012000, 1419015600, 
    1419019200, 1419022800, 1419026400, 1419030000, 1419033600, 1419037200, 
    1419040800, 1419044400, 1419048000, 1419051600, 1419055200, 1419058800, 
    1419062400, 1419066000, 1419069600, 1419073200, 1419076800, 1419080400, 
    1419084000, 1419087600, 1419091200, 1419094800, 1419098400, 1419102000, 
    1419105600, 1419109200, 1419112800, 1419116400, 1419120000, 1419123600, 
    1419127200, 1419130800, 1419134400, 1419138000, 1419141600, 1419145200, 
    1419148800, 1419152400, 1419156000, 1419159600, 1419163200, 1419166800, 
    1419170400, 1419174000, 1419177600, 1419181200, 1419184800, 1419188400, 
    1419192000, 1419195600, 1419199200, 1419202800, 1419206400, 1419210000, 
    1419213600, 1419217200, 1419220800, 1419224400, 1419228000, 1419231600, 
    1419235200, 1419238800, 1419242400, 1419246000, 1419249600, 1419253200, 
    1419256800, 1419260400, 1419264000, 1419267600, 1419271200, 1419274800, 
    1419278400, 1419282000, 1419285600, 1419289200, 1419292800, 1419296400, 
    1419300000, 1419303600, 1419307200, 1419310800, 1419314400, 1419318000, 
    1419321600, 1419325200, 1419328800, 1419332400, 1419336000, 1419339600, 
    1419343200, 1419346800, 1419350400, 1419354000, 1419357600, 1419361200, 
    1419364800, 1419368400, 1419372000, 1419375600, 1419379200, 1419382800, 
    1419386400, 1419390000, 1419393600, 1419397200, 1419400800, 1419404400, 
    1419408000, 1419411600, 1419415200, 1419418800, 1419422400, 1419426000, 
    1419429600, 1419433200, 1419436800, 1419440400, 1419444000, 1419447600, 
    1419451200, 1419454800, 1419458400, 1419462000, 1419465600, 1419469200, 
    1419472800, 1419476400, 1419480000, 1419483600, 1419487200, 1419490800, 
    1419494400, 1419498000, 1419501600, 1419505200, 1419508800, 1419512400, 
    1419516000, 1419519600, 1419523200, 1419526800, 1419530400, 1419534000, 
    1419537600, 1419541200, 1419544800, 1419548400, 1419552000, 1419555600, 
    1419559200, 1419562800, 1419566400, 1419570000, 1419573600, 1419577200, 
    1419580800, 1419584400, 1419588000, 1419591600, 1419595200, 1419598800, 
    1419602400, 1419606000, 1419609600, 1419613200, 1419616800, 1419620400, 
    1419624000, 1419627600, 1419631200, 1419634800, 1419638400, 1419642000, 
    1419645600, 1419649200, 1419652800, 1419656400, 1419660000, 1419663600, 
    1419667200, 1419670800, 1419674400, 1419678000, 1419681600, 1419685200, 
    1419688800, 1419692400, 1419696000, 1419699600, 1419703200, 1419706800, 
    1419710400, 1419714000, 1419717600, 1419721200, 1419724800, 1419728400, 
    1419732000, 1419735600, 1419739200, 1419742800, 1419746400, 1419750000, 
    1419753600, 1419757200, 1419760800, 1419764400, 1419768000, 1419771600, 
    1419775200, 1419778800, 1419782400, 1419786000, 1419789600, 1419793200, 
    1419796800, 1419800400, 1419804000, 1419807600, 1419811200, 1419814800, 
    1419818400, 1419822000, 1419825600, 1419829200, 1419832800, 1419836400, 
    1419840000, 1419843600, 1419847200, 1419850800, 1419854400, 1419858000, 
    1419861600, 1419865200, 1419868800, 1419872400, 1419876000, 1419879600, 
    1419883200, 1419886800, 1419890400, 1419894000, 1419897600, 1419901200, 
    1419904800, 1419908400, 1419912000, 1419915600, 1419919200, 1419922800, 
    1419926400, 1419930000, 1419933600, 1419937200, 1419940800, 1419944400, 
    1419948000, 1419951600, 1419955200, 1419958800, 1419962400, 1419966000, 
    1419969600, 1419973200, 1419976800, 1419980400, 1419984000, 1419987600, 
    1419991200, 1419994800, 1419998400, 1420002000, 1420005600, 1420009200, 
    1420012800, 1420016400, 1420020000, 1420023600, 1420027200, 1420030800, 
    1420034400, 1420038000, 1420041600, 1420045200, 1420048800, 1420052400, 
    1420056000, 1420059600, 1420063200, 1420066800, 1420070400, 1420074000, 
    1420077600, 1420081200, 1420084800, 1420088400, 1420092000, 1420095600, 
    1420099200, 1420102800, 1420106400, 1420110000, 1420113600, 1420117200, 
    1420120800, 1420124400, 1420128000, 1420131600, 1420135200, 1420138800, 
    1420142400, 1420146000, 1420149600, 1420153200, 1420156800, 1420160400, 
    1420164000, 1420167600, 1420171200, 1420174800, 1420178400, 1420182000, 
    1420185600, 1420189200, 1420192800, 1420196400, 1420200000, 1420203600, 
    1420207200, 1420210800, 1420214400, 1420218000, 1420221600, 1420225200, 
    1420228800, 1420232400, 1420236000, 1420239600, 1420243200, 1420246800, 
    1420250400, 1420254000, 1420257600, 1420261200, 1420264800, 1420268400, 
    1420272000, 1420275600, 1420279200, 1420282800, 1420286400, 1420290000, 
    1420293600, 1420297200, 1420300800, 1420304400, 1420308000, 1420311600, 
    1420315200, 1420318800, 1420322400, 1420326000, 1420329600, 1420333200, 
    1420336800, 1420340400, 1420344000, 1420347600, 1420351200, 1420354800, 
    1420358400, 1420362000, 1420365600, 1420369200, 1420372800, 1420376400, 
    1420380000, 1420383600, 1420387200, 1420390800, 1420394400, 1420398000, 
    1420401600, 1420405200, 1420408800, 1420412400, 1420416000, 1420419600, 
    1420423200, 1420426800, 1420430400, 1420434000, 1420437600, 1420441200, 
    1420444800, 1420448400, 1420452000, 1420455600, 1420459200, 1420462800, 
    1420466400, 1420470000, 1420473600, 1420477200, 1420480800, 1420484400, 
    1420488000, 1420491600, 1420495200, 1420498800, 1420502400, 1420506000, 
    1420509600, 1420513200, 1420516800, 1420520400, 1420524000, 1420527600, 
    1420531200, 1420534800, 1420538400, 1420542000, 1420545600, 1420549200, 
    1420552800, 1420556400, 1420560000, 1420563600, 1420567200, 1420570800, 
    1420574400, 1420578000, 1420581600, 1420585200, 1420588800, 1420592400, 
    1420596000, 1420599600, 1420603200, 1420606800, 1420610400, 1420614000, 
    1420617600, 1420621200, 1420624800, 1420628400, 1420632000, 1420635600, 
    1420639200, 1420642800, 1420646400, 1420650000, 1420653600, 1420657200, 
    1420660800, 1420664400, 1420668000, 1420671600, 1420675200, 1420678800, 
    1420682400, 1420686000, 1420689600, 1420693200, 1420696800, 1420700400, 
    1420704000, 1420707600, 1420711200, 1420714800, 1420718400, 1420722000, 
    1420725600, 1420729200, 1420732800, 1420736400, 1420740000, 1420743600, 
    1420747200, 1420750800, 1420754400, 1420758000, 1420761600, 1420765200, 
    1420768800, 1420772400, 1420776000, 1420779600, 1420783200, 1420786800, 
    1420790400, 1420794000, 1420797600, 1420801200, 1420804800, 1420808400, 
    1420812000, 1420815600, 1420819200, 1420822800, 1420826400, 1420830000, 
    1420833600, 1420837200, 1420840800, 1420844400, 1420848000, 1420851600, 
    1420855200, 1420858800, 1420862400, 1420866000, 1420869600, 1420873200, 
    1420876800, 1420880400, 1420884000, 1420887600, 1420891200, 1420894800, 
    1420898400, 1420902000, 1420905600, 1420909200, 1420912800, 1420916400, 
    1420920000, 1420923600, 1420927200, 1420930800, 1420934400, 1420938000, 
    1420941600, 1420945200, 1420948800, 1420952400, 1420956000, 1420959600, 
    1420963200, 1420966800, 1420970400, 1420974000, 1420977600, 1420981200, 
    1420984800, 1420988400, 1420992000, 1420995600, 1420999200, 1421002800, 
    1421006400, 1421010000, 1421013600, 1421017200, 1421020800, 1421024400, 
    1421028000, 1421031600, 1421035200, 1421038800, 1421042400, 1421046000, 
    1421049600, 1421053200, 1421056800, 1421060400, 1421064000, 1421067600, 
    1421071200, 1421074800, 1421078400, 1421082000, 1421085600, 1421089200, 
    1421092800, 1421096400, 1421100000, 1421103600, 1421107200, 1421110800, 
    1421114400, 1421118000, 1421121600, 1421125200, 1421128800, 1421132400, 
    1421136000, 1421139600, 1421143200, 1421146800, 1421150400, 1421154000, 
    1421157600, 1421161200, 1421164800, 1421168400, 1421172000, 1421175600, 
    1421179200, 1421182800, 1421186400, 1421190000, 1421193600, 1421197200, 
    1421200800, 1421204400, 1421208000, 1421211600, 1421215200, 1421218800, 
    1421222400, 1421226000, 1421229600, 1421233200, 1421236800, 1421240400, 
    1421244000, 1421247600, 1421251200, 1421254800, 1421258400, 1421262000, 
    1421265600, 1421269200, 1421272800, 1421276400, 1421280000, 1421283600, 
    1421287200, 1421290800, 1421294400, 1421298000, 1421301600, 1421305200, 
    1421308800, 1421312400, 1421316000, 1421319600, 1421323200, 1421326800, 
    1421330400, 1421334000, 1421337600, 1421341200, 1421344800, 1421348400, 
    1421352000, 1421355600, 1421359200, 1421362800, 1421366400, 1421370000, 
    1421373600, 1421377200, 1421380800, 1421384400, 1421388000, 1421391600, 
    1421395200, 1421398800, 1421402400, 1421406000, 1421409600, 1421413200, 
    1421416800, 1421420400, 1421424000, 1421427600, 1421431200, 1421434800, 
    1421438400, 1421442000, 1421445600, 1421449200, 1421452800, 1421456400, 
    1421460000, 1421463600, 1421467200, 1421470800, 1421474400, 1421478000, 
    1421481600, 1421485200, 1421488800, 1421492400, 1421496000, 1421499600, 
    1421503200, 1421506800, 1421510400, 1421514000, 1421517600, 1421521200, 
    1421524800, 1421528400, 1421532000, 1421535600, 1421539200, 1421542800, 
    1421546400, 1421550000, 1421553600, 1421557200, 1421560800, 1421564400, 
    1421568000, 1421571600, 1421575200, 1421578800, 1421582400, 1421586000, 
    1421589600, 1421593200, 1421596800, 1421600400, 1421604000, 1421607600, 
    1421611200, 1421614800, 1421618400, 1421622000, 1421625600, 1421629200, 
    1421632800, 1421636400, 1421640000, 1421643600, 1421647200, 1421650800, 
    1421654400, 1421658000, 1421661600, 1421665200, 1421668800, 1421672400, 
    1421676000, 1421679600, 1421683200, 1421686800, 1421690400, 1421694000, 
    1421697600, 1421701200, 1421704800, 1421708400, 1421712000, 1421715600, 
    1421719200, 1421722800, 1421726400, 1421730000, 1421733600, 1421737200, 
    1421740800, 1421744400, 1421748000, 1421751600, 1421755200, 1421758800, 
    1421762400, 1421766000, 1421769600, 1421773200, 1421776800, 1421780400, 
    1421784000, 1421787600, 1421791200, 1421794800, 1421798400, 1421802000, 
    1421805600, 1421809200, 1421812800, 1421816400, 1421820000, 1421823600, 
    1421827200, 1421830800, 1421834400, 1421838000, 1421841600, 1421845200, 
    1421848800, 1421852400, 1421856000, 1421859600, 1421863200, 1421866800, 
    1421870400, 1421874000, 1421877600, 1421881200, 1421884800, 1421888400, 
    1421892000, 1421895600, 1421899200, 1421902800, 1421906400, 1421910000, 
    1421913600, 1421917200, 1421920800, 1421924400, 1421928000, 1421931600, 
    1421935200, 1421938800, 1421942400, 1421946000, 1421949600, 1421953200, 
    1421956800, 1421960400, 1421964000, 1421967600, 1421971200, 1421974800, 
    1421978400, 1421982000, 1421985600, 1421989200, 1421992800, 1421996400, 
    1422000000, 1422003600, 1422007200, 1422010800, 1422014400, 1422018000, 
    1422021600, 1422025200, 1422028800, 1422032400, 1422036000, 1422039600, 
    1422043200, 1422046800, 1422050400, 1422054000, 1422057600, 1422061200, 
    1422064800, 1422068400, 1422072000, 1422075600, 1422079200, 1422082800, 
    1422086400, 1422090000, 1422093600, 1422097200, 1422100800, 1422104400, 
    1422108000, 1422111600, 1422115200, 1422118800, 1422122400, 1422126000, 
    1422129600, 1422133200, 1422136800, 1422140400, 1422144000, 1422147600, 
    1422151200, 1422154800, 1422158400, 1422162000, 1422165600, 1422169200, 
    1422172800, 1422176400, 1422180000, 1422183600, 1422187200, 1422190800, 
    1422194400, 1422198000, 1422201600, 1422205200, 1422208800, 1422212400, 
    1422216000, 1422219600, 1422223200, 1422226800, 1422230400, 1422234000, 
    1422237600, 1422241200, 1422244800, 1422248400, 1422252000, 1422255600, 
    1422259200, 1422262800, 1422266400, 1422270000, 1422273600, 1422277200, 
    1422280800, 1422284400, 1422288000, 1422291600, 1422295200, 1422298800, 
    1422302400, 1422306000, 1422309600, 1422313200, 1422316800, 1422320400, 
    1422324000, 1422327600, 1422331200, 1422334800, 1422338400, 1422342000, 
    1422345600, 1422349200, 1422352800, 1422356400, 1422360000, 1422363600, 
    1422367200, 1422370800, 1422374400, 1422378000, 1422381600, 1422385200, 
    1422388800, 1422392400, 1422396000, 1422399600, 1422403200, 1422406800, 
    1422410400, 1422414000, 1422417600, 1422421200, 1422424800, 1422428400, 
    1422432000, 1422435600, 1422439200, 1422442800, 1422446400, 1422450000, 
    1422453600, 1422457200, 1422460800, 1422464400, 1422468000, 1422471600, 
    1422475200, 1422478800, 1422482400, 1422486000, 1422489600, 1422493200, 
    1422496800, 1422500400, 1422504000, 1422507600, 1422511200, 1422514800, 
    1422518400, 1422522000, 1422525600, 1422529200, 1422532800, 1422536400, 
    1422540000, 1422543600, 1422547200, 1422550800, 1422554400, 1422558000, 
    1422561600, 1422565200, 1422568800, 1422572400, 1422576000, 1422579600, 
    1422583200, 1422586800, 1422590400, 1422594000, 1422597600, 1422601200, 
    1422604800, 1422608400, 1422612000, 1422615600, 1422619200, 1422622800, 
    1422626400, 1422630000, 1422633600, 1422637200, 1422640800, 1422644400, 
    1422648000, 1422651600, 1422655200, 1422658800, 1422662400, 1422666000, 
    1422669600, 1422673200, 1422676800, 1422680400, 1422684000, 1422687600, 
    1422691200, 1422694800, 1422698400, 1422702000, 1422705600, 1422709200, 
    1422712800, 1422716400, 1422720000, 1422723600, 1422727200, 1422730800, 
    1422734400, 1422738000, 1422741600, 1422745200, 1422748800, 1422752400, 
    1422756000, 1422759600, 1422763200, 1422766800, 1422770400, 1422774000, 
    1422777600, 1422781200, 1422784800, 1422788400, 1422792000, 1422795600, 
    1422799200, 1422802800, 1422806400, 1422810000, 1422813600, 1422817200, 
    1422820800, 1422824400, 1422828000, 1422831600, 1422835200, 1422838800, 
    1422842400, 1422846000, 1422849600, 1422853200, 1422856800, 1422860400, 
    1422864000, 1422867600, 1422871200, 1422874800, 1422878400, 1422882000, 
    1422885600, 1422889200, 1422892800, 1422896400, 1422900000, 1422903600, 
    1422907200, 1422910800, 1422914400, 1422918000, 1422921600, 1422925200, 
    1422928800, 1422932400, 1422936000, 1422939600, 1422943200, 1422946800, 
    1422950400, 1422954000, 1422957600, 1422961200, 1422964800, 1422968400, 
    1422972000, 1422975600, 1422979200, 1422982800, 1422986400, 1422990000, 
    1422993600, 1422997200, 1423000800, 1423004400, 1423008000, 1423011600, 
    1423015200, 1423018800, 1423022400, 1423026000, 1423029600, 1423033200, 
    1423036800, 1423040400, 1423044000, 1423047600, 1423051200, 1423054800, 
    1423058400, 1423062000, 1423065600, 1423069200, 1423072800, 1423076400, 
    1423080000, 1423083600, 1423087200, 1423090800, 1423094400, 1423098000, 
    1423101600, 1423105200, 1423108800, 1423112400, 1423116000, 1423119600, 
    1423123200, 1423126800, 1423130400, 1423134000, 1423137600, 1423141200, 
    1423144800, 1423148400, 1423152000, 1423155600, 1423159200, 1423162800, 
    1423166400, 1423170000, 1423173600, 1423177200, 1423180800, 1423184400, 
    1423188000, 1423191600, 1423195200, 1423198800, 1423202400, 1423206000, 
    1423209600, 1423213200, 1423216800, 1423220400, 1423224000, 1423227600, 
    1423231200, 1423234800, 1423238400, 1423242000, 1423245600, 1423249200, 
    1423252800, 1423256400, 1423260000, 1423263600, 1423267200, 1423270800, 
    1423274400, 1423278000, 1423281600, 1423285200, 1423288800, 1423292400, 
    1423296000, 1423299600, 1423303200, 1423306800, 1423310400, 1423314000, 
    1423317600, 1423321200, 1423324800, 1423328400, 1423332000, 1423335600, 
    1423339200, 1423342800, 1423346400, 1423350000, 1423353600, 1423357200, 
    1423360800, 1423364400, 1423368000, 1423371600, 1423375200, 1423378800, 
    1423382400, 1423386000, 1423389600, 1423393200, 1423396800, 1423400400, 
    1423404000, 1423407600, 1423411200, 1423414800, 1423418400, 1423422000, 
    1423425600, 1423429200, 1423432800, 1423436400, 1423440000, 1423443600, 
    1423447200, 1423450800, 1423454400, 1423458000, 1423461600, 1423465200, 
    1423468800, 1423472400, 1423476000, 1423479600, 1423483200, 1423486800, 
    1423490400, 1423494000, 1423497600, 1423501200, 1423504800, 1423508400, 
    1423512000, 1423515600, 1423519200, 1423522800, 1423526400, 1423530000, 
    1423533600, 1423537200, 1423540800, 1423544400, 1423548000, 1423551600, 
    1423555200, 1423558800, 1423562400, 1423566000, 1423569600, 1423573200, 
    1423576800, 1423580400, 1423584000, 1423587600, 1423591200, 1423594800, 
    1423598400, 1423602000, 1423605600, 1423609200, 1423612800, 1423616400, 
    1423620000, 1423623600, 1423627200, 1423630800, 1423634400, 1423638000, 
    1423641600, 1423645200, 1423648800, 1423652400, 1423656000, 1423659600, 
    1423663200, 1423666800, 1423670400, 1423674000, 1423677600, 1423681200, 
    1423684800, 1423688400, 1423692000, 1423695600, 1423699200, 1423702800, 
    1423706400, 1423710000, 1423713600, 1423717200, 1423720800, 1423724400, 
    1423728000, 1423731600, 1423735200, 1423738800, 1423742400, 1423746000, 
    1423749600, 1423753200, 1423756800, 1423760400, 1423764000, 1423767600, 
    1423771200, 1423774800, 1423778400, 1423782000, 1423785600, 1423789200, 
    1423792800, 1423796400, 1423800000, 1423803600, 1423807200, 1423810800, 
    1423814400, 1423818000, 1423821600, 1423825200, 1423828800, 1423832400, 
    1423836000, 1423839600, 1423843200, 1423846800, 1423850400, 1423854000, 
    1423857600, 1423861200, 1423864800, 1423868400, 1423872000, 1423875600, 
    1423879200, 1423882800, 1423886400, 1423890000, 1423893600, 1423897200, 
    1423900800, 1423904400, 1423908000, 1423911600, 1423915200, 1423918800, 
    1423922400, 1423926000, 1423929600, 1423933200, 1423936800, 1423940400, 
    1423944000, 1423947600, 1423951200, 1423954800, 1423958400, 1423962000, 
    1423965600, 1423969200, 1423972800, 1423976400, 1423980000, 1423983600, 
    1423987200, 1423990800, 1423994400, 1423998000, 1424001600, 1424005200, 
    1424008800, 1424012400, 1424016000, 1424019600, 1424023200, 1424026800, 
    1424030400, 1424034000, 1424037600, 1424041200, 1424044800, 1424048400, 
    1424052000, 1424055600, 1424059200, 1424062800, 1424066400, 1424070000, 
    1424073600, 1424077200, 1424080800, 1424084400, 1424088000, 1424091600, 
    1424095200, 1424098800, 1424102400, 1424106000, 1424109600, 1424113200, 
    1424116800, 1424120400, 1424124000, 1424127600, 1424131200, 1424134800, 
    1424138400, 1424142000, 1424145600, 1424149200, 1424152800, 1424156400, 
    1424160000, 1424163600, 1424167200, 1424170800, 1424174400, 1424178000, 
    1424181600, 1424185200, 1424188800, 1424192400, 1424196000, 1424199600, 
    1424203200, 1424206800, 1424210400, 1424214000, 1424217600, 1424221200, 
    1424224800, 1424228400, 1424232000, 1424235600, 1424239200, 1424242800, 
    1424246400, 1424250000, 1424253600, 1424257200, 1424260800, 1424264400, 
    1424268000, 1424271600, 1424275200, 1424278800, 1424282400, 1424286000, 
    1424289600, 1424293200, 1424296800, 1424300400, 1424304000, 1424307600, 
    1424311200, 1424314800, 1424318400, 1424322000, 1424325600, 1424329200, 
    1424332800, 1424336400, 1424340000, 1424343600, 1424347200, 1424350800, 
    1424354400, 1424358000, 1424361600, 1424365200, 1424368800, 1424372400, 
    1424376000, 1424379600, 1424383200, 1424386800, 1424390400, 1424394000, 
    1424397600, 1424401200, 1424404800, 1424408400, 1424412000, 1424415600, 
    1424419200, 1424422800, 1424426400, 1424430000, 1424433600, 1424437200, 
    1424440800, 1424444400, 1424448000, 1424451600, 1424455200, 1424458800, 
    1424462400, 1424466000, 1424469600, 1424473200, 1424476800, 1424480400, 
    1424484000, 1424487600, 1424491200, 1424494800, 1424498400, 1424502000, 
    1424505600, 1424509200, 1424512800, 1424516400, 1424520000, 1424523600, 
    1424527200, 1424530800, 1424534400, 1424538000, 1424541600, 1424545200, 
    1424548800, 1424552400, 1424556000, 1424559600, 1424563200, 1424566800, 
    1424570400, 1424574000, 1424577600, 1424581200, 1424584800, 1424588400, 
    1424592000, 1424595600, 1424599200, 1424602800, 1424606400, 1424610000, 
    1424613600, 1424617200, 1424620800, 1424624400, 1424628000, 1424631600, 
    1424635200, 1424638800, 1424642400, 1424646000, 1424649600, 1424653200, 
    1424656800, 1424660400, 1424664000, 1424667600, 1424671200, 1424674800, 
    1424678400, 1424682000, 1424685600, 1424689200, 1424692800, 1424696400, 
    1424700000, 1424703600, 1424707200, 1424710800, 1424714400, 1424718000, 
    1424721600, 1424725200, 1424728800, 1424732400, 1424736000, 1424739600, 
    1424743200, 1424746800, 1424750400, 1424754000, 1424757600, 1424761200, 
    1424764800, 1424768400, 1424772000, 1424775600, 1424779200, 1424782800, 
    1424786400, 1424790000, 1424793600, 1424797200, 1424800800, 1424804400, 
    1424808000, 1424811600, 1424815200, 1424818800, 1424822400, 1424826000, 
    1424829600, 1424833200, 1424836800, 1424840400, 1424844000, 1424847600, 
    1424851200, 1424854800, 1424858400, 1424862000, 1424865600, 1424869200, 
    1424872800, 1424876400, 1424880000, 1424883600, 1424887200, 1424890800, 
    1424894400, 1424898000, 1424901600, 1424905200, 1424908800, 1424912400, 
    1424916000, 1424919600, 1424923200, 1424926800, 1424930400, 1424934000, 
    1424937600, 1424941200, 1424944800, 1424948400, 1424952000, 1424955600, 
    1424959200, 1424962800, 1424966400, 1424970000, 1424973600, 1424977200, 
    1424980800, 1424984400, 1424988000, 1424991600, 1424995200, 1424998800, 
    1425002400, 1425006000, 1425009600, 1425013200, 1425016800, 1425020400, 
    1425024000, 1425027600, 1425031200, 1425034800, 1425038400, 1425042000, 
    1425045600, 1425049200, 1425052800, 1425056400, 1425060000, 1425063600, 
    1425067200, 1425070800, 1425074400, 1425078000, 1425081600, 1425085200, 
    1425088800, 1425092400, 1425096000, 1425099600, 1425103200, 1425106800, 
    1425110400, 1425114000, 1425117600, 1425121200, 1425124800, 1425128400, 
    1425132000, 1425135600, 1425139200, 1425142800, 1425146400, 1425150000, 
    1425153600, 1425157200, 1425160800, 1425164400, 1425168000, 1425171600, 
    1425175200, 1425178800, 1425182400, 1425186000, 1425189600, 1425193200, 
    1425196800, 1425200400, 1425204000, 1425207600, 1425211200, 1425214800, 
    1425218400, 1425222000, 1425225600, 1425229200, 1425232800, 1425236400, 
    1425240000, 1425243600, 1425247200, 1425250800, 1425254400, 1425258000, 
    1425261600, 1425265200, 1425268800, 1425272400, 1425276000, 1425279600, 
    1425283200, 1425286800, 1425290400, 1425294000, 1425297600, 1425301200, 
    1425304800, 1425308400, 1425312000, 1425315600, 1425319200, 1425322800, 
    1425326400, 1425330000, 1425333600, 1425337200, 1425340800, 1425344400, 
    1425348000, 1425351600, 1425355200, 1425358800, 1425362400, 1425366000, 
    1425369600, 1425373200, 1425376800, 1425380400, 1425384000, 1425387600, 
    1425391200, 1425394800, 1425398400, 1425402000, 1425405600, 1425409200, 
    1425412800, 1425416400, 1425420000, 1425423600, 1425427200, 1425430800, 
    1425434400, 1425438000, 1425441600, 1425445200, 1425448800, 1425452400, 
    1425456000, 1425459600, 1425463200, 1425466800, 1425470400, 1425474000, 
    1425477600, 1425481200, 1425484800, 1425488400, 1425492000, 1425495600, 
    1425499200, 1425502800, 1425506400, 1425510000, 1425513600, 1425517200, 
    1425520800, 1425524400, 1425528000, 1425531600, 1425535200, 1425538800, 
    1425542400, 1425546000, 1425549600, 1425553200, 1425556800, 1425560400, 
    1425564000, 1425567600, 1425571200, 1425574800, 1425578400, 1425582000, 
    1425585600, 1425589200, 1425592800, 1425596400, 1425600000, 1425603600, 
    1425607200, 1425610800, 1425614400, 1425618000, 1425621600, 1425625200, 
    1425628800, 1425632400, 1425636000, 1425639600, 1425643200, 1425646800, 
    1425650400, 1425654000, 1425657600, 1425661200, 1425664800, 1425668400, 
    1425672000, 1425675600, 1425679200, 1425682800, 1425686400, 1425690000, 
    1425693600, 1425697200, 1425700800, 1425704400, 1425708000, 1425711600, 
    1425715200, 1425718800, 1425722400, 1425726000, 1425729600, 1425733200, 
    1425736800, 1425740400, 1425744000, 1425747600, 1425751200, 1425754800, 
    1425758400, 1425762000, 1425765600, 1425769200, 1425772800, 1425776400, 
    1425780000, 1425783600, 1425787200, 1425790800, 1425794400, 1425798000, 
    1425801600, 1425805200, 1425808800, 1425812400, 1425816000, 1425819600, 
    1425823200, 1425826800, 1425830400, 1425834000, 1425837600, 1425841200, 
    1425844800, 1425848400, 1425852000, 1425855600, 1425859200, 1425862800, 
    1425866400, 1425870000, 1425873600, 1425877200, 1425880800, 1425884400, 
    1425888000, 1425891600, 1425895200, 1425898800, 1425902400, 1425906000, 
    1425909600, 1425913200, 1425916800, 1425920400, 1425924000, 1425927600, 
    1425931200, 1425934800, 1425938400, 1425942000, 1425945600, 1425949200, 
    1425952800, 1425956400, 1425960000, 1425963600, 1425967200, 1425970800, 
    1425974400, 1425981600, 1425985200, 1425988800, 1425992400, 1425996000, 
    1425999600, 1426003200, 1426006800, 1426010400, 1426014000, 1426017600, 
    1426021200, 1426024800, 1426028400, 1426032000, 1426035600, 1426039200, 
    1426042800, 1426046400, 1426050000, 1426053600, 1426057200, 1426060800, 
    1426064400, 1426068000, 1426071600, 1426075200, 1426078800, 1426082400, 
    1426086000, 1426089600, 1426093200, 1426096800, 1426100400, 1426104000, 
    1426107600, 1426111200, 1426114800, 1426118400, 1426122000, 1426125600, 
    1426129200, 1426132800, 1426136400, 1426140000, 1426143600, 1426147200, 
    1426150800, 1426154400, 1426158000, 1426161600, 1426165200, 1426168800, 
    1426172400, 1426176000, 1426179600, 1426183200, 1426186800, 1426190400, 
    1426194000, 1426197600, 1426201200, 1426204800, 1426208400, 1426212000, 
    1426215600, 1426219200, 1426222800, 1426226400, 1426230000, 1426233600, 
    1426237200, 1426240800, 1426244400, 1426248000, 1426251600, 1426255200, 
    1426258800, 1426262400, 1426266000, 1426269600, 1426273200, 1426276800, 
    1426280400, 1426284000, 1426287600, 1426291200, 1426294800, 1426298400, 
    1426302000, 1426305600, 1426309200, 1426312800, 1426316400, 1426320000, 
    1426323600, 1426327200, 1426330800, 1426334400, 1426338000, 1426341600, 
    1426345200, 1426348800, 1426352400, 1426356000, 1426359600, 1426363200, 
    1426366800, 1426370400, 1426374000, 1426377600, 1426381200, 1426384800, 
    1426388400, 1426392000, 1426395600, 1426399200, 1426402800, 1426406400, 
    1426410000, 1426413600, 1426417200, 1426420800, 1426424400, 1426428000, 
    1426431600, 1426435200, 1426438800, 1426442400, 1426446000, 1426449600, 
    1426453200, 1426456800, 1426460400, 1426464000, 1426467600, 1426471200, 
    1426474800, 1426478400, 1426482000, 1426485600, 1426489200, 1426492800, 
    1426496400, 1426500000, 1426503600, 1426507200, 1426510800, 1426514400, 
    1426518000, 1426521600, 1426525200, 1426528800, 1426532400, 1426536000, 
    1426539600, 1426543200, 1426546800, 1426550400, 1426554000, 1426557600, 
    1426561200, 1426564800, 1426568400, 1426572000, 1426575600, 1426579200, 
    1426582800, 1426586400, 1426590000, 1426593600, 1426597200, 1426600800, 
    1426604400, 1426608000, 1426611600, 1426615200, 1426618800, 1426622400, 
    1426626000, 1426629600, 1426633200, 1426636800, 1426640400, 1426644000, 
    1426647600, 1426651200, 1426654800, 1426658400, 1426662000, 1426665600, 
    1426669200, 1426672800, 1426676400, 1426680000, 1426683600, 1426687200, 
    1426690800, 1426694400, 1426698000, 1426701600, 1426705200, 1426708800, 
    1426712400, 1426716000, 1426719600, 1426723200, 1426726800, 1426730400, 
    1426734000, 1426737600, 1426741200, 1426744800, 1426748400, 1426752000, 
    1426755600, 1426759200, 1426762800, 1426766400, 1426770000, 1426773600, 
    1426777200, 1426780800, 1426784400, 1426788000, 1426791600, 1426795200, 
    1426798800, 1426802400, 1426806000, 1426809600, 1426813200, 1426816800, 
    1426820400, 1426824000, 1426827600, 1426831200, 1426834800, 1426838400, 
    1426842000, 1426845600, 1426849200, 1426852800, 1426856400, 1426860000, 
    1426863600, 1426867200, 1426870800, 1426874400, 1426878000, 1426881600, 
    1426885200, 1426888800, 1426892400, 1426896000, 1426899600, 1426903200, 
    1426906800, 1426910400, 1426914000, 1426917600, 1426921200, 1426924800, 
    1426928400, 1426932000, 1426935600, 1426939200, 1426942800, 1426946400, 
    1426950000, 1426953600, 1426957200, 1426960800, 1426964400, 1426968000, 
    1426971600, 1426975200, 1426978800, 1426982400, 1426986000, 1426989600, 
    1426993200, 1426996800, 1427000400, 1427004000, 1427007600, 1427011200, 
    1427014800, 1427018400, 1427022000, 1427025600, 1427029200, 1427032800, 
    1427036400, 1427040000, 1427043600, 1427047200, 1427050800, 1427054400, 
    1427058000, 1427061600, 1427065200, 1427068800, 1427072400, 1427076000, 
    1427079600, 1427083200, 1427086800, 1427090400, 1427094000, 1427097600, 
    1427101200, 1427104800, 1427108400, 1427112000, 1427115600, 1427119200, 
    1427122800, 1427126400, 1427130000, 1427133600, 1427137200, 1427140800, 
    1427144400, 1427148000, 1427151600, 1427155200, 1427158800, 1427162400, 
    1427166000, 1427169600, 1427173200, 1427176800, 1427180400, 1427184000, 
    1427187600, 1427191200, 1427194800, 1427198400, 1427202000, 1427205600, 
    1427209200, 1427212800, 1427216400, 1427220000, 1427223600, 1427227200, 
    1427230800, 1427234400, 1427238000, 1427252400, 1427256000, 1427259600, 
    1427263200, 1427266800, 1427270400, 1427274000, 1427277600, 1427281200, 
    1427284800, 1427288400, 1427292000, 1427295600, 1427299200, 1427302800, 
    1427306400, 1427310000, 1427313600, 1427317200, 1427320800, 1427324400, 
    1427328000, 1427331600, 1427335200, 1427338800, 1427342400, 1427346000, 
    1427349600, 1427353200, 1427356800, 1427360400, 1427364000, 1427367600, 
    1427371200, 1427374800, 1427378400, 1427382000, 1427385600, 1427389200, 
    1427392800, 1427396400, 1427400000, 1427403600, 1427407200, 1427410800, 
    1427414400, 1427418000, 1427421600, 1427425200, 1427428800, 1427432400, 
    1427436000, 1427439600, 1427443200, 1427446800, 1427450400, 1427454000, 
    1427457600, 1427461200, 1427464800, 1427468400, 1427472000, 1427475600, 
    1427479200, 1427482800, 1427486400, 1427490000, 1427493600, 1427497200, 
    1427500800, 1427504400, 1427508000, 1427511600, 1427515200, 1427518800, 
    1427522400, 1427526000, 1427529600, 1427533200, 1427536800, 1427540400, 
    1427544000, 1427547600, 1427551200, 1427554800, 1427558400, 1427562000, 
    1427565600, 1427569200, 1427572800, 1427576400, 1427580000, 1427583600, 
    1427587200, 1427590800, 1427594400, 1427598000, 1427601600, 1427605200, 
    1427608800, 1427612400, 1427616000, 1427619600, 1427623200, 1427626800, 
    1427630400, 1427634000, 1427637600, 1427641200, 1427644800, 1427648400, 
    1427652000, 1427655600, 1427659200, 1427662800, 1427666400, 1427670000, 
    1427673600, 1427677200, 1427680800, 1427684400, 1427688000, 1427691600, 
    1427695200, 1427698800, 1427702400, 1427706000, 1427709600, 1427713200, 
    1427716800, 1427720400, 1427724000, 1427727600, 1427731200, 1427734800, 
    1427738400, 1427742000, 1427745600, 1427749200, 1427752800, 1427756400, 
    1427760000, 1427763600, 1427767200, 1427770800, 1427774400, 1427778000, 
    1427781600, 1427785200, 1427788800, 1427792400, 1427796000, 1427799600, 
    1427803200, 1427806800, 1427810400, 1427814000, 1427817600, 1427821200, 
    1427824800, 1427828400, 1427832000, 1427835600, 1427839200, 1427842800, 
    1427846400, 1427850000, 1427853600, 1427857200, 1427860800, 1427864400, 
    1427868000, 1427871600, 1427875200, 1427878800, 1427882400, 1427886000, 
    1427889600, 1427893200, 1427896800, 1427900400, 1427904000, 1427907600, 
    1427911200, 1427914800, 1427918400, 1427922000, 1427925600, 1427929200, 
    1427932800, 1427936400, 1427940000, 1427943600, 1427947200, 1427950800, 
    1427954400, 1427958000, 1427961600, 1427965200, 1427968800, 1427972400, 
    1427976000, 1427979600, 1427983200, 1427986800, 1427990400, 1427994000, 
    1427997600, 1428001200, 1428004800, 1428008400, 1428012000, 1428015600, 
    1428019200, 1428022800, 1428026400, 1428030000, 1428033600, 1428037200, 
    1428040800, 1428044400, 1428048000, 1428051600, 1428055200, 1428058800, 
    1428062400, 1428066000, 1428069600, 1428073200, 1428076800, 1428080400, 
    1428084000, 1428087600, 1428091200, 1428094800, 1428098400, 1428102000, 
    1428105600, 1428109200, 1428112800, 1428116400, 1428120000, 1428123600, 
    1428127200, 1428130800, 1428134400, 1428138000, 1428141600, 1428145200, 
    1428148800, 1428152400, 1428156000, 1428159600, 1428163200, 1428166800, 
    1428170400, 1428174000, 1428177600, 1428181200, 1428184800, 1428188400, 
    1428192000, 1428195600, 1428199200, 1428202800, 1428206400, 1428210000, 
    1428213600, 1428217200, 1428220800, 1428224400, 1428228000, 1428231600, 
    1428235200, 1428238800, 1428242400, 1428246000, 1428249600, 1428253200, 
    1428256800, 1428260400, 1428264000, 1428267600, 1428271200, 1428274800, 
    1428278400, 1428282000, 1428285600, 1428289200, 1428292800, 1428296400, 
    1428300000, 1428303600, 1428307200, 1428310800, 1428314400, 1428318000, 
    1428321600, 1428325200, 1428328800, 1428332400, 1428336000, 1428339600, 
    1428343200, 1428346800, 1428350400, 1428354000, 1428357600, 1428361200, 
    1428364800, 1428368400, 1428372000, 1428375600, 1428379200, 1428382800, 
    1428386400, 1428390000, 1428393600, 1428397200, 1428400800, 1428404400, 
    1428408000, 1428411600, 1428415200, 1428418800, 1428422400, 1428426000, 
    1428429600, 1428433200, 1428436800, 1428440400, 1428444000, 1428447600, 
    1428451200, 1428454800, 1428458400, 1428462000, 1428465600, 1428469200, 
    1428472800, 1428476400, 1428480000, 1428483600, 1428487200, 1428490800, 
    1428494400, 1428498000, 1428501600, 1428505200, 1428508800, 1428512400, 
    1428516000, 1428519600, 1428523200, 1428526800, 1428530400, 1428534000, 
    1428537600, 1428541200, 1428544800, 1428548400, 1428552000, 1428555600, 
    1428559200, 1428562800, 1428566400, 1428570000, 1428573600, 1428577200, 
    1428580800, 1428584400, 1428588000, 1428591600, 1428595200, 1428598800, 
    1428602400, 1428606000, 1428609600, 1428613200, 1428616800, 1428620400, 
    1428624000, 1428627600, 1428631200, 1428634800, 1428638400, 1428642000, 
    1428645600, 1428649200, 1428652800, 1428656400, 1428660000, 1428663600, 
    1428667200, 1428670800, 1428674400, 1428678000, 1428681600, 1428685200, 
    1428688800, 1428692400, 1428696000, 1428699600, 1428703200, 1428706800, 
    1428710400, 1428714000, 1428717600, 1428721200, 1428724800, 1428728400, 
    1428732000, 1428735600, 1428742800, 1428746400, 1428750000, 1428753600, 
    1428757200, 1428760800, 1428764400, 1428768000, 1428771600, 1428775200, 
    1428778800, 1428782400, 1428786000, 1428789600, 1428793200, 1428796800, 
    1428800400, 1428804000, 1428807600, 1428811200, 1428814800, 1428818400, 
    1428822000, 1428825600, 1428829200, 1428832800, 1428836400, 1428840000, 
    1428843600, 1428847200, 1428850800, 1428854400, 1428858000, 1428861600, 
    1428865200, 1428868800, 1428872400, 1428876000, 1428879600, 1428883200, 
    1428886800, 1428890400, 1428894000, 1428897600, 1428901200, 1428904800, 
    1428908400, 1428912000, 1428915600, 1428919200, 1428922800, 1428926400, 
    1428930000, 1428933600, 1428937200, 1428940800, 1428944400, 1428948000, 
    1428951600, 1428955200, 1428958800, 1428962400, 1428966000, 1428969600, 
    1428973200, 1428976800, 1428980400, 1428984000, 1428987600, 1428991200, 
    1428994800, 1428998400, 1429002000, 1429005600, 1429009200, 1429012800, 
    1429016400, 1429020000, 1429023600, 1429027200, 1429030800, 1429034400, 
    1429038000, 1429041600, 1429045200, 1429048800, 1429052400, 1429056000, 
    1429059600, 1429063200, 1429066800, 1429070400, 1429074000, 1429077600, 
    1429088400, 1429092000, 1429095600, 1429099200, 1429102800, 1429185600, 
    1429189200, 1429192800, 1429196400, 1429200000, 1429203600, 1429207200, 
    1429210800, 1429214400, 1429218000, 1429221600, 1429225200, 1429228800, 
    1429232400, 1429236000, 1429239600, 1429243200, 1429246800, 1429250400, 
    1429254000, 1429261200, 1429264800, 1429268400, 1429272000, 1429275600, 
    1429279200, 1429282800, 1429286400, 1429290000, 1429293600, 1429297200, 
    1429300800, 1429304400, 1429308000, 1429311600, 1429315200, 1429318800, 
    1429322400, 1429326000, 1429329600, 1429333200, 1429336800, 1429344000, 
    1429347600, 1429351200, 1429354800, 1429358400, 1429362000, 1429365600, 
    1429369200, 1429372800, 1429376400, 1429380000, 1429383600, 1429387200, 
    1429390800, 1429394400, 1429398000, 1429401600, 1429405200, 1429408800, 
    1429412400, 1429416000, 1429419600, 1429423200, 1429426800, 1429430400, 
    1429434000, 1429437600, 1429441200, 1429444800, 1429448400, 1429452000, 
    1429455600, 1429459200, 1429462800, 1429466400, 1429470000, 1429473600, 
    1429477200, 1429480800, 1429484400, 1429488000, 1429491600, 1429495200, 
    1429498800, 1429502400, 1429506000, 1429509600, 1429513200, 1429516800, 
    1429520400, 1429524000, 1429527600, 1429531200, 1429534800, 1429538400, 
    1429542000, 1429545600, 1429549200, 1429552800, 1429556400, 1429560000, 
    1429563600, 1429567200, 1429570800, 1429574400, 1429578000, 1429581600, 
    1429585200, 1429588800, 1429592400, 1429596000, 1429599600, 1429603200, 
    1429606800, 1429614000, 1429621200, 1429624800, 1429628400, 1429635600, 
    1429642800, 1429646400, 1429650000, 1429653600, 1429664400, 1429668000, 
    1429671600, 1429675200, 1429678800, 1429682400, 1429686000, 1429689600, 
    1429693200, 1429700400, 1429704000, 1429707600, 1429711200, 1429725600, 
    1429729200, 1429732800, 1429740000, 1429743600, 1429754400, 1429758000, 
    1429761600, 1429765200, 1429772400, 1429776000, 1429783200, 1429786800, 
    1429794000, 1429804800, 1429808400, 1429812000, 1429819200, 1429826400, 
    1429830000, 1429833600, 1429837200, 1429848000, 1429851600, 1429855200, 
    1429862400, 1429866000, 1429869600, 1429873200, 1429884000, 1429887600, 
    1429894800, 1429898400, 1429902000, 1429905600, 1429909200, 1429912800, 
    1429916400, 1429920000, 1429923600, 1429927200, 1429930800, 1429934400, 
    1429938000, 1429941600, 1429948800, 1429966800, 1429974000, 1429984800, 
    1430013600, 1430017200, 1430020800, 1430024400, 1430028000, 1430031600, 
    1430035200, 1430038800, 1430042400, 1430049600, 1430053200, 1430056800, 
    1430060400, 1430064000, 1430067600, 1430074800, 1430085600, 1430103600, 
    1430107200, 1430114400, 1430118000, 1430121600, 1430125200, 1430128800, 
    1430132400, 1430136000, 1430139600, 1430146800, 1430150400, 1430161200, 
    1430164800, 1430168400, 1430172000, 1430175600, 1430182800, 1430186400, 
    1430190000, 1430193600, 1430197200, 1430200800, 1430204400, 1430208000, 
    1430211600, 1430215200, 1430226000, 1430229600, 1430236800, 1430244000, 
    1430247600, 1430254800, 1430258400, 1430262000, 1430272800, 1430283600, 
    1430287200, 1430290800, 1430294400, 1430298000, 1430301600, 1430305200, 
    1430312400, 1430316000, 1430319600, 1430326800, 1430330400, 1430334000, 
    1430337600, 1430341200, 1430344800, 1430348400, 1430352000, 1430355600, 
    1430359200, 1430362800, 1430366400, 1430370000, 1430373600, 1430377200, 
    1430380800, 1430395200, 1430398800, 1430402400, 1430406000, 1430409600, 
    1430413200, 1430416800, 1430427600, 1430434800, 1430438400, 1430445600, 
    1430449200, 1430456400, 1430460000, 1430467200, 1430478000, 1430485200, 
    1430492400, 1430496000, 1430499600, 1430503200, 1430506800, 1430510400, 
    1430514000, 1430546400, 1430550000, 1430553600, 1430557200, 1430564400, 
    1430568000, 1430571600, 1430575200, 1430578800, 1430582400, 1430586000, 
    1430589600, 1430593200, 1430596800, 1430600400, 1430604000, 1430607600, 
    1430611200, 1430614800, 1430618400, 1430622000, 1430625600, 1430629200, 
    1430632800, 1430636400, 1430640000, 1430643600, 1430647200, 1430650800, 
    1430654400, 1430658000, 1430661600, 1430665200, 1430668800, 1430672400, 
    1430722800, 1430726400, 1430730000, 1430733600, 1430737200, 1430740800, 
    1430744400, 1430748000, 1430751600, 1430755200, 1430758800, 1430762400, 
    1430766000, 1430769600, 1430773200, 1430776800, 1430780400, 1430784000, 
    1430787600, 1430791200, 1430794800, 1430798400, 1430802000, 1430805600, 
    1430809200, 1430812800, 1430816400, 1430820000, 1430823600, 1430827200, 
    1430830800, 1430834400, 1430838000, 1430841600, 1430845200, 1430848800, 
    1430852400, 1430856000, 1430859600, 1430863200, 1430866800, 1430870400, 
    1430874000, 1430877600, 1430881200, 1430884800, 1430888400, 1430892000, 
    1430895600, 1430899200, 1430902800, 1430906400, 1430910000, 1430913600, 
    1430917200, 1430920800, 1430924400, 1430928000, 1430931600, 1430935200, 
    1430938800, 1430942400, 1430946000, 1430949600, 1430953200, 1430956800, 
    1430960400, 1430964000, 1430967600, 1430971200, 1430974800, 1430978400, 
    1430982000, 1430985600, 1430989200, 1430992800, 1430996400, 1431000000, 
    1431003600, 1431007200, 1431010800, 1431014400, 1431018000, 1431021600, 
    1431025200, 1431028800, 1431032400, 1431036000, 1431039600, 1431043200, 
    1431046800, 1431050400, 1431054000, 1431057600, 1431061200, 1431064800, 
    1431068400, 1431072000, 1431075600, 1431079200, 1431082800, 1431086400, 
    1431090000, 1431093600, 1431097200, 1431100800, 1431104400, 1431108000, 
    1431111600, 1431115200, 1431118800, 1431122400, 1431126000, 1431129600, 
    1431133200, 1431136800, 1431140400, 1431144000, 1431147600, 1431151200, 
    1431154800, 1431158400, 1431162000, 1431165600, 1431169200, 1431172800, 
    1431176400, 1431180000, 1431183600, 1431187200, 1431190800, 1431194400, 
    1431201600, 1431205200, 1431208800, 1431212400, 1431216000, 1431219600, 
    1431223200, 1431226800, 1431230400, 1431234000, 1431237600, 1431241200, 
    1431244800, 1431248400, 1431252000, 1431255600, 1431259200, 1431262800, 
    1431266400, 1431270000, 1431273600, 1431277200, 1431280800, 1431284400, 
    1431288000, 1431291600, 1431295200, 1431298800, 1431302400, 1431306000, 
    1431309600, 1431313200, 1431316800, 1431320400, 1431324000, 1431327600, 
    1431331200, 1431334800, 1431338400, 1431342000, 1431345600, 1431349200, 
    1431352800, 1431356400, 1431360000, 1431363600, 1431367200, 1431370800, 
    1431374400, 1431378000, 1431381600, 1431385200, 1431388800, 1431392400, 
    1431396000, 1431399600, 1431403200, 1431406800, 1431410400, 1431414000, 
    1431417600, 1431421200, 1431424800, 1431428400, 1431435600, 1431439200, 
    1431442800, 1431446400, 1431450000, 1431453600, 1431457200, 1431460800, 
    1431464400, 1431471600, 1431475200, 1431478800, 1431482400, 1431486000, 
    1431489600, 1431493200, 1431496800, 1431500400, 1431504000, 1431507600, 
    1431511200, 1431514800, 1431518400, 1431522000, 1431525600, 1431529200, 
    1431532800, 1431536400, 1431540000, 1431543600, 1431547200, 1431550800, 
    1431554400, 1431558000, 1431561600, 1431565200, 1431568800, 1431572400, 
    1431576000, 1431579600, 1431583200, 1431586800, 1431590400, 1431594000, 
    1431597600, 1431601200, 1431604800, 1431608400, 1431612000, 1431615600, 
    1431619200, 1431622800, 1431626400, 1431630000, 1431633600, 1431637200, 
    1431640800, 1431644400, 1431648000, 1431651600, 1431655200, 1431658800, 
    1431662400, 1431666000, 1431669600, 1431673200, 1431676800, 1431680400, 
    1431684000, 1431687600, 1431691200, 1431694800, 1431698400, 1431702000, 
    1431705600, 1431709200, 1431712800, 1431716400, 1431720000, 1431723600, 
    1431727200, 1431730800, 1431734400, 1431738000, 1431741600, 1431745200, 
    1431748800, 1431752400, 1431756000, 1431759600, 1431763200, 1431766800, 
    1431770400, 1431774000, 1431777600, 1431781200, 1431784800, 1431788400, 
    1431792000, 1431795600, 1431799200, 1431802800, 1431806400, 1431813600, 
    1431817200, 1431820800, 1431824400, 1431828000, 1431831600, 1431835200, 
    1431838800, 1431842400, 1431846000, 1431849600, 1431853200, 1431856800, 
    1431860400, 1431864000, 1431867600, 1431871200, 1431874800, 1431878400, 
    1431882000, 1431885600, 1431889200, 1431892800, 1431896400, 1431900000, 
    1431903600, 1431907200, 1431910800, 1431914400, 1431918000, 1431921600, 
    1431925200, 1431928800, 1431932400, 1431936000, 1431939600, 1431943200, 
    1431946800, 1431950400, 1431954000, 1431957600, 1431961200, 1431964800, 
    1431968400, 1431972000, 1431975600, 1431979200, 1431982800, 1431986400, 
    1431990000, 1431993600, 1431997200, 1432000800, 1432004400, 1432008000, 
    1432011600, 1432015200, 1432018800, 1432022400, 1432026000, 1432029600, 
    1432033200, 1432036800, 1432040400, 1432044000, 1432047600, 1432051200, 
    1432058400, 1432062000, 1432065600, 1432069200, 1432072800, 1432076400, 
    1432080000, 1432083600, 1432087200, 1432090800, 1432094400, 1432098000, 
    1432101600, 1432105200, 1432108800, 1432112400, 1432116000, 1432119600, 
    1432123200, 1432126800, 1432130400, 1432134000, 1432137600, 1432141200, 
    1432144800, 1432148400, 1432152000, 1432155600, 1432159200, 1432162800, 
    1432166400, 1432170000, 1432173600, 1432177200, 1432180800, 1432184400, 
    1432188000, 1432191600, 1432195200, 1432198800, 1432202400, 1432206000, 
    1432209600, 1432213200, 1432216800, 1432220400, 1432224000, 1432227600, 
    1432231200, 1432234800, 1432238400, 1432242000, 1432245600, 1432249200, 
    1432252800, 1432256400, 1432260000, 1432263600, 1432267200, 1432270800, 
    1432274400, 1432278000, 1432281600, 1432285200, 1432288800, 1432292400, 
    1432296000, 1432299600, 1432303200, 1432306800, 1432310400, 1432314000, 
    1432317600, 1432321200, 1432324800, 1432328400, 1432332000, 1432335600, 
    1432339200, 1432342800, 1432346400, 1432350000, 1432357200, 1432360800, 
    1432364400, 1432368000, 1432371600, 1432375200, 1432378800, 1432382400, 
    1432386000, 1432389600, 1432393200, 1432396800, 1432400400, 1432404000, 
    1432407600, 1432411200, 1432414800, 1432418400, 1432422000, 1432425600, 
    1432429200, 1432432800, 1432436400, 1432458000, 1432461600, 1432465200, 
    1432468800, 1432472400, 1432476000, 1432483200, 1432486800, 1432490400, 
    1432494000, 1432497600, 1432501200, 1432504800, 1432508400, 1432512000, 
    1432515600, 1432519200, 1432526400, 1432530000, 1432537200, 1432544400, 
    1432551600, 1432555200, 1432558800, 1432562400, 1432566000, 1432573200, 
    1432576800, 1432580400, 1432584000, 1432587600, 1432591200, 1432594800, 
    1432598400, 1432605600, 1432616400, 1432620000, 1432623600, 1432627200, 
    1432630800, 1432634400, 1432638000, 1432641600, 1432645200, 1432648800, 
    1432652400, 1432656000, 1432659600, 1432663200, 1432666800, 1432670400, 
    1432674000, 1432677600, 1432681200, 1432684800, 1432688400, 1432692000, 
    1432695600, 1432699200, 1432702800, 1432706400, 1432710000, 1432713600, 
    1432717200, 1432720800, 1432724400, 1432728000, 1432731600, 1432735200, 
    1432738800, 1432742400, 1432746000, 1432749600, 1432753200, 1432756800, 
    1432760400, 1432764000, 1432767600, 1432771200, 1432774800, 1432778400, 
    1432782000, 1432785600, 1432789200, 1432792800, 1432796400, 1432800000, 
    1432803600, 1432807200, 1432810800, 1432814400, 1432818000, 1432821600, 
    1432825200, 1432828800, 1432832400, 1432836000, 1432839600, 1432843200, 
    1432846800, 1432850400, 1432854000, 1432857600, 1432861200, 1432864800, 
    1432868400, 1432872000, 1432875600, 1432879200, 1432882800, 1432886400, 
    1432890000, 1432893600, 1432897200, 1432900800, 1432904400, 1432908000, 
    1432911600, 1432915200, 1432918800, 1432922400, 1432926000, 1432929600, 
    1432933200, 1432936800, 1432940400, 1432944000, 1432947600, 1432951200, 
    1432954800, 1432958400, 1432962000, 1432965600, 1432969200, 1432972800, 
    1432976400, 1432980000, 1432983600, 1432987200, 1432990800, 1432994400, 
    1432998000, 1433001600, 1433005200, 1433008800, 1433012400, 1433016000, 
    1433019600, 1433023200, 1433026800, 1433030400, 1433034000, 1433037600, 
    1433041200, 1433044800, 1433048400, 1433052000, 1433055600, 1433059200, 
    1433062800, 1433066400, 1433070000, 1433073600, 1433077200, 1433080800, 
    1433084400, 1433088000, 1433091600, 1433095200, 1433098800, 1433102400, 
    1433106000, 1433109600, 1433113200, 1433116800, 1433120400, 1433124000, 
    1433127600, 1433131200, 1433134800, 1433138400, 1433142000, 1433145600, 
    1433149200, 1433152800, 1433156400, 1433160000, 1433163600, 1433167200, 
    1433170800, 1433174400, 1433178000, 1433181600, 1433185200, 1433188800, 
    1433192400, 1433196000, 1433199600, 1433203200, 1433206800, 1433210400, 
    1433214000, 1433217600, 1433221200, 1433224800, 1433228400, 1433232000, 
    1433235600, 1433239200, 1433242800, 1433246400, 1433250000, 1433253600, 
    1433257200, 1433260800, 1433264400, 1433268000, 1433271600, 1433275200, 
    1433278800, 1433282400, 1433286000, 1433289600, 1433293200, 1433296800, 
    1433300400, 1433304000, 1433307600, 1433311200, 1433314800, 1433318400, 
    1433322000, 1433325600, 1433329200, 1433332800, 1433336400, 1433340000, 
    1433343600, 1433347200, 1433350800, 1433354400, 1433358000, 1433361600, 
    1433365200, 1433368800, 1433372400, 1433376000, 1433379600, 1433383200, 
    1433386800, 1433390400, 1433394000, 1433397600, 1433401200, 1433404800, 
    1433408400, 1433412000, 1433415600, 1433419200, 1433422800, 1433426400, 
    1433430000, 1433433600, 1433437200, 1433440800, 1433444400, 1433448000, 
    1433451600, 1433455200, 1433458800, 1433462400, 1433466000, 1433469600, 
    1433473200, 1433476800, 1433480400, 1433484000, 1433487600, 1433491200, 
    1433494800, 1433498400, 1433502000, 1433505600, 1433509200, 1433512800, 
    1433516400, 1433520000, 1433523600, 1433527200, 1433530800, 1433534400, 
    1433538000, 1433541600, 1433545200, 1433548800, 1433552400, 1433556000, 
    1433559600, 1433563200, 1433566800, 1433570400, 1433574000, 1433577600, 
    1433581200, 1433584800, 1433588400, 1433592000, 1433595600, 1433599200, 
    1433602800, 1433606400, 1433610000, 1433613600, 1433617200, 1433620800, 
    1433624400, 1433628000, 1433631600, 1433635200, 1433638800, 1433642400, 
    1433646000, 1433649600, 1433653200, 1433656800, 1433660400, 1433664000, 
    1433667600, 1433671200, 1433674800, 1433678400, 1433682000, 1433685600, 
    1433689200, 1433692800, 1433696400, 1433700000, 1433703600, 1433707200, 
    1433710800, 1433714400, 1433718000, 1433721600, 1433725200, 1433728800, 
    1433732400, 1433736000, 1433739600, 1433743200, 1433746800, 1433750400, 
    1433754000, 1433757600, 1433761200, 1433764800, 1433768400, 1433772000, 
    1433775600, 1433779200, 1433782800, 1433786400, 1433790000, 1433793600, 
    1433797200, 1433800800, 1433804400, 1433808000, 1433811600, 1433815200, 
    1433818800, 1433822400, 1433826000, 1433829600, 1433833200, 1433836800, 
    1433840400, 1433844000, 1433847600, 1433851200, 1433854800, 1433858400, 
    1433862000, 1433865600, 1433869200, 1433872800, 1433876400, 1433880000, 
    1433883600, 1433887200, 1433890800, 1433894400, 1433898000, 1433901600, 
    1433905200, 1433908800, 1433912400, 1433916000, 1433919600, 1433923200, 
    1433926800, 1433930400, 1433934000, 1433937600, 1433941200, 1433944800, 
    1433948400, 1433952000, 1433955600, 1433959200, 1433962800, 1433966400, 
    1433970000, 1433973600, 1433977200, 1433980800, 1433984400, 1433988000, 
    1433991600, 1433995200, 1433998800, 1434002400, 1434006000, 1434009600, 
    1434013200, 1434016800, 1434020400, 1434024000, 1434027600, 1434031200, 
    1434034800, 1434038400, 1434042000, 1434045600, 1434049200, 1434052800, 
    1434056400, 1434060000, 1434063600, 1434067200, 1434070800, 1434074400, 
    1434078000, 1434081600, 1434085200, 1434088800, 1434092400, 1434096000, 
    1434099600, 1434103200, 1434106800, 1434110400, 1434114000, 1434117600, 
    1434121200, 1434124800, 1434128400, 1434132000, 1434135600, 1434139200, 
    1434142800, 1434146400, 1434150000, 1434153600, 1434157200, 1434160800, 
    1434164400, 1434168000, 1434171600, 1434175200, 1434178800, 1434182400, 
    1434186000, 1434189600, 1434193200, 1434196800, 1434200400, 1434204000, 
    1434207600, 1434211200, 1434214800, 1434218400, 1434222000, 1434225600, 
    1434229200, 1434232800, 1434236400, 1434240000, 1434243600, 1434247200, 
    1434250800, 1434254400, 1434258000, 1434261600, 1434265200, 1434268800, 
    1434272400, 1434276000, 1434279600, 1434283200, 1434286800, 1434290400, 
    1434294000, 1434297600, 1434301200, 1434304800, 1434308400, 1434312000, 
    1434315600, 1434319200, 1434322800, 1434326400, 1434330000, 1434333600, 
    1434337200, 1434340800, 1434344400, 1434348000, 1434351600, 1434355200, 
    1434358800, 1434362400, 1434366000, 1434369600, 1434373200, 1434376800, 
    1434380400, 1434384000, 1434387600, 1434391200, 1434394800, 1434398400, 
    1434402000, 1434405600, 1434409200, 1434412800, 1434416400, 1434420000, 
    1434423600, 1434427200, 1434430800, 1434434400, 1434438000, 1434441600, 
    1434445200, 1434448800, 1434452400, 1434456000, 1434459600, 1434463200, 
    1434466800, 1434470400, 1434474000, 1434477600, 1434481200, 1434484800, 
    1434488400, 1434492000, 1434495600, 1434499200, 1434502800, 1434506400, 
    1434510000, 1434513600, 1434517200, 1434520800, 1434524400, 1434528000, 
    1434531600, 1434535200, 1434538800, 1434542400, 1434546000, 1434549600, 
    1434553200, 1434556800, 1434560400, 1434564000, 1434567600, 1434571200, 
    1434574800, 1434578400, 1434582000, 1434585600, 1434589200, 1434592800, 
    1434596400, 1434600000, 1434603600, 1434607200, 1434610800, 1434614400, 
    1434618000, 1434621600, 1434625200, 1434628800, 1434632400, 1434636000, 
    1434639600, 1434643200, 1434646800, 1434650400, 1434654000, 1434657600, 
    1434661200, 1434664800, 1434668400, 1434672000, 1434675600, 1434679200, 
    1434682800, 1434686400, 1434690000, 1434693600, 1434697200, 1434700800, 
    1434704400, 1434708000, 1434711600, 1434715200, 1434718800, 1434722400, 
    1434726000, 1434729600, 1434733200, 1434736800, 1434740400, 1434744000, 
    1434747600, 1434751200, 1434754800, 1434758400, 1434762000, 1434765600, 
    1434769200, 1434772800, 1434776400, 1434780000, 1434783600, 1434787200, 
    1434790800, 1434794400, 1434798000, 1434801600, 1434805200, 1434808800, 
    1434812400, 1434816000, 1434819600, 1434823200, 1434826800, 1434830400, 
    1434834000, 1434837600, 1434841200, 1434844800, 1434848400, 1434852000, 
    1434855600, 1434859200, 1434862800, 1434866400, 1434870000, 1434873600, 
    1434877200, 1434880800, 1434884400, 1434888000, 1434891600, 1434895200, 
    1434898800, 1434902400, 1434906000, 1434909600, 1434913200, 1434916800, 
    1434920400, 1434924000, 1434927600, 1434931200, 1434934800, 1434938400, 
    1434942000, 1434945600, 1434949200, 1434952800, 1434956400, 1434960000, 
    1434963600, 1434967200, 1434970800, 1434974400, 1434978000, 1434981600, 
    1434985200, 1434988800, 1434992400, 1434996000, 1434999600, 1435003200, 
    1435006800, 1435010400, 1435014000, 1435017600, 1435021200, 1435024800, 
    1435028400, 1435032000, 1435035600, 1435039200, 1435042800, 1435046400, 
    1435050000, 1435053600, 1435057200, 1435060800, 1435064400, 1435068000, 
    1435071600, 1435075200, 1435078800, 1435082400, 1435086000, 1435089600, 
    1435093200, 1435096800, 1435100400, 1435104000, 1435107600, 1435111200, 
    1435114800, 1435118400, 1435122000, 1435125600, 1435129200, 1435132800, 
    1435136400, 1435140000, 1435143600, 1435147200, 1435150800, 1435154400, 
    1435158000, 1435161600, 1435165200, 1435168800, 1435172400, 1435176000, 
    1435179600, 1435183200, 1435186800, 1435190400, 1435194000, 1435197600, 
    1435201200, 1435204800, 1435208400, 1435212000, 1435215600, 1435219200, 
    1435222800, 1435226400, 1435230000, 1435233600, 1435237200, 1435240800, 
    1435244400, 1435248000, 1435251600, 1435255200, 1435258800, 1435262400, 
    1435266000, 1435269600, 1435273200, 1435276800, 1435280400, 1435284000, 
    1435287600, 1435291200, 1435294800, 1435298400, 1435302000, 1435305600, 
    1435309200, 1435312800, 1435316400, 1435320000, 1435323600, 1435327200, 
    1435330800, 1435334400, 1435338000, 1435341600, 1435345200, 1435348800, 
    1435352400, 1435356000, 1435359600, 1435363200, 1435366800, 1435370400, 
    1435374000, 1435377600, 1435381200, 1435384800, 1435388400, 1435392000, 
    1435395600, 1435399200, 1435402800, 1435406400, 1435410000, 1435413600, 
    1435417200, 1435420800, 1435424400, 1435428000, 1435431600, 1435435200, 
    1435438800, 1435442400, 1435446000, 1435449600, 1435453200, 1435456800, 
    1435460400, 1435464000, 1435467600, 1435471200, 1435474800, 1435478400, 
    1435482000, 1435485600, 1435489200, 1435492800, 1435496400, 1435500000, 
    1435503600, 1435507200, 1435510800, 1435514400, 1435518000, 1435521600, 
    1435525200, 1435528800, 1435532400, 1435536000, 1435539600, 1435543200, 
    1435546800, 1435550400, 1435554000, 1435557600, 1435561200, 1435564800, 
    1435568400, 1435572000, 1435575600, 1435579200, 1435582800, 1435586400, 
    1435590000, 1435593600, 1435597200, 1435600800, 1435604400, 1435608000, 
    1435611600, 1435615200, 1435618800, 1435622400, 1435626000, 1435629600, 
    1435633200, 1435636800, 1435640400, 1435644000, 1435647600, 1435651200, 
    1435654800, 1435658400, 1435662000, 1435665600, 1435669200, 1435672800, 
    1435676400, 1435680000, 1435683600, 1435687200, 1435690800, 1435694400, 
    1435698000, 1435701600, 1435705200, 1435708800, 1435712400, 1435716000, 
    1435719600, 1435723200, 1435726800, 1435730400, 1435734000, 1435737600, 
    1435741200, 1435744800, 1435748400, 1435752000, 1435755600, 1435759200, 
    1435762800, 1435766400, 1435770000, 1435773600, 1435777200, 1435780800, 
    1435784400, 1435788000, 1435791600, 1435795200, 1435798800, 1435802400, 
    1435806000, 1435809600, 1435813200, 1435816800, 1435820400, 1435824000, 
    1435827600, 1435831200, 1435834800, 1435838400, 1435842000, 1435845600, 
    1435849200, 1435852800, 1435856400, 1435860000, 1435863600, 1435867200, 
    1435870800, 1435874400, 1435878000, 1435881600, 1435885200, 1435888800, 
    1435892400, 1435896000, 1435899600, 1435903200, 1435906800, 1435910400, 
    1435914000, 1435917600, 1435921200, 1435924800, 1435928400, 1435932000, 
    1435935600, 1435939200, 1435942800, 1435946400, 1435950000, 1435953600, 
    1435957200, 1435960800, 1435964400, 1435968000, 1435971600, 1435975200, 
    1435978800, 1435982400, 1435986000, 1435989600, 1435993200, 1435996800, 
    1436000400, 1436004000, 1436007600, 1436011200, 1436014800, 1436018400, 
    1436022000, 1436025600, 1436029200, 1436032800, 1436036400, 1436040000, 
    1436043600, 1436047200, 1436050800, 1436054400, 1436058000, 1436061600, 
    1436065200, 1436068800, 1436072400, 1436076000, 1436079600, 1436083200, 
    1436086800, 1436090400, 1436094000, 1436097600, 1436101200, 1436104800, 
    1436108400, 1436112000, 1436115600, 1436119200, 1436122800, 1436126400, 
    1436130000, 1436133600, 1436137200, 1436140800, 1436144400, 1436148000, 
    1436151600, 1436155200, 1436158800, 1436162400, 1436166000, 1436169600, 
    1436173200, 1436176800, 1436180400, 1436184000, 1436187600, 1436191200, 
    1436194800, 1436198400, 1436202000, 1436205600, 1436209200, 1436212800, 
    1436216400, 1436220000, 1436223600, 1436227200, 1436230800, 1436234400, 
    1436238000, 1436241600, 1436245200, 1436248800, 1436252400, 1436256000, 
    1436259600, 1436263200, 1436266800, 1436270400, 1436274000, 1436277600, 
    1436281200, 1436284800, 1436288400, 1436292000, 1436295600, 1436299200, 
    1436302800, 1436306400, 1436310000, 1436313600, 1436317200, 1436320800, 
    1436324400, 1436328000, 1436331600, 1436335200, 1436338800, 1436342400, 
    1436346000, 1436349600, 1436353200, 1436356800, 1436360400, 1436364000, 
    1436367600, 1436371200, 1436374800, 1436378400, 1436382000, 1436385600, 
    1436389200, 1436392800, 1436396400, 1436400000, 1436403600, 1436407200, 
    1436410800, 1436414400, 1436418000, 1436421600, 1436425200, 1436428800, 
    1436432400, 1436436000, 1436439600, 1436443200, 1436446800, 1436450400, 
    1436454000, 1436457600, 1436461200, 1436464800, 1436468400, 1436472000, 
    1436475600, 1436479200, 1436482800, 1436486400, 1436490000, 1436493600, 
    1436497200, 1436500800, 1436504400, 1436508000, 1436511600, 1436515200, 
    1436518800, 1436522400, 1436526000, 1436529600, 1436533200, 1436536800, 
    1436540400, 1436544000, 1436547600, 1436551200, 1436554800, 1436558400, 
    1436562000, 1436565600, 1436569200, 1436572800, 1436576400, 1436580000, 
    1436583600, 1436587200, 1436590800, 1436594400, 1436598000, 1436601600, 
    1436605200, 1436608800, 1436612400, 1436616000, 1436619600, 1436623200, 
    1436626800, 1436630400, 1436634000, 1436637600, 1436641200, 1436644800, 
    1436648400, 1436652000, 1436655600, 1436659200, 1436662800, 1436666400, 
    1436670000, 1436673600, 1436677200, 1436680800, 1436684400, 1436688000, 
    1436691600, 1436695200, 1436698800, 1436702400, 1436706000, 1436709600, 
    1436713200, 1436716800, 1436720400, 1436724000, 1436727600, 1436731200, 
    1436734800, 1436738400, 1436742000, 1436745600, 1436749200, 1436752800, 
    1436756400, 1436760000, 1436763600, 1436767200, 1436770800, 1436774400, 
    1436778000, 1436781600, 1436785200, 1436788800, 1436792400, 1436796000, 
    1436799600, 1436803200, 1436806800, 1436810400, 1436814000, 1436817600, 
    1436821200, 1436824800, 1436828400, 1436832000, 1436835600, 1436839200, 
    1436842800, 1436846400, 1436850000, 1436853600, 1436857200, 1436860800, 
    1436864400, 1436868000, 1436871600, 1436875200, 1436878800, 1436882400, 
    1436886000, 1436889600, 1436893200, 1436896800, 1436900400, 1436904000, 
    1436907600, 1436911200, 1436914800, 1436918400, 1436922000, 1436925600, 
    1436929200, 1436932800, 1436936400, 1436940000, 1436943600, 1436947200, 
    1436950800, 1436954400, 1436958000, 1436961600, 1436965200, 1436968800, 
    1436972400, 1436976000, 1436979600, 1436983200, 1436986800, 1436990400, 
    1436994000, 1436997600, 1437001200, 1437004800, 1437008400, 1437012000, 
    1437015600, 1437019200, 1437022800, 1437026400, 1437030000, 1437033600, 
    1437037200, 1437040800, 1437044400, 1437048000, 1437051600, 1437055200, 
    1437058800, 1437062400, 1437066000, 1437069600, 1437073200, 1437076800, 
    1437080400, 1437084000, 1437087600, 1437091200, 1437094800, 1437098400, 
    1437102000, 1437105600, 1437109200, 1437112800, 1437116400, 1437120000, 
    1437123600, 1437127200, 1437130800, 1437134400, 1437138000, 1437141600, 
    1437145200, 1437148800, 1437152400, 1437156000, 1437159600, 1437163200, 
    1437166800, 1437170400, 1437174000, 1437177600, 1437181200, 1437184800, 
    1437188400, 1437192000, 1437195600, 1437199200, 1437202800, 1437206400, 
    1437210000, 1437213600, 1437217200, 1437220800, 1437224400, 1437228000, 
    1437231600, 1437235200, 1437238800, 1437242400, 1437246000, 1437249600, 
    1437253200, 1437256800, 1437260400, 1437264000, 1437267600, 1437271200, 
    1437274800, 1437278400, 1437282000, 1437285600, 1437289200, 1437292800, 
    1437296400, 1437300000, 1437303600, 1437307200, 1437310800, 1437314400, 
    1437318000, 1437321600, 1437325200, 1437328800, 1437332400, 1437336000, 
    1437339600, 1437343200, 1437346800, 1437350400, 1437354000, 1437357600, 
    1437361200, 1437364800, 1437368400, 1437372000, 1437375600, 1437379200, 
    1437382800, 1437386400, 1437390000, 1437393600, 1437397200, 1437400800, 
    1437404400, 1437408000, 1437411600, 1437415200, 1437418800, 1437422400, 
    1437426000, 1437429600, 1437433200, 1437436800, 1437440400, 1437444000, 
    1437447600, 1437451200, 1437454800, 1437458400, 1437462000, 1437465600, 
    1437469200, 1437472800, 1437476400, 1437480000, 1437483600, 1437487200, 
    1437490800, 1437494400, 1437498000, 1437501600, 1437505200, 1437508800, 
    1437512400, 1437516000, 1437519600, 1437523200, 1437526800, 1437530400, 
    1437534000, 1437537600, 1437541200, 1437544800, 1437548400, 1437552000, 
    1437555600, 1437559200, 1437562800, 1437566400, 1437570000, 1437573600, 
    1437577200, 1437580800, 1437584400, 1437588000, 1437591600, 1437595200, 
    1437598800, 1437602400, 1437606000, 1437609600, 1437613200, 1437616800, 
    1437620400, 1437624000, 1437627600, 1437631200, 1437634800, 1437638400, 
    1437642000, 1437645600, 1437649200, 1437652800, 1437656400, 1437660000, 
    1437663600, 1437667200, 1437670800, 1437674400, 1437678000, 1437681600, 
    1437685200, 1437688800, 1437692400, 1437696000, 1437699600, 1437703200, 
    1437706800, 1437710400, 1437714000, 1437717600, 1437721200, 1437724800, 
    1437728400, 1437732000, 1437735600, 1437739200, 1437742800, 1437746400, 
    1437750000, 1437753600, 1437757200, 1437760800, 1437764400, 1437768000, 
    1437771600, 1437775200, 1437778800, 1437782400, 1437786000, 1437789600, 
    1437793200, 1437796800, 1437800400, 1437804000, 1437807600, 1437811200, 
    1437814800, 1437818400, 1437822000, 1437825600, 1437829200, 1437832800, 
    1437836400, 1437840000, 1437843600, 1437847200, 1437850800, 1437854400, 
    1437858000, 1437861600, 1437865200, 1437868800, 1437872400, 1437876000, 
    1437879600, 1437883200, 1437886800, 1437890400, 1437894000, 1437897600, 
    1437901200, 1437904800, 1437908400, 1437912000, 1437915600, 1437919200, 
    1437922800, 1437926400, 1437930000, 1437933600, 1437937200, 1437940800, 
    1437944400, 1437948000, 1437951600, 1437955200, 1437958800, 1437962400, 
    1437966000, 1437969600, 1437973200, 1437976800, 1437980400, 1437984000, 
    1437987600, 1437991200, 1437994800, 1437998400, 1438002000, 1438005600, 
    1438009200, 1438012800, 1438016400, 1438020000, 1438023600, 1438027200, 
    1438030800, 1438034400, 1438038000, 1438041600, 1438045200, 1438048800, 
    1438052400, 1438056000, 1438059600, 1438063200, 1438066800, 1438070400, 
    1438074000, 1438077600, 1438081200, 1438084800, 1438088400, 1438092000, 
    1438095600, 1438099200, 1438102800, 1438106400, 1438110000, 1438113600, 
    1438117200, 1438120800, 1438124400, 1438128000, 1438131600, 1438135200, 
    1438138800, 1438142400, 1438146000, 1438149600, 1438153200, 1438156800, 
    1438160400, 1438164000, 1438167600, 1438171200, 1438174800, 1438178400, 
    1438182000, 1438185600, 1438189200, 1438192800, 1438196400, 1438200000, 
    1438203600, 1438207200, 1438210800, 1438214400, 1438218000, 1438221600, 
    1438225200, 1438228800, 1438232400, 1438236000, 1438239600, 1438243200, 
    1438246800, 1438250400, 1438254000, 1438257600, 1438261200, 1438264800, 
    1438268400, 1438272000, 1438275600, 1438279200, 1438282800, 1438286400, 
    1438290000, 1438293600, 1438297200, 1438300800, 1438304400, 1438308000, 
    1438311600, 1438315200, 1438318800, 1438322400, 1438326000, 1438329600, 
    1438333200, 1438336800, 1438340400, 1438344000, 1438347600, 1438351200, 
    1438354800, 1438358400, 1438362000, 1438365600, 1438369200, 1438372800, 
    1438376400, 1438380000, 1438383600, 1438387200, 1438390800, 1438394400, 
    1438398000, 1438401600, 1438405200, 1438408800, 1438412400, 1438416000, 
    1438419600, 1438423200, 1438426800, 1438430400, 1438434000, 1438437600, 
    1438441200, 1438444800, 1438448400, 1438452000, 1438455600, 1438459200, 
    1438462800, 1438466400, 1438470000, 1438473600, 1438477200, 1438480800, 
    1438484400, 1438488000, 1438491600, 1438495200, 1438498800, 1438502400, 
    1438506000, 1438509600, 1438513200, 1438516800, 1438520400, 1438524000, 
    1438527600, 1438531200, 1438534800, 1438538400, 1438542000, 1438545600, 
    1438549200, 1438552800, 1438556400, 1438560000, 1438563600, 1438567200, 
    1438570800, 1438574400, 1438578000, 1438581600, 1438585200, 1438588800, 
    1438592400, 1438596000, 1438599600, 1438603200, 1438606800, 1438610400, 
    1438614000, 1438617600, 1438621200, 1438624800, 1438628400, 1438632000, 
    1438635600, 1438639200, 1438642800, 1438646400, 1438650000, 1438653600, 
    1438657200, 1438660800, 1438664400, 1438668000, 1438671600, 1438675200, 
    1438678800, 1438682400, 1438686000, 1438689600, 1438693200, 1438696800, 
    1438700400, 1438704000, 1438707600, 1438711200, 1438714800, 1438718400, 
    1438722000, 1438725600, 1438729200, 1438732800, 1438736400, 1438740000, 
    1438743600, 1438747200, 1438750800, 1438754400, 1438758000, 1438761600, 
    1438765200, 1438768800, 1438772400, 1438776000, 1438779600, 1438783200, 
    1438786800, 1438790400, 1438794000, 1438797600, 1438801200, 1438804800, 
    1438808400, 1438812000, 1438815600, 1438819200, 1438822800, 1438826400, 
    1438830000, 1438833600, 1438837200, 1438840800, 1438844400, 1438848000, 
    1438851600, 1438855200, 1438858800, 1438862400, 1438866000, 1438869600, 
    1438873200, 1438876800, 1438880400, 1438884000, 1438887600, 1438891200, 
    1438894800, 1438898400, 1438902000, 1438905600, 1438909200, 1438912800, 
    1438916400, 1438920000, 1438923600, 1438927200, 1438930800, 1438934400, 
    1438938000, 1438941600, 1438945200, 1438948800, 1438952400, 1438956000, 
    1438959600, 1438963200, 1438966800, 1438970400, 1438974000, 1438977600, 
    1438981200, 1438984800, 1438988400, 1438992000, 1438995600, 1438999200, 
    1439002800, 1439006400, 1439010000, 1439013600, 1439017200, 1439020800, 
    1439024400, 1439028000, 1439031600, 1439035200, 1439038800, 1439042400, 
    1439046000, 1439049600, 1439053200, 1439056800, 1439060400, 1439064000, 
    1439067600, 1439071200, 1439074800, 1439078400, 1439082000, 1439085600, 
    1439089200, 1439092800, 1439096400, 1439100000, 1439103600, 1439107200, 
    1439110800, 1439114400, 1439118000, 1439121600, 1439125200, 1439128800, 
    1439132400, 1439136000, 1439139600, 1439143200, 1439146800, 1439150400, 
    1439154000, 1439157600, 1439161200, 1439164800, 1439168400, 1439172000, 
    1439175600, 1439179200, 1439182800, 1439186400, 1439190000, 1439193600, 
    1439197200, 1439200800, 1439204400, 1439208000, 1439211600, 1439215200, 
    1439218800, 1439222400, 1439226000, 1439229600, 1439233200, 1439236800, 
    1439240400, 1439244000, 1439247600, 1439251200, 1439254800, 1439258400, 
    1439262000, 1439265600, 1439269200, 1439272800, 1439276400, 1439280000, 
    1439283600, 1439287200, 1439290800, 1439294400, 1439298000, 1439301600, 
    1439305200, 1439308800, 1439312400, 1439316000, 1439319600, 1439323200, 
    1439326800, 1439330400, 1439334000, 1439337600, 1439341200, 1439344800, 
    1439348400, 1439352000, 1439355600, 1439359200, 1439362800, 1439366400, 
    1439370000, 1439373600, 1439377200, 1439380800, 1439384400, 1439388000, 
    1439391600, 1439395200, 1439398800, 1439402400, 1439406000, 1439409600, 
    1439413200, 1439416800, 1439420400, 1439424000, 1439427600, 1439431200, 
    1439434800, 1439438400, 1439442000, 1439445600, 1439449200, 1439452800, 
    1439456400, 1439460000, 1439463600, 1439467200, 1439470800, 1439474400, 
    1439478000, 1439481600, 1439485200, 1439488800, 1439492400, 1439496000, 
    1439499600, 1439503200, 1439506800, 1439510400, 1439514000, 1439517600, 
    1439521200, 1439524800, 1439528400, 1439532000, 1439535600, 1439539200, 
    1439542800, 1439546400, 1439550000, 1439553600, 1439557200, 1439560800, 
    1439564400, 1439568000, 1439571600, 1439575200, 1439578800, 1439582400, 
    1439586000, 1439589600, 1439593200, 1439596800, 1439600400, 1439604000, 
    1439607600, 1439611200, 1439614800, 1439618400, 1439622000, 1439625600, 
    1439629200, 1439632800, 1439636400, 1439640000, 1439643600, 1439647200, 
    1439650800, 1439654400, 1439658000, 1439661600, 1439665200, 1439668800, 
    1439672400, 1439676000, 1439679600, 1439683200, 1439686800, 1439690400, 
    1439694000, 1439697600, 1439701200, 1439704800, 1439708400, 1439712000, 
    1439715600, 1439719200, 1439722800, 1439726400, 1439730000, 1439733600, 
    1439737200, 1439740800, 1439744400, 1439748000, 1439751600, 1439755200, 
    1439758800, 1439762400, 1439766000, 1439769600, 1439773200, 1439776800, 
    1439780400, 1439784000, 1439787600, 1439791200, 1439794800, 1439798400, 
    1439802000, 1439805600, 1439809200, 1439812800, 1439816400, 1439820000, 
    1439823600, 1439827200, 1439830800, 1439834400, 1439838000, 1439841600, 
    1439845200, 1439848800, 1439852400, 1439856000, 1439859600, 1439863200, 
    1439866800, 1439870400, 1439874000, 1439877600, 1439881200, 1439884800, 
    1439888400, 1439892000, 1439895600, 1439899200, 1439902800, 1439906400, 
    1439910000, 1439913600, 1439917200, 1439920800, 1439924400, 1439928000, 
    1439931600, 1439935200, 1439938800, 1439942400, 1439946000, 1439949600, 
    1439953200, 1439956800, 1439960400, 1439964000, 1439967600, 1439971200, 
    1439974800, 1439978400, 1439982000, 1439985600, 1439989200, 1439992800, 
    1439996400, 1440000000, 1440003600, 1440007200, 1440010800, 1440014400, 
    1440018000, 1440021600, 1440025200, 1440028800, 1440032400, 1440036000, 
    1440039600, 1440043200, 1440046800, 1440050400, 1440054000, 1440057600, 
    1440061200, 1440064800, 1440068400, 1440072000, 1440075600, 1440079200, 
    1440082800, 1440086400, 1440090000, 1440093600, 1440097200, 1440100800, 
    1440104400, 1440108000, 1440111600, 1440115200, 1440118800, 1440122400, 
    1440126000, 1440129600, 1440133200, 1440136800, 1440140400, 1440144000, 
    1440147600, 1440151200, 1440154800, 1440158400, 1440162000, 1440165600, 
    1440169200, 1440172800, 1440176400, 1440180000, 1440183600, 1440187200, 
    1440190800, 1440194400, 1440198000, 1440201600, 1440205200, 1440208800, 
    1440212400, 1440216000, 1440219600, 1440223200, 1440226800, 1440230400, 
    1440234000, 1440237600, 1440241200, 1440244800, 1440248400, 1440252000, 
    1440255600, 1440259200, 1440262800, 1440266400, 1440270000, 1440273600, 
    1440277200, 1440280800, 1440284400, 1440288000, 1440291600, 1440295200, 
    1440298800, 1440302400, 1440306000, 1440309600, 1440313200, 1440316800, 
    1440320400, 1440324000, 1440327600, 1440331200, 1440334800, 1440338400, 
    1440342000, 1440345600, 1440349200, 1440352800, 1440356400, 1440360000, 
    1440363600, 1440367200, 1440370800, 1440374400, 1440378000, 1440381600, 
    1440385200, 1440388800, 1440392400, 1440396000, 1440399600, 1440403200, 
    1440406800, 1440410400, 1440414000, 1440417600, 1440421200, 1440424800, 
    1440428400, 1440432000, 1440435600, 1440439200, 1440442800, 1440446400, 
    1440450000, 1440453600, 1440457200, 1440460800, 1440464400, 1440468000, 
    1440471600, 1440475200, 1440478800, 1440482400, 1440486000, 1440489600, 
    1440493200, 1440496800, 1440500400, 1440504000, 1440507600, 1440511200, 
    1440514800, 1440518400, 1440522000, 1440525600, 1440529200, 1440532800, 
    1440536400, 1440540000, 1440543600, 1440547200, 1440550800, 1440554400, 
    1440558000, 1440561600, 1440565200, 1440568800, 1440572400, 1440576000, 
    1440579600, 1440583200, 1440586800, 1440590400, 1440594000, 1440597600, 
    1440601200, 1440604800, 1440608400, 1440612000, 1440615600, 1440619200, 
    1440622800, 1440626400, 1440630000, 1440633600, 1440637200, 1440640800, 
    1440644400, 1440648000, 1440651600, 1440655200, 1440658800, 1440662400, 
    1440666000, 1440669600, 1440673200, 1440676800, 1440680400, 1440684000, 
    1440687600, 1440691200, 1440694800, 1440698400, 1440702000, 1440705600, 
    1440709200, 1440712800, 1440716400, 1440720000, 1440723600, 1440727200, 
    1440730800, 1440734400, 1440738000, 1440741600, 1440745200, 1440748800, 
    1440752400, 1440756000, 1440759600, 1440763200, 1440766800, 1440770400, 
    1440774000, 1440777600, 1440781200, 1440784800, 1440788400, 1440792000, 
    1440795600, 1440799200, 1440802800, 1440806400, 1440810000, 1440813600, 
    1440817200, 1440820800, 1440824400, 1440828000, 1440831600, 1440835200, 
    1440838800, 1440842400, 1440846000, 1440849600, 1440853200, 1440856800, 
    1440860400, 1440864000, 1440867600, 1440871200, 1440874800, 1440878400, 
    1440882000, 1440885600, 1440889200, 1440892800, 1440896400, 1440900000, 
    1440903600, 1440907200, 1440910800, 1440914400, 1440918000, 1440921600, 
    1440925200, 1440928800, 1440932400, 1440936000, 1440939600, 1440943200, 
    1440946800, 1440950400, 1440954000, 1440957600, 1440961200, 1440964800, 
    1440968400, 1440972000, 1440975600, 1440979200, 1440982800, 1440986400, 
    1440990000, 1440993600, 1440997200, 1441000800, 1441004400, 1441008000, 
    1441011600, 1441015200, 1441018800, 1441022400, 1441026000, 1441029600, 
    1441033200, 1441036800, 1441040400, 1441044000, 1441047600, 1441051200, 
    1441054800, 1441058400, 1441062000, 1441065600, 1441069200, 1441072800, 
    1441076400, 1441080000, 1441083600, 1441087200, 1441090800, 1441094400, 
    1441098000, 1441101600, 1441105200, 1441108800, 1441112400, 1441116000, 
    1441119600, 1441123200, 1441126800, 1441130400, 1441134000, 1441137600, 
    1441141200, 1441144800, 1441148400, 1441152000, 1441155600, 1441159200, 
    1441162800, 1441166400, 1441170000, 1441173600, 1441177200, 1441180800, 
    1441184400, 1441188000, 1441191600, 1441195200, 1441198800, 1441202400, 
    1441206000, 1441209600, 1441213200, 1441216800, 1441220400, 1441224000, 
    1441227600, 1441231200, 1441234800, 1441238400, 1441242000, 1441245600, 
    1441249200, 1441252800, 1441256400, 1441260000, 1441263600, 1441267200, 
    1441270800, 1441274400, 1441278000, 1441281600, 1441285200, 1441288800, 
    1441292400, 1441296000, 1441299600, 1441303200, 1441306800, 1441310400, 
    1441314000, 1441317600, 1441321200, 1441324800, 1441328400, 1441332000, 
    1441335600, 1441339200, 1441342800, 1441346400, 1441350000, 1441353600, 
    1441357200, 1441360800, 1441364400, 1441368000, 1441371600, 1441375200, 
    1441378800, 1441382400, 1441386000, 1441389600, 1441393200, 1441396800, 
    1441400400, 1441404000, 1441407600, 1441411200, 1441414800, 1441418400, 
    1441422000, 1441425600, 1441429200, 1441432800, 1441436400, 1441440000, 
    1441443600, 1441447200, 1441450800, 1441454400, 1441458000, 1441461600, 
    1441465200, 1441468800, 1441472400, 1441476000, 1441479600, 1441483200, 
    1441486800, 1441490400, 1441494000, 1441497600, 1441501200, 1441504800, 
    1441508400, 1441512000, 1441515600, 1441519200, 1441522800, 1441526400, 
    1441530000, 1441533600, 1441537200, 1441540800, 1441544400, 1441548000, 
    1441551600, 1441555200, 1441558800, 1441562400, 1441566000, 1441569600, 
    1441573200, 1441576800, 1441580400, 1441584000, 1441587600, 1441591200, 
    1441594800, 1441598400, 1441602000, 1441605600, 1441609200, 1441612800, 
    1441616400, 1441620000, 1441623600, 1441627200, 1441630800, 1441634400, 
    1441638000, 1441641600, 1441645200, 1441648800, 1441652400, 1441656000, 
    1441659600, 1441663200, 1441666800, 1441670400, 1441674000, 1441677600, 
    1441681200, 1441684800, 1441688400, 1441692000, 1441695600, 1441699200, 
    1441702800, 1441706400, 1441710000, 1441713600, 1441717200, 1441720800, 
    1441724400, 1441728000, 1441731600, 1441735200, 1441738800, 1441742400, 
    1441746000, 1441749600, 1441753200, 1441756800, 1441760400, 1441764000, 
    1441767600, 1441771200, 1441774800, 1441778400, 1441782000, 1441785600, 
    1441789200, 1441792800, 1441796400, 1441800000, 1441803600, 1441807200, 
    1441810800, 1441814400, 1441818000, 1441821600, 1441825200, 1441828800, 
    1441832400, 1441836000, 1441839600, 1441843200, 1441846800, 1441850400, 
    1441854000, 1441857600, 1441861200, 1441864800, 1441868400, 1441872000, 
    1441875600, 1441879200, 1441882800, 1441886400, 1441890000, 1441893600, 
    1441897200, 1441900800, 1441904400, 1441908000, 1441911600, 1441915200, 
    1441918800, 1441922400, 1441926000, 1441929600, 1441933200, 1441936800, 
    1441940400, 1441944000, 1441947600, 1441951200, 1441954800, 1441958400, 
    1441962000, 1441965600, 1441969200, 1441972800, 1441976400, 1441980000, 
    1441983600, 1441987200, 1441990800, 1441994400, 1441998000, 1442001600, 
    1442005200, 1442008800, 1442012400, 1442016000, 1442019600, 1442023200, 
    1442026800, 1442030400, 1442034000, 1442037600, 1442041200, 1442044800, 
    1442048400, 1442052000, 1442055600, 1442059200, 1442062800, 1442066400, 
    1442070000, 1442073600, 1442077200, 1442080800, 1442084400, 1442088000, 
    1442091600, 1442095200, 1442098800, 1442102400, 1442106000, 1442109600, 
    1442113200, 1442116800, 1442120400, 1442124000, 1442127600, 1442131200, 
    1442134800, 1442138400, 1442142000, 1442145600, 1442149200, 1442152800, 
    1442156400, 1442160000, 1442163600, 1442167200, 1442170800, 1442174400, 
    1442178000, 1442181600, 1442185200, 1442188800, 1442192400, 1442196000, 
    1442199600, 1442203200, 1442206800, 1442210400, 1442214000, 1442217600, 
    1442221200, 1442224800, 1442228400, 1442232000, 1442235600, 1442239200, 
    1442242800, 1442246400, 1442250000, 1442253600, 1442257200, 1442260800, 
    1442264400, 1442268000, 1442271600, 1442275200, 1442278800, 1442282400, 
    1442286000, 1442289600, 1442293200, 1442296800, 1442300400, 1442304000, 
    1442307600, 1442311200, 1442314800, 1442318400, 1442322000, 1442325600, 
    1442329200, 1442332800, 1442336400, 1442340000, 1442343600, 1442347200, 
    1442350800, 1442354400, 1442358000, 1442361600, 1442365200, 1442368800, 
    1442372400, 1442376000, 1442379600, 1442383200, 1442386800, 1442390400, 
    1442394000, 1442397600, 1442401200, 1442404800, 1442408400, 1442412000, 
    1442415600, 1442419200, 1442422800, 1442426400, 1442430000, 1442433600, 
    1442437200, 1442440800, 1442444400, 1442448000, 1442451600, 1442455200, 
    1442458800, 1442462400, 1442466000, 1442469600, 1442473200, 1442476800, 
    1442480400, 1442484000, 1442487600, 1442491200, 1442494800, 1442498400, 
    1442502000, 1442505600, 1442509200, 1442512800, 1442516400, 1442520000, 
    1442523600, 1442527200, 1442530800, 1442534400, 1442538000, 1442541600, 
    1442545200, 1442548800, 1442552400, 1442556000, 1442559600, 1442563200, 
    1442566800, 1442570400, 1442574000, 1442577600, 1442581200, 1442584800, 
    1442588400, 1442592000, 1442595600, 1442599200, 1442602800, 1442606400, 
    1442610000, 1442613600, 1442617200, 1442620800, 1442624400, 1442628000, 
    1442631600, 1442635200, 1442638800, 1442642400, 1442646000, 1442649600, 
    1442653200, 1442656800, 1442660400, 1442664000, 1442667600, 1442671200, 
    1442674800, 1442678400, 1442682000, 1442685600, 1442689200, 1442692800, 
    1442696400, 1442700000, 1442703600, 1442707200, 1442710800, 1442714400, 
    1442718000, 1442721600, 1442725200, 1442728800, 1442732400, 1442736000, 
    1442739600, 1442743200, 1442746800, 1442750400, 1442754000, 1442757600, 
    1442761200, 1442764800, 1442768400, 1442772000, 1442775600, 1442779200, 
    1442782800, 1442786400, 1442790000, 1442793600, 1442797200, 1442800800, 
    1442804400, 1442808000, 1442811600, 1442815200, 1442818800, 1442822400, 
    1442826000, 1442829600, 1442833200, 1442836800, 1442840400, 1442844000, 
    1442847600, 1442851200, 1442854800, 1442858400, 1442862000, 1442865600, 
    1442869200, 1442872800, 1442876400, 1442880000, 1442883600, 1442887200, 
    1442890800, 1442894400, 1442898000, 1442901600, 1442905200, 1442908800, 
    1442912400, 1442916000, 1442919600, 1442923200, 1442926800, 1442930400, 
    1442934000, 1442937600, 1442941200, 1442944800, 1442948400, 1442952000, 
    1442955600, 1442959200, 1442962800, 1442966400, 1442970000, 1442973600, 
    1442977200, 1442980800, 1442984400, 1442988000, 1442991600, 1442995200, 
    1442998800, 1443002400, 1443006000, 1443009600, 1443013200, 1443016800, 
    1443020400, 1443024000, 1443027600, 1443031200, 1443034800, 1443038400, 
    1443042000, 1443045600, 1443049200, 1443052800, 1443056400, 1443060000, 
    1443063600, 1443067200, 1443070800, 1443074400, 1443078000, 1443081600, 
    1443085200, 1443088800, 1443092400, 1443096000, 1443099600, 1443103200, 
    1443106800, 1443110400, 1443114000, 1443117600, 1443121200, 1443124800, 
    1443128400, 1443132000, 1443135600, 1443139200, 1443142800, 1443146400, 
    1443150000, 1443153600, 1443157200, 1443160800, 1443164400, 1443168000, 
    1443171600, 1443175200, 1443178800, 1443182400, 1443186000, 1443189600, 
    1443193200, 1443196800, 1443200400, 1443204000, 1443207600, 1443211200, 
    1443214800, 1443218400, 1443222000, 1443225600, 1443229200, 1443232800, 
    1443236400, 1443240000, 1443243600, 1443247200, 1443250800, 1443254400, 
    1443258000, 1443261600, 1443265200, 1443268800, 1443272400, 1443276000, 
    1443279600, 1443283200, 1443286800, 1443290400, 1443294000, 1443297600, 
    1443301200, 1443304800, 1443308400, 1443312000, 1443315600, 1443319200, 
    1443322800, 1443326400, 1443330000, 1443333600, 1443337200, 1443340800, 
    1443344400, 1443348000, 1443351600, 1443355200, 1443358800, 1443362400, 
    1443366000, 1443369600, 1443373200, 1443376800, 1443380400, 1443384000, 
    1443387600, 1443391200, 1443394800, 1443398400, 1443402000, 1443405600, 
    1443409200, 1443412800, 1443416400, 1443420000, 1443423600, 1443427200, 
    1443430800, 1443434400, 1443438000, 1443441600, 1443445200, 1443448800, 
    1443452400, 1443456000, 1443459600, 1443463200, 1443466800, 1443470400, 
    1443474000, 1443477600, 1443481200, 1443484800, 1443488400, 1443492000, 
    1443495600, 1443499200, 1443502800, 1443506400, 1443510000, 1443513600, 
    1443517200, 1443520800, 1443524400, 1443528000, 1443531600, 1443535200, 
    1443538800, 1443542400, 1443546000, 1443549600, 1443553200, 1443556800, 
    1443560400, 1443564000, 1443567600, 1443571200, 1443574800, 1443578400, 
    1443582000, 1443585600, 1443589200, 1443592800, 1443596400, 1443600000, 
    1443603600, 1443607200, 1443610800, 1443614400, 1443618000, 1443621600, 
    1443625200, 1443628800, 1443632400, 1443636000, 1443639600, 1443643200, 
    1443646800, 1443650400, 1443654000, 1443657600, 1443661200, 1443664800, 
    1443668400, 1443672000, 1443675600, 1443679200, 1443682800, 1443686400, 
    1443690000, 1443693600, 1443697200, 1443700800, 1443704400, 1443708000, 
    1443711600, 1443715200, 1443718800, 1443722400, 1443726000, 1443729600, 
    1443733200, 1443736800, 1443740400, 1443744000, 1443747600, 1443751200, 
    1443754800, 1443758400, 1443762000, 1443765600, 1443769200, 1443772800, 
    1443776400, 1443780000, 1443783600, 1443787200, 1443790800, 1443794400, 
    1443798000, 1443801600, 1443805200, 1443808800, 1443812400, 1443816000, 
    1443819600, 1443823200, 1443826800, 1443830400, 1443834000, 1443837600, 
    1443841200, 1443844800, 1443848400, 1443852000, 1443855600, 1443859200, 
    1443862800, 1443866400, 1443870000, 1443873600, 1443877200, 1443880800, 
    1443884400, 1443888000, 1443891600, 1443895200, 1443898800, 1443902400, 
    1443906000, 1443909600, 1443913200, 1443916800, 1443920400, 1443924000, 
    1443927600, 1443931200, 1443934800, 1443938400, 1443942000, 1443945600, 
    1443949200, 1443952800, 1443956400, 1443960000, 1443963600, 1443967200, 
    1443970800, 1443974400, 1443978000, 1443981600, 1443985200, 1443988800, 
    1443992400, 1443996000, 1443999600, 1444003200, 1444006800, 1444010400, 
    1444014000, 1444017600, 1444021200, 1444024800, 1444028400, 1444032000, 
    1444035600, 1444039200, 1444042800, 1444046400, 1444050000, 1444053600, 
    1444057200, 1444060800, 1444064400, 1444068000, 1444071600, 1444075200, 
    1444078800, 1444082400, 1444086000, 1444089600, 1444093200, 1444096800, 
    1444100400, 1444104000, 1444107600, 1444111200, 1444114800, 1444118400, 
    1444122000, 1444125600, 1444129200, 1444132800, 1444136400, 1444140000, 
    1444143600, 1444147200, 1444150800, 1444154400, 1444158000, 1444161600, 
    1444165200, 1444168800, 1444172400, 1444176000, 1444179600, 1444183200, 
    1444186800, 1444190400, 1444194000, 1444197600, 1444201200, 1444204800, 
    1444208400, 1444212000, 1444215600, 1444219200, 1444222800, 1444226400, 
    1444230000, 1444233600, 1444237200, 1444240800, 1444244400, 1444248000, 
    1444251600, 1444255200, 1444258800, 1444262400, 1444266000, 1444269600, 
    1444273200, 1444276800, 1444280400, 1444284000, 1444287600, 1444291200, 
    1444294800, 1444298400, 1444302000, 1444305600, 1444309200, 1444312800, 
    1444316400, 1444320000, 1444323600, 1444327200, 1444330800, 1444334400, 
    1444338000, 1444341600, 1444345200, 1444348800, 1444352400, 1444356000, 
    1444359600, 1444363200, 1444366800, 1444370400, 1444374000, 1444377600, 
    1444381200, 1444384800, 1444388400, 1444392000, 1444395600, 1444399200, 
    1444402800, 1444406400, 1444410000, 1444413600, 1444417200, 1444420800, 
    1444424400, 1444428000, 1444431600, 1444435200, 1444438800, 1444442400, 
    1444446000, 1444449600, 1444453200, 1444456800, 1444460400, 1444464000, 
    1444467600, 1444471200, 1444474800, 1444478400, 1444482000, 1444485600, 
    1444489200, 1444492800, 1444496400, 1444500000, 1444503600, 1444507200, 
    1444510800, 1444514400, 1444518000, 1444521600, 1444525200, 1444528800, 
    1444532400, 1444536000, 1444539600, 1444543200, 1444546800, 1444550400, 
    1444554000, 1444557600, 1444561200, 1444564800, 1444568400, 1444572000, 
    1444575600, 1444579200, 1444582800, 1444586400, 1444590000, 1444593600, 
    1444597200, 1444600800, 1444604400, 1444608000, 1444611600, 1444615200, 
    1444618800, 1444622400, 1444626000, 1444629600, 1444633200, 1444636800, 
    1444640400, 1444644000, 1444647600, 1444651200, 1444654800, 1444658400, 
    1444662000, 1444665600, 1444669200, 1444672800, 1444676400, 1444680000, 
    1444683600, 1444687200, 1444690800, 1444694400, 1444698000, 1444701600, 
    1444705200, 1444708800, 1444712400, 1444716000, 1444719600, 1444723200, 
    1444726800, 1444730400, 1444734000, 1444737600, 1444741200, 1444744800, 
    1444748400, 1444752000, 1444755600, 1444759200, 1444762800, 1444766400, 
    1444770000, 1444773600, 1444777200, 1444780800, 1444784400, 1444788000, 
    1444791600, 1444795200, 1444798800, 1444802400, 1444806000, 1444809600, 
    1444813200, 1444816800, 1444820400, 1444824000, 1444827600, 1444831200, 
    1444834800, 1444838400, 1444842000, 1444845600, 1444849200, 1444852800, 
    1444856400, 1444860000, 1444863600, 1444867200, 1444870800, 1444874400, 
    1444878000, 1444881600, 1444885200, 1444888800, 1444892400, 1444896000, 
    1444899600, 1444903200, 1444906800, 1444910400, 1444914000, 1444917600, 
    1444921200, 1444924800, 1444928400, 1444932000, 1444935600, 1444939200, 
    1444942800, 1444946400, 1444950000, 1444953600, 1444957200, 1444960800, 
    1444964400, 1444968000, 1444971600, 1444975200, 1444978800, 1444982400, 
    1444986000, 1444989600, 1444993200, 1444996800, 1445000400, 1445004000, 
    1445007600, 1445011200, 1445014800, 1445018400, 1445022000, 1445025600, 
    1445029200, 1445032800, 1445036400, 1445040000, 1445043600, 1445047200, 
    1445050800, 1445054400, 1445058000, 1445061600, 1445065200, 1445068800, 
    1445072400, 1445076000, 1445079600, 1445083200, 1445086800, 1445090400, 
    1445094000, 1445097600, 1445101200, 1445104800, 1445108400, 1445112000, 
    1445115600, 1445119200, 1445122800, 1445126400, 1445130000, 1445133600, 
    1445137200, 1445140800, 1445144400, 1445148000, 1445151600, 1445155200, 
    1445158800, 1445162400, 1445166000, 1445169600, 1445173200, 1445176800, 
    1445180400, 1445184000, 1445187600, 1445191200, 1445194800, 1445198400, 
    1445202000, 1445205600, 1445209200, 1445212800, 1445216400, 1445220000, 
    1445223600, 1445227200, 1445230800, 1445234400, 1445238000, 1445241600, 
    1445245200, 1445248800, 1445252400, 1445256000, 1445259600, 1445263200, 
    1445266800, 1445270400, 1445274000, 1445277600, 1445281200, 1445284800, 
    1445288400, 1445292000, 1445295600, 1445299200, 1445302800, 1445306400, 
    1445310000, 1445313600, 1445317200, 1445320800, 1445324400, 1445328000, 
    1445331600, 1445335200, 1445338800, 1445342400, 1445346000, 1445349600, 
    1445353200, 1445356800, 1445360400, 1445364000, 1445367600, 1445371200, 
    1445374800, 1445378400, 1445382000, 1445385600, 1445389200, 1445392800, 
    1445396400, 1445400000, 1445403600, 1445407200, 1445410800, 1445414400, 
    1445418000, 1445421600, 1445425200, 1445428800, 1445432400, 1445436000, 
    1445439600, 1445443200, 1445446800, 1445450400, 1445454000, 1445457600, 
    1445461200, 1445464800, 1445468400, 1445472000, 1445475600, 1445479200, 
    1445482800, 1445486400, 1445490000, 1445493600, 1445497200, 1445500800, 
    1445504400, 1445508000, 1445511600, 1445515200, 1445518800, 1445522400, 
    1445526000, 1445529600, 1445533200, 1445536800, 1445540400, 1445544000, 
    1445547600, 1445551200, 1445554800, 1445558400, 1445562000, 1445565600, 
    1445569200, 1445572800, 1445576400, 1445580000, 1445583600, 1445587200, 
    1445590800, 1445594400, 1445598000, 1445601600, 1445605200, 1445608800, 
    1445612400, 1445616000, 1445619600, 1445623200, 1445626800, 1445630400, 
    1445634000, 1445637600, 1445641200, 1445644800, 1445648400, 1445652000, 
    1445655600, 1445659200, 1445662800, 1445666400, 1445670000, 1445673600, 
    1445677200, 1445680800, 1445684400, 1445688000, 1445691600, 1445695200, 
    1445698800, 1445702400, 1445706000, 1445709600, 1445713200, 1445716800, 
    1445720400, 1445724000, 1445727600, 1445731200, 1445734800, 1445738400, 
    1445742000, 1445745600, 1445749200, 1445752800, 1445756400, 1445760000, 
    1445763600, 1445767200, 1445770800, 1445774400, 1445778000, 1445781600, 
    1445785200, 1445788800, 1445792400, 1445796000, 1445799600, 1445803200, 
    1445806800, 1445810400, 1445814000, 1445817600, 1445821200, 1445824800, 
    1445828400, 1445832000, 1445835600, 1445839200, 1445842800, 1445846400, 
    1445850000, 1445853600, 1445857200, 1445860800, 1445864400, 1445868000, 
    1445871600, 1445875200, 1445878800, 1445882400, 1445886000, 1445889600, 
    1445893200, 1445896800, 1445900400, 1445904000, 1445907600, 1445911200, 
    1445914800, 1445918400, 1445922000, 1445925600, 1445929200, 1445932800, 
    1445936400, 1445940000, 1445943600, 1445947200, 1445950800, 1445954400, 
    1445958000, 1445961600, 1445965200, 1445968800, 1445972400, 1445976000, 
    1445979600, 1445983200, 1445986800, 1445990400, 1445994000, 1445997600, 
    1446001200, 1446004800, 1446008400, 1446012000, 1446015600, 1446019200, 
    1446022800, 1446026400, 1446030000, 1446033600, 1446037200, 1446040800, 
    1446044400, 1446048000, 1446051600, 1446055200, 1446058800, 1446062400, 
    1446066000, 1446069600, 1446073200, 1446076800, 1446080400, 1446084000, 
    1446087600, 1446091200, 1446094800, 1446098400, 1446102000, 1446105600, 
    1446109200, 1446112800, 1446116400, 1446120000, 1446123600, 1446127200, 
    1446130800, 1446134400, 1446138000, 1446141600, 1446145200, 1446148800, 
    1446152400, 1446156000, 1446159600, 1446163200, 1446166800, 1446170400, 
    1446174000, 1446177600, 1446181200, 1446184800, 1446188400, 1446192000, 
    1446195600, 1446199200, 1446202800, 1446206400, 1446210000, 1446213600, 
    1446217200, 1446220800, 1446224400, 1446228000, 1446231600, 1446235200, 
    1446238800, 1446242400, 1446246000, 1446249600, 1446253200, 1446256800, 
    1446260400, 1446264000, 1446267600, 1446271200, 1446274800, 1446278400, 
    1446282000, 1446285600, 1446289200, 1446292800, 1446296400, 1446300000, 
    1446303600, 1446307200, 1446310800, 1446314400, 1446318000, 1446321600, 
    1446325200, 1446328800, 1446332400, 1446336000, 1446339600, 1446343200, 
    1446346800, 1446350400, 1446354000, 1446357600, 1446361200, 1446364800, 
    1446368400, 1446372000, 1446375600, 1446379200, 1446382800, 1446386400, 
    1446390000, 1446393600, 1446397200, 1446400800, 1446404400, 1446408000, 
    1446411600, 1446415200, 1446418800, 1446422400, 1446426000, 1446429600, 
    1446433200, 1446436800, 1446440400, 1446444000, 1446447600, 1446451200, 
    1446454800, 1446458400, 1446462000, 1446465600, 1446469200, 1446472800, 
    1446476400, 1446480000, 1446483600, 1446487200, 1446490800, 1446494400, 
    1446498000, 1446501600, 1446505200, 1446508800, 1446512400, 1446516000, 
    1446519600, 1446523200, 1446526800, 1446530400, 1446534000, 1446537600, 
    1446541200, 1446544800, 1446548400, 1446552000, 1446555600, 1446559200, 
    1446562800, 1446566400, 1446570000, 1446573600, 1446577200, 1446580800, 
    1446584400, 1446588000, 1446591600, 1446595200, 1446598800, 1446602400, 
    1446606000, 1446609600, 1446613200, 1446616800, 1446620400, 1446624000, 
    1446627600, 1446631200, 1446634800, 1446638400, 1446642000, 1446645600, 
    1446649200, 1446652800, 1446656400, 1446660000, 1446663600, 1446667200, 
    1446670800, 1446674400, 1446678000, 1446681600, 1446685200, 1446688800, 
    1446692400, 1446696000, 1446699600, 1446703200, 1446706800, 1446710400, 
    1446714000, 1446717600, 1446721200, 1446724800, 1446728400, 1446732000, 
    1446735600, 1446739200, 1446742800, 1446746400, 1446750000, 1446753600, 
    1446757200, 1446760800, 1446764400, 1446768000, 1446771600, 1446775200, 
    1446778800, 1446782400, 1446786000, 1446789600, 1446793200, 1446796800, 
    1446800400, 1446804000, 1446807600, 1446811200, 1446814800, 1446818400, 
    1446822000, 1446825600, 1446829200, 1446832800, 1446836400, 1446840000, 
    1446843600, 1446847200, 1446850800, 1446854400, 1446858000, 1446861600, 
    1446865200, 1446868800, 1446872400, 1446876000, 1446879600, 1446883200, 
    1446886800, 1446890400, 1446894000, 1446897600, 1446901200, 1446904800, 
    1446908400, 1446912000, 1446915600, 1446919200, 1446922800, 1446926400, 
    1446930000, 1446933600, 1446937200, 1446940800, 1446944400, 1446948000, 
    1446951600, 1446955200, 1446958800, 1446962400, 1446966000, 1446969600, 
    1446973200, 1446976800, 1446980400, 1446984000, 1446987600, 1446991200, 
    1446994800, 1446998400, 1447002000, 1447005600, 1447009200, 1447012800, 
    1447016400, 1447020000, 1447023600, 1447027200, 1447030800, 1447034400, 
    1447038000, 1447041600, 1447045200, 1447048800, 1447052400, 1447056000, 
    1447059600, 1447063200, 1447066800, 1447070400, 1447074000, 1447077600, 
    1447081200, 1447084800, 1447088400, 1447092000, 1447095600, 1447099200, 
    1447102800, 1447106400, 1447110000, 1447113600, 1447117200, 1447120800, 
    1447124400, 1447128000, 1447131600, 1447135200, 1447138800, 1447142400, 
    1447146000, 1447149600, 1447153200, 1447156800, 1447160400, 1447164000, 
    1447167600, 1447171200, 1447174800, 1447178400, 1447182000, 1447185600, 
    1447189200, 1447192800, 1447196400, 1447200000, 1447203600, 1447207200, 
    1447210800, 1447214400, 1447218000, 1447221600, 1447225200, 1447228800, 
    1447232400, 1447236000, 1447239600, 1447243200, 1447246800, 1447250400, 
    1447254000, 1447257600, 1447261200, 1447264800, 1447268400, 1447272000, 
    1447275600, 1447279200, 1447282800, 1447286400, 1447290000, 1447293600, 
    1447297200, 1447300800, 1447304400, 1447308000, 1447311600, 1447315200, 
    1447318800, 1447322400, 1447326000, 1447329600, 1447333200, 1447336800, 
    1447340400, 1447344000, 1447347600, 1447351200, 1447354800, 1447358400, 
    1447362000, 1447365600, 1447369200, 1447372800, 1447376400, 1447380000, 
    1447383600, 1447387200, 1447390800, 1447394400, 1447398000, 1447401600, 
    1447405200, 1447408800, 1447412400, 1447416000, 1447419600, 1447423200, 
    1447426800, 1447430400, 1447434000, 1447437600, 1447441200, 1447444800, 
    1447448400, 1447452000, 1447455600, 1447459200, 1447462800, 1447466400, 
    1447470000, 1447473600, 1447477200, 1447480800, 1447484400, 1447488000, 
    1447491600, 1447495200, 1447498800, 1447502400, 1447506000, 1447509600, 
    1447513200, 1447516800, 1447520400, 1447524000, 1447527600, 1447531200, 
    1447534800, 1447538400, 1447542000, 1447545600, 1447549200, 1447552800, 
    1447556400, 1447560000, 1447563600, 1447567200, 1447570800, 1447574400, 
    1447578000, 1447581600, 1447585200, 1447588800, 1447592400, 1447596000, 
    1447599600, 1447603200, 1447606800, 1447610400, 1447614000, 1447617600, 
    1447621200, 1447624800, 1447628400, 1447632000, 1447635600, 1447639200, 
    1447642800, 1447646400, 1447650000, 1447653600, 1447657200, 1447660800, 
    1447664400, 1447668000, 1447671600, 1447675200, 1447678800, 1447682400, 
    1447686000, 1447689600, 1447693200, 1447696800, 1447700400, 1447704000, 
    1447707600, 1447711200, 1447714800, 1447718400, 1447722000, 1447725600, 
    1447729200, 1447732800, 1447736400, 1447740000, 1447743600, 1447747200, 
    1447750800, 1447754400, 1447758000, 1447761600, 1447765200, 1447768800, 
    1447772400, 1447776000, 1447779600, 1447783200, 1447786800, 1447790400, 
    1447794000, 1447797600, 1447801200, 1447804800, 1447808400, 1447812000, 
    1447815600, 1447819200, 1447822800, 1447826400, 1447830000, 1447833600, 
    1447837200, 1447840800, 1447844400, 1447848000, 1447851600, 1447855200, 
    1447858800, 1447862400, 1447866000, 1447869600, 1447873200, 1447876800, 
    1447880400, 1447884000, 1447887600, 1447891200, 1447894800, 1447898400, 
    1447902000, 1447905600, 1447909200, 1447912800, 1447916400, 1447920000, 
    1447923600, 1447927200, 1447930800, 1447934400, 1447938000, 1447941600, 
    1447945200, 1447948800, 1447952400, 1447956000, 1447959600, 1447963200, 
    1447966800, 1447970400, 1447974000, 1447977600, 1447981200, 1447984800, 
    1447988400, 1447992000, 1447995600, 1447999200, 1448002800, 1448006400, 
    1448010000, 1448013600, 1448017200, 1448020800, 1448024400, 1448028000, 
    1448031600, 1448035200, 1448038800, 1448042400, 1448046000, 1448049600, 
    1448053200, 1448056800, 1448060400, 1448064000, 1448067600, 1448071200, 
    1448074800, 1448078400, 1448082000, 1448085600, 1448089200, 1448092800, 
    1448096400, 1448100000, 1448103600, 1448107200, 1448110800, 1448114400, 
    1448118000, 1448121600, 1448125200, 1448128800, 1448132400, 1448136000, 
    1448139600, 1448143200, 1448146800, 1448150400, 1448154000, 1448157600, 
    1448161200, 1448164800, 1448168400, 1448172000, 1448175600, 1448179200, 
    1448182800, 1448186400, 1448190000, 1448193600, 1448197200, 1448200800, 
    1448204400, 1448208000, 1448211600, 1448215200, 1448218800, 1448222400, 
    1448226000, 1448229600, 1448233200, 1448236800, 1448240400, 1448244000, 
    1448247600, 1448251200, 1448254800, 1448258400, 1448262000, 1448265600, 
    1448269200, 1448272800, 1448276400, 1448280000, 1448283600, 1448287200, 
    1448290800, 1448294400, 1448298000, 1448301600, 1448305200, 1448308800, 
    1448312400, 1448316000, 1448319600, 1448323200, 1448326800, 1448330400, 
    1448334000, 1448337600, 1448341200, 1448344800, 1448348400, 1448352000, 
    1448355600, 1448359200, 1448362800, 1448366400, 1448370000, 1448373600, 
    1448377200, 1448380800, 1448384400, 1448388000, 1448391600, 1448395200, 
    1448398800, 1448402400, 1448406000, 1448409600, 1448413200, 1448416800, 
    1448420400, 1448424000, 1448427600, 1448431200, 1448434800, 1448438400, 
    1448442000, 1448445600, 1448449200, 1448452800, 1448456400, 1448460000, 
    1448463600, 1448467200, 1448470800, 1448474400, 1448478000, 1448481600, 
    1448485200, 1448488800, 1448492400, 1448496000, 1448499600, 1448503200, 
    1448506800, 1448510400, 1448514000, 1448517600, 1448521200, 1448524800, 
    1448528400, 1448532000, 1448535600, 1448539200, 1448542800, 1448546400, 
    1448550000, 1448553600, 1448557200, 1448560800, 1448564400, 1448568000, 
    1448571600, 1448575200, 1448578800, 1448582400, 1448586000, 1448589600, 
    1448593200, 1448596800, 1448600400, 1448604000, 1448607600, 1448611200, 
    1448614800, 1448618400, 1448622000, 1448625600, 1448629200, 1448632800, 
    1448636400, 1448640000, 1448643600, 1448647200, 1448650800, 1448654400, 
    1448658000, 1448661600, 1448665200, 1448668800, 1448672400, 1448676000, 
    1448679600, 1448683200, 1448686800, 1448690400, 1448694000, 1448697600, 
    1448701200, 1448704800, 1448708400, 1448712000, 1448715600, 1448719200, 
    1448722800, 1448726400, 1448730000, 1448733600, 1448737200, 1448740800, 
    1448744400, 1448748000, 1448751600, 1448755200, 1448758800, 1448762400, 
    1448766000, 1448769600, 1448773200, 1448776800, 1448780400, 1448784000, 
    1448787600, 1448791200, 1448794800, 1448798400, 1448802000, 1448805600, 
    1448809200, 1448812800, 1448816400, 1448820000, 1448823600, 1448827200, 
    1448830800, 1448834400, 1448838000, 1448841600, 1448845200, 1448848800, 
    1448852400, 1448856000, 1448859600, 1448863200, 1448866800, 1448870400, 
    1448874000, 1448877600, 1448881200, 1448884800, 1448888400, 1448892000, 
    1448895600, 1448899200, 1448902800, 1448906400, 1448910000, 1448913600, 
    1448917200, 1448920800, 1448924400, 1448928000, 1448931600, 1448935200, 
    1448938800, 1448942400, 1448946000, 1448949600, 1448953200, 1448956800, 
    1448960400, 1448964000, 1448967600, 1448971200, 1448974800, 1448978400, 
    1448982000, 1448985600, 1448989200, 1448992800, 1448996400, 1449000000, 
    1449003600, 1449007200, 1449010800, 1449014400, 1449018000, 1449021600, 
    1449025200, 1449028800, 1449032400, 1449036000, 1449039600, 1449043200, 
    1449046800, 1449050400, 1449054000, 1449057600, 1449061200, 1449064800, 
    1449068400, 1449072000, 1449075600, 1449079200, 1449082800, 1449086400, 
    1449090000, 1449093600, 1449097200, 1449100800, 1449104400, 1449108000, 
    1449111600, 1449115200, 1449118800, 1449122400, 1449126000, 1449129600, 
    1449133200, 1449136800, 1449140400, 1449144000, 1449147600, 1449151200, 
    1449154800, 1449158400, 1449162000, 1449165600, 1449169200, 1449172800, 
    1449176400, 1449180000, 1449183600, 1449187200, 1449190800, 1449194400, 
    1449198000, 1449201600, 1449205200, 1449208800, 1449212400, 1449216000, 
    1449219600, 1449223200, 1449226800, 1449230400, 1449234000, 1449237600, 
    1449241200, 1449244800, 1449248400, 1449252000, 1449255600, 1449259200, 
    1449262800, 1449266400, 1449270000, 1449273600, 1449277200, 1449280800, 
    1449284400, 1449288000, 1449291600, 1449295200, 1449298800, 1449302400, 
    1449306000, 1449309600, 1449313200, 1449316800, 1449320400, 1449324000, 
    1449327600, 1449331200, 1449334800, 1449338400, 1449342000, 1449345600, 
    1449349200, 1449352800, 1449356400, 1449360000, 1449363600, 1449367200, 
    1449370800, 1449374400, 1449378000, 1449381600, 1449385200, 1449388800, 
    1449392400, 1449396000, 1449399600, 1449403200, 1449406800, 1449410400, 
    1449414000, 1449417600, 1449421200, 1449424800, 1449428400, 1449432000, 
    1449435600, 1449439200, 1449442800, 1449446400, 1449450000, 1449453600, 
    1449457200, 1449460800, 1449464400, 1449468000, 1449471600, 1449475200, 
    1449478800, 1449482400, 1449486000, 1449489600, 1449493200, 1449496800, 
    1449500400, 1449504000, 1449507600, 1449511200, 1449514800, 1449518400, 
    1449522000, 1449525600, 1449529200, 1449532800, 1449536400, 1449540000, 
    1449543600, 1449547200, 1449550800, 1449554400, 1449558000, 1449561600, 
    1449565200, 1449568800, 1449572400, 1449576000, 1449579600, 1449583200, 
    1449586800, 1449590400, 1449594000, 1449597600, 1449601200, 1449604800, 
    1449608400, 1449612000, 1449615600, 1449619200, 1449622800, 1449626400, 
    1449630000, 1449633600, 1449637200, 1449640800, 1449644400, 1449648000, 
    1449651600, 1449655200, 1449658800, 1449662400, 1449666000, 1449669600, 
    1449673200, 1449676800, 1449680400, 1449684000, 1449687600, 1449691200, 
    1449694800, 1449698400, 1449702000, 1449705600, 1449709200, 1449712800, 
    1449716400, 1449720000, 1449723600, 1449727200, 1449730800, 1449734400, 
    1449738000, 1449741600, 1449745200, 1449748800, 1449752400, 1449756000, 
    1449759600, 1449763200, 1449766800, 1449770400, 1449774000, 1449777600, 
    1449781200, 1449784800, 1449788400, 1449792000, 1449795600, 1449799200, 
    1449802800, 1449806400, 1449810000, 1449813600, 1449817200, 1449820800, 
    1449824400, 1449828000, 1449831600, 1449835200, 1449838800, 1449842400, 
    1449846000, 1449849600, 1449853200, 1449856800, 1449860400, 1449864000, 
    1449867600, 1449871200, 1449874800, 1449878400, 1449882000, 1449885600, 
    1449889200, 1449892800, 1449896400, 1449900000, 1449903600, 1449907200, 
    1449910800, 1449914400, 1449918000, 1449921600, 1449925200, 1449928800, 
    1449932400, 1449936000, 1449939600, 1449943200, 1449946800, 1449950400, 
    1449954000, 1449957600, 1449961200, 1449964800, 1449968400, 1449972000, 
    1449975600, 1449979200, 1449982800, 1449986400, 1449990000, 1449993600, 
    1449997200, 1450000800, 1450004400, 1450008000, 1450011600, 1450015200, 
    1450018800, 1450022400, 1450026000, 1450029600, 1450033200, 1450036800, 
    1450040400, 1450044000, 1450047600, 1450051200, 1450054800, 1450058400, 
    1450062000, 1450065600, 1450069200, 1450072800, 1450076400, 1450080000, 
    1450083600, 1450087200, 1450090800, 1450094400, 1450098000, 1450101600, 
    1450105200, 1450108800, 1450112400, 1450116000, 1450119600, 1450123200, 
    1450126800, 1450130400, 1450134000, 1450137600, 1450141200, 1450144800, 
    1450148400, 1450152000, 1450155600, 1450159200, 1450162800, 1450166400, 
    1450170000, 1450173600, 1450177200, 1450180800, 1450184400, 1450188000, 
    1450191600, 1450195200, 1450198800, 1450202400, 1450206000, 1450209600, 
    1450213200, 1450216800, 1450220400, 1450224000, 1450227600, 1450231200, 
    1450234800, 1450238400, 1450242000, 1450245600, 1450249200, 1450252800, 
    1450256400, 1450260000, 1450263600, 1450267200, 1450270800, 1450274400, 
    1450278000, 1450281600, 1450285200, 1450288800, 1450292400, 1450296000, 
    1450299600, 1450303200, 1450306800, 1450310400, 1450314000, 1450317600, 
    1450321200, 1450324800, 1450328400, 1450332000, 1450335600, 1450339200, 
    1450342800, 1450346400, 1450350000, 1450353600, 1450357200, 1450360800, 
    1450364400, 1450368000, 1450371600, 1450375200, 1450378800, 1450382400, 
    1450386000, 1450389600, 1450393200, 1450396800, 1450400400, 1450404000, 
    1450407600, 1450411200, 1450414800, 1450418400, 1450422000, 1450425600, 
    1450429200, 1450432800, 1450436400, 1450440000, 1450443600, 1450447200, 
    1450450800, 1450454400, 1450458000, 1450461600, 1450465200, 1450468800, 
    1450472400, 1450476000, 1450479600, 1450483200, 1450486800, 1450490400, 
    1450494000, 1450497600, 1450501200, 1450504800, 1450508400, 1450512000, 
    1450515600, 1450519200, 1450522800, 1450526400, 1450530000, 1450533600, 
    1450537200, 1450540800, 1450544400, 1450548000, 1450551600, 1450555200, 
    1450558800, 1450562400, 1450566000, 1450569600, 1450573200, 1450576800, 
    1450580400, 1450584000, 1450587600, 1450591200, 1450594800, 1450598400, 
    1450602000, 1450605600, 1450609200, 1450612800, 1450616400, 1450620000, 
    1450623600, 1450627200, 1450630800, 1450634400, 1450638000, 1450641600, 
    1450645200, 1450648800, 1450652400, 1450656000, 1450659600, 1450663200, 
    1450666800, 1450670400, 1450674000, 1450677600, 1450681200, 1450684800, 
    1450688400, 1450692000, 1450695600, 1450699200, 1450702800, 1450706400, 
    1450710000, 1450713600, 1450717200, 1450720800, 1450724400, 1450728000, 
    1450731600, 1450735200, 1450738800, 1450742400, 1450746000, 1450749600, 
    1450753200, 1450756800, 1450760400, 1450764000, 1450767600, 1450771200, 
    1450774800, 1450778400, 1450782000, 1450785600, 1450789200, 1450792800, 
    1450796400, 1450800000, 1450803600, 1450807200, 1450810800, 1450814400, 
    1450818000, 1450821600, 1450825200, 1450828800, 1450832400, 1450836000, 
    1450839600, 1450843200, 1450846800, 1450850400, 1450854000, 1450857600, 
    1450861200, 1450864800, 1450868400, 1450872000, 1450875600, 1450879200, 
    1450882800, 1450886400, 1450890000, 1450893600, 1450897200, 1450900800, 
    1450904400, 1450908000, 1450911600, 1450915200, 1450918800, 1450922400, 
    1450926000, 1450929600, 1450933200, 1450936800, 1450940400, 1450944000, 
    1450947600, 1450951200, 1450954800, 1450958400, 1450962000, 1450965600, 
    1450969200, 1450972800, 1450976400, 1450980000, 1450983600, 1450987200, 
    1450990800, 1450994400, 1450998000, 1451001600, 1451005200, 1451008800, 
    1451012400, 1451016000, 1451019600, 1451023200, 1451026800, 1451030400, 
    1451034000, 1451037600, 1451041200, 1451044800, 1451048400, 1451052000, 
    1451055600, 1451059200, 1451062800, 1451066400, 1451070000, 1451073600, 
    1451077200, 1451080800, 1451084400, 1451088000, 1451091600, 1451095200, 
    1451098800, 1451102400, 1451106000, 1451109600, 1451113200, 1451116800, 
    1451120400, 1451124000, 1451127600, 1451131200, 1451134800, 1451138400, 
    1451142000, 1451145600, 1451149200, 1451152800, 1451156400, 1451160000, 
    1451163600, 1451167200, 1451170800, 1451174400, 1451178000, 1451181600, 
    1451185200, 1451188800, 1451192400, 1451196000, 1451199600, 1451203200, 
    1451206800, 1451210400, 1451214000, 1451217600, 1451221200, 1451224800, 
    1451228400, 1451232000, 1451235600, 1451239200, 1451242800, 1451246400, 
    1451250000, 1451253600, 1451257200, 1451260800, 1451264400, 1451268000, 
    1451271600, 1451275200, 1451278800, 1451282400, 1451286000, 1451289600, 
    1451293200, 1451296800, 1451300400, 1451304000, 1451307600, 1451311200, 
    1451314800, 1451318400, 1451322000, 1451325600, 1451329200, 1451332800, 
    1451336400, 1451340000, 1451343600, 1451347200, 1451350800, 1451354400, 
    1451358000, 1451361600, 1451365200, 1451368800, 1451372400, 1451376000, 
    1451379600, 1451383200, 1451386800, 1451390400, 1451394000, 1451397600, 
    1451401200, 1451404800, 1451408400, 1451412000, 1451415600, 1451419200, 
    1451422800, 1451426400, 1451430000, 1451433600, 1451437200, 1451440800, 
    1451444400, 1451448000, 1451451600, 1451455200, 1451458800, 1451462400, 
    1451466000, 1451469600, 1451473200, 1451476800, 1451480400, 1451484000, 
    1451487600, 1451491200, 1451494800, 1451498400, 1451502000, 1451505600, 
    1451509200, 1451512800, 1451516400, 1451520000, 1451523600, 1451527200, 
    1451530800, 1451534400, 1451548800, 1451552400, 1451566800, 1451570400, 
    1451574000, 1451577600, 1451592000, 1451602800, 1451606400, 1451610000, 
    1451613600, 1451617200, 1451620800, 1451624400, 1451628000, 1451631600, 
    1451635200, 1451638800, 1451642400, 1451646000, 1451649600, 1451653200, 
    1451656800, 1451660400, 1451664000, 1451667600, 1451671200, 1451674800, 
    1451678400, 1451682000, 1451685600, 1451689200, 1451692800, 1451696400, 
    1451700000, 1451703600, 1451707200, 1451710800, 1451714400, 1451718000, 
    1451721600, 1451725200, 1451728800, 1451732400, 1451736000, 1451739600, 
    1451743200, 1451746800, 1451750400, 1451754000, 1451757600, 1451761200, 
    1451764800, 1451768400, 1451772000, 1451775600, 1451779200, 1451782800, 
    1451786400, 1451790000, 1451793600, 1451797200, 1451800800, 1451804400, 
    1451808000, 1451811600, 1451815200, 1451818800, 1451822400, 1451826000, 
    1451829600, 1451833200, 1451836800, 1451840400, 1451844000, 1451847600, 
    1451851200, 1451854800, 1451858400, 1451862000, 1451865600, 1451869200, 
    1451872800, 1451876400, 1451880000, 1451883600, 1451887200, 1451890800, 
    1451894400, 1451898000, 1451901600, 1451905200, 1451908800, 1451912400, 
    1451916000, 1451919600, 1451923200, 1451926800, 1451930400, 1451934000, 
    1451937600, 1451941200, 1451944800, 1451948400, 1451952000, 1451955600, 
    1451959200, 1451962800, 1451966400, 1451970000, 1451973600, 1451977200, 
    1451980800, 1451984400, 1451988000, 1451991600, 1451995200, 1451998800, 
    1452002400, 1452006000, 1452009600, 1452013200, 1452016800, 1452020400, 
    1452024000, 1452027600, 1452031200, 1452034800, 1452038400, 1452042000, 
    1452045600, 1452049200, 1452052800, 1452056400, 1452060000, 1452063600, 
    1452067200, 1452070800, 1452074400, 1452078000, 1452081600, 1452085200, 
    1452088800, 1452092400, 1452096000, 1452099600, 1452103200, 1452106800, 
    1452110400, 1452114000, 1452117600, 1452121200, 1452124800, 1452128400, 
    1452132000, 1452135600, 1452139200, 1452142800, 1452146400, 1452150000, 
    1452153600, 1452157200, 1452160800, 1452164400, 1452168000, 1452171600, 
    1452175200, 1452178800, 1452182400, 1452186000, 1452189600, 1452193200, 
    1452196800, 1452200400, 1452204000, 1452207600, 1452211200, 1452214800, 
    1452218400, 1452222000, 1452225600, 1452229200, 1452232800, 1452236400, 
    1452240000, 1452243600, 1452247200, 1452250800, 1452254400, 1452258000, 
    1452261600, 1452265200, 1452268800, 1452272400, 1452276000, 1452279600, 
    1452283200, 1452286800, 1452290400, 1452294000, 1452297600, 1452301200, 
    1452304800, 1452308400, 1452312000, 1452315600, 1452319200, 1452322800, 
    1452326400, 1452330000, 1452333600, 1452337200, 1452340800, 1452344400, 
    1452348000, 1452351600, 1452355200, 1452358800, 1452362400, 1452366000, 
    1452369600, 1452373200, 1452376800, 1452380400, 1452384000, 1452387600, 
    1452391200, 1452394800, 1452398400, 1452402000, 1452405600, 1452409200, 
    1452412800, 1452416400, 1452420000, 1452423600, 1452427200, 1452430800, 
    1452434400, 1452438000, 1452441600, 1452445200, 1452448800, 1452452400, 
    1452456000, 1452459600, 1452463200, 1452466800, 1452470400, 1452474000, 
    1452477600, 1452481200, 1452484800, 1452488400, 1452492000, 1452495600, 
    1452499200, 1452502800, 1452506400, 1452510000, 1452513600, 1452517200, 
    1452520800, 1452524400, 1452528000, 1452531600, 1452535200, 1452538800, 
    1452542400, 1452546000, 1452549600, 1452553200, 1452556800, 1452560400, 
    1452564000, 1452567600, 1452571200, 1452574800, 1452578400, 1452582000, 
    1452585600, 1452589200, 1452592800, 1452596400, 1452600000, 1452603600, 
    1452607200, 1452610800, 1452614400, 1452618000, 1452621600, 1452625200, 
    1452628800, 1452632400, 1452636000, 1452639600, 1452643200, 1452646800, 
    1452650400, 1452654000, 1452657600, 1452661200, 1452664800, 1452668400, 
    1452672000, 1452675600, 1452679200, 1452682800, 1452686400, 1452690000, 
    1452693600, 1452697200, 1452700800, 1452704400, 1452708000, 1452711600, 
    1452715200, 1452718800, 1452722400, 1452726000, 1452729600, 1452733200, 
    1452736800, 1452740400, 1452744000, 1452747600, 1452751200, 1452754800, 
    1452758400, 1452762000, 1452765600, 1452769200, 1452772800, 1452776400, 
    1452780000, 1452783600, 1452787200, 1452790800, 1452794400, 1452798000, 
    1452801600, 1452805200, 1452808800, 1452812400, 1452816000, 1452819600, 
    1452823200, 1452826800, 1452830400, 1452834000, 1452837600, 1452841200, 
    1452844800, 1452848400, 1452852000, 1452855600, 1452859200, 1452862800, 
    1452866400, 1452870000, 1452873600, 1452877200, 1452880800, 1452884400, 
    1452888000, 1452891600, 1452895200, 1452898800, 1452902400, 1452906000, 
    1452909600, 1452913200, 1452916800, 1452920400, 1452924000, 1452927600, 
    1452931200, 1452934800, 1452938400, 1452942000, 1452945600, 1452949200, 
    1452952800, 1452956400, 1452960000, 1452963600, 1452967200, 1452970800, 
    1452974400, 1452978000, 1452981600, 1452985200, 1452988800, 1452992400, 
    1452996000, 1452999600, 1453003200, 1453006800, 1453010400, 1453014000, 
    1453017600, 1453021200, 1453024800, 1453028400, 1453032000, 1453035600, 
    1453039200, 1453042800, 1453046400, 1453050000, 1453053600, 1453057200, 
    1453060800, 1453064400, 1453068000, 1453071600, 1453075200, 1453078800, 
    1453082400, 1453086000, 1453089600, 1453093200, 1453096800, 1453100400, 
    1453104000, 1453107600, 1453111200, 1453114800, 1453118400, 1453122000, 
    1453125600, 1453129200, 1453132800, 1453136400, 1453140000, 1453143600, 
    1453147200, 1453150800, 1453154400, 1453158000, 1453161600, 1453165200, 
    1453168800, 1453172400, 1453176000, 1453179600, 1453183200, 1453186800, 
    1453190400, 1453194000, 1453197600, 1453201200, 1453204800, 1453208400, 
    1453212000, 1453215600, 1453219200, 1453222800, 1453226400, 1453230000, 
    1453233600, 1453237200, 1453240800, 1453244400, 1453248000, 1453251600, 
    1453255200, 1453258800, 1453262400, 1453266000, 1453269600, 1453273200, 
    1453276800, 1453280400, 1453284000, 1453287600, 1453291200, 1453294800, 
    1453298400, 1453302000, 1453305600, 1453309200, 1453312800, 1453316400, 
    1453320000, 1453323600, 1453327200, 1453330800, 1453334400, 1453338000, 
    1453341600, 1453345200, 1453348800, 1453352400, 1453356000, 1453359600, 
    1453363200, 1453366800, 1453370400, 1453374000, 1453377600, 1453381200, 
    1453384800, 1453388400, 1453392000, 1453395600, 1453399200, 1453402800, 
    1453406400, 1453410000, 1453413600, 1453417200, 1453420800, 1453424400, 
    1453428000, 1453431600, 1453435200, 1453438800, 1453442400, 1453446000, 
    1453449600, 1453453200, 1453456800, 1453460400, 1453464000, 1453467600, 
    1453471200, 1453474800, 1453478400, 1453482000, 1453485600, 1453489200, 
    1453492800, 1453496400, 1453500000, 1453503600, 1453507200, 1453510800, 
    1453514400, 1453518000, 1453521600, 1453525200, 1453528800, 1453532400, 
    1453536000, 1453539600, 1453543200, 1453546800, 1453550400, 1453554000, 
    1453557600, 1453561200, 1453564800, 1453568400, 1453572000, 1453575600, 
    1453579200, 1453582800, 1453586400, 1453590000, 1453593600, 1453597200, 
    1453600800, 1453604400, 1453608000, 1453611600, 1453615200, 1453618800, 
    1453622400, 1453626000, 1453629600, 1453633200, 1453636800, 1453640400, 
    1453644000, 1453647600, 1453651200, 1453654800, 1453658400, 1453662000, 
    1453665600, 1453669200, 1453672800, 1453676400, 1453680000, 1453683600, 
    1453687200, 1453690800, 1453694400, 1453698000, 1453701600, 1453705200, 
    1453708800, 1453712400, 1453716000, 1453719600, 1453723200, 1453726800, 
    1453730400, 1453734000, 1453737600, 1453741200, 1453744800, 1453748400, 
    1453752000, 1453755600, 1453759200, 1453762800, 1453766400, 1453770000, 
    1453773600, 1453777200, 1453780800, 1453784400, 1453788000, 1453791600, 
    1453795200, 1453798800, 1453802400, 1453806000, 1453809600, 1453813200, 
    1453816800, 1453820400, 1453824000, 1453827600, 1453831200, 1453834800, 
    1453838400, 1453842000, 1453845600, 1453849200, 1453852800, 1453856400, 
    1453860000, 1453863600, 1453867200, 1453870800, 1453874400, 1453878000, 
    1453881600, 1453885200, 1453888800, 1453892400, 1453896000, 1453899600, 
    1453903200, 1453906800, 1453910400, 1453914000, 1453917600, 1453921200, 
    1453924800, 1453928400, 1453932000, 1453935600, 1453939200, 1453942800, 
    1453946400, 1453950000, 1453953600, 1453957200, 1453960800, 1453964400, 
    1453968000, 1453971600, 1453975200, 1453978800, 1453982400, 1453986000, 
    1453989600, 1453993200, 1453996800, 1454000400, 1454004000, 1454007600, 
    1454011200, 1454014800, 1454018400, 1454022000, 1454025600, 1454029200, 
    1454032800, 1454036400, 1454040000, 1454043600, 1454047200, 1454050800, 
    1454054400, 1454058000, 1454061600, 1454065200, 1454068800, 1454072400, 
    1454076000, 1454079600, 1454083200, 1454086800, 1454090400, 1454094000, 
    1454097600, 1454101200, 1454104800, 1454108400, 1454112000, 1454115600, 
    1454119200, 1454122800, 1454126400, 1454130000, 1454133600, 1454137200, 
    1454140800, 1454144400, 1454148000, 1454151600, 1454155200, 1454158800, 
    1454162400, 1454166000, 1454169600, 1454173200, 1454176800, 1454180400, 
    1454184000, 1454187600, 1454191200, 1454194800, 1454198400, 1454202000, 
    1454205600, 1454209200, 1454212800, 1454216400, 1454220000, 1454223600, 
    1454227200, 1454230800, 1454234400, 1454238000, 1454241600, 1454245200, 
    1454248800, 1454252400, 1454256000, 1454259600, 1454263200, 1454266800, 
    1454270400, 1454274000, 1454277600, 1454281200, 1454284800, 1454288400, 
    1454292000, 1454295600, 1454299200, 1454302800, 1454306400, 1454310000, 
    1454313600, 1454317200, 1454320800, 1454324400, 1454328000, 1454331600, 
    1454335200, 1454338800, 1454342400, 1454346000, 1454349600, 1454353200, 
    1454356800, 1454360400, 1454364000, 1454367600, 1454371200, 1454374800, 
    1454378400, 1454382000, 1454385600, 1454389200, 1454392800, 1454396400, 
    1454400000, 1454403600, 1454407200, 1454410800, 1454414400, 1454418000, 
    1454421600, 1454425200, 1454428800, 1454432400, 1454436000, 1454439600, 
    1454443200, 1454446800, 1454450400, 1454454000, 1454457600, 1454461200, 
    1454464800, 1454468400, 1454472000, 1454475600, 1454479200, 1454482800, 
    1454486400, 1454490000, 1454493600, 1454497200, 1454500800, 1454504400, 
    1454508000, 1454511600, 1454515200, 1454518800, 1454522400, 1454526000, 
    1454529600, 1454533200, 1454536800, 1454540400, 1454544000, 1454547600, 
    1454551200, 1454554800, 1454558400, 1454562000, 1454565600, 1454569200, 
    1454572800, 1454576400, 1454580000, 1454583600, 1454587200, 1454590800, 
    1454594400, 1454598000, 1454601600, 1454605200, 1454608800, 1454612400, 
    1454616000, 1454619600, 1454623200, 1454626800, 1454630400, 1454634000, 
    1454637600, 1454641200, 1454644800, 1454648400, 1454652000, 1454655600, 
    1454659200, 1454662800, 1454666400, 1454670000, 1454673600, 1454677200, 
    1454680800, 1454684400, 1454688000, 1454691600, 1454695200, 1454698800, 
    1454702400, 1454706000, 1454709600, 1454713200, 1454716800, 1454720400, 
    1454724000, 1454727600, 1454731200, 1454734800, 1454738400, 1454742000, 
    1454745600, 1454749200, 1454752800, 1454756400, 1454760000, 1454763600, 
    1454767200, 1454770800, 1454774400, 1454778000, 1454781600, 1454785200, 
    1454788800, 1454792400, 1454796000, 1454799600, 1454803200, 1454806800, 
    1454810400, 1454814000, 1454817600, 1454821200, 1454824800, 1454828400, 
    1454832000, 1454835600, 1454839200, 1454842800, 1454846400, 1454850000, 
    1454853600, 1454857200, 1454860800, 1454864400, 1454868000, 1454871600, 
    1454875200, 1454878800, 1454882400, 1454886000, 1454889600, 1454893200, 
    1454896800, 1454900400, 1454904000, 1454907600, 1454911200, 1454914800, 
    1454918400, 1454922000, 1454925600, 1454929200, 1454932800, 1454936400, 
    1454940000, 1454943600, 1454947200, 1454950800, 1454954400, 1454958000, 
    1454961600, 1454965200, 1454968800, 1454972400, 1454976000, 1454979600, 
    1454983200, 1454986800, 1454990400, 1454994000, 1454997600, 1455001200, 
    1455004800, 1455008400, 1455012000, 1455015600, 1455019200, 1455022800, 
    1455026400, 1455030000, 1455033600, 1455037200, 1455040800, 1455044400, 
    1455048000, 1455051600, 1455055200, 1455058800, 1455062400, 1455066000, 
    1455069600, 1455073200, 1455076800, 1455080400, 1455084000, 1455087600, 
    1455091200, 1455094800, 1455098400, 1455102000, 1455105600, 1455109200, 
    1455112800, 1455116400, 1455120000, 1455123600, 1455127200, 1455130800, 
    1455134400, 1455138000, 1455141600, 1455145200, 1455148800, 1455152400, 
    1455156000, 1455159600, 1455163200, 1455166800, 1455170400, 1455174000, 
    1455177600, 1455181200, 1455184800, 1455188400, 1455192000, 1455195600, 
    1455199200, 1455202800, 1455206400, 1455210000, 1455213600, 1455217200, 
    1455220800, 1455224400, 1455228000, 1455231600, 1455235200, 1455238800, 
    1455242400, 1455246000, 1455249600, 1455253200, 1455256800, 1455260400, 
    1455264000, 1455267600, 1455271200, 1455274800, 1455278400, 1455282000, 
    1455285600, 1455289200, 1455292800, 1455296400, 1455300000, 1455303600, 
    1455307200, 1455310800, 1455314400, 1455318000, 1455321600, 1455325200, 
    1455328800, 1455332400, 1455336000, 1455339600, 1455343200, 1455346800, 
    1455350400, 1455354000, 1455357600, 1455361200, 1455364800, 1455368400, 
    1455372000, 1455375600, 1455379200, 1455382800, 1455386400, 1455390000, 
    1455393600, 1455397200, 1455400800, 1455404400, 1455408000, 1455411600, 
    1455415200, 1455418800, 1455422400, 1455426000, 1455429600, 1455433200, 
    1455436800, 1455440400, 1455444000, 1455447600, 1455451200, 1455454800, 
    1455458400, 1455462000, 1455465600, 1455469200, 1455472800, 1455476400, 
    1455480000, 1455483600, 1455487200, 1455490800, 1455494400, 1455498000, 
    1455501600, 1455505200, 1455508800, 1455512400, 1455516000, 1455519600, 
    1455523200, 1455526800, 1455530400, 1455534000, 1455537600, 1455541200, 
    1455544800, 1455548400, 1455552000, 1455555600, 1455559200, 1455562800, 
    1455566400, 1455570000, 1455573600, 1455577200, 1455580800, 1455584400, 
    1455588000, 1455591600, 1455595200, 1455598800, 1455602400, 1455606000, 
    1455609600, 1455613200, 1455616800, 1455620400, 1455624000, 1455627600, 
    1455631200, 1455634800, 1455638400, 1455642000, 1455645600, 1455649200, 
    1455652800, 1455656400, 1455660000, 1455663600, 1455667200, 1455670800, 
    1455674400, 1455678000, 1455681600, 1455685200, 1455688800, 1455692400, 
    1455696000, 1455699600, 1455703200, 1455706800, 1455710400, 1455714000, 
    1455717600, 1455721200, 1455724800, 1455728400, 1455732000, 1455735600, 
    1455739200, 1455742800, 1455746400, 1455750000, 1455753600, 1455757200, 
    1455760800, 1455764400, 1455768000, 1455771600, 1455775200, 1455778800, 
    1455782400, 1455786000, 1455789600, 1455793200, 1455796800, 1455800400, 
    1455804000, 1455807600, 1455811200, 1455814800, 1455818400, 1455822000, 
    1455825600, 1455829200, 1455832800, 1455836400, 1455840000, 1455843600, 
    1455847200, 1455850800, 1455854400, 1455858000, 1455861600, 1455865200, 
    1455868800, 1455872400, 1455876000, 1455879600, 1455883200, 1455886800, 
    1455890400, 1455894000, 1455897600, 1455901200, 1455904800, 1455908400, 
    1455912000, 1455915600, 1455919200, 1455922800, 1455926400, 1455930000, 
    1455933600, 1455937200, 1455940800, 1455944400, 1455948000, 1455951600, 
    1455955200, 1455958800, 1455962400, 1455966000, 1455969600, 1455973200, 
    1455976800, 1455980400, 1455984000, 1455987600, 1455991200, 1455994800, 
    1455998400, 1456002000, 1456005600, 1456009200, 1456012800, 1456016400, 
    1456020000, 1456023600, 1456027200, 1456030800, 1456034400, 1456038000, 
    1456041600, 1456045200, 1456048800, 1456052400, 1456056000, 1456059600, 
    1456063200, 1456066800, 1456070400, 1456074000, 1456077600, 1456081200, 
    1456084800, 1456088400, 1456092000, 1456095600, 1456099200, 1456102800, 
    1456106400, 1456110000, 1456113600, 1456117200, 1456120800, 1456124400, 
    1456128000, 1456131600, 1456135200, 1456138800, 1456142400, 1456146000, 
    1456149600, 1456153200, 1456156800, 1456160400, 1456164000, 1456167600, 
    1456171200, 1456174800, 1456178400, 1456182000, 1456185600, 1456189200, 
    1456192800, 1456196400, 1456200000, 1456203600, 1456207200, 1456210800, 
    1456214400, 1456218000, 1456221600, 1456225200, 1456228800, 1456232400, 
    1456236000, 1456239600, 1456243200, 1456246800, 1456250400, 1456254000, 
    1456257600, 1456261200, 1456264800, 1456268400, 1456272000, 1456275600, 
    1456279200, 1456282800, 1456286400, 1456290000, 1456293600, 1456297200, 
    1456300800, 1456304400, 1456308000, 1456311600, 1456315200, 1456318800, 
    1456322400, 1456326000, 1456329600, 1456333200, 1456336800, 1456340400, 
    1456344000, 1456347600, 1456351200, 1456354800, 1456358400, 1456362000, 
    1456365600, 1456369200, 1456372800, 1456376400, 1456380000, 1456383600, 
    1456387200, 1456390800, 1456394400, 1456398000, 1456401600, 1456405200, 
    1456408800, 1456412400, 1456416000, 1456419600, 1456423200, 1456426800, 
    1456430400, 1456434000, 1456437600, 1456441200, 1456444800, 1456448400, 
    1456452000, 1456455600, 1456459200, 1456462800, 1456466400, 1456470000, 
    1456473600, 1456477200, 1456480800, 1456484400, 1456488000, 1456491600, 
    1456495200, 1456498800, 1456502400, 1456506000, 1456509600, 1456513200, 
    1456516800, 1456520400, 1456524000, 1456527600, 1456531200, 1456534800, 
    1456538400, 1456542000, 1456545600, 1456549200, 1456552800, 1456556400, 
    1456560000, 1456563600, 1456567200, 1456570800, 1456574400, 1456578000, 
    1456581600, 1456585200, 1456588800, 1456592400, 1456596000, 1456599600, 
    1456603200, 1456606800, 1456610400, 1456614000, 1456617600, 1456621200, 
    1456624800, 1456628400, 1456632000, 1456635600, 1456639200, 1456642800, 
    1456646400, 1456650000, 1456653600, 1456657200, 1456660800, 1456664400, 
    1456668000, 1456671600, 1456675200, 1456678800, 1456682400, 1456686000, 
    1456689600, 1456693200, 1456696800, 1456700400, 1456704000, 1456707600, 
    1456711200, 1456714800, 1456718400, 1456722000, 1456725600, 1456729200, 
    1456732800, 1456736400, 1456740000, 1456743600, 1456747200, 1456750800, 
    1456754400, 1456758000, 1456761600, 1456765200, 1456768800, 1456772400, 
    1456776000, 1456779600, 1456783200, 1456786800, 1456790400, 1456794000, 
    1456797600, 1456801200, 1456804800, 1456808400, 1456812000, 1456815600, 
    1456819200, 1456822800, 1456826400, 1456830000, 1456833600, 1456837200, 
    1456840800, 1456844400, 1456848000, 1456851600, 1456855200, 1456858800, 
    1456862400, 1456866000, 1456869600, 1456873200, 1456876800, 1456880400, 
    1456884000, 1456887600, 1456891200, 1456894800, 1456898400, 1456902000, 
    1456905600, 1456909200, 1456912800, 1456916400, 1456920000, 1456923600, 
    1456927200, 1456930800, 1456934400, 1456938000, 1456941600, 1456945200, 
    1456948800, 1456952400, 1456956000, 1456959600, 1456963200, 1456966800, 
    1456970400, 1456974000, 1456977600, 1456981200, 1456984800, 1456988400, 
    1456992000, 1456995600, 1456999200, 1457002800, 1457006400, 1457010000, 
    1457013600, 1457017200, 1457020800, 1457024400, 1457028000, 1457031600, 
    1457035200, 1457038800, 1457042400, 1457046000, 1457049600, 1457053200, 
    1457056800, 1457060400, 1457064000, 1457067600, 1457071200, 1457074800, 
    1457078400, 1457082000, 1457085600, 1457089200, 1457092800, 1457096400, 
    1457100000, 1457103600, 1457107200, 1457110800, 1457114400, 1457118000, 
    1457121600, 1457125200, 1457128800, 1457132400, 1457136000, 1457139600, 
    1457143200, 1457146800, 1457150400, 1457154000, 1457157600, 1457161200, 
    1457164800, 1457168400, 1457172000, 1457175600, 1457179200, 1457182800, 
    1457186400, 1457190000, 1457193600, 1457197200, 1457200800, 1457204400, 
    1457208000, 1457211600, 1457215200, 1457218800, 1457222400, 1457226000, 
    1457229600, 1457233200, 1457236800, 1457240400, 1457244000, 1457247600, 
    1457251200, 1457254800, 1457258400, 1457262000, 1457265600, 1457269200, 
    1457272800, 1457276400, 1457280000, 1457283600, 1457287200, 1457290800, 
    1457294400, 1457298000, 1457301600, 1457305200, 1457308800, 1457312400, 
    1457316000, 1457319600, 1457323200, 1457326800, 1457330400, 1457334000, 
    1457337600, 1457341200, 1457344800, 1457348400, 1457352000, 1457355600, 
    1457359200, 1457362800, 1457366400, 1457370000, 1457373600, 1457377200, 
    1457380800, 1457384400, 1457388000, 1457391600, 1457395200, 1457398800, 
    1457402400, 1457406000, 1457409600, 1457413200, 1457416800, 1457420400, 
    1457424000, 1457427600, 1457431200, 1457434800, 1457438400, 1457442000, 
    1457445600, 1457449200, 1457452800, 1457456400, 1457460000, 1457463600, 
    1457467200, 1457470800, 1457474400, 1457478000, 1457481600, 1457485200, 
    1457488800, 1457492400, 1457496000, 1457499600, 1457503200, 1457506800, 
    1457510400, 1457514000, 1457517600, 1457521200, 1457524800, 1457528400, 
    1457532000, 1457535600, 1457539200, 1457542800, 1457546400, 1457550000, 
    1457553600, 1457557200, 1457560800, 1457564400, 1457568000, 1457571600, 
    1457575200, 1457578800, 1457582400, 1457586000, 1457589600, 1457593200, 
    1457596800, 1457600400, 1457604000, 1457607600, 1457611200, 1457614800, 
    1457618400, 1457622000, 1457625600, 1457629200, 1457632800, 1457636400, 
    1457640000, 1457643600, 1457647200, 1457650800, 1457654400, 1457658000, 
    1457661600, 1457665200, 1457668800, 1457672400, 1457676000, 1457679600, 
    1457683200, 1457686800, 1457690400, 1457694000, 1457697600, 1457701200, 
    1457704800, 1457708400, 1457712000, 1457715600, 1457719200, 1457722800, 
    1457726400, 1457730000, 1457733600, 1457737200, 1457740800, 1457744400, 
    1457748000, 1457751600, 1457755200, 1457758800, 1457762400, 1457766000, 
    1457769600, 1457773200, 1457776800, 1457780400, 1457784000, 1457787600, 
    1457791200, 1457794800, 1457798400, 1457802000, 1457805600, 1457809200, 
    1457812800, 1457816400, 1457820000, 1457823600, 1457827200, 1457830800, 
    1457834400, 1457838000, 1457841600, 1457845200, 1457848800, 1457852400, 
    1457856000, 1457859600, 1457863200, 1457866800, 1457870400, 1457874000, 
    1457877600, 1457881200, 1457884800, 1457888400, 1457892000, 1457895600, 
    1457899200, 1457902800, 1457906400, 1457910000, 1457913600, 1457917200, 
    1457920800, 1457924400, 1457928000, 1457931600, 1457935200, 1457938800, 
    1457942400, 1457946000, 1457949600, 1457953200, 1457956800, 1457960400, 
    1457964000, 1457967600, 1457971200, 1457974800, 1457978400, 1457982000, 
    1457985600, 1457989200, 1457992800, 1457996400, 1458000000, 1458003600, 
    1458007200, 1458010800, 1458014400, 1458018000, 1458021600, 1458025200, 
    1458028800, 1458032400, 1458036000, 1458039600, 1458043200, 1458046800, 
    1458050400, 1458054000, 1458057600, 1458061200, 1458064800, 1458068400, 
    1458072000, 1458075600, 1458079200, 1458082800, 1458086400, 1458090000, 
    1458093600, 1458097200, 1458100800, 1458104400, 1458108000, 1458111600, 
    1458115200, 1458118800, 1458122400, 1458126000, 1458129600, 1458133200, 
    1458136800, 1458140400, 1458144000, 1458147600, 1458151200, 1458154800, 
    1458158400, 1458162000, 1458165600, 1458169200, 1458172800, 1458176400, 
    1458180000, 1458183600, 1458187200, 1458190800, 1458194400, 1458198000, 
    1458201600, 1458205200, 1458208800, 1458212400, 1458216000, 1458219600, 
    1458223200, 1458226800, 1458230400, 1458234000, 1458237600, 1458241200, 
    1458244800, 1458248400, 1458252000, 1458255600, 1458259200, 1458262800, 
    1458266400, 1458270000, 1458273600, 1458277200, 1458280800, 1458284400, 
    1458288000, 1458291600, 1458295200, 1458298800, 1458302400, 1458306000, 
    1458309600, 1458313200, 1458316800, 1458320400, 1458324000, 1458327600, 
    1458331200, 1458334800, 1458338400, 1458342000, 1458345600, 1458349200, 
    1458352800, 1458356400, 1458360000, 1458363600, 1458367200, 1458370800, 
    1458374400, 1458378000, 1458381600, 1458385200, 1458388800, 1458392400, 
    1458396000, 1458399600, 1458403200, 1458406800, 1458410400, 1458414000, 
    1458417600, 1458421200, 1458424800, 1458428400, 1458432000, 1458435600, 
    1458439200, 1458442800, 1458446400, 1458450000, 1458453600, 1458457200, 
    1458460800, 1458464400, 1458468000, 1458471600, 1458475200, 1458478800, 
    1458482400, 1458486000, 1458489600, 1458493200, 1458496800, 1458500400, 
    1458504000, 1458507600, 1458511200, 1458514800, 1458518400, 1458522000, 
    1458525600, 1458529200, 1458532800, 1458536400, 1458540000, 1458543600, 
    1458547200, 1458550800, 1458554400, 1458558000, 1458561600, 1458565200, 
    1458568800, 1458572400, 1458576000, 1458579600, 1458583200, 1458586800, 
    1458590400, 1458594000, 1458597600, 1458601200, 1458604800, 1458608400, 
    1458612000, 1458615600, 1458619200, 1458622800, 1458626400, 1458630000, 
    1458633600, 1458637200, 1458640800, 1458644400, 1458648000, 1458651600, 
    1458655200, 1458658800, 1458662400, 1458666000, 1458669600, 1458673200, 
    1458676800, 1458680400, 1458684000, 1458687600, 1458691200, 1458694800, 
    1458698400, 1458702000, 1458705600, 1458709200, 1458712800, 1458716400, 
    1458720000, 1458723600, 1458727200, 1458730800, 1458734400, 1458738000, 
    1458741600, 1458745200, 1458748800, 1458752400, 1458756000, 1458759600, 
    1458763200, 1458766800, 1458770400, 1458774000, 1458777600, 1458781200, 
    1458784800, 1458788400, 1458792000, 1458795600, 1458799200, 1458802800, 
    1458806400, 1458810000, 1458813600, 1458817200, 1458820800, 1458824400, 
    1458828000, 1458831600, 1458835200, 1458838800, 1458842400, 1458846000, 
    1458849600, 1458853200, 1458856800, 1458860400, 1458864000, 1458867600, 
    1458871200, 1458874800, 1458878400, 1458882000, 1458885600, 1458889200, 
    1458892800, 1458896400, 1458900000, 1458903600, 1458907200, 1458910800, 
    1458914400, 1458918000, 1458921600, 1458925200, 1458928800, 1458932400, 
    1458936000, 1458939600, 1458943200, 1458946800, 1458950400, 1458954000, 
    1458957600, 1458961200, 1458964800, 1458968400, 1458972000, 1458975600, 
    1458979200, 1458982800, 1458986400, 1458990000, 1458993600, 1458997200, 
    1459000800, 1459004400, 1459008000, 1459011600, 1459015200, 1459018800, 
    1459022400, 1459026000, 1459029600, 1459033200, 1459036800, 1459040400, 
    1459044000, 1459047600, 1459051200, 1459054800, 1459058400, 1459062000, 
    1459065600, 1459069200, 1459072800, 1459076400, 1459080000, 1459083600, 
    1459087200, 1459090800, 1459094400, 1459098000, 1459101600, 1459105200, 
    1459108800, 1459112400, 1459116000, 1459119600, 1459123200, 1459126800, 
    1459130400, 1459134000, 1459137600, 1459141200, 1459144800, 1459148400, 
    1459152000, 1459155600, 1459159200, 1459162800, 1459166400, 1459170000, 
    1459173600, 1459177200, 1459180800, 1459184400, 1459188000, 1459191600, 
    1459195200, 1459198800, 1459202400, 1459206000, 1459209600, 1459213200, 
    1459216800, 1459220400, 1459224000, 1459227600, 1459231200, 1459234800, 
    1459238400, 1459242000, 1459245600, 1459249200, 1459252800, 1459256400, 
    1459260000, 1459263600, 1459267200, 1459270800, 1459274400, 1459278000, 
    1459281600, 1459285200, 1459288800, 1459292400, 1459296000, 1459299600, 
    1459303200, 1459306800, 1459310400, 1459314000, 1459317600, 1459321200, 
    1459324800, 1459328400, 1459332000, 1459335600, 1459339200, 1459342800, 
    1459346400, 1459350000, 1459353600, 1459357200, 1459360800, 1459364400, 
    1459368000, 1459371600, 1459375200, 1459378800, 1459382400, 1459386000, 
    1459389600, 1459393200, 1459396800, 1459400400, 1459404000, 1459407600, 
    1459411200, 1459414800, 1459418400, 1459422000, 1459425600, 1459429200, 
    1459432800, 1459436400, 1459440000, 1459443600, 1459447200, 1459450800, 
    1459454400, 1459458000, 1459461600, 1459465200, 1459468800, 1459472400, 
    1459476000, 1459479600, 1459483200, 1459486800, 1459490400, 1459494000, 
    1459497600, 1459501200, 1459504800, 1459508400, 1459512000, 1459515600, 
    1459519200, 1459522800, 1459526400, 1459530000, 1459533600, 1459537200, 
    1459540800, 1459544400, 1459548000, 1459551600, 1459555200, 1459558800, 
    1459562400, 1459566000, 1459569600, 1459573200, 1459576800, 1459580400, 
    1459584000, 1459587600, 1459591200, 1459594800, 1459598400, 1459602000, 
    1459605600, 1459609200, 1459612800, 1459616400, 1459620000, 1459623600, 
    1459627200, 1459630800, 1459634400, 1459638000, 1459641600, 1459645200, 
    1459648800, 1459652400, 1459656000, 1459659600, 1459663200, 1459666800, 
    1459670400, 1459674000, 1459677600, 1459681200, 1459684800, 1459688400, 
    1459692000, 1459695600, 1459699200, 1459702800, 1459706400, 1459710000, 
    1459713600, 1459717200, 1459720800, 1459724400, 1459728000, 1459731600, 
    1459735200, 1459738800, 1459742400, 1459746000, 1459749600, 1459753200, 
    1459756800, 1459760400, 1459764000, 1459767600, 1459771200, 1459774800, 
    1459778400, 1459782000, 1459785600, 1459789200, 1459792800, 1459796400, 
    1459800000, 1459803600, 1459807200, 1459810800, 1459814400, 1459818000, 
    1459821600, 1459825200, 1459828800, 1459832400, 1459836000, 1459839600, 
    1459843200, 1459846800, 1459850400, 1459854000, 1459857600, 1459861200, 
    1459864800, 1459868400, 1459872000, 1459875600, 1459879200, 1459882800, 
    1459886400, 1459890000, 1459893600, 1459897200, 1459900800, 1459904400, 
    1459908000, 1459911600, 1459915200, 1459918800, 1459922400, 1459926000, 
    1459929600, 1459933200, 1459936800, 1459940400, 1459944000, 1459947600, 
    1459951200, 1459954800, 1459958400, 1459962000, 1459965600, 1459969200, 
    1459972800, 1459976400, 1459980000, 1459983600, 1459987200, 1459990800, 
    1459994400, 1459998000, 1460001600, 1460005200, 1460008800, 1460012400, 
    1460016000, 1460019600, 1460023200, 1460026800, 1460030400, 1460034000, 
    1460037600, 1460041200, 1460044800, 1460048400, 1460052000, 1460055600, 
    1460059200, 1460062800, 1460066400, 1460070000, 1460073600, 1460077200, 
    1460080800, 1460084400, 1460088000, 1460091600, 1460095200, 1460098800, 
    1460102400, 1460106000, 1460109600, 1460113200, 1460116800, 1460120400, 
    1460124000, 1460127600, 1460131200, 1460134800, 1460138400, 1460142000, 
    1460145600, 1460149200, 1460152800, 1460156400, 1460160000, 1460163600, 
    1460167200, 1460170800, 1460174400, 1460178000, 1460181600, 1460185200, 
    1460188800, 1460192400, 1460196000, 1460199600, 1460203200, 1460206800, 
    1460210400, 1460214000, 1460217600, 1460221200, 1460224800, 1460228400, 
    1460232000, 1460235600, 1460239200, 1460242800, 1460246400, 1460250000, 
    1460253600, 1460257200, 1460260800, 1460264400, 1460268000, 1460271600, 
    1460275200, 1460278800, 1460282400, 1460286000, 1460289600, 1460293200, 
    1460296800, 1460300400, 1460304000, 1460307600, 1460311200, 1460314800, 
    1460318400, 1460322000, 1460325600, 1460329200, 1460332800, 1460336400, 
    1460340000, 1460343600, 1460347200, 1460350800, 1460354400, 1460358000, 
    1460361600, 1460365200, 1460368800, 1460372400, 1460376000, 1460379600, 
    1460383200, 1460386800, 1460390400, 1460394000, 1460397600, 1460401200, 
    1460404800, 1460408400, 1460412000, 1460415600, 1460419200, 1460422800, 
    1460426400, 1460430000, 1460433600, 1460437200, 1460440800, 1460444400, 
    1460448000, 1460451600, 1460455200, 1460458800, 1460462400, 1460466000, 
    1460469600, 1460473200, 1460476800, 1460480400, 1460484000, 1460487600, 
    1460491200, 1460494800, 1460498400, 1460502000, 1460505600, 1460509200, 
    1460512800, 1460516400, 1460520000, 1460523600, 1460527200, 1460530800, 
    1460534400, 1460538000, 1460541600, 1460545200, 1460548800, 1460552400, 
    1460556000, 1460559600, 1460563200, 1460566800, 1460570400, 1460574000, 
    1460577600, 1460581200, 1460584800, 1460588400, 1460592000, 1460595600, 
    1460599200, 1460602800, 1460606400, 1460610000, 1460613600, 1460617200, 
    1460620800, 1460624400, 1460628000, 1460631600, 1460635200, 1460638800, 
    1460642400, 1460646000, 1460649600, 1460653200, 1460656800, 1460660400, 
    1460664000, 1460667600, 1460671200, 1460674800, 1460678400, 1460682000, 
    1460685600, 1460689200, 1460692800, 1460696400, 1460700000, 1460703600, 
    1460707200, 1460710800, 1460714400, 1460718000, 1460721600, 1460725200, 
    1460728800, 1460732400, 1460736000, 1460739600, 1460743200, 1460746800, 
    1460750400, 1460754000, 1460757600, 1460761200, 1460764800, 1460768400, 
    1460772000, 1460775600, 1460779200, 1460782800, 1460786400, 1460790000, 
    1460793600, 1460797200, 1460800800, 1460804400, 1460808000, 1460811600, 
    1460815200, 1460818800, 1460822400, 1460826000, 1460829600, 1460833200, 
    1460836800, 1460840400, 1460844000, 1460847600, 1460851200, 1460854800, 
    1460858400, 1460862000, 1460865600, 1460869200, 1460872800, 1460876400, 
    1460880000, 1460883600, 1460887200, 1460890800, 1460894400, 1460898000, 
    1460901600, 1460905200, 1460908800, 1460912400, 1460916000, 1460919600, 
    1460923200, 1460926800, 1460930400, 1460934000, 1460937600, 1460941200, 
    1460944800, 1460948400, 1460952000, 1460955600, 1460959200, 1460962800, 
    1460966400, 1460970000, 1460973600, 1460977200, 1460980800, 1460984400, 
    1460988000, 1460991600, 1460995200, 1460998800, 1461002400, 1461006000, 
    1461009600, 1461013200, 1461016800, 1461020400, 1461024000, 1461027600, 
    1461031200, 1461034800, 1461038400, 1461042000, 1461045600, 1461049200, 
    1461052800, 1461056400, 1461060000, 1461063600, 1461067200, 1461070800, 
    1461074400, 1461078000, 1461081600, 1461085200, 1461088800, 1461092400, 
    1461096000, 1461099600, 1461103200, 1461106800, 1461110400, 1461114000, 
    1461117600, 1461121200, 1461124800, 1461128400, 1461132000, 1461135600, 
    1461139200, 1461142800, 1461146400, 1461150000, 1461153600, 1461157200, 
    1461160800, 1461164400, 1461168000, 1461171600, 1461175200, 1461178800, 
    1461182400, 1461186000, 1461189600, 1461193200, 1461196800, 1461200400, 
    1461204000, 1461207600, 1461211200, 1461214800, 1461218400, 1461222000, 
    1461225600, 1461229200, 1461232800, 1461236400, 1461240000, 1461243600, 
    1461247200, 1461250800, 1461254400, 1461258000, 1461261600, 1461265200, 
    1461268800, 1461272400, 1461276000, 1461279600, 1461283200, 1461286800, 
    1461290400, 1461294000, 1461297600, 1461301200, 1461304800, 1461308400, 
    1461312000, 1461315600, 1461319200, 1461322800, 1461326400, 1461330000, 
    1461333600, 1461337200, 1461340800, 1461344400, 1461348000, 1461351600, 
    1461355200, 1461358800, 1461362400, 1461366000, 1461369600, 1461373200, 
    1461376800, 1461380400, 1461384000, 1461387600, 1461391200, 1461394800, 
    1461398400, 1461402000, 1461405600, 1461409200, 1461412800, 1461416400, 
    1461420000, 1461423600, 1461427200, 1461430800, 1461434400, 1461438000, 
    1461441600, 1461445200, 1461448800, 1461452400, 1461456000, 1461459600, 
    1461463200, 1461466800, 1461470400, 1461474000, 1461477600, 1461481200, 
    1461484800, 1461488400, 1461492000, 1461495600, 1461499200, 1461502800, 
    1461506400, 1461510000, 1461513600, 1461517200, 1461520800, 1461524400, 
    1461528000, 1461531600, 1461535200, 1461538800, 1461542400, 1461546000, 
    1461549600, 1461553200, 1461556800, 1461560400, 1461564000, 1461567600, 
    1461571200, 1461574800, 1461578400, 1461582000, 1461585600, 1461589200, 
    1461592800, 1461596400, 1461600000, 1461603600, 1461607200, 1461610800, 
    1461614400, 1461618000, 1461621600, 1461625200, 1461628800, 1461632400, 
    1461636000, 1461639600, 1461643200, 1461646800, 1461650400, 1461654000, 
    1461657600, 1461661200, 1461664800, 1461668400, 1461672000, 1461675600, 
    1461679200, 1461682800, 1461686400, 1461690000, 1461693600, 1461697200, 
    1461700800, 1461704400, 1461708000, 1461711600, 1461715200, 1461718800, 
    1461722400, 1461726000, 1461729600, 1461733200, 1461736800, 1461740400, 
    1461744000, 1461747600, 1461751200, 1461754800, 1461758400, 1461762000, 
    1461765600, 1461769200, 1461772800, 1461776400, 1461780000, 1461783600, 
    1461787200, 1461790800, 1461794400, 1461798000, 1461801600, 1461805200, 
    1461808800, 1461812400, 1461816000, 1461819600, 1461823200, 1461826800, 
    1461830400, 1461834000, 1461837600, 1461841200, 1461844800, 1461848400, 
    1461852000, 1461855600, 1461859200, 1461862800, 1461866400, 1461870000, 
    1461873600, 1461877200, 1461880800, 1461884400, 1461888000, 1461891600, 
    1461895200, 1461898800, 1461902400, 1461906000, 1461909600, 1461913200, 
    1461916800, 1461920400, 1461924000, 1461927600, 1461931200, 1461934800, 
    1461938400, 1461942000, 1461945600, 1461949200, 1461952800, 1461956400, 
    1461960000, 1461963600, 1461967200, 1461970800, 1461974400, 1461978000, 
    1461981600, 1461985200, 1461988800, 1461992400, 1461996000, 1461999600, 
    1462003200, 1462006800, 1462010400, 1462014000, 1462017600, 1462021200, 
    1462024800, 1462028400, 1462032000, 1462035600, 1462039200, 1462042800, 
    1462046400, 1462050000, 1462053600, 1462057200, 1462060800, 1462064400, 
    1462068000, 1462071600, 1462075200, 1462078800, 1462082400, 1462086000, 
    1462089600, 1462093200, 1462096800, 1462100400, 1462104000, 1462107600, 
    1462111200, 1462114800, 1462118400, 1462122000, 1462125600, 1462129200, 
    1462132800, 1462136400, 1462140000, 1462143600, 1462147200, 1462150800, 
    1462154400, 1462158000, 1462161600, 1462165200, 1462168800, 1462172400, 
    1462176000, 1462179600, 1462183200, 1462186800, 1462190400, 1462194000, 
    1462197600, 1462201200, 1462204800, 1462208400, 1462212000, 1462215600, 
    1462219200, 1462222800, 1462226400, 1462230000, 1462233600, 1462237200, 
    1462240800, 1462244400, 1462248000, 1462251600, 1462255200, 1462258800, 
    1462262400, 1462266000, 1462269600, 1462273200, 1462276800, 1462280400, 
    1462284000, 1462287600, 1462291200, 1462294800, 1462298400, 1462302000, 
    1462305600, 1462309200, 1462312800, 1462316400, 1462320000, 1462323600, 
    1462327200, 1462330800, 1462334400, 1462338000, 1462341600, 1462345200, 
    1462348800, 1462352400, 1462356000, 1462359600, 1462363200, 1462366800, 
    1462370400, 1462374000, 1462377600, 1462381200, 1462384800, 1462388400, 
    1462392000, 1462395600, 1462399200, 1462402800, 1462406400, 1462410000, 
    1462413600, 1462417200, 1462420800, 1462424400, 1462428000, 1462431600, 
    1462435200, 1462438800, 1462442400, 1462446000, 1462449600, 1462453200, 
    1462456800, 1462460400, 1462464000, 1462467600, 1462471200, 1462474800, 
    1462478400, 1462482000, 1462485600, 1462489200, 1462492800, 1462496400, 
    1462500000, 1462503600, 1462507200, 1462510800, 1462514400, 1462518000, 
    1462521600, 1462525200, 1462528800, 1462532400, 1462536000, 1462539600, 
    1462543200, 1462546800, 1462550400, 1462554000, 1462557600, 1462561200, 
    1462564800, 1462568400, 1462572000, 1462575600, 1462579200, 1462582800, 
    1462586400, 1462590000, 1462593600, 1462597200, 1462600800, 1462604400, 
    1462608000, 1462611600, 1462615200, 1462618800, 1462622400, 1462626000, 
    1462629600, 1462633200, 1462636800, 1462640400, 1462644000, 1462647600, 
    1462651200, 1462654800, 1462658400, 1462662000, 1462665600, 1462669200, 
    1462672800, 1462676400, 1462680000, 1462683600, 1462687200, 1462690800, 
    1462694400, 1462698000, 1462701600, 1462705200, 1462708800, 1462712400, 
    1462716000, 1462719600, 1462723200, 1462726800, 1462730400, 1462734000, 
    1462737600, 1462741200, 1462744800, 1462748400, 1462752000, 1462755600, 
    1462759200, 1462762800, 1462766400, 1462770000, 1462773600, 1462777200, 
    1462780800, 1462784400, 1462788000, 1462791600, 1462795200, 1462798800, 
    1462802400, 1462806000, 1462809600, 1462813200, 1462816800, 1462820400, 
    1462824000, 1462827600, 1462831200, 1462834800, 1462838400, 1462842000, 
    1462845600, 1462849200, 1462852800, 1462856400, 1462860000, 1462863600, 
    1462867200, 1462870800, 1462874400, 1462878000, 1462881600, 1462885200, 
    1462888800, 1462892400, 1462896000, 1462899600, 1462903200, 1462906800, 
    1462910400, 1462914000, 1462917600, 1462921200, 1462924800, 1462928400, 
    1462932000, 1462935600, 1462939200, 1462942800, 1462946400, 1462950000, 
    1462953600, 1462957200, 1462960800, 1462964400, 1462968000, 1462971600, 
    1462975200, 1462978800, 1462982400, 1462986000, 1462989600, 1462993200, 
    1462996800, 1463000400, 1463004000, 1463007600, 1463011200, 1463014800, 
    1463018400, 1463022000, 1463025600, 1463029200, 1463032800, 1463036400, 
    1463040000, 1463043600, 1463047200, 1463050800, 1463054400, 1463058000, 
    1463061600, 1463065200, 1463068800, 1463072400, 1463076000, 1463079600, 
    1463083200, 1463086800, 1463090400, 1463094000, 1463097600, 1463101200, 
    1463104800, 1463108400, 1463112000, 1463115600, 1463119200, 1463122800, 
    1463126400, 1463130000, 1463133600, 1463137200, 1463140800, 1463144400, 
    1463148000, 1463151600, 1463155200, 1463158800, 1463162400, 1463166000, 
    1463169600, 1463173200, 1463176800, 1463180400, 1463184000, 1463187600, 
    1463191200, 1463194800, 1463198400, 1463202000, 1463205600, 1463209200, 
    1463212800, 1463216400, 1463220000, 1463223600, 1463227200, 1463230800, 
    1463234400, 1463238000, 1463241600, 1463245200, 1463248800, 1463252400, 
    1463256000, 1463259600, 1463263200, 1463266800, 1463270400, 1463274000, 
    1463277600, 1463281200, 1463284800, 1463288400, 1463292000, 1463295600, 
    1463299200, 1463302800, 1463306400, 1463310000, 1463313600, 1463317200, 
    1463320800, 1463324400, 1463328000, 1463331600, 1463335200, 1463338800, 
    1463342400, 1463346000, 1463349600, 1463353200, 1463356800, 1463360400, 
    1463364000, 1463367600, 1463371200, 1463374800, 1463378400, 1463382000, 
    1463385600, 1463389200, 1463392800, 1463396400, 1463400000, 1463403600, 
    1463407200, 1463410800, 1463414400, 1463418000, 1463421600, 1463425200, 
    1463428800, 1463432400, 1463436000, 1463439600, 1463443200, 1463446800, 
    1463450400, 1463454000, 1463457600, 1463461200, 1463464800, 1463468400, 
    1463472000, 1463475600, 1463479200, 1463482800, 1463486400, 1463490000, 
    1463493600, 1463497200, 1463500800, 1463504400, 1463508000, 1463511600, 
    1463515200, 1463518800, 1463522400, 1463526000, 1463529600, 1463533200, 
    1463536800, 1463540400, 1463544000, 1463547600, 1463551200, 1463554800, 
    1463558400, 1463562000, 1463565600, 1463569200, 1463572800, 1463576400, 
    1463580000, 1463583600, 1463587200, 1463590800, 1463594400, 1463598000, 
    1463601600, 1463605200, 1463608800, 1463612400, 1463616000, 1463619600, 
    1463623200, 1463626800, 1463630400, 1463634000, 1463637600, 1463641200, 
    1463644800, 1463648400, 1463652000, 1463655600, 1463659200, 1463662800, 
    1463666400, 1463670000, 1463673600, 1463677200, 1463680800, 1463684400, 
    1463688000, 1463691600, 1463695200, 1463698800, 1463702400, 1463706000, 
    1463709600, 1463713200, 1463716800, 1463720400, 1463724000, 1463727600, 
    1463731200, 1463734800, 1463738400, 1463742000, 1463745600, 1463749200, 
    1463752800, 1463756400, 1463760000, 1463763600, 1463767200, 1463770800, 
    1463774400, 1463778000, 1463781600, 1463785200, 1463788800, 1463792400, 
    1463796000, 1463799600, 1463803200, 1463806800, 1463810400, 1463814000, 
    1463817600, 1463821200, 1463824800, 1463828400, 1463832000, 1463835600, 
    1463839200, 1463842800, 1463846400, 1463850000, 1463853600, 1463857200, 
    1463860800, 1463864400, 1463868000, 1463871600, 1463875200, 1463878800, 
    1463882400, 1463886000, 1463889600, 1463893200, 1463896800, 1463900400, 
    1463904000, 1463907600, 1463911200, 1463914800, 1463918400, 1463922000, 
    1463925600, 1463929200, 1463932800, 1463936400, 1463940000, 1463943600, 
    1463947200, 1463950800, 1463954400, 1463958000, 1463961600, 1463965200, 
    1463968800, 1463972400, 1463976000, 1463979600, 1463983200, 1463986800, 
    1463990400, 1463994000, 1463997600, 1464001200, 1464004800, 1464008400, 
    1464012000, 1464015600, 1464019200, 1464022800, 1464026400, 1464030000, 
    1464033600, 1464037200, 1464040800, 1464044400, 1464048000, 1464051600, 
    1464055200, 1464058800, 1464062400, 1464066000, 1464069600, 1464073200, 
    1464076800, 1464080400, 1464084000, 1464087600, 1464091200, 1464094800, 
    1464098400, 1464102000, 1464105600, 1464109200, 1464112800, 1464116400, 
    1464120000, 1464123600, 1464127200, 1464130800, 1464134400, 1464138000, 
    1464141600, 1464145200, 1464148800, 1464152400, 1464156000, 1464159600, 
    1464163200, 1464166800, 1464170400, 1464174000, 1464177600, 1464181200, 
    1464184800, 1464188400, 1464192000, 1464195600, 1464199200, 1464202800, 
    1464206400, 1464210000, 1464213600, 1464217200, 1464220800, 1464224400, 
    1464228000, 1464231600, 1464235200, 1464238800, 1464242400, 1464246000, 
    1464249600, 1464253200, 1464256800, 1464260400, 1464264000, 1464267600, 
    1464271200, 1464274800, 1464278400, 1464282000, 1464285600, 1464289200, 
    1464292800, 1464296400, 1464300000, 1464303600, 1464307200, 1464310800, 
    1464314400, 1464318000, 1464321600, 1464325200, 1464328800, 1464332400, 
    1464336000, 1464339600, 1464343200, 1464346800, 1464350400, 1464354000, 
    1464357600, 1464361200, 1464364800, 1464368400, 1464372000, 1464375600, 
    1464379200, 1464382800, 1464386400, 1464390000, 1464393600, 1464397200, 
    1464400800, 1464404400, 1464408000, 1464411600, 1464415200, 1464418800, 
    1464422400, 1464426000, 1464429600, 1464433200, 1464436800, 1464440400, 
    1464444000, 1464447600, 1464451200, 1464454800, 1464458400, 1464462000, 
    1464465600, 1464469200, 1464472800, 1464476400, 1464480000, 1464483600, 
    1464487200, 1464490800, 1464494400, 1464498000, 1464501600, 1464505200, 
    1464508800, 1464512400, 1464516000, 1464519600, 1464523200, 1464526800, 
    1464530400, 1464534000, 1464537600, 1464541200, 1464544800, 1464548400, 
    1464552000, 1464555600, 1464559200, 1464562800, 1464566400, 1464570000, 
    1464573600, 1464577200, 1464580800, 1464584400, 1464588000, 1464591600, 
    1464595200, 1464598800, 1464602400, 1464606000, 1464609600, 1464613200, 
    1464616800, 1464620400, 1464624000, 1464627600, 1464631200, 1464634800, 
    1464638400, 1464642000, 1464645600, 1464649200, 1464652800, 1464656400, 
    1464660000, 1464663600, 1464667200, 1464670800, 1464674400, 1464678000, 
    1464681600, 1464685200, 1464688800, 1464692400, 1464696000, 1464699600, 
    1464703200, 1464706800, 1464710400, 1464714000, 1464717600, 1464721200, 
    1464724800, 1464728400, 1464732000, 1464735600, 1464739200, 1464742800, 
    1464746400, 1464750000, 1464753600, 1464757200, 1464760800, 1464764400, 
    1464768000, 1464771600, 1464775200, 1464778800, 1464782400, 1464786000, 
    1464789600, 1464793200, 1464796800, 1464800400, 1464804000, 1464807600, 
    1464811200, 1464814800, 1464818400, 1464822000, 1464825600, 1464829200, 
    1464832800, 1464836400, 1464840000, 1464843600, 1464847200, 1464850800, 
    1464854400, 1464858000, 1464861600, 1464865200, 1464868800, 1464872400, 
    1464876000, 1464879600, 1464883200, 1464886800, 1464890400, 1464894000, 
    1464897600, 1464901200, 1464904800, 1464908400, 1464912000, 1464915600, 
    1464919200, 1464922800, 1464926400, 1464930000, 1464933600, 1464937200, 
    1464940800, 1464944400, 1464948000, 1464951600, 1464955200, 1464958800, 
    1464962400, 1464966000, 1464969600, 1464973200, 1464976800, 1464980400, 
    1464984000, 1464987600, 1464991200, 1464994800, 1464998400, 1465002000, 
    1465005600, 1465009200, 1465012800, 1465016400, 1465020000, 1465023600, 
    1465027200, 1465030800, 1465034400, 1465038000, 1465041600, 1465045200, 
    1465048800, 1465052400, 1465056000, 1465059600, 1465063200, 1465066800, 
    1465070400, 1465074000, 1465077600, 1465081200, 1465084800, 1465088400, 
    1465092000, 1465095600, 1465099200, 1465102800, 1465106400, 1465110000, 
    1465113600, 1465117200, 1465120800, 1465124400, 1465128000, 1465131600, 
    1465135200, 1465138800, 1465142400, 1465146000, 1465149600, 1465153200, 
    1465156800, 1465160400, 1465164000, 1465167600, 1465171200, 1465174800, 
    1465178400, 1465182000, 1465185600, 1465189200, 1465192800, 1465196400, 
    1465200000, 1465203600, 1465207200, 1465210800, 1465214400, 1465218000, 
    1465221600, 1465225200, 1465228800, 1465232400, 1465236000, 1465239600, 
    1465243200, 1465246800, 1465250400, 1465254000, 1465257600, 1465261200, 
    1465264800, 1465268400, 1465272000, 1465275600, 1465279200, 1465282800, 
    1465286400, 1465290000, 1465293600, 1465297200, 1465300800, 1465304400, 
    1465308000, 1465311600, 1465315200, 1465318800, 1465322400, 1465326000, 
    1465329600, 1465333200, 1465336800, 1465340400, 1465344000, 1465347600, 
    1465351200, 1465354800, 1465358400, 1465362000, 1465365600, 1465369200, 
    1465372800, 1465376400, 1465380000, 1465383600, 1465387200, 1465390800, 
    1465394400, 1465398000, 1465401600, 1465405200, 1465408800, 1465412400, 
    1465416000, 1465419600, 1465423200, 1465426800, 1465430400, 1465434000, 
    1465437600, 1465441200, 1465444800, 1465448400, 1465452000, 1465455600, 
    1465459200, 1465462800, 1465466400, 1465470000, 1465473600, 1465477200, 
    1465480800, 1465484400, 1465488000, 1465491600, 1465495200, 1465498800, 
    1465502400, 1465506000, 1465509600, 1465513200, 1465516800, 1465520400, 
    1465524000, 1465527600, 1465531200, 1465534800, 1465538400, 1465542000, 
    1465545600, 1465549200, 1465552800, 1465556400, 1465560000, 1465563600, 
    1465567200, 1465570800, 1465574400, 1465578000, 1465581600, 1465585200, 
    1465588800, 1465592400, 1465596000, 1465599600, 1465603200, 1465606800, 
    1465610400, 1465614000, 1465617600, 1465621200, 1465624800, 1465628400, 
    1465632000, 1465635600, 1465639200, 1465642800, 1465646400, 1465650000, 
    1465653600, 1465657200, 1465660800, 1465664400, 1465668000, 1465671600, 
    1465675200, 1465678800, 1465682400, 1465686000, 1465689600, 1465693200, 
    1465696800, 1465700400, 1465704000, 1465707600, 1465711200, 1465714800, 
    1465718400, 1465722000, 1465725600, 1465729200, 1465732800, 1465736400, 
    1465740000, 1465743600, 1465747200, 1465750800, 1465754400, 1465758000, 
    1465761600, 1465765200, 1465768800, 1465772400, 1465776000, 1465779600, 
    1465783200, 1465786800, 1465790400, 1465794000, 1465797600, 1465801200, 
    1465804800, 1465808400, 1465812000, 1465815600, 1465819200, 1465822800, 
    1465826400, 1465830000, 1465833600, 1465837200, 1465840800, 1465844400, 
    1465848000, 1465851600, 1465855200, 1465858800, 1465862400, 1465866000, 
    1465869600, 1465873200, 1465876800, 1465880400, 1465884000, 1465887600, 
    1465891200, 1465894800, 1465898400, 1465902000, 1465905600, 1465909200, 
    1465912800, 1465916400, 1465920000, 1465923600, 1465927200, 1465930800, 
    1465934400, 1465938000, 1465941600, 1465945200, 1465948800, 1465952400, 
    1465956000, 1465959600, 1465963200, 1465966800, 1465970400, 1465974000, 
    1465977600, 1465981200, 1465984800, 1465988400, 1465992000, 1465995600, 
    1465999200, 1466002800, 1466006400, 1466010000, 1466013600, 1466017200, 
    1466020800, 1466024400, 1466028000, 1466031600, 1466035200, 1466038800, 
    1466042400, 1466046000, 1466049600, 1466053200, 1466056800, 1466060400, 
    1466064000, 1466067600, 1466071200, 1466074800, 1466078400, 1466082000, 
    1466085600, 1466089200, 1466092800, 1466096400, 1466100000, 1466103600, 
    1466107200, 1466110800, 1466114400, 1466118000, 1466121600, 1466125200, 
    1466128800, 1466132400, 1466136000, 1466139600, 1466143200, 1466146800, 
    1466150400, 1466154000, 1466157600, 1466161200, 1466164800, 1466168400, 
    1466172000, 1466175600, 1466179200, 1466182800, 1466186400, 1466190000, 
    1466193600, 1466197200, 1466200800, 1466204400, 1466208000, 1466211600, 
    1466215200, 1466218800, 1466222400, 1466226000, 1466229600, 1466233200, 
    1466236800, 1466240400, 1466244000, 1466247600, 1466251200, 1466254800, 
    1466258400, 1466262000, 1466265600, 1466269200, 1466272800, 1466276400, 
    1466280000, 1466283600, 1466287200, 1466290800, 1466294400, 1466298000, 
    1466301600, 1466305200, 1466308800, 1466312400, 1466316000, 1466319600, 
    1466323200, 1466326800, 1466330400, 1466334000, 1466337600, 1466341200, 
    1466344800, 1466348400, 1466352000, 1466355600, 1466359200, 1466362800, 
    1466366400, 1466370000, 1466373600, 1466377200, 1466380800, 1466384400, 
    1466388000, 1466391600, 1466395200, 1466398800, 1466402400, 1466406000, 
    1466409600, 1466413200, 1466416800, 1466420400, 1466424000, 1466427600, 
    1466431200, 1466434800, 1466438400, 1466442000, 1466445600, 1466449200, 
    1466452800, 1466456400, 1466460000, 1466463600, 1466467200, 1466470800, 
    1466474400, 1466478000, 1466481600, 1466485200, 1466488800, 1466492400, 
    1466496000, 1466499600, 1466503200, 1466506800, 1466510400, 1466514000, 
    1466517600, 1466521200, 1466524800, 1466528400, 1466532000, 1466535600, 
    1466539200, 1466542800, 1466546400, 1466550000, 1466553600, 1466557200, 
    1466560800, 1466564400, 1466568000, 1466571600, 1466575200, 1466578800, 
    1466582400, 1466586000, 1466589600, 1466593200, 1466596800, 1466600400, 
    1466604000, 1466607600, 1466611200, 1466614800, 1466618400, 1466622000, 
    1466625600, 1466629200, 1466632800, 1466636400, 1466640000, 1466643600, 
    1466647200, 1466650800, 1466654400, 1466658000, 1466661600, 1466665200, 
    1466668800, 1466672400, 1466676000, 1466679600, 1466683200, 1466686800, 
    1466690400, 1466694000, 1466697600, 1466701200, 1466704800, 1466708400, 
    1466712000, 1466715600, 1466719200, 1466722800, 1466726400, 1466730000, 
    1466733600, 1466737200, 1466740800, 1466744400, 1466748000, 1466751600, 
    1466755200, 1466758800, 1466762400, 1466766000, 1466769600, 1466773200, 
    1466776800, 1466780400, 1466784000, 1466787600, 1466791200, 1466794800, 
    1466798400, 1466802000, 1466805600, 1466809200, 1466812800, 1466816400, 
    1466820000, 1466823600, 1466827200, 1466830800, 1466834400, 1466838000, 
    1466841600, 1466845200, 1466848800, 1466852400, 1466856000, 1466859600, 
    1466863200, 1466866800, 1466870400, 1466874000, 1466877600, 1466881200, 
    1466884800, 1466888400, 1466892000, 1466895600, 1466899200, 1466902800, 
    1466906400, 1466910000, 1466913600, 1466917200, 1466920800, 1466924400, 
    1466928000, 1466931600, 1466935200, 1466938800, 1466942400, 1466946000, 
    1466949600, 1466953200, 1466956800, 1466960400, 1466964000, 1466967600, 
    1466971200, 1466974800, 1466978400, 1466982000, 1466985600, 1466989200, 
    1466992800, 1466996400, 1467000000, 1467003600, 1467007200, 1467010800, 
    1467014400, 1467018000, 1467021600, 1467025200, 1467028800, 1467032400, 
    1467036000, 1467039600, 1467043200, 1467046800, 1467050400, 1467054000, 
    1467057600, 1467061200, 1467064800, 1467068400, 1467072000, 1467075600, 
    1467079200, 1467082800, 1467086400, 1467090000, 1467093600, 1467097200, 
    1467100800, 1467104400, 1467108000, 1467111600, 1467115200, 1467118800, 
    1467122400, 1467126000, 1467129600, 1467133200, 1467136800, 1467140400, 
    1467144000, 1467147600, 1467151200, 1467154800, 1467158400, 1467162000, 
    1467165600, 1467169200, 1467172800, 1467176400, 1467180000, 1467183600, 
    1467187200, 1467190800, 1467194400, 1467198000, 1467201600, 1467205200, 
    1467208800, 1467212400, 1467216000, 1467219600, 1467223200, 1467226800, 
    1467230400, 1467234000, 1467237600, 1467241200, 1467244800, 1467248400, 
    1467252000, 1467255600, 1467259200, 1467262800, 1467266400, 1467270000, 
    1467273600, 1467277200, 1467280800, 1467284400, 1467288000, 1467291600, 
    1467295200, 1467298800, 1467302400, 1467306000, 1467309600, 1467313200, 
    1467316800, 1467320400, 1467324000, 1467327600, 1467331200, 1467334800, 
    1467338400, 1467342000, 1467345600, 1467349200, 1467352800, 1467356400, 
    1467360000, 1467363600, 1467367200, 1467370800, 1467374400, 1467378000, 
    1467381600, 1467385200, 1467388800, 1467392400, 1467396000, 1467399600, 
    1467403200, 1467406800, 1467410400, 1467414000, 1467417600, 1467421200, 
    1467424800, 1467428400, 1467432000, 1467435600, 1467439200, 1467442800, 
    1467446400, 1467450000, 1467453600, 1467457200, 1467460800, 1467464400, 
    1467468000, 1467471600, 1467475200, 1467478800, 1467482400, 1467486000, 
    1467489600, 1467493200, 1467496800, 1467500400, 1467504000, 1467507600, 
    1467511200, 1467514800, 1467518400, 1467522000, 1467525600, 1467529200, 
    1467532800, 1467536400, 1467540000, 1467543600, 1467547200, 1467550800, 
    1467554400, 1467558000, 1467561600, 1467565200, 1467568800, 1467572400, 
    1467576000, 1467579600, 1467583200, 1467586800, 1467590400, 1467594000, 
    1467597600, 1467601200, 1467604800, 1467608400, 1467612000, 1467615600, 
    1467619200, 1467622800, 1467626400, 1467630000, 1467633600, 1467637200, 
    1467640800, 1467644400, 1467648000, 1467651600, 1467655200, 1467658800, 
    1467662400, 1467666000, 1467669600, 1467673200, 1467676800, 1467680400, 
    1467684000, 1467687600, 1467691200, 1467694800, 1467698400, 1467702000, 
    1467705600, 1467709200, 1467712800, 1467716400, 1467720000, 1467723600, 
    1467727200, 1467730800, 1467734400, 1467738000, 1467741600, 1467745200, 
    1467748800, 1467752400, 1467756000, 1467759600, 1467763200, 1467766800, 
    1467770400, 1467774000, 1467777600, 1467781200, 1467784800, 1467788400, 
    1467792000, 1467795600, 1467799200, 1467802800, 1467806400, 1467810000, 
    1467813600, 1467817200, 1467820800, 1467824400, 1467828000, 1467831600, 
    1467835200, 1467838800, 1467842400, 1467846000, 1467849600, 1467853200, 
    1467856800, 1467860400, 1467864000, 1467867600, 1467871200, 1467874800, 
    1467878400, 1467882000, 1467885600, 1467889200, 1467892800, 1467896400, 
    1467900000, 1467903600, 1467907200, 1467910800, 1467914400, 1467918000, 
    1467921600, 1467925200, 1467928800, 1467932400, 1467936000, 1467939600, 
    1467943200, 1467946800, 1467950400, 1467954000, 1467957600, 1467961200, 
    1467964800, 1467968400, 1467972000, 1467975600, 1467979200, 1467982800, 
    1467986400, 1467990000, 1467993600, 1467997200, 1468000800, 1468004400, 
    1468008000, 1468011600, 1468015200, 1468018800, 1468022400, 1468026000, 
    1468029600, 1468033200, 1468036800, 1468040400, 1468044000, 1468047600, 
    1468051200, 1468054800, 1468058400, 1468062000, 1468065600, 1468069200, 
    1468072800, 1468076400, 1468080000, 1468083600, 1468087200, 1468090800, 
    1468094400, 1468098000, 1468101600, 1468105200, 1468108800, 1468112400, 
    1468116000, 1468119600, 1468123200, 1468126800, 1468130400, 1468134000, 
    1468137600, 1468141200, 1468144800, 1468148400, 1468152000, 1468155600, 
    1468159200, 1468162800, 1468166400, 1468170000, 1468173600, 1468177200, 
    1468180800, 1468184400, 1468188000, 1468191600, 1468195200, 1468198800, 
    1468202400, 1468206000, 1468209600, 1468213200, 1468216800, 1468220400, 
    1468224000, 1468227600, 1468231200, 1468234800, 1468238400, 1468242000, 
    1468245600, 1468249200, 1468252800, 1468256400, 1468260000, 1468263600, 
    1468267200, 1468270800, 1468274400, 1468278000, 1468281600, 1468285200, 
    1468288800, 1468292400, 1468296000, 1468299600, 1468303200, 1468306800, 
    1468310400, 1468314000, 1468317600, 1468321200, 1468324800, 1468328400, 
    1468332000, 1468335600, 1468339200, 1468342800, 1468346400, 1468350000, 
    1468353600, 1468357200, 1468360800, 1468364400, 1468368000, 1468371600, 
    1468375200, 1468378800, 1468382400, 1468386000, 1468389600, 1468393200, 
    1468396800, 1468400400, 1468404000, 1468407600, 1468411200, 1468414800, 
    1468418400, 1468422000, 1468425600, 1468429200, 1468432800, 1468436400, 
    1468440000, 1468443600, 1468447200, 1468450800, 1468454400, 1468458000, 
    1468461600, 1468465200, 1468468800, 1468472400, 1468476000, 1468479600, 
    1468483200, 1468486800, 1468490400, 1468494000, 1468497600, 1468501200, 
    1468504800, 1468508400, 1468512000, 1468515600, 1468519200, 1468522800, 
    1468526400, 1468530000, 1468533600, 1468537200, 1468540800, 1468544400, 
    1468548000, 1468551600, 1468555200, 1468558800, 1468562400, 1468566000, 
    1468569600, 1468573200, 1468576800, 1468580400, 1468584000, 1468587600, 
    1468591200, 1468594800, 1468598400, 1468602000, 1468605600, 1468609200, 
    1468612800, 1468616400, 1468620000, 1468623600, 1468627200, 1468630800, 
    1468634400, 1468638000, 1468641600, 1468645200, 1468648800, 1468652400, 
    1468656000, 1468659600, 1468663200, 1468666800, 1468670400, 1468674000, 
    1468677600, 1468681200, 1468684800, 1468688400, 1468692000, 1468695600, 
    1468699200, 1468702800, 1468706400, 1468710000, 1468713600, 1468717200, 
    1468720800, 1468724400, 1468728000, 1468731600, 1468735200, 1468738800, 
    1468742400, 1468746000, 1468749600, 1468753200, 1468756800, 1468760400, 
    1468764000, 1468767600, 1468771200, 1468774800, 1468778400, 1468782000, 
    1468785600, 1468789200, 1468792800, 1468796400, 1468800000, 1468803600, 
    1468807200, 1468810800, 1468814400, 1468818000, 1468821600, 1468825200, 
    1468828800, 1468832400, 1468836000, 1468839600, 1468843200, 1468846800, 
    1468850400, 1468854000, 1468857600, 1468861200, 1468864800, 1468868400, 
    1468872000, 1468875600, 1468879200, 1468882800, 1468886400, 1468890000, 
    1468893600, 1468897200, 1468900800, 1468904400, 1468908000, 1468911600, 
    1468915200, 1468918800, 1468922400, 1468926000, 1468929600, 1468933200, 
    1468936800, 1468940400, 1468944000, 1468947600, 1468951200, 1468954800, 
    1468958400, 1468962000, 1468965600, 1468969200, 1468972800, 1468976400, 
    1468980000, 1468983600, 1468987200, 1468990800, 1468994400, 1468998000, 
    1469001600, 1469005200, 1469008800, 1469012400, 1469016000, 1469019600, 
    1469023200, 1469026800, 1469030400, 1469034000, 1469037600, 1469041200, 
    1469044800, 1469048400, 1469052000, 1469055600, 1469059200, 1469062800, 
    1469066400, 1469070000, 1469073600, 1469077200, 1469080800, 1469084400, 
    1469088000, 1469091600, 1469095200, 1469098800, 1469102400, 1469106000, 
    1469109600, 1469113200, 1469116800, 1469120400, 1469124000, 1469127600, 
    1469131200, 1469134800, 1469138400, 1469142000, 1469145600, 1469149200, 
    1469152800, 1469156400, 1469160000, 1469163600, 1469167200, 1469170800, 
    1469174400, 1469178000, 1469181600, 1469185200, 1469188800, 1469192400, 
    1469196000, 1469199600, 1469203200, 1469206800, 1469210400, 1469214000, 
    1469217600, 1469221200, 1469224800, 1469228400, 1469232000, 1469235600, 
    1469239200, 1469242800, 1469246400, 1469250000, 1469253600, 1469257200, 
    1469260800, 1469264400, 1469268000, 1469271600, 1469275200, 1469278800, 
    1469282400, 1469286000, 1469289600, 1469293200, 1469296800, 1469300400, 
    1469304000, 1469307600, 1469311200, 1469314800, 1469318400, 1469322000, 
    1469325600, 1469329200, 1469332800, 1469336400, 1469340000, 1469343600, 
    1469347200, 1469350800, 1469354400, 1469358000, 1469361600, 1469365200, 
    1469368800, 1469372400, 1469376000, 1469379600, 1469383200, 1469386800, 
    1469390400, 1469394000, 1469397600, 1469401200, 1469404800, 1469408400, 
    1469412000, 1469415600, 1469419200, 1469422800, 1469426400, 1469430000, 
    1469433600, 1469437200, 1469440800, 1469444400, 1469448000, 1469451600, 
    1469455200, 1469458800, 1469462400, 1469466000, 1469469600, 1469473200, 
    1469476800, 1469480400, 1469484000, 1469487600, 1469491200, 1469494800, 
    1469498400, 1469502000, 1469505600, 1469509200, 1469512800, 1469516400, 
    1469520000, 1469523600, 1469527200, 1469530800, 1469534400, 1469538000, 
    1469541600, 1469545200, 1469548800, 1469552400, 1469556000, 1469559600, 
    1469563200, 1469566800, 1469570400, 1469574000, 1469577600, 1469581200, 
    1469584800, 1469588400, 1469592000, 1469595600, 1469599200, 1469602800, 
    1469606400, 1469610000, 1469613600, 1469617200, 1469620800, 1469624400, 
    1469628000, 1469631600, 1469635200, 1469638800, 1469642400, 1469646000, 
    1469649600, 1469653200, 1469656800, 1469660400, 1469664000, 1469667600, 
    1469671200, 1469674800, 1469678400, 1469682000, 1469685600, 1469689200, 
    1469692800, 1469696400, 1469700000, 1469703600, 1469707200, 1469710800, 
    1469714400, 1469718000, 1469721600, 1469725200, 1469728800, 1469732400, 
    1469736000, 1469739600, 1469743200, 1469746800, 1469750400, 1469754000, 
    1469757600, 1469761200, 1469764800, 1469768400, 1469772000, 1469775600, 
    1469779200, 1469782800, 1469786400, 1469790000, 1469793600, 1469797200, 
    1469800800, 1469804400, 1469808000, 1469811600, 1469815200, 1469818800, 
    1469822400, 1469826000, 1469829600, 1469833200, 1469836800, 1469840400, 
    1469844000, 1469847600, 1469851200, 1469854800, 1469858400, 1469862000, 
    1469865600, 1469869200, 1469872800, 1469876400, 1469880000, 1469883600, 
    1469887200, 1469890800, 1469894400, 1469898000, 1469901600, 1469905200, 
    1469908800, 1469912400, 1469916000, 1469919600, 1469923200, 1469926800, 
    1469930400, 1469934000, 1469937600, 1469941200, 1469944800, 1469948400, 
    1469952000, 1469955600, 1469959200, 1469962800, 1469966400, 1469970000, 
    1469973600, 1469977200, 1469980800, 1469984400, 1469988000, 1469991600, 
    1469995200, 1469998800, 1470002400, 1470006000, 1470009600, 1470013200, 
    1470016800, 1470020400, 1470024000, 1470027600, 1470031200, 1470034800, 
    1470038400, 1470042000, 1470045600, 1470049200, 1470052800, 1470056400, 
    1470060000, 1470063600, 1470067200, 1470070800, 1470074400, 1470078000, 
    1470081600, 1470085200, 1470088800, 1470092400, 1470096000, 1470099600, 
    1470103200, 1470106800, 1470110400, 1470114000, 1470117600, 1470121200, 
    1470124800, 1470128400, 1470132000, 1470135600, 1470139200, 1470142800, 
    1470146400, 1470150000, 1470153600, 1470157200, 1470160800, 1470164400, 
    1470168000, 1470171600, 1470175200, 1470178800, 1470182400, 1470186000, 
    1470189600, 1470193200, 1470196800, 1470200400, 1470204000, 1470207600, 
    1470211200, 1470214800, 1470218400, 1470222000, 1470225600, 1470229200, 
    1470232800, 1470236400, 1470240000, 1470243600, 1470247200, 1470250800, 
    1470254400, 1470258000, 1470261600, 1470265200, 1470268800, 1470272400, 
    1470276000, 1470279600, 1470283200, 1470286800, 1470290400, 1470294000, 
    1470297600, 1470301200, 1470304800, 1470308400, 1470312000, 1470315600, 
    1470319200, 1470322800, 1470326400, 1470330000, 1470333600, 1470337200, 
    1470340800, 1470344400, 1470348000, 1470351600, 1470355200, 1470358800, 
    1470362400, 1470366000, 1470369600, 1470373200, 1470376800, 1470380400, 
    1470384000, 1470387600, 1470391200, 1470394800, 1470398400, 1470402000, 
    1470405600, 1470409200, 1470412800, 1470416400, 1470420000, 1470423600, 
    1470427200, 1470430800, 1470434400, 1470438000, 1470441600, 1470445200, 
    1470448800, 1470452400, 1470456000, 1470459600, 1470463200, 1470466800, 
    1470470400, 1470474000, 1470477600, 1470481200, 1470484800, 1470488400, 
    1470492000, 1470495600, 1470499200, 1470502800, 1470506400, 1470510000, 
    1470513600, 1470517200, 1470520800, 1470524400, 1470528000, 1470531600, 
    1470535200, 1470538800, 1470542400, 1470546000, 1470549600, 1470553200, 
    1470556800, 1470560400, 1470564000, 1470567600, 1470571200, 1470574800, 
    1470578400, 1470582000, 1470585600, 1470589200, 1470592800, 1470596400, 
    1470600000, 1470603600, 1470607200, 1470610800, 1470614400, 1470618000, 
    1470621600, 1470625200, 1470628800, 1470632400, 1470636000, 1470639600, 
    1470643200, 1470646800, 1470650400, 1470654000, 1470657600, 1470661200, 
    1470664800, 1470668400, 1470672000, 1470675600, 1470679200, 1470682800, 
    1470686400, 1470690000, 1470693600, 1470697200, 1470700800, 1470704400, 
    1470708000, 1470711600, 1470715200, 1470718800, 1470722400, 1470726000, 
    1470729600, 1470733200, 1470736800, 1470740400, 1470744000, 1470747600, 
    1470751200, 1470754800, 1470758400, 1470762000, 1470765600, 1470769200, 
    1470772800, 1470776400, 1470780000, 1470783600, 1470787200, 1470790800, 
    1470794400, 1470798000, 1470801600, 1470805200, 1470808800, 1470812400, 
    1470816000, 1470819600, 1470823200, 1470826800, 1470830400, 1470834000, 
    1470837600, 1470841200, 1470844800, 1470848400, 1470852000, 1470855600, 
    1470859200, 1470862800, 1470866400, 1470870000, 1470873600, 1470877200, 
    1470880800, 1470884400, 1470888000, 1470891600, 1470895200, 1470898800, 
    1470902400, 1470906000, 1470909600, 1470913200, 1470916800, 1470920400, 
    1470924000, 1470927600, 1470931200, 1470934800, 1470938400, 1470942000, 
    1470945600, 1470949200, 1470952800, 1470956400, 1470960000, 1470963600, 
    1470967200, 1470970800, 1470974400, 1470978000, 1470981600, 1470985200, 
    1470988800, 1470992400, 1470996000, 1470999600, 1471003200, 1471006800, 
    1471010400, 1471014000, 1471017600, 1471021200, 1471024800, 1471028400, 
    1471032000, 1471035600, 1471039200, 1471042800, 1471046400, 1471050000, 
    1471053600, 1471057200, 1471060800, 1471064400, 1471068000, 1471071600, 
    1471075200, 1471078800, 1471082400, 1471086000, 1471089600, 1471093200, 
    1471096800, 1471100400, 1471104000, 1471107600, 1471111200, 1471114800, 
    1471118400, 1471122000, 1471125600, 1471129200, 1471132800, 1471136400, 
    1471140000, 1471143600, 1471147200, 1471150800, 1471154400, 1471158000, 
    1471161600, 1471165200, 1471168800, 1471172400, 1471176000, 1471179600, 
    1471183200, 1471186800, 1471190400, 1471194000, 1471197600, 1471201200, 
    1471204800, 1471208400, 1471212000, 1471215600, 1471219200, 1471222800, 
    1471226400, 1471230000, 1471233600, 1471237200, 1471240800, 1471244400, 
    1471248000, 1471251600, 1471255200, 1471258800, 1471262400, 1471266000, 
    1471269600, 1471273200, 1471276800, 1471280400, 1471284000, 1471287600, 
    1471291200, 1471294800, 1471298400, 1471302000, 1471305600, 1471309200, 
    1471312800, 1471316400, 1471320000, 1471323600, 1471327200, 1471330800, 
    1471334400, 1471338000, 1471341600, 1471345200, 1471348800, 1471352400, 
    1471356000, 1471359600, 1471363200, 1471366800, 1471370400, 1471374000, 
    1471377600, 1471381200, 1471384800, 1471388400, 1471392000, 1471395600, 
    1471399200, 1471402800, 1471406400, 1471410000, 1471413600, 1471417200, 
    1471420800, 1471424400, 1471428000, 1471431600, 1471435200, 1471438800, 
    1471442400, 1471446000, 1471449600, 1471453200, 1471456800, 1471460400, 
    1471464000, 1471467600, 1471471200, 1471474800, 1471478400, 1471482000, 
    1471485600, 1471489200, 1471492800, 1471496400, 1471500000, 1471503600, 
    1471507200, 1471510800, 1471514400, 1471518000, 1471521600, 1471525200, 
    1471528800, 1471532400, 1471536000, 1471539600, 1471543200, 1471546800, 
    1471550400, 1471554000, 1471557600, 1471561200, 1471564800, 1471568400, 
    1471572000, 1471575600, 1471579200, 1471582800, 1471586400, 1471590000, 
    1471593600, 1471597200, 1471600800, 1471604400, 1471608000, 1471611600, 
    1471615200, 1471618800, 1471622400, 1471626000, 1471629600, 1471633200, 
    1471636800, 1471640400, 1471644000, 1471647600, 1471651200, 1471654800, 
    1471658400, 1471662000, 1471665600, 1471669200, 1471672800, 1471676400, 
    1471680000, 1471683600, 1471687200, 1471690800, 1471694400, 1471698000, 
    1471701600, 1471705200, 1471708800, 1471712400, 1471716000, 1471719600, 
    1471723200, 1471726800, 1471730400, 1471734000, 1471737600, 1471741200, 
    1471744800, 1471748400, 1471752000, 1471755600, 1471759200, 1471762800, 
    1471766400, 1471770000, 1471773600, 1471777200, 1471780800, 1471784400, 
    1471788000, 1471791600, 1471795200, 1471798800, 1471802400, 1471806000, 
    1471809600, 1471813200, 1471816800, 1471820400, 1471824000, 1471827600, 
    1471831200, 1471834800, 1471838400, 1471842000, 1471845600, 1471849200, 
    1471852800, 1471856400, 1471860000, 1471863600, 1471867200, 1471870800, 
    1471874400, 1471878000, 1471881600, 1471885200, 1471888800, 1471892400, 
    1471896000, 1471899600, 1471903200, 1471906800, 1471910400, 1471914000, 
    1471917600, 1471921200, 1471924800, 1471928400, 1471932000, 1471935600, 
    1471939200, 1471942800, 1471946400, 1471950000, 1471953600, 1471957200, 
    1471960800, 1471964400, 1471968000, 1471971600, 1471975200, 1471978800, 
    1471982400, 1471986000, 1471989600, 1471993200, 1471996800, 1472000400, 
    1472004000, 1472007600, 1472011200, 1472014800, 1472018400, 1472022000, 
    1472025600, 1472029200, 1472032800, 1472036400, 1472040000, 1472043600, 
    1472047200, 1472050800, 1472054400, 1472058000, 1472061600, 1472065200, 
    1472068800, 1472072400, 1472076000, 1472079600, 1472083200, 1472086800, 
    1472090400, 1472094000, 1472097600, 1472101200, 1472104800, 1472108400, 
    1472112000, 1472115600, 1472119200, 1472122800, 1472126400, 1472130000, 
    1472133600, 1472137200, 1472140800, 1472144400, 1472148000, 1472151600, 
    1472155200, 1472158800, 1472162400, 1472166000, 1472169600, 1472173200, 
    1472176800, 1472180400, 1472184000, 1472187600, 1472191200, 1472194800, 
    1472198400, 1472202000, 1472205600, 1472209200, 1472212800, 1472216400, 
    1472220000, 1472223600, 1472227200, 1472230800, 1472234400, 1472238000, 
    1472241600, 1472245200, 1472248800, 1472252400, 1472256000, 1472259600, 
    1472263200, 1472266800, 1472270400, 1472274000, 1472277600, 1472281200, 
    1472284800, 1472288400, 1472292000, 1472295600, 1472299200, 1472302800, 
    1472306400, 1472310000, 1472313600, 1472317200, 1472320800, 1472324400, 
    1472328000, 1472331600, 1472335200, 1472338800, 1472342400, 1472346000, 
    1472349600, 1472353200, 1472356800, 1472360400, 1472364000, 1472367600, 
    1472371200, 1472374800, 1472378400, 1472382000, 1472385600, 1472389200, 
    1472392800, 1472396400, 1472400000, 1472403600, 1472407200, 1472410800, 
    1472414400, 1472418000, 1472421600, 1472425200, 1472428800, 1472432400, 
    1472436000, 1472439600, 1472443200, 1472446800, 1472450400, 1472454000, 
    1472457600, 1472461200, 1472464800, 1472468400, 1472472000, 1472475600, 
    1472479200, 1472482800, 1472486400, 1472490000, 1472493600, 1472497200, 
    1472500800, 1472504400, 1472508000, 1472511600, 1472515200, 1472518800, 
    1472522400, 1472526000, 1472529600, 1472533200, 1472536800, 1472540400, 
    1472544000, 1472547600, 1472551200, 1472554800, 1472558400, 1472562000, 
    1472565600, 1472569200, 1472572800, 1472576400, 1472580000, 1472583600, 
    1472587200, 1472590800, 1472594400, 1472598000, 1472601600, 1472605200, 
    1472608800, 1472612400, 1472616000, 1472619600, 1472623200, 1472626800, 
    1472630400, 1472634000, 1472637600, 1472641200, 1472644800, 1472648400, 
    1472652000, 1472655600, 1472659200, 1472662800, 1472666400, 1472670000, 
    1472673600, 1472677200, 1472680800, 1472684400, 1472688000, 1472691600, 
    1472695200, 1472698800, 1472702400, 1472706000, 1472709600, 1472713200, 
    1472716800, 1472720400, 1472724000, 1472727600, 1472731200, 1472734800, 
    1472738400, 1472742000, 1472745600, 1472749200, 1472752800, 1472756400, 
    1472760000, 1472763600, 1472767200, 1472770800, 1472774400, 1472778000, 
    1472781600, 1472785200, 1472788800, 1472792400, 1472796000, 1472799600, 
    1472803200, 1472806800, 1472810400, 1472814000, 1472817600, 1472821200, 
    1472824800, 1472828400, 1472832000, 1472835600, 1472839200, 1472842800, 
    1472846400, 1472850000, 1472853600, 1472857200, 1472860800, 1472864400, 
    1472868000, 1472871600, 1472875200, 1472878800, 1472882400, 1472886000, 
    1472889600, 1472893200, 1472896800, 1472900400, 1472904000, 1472907600, 
    1472911200, 1472914800, 1472918400, 1472922000, 1472925600, 1472929200, 
    1472932800, 1472936400, 1472940000, 1472943600, 1472947200, 1472950800, 
    1472954400, 1472958000, 1472961600, 1472965200, 1472968800, 1472972400, 
    1472976000, 1472979600, 1472983200, 1472986800, 1472990400, 1472994000, 
    1472997600, 1473001200, 1473004800, 1473008400, 1473012000, 1473015600, 
    1473019200, 1473022800, 1473026400, 1473030000, 1473033600, 1473037200, 
    1473040800, 1473044400, 1473048000, 1473051600, 1473055200, 1473058800, 
    1473062400, 1473066000, 1473069600, 1473073200, 1473076800, 1473080400, 
    1473084000, 1473087600, 1473091200, 1473094800, 1473098400, 1473102000, 
    1473105600, 1473109200, 1473112800, 1473116400, 1473120000, 1473123600, 
    1473127200, 1473130800, 1473134400, 1473138000, 1473141600, 1473145200, 
    1473148800, 1473152400, 1473156000, 1473159600, 1473163200, 1473166800, 
    1473170400, 1473174000, 1473177600, 1473181200, 1473184800, 1473188400, 
    1473192000, 1473195600, 1473199200, 1473202800, 1473206400, 1473210000, 
    1473213600, 1473217200, 1473220800, 1473224400, 1473228000, 1473231600, 
    1473235200, 1473238800, 1473242400, 1473246000, 1473249600, 1473253200, 
    1473256800, 1473260400, 1473264000, 1473267600, 1473271200, 1473274800, 
    1473278400, 1473282000, 1473285600, 1473289200, 1473292800, 1473296400, 
    1473300000, 1473303600, 1473307200, 1473310800, 1473314400, 1473318000, 
    1473321600, 1473325200, 1473328800, 1473332400, 1473336000, 1473339600, 
    1473343200, 1473346800, 1473350400, 1473354000, 1473357600, 1473361200, 
    1473364800, 1473368400, 1473372000, 1473375600, 1473379200, 1473382800, 
    1473386400, 1473390000, 1473393600, 1473397200, 1473400800, 1473404400, 
    1473408000, 1473411600, 1473415200, 1473418800, 1473422400, 1473426000, 
    1473429600, 1473433200, 1473436800, 1473440400, 1473444000, 1473447600, 
    1473451200, 1473454800, 1473458400, 1473462000, 1473465600, 1473469200, 
    1473472800, 1473476400, 1473480000, 1473483600, 1473487200, 1473490800, 
    1473494400, 1473498000, 1473501600, 1473505200, 1473508800, 1473512400, 
    1473516000, 1473519600, 1473523200, 1473526800, 1473530400, 1473534000, 
    1473537600, 1473541200, 1473544800, 1473548400, 1473552000, 1473555600, 
    1473559200, 1473562800, 1473566400, 1473570000, 1473573600, 1473577200, 
    1473580800, 1473584400, 1473588000, 1473591600, 1473595200, 1473598800, 
    1473602400, 1473606000, 1473609600, 1473613200, 1473616800, 1473620400, 
    1473624000, 1473627600, 1473631200, 1473634800, 1473638400, 1473642000, 
    1473645600, 1473649200, 1473652800, 1473656400, 1473660000, 1473663600, 
    1473667200, 1473670800, 1473674400, 1473678000, 1473681600, 1473685200, 
    1473688800, 1473692400, 1473696000, 1473699600, 1473703200, 1473706800, 
    1473710400, 1473714000, 1473717600, 1473721200, 1473724800, 1473728400, 
    1473732000, 1473735600, 1473739200, 1473742800, 1473746400, 1473750000, 
    1473753600, 1473757200, 1473760800, 1473764400, 1473768000, 1473771600, 
    1473775200, 1473778800, 1473782400, 1473786000, 1473789600, 1473793200, 
    1473796800, 1473800400, 1473804000, 1473807600, 1473811200, 1473814800, 
    1473818400, 1473822000, 1473825600, 1473829200, 1473832800, 1473836400, 
    1473840000, 1473843600, 1473847200, 1473850800, 1473854400, 1473858000, 
    1473861600, 1473865200, 1473868800, 1473872400, 1473876000, 1473879600, 
    1473883200, 1473886800, 1473890400, 1473894000, 1473897600, 1473901200, 
    1473904800, 1473908400, 1473912000, 1473915600, 1473919200, 1473922800, 
    1473926400, 1473930000, 1473933600, 1473937200, 1473940800, 1473944400, 
    1473948000, 1473951600, 1473955200, 1473958800, 1473962400, 1473966000, 
    1473969600, 1473973200, 1473976800, 1473980400, 1473984000, 1473987600, 
    1473991200, 1473994800, 1473998400, 1474002000, 1474005600, 1474009200, 
    1474012800, 1474016400, 1474020000, 1474023600, 1474027200, 1474030800, 
    1474034400, 1474038000, 1474041600, 1474045200, 1474048800, 1474052400, 
    1474056000, 1474059600, 1474063200, 1474066800, 1474070400, 1474074000, 
    1474077600, 1474081200, 1474084800, 1474088400, 1474092000, 1474095600, 
    1474099200, 1474102800, 1474106400, 1474110000, 1474113600, 1474117200, 
    1474120800, 1474124400, 1474128000, 1474131600, 1474135200, 1474138800, 
    1474142400, 1474146000, 1474149600, 1474153200, 1474156800, 1474160400, 
    1474164000, 1474167600, 1474171200, 1474174800, 1474178400, 1474182000, 
    1474185600, 1474189200, 1474192800, 1474196400, 1474200000, 1474203600, 
    1474207200, 1474210800, 1474214400, 1474218000, 1474221600, 1474225200, 
    1474228800, 1474232400, 1474236000, 1474239600, 1474243200, 1474246800, 
    1474250400, 1474254000, 1474257600, 1474261200, 1474264800, 1474268400, 
    1474272000, 1474275600, 1474279200, 1474282800, 1474286400, 1474290000, 
    1474293600, 1474297200, 1474300800, 1474304400, 1474308000, 1474311600, 
    1474315200, 1474318800, 1474322400, 1474326000, 1474329600, 1474333200, 
    1474336800, 1474340400, 1474344000, 1474347600, 1474351200, 1474354800, 
    1474358400, 1474362000, 1474365600, 1474369200, 1474372800, 1474376400, 
    1474380000, 1474383600, 1474387200, 1474390800, 1474394400, 1474398000, 
    1474401600, 1474405200, 1474408800, 1474412400, 1474416000, 1474419600, 
    1474423200, 1474426800, 1474430400, 1474434000, 1474437600, 1474441200, 
    1474444800, 1474448400, 1474452000, 1474455600, 1474459200, 1474462800, 
    1474466400, 1474470000, 1474473600, 1474477200, 1474480800, 1474484400, 
    1474488000, 1474491600, 1474495200, 1474498800, 1474502400, 1474506000, 
    1474509600, 1474513200, 1474516800, 1474520400, 1474524000, 1474527600, 
    1474531200, 1474534800, 1474538400, 1474542000, 1474545600, 1474549200, 
    1474552800, 1474556400, 1474560000, 1474563600, 1474567200, 1474570800, 
    1474574400, 1474578000, 1474581600, 1474585200, 1474588800, 1474592400, 
    1474596000, 1474599600, 1474603200, 1474606800, 1474610400, 1474614000, 
    1474617600, 1474621200, 1474624800, 1474628400, 1474632000, 1474635600, 
    1474639200, 1474642800, 1474646400, 1474650000, 1474653600, 1474657200, 
    1474660800, 1474664400, 1474668000, 1474671600, 1474675200, 1474678800, 
    1474682400, 1474686000, 1474689600, 1474693200, 1474696800, 1474700400, 
    1474704000, 1474707600, 1474711200, 1474714800, 1474718400, 1474722000, 
    1474725600, 1474729200, 1474732800, 1474736400, 1474740000, 1474743600, 
    1474747200, 1474750800, 1474754400, 1474758000, 1474761600, 1474765200, 
    1474768800, 1474772400, 1474776000, 1474779600, 1474783200, 1474786800, 
    1474790400, 1474794000, 1474797600, 1474801200, 1474804800, 1474808400, 
    1474812000, 1474815600, 1474819200, 1474822800, 1474826400, 1474830000, 
    1474833600, 1474837200, 1474840800, 1474844400, 1474848000, 1474851600, 
    1474855200, 1474858800, 1474862400, 1474866000, 1474869600, 1474873200, 
    1474876800, 1474880400, 1474884000, 1474887600, 1474891200, 1474894800, 
    1474898400, 1474902000, 1474905600, 1474909200, 1474912800, 1474916400, 
    1474920000, 1474923600, 1474927200, 1474930800, 1474934400, 1474938000, 
    1474941600, 1474945200, 1474948800, 1474952400, 1474956000, 1474959600, 
    1474963200, 1474966800, 1474970400, 1474974000, 1474977600, 1474981200, 
    1474984800, 1474988400, 1474992000, 1474995600, 1474999200, 1475002800, 
    1475006400, 1475010000, 1475013600, 1475017200, 1475020800, 1475024400, 
    1475028000, 1475031600, 1475035200, 1475038800, 1475042400, 1475046000, 
    1475049600, 1475053200, 1475056800, 1475060400, 1475064000, 1475067600, 
    1475071200, 1475074800, 1475078400, 1475082000, 1475085600, 1475089200, 
    1475092800, 1475096400, 1475100000, 1475103600, 1475107200, 1475110800, 
    1475114400, 1475118000, 1475121600, 1475125200, 1475128800, 1475132400, 
    1475136000, 1475139600, 1475143200, 1475146800, 1475150400, 1475154000, 
    1475157600, 1475161200, 1475164800, 1475168400, 1475172000, 1475175600, 
    1475179200, 1475182800, 1475186400, 1475190000, 1475193600, 1475197200, 
    1475200800, 1475204400, 1475208000, 1475211600, 1475215200, 1475218800, 
    1475222400, 1475226000, 1475229600, 1475233200, 1475236800, 1475240400, 
    1475244000, 1475247600, 1475251200, 1475254800, 1475258400, 1475262000, 
    1475265600, 1475269200, 1475272800, 1475276400, 1475280000, 1475283600, 
    1475287200, 1475290800, 1475294400, 1475298000, 1475301600, 1475305200, 
    1475308800, 1475312400, 1475316000, 1475319600, 1475323200, 1475326800, 
    1475330400, 1475334000, 1475337600, 1475341200, 1475344800, 1475348400, 
    1475352000, 1475355600, 1475359200, 1475362800, 1475366400, 1475370000, 
    1475373600, 1475377200, 1475380800, 1475384400, 1475388000, 1475391600, 
    1475395200, 1475398800, 1475402400, 1475406000, 1475409600, 1475413200, 
    1475416800, 1475420400, 1475424000, 1475427600, 1475431200, 1475434800, 
    1475438400, 1475442000, 1475445600, 1475449200, 1475452800, 1475456400, 
    1475460000, 1475463600, 1475467200, 1475470800, 1475474400, 1475478000, 
    1475481600, 1475485200, 1475488800, 1475492400, 1475496000, 1475499600, 
    1475503200, 1475506800, 1475510400, 1475514000, 1475517600, 1475521200, 
    1475524800, 1475528400, 1475532000, 1475535600, 1475539200, 1475542800, 
    1475546400, 1475550000, 1475553600, 1475557200, 1475560800, 1475564400, 
    1475568000, 1475571600, 1475575200, 1475578800, 1475582400, 1475586000, 
    1475589600, 1475593200, 1475596800, 1475600400, 1475604000, 1475607600, 
    1475611200, 1475614800, 1475618400, 1475622000, 1475625600, 1475629200, 
    1475632800, 1475636400, 1475640000, 1475643600, 1475647200, 1475650800, 
    1475654400, 1475658000, 1475661600, 1475665200, 1475668800, 1475672400, 
    1475676000, 1475679600, 1475683200, 1475686800, 1475690400, 1475694000, 
    1475697600, 1475701200, 1475704800, 1475708400, 1475712000, 1475715600, 
    1475719200, 1475722800, 1475726400, 1475730000, 1475733600, 1475737200, 
    1475740800, 1475744400, 1475748000, 1475751600, 1475755200, 1475758800, 
    1475762400, 1475766000, 1475769600, 1475773200, 1475776800, 1475780400, 
    1475784000, 1475787600, 1475791200, 1475794800, 1475798400, 1475802000, 
    1475805600, 1475809200, 1475812800, 1475816400, 1475820000, 1475823600, 
    1475827200, 1475830800, 1475834400, 1475838000, 1475841600, 1475845200, 
    1475848800, 1475852400, 1475856000, 1475859600, 1475863200, 1475866800, 
    1475870400, 1475874000, 1475877600, 1475881200, 1475884800, 1475888400, 
    1475892000, 1475895600, 1475899200, 1475902800, 1475906400, 1475910000, 
    1475913600, 1475917200, 1475920800, 1475924400, 1475928000, 1475931600, 
    1475935200, 1475938800, 1475942400, 1475946000, 1475949600, 1475953200, 
    1475956800, 1475960400, 1475964000, 1475967600, 1475971200, 1475974800, 
    1475978400, 1475982000, 1475985600, 1475989200, 1475992800, 1475996400, 
    1476000000, 1476003600, 1476007200, 1476010800, 1476014400, 1476018000, 
    1476021600, 1476025200, 1476028800, 1476032400, 1476036000, 1476039600, 
    1476043200, 1476046800, 1476050400, 1476054000, 1476057600, 1476061200, 
    1476064800, 1476068400, 1476072000, 1476075600, 1476079200, 1476082800, 
    1476086400, 1476090000, 1476093600, 1476097200, 1476100800, 1476104400, 
    1476108000, 1476111600, 1476115200, 1476118800, 1476122400, 1476126000, 
    1476129600, 1476133200, 1476136800, 1476140400, 1476144000, 1476147600, 
    1476151200, 1476154800, 1476158400, 1476162000, 1476165600, 1476169200, 
    1476172800, 1476176400, 1476180000, 1476183600, 1476187200, 1476190800, 
    1476194400, 1476198000, 1476201600, 1476205200, 1476208800, 1476212400, 
    1476216000, 1476219600, 1476223200, 1476226800, 1476230400, 1476234000, 
    1476237600, 1476241200, 1476244800, 1476248400, 1476252000, 1476255600, 
    1476259200, 1476262800, 1476266400, 1476270000, 1476273600, 1476277200, 
    1476280800, 1476284400, 1476288000, 1476291600, 1476295200, 1476298800, 
    1476302400, 1476306000, 1476309600, 1476313200, 1476316800, 1476320400, 
    1476324000, 1476327600, 1476331200, 1476334800, 1476338400, 1476342000, 
    1476345600, 1476349200, 1476352800, 1476356400, 1476360000, 1476363600, 
    1476367200, 1476370800, 1476374400, 1476378000, 1476381600, 1476385200, 
    1476388800, 1476392400, 1476396000, 1476399600, 1476403200, 1476406800, 
    1476410400, 1476414000, 1476417600, 1476421200, 1476424800, 1476428400, 
    1476432000, 1476435600, 1476439200, 1476442800, 1476446400, 1476450000, 
    1476453600, 1476457200, 1476460800, 1476464400, 1476468000, 1476471600, 
    1476475200, 1476478800, 1476482400, 1476486000, 1476489600, 1476493200, 
    1476496800, 1476500400, 1476504000, 1476507600, 1476511200, 1476514800, 
    1476518400, 1476522000, 1476525600, 1476529200, 1476532800, 1476536400, 
    1476540000, 1476543600, 1476547200, 1476550800, 1476554400, 1476558000, 
    1476561600, 1476565200, 1476568800, 1476572400, 1476576000, 1476579600, 
    1476583200, 1476586800, 1476590400, 1476594000, 1476597600, 1476601200, 
    1476604800, 1476608400, 1476612000, 1476615600, 1476619200, 1476622800, 
    1476626400, 1476630000, 1476633600, 1476637200, 1476640800, 1476644400, 
    1476648000, 1476651600, 1476655200, 1476658800, 1476662400, 1476666000, 
    1476669600, 1476673200, 1476676800, 1476680400, 1476684000, 1476687600, 
    1476691200, 1476694800, 1476698400, 1476702000, 1476705600, 1476709200, 
    1476712800, 1476716400, 1476720000, 1476723600, 1476727200, 1476730800, 
    1476734400, 1476738000, 1476741600, 1476745200, 1476748800, 1476752400, 
    1476756000, 1476759600, 1476763200, 1476766800, 1476770400, 1476774000, 
    1476777600, 1476781200, 1476784800, 1476788400, 1476792000, 1476795600, 
    1476799200, 1476802800, 1476806400, 1476810000, 1476813600, 1476817200, 
    1476820800, 1476824400, 1476828000, 1476831600, 1476835200, 1476838800, 
    1476842400, 1476846000, 1476849600, 1476853200, 1476856800, 1476860400, 
    1476864000, 1476867600, 1476871200, 1476874800, 1476878400, 1476882000, 
    1476885600, 1476889200, 1476892800, 1476896400, 1476900000, 1476903600, 
    1476907200, 1476910800, 1476914400, 1476918000, 1476921600, 1476925200, 
    1476928800, 1476932400, 1476936000, 1476939600, 1476943200, 1476946800, 
    1476950400, 1476954000, 1476957600, 1476961200, 1476964800, 1476968400, 
    1476972000, 1476975600, 1476979200, 1476982800, 1476986400, 1476990000, 
    1476993600, 1476997200, 1477000800, 1477004400, 1477008000, 1477011600, 
    1477015200, 1477018800, 1477022400, 1477026000, 1477029600, 1477033200, 
    1477036800, 1477040400, 1477044000, 1477047600, 1477051200, 1477054800, 
    1477058400, 1477062000, 1477065600, 1477069200, 1477072800, 1477076400, 
    1477080000, 1477083600, 1477087200, 1477090800, 1477094400, 1477098000, 
    1477101600, 1477105200, 1477108800, 1477112400, 1477116000, 1477119600, 
    1477123200, 1477126800, 1477130400, 1477134000, 1477137600, 1477141200, 
    1477144800, 1477148400, 1477152000, 1477155600, 1477159200, 1477162800, 
    1477166400, 1477170000, 1477173600, 1477177200, 1477180800, 1477184400, 
    1477188000, 1477191600, 1477195200, 1477198800, 1477202400, 1477206000, 
    1477209600, 1477213200, 1477216800, 1477220400, 1477224000, 1477227600, 
    1477231200, 1477234800, 1477238400, 1477242000, 1477245600, 1477249200, 
    1477252800, 1477256400, 1477260000, 1477263600, 1477267200, 1477270800, 
    1477274400, 1477278000, 1477281600, 1477285200, 1477288800, 1477292400, 
    1477296000, 1477299600, 1477303200, 1477306800, 1477310400, 1477314000, 
    1477317600, 1477321200, 1477324800, 1477328400, 1477332000, 1477335600, 
    1477339200, 1477342800, 1477346400, 1477350000, 1477353600, 1477357200, 
    1477360800, 1477364400, 1477368000, 1477371600, 1477375200, 1477378800, 
    1477382400, 1477386000, 1477389600, 1477393200, 1477396800, 1477400400, 
    1477404000, 1477407600, 1477411200, 1477414800, 1477418400, 1477422000, 
    1477425600, 1477429200, 1477432800, 1477436400, 1477440000, 1477443600, 
    1477447200, 1477450800, 1477454400, 1477458000, 1477461600, 1477465200, 
    1477468800, 1477472400, 1477476000, 1477479600, 1477483200, 1477486800, 
    1477490400, 1477494000, 1477497600, 1477501200, 1477504800, 1477508400, 
    1477512000, 1477515600, 1477519200, 1477522800, 1477526400, 1477530000, 
    1477533600, 1477537200, 1477540800, 1477544400, 1477548000, 1477551600, 
    1477555200, 1477558800, 1477562400, 1477566000, 1477569600, 1477573200, 
    1477576800, 1477580400, 1477584000, 1477587600, 1477591200, 1477594800, 
    1477598400, 1477602000, 1477605600, 1477609200, 1477612800, 1477616400, 
    1477620000, 1477623600, 1477627200, 1477630800, 1477634400, 1477638000, 
    1477641600, 1477645200, 1477648800, 1477652400, 1477656000, 1477659600, 
    1477663200, 1477666800, 1477670400, 1477674000, 1477677600, 1477681200, 
    1477684800, 1477688400, 1477692000, 1477695600, 1477699200, 1477702800, 
    1477706400, 1477710000, 1477713600, 1477717200, 1477720800, 1477724400, 
    1477728000, 1477731600, 1477735200, 1477738800, 1477742400, 1477746000, 
    1477749600, 1477753200, 1477756800, 1477760400, 1477764000, 1477767600, 
    1477771200, 1477774800, 1477778400, 1477782000, 1477785600, 1477789200, 
    1477792800, 1477796400, 1477800000, 1477803600, 1477807200, 1477810800, 
    1477814400, 1477818000, 1477821600, 1477825200, 1477828800, 1477832400, 
    1477836000, 1477839600, 1477843200, 1477846800, 1477850400, 1477854000, 
    1477857600, 1477861200, 1477864800, 1477868400, 1477872000, 1477875600, 
    1477879200, 1477882800, 1477886400, 1477890000, 1477893600, 1477897200, 
    1477900800, 1477904400, 1477908000, 1477911600, 1477915200, 1477918800, 
    1477922400, 1477926000, 1477929600, 1477933200, 1477936800, 1477940400, 
    1477944000, 1477947600, 1477951200, 1477954800, 1477958400, 1477962000, 
    1477965600, 1477969200, 1477972800, 1477976400, 1477980000, 1477983600, 
    1477987200, 1477990800, 1477994400, 1477998000, 1478001600, 1478005200, 
    1478008800, 1478012400, 1478016000, 1478019600, 1478023200, 1478026800, 
    1478030400, 1478034000, 1478037600, 1478041200, 1478044800, 1478048400, 
    1478052000, 1478055600, 1478059200, 1478062800, 1478066400, 1478070000, 
    1478073600, 1478077200, 1478080800, 1478084400, 1478088000, 1478091600, 
    1478095200, 1478098800, 1478102400, 1478106000, 1478109600, 1478113200, 
    1478116800, 1478120400, 1478124000, 1478127600, 1478131200, 1478134800, 
    1478138400, 1478142000, 1478145600, 1478149200, 1478152800, 1478156400, 
    1478160000, 1478163600, 1478167200, 1478170800, 1478174400, 1478178000, 
    1478181600, 1478185200, 1478188800, 1478192400, 1478196000, 1478199600, 
    1478203200, 1478206800, 1478210400, 1478214000, 1478217600, 1478221200, 
    1478224800, 1478228400, 1478232000, 1478235600, 1478239200, 1478242800, 
    1478246400, 1478250000, 1478253600, 1478257200, 1478260800, 1478264400, 
    1478268000, 1478271600, 1478275200, 1478278800, 1478282400, 1478286000, 
    1478289600, 1478293200, 1478296800, 1478300400, 1478304000, 1478307600, 
    1478311200, 1478314800, 1478318400, 1478322000, 1478325600, 1478329200, 
    1478332800, 1478336400, 1478340000, 1478343600, 1478347200, 1478350800, 
    1478354400, 1478358000, 1478361600, 1478365200, 1478368800, 1478372400, 
    1478376000, 1478379600, 1478383200, 1478386800, 1478390400, 1478394000, 
    1478397600, 1478401200, 1478404800, 1478408400, 1478412000, 1478415600, 
    1478419200, 1478422800, 1478426400, 1478430000, 1478433600, 1478437200, 
    1478440800, 1478444400, 1478448000, 1478451600, 1478455200, 1478458800, 
    1478462400, 1478466000, 1478469600, 1478473200, 1478476800, 1478480400, 
    1478484000, 1478487600, 1478491200, 1478494800, 1478498400, 1478502000, 
    1478505600, 1478509200, 1478512800, 1478516400, 1478520000, 1478523600, 
    1478527200, 1478530800, 1478534400, 1478538000, 1478541600, 1478545200, 
    1478548800, 1478552400, 1478556000, 1478559600, 1478563200, 1478566800, 
    1478570400, 1478574000, 1478577600, 1478581200, 1478584800, 1478588400, 
    1478592000, 1478595600, 1478599200, 1478602800, 1478606400, 1478610000, 
    1478613600, 1478617200, 1478620800, 1478624400, 1478628000, 1478631600, 
    1478635200, 1478638800, 1478642400, 1478646000, 1478649600, 1478653200, 
    1478656800, 1478660400, 1478664000, 1478667600, 1478671200, 1478674800, 
    1478678400, 1478682000, 1478685600, 1478689200, 1478692800, 1478696400, 
    1478700000, 1478703600, 1478707200, 1478710800, 1478714400, 1478718000, 
    1478721600, 1478725200, 1478728800, 1478732400, 1478736000, 1478739600, 
    1478743200, 1478746800, 1478750400, 1478754000, 1478757600, 1478761200, 
    1478764800, 1478768400, 1478772000, 1478775600, 1478779200, 1478782800, 
    1478786400, 1478790000, 1478793600, 1478797200, 1478800800, 1478804400, 
    1478808000, 1478811600, 1478815200, 1478818800, 1478822400, 1478826000, 
    1478829600, 1478833200, 1478836800, 1478840400, 1478844000, 1478847600, 
    1478851200, 1478854800, 1478858400, 1478862000, 1478865600, 1478869200, 
    1478872800, 1478876400, 1478880000, 1478883600, 1478887200, 1478890800, 
    1478894400, 1478898000, 1478901600, 1478905200, 1478908800, 1478912400, 
    1478916000, 1478919600, 1478923200, 1478926800, 1478930400, 1478934000, 
    1478937600, 1478941200, 1478944800, 1478948400, 1478952000, 1478955600, 
    1478959200, 1478962800, 1478966400, 1478970000, 1478973600, 1478977200, 
    1478980800, 1478984400, 1478988000, 1478991600, 1478995200, 1478998800, 
    1479002400, 1479006000, 1479009600, 1479013200, 1479016800, 1479020400, 
    1479024000, 1479027600, 1479031200, 1479034800, 1479038400, 1479042000, 
    1479045600, 1479049200, 1479052800, 1479056400, 1479060000, 1479063600, 
    1479067200, 1479070800, 1479074400, 1479078000, 1479081600, 1479085200, 
    1479088800, 1479092400, 1479096000, 1479099600, 1479103200, 1479106800, 
    1479110400, 1479114000, 1479117600, 1479121200, 1479124800, 1479128400, 
    1479132000, 1479135600, 1479139200, 1479142800, 1479146400, 1479150000, 
    1479153600, 1479157200, 1479160800, 1479164400, 1479168000, 1479171600, 
    1479175200, 1479178800, 1479182400, 1479186000, 1479189600, 1479193200, 
    1479196800, 1479200400, 1479204000, 1479207600, 1479211200, 1479214800, 
    1479218400, 1479222000, 1479225600, 1479229200, 1479232800, 1479236400, 
    1479240000, 1479243600, 1479247200, 1479250800, 1479254400, 1479258000, 
    1479261600, 1479265200, 1479268800, 1479272400, 1479276000, 1479279600, 
    1479283200, 1479286800, 1479290400, 1479294000, 1479297600, 1479301200, 
    1479304800, 1479308400, 1479312000, 1479315600, 1479319200, 1479322800, 
    1479326400, 1479330000, 1479333600, 1479337200, 1479340800, 1479344400, 
    1479348000, 1479351600, 1479355200, 1479358800, 1479362400, 1479366000, 
    1479369600, 1479373200, 1479376800, 1479380400, 1479384000, 1479387600, 
    1479391200, 1479394800, 1479398400, 1479402000, 1479405600, 1479409200, 
    1479412800, 1479416400, 1479420000, 1479423600, 1479427200, 1479430800, 
    1479434400, 1479438000, 1479441600, 1479445200, 1479448800, 1479452400, 
    1479456000, 1479459600, 1479463200, 1479466800, 1479470400, 1479474000, 
    1479477600, 1479481200, 1479484800, 1479488400, 1479492000, 1479495600, 
    1479499200, 1479502800, 1479506400, 1479510000, 1479513600, 1479517200, 
    1479520800, 1479524400, 1479528000, 1479531600, 1479535200, 1479538800, 
    1479542400, 1479546000, 1479549600, 1479553200, 1479556800, 1479560400, 
    1479564000, 1479567600, 1479571200, 1479574800, 1479578400, 1479582000, 
    1479585600, 1479589200, 1479592800, 1479596400, 1479600000, 1479603600, 
    1479607200, 1479610800, 1479614400, 1479618000, 1479621600, 1479625200, 
    1479628800, 1479632400, 1479636000, 1479639600, 1479643200, 1479646800, 
    1479650400, 1479654000, 1479657600, 1479661200, 1479664800, 1479668400, 
    1479672000, 1479675600, 1479679200, 1479682800, 1479686400, 1479690000, 
    1479693600, 1479697200, 1479700800, 1479704400, 1479708000, 1479711600, 
    1479715200, 1479718800, 1479722400, 1479726000, 1479729600, 1479733200, 
    1479736800, 1479740400, 1479744000, 1479747600, 1479751200, 1479754800, 
    1479758400, 1479762000, 1479765600, 1479769200, 1479772800, 1479776400, 
    1479780000, 1479783600, 1479787200, 1479790800, 1479794400, 1479798000, 
    1479801600, 1479805200, 1479808800, 1479812400, 1479816000, 1479819600, 
    1479823200, 1479826800, 1479830400, 1479834000, 1479837600, 1479841200, 
    1479844800, 1479848400, 1479852000, 1479855600, 1479859200, 1479862800, 
    1479866400, 1479870000, 1479873600, 1479877200, 1479880800, 1479884400, 
    1479888000, 1479891600, 1479895200, 1479898800, 1479902400, 1479906000, 
    1479909600, 1479913200, 1479916800, 1479920400, 1479924000, 1479927600, 
    1479931200, 1479934800, 1479938400, 1479942000, 1479945600, 1479949200, 
    1479952800, 1479956400, 1479960000, 1479963600, 1479967200, 1479970800, 
    1479974400, 1479978000, 1479981600, 1479985200, 1479988800, 1479992400, 
    1479996000, 1479999600, 1480003200, 1480006800, 1480010400, 1480014000, 
    1480017600, 1480021200, 1480024800, 1480028400, 1480032000, 1480035600, 
    1480039200, 1480042800, 1480046400, 1480050000, 1480053600, 1480057200, 
    1480060800, 1480064400, 1480068000, 1480071600, 1480075200, 1480078800, 
    1480082400, 1480086000, 1480089600, 1480093200, 1480096800, 1480100400, 
    1480104000, 1480107600, 1480111200, 1480114800, 1480118400, 1480122000, 
    1480125600, 1480129200, 1480132800, 1480136400, 1480140000, 1480143600, 
    1480147200, 1480150800, 1480154400, 1480158000, 1480161600, 1480165200, 
    1480168800, 1480172400, 1480176000, 1480179600, 1480183200, 1480186800, 
    1480190400, 1480194000, 1480197600, 1480201200, 1480204800, 1480208400, 
    1480212000, 1480215600, 1480219200, 1480222800, 1480226400, 1480230000, 
    1480233600, 1480237200, 1480240800, 1480244400, 1480248000, 1480251600, 
    1480255200, 1480258800, 1480262400, 1480266000, 1480269600, 1480273200, 
    1480276800, 1480280400, 1480284000, 1480287600, 1480291200, 1480294800, 
    1480298400, 1480302000, 1480305600, 1480309200, 1480312800, 1480316400, 
    1480320000, 1480323600, 1480327200, 1480330800, 1480334400, 1480338000, 
    1480341600, 1480345200, 1480348800, 1480352400, 1480356000, 1480359600, 
    1480363200, 1480366800, 1480370400, 1480374000, 1480377600, 1480381200, 
    1480384800, 1480388400, 1480392000, 1480395600, 1480399200, 1480402800, 
    1480406400, 1480410000, 1480413600, 1480417200, 1480420800, 1480424400, 
    1480428000, 1480431600, 1480435200, 1480438800, 1480442400, 1480446000, 
    1480449600, 1480453200, 1480456800, 1480460400, 1480464000, 1480467600, 
    1480471200, 1480474800, 1480478400, 1480482000, 1480485600, 1480489200, 
    1480492800, 1480496400, 1480500000, 1480503600, 1480507200, 1480510800, 
    1480514400, 1480518000, 1480521600, 1480525200, 1480528800, 1480532400, 
    1480536000, 1480539600, 1480543200, 1480546800, 1480550400, 1480554000, 
    1480557600, 1480561200, 1480564800, 1480568400, 1480572000, 1480575600, 
    1480579200, 1480582800, 1480586400, 1480590000, 1480593600, 1480597200, 
    1480600800, 1480604400, 1480608000, 1480611600, 1480615200, 1480618800, 
    1480622400, 1480626000, 1480629600, 1480633200, 1480636800, 1480640400, 
    1480644000, 1480647600, 1480651200, 1480654800, 1480658400, 1480662000, 
    1480665600, 1480669200, 1480672800, 1480676400, 1480680000, 1480683600, 
    1480687200, 1480690800, 1480694400, 1480698000, 1480701600, 1480705200, 
    1480708800, 1480712400, 1480716000, 1480719600, 1480723200, 1480726800, 
    1480730400, 1480734000, 1480737600, 1480741200, 1480744800, 1480748400, 
    1480752000, 1480755600, 1480759200, 1480762800, 1480766400, 1480770000, 
    1480773600, 1480777200, 1480780800, 1480784400, 1480788000, 1480791600, 
    1480795200, 1480798800, 1480802400, 1480806000, 1480809600, 1480813200, 
    1480816800, 1480820400, 1480824000, 1480827600, 1480831200, 1480834800, 
    1480838400, 1480842000, 1480845600, 1480849200, 1480852800, 1480856400, 
    1480860000, 1480863600, 1480867200, 1480870800, 1480874400, 1480878000, 
    1480881600, 1480885200, 1480888800, 1480892400, 1480896000, 1480899600, 
    1480903200, 1480906800, 1480910400, 1480914000, 1480917600, 1480921200, 
    1480924800, 1480928400, 1480932000, 1480935600, 1480939200, 1480942800, 
    1480946400, 1480950000, 1480953600, 1480957200, 1480960800, 1480964400, 
    1480968000, 1480971600, 1480975200, 1480978800, 1480982400, 1480986000, 
    1480989600, 1480993200, 1480996800, 1481000400, 1481004000, 1481007600, 
    1481011200, 1481014800, 1481018400, 1481022000, 1481025600, 1481029200, 
    1481032800, 1481036400, 1481040000, 1481043600, 1481047200, 1481050800, 
    1481054400, 1481058000, 1481061600, 1481065200, 1481068800, 1481072400, 
    1481076000, 1481079600, 1481083200, 1481086800, 1481090400, 1481094000, 
    1481097600, 1481101200, 1481104800, 1481108400, 1481112000, 1481115600, 
    1481119200, 1481122800, 1481126400, 1481130000, 1481133600, 1481137200, 
    1481140800, 1481144400, 1481148000, 1481151600, 1481155200, 1481158800, 
    1481162400, 1481166000, 1481169600, 1481173200, 1481176800, 1481180400, 
    1481184000, 1481187600, 1481191200, 1481194800, 1481198400, 1481202000, 
    1481205600, 1481209200, 1481212800, 1481216400, 1481220000, 1481223600, 
    1481227200, 1481230800, 1481234400, 1481238000, 1481241600, 1481245200, 
    1481248800, 1481252400, 1481256000, 1481259600, 1481263200, 1481266800, 
    1481270400, 1481274000, 1481277600, 1481281200, 1481284800, 1481288400, 
    1481292000, 1481295600, 1481299200, 1481302800, 1481306400, 1481310000, 
    1481313600, 1481317200, 1481320800, 1481324400, 1481328000, 1481331600, 
    1481335200, 1481338800, 1481342400, 1481346000, 1481349600, 1481353200, 
    1481356800, 1481360400, 1481364000, 1481367600, 1481371200, 1481374800, 
    1481378400, 1481382000, 1481385600, 1481389200, 1481392800, 1481396400, 
    1481400000, 1481403600, 1481407200, 1481410800, 1481414400, 1481418000, 
    1481421600, 1481425200, 1481428800, 1481432400, 1481436000, 1481439600, 
    1481443200, 1481446800, 1481450400, 1481454000, 1481457600, 1481461200, 
    1481464800, 1481468400, 1481472000, 1481475600, 1481479200, 1481482800, 
    1481486400, 1481490000, 1481493600, 1481497200, 1481500800, 1481504400, 
    1481508000, 1481511600, 1481515200, 1481518800, 1481522400, 1481526000, 
    1481529600, 1481533200, 1481536800, 1481540400, 1481544000, 1481547600, 
    1481551200, 1481554800, 1481558400, 1481562000, 1481565600, 1481569200, 
    1481572800, 1481576400, 1481580000, 1481583600, 1481587200, 1481590800, 
    1481594400, 1481598000, 1481601600, 1481605200, 1481608800, 1481612400, 
    1481616000, 1481619600, 1481623200, 1481626800, 1481630400, 1481634000, 
    1481637600, 1481641200, 1481644800, 1481648400, 1481652000, 1481655600, 
    1481659200, 1481662800, 1481666400, 1481670000, 1481673600, 1481677200, 
    1481680800, 1481684400, 1481688000, 1481691600, 1481695200, 1481698800, 
    1481702400, 1481706000, 1481709600, 1481713200, 1481716800, 1481720400, 
    1481724000, 1481727600, 1481731200, 1481734800, 1481738400, 1481742000, 
    1481745600, 1481749200, 1481752800, 1481756400, 1481760000, 1481763600, 
    1481767200, 1481770800, 1481774400, 1481778000, 1481781600, 1481785200, 
    1481788800, 1481792400, 1481796000, 1481799600, 1481803200, 1481806800, 
    1481810400, 1481814000, 1481817600, 1481821200, 1481824800, 1481828400, 
    1481832000, 1481835600, 1481839200, 1481842800, 1481846400, 1481850000, 
    1481853600, 1481857200, 1481860800, 1481864400, 1481868000, 1481871600, 
    1481875200, 1481878800, 1481882400, 1481886000, 1481889600, 1481893200, 
    1481896800, 1481900400, 1481904000, 1481907600, 1481911200, 1481914800, 
    1481918400, 1481922000, 1481925600, 1481929200, 1481932800, 1481936400, 
    1481940000, 1481943600, 1481947200, 1481950800, 1481954400, 1481958000, 
    1481961600, 1481965200, 1481968800, 1481972400, 1481976000, 1481979600, 
    1481983200, 1481986800, 1481990400, 1481994000, 1481997600, 1482001200, 
    1482004800, 1482008400, 1482012000, 1482015600, 1482019200, 1482022800, 
    1482026400, 1482030000, 1482033600, 1482037200, 1482040800, 1482044400, 
    1482048000, 1482051600, 1482055200, 1482058800, 1482062400, 1482066000, 
    1482069600, 1482073200, 1482076800, 1482080400, 1482084000, 1482087600, 
    1482091200, 1482094800, 1482098400, 1482102000, 1482105600, 1482109200, 
    1482112800, 1482116400, 1482120000, 1482123600, 1482127200, 1482130800, 
    1482134400, 1482138000, 1482141600, 1482145200, 1482148800, 1482152400, 
    1482156000, 1482159600, 1482163200, 1482166800, 1482170400, 1482174000, 
    1482177600, 1482181200, 1482184800, 1482188400, 1482192000, 1482195600, 
    1482199200, 1482202800, 1482206400, 1482210000, 1482213600, 1482217200, 
    1482220800, 1482224400, 1482228000, 1482231600, 1482235200, 1482238800, 
    1482242400, 1482246000, 1482249600, 1482253200, 1482256800, 1482260400, 
    1482264000, 1482267600, 1482271200, 1482274800, 1482278400, 1482282000, 
    1482285600, 1482289200, 1482292800, 1482296400, 1482300000, 1482303600, 
    1482307200, 1482310800, 1482314400, 1482318000, 1482321600, 1482325200, 
    1482328800, 1482332400, 1482336000, 1482339600, 1482343200, 1482346800, 
    1482350400, 1482354000, 1482357600, 1482361200, 1482364800, 1482368400, 
    1482372000, 1482375600, 1482379200, 1482382800, 1482386400, 1482390000, 
    1482393600, 1482397200, 1482400800, 1482404400, 1482408000, 1482411600, 
    1482415200, 1482418800, 1482422400, 1482426000, 1482429600, 1482433200, 
    1482436800, 1482440400, 1482444000, 1482447600, 1482451200, 1482454800, 
    1482458400, 1482462000, 1482465600, 1482469200, 1482472800, 1482476400, 
    1482480000, 1482483600, 1482487200, 1482490800, 1482494400, 1482498000, 
    1482501600, 1482505200, 1482508800, 1482512400, 1482516000, 1482519600, 
    1482523200, 1482526800, 1482530400, 1482534000, 1482537600, 1482541200, 
    1482544800, 1482548400, 1482552000, 1482555600, 1482559200, 1482562800, 
    1482566400, 1482570000, 1482573600, 1482577200, 1482580800, 1482584400, 
    1482588000, 1482591600, 1482595200, 1482598800, 1482602400, 1482606000, 
    1482609600, 1482613200, 1482616800, 1482620400, 1482624000, 1482627600, 
    1482631200, 1482634800, 1482638400, 1482642000, 1482645600, 1482649200, 
    1482652800, 1482656400, 1482660000, 1482663600, 1482667200, 1482670800, 
    1482674400, 1482678000, 1482681600, 1482685200, 1482688800, 1482692400, 
    1482696000, 1482699600, 1482703200, 1482706800, 1482710400, 1482714000, 
    1482717600, 1482721200, 1482724800, 1482728400, 1482732000, 1482735600, 
    1482739200, 1482742800, 1482746400, 1482750000, 1482753600, 1482757200, 
    1482760800, 1482764400, 1482768000, 1482771600, 1482775200, 1482778800, 
    1482782400, 1482786000, 1482789600, 1482793200, 1482796800, 1482800400, 
    1482804000, 1482807600, 1482811200, 1482814800, 1482818400, 1482822000, 
    1482825600, 1482829200, 1482832800, 1482836400, 1482840000, 1482843600, 
    1482847200, 1482850800, 1482854400, 1482858000, 1482861600, 1482865200, 
    1482868800, 1482872400, 1482876000, 1482879600, 1482883200, 1482886800, 
    1482890400, 1482894000, 1482897600, 1482901200, 1482904800, 1482908400, 
    1482912000, 1482915600, 1482919200, 1482922800, 1482926400, 1482930000, 
    1482933600, 1482937200, 1482940800, 1482944400, 1482948000, 1482951600, 
    1482955200, 1482958800, 1482962400, 1482966000, 1482969600, 1482973200, 
    1482976800, 1482980400, 1482984000, 1482987600, 1482991200, 1482994800, 
    1482998400, 1483002000, 1483005600, 1483009200, 1483012800, 1483016400, 
    1483020000, 1483023600, 1483027200, 1483030800, 1483034400, 1483038000, 
    1483041600, 1483045200, 1483048800, 1483052400, 1483056000, 1483059600, 
    1483063200, 1483066800, 1483070400, 1483074000, 1483077600, 1483081200, 
    1483084800, 1483088400, 1483092000, 1483095600, 1483099200, 1483102800, 
    1483106400, 1483110000, 1483113600, 1483117200, 1483120800, 1483124400, 
    1483128000, 1483131600, 1483135200, 1483138800, 1483142400, 1483146000, 
    1483149600, 1483153200, 1483156800, 1483160400, 1483164000, 1483167600, 
    1483171200, 1483174800, 1483178400, 1483182000, 1483185600, 1483189200, 
    1483192800, 1483196400, 1483200000, 1483203600, 1483207200, 1483210800, 
    1483214400, 1483218000, 1483221600, 1483225200, 1483228800, 1483232400, 
    1483236000, 1483239600, 1483243200, 1483246800, 1483250400, 1483254000, 
    1483257600, 1483261200, 1483264800, 1483268400, 1483272000, 1483275600, 
    1483279200, 1483282800, 1483286400, 1483290000, 1483293600, 1483297200, 
    1483300800, 1483304400, 1483308000, 1483311600, 1483315200, 1483318800, 
    1483322400, 1483326000, 1483329600, 1483333200, 1483336800, 1483340400, 
    1483344000, 1483347600, 1483351200, 1483354800, 1483358400, 1483362000, 
    1483365600, 1483369200, 1483372800, 1483376400, 1483380000, 1483383600, 
    1483387200, 1483390800, 1483394400, 1483398000, 1483401600, 1483405200, 
    1483408800, 1483412400, 1483416000, 1483419600, 1483423200, 1483426800, 
    1483430400, 1483434000, 1483437600, 1483441200, 1483444800, 1483448400, 
    1483452000, 1483455600, 1483459200, 1483462800, 1483466400, 1483470000, 
    1483473600, 1483477200, 1483480800, 1483484400, 1483488000, 1483491600, 
    1483495200, 1483498800, 1483502400, 1483506000, 1483509600, 1483513200, 
    1483516800, 1483520400, 1483524000, 1483527600, 1483531200, 1483534800, 
    1483538400, 1483542000, 1483545600, 1483549200, 1483552800, 1483556400, 
    1483560000, 1483563600, 1483567200, 1483570800, 1483574400, 1483578000, 
    1483581600, 1483585200, 1483588800, 1483592400, 1483596000, 1483599600, 
    1483603200, 1483606800, 1483610400, 1483614000, 1483617600, 1483621200, 
    1483624800, 1483628400, 1483632000, 1483635600, 1483639200, 1483642800, 
    1483646400, 1483650000, 1483653600, 1483657200, 1483660800, 1483664400, 
    1483668000, 1483671600, 1483675200, 1483678800, 1483682400, 1483686000, 
    1483689600, 1483693200, 1483696800, 1483700400, 1483704000, 1483707600, 
    1483711200, 1483714800, 1483718400, 1483722000, 1483725600, 1483729200, 
    1483732800, 1483736400, 1483740000, 1483743600, 1483747200, 1483750800, 
    1483754400, 1483758000, 1483761600, 1483765200, 1483768800, 1483772400, 
    1483776000, 1483779600, 1483783200, 1483786800, 1483790400, 1483794000, 
    1483797600, 1483801200, 1483804800, 1483808400, 1483812000, 1483815600, 
    1483819200, 1483822800, 1483826400, 1483830000, 1483833600, 1483837200, 
    1483840800, 1483844400, 1483848000, 1483851600, 1483855200, 1483858800, 
    1483862400, 1483866000, 1483869600, 1483873200, 1483876800, 1483880400, 
    1483884000, 1483887600, 1483891200, 1483894800, 1483898400, 1483902000, 
    1483905600, 1483909200, 1483912800, 1483916400, 1483920000, 1483923600, 
    1483927200, 1483930800, 1483934400, 1483938000, 1483941600, 1483945200, 
    1483948800, 1483952400, 1483956000, 1483959600, 1483963200, 1483966800, 
    1483970400, 1483974000, 1483977600, 1483981200, 1483984800, 1483988400, 
    1483992000, 1483995600, 1483999200, 1484002800, 1484006400, 1484010000, 
    1484013600, 1484017200, 1484020800, 1484024400, 1484028000, 1484031600, 
    1484035200, 1484038800, 1484042400, 1484046000, 1484049600, 1484053200, 
    1484056800, 1484060400, 1484064000, 1484067600, 1484071200, 1484074800, 
    1484078400, 1484082000, 1484085600, 1484089200, 1484092800, 1484096400, 
    1484100000, 1484103600, 1484107200, 1484110800, 1484114400, 1484118000, 
    1484121600, 1484125200, 1484128800, 1484132400, 1484136000, 1484139600, 
    1484143200, 1484146800, 1484150400, 1484154000, 1484157600, 1484161200, 
    1484164800, 1484168400, 1484172000, 1484175600, 1484179200, 1484182800, 
    1484186400, 1484190000, 1484193600, 1484197200, 1484200800, 1484204400, 
    1484208000, 1484211600, 1484215200, 1484218800, 1484222400, 1484226000, 
    1484229600, 1484233200, 1484236800, 1484240400, 1484244000, 1484247600, 
    1484251200, 1484254800, 1484258400, 1484262000, 1484265600, 1484269200, 
    1484272800, 1484276400, 1484280000, 1484283600, 1484287200, 1484290800, 
    1484294400, 1484298000, 1484301600, 1484305200, 1484308800, 1484312400, 
    1484316000, 1484319600, 1484323200, 1484326800, 1484330400, 1484334000, 
    1484337600, 1484341200, 1484344800, 1484348400, 1484352000, 1484355600, 
    1484359200, 1484362800, 1484366400, 1484370000, 1484373600, 1484377200, 
    1484380800, 1484384400, 1484388000, 1484391600, 1484395200, 1484398800, 
    1484402400, 1484406000, 1484409600, 1484413200, 1484416800, 1484420400, 
    1484424000, 1484427600, 1484431200, 1484434800, 1484438400, 1484442000, 
    1484445600, 1484449200, 1484452800, 1484456400, 1484460000, 1484463600, 
    1484467200, 1484470800, 1484474400, 1484478000, 1484481600, 1484485200, 
    1484488800, 1484492400, 1484496000, 1484499600, 1484503200, 1484506800, 
    1484510400, 1484514000, 1484517600, 1484521200, 1484524800, 1484528400, 
    1484532000, 1484535600, 1484539200, 1484542800, 1484546400, 1484550000, 
    1484553600, 1484557200, 1484560800, 1484564400, 1484568000, 1484571600, 
    1484575200, 1484578800, 1484582400, 1484586000, 1484589600, 1484593200, 
    1484596800, 1484600400, 1484604000, 1484607600, 1484611200, 1484614800, 
    1484618400, 1484622000, 1484625600, 1484629200, 1484632800, 1484636400, 
    1484640000, 1484643600, 1484647200, 1484650800, 1484654400, 1484658000, 
    1484661600, 1484665200, 1484668800, 1484672400, 1484676000, 1484679600, 
    1484683200, 1484686800, 1484690400, 1484694000, 1484697600, 1484701200, 
    1484704800, 1484708400, 1484712000, 1484715600, 1484719200, 1484722800, 
    1484726400, 1484730000, 1484733600, 1484737200, 1484740800, 1484744400, 
    1484748000, 1484751600, 1484755200, 1484758800, 1484762400, 1484766000, 
    1484769600, 1484773200, 1484776800, 1484780400, 1484784000, 1484787600, 
    1484791200, 1484794800, 1484798400, 1484802000, 1484805600, 1484809200, 
    1484812800, 1484816400, 1484820000, 1484823600, 1484827200, 1484830800, 
    1484834400, 1484838000, 1484841600, 1484845200, 1484848800, 1484852400, 
    1484856000, 1484859600, 1484863200, 1484866800, 1484870400, 1484874000, 
    1484877600, 1484881200, 1484884800, 1484888400, 1484892000, 1484895600, 
    1484899200, 1484902800, 1484906400, 1484910000, 1484913600, 1484917200, 
    1484920800, 1484924400, 1484928000, 1484931600, 1484935200, 1484938800, 
    1484942400, 1484946000, 1484949600, 1484953200, 1484956800, 1484960400, 
    1484964000, 1484967600, 1484971200, 1484974800, 1484978400, 1484982000, 
    1484985600, 1484989200, 1484992800, 1484996400, 1485000000, 1485003600, 
    1485007200, 1485010800, 1485014400, 1485018000, 1485021600, 1485025200, 
    1485028800, 1485032400, 1485036000, 1485039600, 1485043200, 1485046800, 
    1485050400, 1485054000, 1485057600, 1485061200, 1485064800, 1485068400, 
    1485072000, 1485075600, 1485079200, 1485082800, 1485086400, 1485090000, 
    1485093600, 1485097200, 1485100800, 1485104400, 1485108000, 1485111600, 
    1485115200, 1485118800, 1485122400, 1485126000, 1485129600, 1485133200, 
    1485136800, 1485140400, 1485144000, 1485147600, 1485151200, 1485154800, 
    1485158400, 1485162000, 1485165600, 1485169200, 1485172800, 1485176400, 
    1485180000, 1485183600, 1485187200, 1485190800, 1485194400, 1485198000, 
    1485201600, 1485205200, 1485208800, 1485212400, 1485216000, 1485219600, 
    1485223200, 1485226800, 1485230400, 1485234000, 1485237600, 1485241200, 
    1485244800, 1485248400, 1485252000, 1485255600, 1485259200, 1485262800, 
    1485266400, 1485270000, 1485273600, 1485277200, 1485280800, 1485284400, 
    1485288000, 1485291600, 1485295200, 1485298800, 1485302400, 1485306000, 
    1485309600, 1485313200, 1485316800, 1485320400, 1485324000, 1485327600, 
    1485331200, 1485334800, 1485338400, 1485342000, 1485345600, 1485349200, 
    1485352800, 1485356400, 1485360000, 1485363600, 1485367200, 1485370800, 
    1485374400, 1485378000, 1485381600, 1485385200, 1485388800, 1485392400, 
    1485396000, 1485399600, 1485403200, 1485406800, 1485410400, 1485414000, 
    1485417600, 1485421200, 1485424800, 1485428400, 1485432000, 1485435600, 
    1485439200, 1485442800, 1485446400, 1485450000, 1485453600, 1485457200, 
    1485460800, 1485464400, 1485468000, 1485471600, 1485475200, 1485478800, 
    1485482400, 1485486000, 1485489600, 1485493200, 1485496800, 1485500400, 
    1485504000, 1485507600, 1485511200, 1485514800, 1485518400, 1485522000, 
    1485525600, 1485529200, 1485532800, 1485536400, 1485540000, 1485543600, 
    1485547200, 1485550800, 1485554400, 1485558000, 1485561600, 1485565200, 
    1485568800, 1485572400, 1485576000, 1485579600, 1485583200, 1485586800, 
    1485590400, 1485594000, 1485597600, 1485601200, 1485604800, 1485608400, 
    1485612000, 1485615600, 1485619200, 1485622800, 1485626400, 1485630000, 
    1485633600, 1485637200, 1485640800, 1485644400, 1485648000, 1485651600, 
    1485655200, 1485658800, 1485662400, 1485666000, 1485669600, 1485673200, 
    1485676800, 1485680400, 1485684000, 1485687600, 1485691200, 1485694800, 
    1485698400, 1485702000, 1485705600, 1485709200, 1485712800, 1485716400, 
    1485720000, 1485723600, 1485727200, 1485730800, 1485734400, 1485738000, 
    1485741600, 1485745200, 1485748800, 1485752400, 1485756000, 1485759600, 
    1485763200, 1485766800, 1485770400, 1485774000, 1485777600, 1485781200, 
    1485784800, 1485788400, 1485792000, 1485795600, 1485799200, 1485802800, 
    1485806400, 1485810000, 1485813600, 1485817200, 1485820800, 1485824400, 
    1485828000, 1485831600, 1485835200, 1485838800, 1485842400, 1485846000, 
    1485849600, 1485853200, 1485856800, 1485860400, 1485864000, 1485867600, 
    1485871200, 1485874800, 1485878400, 1485882000, 1485885600, 1485889200, 
    1485892800, 1485896400, 1485900000, 1485903600, 1485907200, 1485910800, 
    1485914400, 1485918000, 1485921600, 1485925200, 1485928800, 1485932400, 
    1485936000, 1485939600, 1485943200, 1485946800, 1485950400, 1485954000, 
    1485957600, 1485961200, 1485964800, 1485968400, 1485972000, 1485975600, 
    1485979200, 1485982800, 1485986400, 1485990000, 1485993600, 1485997200, 
    1486000800, 1486004400, 1486008000, 1486011600, 1486015200, 1486018800, 
    1486022400, 1486026000, 1486029600, 1486033200, 1486036800, 1486040400, 
    1486044000, 1486047600, 1486051200, 1486054800, 1486058400, 1486062000, 
    1486065600, 1486069200, 1486072800, 1486076400, 1486080000, 1486083600, 
    1486087200, 1486090800, 1486094400, 1486098000, 1486101600, 1486105200, 
    1486108800, 1486112400, 1486116000, 1486119600, 1486123200, 1486126800, 
    1486130400, 1486134000, 1486137600, 1486141200, 1486144800, 1486148400, 
    1486152000, 1486155600, 1486159200, 1486162800, 1486166400, 1486170000, 
    1486173600, 1486177200, 1486180800, 1486184400, 1486188000, 1486191600, 
    1486195200, 1486198800, 1486202400, 1486206000, 1486209600, 1486213200, 
    1486216800, 1486220400, 1486224000, 1486227600, 1486231200, 1486234800, 
    1486238400, 1486242000, 1486245600, 1486249200, 1486252800, 1486256400, 
    1486260000, 1486263600, 1486267200, 1486270800, 1486274400, 1486278000, 
    1486281600, 1486285200, 1486288800, 1486292400, 1486296000, 1486299600, 
    1486303200, 1486306800, 1486310400, 1486314000, 1486317600, 1486321200, 
    1486324800, 1486328400, 1486332000, 1486335600, 1486339200, 1486342800, 
    1486346400, 1486350000, 1486353600, 1486357200, 1486360800, 1486364400, 
    1486368000, 1486371600, 1486375200, 1486378800, 1486382400, 1486386000, 
    1486389600, 1486393200, 1486396800, 1486400400, 1486404000, 1486407600, 
    1486411200, 1486414800, 1486418400, 1486422000, 1486425600, 1486429200, 
    1486432800, 1486436400, 1486440000, 1486443600, 1486447200, 1486450800, 
    1486454400, 1486458000, 1486461600, 1486465200, 1486468800, 1486472400, 
    1486476000, 1486479600, 1486483200, 1486486800, 1486490400, 1486494000, 
    1486497600, 1486501200, 1486504800, 1486508400, 1486512000, 1486515600, 
    1486519200, 1486522800, 1486526400, 1486530000, 1486533600, 1486537200, 
    1486540800, 1486544400, 1486548000, 1486551600, 1486555200, 1486558800, 
    1486562400, 1486566000, 1486569600, 1486573200, 1486576800, 1486580400, 
    1486584000, 1486587600, 1486591200, 1486594800, 1486598400, 1486602000, 
    1486605600, 1486609200, 1486612800, 1486616400, 1486620000, 1486623600, 
    1486627200, 1486630800, 1486634400, 1486638000, 1486641600, 1486645200, 
    1486648800, 1486652400, 1486656000, 1486659600, 1486663200, 1486666800, 
    1486670400, 1486674000, 1486677600, 1486681200, 1486684800, 1486688400, 
    1486692000, 1486695600, 1486699200, 1486702800, 1486706400, 1486710000, 
    1486713600, 1486717200, 1486720800, 1486724400, 1486728000, 1486731600, 
    1486735200, 1486738800, 1486742400, 1486746000, 1486749600, 1486753200, 
    1486756800, 1486760400, 1486764000, 1486767600, 1486771200, 1486774800, 
    1486778400, 1486782000, 1486785600, 1486789200, 1486792800, 1486796400, 
    1486800000, 1486803600, 1486807200, 1486810800, 1486814400, 1486818000, 
    1486821600, 1486825200, 1486828800, 1486832400, 1486836000, 1486839600, 
    1486843200, 1486846800, 1486850400, 1486854000, 1486857600, 1486861200, 
    1486864800, 1486868400, 1486872000, 1486875600, 1486879200, 1486882800, 
    1486886400, 1486890000, 1486893600, 1486897200, 1486900800, 1486904400, 
    1486908000, 1486911600, 1486915200, 1486918800, 1486922400, 1486926000, 
    1486929600, 1486933200, 1486936800, 1486940400, 1486944000, 1486947600, 
    1486951200, 1486954800, 1486958400, 1486962000, 1486965600, 1486969200, 
    1486972800, 1486976400, 1486980000, 1486983600, 1486987200, 1486990800, 
    1486994400, 1486998000, 1487001600, 1487005200, 1487008800, 1487012400, 
    1487016000, 1487019600, 1487023200, 1487026800, 1487030400, 1487034000, 
    1487037600, 1487041200, 1487044800, 1487048400, 1487052000, 1487055600, 
    1487059200, 1487062800, 1487066400, 1487070000, 1487073600, 1487077200, 
    1487080800, 1487084400, 1487088000, 1487091600, 1487095200, 1487098800, 
    1487102400, 1487106000, 1487109600, 1487113200, 1487116800, 1487120400, 
    1487124000, 1487127600, 1487131200, 1487134800, 1487138400, 1487142000, 
    1487145600, 1487149200, 1487152800, 1487156400, 1487160000, 1487163600, 
    1487167200, 1487170800, 1487174400, 1487178000, 1487181600, 1487185200, 
    1487188800, 1487192400, 1487196000, 1487199600, 1487203200, 1487206800, 
    1487210400, 1487214000, 1487217600, 1487221200, 1487224800, 1487228400, 
    1487232000, 1487235600, 1487239200, 1487242800, 1487246400, 1487250000, 
    1487253600, 1487257200, 1487260800, 1487264400, 1487268000, 1487271600, 
    1487275200, 1487278800, 1487282400, 1487286000, 1487289600, 1487293200, 
    1487296800, 1487300400, 1487304000, 1487307600, 1487311200, 1487314800, 
    1487318400, 1487322000, 1487325600, 1487329200, 1487332800, 1487336400, 
    1487340000, 1487343600, 1487347200, 1487350800, 1487354400, 1487358000, 
    1487361600, 1487365200, 1487368800, 1487372400, 1487376000, 1487379600, 
    1487383200, 1487386800, 1487390400, 1487394000, 1487397600, 1487401200, 
    1487404800, 1487408400, 1487412000, 1487415600, 1487419200, 1487422800, 
    1487426400, 1487430000, 1487433600, 1487437200, 1487440800, 1487444400, 
    1487448000, 1487451600, 1487455200, 1487458800, 1487462400, 1487466000, 
    1487469600, 1487473200, 1487476800, 1487480400, 1487484000, 1487487600, 
    1487491200, 1487494800, 1487498400, 1487502000, 1487505600, 1487509200, 
    1487512800, 1487516400, 1487520000, 1487523600, 1487527200, 1487530800, 
    1487534400, 1487538000, 1487541600, 1487545200, 1487548800, 1487552400, 
    1487556000, 1487559600, 1487563200, 1487566800, 1487570400, 1487574000, 
    1487577600, 1487581200, 1487584800, 1487588400, 1487592000, 1487595600, 
    1487599200, 1487602800, 1487606400, 1487610000, 1487613600, 1487617200, 
    1487620800, 1487624400, 1487628000, 1487631600, 1487635200, 1487638800, 
    1487642400, 1487646000, 1487649600, 1487653200, 1487656800, 1487660400, 
    1487664000, 1487667600, 1487671200, 1487674800, 1487678400, 1487682000, 
    1487685600, 1487689200, 1487692800, 1487696400, 1487700000, 1487703600, 
    1487707200, 1487710800, 1487714400, 1487718000, 1487721600, 1487725200, 
    1487728800, 1487732400, 1487736000, 1487739600, 1487743200, 1487746800, 
    1487750400, 1487754000, 1487757600, 1487761200, 1487764800, 1487768400, 
    1487772000, 1487775600, 1487779200, 1487782800, 1487786400, 1487790000, 
    1487793600, 1487797200, 1487800800, 1487804400, 1487808000, 1487811600, 
    1487815200, 1487818800, 1487822400, 1487826000, 1487829600, 1487833200, 
    1487836800, 1487840400, 1487844000, 1487847600, 1487851200, 1487854800, 
    1487858400, 1487862000, 1487865600, 1487869200, 1487872800, 1487876400, 
    1487880000, 1487883600, 1487887200, 1487890800, 1487894400, 1487898000, 
    1487901600, 1487905200, 1487908800, 1487912400, 1487916000, 1487919600, 
    1487923200, 1487926800, 1487930400, 1487934000, 1487937600, 1487941200, 
    1487944800, 1487948400, 1487952000, 1487955600, 1487959200, 1487962800, 
    1487966400, 1487970000, 1487973600, 1487977200, 1487980800, 1487984400, 
    1487988000, 1487991600, 1487995200, 1487998800, 1488002400, 1488006000, 
    1488009600, 1488013200, 1488016800, 1488020400, 1488024000, 1488027600, 
    1488031200, 1488034800, 1488038400, 1488042000, 1488045600, 1488049200, 
    1488052800, 1488056400, 1488060000, 1488063600, 1488067200, 1488070800, 
    1488074400, 1488078000, 1488081600, 1488085200, 1488088800, 1488092400, 
    1488096000, 1488099600, 1488103200, 1488106800, 1488110400, 1488114000, 
    1488117600, 1488121200, 1488124800, 1488128400, 1488132000, 1488135600, 
    1488139200, 1488142800, 1488146400, 1488150000, 1488153600, 1488157200, 
    1488160800, 1488164400, 1488168000, 1488171600, 1488175200, 1488178800, 
    1488182400, 1488186000, 1488189600, 1488193200, 1488196800, 1488200400, 
    1488204000, 1488207600, 1488211200, 1488214800, 1488218400, 1488222000, 
    1488225600, 1488229200, 1488232800, 1488236400, 1488240000, 1488243600, 
    1488247200, 1488250800, 1488254400, 1488258000, 1488261600, 1488265200, 
    1488268800, 1488272400, 1488276000, 1488279600, 1488283200, 1488286800, 
    1488290400, 1488294000, 1488297600, 1488301200, 1488304800, 1488308400, 
    1488312000, 1488315600, 1488319200, 1488322800, 1488326400, 1488330000, 
    1488333600, 1488337200, 1488340800, 1488344400, 1488348000, 1488351600, 
    1488355200, 1488358800, 1488362400, 1488366000, 1488369600, 1488373200, 
    1488376800, 1488380400, 1488384000, 1488387600, 1488391200, 1488394800, 
    1488398400, 1488402000, 1488405600, 1488409200, 1488412800, 1488416400, 
    1488420000, 1488423600, 1488427200, 1488430800, 1488434400, 1488438000, 
    1488441600, 1488445200, 1488448800, 1488452400, 1488456000, 1488459600, 
    1488463200, 1488466800, 1488470400, 1488474000, 1488477600, 1488481200, 
    1488484800, 1488488400, 1488492000, 1488495600, 1488499200, 1488502800, 
    1488506400, 1488510000, 1488513600, 1488517200, 1488520800, 1488524400, 
    1488528000, 1488531600, 1488535200, 1488538800, 1488542400, 1488546000, 
    1488549600, 1488553200, 1488556800, 1488560400, 1488564000, 1488567600, 
    1488571200, 1488574800, 1488578400, 1488582000, 1488585600, 1488589200, 
    1488592800, 1488596400, 1488600000, 1488603600, 1488607200, 1488610800, 
    1488614400, 1488618000, 1488621600, 1488625200, 1488628800, 1488632400, 
    1488636000, 1488639600, 1488643200, 1488646800, 1488650400, 1488654000, 
    1488657600, 1488661200, 1488664800, 1488668400, 1488672000, 1488675600, 
    1488679200, 1488682800, 1488686400, 1488690000, 1488693600, 1488697200, 
    1488700800, 1488704400, 1488708000, 1488711600, 1488715200, 1488718800, 
    1488722400, 1488726000, 1488729600, 1488733200, 1488736800, 1488740400, 
    1488744000, 1488747600, 1488751200, 1488754800, 1488758400, 1488762000, 
    1488765600, 1488769200, 1488772800, 1488776400, 1488780000, 1488783600, 
    1488787200, 1488790800, 1488794400, 1488798000, 1488801600, 1488805200, 
    1488808800, 1488812400, 1488816000, 1488819600, 1488823200, 1488826800, 
    1488830400, 1488834000, 1488837600, 1488841200, 1488844800, 1488848400, 
    1488852000, 1488855600, 1488859200, 1488862800, 1488866400, 1488870000, 
    1488873600, 1488877200, 1488880800, 1488884400, 1488888000, 1488891600, 
    1488895200, 1488898800, 1488902400, 1488906000, 1488909600, 1488913200, 
    1488916800, 1488920400, 1488924000, 1488927600, 1488931200, 1488934800, 
    1488938400, 1488942000, 1488945600, 1488949200, 1488952800, 1488956400, 
    1488960000, 1488963600, 1488967200, 1488970800, 1488974400, 1488978000, 
    1488981600, 1488985200, 1488988800, 1488992400, 1488996000, 1488999600, 
    1489003200, 1489006800, 1489010400, 1489014000, 1489017600, 1489021200, 
    1489024800, 1489028400, 1489032000, 1489035600, 1489039200, 1489042800, 
    1489046400, 1489050000, 1489053600, 1489057200, 1489060800, 1489064400, 
    1489068000, 1489071600, 1489075200, 1489078800, 1489082400, 1489086000, 
    1489089600, 1489093200, 1489096800, 1489100400, 1489104000, 1489107600, 
    1489111200, 1489114800, 1489118400, 1489122000, 1489125600, 1489129200, 
    1489132800, 1489136400, 1489140000, 1489143600, 1489147200, 1489150800, 
    1489154400, 1489158000, 1489161600, 1489165200, 1489168800, 1489172400, 
    1489176000, 1489179600, 1489183200, 1489186800, 1489190400, 1489194000, 
    1489197600, 1489201200, 1489204800, 1489208400, 1489212000, 1489215600, 
    1489219200, 1489222800, 1489226400, 1489230000, 1489233600, 1489237200, 
    1489240800, 1489244400, 1489248000, 1489251600, 1489255200, 1489258800, 
    1489262400, 1489266000, 1489269600, 1489273200, 1489276800, 1489280400, 
    1489284000, 1489287600, 1489291200, 1489294800, 1489298400, 1489302000, 
    1489305600, 1489309200, 1489312800, 1489316400, 1489320000, 1489323600, 
    1489327200, 1489330800, 1489334400, 1489338000, 1489341600, 1489345200, 
    1489348800, 1489352400, 1489356000, 1489359600, 1489363200, 1489366800, 
    1489370400, 1489374000, 1489377600, 1489381200, 1489384800, 1489388400, 
    1489392000, 1489395600, 1489399200, 1489402800, 1489406400, 1489410000, 
    1489413600, 1489417200, 1489420800, 1489424400, 1489428000, 1489431600, 
    1489435200, 1489438800, 1489442400, 1489446000, 1489449600, 1489453200, 
    1489456800, 1489460400, 1489464000, 1489467600, 1489471200, 1489474800, 
    1489478400, 1489482000, 1489485600, 1489489200, 1489492800, 1489496400, 
    1489500000, 1489503600, 1489507200, 1489510800, 1489514400, 1489518000, 
    1489521600, 1489525200, 1489528800, 1489532400, 1489536000, 1489539600, 
    1489543200, 1489546800, 1489550400, 1489554000, 1489557600, 1489561200, 
    1489564800, 1489568400, 1489572000, 1489575600, 1489579200, 1489582800, 
    1489586400, 1489590000, 1489593600, 1489597200, 1489600800, 1489604400, 
    1489608000, 1489611600, 1489615200, 1489618800, 1489622400, 1489626000, 
    1489629600, 1489633200, 1489636800, 1489640400, 1489644000, 1489647600, 
    1489651200, 1489654800, 1489658400, 1489662000, 1489665600, 1489669200, 
    1489672800, 1489676400, 1489680000, 1489683600, 1489687200, 1489690800, 
    1489694400, 1489698000, 1489701600, 1489705200, 1489708800, 1489712400, 
    1489716000, 1489719600, 1489723200, 1489726800, 1489730400, 1489734000, 
    1489737600, 1489741200, 1489744800, 1489748400, 1489752000, 1489755600, 
    1489759200, 1489762800, 1489766400, 1489770000, 1489773600, 1489777200, 
    1489780800, 1489784400, 1489788000, 1489791600, 1489795200, 1489798800, 
    1489802400, 1489806000, 1489809600, 1489813200, 1489816800, 1489820400, 
    1489824000, 1489827600, 1489831200, 1489834800, 1489838400, 1489842000, 
    1489845600, 1489849200, 1489852800, 1489856400, 1489860000, 1489863600, 
    1489867200, 1489870800, 1489874400, 1489878000, 1489881600, 1489885200, 
    1489888800, 1489892400, 1489896000, 1489899600, 1489903200, 1489906800, 
    1489910400, 1489914000, 1489917600, 1489921200, 1489924800, 1489928400, 
    1489932000, 1489935600, 1489939200, 1489942800, 1489946400, 1489950000, 
    1489953600, 1489957200, 1489960800, 1489964400, 1489968000, 1489971600, 
    1489975200, 1489978800, 1489982400, 1489986000, 1489989600, 1489993200, 
    1489996800, 1490000400, 1490004000, 1490007600, 1490011200, 1490014800, 
    1490018400, 1490022000, 1490025600, 1490029200, 1490032800, 1490036400, 
    1490040000, 1490043600, 1490047200, 1490050800, 1490054400, 1490058000, 
    1490061600, 1490065200, 1490068800, 1490072400, 1490076000, 1490079600, 
    1490083200, 1490086800, 1490090400, 1490094000, 1490097600, 1490101200, 
    1490104800, 1490108400, 1490112000, 1490115600, 1490119200, 1490122800, 
    1490126400, 1490130000, 1490133600, 1490137200, 1490140800, 1490144400, 
    1490148000, 1490151600, 1490155200, 1490158800, 1490162400, 1490166000, 
    1490169600, 1490173200, 1490176800, 1490180400, 1490184000, 1490187600, 
    1490191200, 1490194800, 1490198400, 1490202000, 1490205600, 1490209200, 
    1490212800, 1490216400, 1490220000, 1490223600, 1490227200, 1490230800, 
    1490234400, 1490238000, 1490241600, 1490245200, 1490248800, 1490252400, 
    1490256000, 1490259600, 1490263200, 1490266800, 1490270400, 1490274000, 
    1490277600, 1490281200, 1490284800, 1490288400, 1490292000, 1490295600, 
    1490299200, 1490302800, 1490306400, 1490310000, 1490313600, 1490317200, 
    1490320800, 1490324400, 1490328000, 1490331600, 1490335200, 1490338800, 
    1490342400, 1490346000, 1490349600, 1490353200, 1490356800, 1490360400, 
    1490364000, 1490367600, 1490371200, 1490374800, 1490378400, 1490382000, 
    1490385600, 1490389200, 1490392800, 1490396400, 1490400000, 1490403600, 
    1490407200, 1490410800, 1490414400, 1490418000, 1490421600, 1490425200, 
    1490428800, 1490432400, 1490436000, 1490439600, 1490443200, 1490446800, 
    1490450400, 1490454000, 1490457600, 1490461200, 1490464800, 1490468400, 
    1490472000, 1490475600, 1490479200, 1490482800, 1490486400, 1490490000, 
    1490493600, 1490497200, 1490500800, 1490504400, 1490508000, 1490511600, 
    1490515200, 1490518800, 1490522400, 1490526000, 1490529600, 1490533200, 
    1490536800, 1490540400, 1490544000, 1490547600, 1490551200, 1490554800, 
    1490558400, 1490562000, 1490565600, 1490569200, 1490572800, 1490576400, 
    1490580000, 1490583600, 1490587200, 1490590800, 1490594400, 1490598000, 
    1490601600, 1490605200, 1490608800, 1490612400, 1490616000, 1490619600, 
    1490623200, 1490626800, 1490630400, 1490634000, 1490637600, 1490641200, 
    1490644800, 1490648400, 1490652000, 1490655600, 1490659200, 1490662800, 
    1490666400, 1490670000, 1490673600, 1490677200, 1490680800, 1490684400, 
    1490688000, 1490691600, 1490695200, 1490698800, 1490702400, 1490706000, 
    1490709600, 1490713200, 1490716800, 1490720400, 1490724000, 1490727600, 
    1490731200, 1490734800, 1490738400, 1490742000, 1490745600, 1490749200, 
    1490752800, 1490756400, 1490760000, 1490763600, 1490767200, 1490770800, 
    1490774400, 1490778000, 1490781600, 1490785200, 1490788800, 1490792400, 
    1490796000, 1490799600, 1490803200, 1490806800, 1490810400, 1490814000, 
    1490817600, 1490821200, 1490824800, 1490828400, 1490832000, 1490835600, 
    1490839200, 1490842800, 1490846400, 1490850000, 1490853600, 1490857200, 
    1490860800, 1490864400, 1490868000, 1490871600, 1490875200, 1490878800, 
    1490882400, 1490886000, 1490889600, 1490893200, 1490896800, 1490900400, 
    1490904000, 1490907600, 1490911200, 1490914800, 1490918400, 1490922000, 
    1490925600, 1490929200, 1490932800, 1490936400, 1490940000, 1490943600, 
    1490947200, 1490950800, 1490954400, 1490958000, 1490961600, 1490965200, 
    1490968800, 1490972400, 1490976000, 1490979600, 1490983200, 1490986800, 
    1490990400, 1490994000, 1490997600, 1491001200, 1491004800, 1491008400, 
    1491012000, 1491015600, 1491019200, 1491022800, 1491026400, 1491030000, 
    1491033600, 1491037200, 1491040800, 1491044400, 1491048000, 1491051600, 
    1491055200, 1491058800, 1491062400, 1491066000, 1491069600, 1491073200, 
    1491076800, 1491080400, 1491084000, 1491087600, 1491091200, 1491094800, 
    1491098400, 1491102000, 1491105600, 1491109200, 1491112800, 1491116400, 
    1491120000, 1491123600, 1491127200, 1491130800, 1491134400, 1491138000, 
    1491141600, 1491145200, 1491148800, 1491152400, 1491156000, 1491159600, 
    1491163200, 1491166800, 1491170400, 1491174000, 1491177600, 1491181200, 
    1491184800, 1491188400, 1491192000, 1491195600, 1491199200, 1491202800, 
    1491206400, 1491210000, 1491213600, 1491217200, 1491220800, 1491224400, 
    1491228000, 1491231600, 1491235200, 1491238800, 1491242400, 1491246000, 
    1491249600, 1491253200, 1491256800, 1491260400, 1491264000, 1491267600, 
    1491271200, 1491274800, 1491278400, 1491282000, 1491285600, 1491289200, 
    1491292800, 1491296400, 1491300000, 1491303600, 1491307200, 1491310800, 
    1491314400, 1491318000, 1491321600, 1491325200, 1491328800, 1491332400, 
    1491336000, 1491339600, 1491343200, 1491346800, 1491350400, 1491354000, 
    1491357600, 1491361200, 1491364800, 1491368400, 1491372000, 1491375600, 
    1491379200, 1491382800, 1491386400, 1491390000, 1491393600, 1491397200, 
    1491400800, 1491404400, 1491408000, 1491411600, 1491415200, 1491418800, 
    1491422400, 1491426000, 1491429600, 1491433200, 1491436800, 1491440400, 
    1491444000, 1491447600, 1491451200, 1491454800, 1491458400, 1491462000, 
    1491465600, 1491469200, 1491472800, 1491476400, 1491480000, 1491483600, 
    1491487200, 1491490800, 1491494400, 1491498000, 1491501600, 1491505200, 
    1491508800, 1491512400, 1491516000, 1491519600, 1491523200, 1491526800, 
    1491530400, 1491534000, 1491537600, 1491541200, 1491544800, 1491548400, 
    1491552000, 1491555600, 1491559200, 1491562800, 1491566400, 1491570000, 
    1491573600, 1491577200, 1491580800, 1491584400, 1491588000, 1491591600, 
    1491595200, 1491598800, 1491602400, 1491606000, 1491609600, 1491613200, 
    1491616800, 1491620400, 1491624000, 1491627600, 1491631200, 1491634800, 
    1491638400, 1491642000, 1491645600, 1491649200, 1491652800, 1491656400, 
    1491660000, 1491663600, 1491667200, 1491670800, 1491674400, 1491678000, 
    1491681600, 1491685200, 1491688800, 1491692400, 1491696000, 1491699600, 
    1491703200, 1491706800, 1491710400, 1491714000, 1491717600, 1491721200, 
    1491724800, 1491728400, 1491732000, 1491735600, 1491739200, 1491742800, 
    1491746400, 1491750000, 1491753600, 1491757200, 1491760800, 1491764400, 
    1491768000, 1491771600, 1491775200, 1491778800, 1491782400, 1491786000, 
    1491789600, 1491793200, 1491796800, 1491800400, 1491804000, 1491807600, 
    1491811200, 1491814800, 1491818400, 1491822000, 1491825600, 1491829200, 
    1491832800, 1491836400, 1491840000, 1491843600, 1491847200, 1491850800, 
    1491854400, 1491858000, 1491861600, 1491865200, 1491868800, 1491872400, 
    1491876000, 1491879600, 1491883200, 1491886800, 1491890400, 1491894000, 
    1491897600, 1491901200, 1491904800, 1491908400, 1491912000, 1491915600, 
    1491919200, 1491922800, 1491926400, 1491930000, 1491933600, 1491937200, 
    1491940800, 1491944400, 1491948000, 1491951600, 1491955200, 1491958800, 
    1491962400, 1491966000, 1491969600, 1491973200, 1491976800, 1491980400, 
    1491984000, 1491987600, 1491991200, 1491994800, 1491998400, 1492002000, 
    1492005600, 1492009200, 1492012800, 1492016400, 1492020000, 1492023600, 
    1492027200, 1492030800, 1492034400, 1492038000, 1492041600, 1492045200, 
    1492048800, 1492052400, 1492056000, 1492059600, 1492063200, 1492066800, 
    1492070400, 1492074000, 1492077600, 1492081200, 1492084800, 1492088400, 
    1492092000, 1492095600, 1492099200, 1492102800, 1492106400, 1492110000, 
    1492113600, 1492117200, 1492120800, 1492124400, 1492128000, 1492131600, 
    1492135200, 1492138800, 1492142400, 1492146000, 1492149600, 1492153200, 
    1492156800, 1492160400, 1492164000, 1492167600, 1492171200, 1492174800, 
    1492178400, 1492182000, 1492185600, 1492189200, 1492192800, 1492196400, 
    1492200000, 1492203600, 1492207200, 1492210800, 1492214400, 1492218000, 
    1492221600, 1492225200, 1492228800, 1492232400, 1492236000, 1492239600, 
    1492243200, 1492246800, 1492250400, 1492254000, 1492257600, 1492261200, 
    1492264800, 1492268400, 1492272000, 1492275600, 1492279200, 1492282800, 
    1492286400, 1492290000, 1492293600, 1492297200, 1492300800, 1492304400, 
    1492308000, 1492311600, 1492315200, 1492318800, 1492322400, 1492326000, 
    1492329600, 1492333200, 1492336800, 1492340400, 1492344000, 1492347600, 
    1492351200, 1492354800, 1492358400, 1492362000, 1492365600, 1492369200, 
    1492372800, 1492376400, 1492380000, 1492383600, 1492387200, 1492390800, 
    1492394400, 1492398000, 1492401600, 1492405200, 1492408800, 1492412400, 
    1492416000, 1492419600, 1492423200, 1492426800, 1492430400, 1492434000, 
    1492437600, 1492441200, 1492444800, 1492448400, 1492452000, 1492455600, 
    1492459200, 1492462800, 1492466400, 1492470000, 1492473600, 1492477200, 
    1492480800, 1492484400, 1492488000, 1492491600, 1492495200, 1492498800, 
    1492502400, 1492506000, 1492509600, 1492513200, 1492516800, 1492520400, 
    1492524000, 1492527600, 1492531200, 1492534800, 1492538400, 1492542000, 
    1492545600, 1492549200, 1492552800, 1492556400, 1492560000, 1492563600, 
    1492567200, 1492570800, 1492574400, 1492578000, 1492581600, 1492585200, 
    1492588800, 1492592400, 1492596000, 1492599600, 1492603200, 1492606800, 
    1492610400, 1492614000, 1492617600, 1492621200, 1492624800, 1492628400, 
    1492632000, 1492635600, 1492639200, 1492642800, 1492646400, 1492650000, 
    1492653600, 1492657200, 1492660800, 1492664400, 1492668000, 1492671600, 
    1492675200, 1492678800, 1492682400, 1492686000, 1492689600, 1492693200, 
    1492696800, 1492700400, 1492704000, 1492707600, 1492711200, 1492714800, 
    1492718400, 1492722000, 1492725600, 1492729200, 1492732800, 1492736400, 
    1492740000, 1492743600, 1492747200, 1492750800, 1492754400, 1492758000, 
    1492761600, 1492765200, 1492768800, 1492772400, 1492776000, 1492779600, 
    1492783200, 1492786800, 1492790400, 1492794000, 1492797600, 1492801200, 
    1492804800, 1492808400, 1492812000, 1492815600, 1492819200, 1492822800, 
    1492826400, 1492830000, 1492833600, 1492837200, 1492840800, 1492844400, 
    1492848000, 1492851600, 1492855200, 1492858800, 1492862400, 1492866000, 
    1492869600, 1492873200, 1492876800, 1492880400, 1492884000, 1492887600, 
    1492891200, 1492894800, 1492898400, 1492902000, 1492905600, 1492909200, 
    1492912800, 1492916400, 1492920000, 1492923600, 1492927200, 1492930800, 
    1492934400, 1492938000, 1492941600, 1492945200, 1492948800, 1492952400, 
    1492956000, 1492959600, 1492963200, 1492966800, 1492970400, 1492974000, 
    1492977600, 1492981200, 1492984800, 1492988400, 1492992000, 1492995600, 
    1492999200, 1493002800, 1493006400, 1493010000, 1493013600, 1493017200, 
    1493020800, 1493024400, 1493028000, 1493031600, 1493035200, 1493038800, 
    1493042400, 1493046000, 1493049600, 1493053200, 1493056800, 1493060400, 
    1493064000, 1493067600, 1493071200, 1493074800, 1493078400, 1493082000, 
    1493085600, 1493089200, 1493092800, 1493096400, 1493100000, 1493103600, 
    1493107200, 1493110800, 1493114400, 1493118000, 1493121600, 1493125200, 
    1493128800, 1493132400, 1493136000, 1493139600, 1493143200, 1493146800, 
    1493150400, 1493154000, 1493157600, 1493161200, 1493164800, 1493168400, 
    1493172000, 1493175600, 1493179200, 1493182800, 1493186400, 1493190000, 
    1493193600, 1493197200, 1493200800, 1493204400, 1493208000, 1493211600, 
    1493215200, 1493218800, 1493222400, 1493226000, 1493229600, 1493233200, 
    1493236800, 1493240400, 1493244000, 1493247600, 1493251200, 1493254800, 
    1493258400, 1493262000, 1493265600, 1493269200, 1493272800, 1493276400, 
    1493280000, 1493283600, 1493287200, 1493290800, 1493294400, 1493298000, 
    1493301600, 1493305200, 1493308800, 1493312400, 1493316000, 1493319600, 
    1493323200, 1493326800, 1493330400, 1493334000, 1493337600, 1493341200, 
    1493344800, 1493348400, 1493352000, 1493355600, 1493359200, 1493362800, 
    1493366400, 1493370000, 1493373600, 1493377200, 1493380800, 1493384400, 
    1493388000, 1493391600, 1493395200, 1493398800, 1493402400, 1493406000, 
    1493409600, 1493413200, 1493416800, 1493420400, 1493424000, 1493427600, 
    1493431200, 1493434800, 1493438400, 1493442000, 1493445600, 1493449200, 
    1493452800, 1493456400, 1493460000, 1493463600, 1493467200, 1493470800, 
    1493474400, 1493478000, 1493481600, 1493485200, 1493488800, 1493492400, 
    1493496000, 1493499600, 1493503200, 1493506800, 1493510400, 1493514000, 
    1493517600, 1493521200, 1493524800, 1493528400, 1493532000, 1493535600, 
    1493539200, 1493542800, 1493546400, 1493550000, 1493553600, 1493557200, 
    1493560800, 1493564400, 1493568000, 1493571600, 1493575200, 1493578800, 
    1493582400, 1493586000, 1493589600, 1493593200, 1493596800, 1493600400, 
    1493604000, 1493607600, 1493611200, 1493614800, 1493618400, 1493622000, 
    1493625600, 1493629200, 1493632800, 1493636400, 1493640000, 1493643600, 
    1493647200, 1493650800, 1493654400, 1493658000, 1493661600, 1493665200, 
    1493668800, 1493672400, 1493676000, 1493679600, 1493683200, 1493686800, 
    1493690400, 1493694000, 1493697600, 1493701200, 1493704800, 1493708400, 
    1493712000, 1493715600, 1493719200, 1493722800, 1493726400, 1493730000, 
    1493733600, 1493737200, 1493740800, 1493744400, 1493748000, 1493751600, 
    1493755200, 1493758800, 1493762400, 1493766000, 1493769600, 1493773200, 
    1493776800, 1493780400, 1493784000, 1493787600, 1493791200, 1493794800, 
    1493798400, 1493802000, 1493805600, 1493809200, 1493812800, 1493816400, 
    1493820000, 1493823600, 1493827200, 1493830800, 1493834400, 1493838000, 
    1493841600, 1493845200, 1493848800, 1493852400, 1493856000, 1493859600, 
    1493863200, 1493866800, 1493870400, 1493874000, 1493877600, 1493881200, 
    1493884800, 1493888400, 1493892000, 1493895600, 1493899200, 1493902800, 
    1493906400, 1493910000, 1493913600, 1493917200, 1493920800, 1493924400, 
    1493928000, 1493931600, 1493935200, 1493938800, 1493942400, 1493946000, 
    1493949600, 1493953200, 1493956800, 1493960400, 1493964000, 1493967600, 
    1493971200, 1493974800, 1493978400, 1493982000, 1493985600, 1493989200, 
    1493992800, 1493996400, 1494000000, 1494003600, 1494007200, 1494010800, 
    1494014400, 1494018000, 1494021600, 1494025200, 1494028800, 1494032400, 
    1494036000, 1494039600, 1494043200, 1494046800, 1494050400, 1494054000, 
    1494057600, 1494061200, 1494064800, 1494068400, 1494072000, 1494075600, 
    1494079200, 1494082800, 1494086400, 1494090000, 1494093600, 1494097200, 
    1494100800, 1494104400, 1494108000, 1494111600, 1494115200, 1494118800, 
    1494122400, 1494126000, 1494129600, 1494133200, 1494136800, 1494140400, 
    1494144000, 1494147600, 1494151200, 1494154800, 1494158400, 1494162000, 
    1494165600, 1494169200, 1494172800, 1494176400, 1494180000, 1494183600, 
    1494187200, 1494190800, 1494194400, 1494198000, 1494201600, 1494205200, 
    1494208800, 1494212400, 1494216000, 1494219600, 1494223200, 1494226800, 
    1494230400, 1494234000, 1494237600, 1494241200, 1494244800, 1494248400, 
    1494252000, 1494255600, 1494259200, 1494262800, 1494266400, 1494270000, 
    1494273600, 1494277200, 1494280800, 1494284400, 1494288000, 1494291600, 
    1494295200, 1494298800, 1494302400, 1494306000, 1494309600, 1494313200, 
    1494316800, 1494320400, 1494324000, 1494327600, 1494331200, 1494334800, 
    1494338400, 1494342000, 1494345600, 1494349200, 1494352800, 1494356400, 
    1494360000, 1494363600, 1494367200, 1494370800, 1494374400, 1494378000, 
    1494381600, 1494385200, 1494388800, 1494392400, 1494396000, 1494399600, 
    1494403200, 1494406800, 1494410400, 1494414000, 1494417600, 1494421200, 
    1494424800, 1494428400, 1494432000, 1494435600, 1494439200, 1494442800, 
    1494446400, 1494450000, 1494453600, 1494457200, 1494460800, 1494464400, 
    1494468000, 1494471600, 1494475200, 1494478800, 1494482400, 1494486000, 
    1494489600, 1494493200, 1494496800, 1494500400, 1494504000, 1494507600, 
    1494511200, 1494514800, 1494518400, 1494522000, 1494525600, 1494529200, 
    1494532800, 1494536400, 1494540000, 1494543600, 1494547200, 1494550800, 
    1494554400, 1494558000, 1494561600, 1494565200, 1494568800, 1494572400, 
    1494576000, 1494579600, 1494583200, 1494586800, 1494590400, 1494594000, 
    1494597600, 1494601200, 1494604800, 1494608400, 1494612000, 1494615600, 
    1494619200, 1494622800, 1494626400, 1494630000, 1494633600, 1494637200, 
    1494640800, 1494644400, 1494648000, 1494651600, 1494655200, 1494658800, 
    1494662400, 1494666000, 1494669600, 1494673200, 1494676800, 1494680400, 
    1494684000, 1494687600, 1494691200, 1494694800, 1494698400, 1494702000, 
    1494705600, 1494709200, 1494712800, 1494716400, 1494720000, 1494723600, 
    1494727200, 1494730800, 1494734400, 1494738000, 1494741600, 1494745200, 
    1494748800, 1494752400, 1494756000, 1494759600, 1494763200, 1494766800, 
    1494770400, 1494774000, 1494777600, 1494781200, 1494784800, 1494788400, 
    1494792000, 1494795600, 1494799200, 1494802800, 1494806400, 1494810000, 
    1494813600, 1494817200, 1494820800, 1494824400, 1494828000, 1494831600, 
    1494835200, 1494838800, 1494842400, 1494846000, 1494849600, 1494853200, 
    1494856800, 1494860400, 1494864000, 1494867600, 1494871200, 1494874800, 
    1494878400, 1494882000, 1494885600, 1494889200, 1494892800, 1494896400, 
    1494900000, 1494903600, 1494907200, 1494910800, 1494914400, 1494918000, 
    1494921600, 1494925200, 1494928800, 1494932400, 1494936000, 1494939600, 
    1494943200, 1494946800, 1494950400, 1494954000, 1494957600, 1494961200, 
    1494964800, 1494968400, 1494972000, 1494975600, 1494979200, 1494982800, 
    1494986400, 1494990000, 1494993600, 1494997200, 1495000800, 1495004400, 
    1495008000, 1495011600, 1495015200, 1495018800, 1495022400, 1495026000, 
    1495029600, 1495033200, 1495036800, 1495040400, 1495044000, 1495047600, 
    1495051200, 1495054800, 1495058400, 1495062000, 1495065600, 1495069200, 
    1495072800, 1495076400, 1495080000, 1495083600, 1495087200, 1495090800, 
    1495094400, 1495098000, 1495101600, 1495105200, 1495108800, 1495112400, 
    1495116000, 1495119600, 1495123200, 1495126800, 1495130400, 1495134000, 
    1495137600, 1495141200, 1495144800, 1495148400, 1495152000, 1495155600, 
    1495159200, 1495162800, 1495166400, 1495170000, 1495173600, 1495177200, 
    1495180800, 1495184400, 1495188000, 1495191600, 1495195200, 1495198800, 
    1495202400, 1495206000, 1495209600, 1495213200, 1495216800, 1495220400, 
    1495224000, 1495227600, 1495231200, 1495234800, 1495238400, 1495242000, 
    1495245600, 1495249200, 1495252800, 1495256400, 1495260000, 1495263600, 
    1495267200, 1495270800, 1495274400, 1495278000, 1495281600, 1495285200, 
    1495288800, 1495292400, 1495296000, 1495299600, 1495303200, 1495306800, 
    1495310400, 1495314000, 1495317600, 1495321200, 1495324800, 1495328400, 
    1495332000, 1495335600, 1495339200, 1495342800, 1495346400, 1495350000, 
    1495353600, 1495357200, 1495360800, 1495364400, 1495368000, 1495371600, 
    1495375200, 1495378800, 1495382400, 1495386000, 1495389600, 1495393200, 
    1495396800, 1495400400, 1495404000, 1495407600, 1495411200, 1495414800, 
    1495418400, 1495422000, 1495425600, 1495429200, 1495432800, 1495436400, 
    1495440000, 1495443600, 1495447200, 1495450800, 1495454400, 1495458000, 
    1495461600, 1495465200, 1495468800, 1495472400, 1495476000, 1495479600, 
    1495483200, 1495486800, 1495490400, 1495494000, 1495497600, 1495501200, 
    1495504800, 1495508400, 1495512000, 1495515600, 1495519200, 1495522800, 
    1495526400, 1495530000, 1495533600, 1495537200, 1495540800, 1495544400, 
    1495548000, 1495551600, 1495555200, 1495558800, 1495562400, 1495566000, 
    1495569600, 1495573200, 1495576800, 1495580400, 1495584000, 1495587600, 
    1495591200, 1495594800, 1495598400, 1495602000, 1495605600, 1495609200, 
    1495612800, 1495616400, 1495620000, 1495623600, 1495627200, 1495630800, 
    1495634400, 1495638000, 1495641600, 1495645200, 1495648800, 1495652400, 
    1495656000, 1495659600, 1495663200, 1495666800, 1495670400, 1495674000, 
    1495677600, 1495681200, 1495684800, 1495688400, 1495692000, 1495695600, 
    1495699200, 1495702800, 1495706400, 1495710000, 1495713600, 1495717200, 
    1495720800, 1495724400, 1495728000, 1495731600, 1495735200, 1495738800, 
    1495742400, 1495746000, 1495749600, 1495753200, 1495756800, 1495760400, 
    1495764000, 1495767600, 1495771200, 1495774800, 1495778400, 1495782000, 
    1495785600, 1495789200, 1495792800, 1495796400, 1495800000, 1495803600, 
    1495807200, 1495810800, 1495814400, 1495818000, 1495821600, 1495825200, 
    1495828800, 1495832400, 1495836000, 1495839600, 1495843200, 1495846800, 
    1495850400, 1495854000, 1495857600, 1495861200, 1495864800, 1495868400, 
    1495872000, 1495875600, 1495879200, 1495882800, 1495886400, 1495890000, 
    1495893600, 1495897200, 1495900800, 1495904400, 1495908000, 1495911600, 
    1495915200, 1495918800, 1495922400, 1495926000, 1495929600, 1495933200, 
    1495936800, 1495940400, 1495944000, 1495947600, 1495951200, 1495954800, 
    1495958400, 1495962000, 1495965600, 1495969200, 1495972800, 1495976400, 
    1495980000, 1495983600, 1495987200, 1495990800, 1495994400, 1495998000, 
    1496001600, 1496005200, 1496008800, 1496012400, 1496016000, 1496019600, 
    1496023200, 1496026800, 1496030400, 1496034000, 1496037600, 1496041200, 
    1496044800, 1496048400, 1496052000, 1496055600, 1496059200, 1496062800, 
    1496066400, 1496070000, 1496073600, 1496077200, 1496080800, 1496084400, 
    1496088000, 1496091600, 1496095200, 1496098800, 1496102400, 1496106000, 
    1496109600, 1496113200, 1496116800, 1496120400, 1496124000, 1496127600, 
    1496131200, 1496134800, 1496138400, 1496142000, 1496145600, 1496149200, 
    1496152800, 1496156400, 1496160000, 1496163600, 1496167200, 1496170800, 
    1496174400, 1496178000, 1496181600, 1496185200, 1496188800, 1496192400, 
    1496196000, 1496199600, 1496203200, 1496206800, 1496210400, 1496214000, 
    1496217600, 1496221200, 1496224800, 1496228400, 1496232000, 1496235600, 
    1496239200, 1496242800, 1496246400, 1496250000, 1496253600, 1496257200, 
    1496260800, 1496264400, 1496268000, 1496271600, 1496275200, 1496278800, 
    1496282400, 1496286000, 1496289600, 1496293200, 1496296800, 1496300400, 
    1496304000, 1496307600, 1496311200, 1496314800, 1496318400, 1496322000, 
    1496325600, 1496329200, 1496332800, 1496336400, 1496340000, 1496343600, 
    1496347200, 1496350800, 1496354400, 1496358000, 1496361600, 1496365200, 
    1496368800, 1496372400, 1496376000, 1496379600, 1496383200, 1496386800, 
    1496390400, 1496394000, 1496397600, 1496401200, 1496404800, 1496408400, 
    1496412000, 1496415600, 1496419200, 1496422800, 1496426400, 1496430000, 
    1496433600, 1496437200, 1496440800, 1496444400, 1496448000, 1496451600, 
    1496455200, 1496458800, 1496462400, 1496466000, 1496469600, 1496473200, 
    1496476800, 1496480400, 1496484000, 1496487600, 1496491200, 1496494800, 
    1496498400, 1496502000, 1496505600, 1496509200, 1496512800, 1496516400, 
    1496520000, 1496523600, 1496527200, 1496530800, 1496534400, 1496538000, 
    1496541600, 1496545200, 1496548800, 1496552400, 1496556000, 1496559600, 
    1496563200, 1496566800, 1496570400, 1496574000, 1496577600, 1496581200, 
    1496584800, 1496588400, 1496592000, 1496595600, 1496599200, 1496602800, 
    1496606400, 1496610000, 1496613600, 1496617200, 1496620800, 1496624400, 
    1496628000, 1496631600, 1496635200, 1496638800, 1496642400, 1496646000, 
    1496649600, 1496653200, 1496656800, 1496660400, 1496664000, 1496667600, 
    1496671200, 1496674800, 1496678400, 1496682000, 1496685600, 1496689200, 
    1496692800, 1496696400, 1496700000, 1496703600, 1496707200, 1496710800, 
    1496714400, 1496718000, 1496721600, 1496725200, 1496728800, 1496732400, 
    1496736000, 1496739600, 1496743200, 1496746800, 1496750400, 1496754000, 
    1496757600, 1496761200, 1496764800, 1496768400, 1496772000, 1496775600, 
    1496779200, 1496782800, 1496786400, 1496790000, 1496793600, 1496797200, 
    1496800800, 1496804400, 1496808000, 1496811600, 1496815200, 1496818800, 
    1496822400, 1496826000, 1496829600, 1496833200, 1496836800, 1496840400, 
    1496844000, 1496847600, 1496851200, 1496854800, 1496858400, 1496862000, 
    1496865600, 1496869200, 1496872800, 1496876400, 1496880000, 1496883600, 
    1496887200, 1496890800, 1496894400, 1496898000, 1496901600, 1496905200, 
    1496908800, 1496912400, 1496916000, 1496919600, 1496923200, 1496926800, 
    1496930400, 1496934000, 1496937600, 1496941200, 1496944800, 1496948400, 
    1496952000, 1496955600, 1496959200, 1496962800, 1496966400, 1496970000, 
    1496973600, 1496977200, 1496980800, 1496984400, 1496988000, 1496991600, 
    1496995200, 1496998800, 1497002400, 1497006000, 1497009600, 1497013200, 
    1497016800, 1497020400, 1497024000, 1497027600, 1497031200, 1497034800, 
    1497038400, 1497042000, 1497045600, 1497049200, 1497052800, 1497056400, 
    1497060000, 1497063600, 1497067200, 1497070800, 1497074400, 1497078000, 
    1497081600, 1497085200, 1497088800, 1497092400, 1497096000, 1497099600, 
    1497103200, 1497106800, 1497110400, 1497114000, 1497117600, 1497121200, 
    1497124800, 1497128400, 1497132000, 1497135600, 1497139200, 1497142800, 
    1497146400, 1497150000, 1497153600, 1497157200, 1497160800, 1497164400, 
    1497168000, 1497171600, 1497175200, 1497178800, 1497182400, 1497186000, 
    1497189600, 1497193200, 1497196800, 1497200400, 1497204000, 1497207600, 
    1497211200, 1497214800, 1497218400, 1497222000, 1497225600, 1497229200, 
    1497232800, 1497236400, 1497240000, 1497243600, 1497247200, 1497250800, 
    1497254400, 1497258000, 1497261600, 1497265200, 1497268800, 1497272400, 
    1497276000, 1497279600, 1497283200, 1497286800, 1497290400, 1497294000, 
    1497297600, 1497301200, 1497304800, 1497308400, 1497312000, 1497315600, 
    1497319200, 1497322800, 1497326400, 1497330000, 1497333600, 1497337200, 
    1497340800, 1497344400, 1497348000, 1497351600, 1497355200, 1497358800, 
    1497362400, 1497366000, 1497369600, 1497373200, 1497376800, 1497380400, 
    1497384000, 1497387600, 1497391200, 1497394800, 1497398400, 1497402000, 
    1497405600, 1497409200, 1497412800, 1497416400, 1497420000, 1497423600, 
    1497427200, 1497430800, 1497434400, 1497438000, 1497441600, 1497445200, 
    1497448800, 1497452400, 1497456000, 1497459600, 1497463200, 1497466800, 
    1497470400, 1497474000, 1497477600, 1497481200, 1497484800, 1497488400, 
    1497492000, 1497495600, 1497499200, 1497502800, 1497506400, 1497510000, 
    1497513600, 1497517200, 1497520800, 1497524400, 1497528000, 1497531600, 
    1497535200, 1497538800, 1497542400, 1497546000, 1497549600, 1497553200, 
    1497556800, 1497560400, 1497564000, 1497567600, 1497571200, 1497574800, 
    1497578400, 1497582000, 1497585600, 1497589200, 1497592800, 1497596400, 
    1497600000, 1497603600, 1497607200, 1497610800, 1497614400, 1497618000, 
    1497621600, 1497625200, 1497628800, 1497632400, 1497636000, 1497639600, 
    1497643200, 1497646800, 1497650400, 1497654000, 1497657600, 1497661200, 
    1497664800, 1497668400, 1497672000, 1497675600, 1497679200, 1497682800, 
    1497686400, 1497690000, 1497693600, 1497697200, 1497700800, 1497704400, 
    1497708000, 1497711600, 1497715200, 1497718800, 1497722400, 1497726000, 
    1497729600, 1497733200, 1497736800, 1497740400, 1497744000, 1497747600, 
    1497751200, 1497754800, 1497758400, 1497762000, 1497765600, 1497769200, 
    1497772800, 1497776400, 1497780000, 1497783600, 1497787200, 1497790800, 
    1497794400, 1497798000, 1497801600, 1497805200, 1497808800, 1497812400, 
    1497816000, 1497819600, 1497823200, 1497826800, 1497830400, 1497834000, 
    1497837600, 1497841200, 1497844800, 1497848400, 1497852000, 1497855600, 
    1497859200, 1497862800, 1497866400, 1497870000, 1497873600, 1497877200, 
    1497880800, 1497884400, 1497888000, 1497891600, 1497895200, 1497898800, 
    1497902400, 1497906000, 1497909600, 1497913200, 1497916800, 1497920400, 
    1497924000, 1497927600, 1497931200, 1497934800, 1497938400, 1497942000, 
    1497945600, 1497949200, 1497952800, 1497956400, 1497960000, 1497963600, 
    1497967200, 1497970800, 1497974400, 1497978000, 1497981600, 1497985200, 
    1497988800, 1497992400, 1497996000, 1497999600, 1498003200, 1498006800, 
    1498010400, 1498014000, 1498017600, 1498021200, 1498024800, 1498028400, 
    1498032000, 1498035600, 1498039200, 1498042800, 1498046400, 1498050000, 
    1498053600, 1498057200, 1498060800, 1498064400, 1498068000, 1498071600, 
    1498075200, 1498078800, 1498082400, 1498086000, 1498089600, 1498093200, 
    1498096800, 1498100400, 1498104000, 1498107600, 1498111200, 1498114800, 
    1498118400, 1498122000, 1498125600, 1498129200, 1498132800, 1498136400, 
    1498140000, 1498143600, 1498147200, 1498150800, 1498154400, 1498158000, 
    1498161600, 1498165200, 1498168800, 1498172400, 1498176000, 1498179600, 
    1498183200, 1498186800, 1498190400, 1498194000, 1498197600, 1498201200, 
    1498204800, 1498208400, 1498212000, 1498215600, 1498219200, 1498222800, 
    1498226400, 1498230000, 1498233600, 1498237200, 1498240800, 1498244400, 
    1498248000, 1498251600, 1498255200, 1498258800, 1498262400, 1498266000, 
    1498269600, 1498273200, 1498276800, 1498280400, 1498284000, 1498287600, 
    1498291200, 1498294800, 1498298400, 1498302000, 1498305600, 1498309200, 
    1498312800, 1498316400, 1498320000, 1498323600, 1498327200, 1498330800, 
    1498334400, 1498338000, 1498341600, 1498345200, 1498348800, 1498352400, 
    1498356000, 1498359600, 1498363200, 1498366800, 1498370400, 1498374000, 
    1498377600, 1498381200, 1498384800, 1498388400, 1498392000, 1498395600, 
    1498399200, 1498402800, 1498406400, 1498410000, 1498413600, 1498417200, 
    1498420800, 1498424400, 1498428000, 1498431600, 1498435200, 1498438800, 
    1498442400, 1498446000, 1498449600, 1498453200, 1498456800, 1498460400, 
    1498464000, 1498467600, 1498471200, 1498474800, 1498478400, 1498482000, 
    1498485600, 1498489200, 1498492800, 1498496400, 1498500000, 1498503600, 
    1498507200, 1498510800, 1498514400, 1498518000, 1498521600, 1498525200, 
    1498528800, 1498532400, 1498536000, 1498539600, 1498543200, 1498546800, 
    1498550400, 1498554000, 1498557600, 1498561200, 1498564800, 1498568400, 
    1498572000, 1498575600, 1498579200, 1498582800, 1498586400, 1498590000, 
    1498593600, 1498597200, 1498600800, 1498604400, 1498608000, 1498611600, 
    1498615200, 1498618800, 1498622400, 1498626000, 1498629600, 1498633200, 
    1498636800, 1498640400, 1498644000, 1498647600, 1498651200, 1498654800, 
    1498658400, 1498662000, 1498665600, 1498669200, 1498672800, 1498676400, 
    1498680000, 1498683600, 1498687200, 1498690800, 1498694400, 1498698000, 
    1498701600, 1498705200, 1498708800, 1498712400, 1498716000, 1498719600, 
    1498723200, 1498726800, 1498730400, 1498734000, 1498737600, 1498741200, 
    1498744800, 1498748400, 1498752000, 1498755600, 1498759200, 1498762800, 
    1498766400, 1498770000, 1498773600, 1498777200, 1498780800, 1498784400, 
    1498788000, 1498791600, 1498795200, 1498798800, 1498802400, 1498806000, 
    1498809600, 1498813200, 1498816800, 1498820400, 1498824000, 1498827600, 
    1498831200, 1498834800, 1498838400, 1498842000, 1498845600, 1498849200, 
    1498852800, 1498856400, 1498860000, 1498863600, 1498867200, 1498870800, 
    1498874400, 1498878000, 1498881600, 1498885200, 1498888800, 1498892400, 
    1498896000, 1498899600, 1498903200, 1498906800, 1498910400, 1498914000, 
    1498917600, 1498921200, 1498924800, 1498928400, 1498932000, 1498935600, 
    1498939200, 1498942800, 1498946400, 1498950000, 1498953600, 1498957200, 
    1498960800, 1498964400, 1498968000, 1498971600, 1498975200, 1498978800, 
    1498982400, 1498986000, 1498989600, 1498993200, 1498996800, 1499000400, 
    1499004000, 1499007600, 1499011200, 1499014800, 1499018400, 1499022000, 
    1499025600, 1499029200, 1499032800, 1499036400, 1499040000, 1499043600, 
    1499047200, 1499050800, 1499054400, 1499058000, 1499061600, 1499065200, 
    1499068800, 1499072400, 1499076000, 1499079600, 1499083200, 1499086800, 
    1499090400, 1499094000, 1499097600, 1499101200, 1499104800, 1499108400, 
    1499112000, 1499115600, 1499119200, 1499122800, 1499126400, 1499130000, 
    1499133600, 1499137200, 1499140800, 1499144400, 1499148000, 1499151600, 
    1499155200, 1499158800, 1499162400, 1499166000, 1499169600, 1499173200, 
    1499176800, 1499180400, 1499184000, 1499187600, 1499191200, 1499194800, 
    1499198400, 1499202000, 1499205600, 1499209200, 1499212800, 1499216400, 
    1499220000, 1499223600, 1499227200, 1499230800, 1499234400, 1499238000, 
    1499241600, 1499245200, 1499248800, 1499252400, 1499256000, 1499259600, 
    1499263200, 1499266800, 1499270400, 1499274000, 1499277600, 1499281200, 
    1499284800, 1499288400, 1499292000, 1499295600, 1499299200, 1499302800, 
    1499306400, 1499310000, 1499313600, 1499317200, 1499320800, 1499324400, 
    1499328000, 1499331600, 1499335200, 1499338800, 1499342400, 1499346000, 
    1499349600, 1499353200, 1499356800, 1499360400, 1499364000, 1499367600, 
    1499371200, 1499374800, 1499378400, 1499382000, 1499385600, 1499389200, 
    1499392800, 1499396400, 1499400000, 1499403600, 1499407200, 1499410800, 
    1499414400, 1499418000, 1499421600, 1499425200, 1499428800, 1499432400, 
    1499436000, 1499439600, 1499443200, 1499446800, 1499450400, 1499454000, 
    1499457600, 1499461200, 1499464800, 1499468400, 1499472000, 1499475600, 
    1499479200, 1499482800, 1499486400, 1499490000, 1499493600, 1499497200, 
    1499500800, 1499504400, 1499508000, 1499511600, 1499515200, 1499518800, 
    1499522400, 1499526000, 1499529600, 1499533200, 1499536800, 1499540400, 
    1499544000, 1499547600, 1499551200, 1499554800, 1499558400, 1499562000, 
    1499565600, 1499569200, 1499572800, 1499576400, 1499580000, 1499583600, 
    1499587200, 1499590800, 1499594400, 1499598000, 1499601600, 1499605200, 
    1499608800, 1499612400, 1499616000, 1499619600, 1499623200, 1499626800, 
    1499630400, 1499634000, 1499637600, 1499641200, 1499644800, 1499648400, 
    1499652000, 1499655600, 1499659200, 1499662800, 1499666400, 1499670000, 
    1499673600, 1499677200, 1499680800, 1499684400, 1499688000, 1499691600, 
    1499695200, 1499698800, 1499702400, 1499706000, 1499709600, 1499713200, 
    1499716800, 1499720400, 1499724000, 1499727600, 1499731200, 1499734800, 
    1499738400, 1499742000, 1499745600, 1499749200, 1499752800, 1499756400, 
    1499760000, 1499763600, 1499767200, 1499770800, 1499774400, 1499778000, 
    1499781600, 1499785200, 1499788800, 1499792400, 1499796000, 1499799600, 
    1499803200, 1499806800, 1499810400, 1499814000, 1499817600, 1499821200, 
    1499824800, 1499828400, 1499832000, 1499835600, 1499839200, 1499842800, 
    1499846400, 1499850000, 1499853600, 1499857200, 1499860800, 1499864400, 
    1499868000, 1499871600, 1499875200, 1499878800, 1499882400, 1499886000, 
    1499889600, 1499893200, 1499896800, 1499900400, 1499904000, 1499907600, 
    1499911200, 1499914800, 1499918400, 1499922000, 1499925600, 1499929200, 
    1499932800, 1499936400, 1499940000, 1499943600, 1499947200, 1499950800, 
    1499954400, 1499958000, 1499961600, 1499965200, 1499968800, 1499972400, 
    1499976000, 1499979600, 1499983200, 1499986800, 1499990400, 1499994000, 
    1499997600, 1500001200, 1500004800, 1500008400, 1500012000, 1500015600, 
    1500019200, 1500022800, 1500026400, 1500030000, 1500033600, 1500037200, 
    1500040800, 1500044400, 1500048000, 1500051600, 1500055200, 1500058800, 
    1500062400, 1500066000, 1500069600, 1500073200, 1500076800, 1500080400, 
    1500084000, 1500087600, 1500091200, 1500094800, 1500098400, 1500102000, 
    1500105600, 1500109200, 1500112800, 1500116400, 1500120000, 1500123600, 
    1500127200, 1500130800, 1500134400, 1500138000, 1500141600, 1500145200, 
    1500148800, 1500152400, 1500156000, 1500159600, 1500163200, 1500166800, 
    1500170400, 1500174000, 1500177600, 1500181200, 1500184800, 1500188400, 
    1500192000, 1500195600, 1500199200, 1500202800, 1500206400, 1500210000, 
    1500213600, 1500217200, 1500220800, 1500224400, 1500228000, 1500231600, 
    1500235200, 1500238800, 1500242400, 1500246000, 1500249600, 1500253200, 
    1500256800, 1500260400, 1500264000, 1500267600, 1500271200, 1500274800, 
    1500278400, 1500282000, 1500285600, 1500289200, 1500292800, 1500296400, 
    1500300000, 1500303600, 1500307200, 1500310800, 1500314400, 1500318000, 
    1500321600, 1500325200, 1500328800, 1500332400, 1500336000, 1500339600, 
    1500343200, 1500346800, 1500350400, 1500354000, 1500357600, 1500361200, 
    1500364800, 1500368400, 1500372000, 1500375600, 1500379200, 1500382800, 
    1500386400, 1500390000, 1500393600, 1500397200, 1500400800, 1500404400, 
    1500408000, 1500411600, 1500415200, 1500418800, 1500422400, 1500426000, 
    1500429600, 1500433200, 1500436800, 1500440400, 1500444000, 1500447600, 
    1500451200, 1500454800, 1500458400, 1500462000, 1500465600, 1500469200, 
    1500472800, 1500476400, 1500480000, 1500483600, 1500487200, 1500490800, 
    1500494400, 1500498000, 1500501600, 1500505200, 1500508800, 1500512400, 
    1500516000, 1500519600, 1500523200, 1500526800, 1500530400, 1500534000, 
    1500537600, 1500541200, 1500544800, 1500548400, 1500552000, 1500555600, 
    1500559200, 1500562800, 1500566400, 1500570000, 1500573600, 1500577200, 
    1500580800, 1500584400, 1500588000, 1500591600, 1500595200, 1500598800, 
    1500602400, 1500606000, 1500609600, 1500613200, 1500616800, 1500620400, 
    1500624000, 1500627600, 1500631200, 1500634800, 1500638400, 1500642000, 
    1500645600, 1500649200, 1500652800, 1500656400, 1500660000, 1500663600, 
    1500667200, 1500670800, 1500674400, 1500678000, 1500681600, 1500685200, 
    1500688800, 1500692400, 1500696000, 1500699600, 1500703200, 1500706800, 
    1500710400, 1500714000, 1500717600, 1500721200, 1500724800, 1500728400, 
    1500732000, 1500735600, 1500739200, 1500742800, 1500746400, 1500750000, 
    1500753600, 1500757200, 1500760800, 1500764400, 1500768000, 1500771600, 
    1500775200, 1500778800, 1500782400, 1500786000, 1500789600, 1500793200, 
    1500796800, 1500800400, 1500804000, 1500807600, 1500811200, 1500814800, 
    1500818400, 1500822000, 1500825600, 1500829200, 1500832800, 1500836400, 
    1500840000, 1500843600, 1500847200, 1500850800, 1500854400, 1500858000, 
    1500861600, 1500865200, 1500868800, 1500872400, 1500876000, 1500879600, 
    1500883200, 1500886800, 1500890400, 1500894000, 1500897600, 1500901200, 
    1500904800, 1500908400, 1500912000, 1500915600, 1500919200, 1500922800, 
    1500926400, 1500930000, 1500933600, 1500937200, 1500940800, 1500944400, 
    1500948000, 1500951600, 1500955200, 1500958800, 1500962400, 1500966000, 
    1500969600, 1500973200, 1500976800, 1500980400, 1500984000, 1500987600, 
    1500991200, 1500994800, 1500998400, 1501002000, 1501005600, 1501009200, 
    1501012800, 1501016400, 1501020000, 1501023600, 1501027200, 1501030800, 
    1501034400, 1501038000, 1501041600, 1501045200, 1501048800, 1501052400, 
    1501056000, 1501059600, 1501063200, 1501066800, 1501070400, 1501074000, 
    1501077600, 1501081200, 1501084800, 1501088400, 1501092000, 1501095600, 
    1501099200, 1501102800, 1501106400, 1501110000, 1501113600, 1501117200, 
    1501120800, 1501124400, 1501128000, 1501131600, 1501135200, 1501138800, 
    1501142400, 1501146000, 1501149600, 1501153200, 1501156800, 1501160400, 
    1501164000, 1501167600, 1501171200, 1501174800, 1501178400, 1501182000, 
    1501185600, 1501189200, 1501192800, 1501196400, 1501200000, 1501203600, 
    1501207200, 1501210800, 1501214400, 1501218000, 1501221600, 1501225200, 
    1501228800, 1501232400, 1501236000, 1501239600, 1501243200, 1501246800, 
    1501250400, 1501254000, 1501257600, 1501261200, 1501264800, 1501268400, 
    1501272000, 1501275600, 1501279200, 1501282800, 1501286400, 1501290000, 
    1501293600, 1501297200, 1501300800, 1501304400, 1501308000, 1501311600, 
    1501315200, 1501318800, 1501322400, 1501326000, 1501329600, 1501333200, 
    1501336800, 1501340400, 1501344000, 1501347600, 1501351200, 1501354800, 
    1501358400, 1501362000, 1501365600, 1501369200, 1501372800, 1501376400, 
    1501380000, 1501383600, 1501387200, 1501390800, 1501394400, 1501398000, 
    1501401600, 1501405200, 1501408800, 1501412400, 1501416000, 1501419600, 
    1501423200, 1501426800, 1501430400, 1501434000, 1501437600, 1501441200, 
    1501444800, 1501448400, 1501452000, 1501455600, 1501459200, 1501462800, 
    1501466400, 1501470000, 1501473600, 1501477200, 1501480800, 1501484400, 
    1501488000, 1501491600, 1501495200, 1501498800, 1501502400, 1501506000, 
    1501509600, 1501513200, 1501516800, 1501520400, 1501524000, 1501527600, 
    1501531200, 1501534800, 1501538400, 1501542000, 1501545600, 1501549200, 
    1501552800, 1501556400, 1501560000, 1501563600, 1501567200, 1501570800, 
    1501574400, 1501578000, 1501581600, 1501585200, 1501588800, 1501592400, 
    1501596000, 1501599600, 1501603200, 1501606800, 1501610400, 1501614000, 
    1501617600, 1501621200, 1501624800, 1501628400, 1501632000, 1501635600, 
    1501639200, 1501642800, 1501646400, 1501650000, 1501653600, 1501657200, 
    1501660800, 1501664400, 1501668000, 1501671600, 1501675200, 1501678800, 
    1501682400, 1501686000, 1501689600, 1501693200, 1501696800, 1501700400, 
    1501704000, 1501707600, 1501711200, 1501714800, 1501718400, 1501722000, 
    1501725600, 1501729200, 1501732800, 1501736400, 1501740000, 1501743600, 
    1501747200, 1501750800, 1501754400, 1501758000, 1501761600, 1501765200, 
    1501768800, 1501772400, 1501776000, 1501779600, 1501783200, 1501786800, 
    1501790400, 1501794000, 1501797600, 1501801200, 1501804800, 1501808400, 
    1501812000, 1501815600, 1501819200, 1501822800, 1501826400, 1501830000, 
    1501833600, 1501837200, 1501840800, 1501844400, 1501848000, 1501851600, 
    1501855200, 1501858800, 1501862400, 1501866000, 1501869600, 1501873200, 
    1501876800, 1501880400, 1501884000, 1501887600, 1501891200, 1501894800, 
    1501898400, 1501902000, 1501905600, 1501909200, 1501912800, 1501916400, 
    1501920000, 1501923600, 1501927200, 1501930800, 1501934400, 1501938000, 
    1501941600, 1501945200, 1501948800, 1501952400, 1501956000, 1501959600, 
    1501963200, 1501966800, 1501970400, 1501974000, 1501977600, 1501981200, 
    1501984800, 1501988400, 1501992000, 1501995600, 1501999200, 1502002800, 
    1502006400, 1502010000, 1502013600, 1502017200, 1502020800, 1502024400, 
    1502028000, 1502031600, 1502035200, 1502038800, 1502042400, 1502046000, 
    1502049600, 1502053200, 1502056800, 1502060400, 1502064000, 1502067600, 
    1502071200, 1502074800, 1502078400, 1502082000, 1502085600, 1502089200, 
    1502092800, 1502096400, 1502100000, 1502103600, 1502107200, 1502110800, 
    1502114400, 1502118000, 1502121600, 1502125200, 1502128800, 1502132400, 
    1502136000, 1502139600, 1502143200, 1502146800, 1502150400, 1502154000, 
    1502157600, 1502161200, 1502164800, 1502168400, 1502172000, 1502175600, 
    1502179200, 1502182800, 1502186400, 1502190000, 1502193600, 1502197200, 
    1502200800, 1502204400, 1502208000, 1502211600, 1502215200, 1502218800, 
    1502222400, 1502226000, 1502229600, 1502233200, 1502236800, 1502240400, 
    1502244000, 1502247600, 1502251200, 1502254800, 1502258400, 1502262000, 
    1502265600, 1502269200, 1502272800, 1502276400, 1502280000, 1502283600, 
    1502287200, 1502290800, 1502294400, 1502298000, 1502301600, 1502305200, 
    1502308800, 1502312400, 1502316000, 1502319600, 1502323200, 1502326800, 
    1502330400, 1502334000, 1502337600, 1502341200, 1502344800, 1502348400, 
    1502352000, 1502355600, 1502359200, 1502362800, 1502366400, 1502370000, 
    1502373600, 1502377200, 1502380800, 1502384400, 1502388000, 1502391600, 
    1502395200, 1502398800, 1502402400, 1502406000, 1502409600, 1502413200, 
    1502416800, 1502420400, 1502424000, 1502427600, 1502431200, 1502434800, 
    1502438400, 1502442000, 1502445600, 1502449200, 1502452800, 1502456400, 
    1502460000, 1502463600, 1502467200, 1502470800, 1502474400, 1502478000, 
    1502481600, 1502485200, 1502488800, 1502492400, 1502496000, 1502499600, 
    1502503200, 1502506800, 1502510400, 1502514000, 1502517600, 1502521200, 
    1502524800, 1502528400, 1502532000, 1502535600, 1502539200, 1502542800, 
    1502546400, 1502550000, 1502553600, 1502557200, 1502560800, 1502564400, 
    1502568000, 1502571600, 1502575200, 1502578800, 1502582400, 1502586000, 
    1502589600, 1502593200, 1502596800, 1502600400, 1502604000, 1502607600, 
    1502611200, 1502614800, 1502618400, 1502622000, 1502625600, 1502629200, 
    1502632800, 1502636400, 1502640000, 1502643600, 1502647200, 1502650800, 
    1502654400, 1502658000, 1502661600, 1502665200, 1502668800, 1502672400, 
    1502676000, 1502679600, 1502683200, 1502686800, 1502690400, 1502694000, 
    1502697600, 1502701200, 1502704800, 1502708400, 1502712000, 1502715600, 
    1502719200, 1502722800, 1502726400, 1502730000, 1502733600, 1502737200, 
    1502740800, 1502744400, 1502748000, 1502751600, 1502755200, 1502758800, 
    1502762400, 1502766000, 1502769600, 1502773200, 1502776800, 1502780400, 
    1502784000, 1502787600, 1502791200, 1502794800, 1502798400, 1502802000, 
    1502805600, 1502809200, 1502812800, 1502816400, 1502820000, 1502823600, 
    1502827200, 1502830800, 1502834400, 1502838000, 1502841600, 1502845200, 
    1502848800, 1502852400, 1502856000, 1502859600, 1502863200, 1502866800, 
    1502870400, 1502874000, 1502877600, 1502881200, 1502884800, 1502888400, 
    1502892000, 1502895600, 1502899200, 1502902800, 1502906400, 1502910000, 
    1502913600, 1502917200, 1502920800, 1502924400, 1502928000, 1502931600, 
    1502935200, 1502938800, 1502942400, 1502946000, 1502949600, 1502953200, 
    1502956800, 1502960400, 1502964000, 1502967600, 1502971200, 1502974800, 
    1502978400, 1502982000, 1502985600, 1502989200, 1502992800, 1502996400, 
    1503000000, 1503003600, 1503007200, 1503010800, 1503014400, 1503018000, 
    1503021600, 1503025200, 1503028800, 1503032400, 1503036000, 1503039600, 
    1503043200, 1503046800, 1503050400, 1503054000, 1503057600, 1503061200, 
    1503064800, 1503068400, 1503072000, 1503075600, 1503079200, 1503082800, 
    1503086400, 1503090000, 1503093600, 1503097200, 1503100800, 1503104400, 
    1503108000, 1503111600, 1503115200, 1503118800, 1503122400, 1503126000, 
    1503129600, 1503133200, 1503136800, 1503140400, 1503144000, 1503147600, 
    1503151200, 1503154800, 1503158400, 1503162000, 1503165600, 1503169200, 
    1503172800, 1503176400, 1503180000, 1503183600, 1503187200, 1503190800, 
    1503194400, 1503198000, 1503201600, 1503205200, 1503208800, 1503212400, 
    1503216000, 1503219600, 1503223200, 1503226800, 1503230400, 1503234000, 
    1503237600, 1503241200, 1503244800, 1503248400, 1503252000, 1503255600, 
    1503259200, 1503262800, 1503266400, 1503270000, 1503273600, 1503277200, 
    1503280800, 1503284400, 1503288000, 1503291600, 1503295200, 1503298800, 
    1503302400, 1503306000, 1503309600, 1503313200, 1503316800, 1503320400, 
    1503324000, 1503327600, 1503331200, 1503334800, 1503338400, 1503342000, 
    1503345600, 1503349200, 1503352800, 1503356400, 1503360000, 1503363600, 
    1503367200, 1503370800, 1503374400, 1503378000, 1503381600, 1503385200, 
    1503388800, 1503392400, 1503396000, 1503399600, 1503403200, 1503406800, 
    1503410400, 1503414000, 1503417600, 1503421200, 1503424800, 1503428400, 
    1503432000, 1503435600, 1503439200, 1503442800, 1503446400, 1503450000, 
    1503453600, 1503457200, 1503460800, 1503464400, 1503468000, 1503471600, 
    1503475200, 1503478800, 1503482400, 1503486000, 1503489600, 1503493200, 
    1503496800, 1503500400, 1503504000, 1503507600, 1503511200, 1503514800, 
    1503518400, 1503522000, 1503525600, 1503529200, 1503532800, 1503536400, 
    1503540000, 1503543600, 1503547200, 1503550800, 1503554400, 1503558000, 
    1503561600, 1503565200, 1503568800, 1503572400, 1503576000, 1503579600, 
    1503583200, 1503586800, 1503590400, 1503594000, 1503597600, 1503601200, 
    1503604800, 1503608400, 1503612000, 1503615600, 1503619200, 1503622800, 
    1503626400, 1503630000, 1503633600, 1503637200, 1503640800, 1503644400, 
    1503648000, 1503651600, 1503655200, 1503658800, 1503662400, 1503666000, 
    1503669600, 1503673200, 1503676800, 1503680400, 1503684000, 1503687600, 
    1503691200, 1503694800, 1503698400, 1503702000, 1503705600, 1503709200, 
    1503712800, 1503716400, 1503720000, 1503723600, 1503727200, 1503730800, 
    1503734400, 1503738000, 1503741600, 1503745200, 1503748800, 1503752400, 
    1503756000, 1503759600, 1503763200, 1503766800, 1503770400, 1503774000, 
    1503777600, 1503781200, 1503784800, 1503788400, 1503792000, 1503795600, 
    1503799200, 1503802800, 1503806400, 1503810000, 1503813600, 1503817200, 
    1503820800, 1503824400, 1503828000, 1503831600, 1503835200, 1503838800, 
    1503842400, 1503846000, 1503849600, 1503853200, 1503856800, 1503860400, 
    1503864000, 1503867600, 1503871200, 1503874800, 1503878400, 1503882000, 
    1503885600, 1503889200, 1503892800, 1503896400, 1503900000, 1503903600, 
    1503907200, 1503910800, 1503914400, 1503918000, 1503921600, 1503925200, 
    1503928800, 1503932400, 1503936000, 1503939600, 1503943200, 1503946800, 
    1503950400, 1503954000, 1503957600, 1503961200, 1503964800, 1503968400, 
    1503972000, 1503975600, 1503979200, 1503982800, 1503986400, 1503990000, 
    1503993600, 1503997200, 1504000800, 1504004400, 1504008000, 1504011600, 
    1504015200, 1504018800, 1504022400, 1504026000, 1504029600, 1504033200, 
    1504036800, 1504040400, 1504044000, 1504047600, 1504051200, 1504054800, 
    1504058400, 1504062000, 1504065600, 1504069200, 1504072800, 1504076400, 
    1504080000, 1504083600, 1504087200, 1504090800, 1504094400, 1504098000, 
    1504101600, 1504105200, 1504108800, 1504112400, 1504116000, 1504119600, 
    1504123200, 1504126800, 1504130400, 1504134000, 1504137600, 1504141200, 
    1504144800, 1504148400, 1504152000, 1504155600, 1504159200, 1504162800, 
    1504166400, 1504170000, 1504173600, 1504177200, 1504180800, 1504184400, 
    1504188000, 1504191600, 1504195200, 1504198800, 1504202400, 1504206000, 
    1504209600, 1504213200, 1504216800, 1504220400, 1504224000, 1504227600, 
    1504231200, 1504234800, 1504238400, 1504242000, 1504245600, 1504249200, 
    1504252800, 1504256400, 1504260000, 1504263600, 1504267200, 1504270800, 
    1504274400, 1504278000, 1504281600, 1504285200, 1504288800, 1504292400, 
    1504296000, 1504299600, 1504303200, 1504306800, 1504310400, 1504314000, 
    1504317600, 1504321200, 1504324800, 1504328400, 1504332000, 1504335600, 
    1504339200, 1504342800, 1504346400, 1504350000, 1504353600, 1504357200, 
    1504360800, 1504364400, 1504368000, 1504371600, 1504375200, 1504378800, 
    1504382400, 1504386000, 1504389600, 1504393200, 1504396800, 1504400400, 
    1504404000, 1504407600, 1504411200, 1504414800, 1504418400, 1504422000, 
    1504425600, 1504429200, 1504432800, 1504436400, 1504440000, 1504443600, 
    1504447200, 1504450800, 1504454400, 1504458000, 1504461600, 1504465200, 
    1504468800, 1504472400, 1504476000, 1504479600, 1504483200, 1504486800, 
    1504490400, 1504494000, 1504497600, 1504501200, 1504504800, 1504508400, 
    1504512000, 1504515600, 1504519200, 1504522800, 1504526400, 1504530000, 
    1504533600, 1504537200, 1504540800, 1504544400, 1504548000, 1504551600, 
    1504555200, 1504558800, 1504562400, 1504566000, 1504569600, 1504573200, 
    1504576800, 1504580400, 1504584000, 1504587600, 1504591200, 1504594800, 
    1504598400, 1504602000, 1504605600, 1504609200, 1504612800, 1504616400, 
    1504620000, 1504623600, 1504627200, 1504630800, 1504634400, 1504638000, 
    1504641600, 1504645200, 1504648800, 1504652400, 1504656000, 1504659600, 
    1504663200, 1504666800, 1504670400, 1504674000, 1504677600, 1504681200, 
    1504684800, 1504688400, 1504692000, 1504695600, 1504699200, 1504702800, 
    1504706400, 1504710000, 1504713600, 1504717200, 1504720800, 1504724400, 
    1504728000, 1504731600, 1504735200, 1504738800, 1504742400, 1504746000, 
    1504749600, 1504753200, 1504756800, 1504760400, 1504764000, 1504767600, 
    1504771200, 1504774800, 1504778400, 1504782000, 1504785600, 1504789200, 
    1504792800, 1504796400, 1504800000, 1504803600, 1504807200, 1504810800, 
    1504814400, 1504818000, 1504821600, 1504825200, 1504828800, 1504832400, 
    1504836000, 1504839600, 1504843200, 1504846800, 1504850400, 1504854000, 
    1504857600, 1504861200, 1504864800, 1504868400, 1504872000, 1504875600, 
    1504879200, 1504882800, 1504886400, 1504890000, 1504893600, 1504897200, 
    1504900800, 1504904400, 1504908000, 1504911600, 1504915200, 1504918800, 
    1504922400, 1504926000, 1504929600, 1504933200, 1504936800, 1504940400, 
    1504944000, 1504947600, 1504951200, 1504954800, 1504958400, 1504962000, 
    1504965600, 1504969200, 1504972800, 1504976400, 1504980000, 1504983600, 
    1504987200, 1504990800, 1504994400, 1504998000, 1505001600, 1505005200, 
    1505008800, 1505012400, 1505016000, 1505019600, 1505023200, 1505026800, 
    1505030400, 1505034000, 1505037600, 1505041200, 1505044800, 1505048400, 
    1505052000, 1505055600, 1505059200, 1505062800, 1505066400, 1505070000, 
    1505073600, 1505077200, 1505080800, 1505084400, 1505088000, 1505091600, 
    1505095200, 1505098800, 1505102400, 1505106000, 1505109600, 1505113200, 
    1505116800, 1505120400, 1505124000, 1505127600, 1505131200, 1505134800, 
    1505138400, 1505142000, 1505145600, 1505149200, 1505152800, 1505156400, 
    1505160000, 1505163600, 1505167200, 1505170800, 1505174400, 1505178000, 
    1505181600, 1505185200, 1505188800, 1505192400, 1505196000, 1505199600, 
    1505203200, 1505206800, 1505210400, 1505214000, 1505217600, 1505221200, 
    1505224800, 1505228400, 1505232000, 1505235600, 1505239200, 1505242800, 
    1505246400, 1505250000, 1505253600, 1505257200, 1505260800, 1505264400, 
    1505268000, 1505271600, 1505275200, 1505278800, 1505282400, 1505286000, 
    1505289600, 1505293200, 1505296800, 1505300400, 1505304000, 1505307600, 
    1505311200, 1505314800, 1505318400, 1505322000, 1505325600, 1505329200, 
    1505332800, 1505336400, 1505340000, 1505343600, 1505347200, 1505350800, 
    1505354400, 1505358000, 1505361600, 1505365200, 1505368800, 1505372400, 
    1505376000, 1505379600, 1505383200, 1505386800, 1505390400, 1505394000, 
    1505397600, 1505401200, 1505404800, 1505408400, 1505412000, 1505415600, 
    1505419200, 1505422800, 1505426400, 1505430000, 1505433600, 1505437200, 
    1505440800, 1505444400, 1505448000, 1505451600, 1505455200, 1505458800, 
    1505462400, 1505466000, 1505469600, 1505473200, 1505476800, 1505480400, 
    1505484000, 1505487600, 1505491200, 1505494800, 1505498400, 1505502000, 
    1505505600, 1505509200, 1505512800, 1505516400, 1505520000, 1505523600, 
    1505527200, 1505530800, 1505534400, 1505538000, 1505541600, 1505545200, 
    1505548800, 1505552400, 1505556000, 1505559600, 1505563200, 1505566800, 
    1505570400, 1505574000, 1505577600, 1505581200, 1505584800, 1505588400, 
    1505592000, 1505595600, 1505599200, 1505602800, 1505606400, 1505610000, 
    1505613600, 1505617200, 1505620800, 1505624400, 1505628000, 1505631600, 
    1505635200, 1505638800, 1505642400, 1505646000, 1505649600, 1505653200, 
    1505656800, 1505660400, 1505664000, 1505667600, 1505671200, 1505674800, 
    1505678400, 1505682000, 1505685600, 1505689200, 1505692800, 1505696400, 
    1505700000, 1505703600, 1505707200, 1505710800, 1505714400, 1505718000, 
    1505721600, 1505725200, 1505728800, 1505732400, 1505736000, 1505739600, 
    1505743200, 1505746800, 1505750400, 1505754000, 1505757600, 1505761200, 
    1505764800, 1505768400, 1505772000, 1505775600, 1505779200, 1505782800, 
    1505786400, 1505790000, 1505793600, 1505797200, 1505800800, 1505804400, 
    1505808000, 1505811600, 1505815200, 1505818800, 1505822400, 1505826000, 
    1505829600, 1505833200, 1505836800, 1505840400, 1505844000, 1505847600, 
    1505851200, 1505854800, 1505858400, 1505862000, 1505865600, 1505869200, 
    1505872800, 1505876400, 1505880000, 1505883600, 1505887200, 1505890800, 
    1505894400, 1505898000, 1505901600, 1505905200, 1505908800, 1505912400, 
    1505916000, 1505919600, 1505923200, 1505926800, 1505930400, 1505934000, 
    1505937600, 1505941200, 1505944800, 1505948400, 1505952000, 1505955600, 
    1505959200, 1505962800, 1505966400, 1505970000, 1505973600, 1505977200, 
    1505980800, 1505984400, 1505988000, 1505991600, 1505995200, 1505998800, 
    1506002400, 1506006000, 1506009600, 1506013200, 1506016800, 1506020400, 
    1506024000, 1506027600, 1506031200, 1506034800, 1506038400, 1506042000, 
    1506045600, 1506049200, 1506052800, 1506056400, 1506060000, 1506063600, 
    1506067200, 1506070800, 1506074400, 1506078000, 1506081600, 1506085200, 
    1506088800, 1506092400, 1506096000, 1506099600, 1506103200, 1506106800, 
    1506110400, 1506114000, 1506117600, 1506121200, 1506124800, 1506128400, 
    1506132000, 1506135600, 1506139200, 1506142800, 1506146400, 1506150000, 
    1506153600, 1506157200, 1506160800, 1506164400, 1506168000, 1506171600, 
    1506175200, 1506178800, 1506182400, 1506186000, 1506189600, 1506193200, 
    1506196800, 1506200400, 1506204000, 1506207600, 1506211200, 1506214800, 
    1506218400, 1506222000, 1506225600, 1506229200, 1506232800, 1506236400, 
    1506240000, 1506243600, 1506247200, 1506250800, 1506254400, 1506258000, 
    1506261600, 1506265200, 1506268800, 1506272400, 1506276000, 1506279600, 
    1506283200, 1506286800, 1506290400, 1506294000, 1506297600, 1506301200, 
    1506304800, 1506308400, 1506312000, 1506315600, 1506319200, 1506322800, 
    1506326400, 1506330000, 1506333600, 1506337200, 1506340800, 1506344400, 
    1506348000, 1506351600, 1506355200, 1506358800, 1506362400, 1506366000, 
    1506369600, 1506373200, 1506376800, 1506380400, 1506384000, 1506387600, 
    1506391200, 1506394800, 1506398400, 1506402000, 1506405600, 1506409200, 
    1506412800, 1506416400, 1506420000, 1506423600, 1506427200, 1506430800, 
    1506434400, 1506438000, 1506441600, 1506445200, 1506448800, 1506452400, 
    1506456000, 1506459600, 1506463200, 1506466800, 1506470400, 1506474000, 
    1506477600, 1506481200, 1506484800, 1506488400, 1506492000, 1506495600, 
    1506499200, 1506502800, 1506506400, 1506510000, 1506513600, 1506517200, 
    1506520800, 1506524400, 1506528000, 1506531600, 1506535200, 1506538800, 
    1506542400, 1506546000, 1506549600, 1506553200, 1506556800, 1506560400, 
    1506564000, 1506567600, 1506571200, 1506574800, 1506578400, 1506582000, 
    1506585600, 1506589200, 1506592800, 1506596400, 1506600000, 1506603600, 
    1506607200, 1506610800, 1506614400, 1506618000, 1506621600, 1506625200, 
    1506628800, 1506632400, 1506636000, 1506639600, 1506643200, 1506646800, 
    1506650400, 1506654000, 1506657600, 1506661200, 1506664800, 1506668400, 
    1506672000, 1506675600, 1506679200, 1506682800, 1506686400, 1506690000, 
    1506693600, 1506697200, 1506700800, 1506704400, 1506708000, 1506711600, 
    1506715200, 1506718800, 1506722400, 1506726000, 1506729600, 1506733200, 
    1506736800, 1506740400, 1506744000, 1506747600, 1506751200, 1506754800, 
    1506758400, 1506762000, 1506765600, 1506769200, 1506772800, 1506776400, 
    1506780000, 1506783600, 1506787200, 1506790800, 1506794400, 1506798000, 
    1506801600, 1506805200, 1506808800, 1506812400, 1506816000, 1506819600, 
    1506823200, 1506826800, 1506830400, 1506834000, 1506837600, 1506841200, 
    1506844800, 1506848400, 1506852000, 1506855600, 1506859200, 1506862800, 
    1506866400, 1506870000, 1506873600, 1506877200, 1506880800, 1506884400, 
    1506888000, 1506891600, 1506895200, 1506898800, 1506902400, 1506906000, 
    1506909600, 1506913200, 1506916800, 1506920400, 1506924000, 1506927600, 
    1506931200, 1506934800, 1506938400, 1506942000, 1506945600, 1506949200, 
    1506952800, 1506956400, 1506960000, 1506963600, 1506967200, 1506970800, 
    1506974400, 1506978000, 1506981600, 1506985200, 1506988800, 1506992400, 
    1506996000, 1506999600, 1507003200, 1507006800, 1507010400, 1507014000, 
    1507017600, 1507021200, 1507024800, 1507028400, 1507032000, 1507035600, 
    1507039200, 1507042800, 1507046400, 1507050000, 1507053600, 1507057200, 
    1507060800, 1507064400, 1507068000, 1507071600, 1507075200, 1507078800, 
    1507082400, 1507086000, 1507089600, 1507093200, 1507096800, 1507100400, 
    1507104000, 1507107600, 1507111200, 1507114800, 1507118400, 1507122000, 
    1507125600, 1507129200, 1507132800, 1507136400, 1507140000, 1507143600, 
    1507147200, 1507150800, 1507154400, 1507158000, 1507161600, 1507165200, 
    1507168800, 1507172400, 1507176000, 1507179600, 1507183200, 1507186800, 
    1507190400, 1507194000, 1507197600, 1507201200, 1507204800, 1507208400, 
    1507212000, 1507215600, 1507219200, 1507222800, 1507226400, 1507230000, 
    1507233600, 1507237200, 1507240800, 1507244400, 1507248000, 1507251600, 
    1507255200, 1507258800, 1507262400, 1507266000, 1507269600, 1507273200, 
    1507276800, 1507280400, 1507284000, 1507287600, 1507291200, 1507294800, 
    1507298400, 1507302000, 1507305600, 1507309200, 1507312800, 1507316400, 
    1507320000, 1507323600, 1507327200, 1507330800, 1507334400, 1507338000, 
    1507341600, 1507345200, 1507348800, 1507352400, 1507356000, 1507359600, 
    1507363200, 1507366800, 1507370400, 1507374000, 1507377600, 1507381200, 
    1507384800, 1507388400, 1507392000, 1507395600, 1507399200, 1507402800, 
    1507406400, 1507410000, 1507413600, 1507417200, 1507420800, 1507424400, 
    1507428000, 1507431600, 1507435200, 1507438800, 1507442400, 1507446000, 
    1507449600, 1507453200, 1507456800, 1507460400, 1507464000, 1507467600, 
    1507471200, 1507474800, 1507478400, 1507482000, 1507485600, 1507489200, 
    1507492800, 1507496400, 1507500000, 1507503600, 1507507200, 1507510800, 
    1507514400, 1507518000, 1507521600, 1507525200, 1507528800, 1507532400, 
    1507536000, 1507539600, 1507543200, 1507546800, 1507550400, 1507554000, 
    1507557600, 1507561200, 1507564800, 1507568400, 1507572000, 1507575600, 
    1507579200, 1507582800, 1507586400, 1507590000, 1507593600, 1507597200, 
    1507600800, 1507604400, 1507608000, 1507611600, 1507615200, 1507618800, 
    1507622400, 1507626000, 1507629600, 1507633200, 1507636800, 1507640400, 
    1507644000, 1507647600, 1507651200, 1507654800, 1507658400, 1507662000, 
    1507665600, 1507669200, 1507672800, 1507676400, 1507680000, 1507683600, 
    1507687200, 1507690800, 1507694400, 1507698000, 1507701600, 1507705200, 
    1507708800, 1507712400, 1507716000, 1507719600, 1507723200, 1507726800, 
    1507730400, 1507734000, 1507737600, 1507741200, 1507744800, 1507748400, 
    1507752000, 1507755600, 1507759200, 1507762800, 1507766400, 1507770000, 
    1507773600, 1507777200, 1507780800, 1507784400, 1507788000, 1507791600, 
    1507795200, 1507798800, 1507802400, 1507806000, 1507809600, 1507813200, 
    1507816800, 1507820400, 1507824000, 1507827600, 1507831200, 1507834800, 
    1507838400, 1507842000, 1507845600, 1507849200, 1507852800, 1507856400, 
    1507860000, 1507863600, 1507867200, 1507870800, 1507874400, 1507878000, 
    1507881600, 1507885200, 1507888800, 1507892400, 1507896000, 1507899600, 
    1507903200, 1507906800, 1507910400, 1507914000, 1507917600, 1507921200, 
    1507924800, 1507928400, 1507932000, 1507935600, 1507939200, 1507942800, 
    1507946400, 1507950000, 1507953600, 1507957200, 1507960800, 1507964400, 
    1507968000, 1507971600, 1507975200, 1507978800, 1507982400, 1507986000, 
    1507989600, 1507993200, 1507996800, 1508000400, 1508004000, 1508007600, 
    1508011200, 1508014800, 1508018400, 1508022000, 1508025600, 1508029200, 
    1508032800, 1508036400, 1508040000, 1508043600, 1508047200, 1508050800, 
    1508054400, 1508058000, 1508061600, 1508065200, 1508068800, 1508072400, 
    1508076000, 1508079600, 1508083200, 1508086800, 1508090400, 1508094000, 
    1508097600, 1508101200, 1508104800, 1508108400, 1508112000, 1508115600, 
    1508119200, 1508122800, 1508126400, 1508130000, 1508133600, 1508137200, 
    1508140800, 1508144400, 1508148000, 1508151600, 1508155200, 1508158800, 
    1508162400, 1508166000, 1508169600, 1508173200, 1508176800, 1508180400, 
    1508184000, 1508187600, 1508191200, 1508194800, 1508198400, 1508202000, 
    1508205600, 1508209200, 1508212800, 1508216400, 1508220000, 1508223600, 
    1508227200, 1508230800, 1508234400, 1508238000, 1508241600, 1508245200, 
    1508248800, 1508252400, 1508256000, 1508259600, 1508263200, 1508266800, 
    1508270400, 1508274000, 1508277600, 1508281200, 1508284800, 1508288400, 
    1508292000, 1508295600, 1508299200, 1508302800, 1508306400, 1508310000, 
    1508313600, 1508317200, 1508320800, 1508324400, 1508328000, 1508331600, 
    1508335200, 1508338800, 1508342400, 1508346000, 1508349600, 1508353200, 
    1508356800, 1508360400, 1508364000, 1508367600, 1508371200, 1508374800, 
    1508378400, 1508382000, 1508385600, 1508389200, 1508392800, 1508396400, 
    1508400000, 1508403600, 1508407200, 1508410800, 1508414400, 1508418000, 
    1508421600, 1508425200, 1508428800, 1508432400, 1508436000, 1508439600, 
    1508443200, 1508446800, 1508450400, 1508454000, 1508457600, 1508461200, 
    1508464800, 1508468400, 1508472000, 1508475600, 1508479200, 1508482800, 
    1508486400, 1508490000, 1508493600, 1508497200, 1508500800, 1508504400, 
    1508508000, 1508511600, 1508515200, 1508518800, 1508522400, 1508526000, 
    1508529600, 1508533200, 1508536800, 1508540400, 1508544000, 1508547600, 
    1508551200, 1508554800, 1508558400, 1508562000, 1508565600, 1508569200, 
    1508572800, 1508576400, 1508580000, 1508583600, 1508587200, 1508590800, 
    1508594400, 1508598000, 1508601600, 1508605200, 1508608800, 1508612400, 
    1508616000, 1508619600, 1508623200, 1508626800, 1508630400, 1508634000, 
    1508637600, 1508641200, 1508644800, 1508648400, 1508652000, 1508655600, 
    1508659200, 1508662800, 1508666400, 1508670000, 1508673600, 1508677200, 
    1508680800, 1508684400, 1508688000, 1508691600, 1508695200, 1508698800, 
    1508702400, 1508706000, 1508709600, 1508713200, 1508716800, 1508720400, 
    1508724000, 1508727600, 1508731200, 1508734800, 1508738400, 1508742000, 
    1508745600, 1508749200, 1508752800, 1508756400, 1508760000, 1508763600, 
    1508767200, 1508770800, 1508774400, 1508778000, 1508781600, 1508785200, 
    1508788800, 1508792400, 1508796000, 1508799600, 1508803200, 1508806800, 
    1508810400, 1508814000, 1508817600, 1508821200, 1508824800, 1508828400, 
    1508832000, 1508835600, 1508839200, 1508842800, 1508846400, 1508850000, 
    1508853600, 1508857200, 1508860800, 1508864400, 1508868000, 1508871600, 
    1508875200, 1508878800, 1508882400, 1508886000, 1508889600, 1508893200, 
    1508896800, 1508900400, 1508904000, 1508907600, 1508911200, 1508914800, 
    1508918400, 1508922000, 1508925600, 1508929200, 1508932800, 1508936400, 
    1508940000, 1508943600, 1508947200, 1508950800, 1508954400, 1508958000, 
    1508961600, 1508965200, 1508968800, 1508972400, 1508976000, 1508979600, 
    1508983200, 1508986800, 1508990400, 1508994000, 1508997600, 1509001200, 
    1509004800, 1509008400, 1509012000, 1509015600, 1509019200, 1509022800, 
    1509026400, 1509030000, 1509033600, 1509037200, 1509040800, 1509044400, 
    1509048000, 1509051600, 1509055200, 1509058800, 1509062400, 1509066000, 
    1509069600, 1509073200, 1509076800, 1509080400, 1509084000, 1509087600, 
    1509091200, 1509094800, 1509098400, 1509102000, 1509105600, 1509109200, 
    1509112800, 1509116400, 1509120000, 1509123600, 1509127200, 1509130800, 
    1509134400, 1509138000, 1509141600, 1509145200, 1509148800, 1509152400, 
    1509156000, 1509159600, 1509163200, 1509166800, 1509170400, 1509174000, 
    1509177600, 1509181200, 1509184800, 1509188400, 1509192000, 1509195600, 
    1509199200, 1509202800, 1509206400, 1509210000, 1509213600, 1509217200, 
    1509220800, 1509224400, 1509228000, 1509231600, 1509235200, 1509238800, 
    1509242400, 1509246000, 1509249600, 1509253200, 1509256800, 1509260400, 
    1509264000, 1509267600, 1509271200, 1509274800, 1509278400, 1509282000, 
    1509285600, 1509289200, 1509292800, 1509296400, 1509300000, 1509303600, 
    1509307200, 1509310800, 1509314400, 1509318000, 1509321600, 1509325200, 
    1509328800, 1509332400, 1509336000, 1509339600, 1509343200, 1509346800, 
    1509350400, 1509354000, 1509357600, 1509361200, 1509364800, 1509368400, 
    1509372000, 1509375600, 1509379200, 1509382800, 1509386400, 1509390000, 
    1509393600, 1509397200, 1509400800, 1509404400, 1509408000, 1509411600, 
    1509415200, 1509418800, 1509422400, 1509426000, 1509429600, 1509433200, 
    1509436800, 1509440400, 1509444000, 1509447600, 1509451200, 1509454800, 
    1509458400, 1509462000, 1509465600, 1509469200, 1509472800, 1509476400, 
    1509480000, 1509483600, 1509487200, 1509490800, 1509494400, 1509498000, 
    1509501600, 1509505200, 1509508800, 1509512400, 1509516000, 1509519600, 
    1509523200, 1509526800, 1509530400, 1509534000, 1509537600, 1509541200, 
    1509544800, 1509548400, 1509552000, 1509555600, 1509559200, 1509562800, 
    1509566400, 1509570000, 1509573600, 1509577200, 1509580800, 1509584400, 
    1509588000, 1509591600, 1509595200, 1509598800, 1509602400, 1509606000, 
    1509609600, 1509613200, 1509616800, 1509620400, 1509624000, 1509627600, 
    1509631200, 1509634800, 1509638400, 1509642000, 1509645600, 1509649200, 
    1509652800, 1509656400, 1509660000, 1509663600, 1509667200, 1509670800, 
    1509674400, 1509678000, 1509681600, 1509685200, 1509688800, 1509692400, 
    1509696000, 1509699600, 1509703200, 1509706800, 1509710400, 1509714000, 
    1509717600, 1509721200, 1509724800, 1509728400, 1509732000, 1509735600, 
    1509739200, 1509742800, 1509746400, 1509750000, 1509753600, 1509757200, 
    1509760800, 1509764400, 1509768000, 1509771600, 1509775200, 1509778800, 
    1509782400, 1509786000, 1509789600, 1509793200, 1509796800, 1509800400, 
    1509804000, 1509807600, 1509811200, 1509814800, 1509818400, 1509822000, 
    1509825600, 1509829200, 1509832800, 1509836400, 1509840000, 1509843600, 
    1509847200, 1509850800, 1509854400, 1509858000, 1509861600, 1509865200, 
    1509868800, 1509872400, 1509876000, 1509879600, 1509883200, 1509886800, 
    1509890400, 1509894000, 1509897600, 1509901200, 1509904800, 1509908400, 
    1509912000, 1509915600, 1509919200, 1509922800, 1509926400, 1509930000, 
    1509933600, 1509937200, 1509940800, 1509944400, 1509948000, 1509951600, 
    1509955200, 1509958800, 1509962400, 1509966000, 1509969600, 1509973200, 
    1509976800, 1509980400, 1509984000, 1509987600, 1509991200, 1509994800, 
    1509998400, 1510002000, 1510005600, 1510009200, 1510012800, 1510016400, 
    1510020000, 1510023600, 1510027200, 1510030800, 1510034400, 1510038000, 
    1510041600, 1510045200, 1510048800, 1510052400, 1510056000, 1510059600, 
    1510063200, 1510066800, 1510070400, 1510074000, 1510077600, 1510081200, 
    1510084800, 1510088400, 1510092000, 1510095600, 1510099200, 1510102800, 
    1510106400, 1510110000, 1510113600, 1510117200, 1510120800, 1510124400, 
    1510128000, 1510131600, 1510135200, 1510138800, 1510142400, 1510146000, 
    1510149600, 1510153200, 1510156800, 1510160400, 1510164000, 1510167600, 
    1510171200, 1510174800, 1510178400, 1510182000, 1510185600, 1510189200, 
    1510192800, 1510196400, 1510200000, 1510203600, 1510207200, 1510210800, 
    1510214400, 1510218000, 1510221600, 1510225200, 1510228800, 1510232400, 
    1510236000, 1510239600, 1510243200, 1510246800, 1510250400, 1510254000, 
    1510257600, 1510261200, 1510264800, 1510268400, 1510272000, 1510275600, 
    1510279200, 1510282800, 1510286400, 1510290000, 1510293600, 1510297200, 
    1510300800, 1510304400, 1510308000, 1510311600, 1510315200, 1510318800, 
    1510322400, 1510326000, 1510329600, 1510333200, 1510336800, 1510340400, 
    1510344000, 1510347600, 1510351200, 1510354800, 1510358400, 1510362000, 
    1510365600, 1510369200, 1510372800, 1510376400, 1510380000, 1510383600, 
    1510387200, 1510390800, 1510394400, 1510398000, 1510401600, 1510405200, 
    1510408800, 1510412400, 1510416000, 1510419600, 1510423200, 1510426800, 
    1510430400, 1510434000, 1510437600, 1510441200, 1510444800, 1510448400, 
    1510452000, 1510455600, 1510459200, 1510462800, 1510466400, 1510470000, 
    1510473600, 1510477200, 1510480800, 1510484400, 1510488000, 1510491600, 
    1510495200, 1510498800, 1510502400, 1510506000, 1510509600, 1510513200, 
    1510516800, 1510520400, 1510524000, 1510527600, 1510531200, 1510534800, 
    1510538400, 1510542000, 1510545600, 1510549200, 1510552800, 1510556400, 
    1510560000, 1510563600, 1510567200, 1510570800, 1510574400, 1510578000, 
    1510581600, 1510585200, 1510588800, 1510592400, 1510596000, 1510599600, 
    1510603200, 1510606800, 1510610400, 1510614000, 1510617600, 1510621200, 
    1510624800, 1510628400, 1510632000, 1510635600, 1510639200, 1510642800, 
    1510646400, 1510650000, 1510653600, 1510657200, 1510660800, 1510664400, 
    1510668000, 1510671600, 1510675200, 1510678800, 1510682400, 1510686000, 
    1510689600, 1510693200, 1510696800, 1510700400, 1510704000, 1510707600, 
    1510711200, 1510714800, 1510718400, 1510722000, 1510725600, 1510729200, 
    1510732800, 1510736400, 1510740000, 1510743600, 1510747200, 1510750800, 
    1510754400, 1510758000, 1510761600, 1510765200, 1510768800, 1510772400, 
    1510776000, 1510779600, 1510783200, 1510786800, 1510790400, 1510794000, 
    1510797600, 1510801200, 1510804800, 1510808400, 1510812000, 1510815600, 
    1510819200, 1510822800, 1510826400, 1510830000, 1510833600, 1510837200, 
    1510840800, 1510844400, 1510848000, 1510851600, 1510855200, 1510858800, 
    1510862400, 1510866000, 1510869600, 1510873200, 1510876800, 1510880400, 
    1510884000, 1510887600, 1510891200, 1510894800, 1510898400, 1510902000, 
    1510905600, 1510909200, 1510912800, 1510916400, 1510920000, 1510923600, 
    1510927200, 1510930800, 1510934400, 1510938000, 1510941600, 1510945200, 
    1510948800, 1510952400, 1510956000, 1510959600, 1510963200, 1510966800, 
    1510970400, 1510974000, 1510977600, 1510981200, 1510984800, 1510988400, 
    1510992000, 1510995600, 1510999200, 1511002800, 1511006400, 1511010000, 
    1511013600, 1511017200, 1511020800, 1511024400, 1511028000, 1511031600, 
    1511035200, 1511038800, 1511042400, 1511046000, 1511049600, 1511053200, 
    1511056800, 1511060400, 1511064000, 1511067600, 1511071200, 1511074800, 
    1511078400, 1511082000, 1511085600, 1511089200, 1511092800, 1511096400, 
    1511100000, 1511103600, 1511107200, 1511110800, 1511114400, 1511118000, 
    1511121600, 1511125200, 1511128800, 1511132400, 1511136000, 1511139600, 
    1511143200, 1511146800, 1511150400, 1511154000, 1511157600, 1511161200, 
    1511164800, 1511168400, 1511172000, 1511175600, 1511179200, 1511182800, 
    1511186400, 1511190000, 1511193600, 1511197200, 1511200800, 1511204400, 
    1511208000, 1511211600, 1511215200, 1511218800, 1511222400, 1511226000, 
    1511229600, 1511233200, 1511236800, 1511240400, 1511244000, 1511247600, 
    1511251200, 1511254800, 1511258400, 1511262000, 1511265600, 1511269200, 
    1511272800, 1511276400, 1511280000, 1511283600, 1511287200, 1511290800, 
    1511294400, 1511298000, 1511301600, 1511305200, 1511308800, 1511312400, 
    1511316000, 1511319600, 1511323200, 1511326800, 1511330400, 1511334000, 
    1511337600, 1511341200, 1511344800, 1511348400, 1511352000, 1511355600, 
    1511359200, 1511362800, 1511366400, 1511370000, 1511373600, 1511377200, 
    1511380800, 1511384400, 1511388000, 1511391600, 1511395200, 1511398800, 
    1511402400, 1511406000, 1511409600, 1511413200, 1511416800, 1511420400, 
    1511424000, 1511427600, 1511431200, 1511434800, 1511438400, 1511442000, 
    1511445600, 1511449200, 1511452800, 1511456400, 1511460000, 1511463600, 
    1511467200, 1511470800, 1511474400, 1511478000, 1511481600, 1511485200, 
    1511488800, 1511492400, 1511496000, 1511499600, 1511503200, 1511506800, 
    1511510400, 1511514000, 1511517600, 1511521200, 1511524800, 1511528400, 
    1511532000, 1511535600, 1511539200, 1511542800, 1511546400, 1511550000, 
    1511553600, 1511557200, 1511560800, 1511564400, 1511568000, 1511571600, 
    1511575200, 1511578800, 1511582400, 1511586000, 1511589600, 1511593200, 
    1511596800, 1511600400, 1511604000, 1511607600, 1511611200, 1511614800, 
    1511618400, 1511622000, 1511625600, 1511629200, 1511632800, 1511636400, 
    1511640000, 1511643600, 1511647200, 1511650800, 1511654400, 1511658000, 
    1511661600, 1511665200, 1511668800, 1511672400, 1511676000, 1511679600, 
    1511683200, 1511686800, 1511690400, 1511694000, 1511697600, 1511701200, 
    1511704800, 1511708400, 1511712000, 1511715600, 1511719200, 1511722800, 
    1511726400, 1511730000, 1511733600, 1511737200, 1511740800, 1511744400, 
    1511748000, 1511751600, 1511755200, 1511758800, 1511762400, 1511766000, 
    1511769600, 1511773200, 1511776800, 1511780400, 1511784000, 1511787600, 
    1511791200, 1511794800, 1511798400, 1511802000, 1511805600, 1511809200, 
    1511812800, 1511816400, 1511820000, 1511823600, 1511827200, 1511830800, 
    1511834400, 1511838000, 1511841600, 1511845200, 1511848800, 1511852400, 
    1511856000, 1511859600, 1511863200, 1511866800, 1511870400, 1511874000, 
    1511877600, 1511881200, 1511884800, 1511888400, 1511892000, 1511895600, 
    1511899200, 1511902800, 1511906400, 1511910000, 1511913600, 1511917200, 
    1511920800, 1511924400, 1511928000, 1511931600, 1511935200, 1511938800, 
    1511942400, 1511946000, 1511949600, 1511953200, 1511956800, 1511960400, 
    1511964000, 1511967600, 1511971200, 1511974800, 1511978400, 1511982000, 
    1511985600, 1511989200, 1511992800, 1511996400, 1512000000, 1512003600, 
    1512007200, 1512010800, 1512014400, 1512018000, 1512021600, 1512025200, 
    1512028800, 1512032400, 1512036000, 1512039600, 1512043200, 1512046800, 
    1512050400, 1512054000, 1512057600, 1512061200, 1512064800, 1512068400, 
    1512072000, 1512075600, 1512079200, 1512082800, 1512086400, 1512090000, 
    1512093600, 1512097200, 1512100800, 1512104400, 1512108000, 1512111600, 
    1512115200, 1512118800, 1512122400, 1512126000, 1512129600, 1512133200, 
    1512136800, 1512140400, 1512144000, 1512147600, 1512151200, 1512154800, 
    1512158400, 1512162000, 1512165600, 1512169200, 1512172800, 1512176400, 
    1512180000, 1512183600, 1512187200, 1512190800, 1512194400, 1512198000, 
    1512201600, 1512205200, 1512208800, 1512212400, 1512216000, 1512219600, 
    1512223200, 1512226800, 1512230400, 1512234000, 1512237600, 1512241200, 
    1512244800, 1512248400, 1512252000, 1512255600, 1512259200, 1512262800, 
    1512266400, 1512270000, 1512273600, 1512277200, 1512280800, 1512284400, 
    1512288000, 1512291600, 1512295200, 1512298800, 1512302400, 1512306000, 
    1512309600, 1512313200, 1512316800, 1512320400, 1512324000, 1512327600, 
    1512331200, 1512334800, 1512338400, 1512342000, 1512345600, 1512349200, 
    1512352800, 1512356400, 1512360000, 1512363600, 1512367200, 1512370800, 
    1512374400, 1512378000, 1512381600, 1512385200, 1512388800, 1512392400, 
    1512396000, 1512399600, 1512403200, 1512406800, 1512410400, 1512414000, 
    1512417600, 1512421200, 1512424800, 1512428400, 1512432000, 1512435600, 
    1512439200, 1512442800, 1512446400, 1512450000, 1512453600, 1512457200, 
    1512460800, 1512464400, 1512468000, 1512471600, 1512475200, 1512478800, 
    1512482400, 1512486000, 1512489600, 1512493200, 1512496800, 1512500400, 
    1512504000, 1512507600, 1512511200, 1512514800, 1512518400, 1512522000, 
    1512525600, 1512529200, 1512532800, 1512536400, 1512540000, 1512543600, 
    1512547200, 1512550800, 1512554400, 1512558000, 1512561600, 1512565200, 
    1512568800, 1512572400, 1512576000, 1512579600, 1512583200, 1512586800, 
    1512590400, 1512594000, 1512597600, 1512601200, 1512604800, 1512608400, 
    1512612000, 1512615600, 1512619200, 1512622800, 1512626400, 1512630000, 
    1512633600, 1512637200, 1512640800, 1512644400, 1512648000, 1512651600, 
    1512655200, 1512658800, 1512662400, 1512666000, 1512669600, 1512673200, 
    1512676800, 1512680400, 1512684000, 1512687600, 1512691200, 1512694800, 
    1512698400, 1512702000, 1512705600, 1512709200, 1512712800, 1512716400, 
    1512720000, 1512723600, 1512727200, 1512730800, 1512734400, 1512738000, 
    1512741600, 1512745200, 1512748800, 1512752400, 1512756000, 1512759600, 
    1512763200, 1512766800, 1512770400, 1512774000, 1512777600, 1512781200, 
    1512784800, 1512788400, 1512792000, 1512795600, 1512799200, 1512802800, 
    1512806400, 1512810000, 1512813600, 1512817200, 1512820800, 1512824400, 
    1512828000, 1512831600, 1512835200, 1512838800, 1512842400, 1512846000, 
    1512849600, 1512853200, 1512856800, 1512860400, 1512864000, 1512867600, 
    1512871200, 1512874800, 1512878400, 1512882000, 1512885600, 1512889200, 
    1512892800, 1512896400, 1512900000, 1512903600, 1512907200, 1512910800, 
    1512914400, 1512918000, 1512921600, 1512925200, 1512928800, 1512932400, 
    1512936000, 1512939600, 1512943200, 1512946800, 1512950400, 1512954000, 
    1512957600, 1512961200, 1512964800, 1512968400, 1512972000, 1512975600, 
    1512979200, 1512982800, 1512986400, 1512990000, 1512993600, 1512997200, 
    1513000800, 1513004400, 1513008000, 1513011600, 1513015200, 1513018800, 
    1513022400, 1513026000, 1513029600, 1513033200, 1513036800, 1513040400, 
    1513044000, 1513047600, 1513051200, 1513054800, 1513058400, 1513062000, 
    1513065600, 1513069200, 1513072800, 1513076400, 1513080000, 1513083600, 
    1513087200, 1513090800, 1513094400, 1513098000, 1513101600, 1513105200, 
    1513108800, 1513112400, 1513116000, 1513119600, 1513123200, 1513126800, 
    1513130400, 1513134000, 1513137600, 1513141200, 1513144800, 1513148400, 
    1513152000, 1513155600, 1513159200, 1513162800, 1513166400, 1513170000, 
    1513173600, 1513177200, 1513180800, 1513184400, 1513188000, 1513191600, 
    1513195200, 1513198800, 1513202400, 1513206000, 1513209600, 1513213200, 
    1513216800, 1513220400, 1513224000, 1513227600, 1513231200, 1513234800, 
    1513238400, 1513242000, 1513245600, 1513249200, 1513252800, 1513256400, 
    1513260000, 1513263600, 1513267200, 1513270800, 1513274400, 1513278000, 
    1513281600, 1513285200, 1513288800, 1513292400, 1513296000, 1513299600, 
    1513303200, 1513306800, 1513310400, 1513314000, 1513317600, 1513321200, 
    1513324800, 1513328400, 1513332000, 1513335600, 1513339200, 1513342800, 
    1513346400, 1513350000, 1513353600, 1513357200, 1513360800, 1513364400, 
    1513368000, 1513371600, 1513375200, 1513378800, 1513382400, 1513386000, 
    1513389600, 1513393200, 1513396800, 1513400400, 1513404000, 1513407600, 
    1513411200, 1513414800, 1513418400, 1513422000, 1513425600, 1513429200, 
    1513432800, 1513436400, 1513440000, 1513443600, 1513447200, 1513450800, 
    1513454400, 1513458000, 1513461600, 1513465200, 1513468800, 1513472400, 
    1513476000, 1513479600, 1513483200, 1513486800, 1513490400, 1513494000, 
    1513497600, 1513501200, 1513504800, 1513508400, 1513512000, 1513515600, 
    1513519200, 1513522800, 1513526400, 1513530000, 1513533600, 1513537200, 
    1513540800, 1513544400, 1513548000, 1513551600, 1513555200, 1513558800, 
    1513562400, 1513566000, 1513569600, 1513573200, 1513576800, 1513580400, 
    1513584000, 1513587600, 1513591200, 1513594800, 1513598400, 1513602000, 
    1513605600, 1513609200, 1513612800, 1513616400, 1513620000, 1513623600, 
    1513627200, 1513630800, 1513634400, 1513638000, 1513641600, 1513645200, 
    1513648800, 1513652400, 1513656000, 1513659600, 1513663200, 1513666800, 
    1513670400, 1513674000, 1513677600, 1513681200, 1513684800, 1513688400, 
    1513692000, 1513695600, 1513699200, 1513702800, 1513706400, 1513710000, 
    1513713600, 1513717200, 1513720800, 1513724400, 1513728000, 1513731600, 
    1513735200, 1513738800, 1513742400, 1513746000, 1513749600, 1513753200, 
    1513756800, 1513760400, 1513764000, 1513767600, 1513771200, 1513774800, 
    1513778400, 1513782000, 1513785600, 1513789200, 1513792800, 1513796400, 
    1513800000, 1513803600, 1513807200, 1513810800, 1513814400, 1513818000, 
    1513821600, 1513825200, 1513828800, 1513832400, 1513836000, 1513839600, 
    1513843200, 1513846800, 1513850400, 1513854000, 1513857600, 1513861200, 
    1513864800, 1513868400, 1513872000, 1513875600, 1513879200, 1513882800, 
    1513886400, 1513890000, 1513893600, 1513897200, 1513900800, 1513904400, 
    1513908000, 1513911600, 1513915200, 1513918800, 1513922400, 1513926000, 
    1513929600, 1513933200, 1513936800, 1513940400, 1513944000, 1513947600, 
    1513951200, 1513954800, 1513958400, 1513962000, 1513965600, 1513969200, 
    1513972800, 1513976400, 1513980000, 1513983600, 1513987200, 1513990800, 
    1513994400, 1513998000, 1514001600, 1514005200, 1514008800, 1514012400, 
    1514016000, 1514019600, 1514023200, 1514026800, 1514030400, 1514034000, 
    1514037600, 1514041200, 1514044800, 1514048400, 1514052000, 1514055600, 
    1514059200, 1514062800, 1514066400, 1514070000, 1514073600, 1514077200, 
    1514080800, 1514084400, 1514088000, 1514091600, 1514095200, 1514098800, 
    1514102400, 1514106000, 1514109600, 1514113200, 1514116800, 1514120400, 
    1514124000, 1514127600, 1514131200, 1514134800, 1514138400, 1514142000, 
    1514145600, 1514149200, 1514152800, 1514156400, 1514160000, 1514163600, 
    1514167200, 1514170800, 1514174400, 1514178000, 1514181600, 1514185200, 
    1514188800, 1514192400, 1514196000, 1514199600, 1514203200, 1514206800, 
    1514210400, 1514214000, 1514217600, 1514221200, 1514224800, 1514228400, 
    1514232000, 1514235600, 1514239200, 1514242800, 1514246400, 1514250000, 
    1514253600, 1514257200, 1514260800, 1514264400, 1514268000, 1514271600, 
    1514275200, 1514278800, 1514282400, 1514286000, 1514289600, 1514293200, 
    1514296800, 1514300400, 1514304000, 1514307600, 1514311200, 1514314800, 
    1514318400, 1514322000, 1514325600, 1514329200, 1514332800, 1514336400, 
    1514340000, 1514343600, 1514347200, 1514350800, 1514354400, 1514358000, 
    1514361600, 1514365200, 1514368800, 1514372400, 1514376000, 1514379600, 
    1514383200, 1514386800, 1514390400, 1514394000, 1514397600, 1514401200, 
    1514404800, 1514408400, 1514412000, 1514415600, 1514419200, 1514422800, 
    1514426400, 1514430000, 1514433600, 1514437200, 1514440800, 1514444400, 
    1514448000, 1514451600, 1514455200, 1514458800, 1514462400, 1514466000, 
    1514469600, 1514473200, 1514476800, 1514480400, 1514484000, 1514487600, 
    1514491200, 1514494800, 1514498400, 1514502000, 1514505600, 1514509200, 
    1514512800, 1514516400, 1514520000, 1514523600, 1514527200, 1514530800, 
    1514534400, 1514538000, 1514541600, 1514545200, 1514548800, 1514552400, 
    1514556000, 1514559600, 1514563200, 1514566800, 1514570400, 1514574000, 
    1514577600, 1514581200, 1514584800, 1514588400, 1514592000, 1514595600, 
    1514599200, 1514602800, 1514606400, 1514610000, 1514613600, 1514617200, 
    1514620800, 1514624400, 1514628000, 1514631600, 1514635200, 1514638800, 
    1514642400, 1514646000, 1514649600, 1514653200, 1514656800, 1514660400, 
    1514664000, 1514667600, 1514671200, 1514674800, 1514678400, 1514682000, 
    1514685600, 1514689200, 1514692800, 1514696400, 1514700000, 1514703600, 
    1514707200, 1514710800, 1514714400, 1514718000, 1514721600, 1514725200, 
    1514728800, 1514732400, 1514736000, 1514739600, 1514743200, 1514746800, 
    1514750400, 1514754000, 1514757600, 1514761200, 1514764800, 1514768400, 
    1514772000, 1514775600, 1514779200, 1514782800, 1514786400, 1514790000, 
    1514793600, 1514797200, 1514800800, 1514804400, 1514808000, 1514811600, 
    1514815200, 1514818800, 1514822400, 1514826000, 1514829600, 1514833200, 
    1514836800, 1514840400, 1514844000, 1514847600, 1514851200, 1514854800, 
    1514858400, 1514862000, 1514865600, 1514869200, 1514872800, 1514876400, 
    1514880000, 1514883600, 1514887200, 1514890800, 1514894400, 1514898000, 
    1514901600, 1514905200, 1514908800, 1514912400, 1514916000, 1514919600, 
    1514923200, 1514926800, 1514930400, 1514934000, 1514937600, 1514941200, 
    1514944800, 1514948400, 1514952000, 1514955600, 1514959200, 1514962800, 
    1514966400, 1514970000, 1514973600, 1514977200, 1514980800, 1514984400, 
    1514988000, 1514991600, 1514995200, 1514998800, 1515002400, 1515006000, 
    1515009600, 1515013200, 1515016800, 1515020400, 1515024000, 1515027600, 
    1515031200, 1515034800, 1515038400, 1515042000, 1515045600, 1515049200, 
    1515052800, 1515056400, 1515060000, 1515063600, 1515067200, 1515070800, 
    1515074400, 1515078000, 1515081600, 1515085200, 1515088800, 1515092400, 
    1515096000, 1515099600, 1515103200, 1515106800, 1515110400, 1515114000, 
    1515117600, 1515121200, 1515124800, 1515128400, 1515132000, 1515135600, 
    1515139200, 1515142800, 1515146400, 1515150000, 1515153600, 1515157200, 
    1515160800, 1515164400, 1515168000, 1515171600, 1515175200, 1515178800, 
    1515182400, 1515186000, 1515189600, 1515193200, 1515196800, 1515200400, 
    1515204000, 1515207600, 1515211200, 1515214800, 1515218400, 1515222000, 
    1515225600, 1515229200, 1515232800, 1515236400, 1515240000, 1515243600, 
    1515247200, 1515250800, 1515254400, 1515258000, 1515261600, 1515265200, 
    1515268800, 1515272400, 1515276000, 1515279600, 1515283200, 1515286800, 
    1515290400, 1515294000, 1515297600, 1515301200, 1515304800, 1515308400, 
    1515312000, 1515315600, 1515319200, 1515322800, 1515326400, 1515330000, 
    1515333600, 1515337200, 1515340800, 1515344400, 1515348000, 1515351600, 
    1515355200, 1515358800, 1515362400, 1515366000, 1515369600, 1515373200, 
    1515376800, 1515380400, 1515384000, 1515387600, 1515391200, 1515394800, 
    1515398400, 1515402000, 1515405600, 1515409200, 1515412800, 1515416400, 
    1515420000, 1515423600, 1515427200, 1515430800, 1515434400, 1515438000, 
    1515441600, 1515445200, 1515448800, 1515452400, 1515456000, 1515459600, 
    1515463200, 1515466800, 1515470400, 1515474000, 1515477600, 1515481200, 
    1515484800, 1515488400, 1515492000, 1515495600, 1515499200, 1515502800, 
    1515506400, 1515510000, 1515513600, 1515517200, 1515520800, 1515524400, 
    1515528000, 1515531600, 1515535200, 1515538800, 1515542400, 1515546000, 
    1515549600, 1515553200, 1515556800, 1515560400, 1515564000, 1515567600, 
    1515571200, 1515574800, 1515578400, 1515582000, 1515585600, 1515589200, 
    1515592800, 1515596400, 1515600000, 1515603600, 1515607200, 1515610800, 
    1515614400, 1515618000, 1515621600, 1515625200, 1515628800, 1515632400, 
    1515636000, 1515639600, 1515643200, 1515646800, 1515650400, 1515654000, 
    1515657600, 1515661200, 1515664800, 1515668400, 1515672000, 1515675600, 
    1515679200, 1515682800, 1515686400, 1515690000, 1515693600, 1515697200, 
    1515700800, 1515704400, 1515708000, 1515711600, 1515715200, 1515718800, 
    1515722400, 1515726000, 1515729600, 1515733200, 1515736800, 1515740400, 
    1515744000, 1515747600, 1515751200, 1515754800, 1515758400, 1515762000, 
    1515765600, 1515769200, 1515772800, 1515776400, 1515780000, 1515783600, 
    1515787200, 1515790800, 1515794400, 1515798000, 1515801600, 1515805200, 
    1515808800, 1515812400, 1515816000, 1515819600, 1515823200, 1515826800, 
    1515830400, 1515834000, 1515837600, 1515841200, 1515844800, 1515848400, 
    1515852000, 1515855600, 1515859200, 1515862800, 1515866400, 1515870000, 
    1515873600, 1515877200, 1515880800, 1515884400, 1515888000, 1515891600, 
    1515895200, 1515898800, 1515902400, 1515906000, 1515909600, 1515913200, 
    1515916800, 1515920400, 1515924000, 1515927600, 1515931200, 1515934800, 
    1515938400, 1515942000, 1515945600, 1515949200, 1515952800, 1515956400, 
    1515960000, 1515963600, 1515967200, 1515970800, 1515974400, 1515978000, 
    1515981600, 1515985200, 1515988800, 1515992400, 1515996000, 1515999600, 
    1516003200, 1516006800, 1516010400, 1516014000, 1516017600, 1516021200, 
    1516024800, 1516028400, 1516032000, 1516035600, 1516039200, 1516042800, 
    1516046400, 1516050000, 1516053600, 1516057200, 1516060800, 1516064400, 
    1516068000, 1516071600, 1516075200, 1516078800, 1516082400, 1516086000, 
    1516089600, 1516093200, 1516096800, 1516100400, 1516104000, 1516107600, 
    1516111200, 1516114800, 1516118400, 1516122000, 1516125600, 1516129200, 
    1516132800, 1516136400, 1516140000, 1516143600, 1516147200, 1516150800, 
    1516154400, 1516158000, 1516161600, 1516165200, 1516168800, 1516172400, 
    1516176000, 1516179600, 1516183200, 1516186800, 1516190400, 1516194000, 
    1516197600, 1516201200, 1516204800, 1516208400, 1516212000, 1516215600, 
    1516219200, 1516222800, 1516226400, 1516230000, 1516233600, 1516237200, 
    1516240800, 1516244400, 1516248000, 1516251600, 1516255200, 1516258800, 
    1516262400, 1516266000, 1516269600, 1516273200, 1516276800, 1516280400, 
    1516284000, 1516287600, 1516291200, 1516294800, 1516298400, 1516302000, 
    1516305600, 1516309200, 1516312800, 1516316400, 1516320000, 1516323600, 
    1516327200, 1516330800, 1516334400, 1516338000, 1516341600, 1516345200, 
    1516348800, 1516352400, 1516356000, 1516359600, 1516363200, 1516366800, 
    1516370400, 1516374000, 1516377600, 1516381200, 1516384800, 1516388400, 
    1516392000, 1516395600, 1516399200, 1516402800, 1516406400, 1516410000, 
    1516413600, 1516417200, 1516420800, 1516424400, 1516428000, 1516431600, 
    1516435200, 1516438800, 1516442400, 1516446000, 1516449600, 1516453200, 
    1516456800, 1516460400, 1516464000, 1516467600, 1516471200, 1516474800, 
    1516478400, 1516482000, 1516485600, 1516489200, 1516492800, 1516496400, 
    1516500000, 1516503600, 1516507200, 1516510800, 1516514400, 1516518000, 
    1516521600, 1516525200, 1516528800, 1516532400, 1516536000, 1516539600, 
    1516543200, 1516546800, 1516550400, 1516554000, 1516557600, 1516561200, 
    1516564800, 1516568400, 1516572000, 1516575600, 1516579200, 1516582800, 
    1516586400, 1516590000, 1516593600, 1516597200, 1516600800, 1516604400, 
    1516608000, 1516611600, 1516615200, 1516618800, 1516622400, 1516626000, 
    1516629600, 1516633200, 1516636800, 1516640400, 1516644000, 1516647600, 
    1516651200, 1516654800, 1516658400, 1516662000, 1516665600, 1516669200, 
    1516672800, 1516676400, 1516680000, 1516683600, 1516687200, 1516690800, 
    1516694400, 1516698000, 1516701600, 1516705200, 1516708800, 1516712400, 
    1516716000, 1516719600, 1516723200, 1516726800, 1516730400, 1516734000, 
    1516737600, 1516741200, 1516744800, 1516748400, 1516752000, 1516755600, 
    1516759200, 1516762800, 1516766400, 1516770000, 1516773600, 1516777200, 
    1516780800, 1516784400, 1516788000, 1516791600, 1516795200, 1516798800, 
    1516802400, 1516806000, 1516809600, 1516813200, 1516816800, 1516820400, 
    1516824000, 1516827600, 1516831200, 1516834800, 1516838400, 1516842000, 
    1516845600, 1516849200, 1516852800, 1516856400, 1516860000, 1516863600, 
    1516867200, 1516870800, 1516874400, 1516878000, 1516881600, 1516885200, 
    1516888800, 1516892400, 1516896000, 1516899600, 1516903200, 1516906800, 
    1516910400, 1516914000, 1516917600, 1516921200, 1516924800, 1516928400, 
    1516932000, 1516935600, 1516939200, 1516942800, 1516946400, 1516950000, 
    1516953600, 1516957200, 1516960800, 1516964400, 1516968000, 1516971600, 
    1516975200, 1516978800, 1516982400, 1516986000, 1516989600, 1516993200, 
    1516996800, 1517000400, 1517004000, 1517007600, 1517011200, 1517014800, 
    1517018400, 1517022000, 1517025600, 1517029200, 1517032800, 1517036400, 
    1517040000, 1517043600, 1517047200, 1517050800, 1517054400, 1517058000, 
    1517061600, 1517065200, 1517068800, 1517072400, 1517076000, 1517079600, 
    1517083200, 1517086800, 1517090400, 1517094000, 1517097600, 1517101200, 
    1517104800, 1517108400, 1517112000, 1517115600, 1517119200, 1517122800, 
    1517126400, 1517130000, 1517133600, 1517137200, 1517140800, 1517144400, 
    1517148000, 1517151600, 1517155200, 1517158800, 1517162400, 1517166000, 
    1517169600, 1517173200, 1517176800, 1517180400, 1517184000, 1517187600, 
    1517191200, 1517194800, 1517198400, 1517202000, 1517205600, 1517209200, 
    1517212800, 1517216400, 1517220000, 1517223600, 1517227200, 1517230800, 
    1517234400, 1517238000, 1517241600, 1517245200, 1517248800, 1517252400, 
    1517256000, 1517259600, 1517263200, 1517266800, 1517270400, 1517274000, 
    1517277600, 1517281200, 1517284800, 1517288400, 1517292000, 1517295600, 
    1517299200, 1517302800, 1517306400, 1517310000, 1517313600, 1517317200, 
    1517320800, 1517324400, 1517328000, 1517331600, 1517335200, 1517338800, 
    1517342400, 1517346000, 1517349600, 1517353200, 1517356800, 1517360400, 
    1517364000, 1517367600, 1517371200, 1517374800, 1517378400, 1517382000, 
    1517385600, 1517389200, 1517392800, 1517396400, 1517400000, 1517403600, 
    1517407200, 1517410800, 1517414400, 1517418000, 1517421600, 1517425200, 
    1517428800, 1517432400, 1517436000, 1517439600, 1517443200, 1517446800, 
    1517450400, 1517454000, 1517457600, 1517461200, 1517464800, 1517468400, 
    1517472000, 1517475600, 1517479200, 1517482800, 1517486400, 1517490000, 
    1517493600, 1517497200, 1517500800, 1517504400, 1517508000, 1517511600, 
    1517515200, 1517518800, 1517522400, 1517526000, 1517529600, 1517533200, 
    1517536800, 1517540400, 1517544000, 1517547600, 1517551200, 1517554800, 
    1517558400, 1517562000, 1517565600, 1517569200, 1517572800, 1517576400, 
    1517580000, 1517583600, 1517587200, 1517590800, 1517594400, 1517598000, 
    1517601600, 1517605200, 1517608800, 1517612400, 1517616000, 1517619600, 
    1517623200, 1517626800, 1517630400, 1517634000, 1517637600, 1517641200, 
    1517644800, 1517648400, 1517652000, 1517655600, 1517659200, 1517662800, 
    1517666400, 1517670000, 1517673600, 1517677200, 1517680800, 1517684400, 
    1517688000, 1517691600, 1517695200, 1517698800, 1517702400, 1517706000, 
    1517709600, 1517713200, 1517716800, 1517720400, 1517724000, 1517727600, 
    1517731200, 1517734800, 1517738400, 1517742000, 1517745600, 1517749200, 
    1517752800, 1517756400, 1517760000, 1517763600, 1517767200, 1517770800, 
    1517774400, 1517778000, 1517781600, 1517785200, 1517788800, 1517792400, 
    1517796000, 1517799600, 1517803200, 1517806800, 1517810400, 1517814000, 
    1517817600, 1517821200, 1517824800, 1517828400, 1517832000, 1517835600, 
    1517839200, 1517842800, 1517846400, 1517850000, 1517853600, 1517857200, 
    1517860800, 1517864400, 1517868000, 1517871600, 1517875200, 1517878800, 
    1517882400, 1517886000, 1517889600, 1517893200, 1517896800, 1517900400, 
    1517904000, 1517907600, 1517911200, 1517914800, 1517918400, 1517922000, 
    1517925600, 1517929200, 1517932800, 1517936400, 1517940000, 1517943600, 
    1517947200, 1517950800, 1517954400, 1517958000, 1517961600, 1517965200, 
    1517968800, 1517972400, 1517976000, 1517979600, 1517983200, 1517986800, 
    1517990400, 1517994000, 1517997600, 1518001200, 1518004800, 1518008400, 
    1518012000, 1518015600, 1518019200, 1518022800, 1518026400, 1518030000, 
    1518033600, 1518037200, 1518040800, 1518044400, 1518048000, 1518051600, 
    1518055200, 1518058800, 1518062400, 1518066000, 1518069600, 1518073200, 
    1518076800, 1518080400, 1518084000, 1518087600, 1518091200, 1518094800, 
    1518098400, 1518102000, 1518105600, 1518109200, 1518112800, 1518116400, 
    1518120000, 1518123600, 1518127200, 1518130800, 1518134400, 1518138000, 
    1518141600, 1518145200, 1518148800, 1518152400, 1518156000, 1518159600, 
    1518163200, 1518166800, 1518170400, 1518174000, 1518177600, 1518181200, 
    1518184800, 1518188400, 1518192000, 1518195600, 1518199200, 1518202800, 
    1518206400, 1518210000, 1518213600, 1518217200, 1518220800, 1518224400, 
    1518228000, 1518231600, 1518235200, 1518238800, 1518242400, 1518246000, 
    1518249600, 1518253200, 1518256800, 1518260400, 1518264000, 1518267600, 
    1518271200, 1518274800, 1518278400, 1518282000, 1518285600, 1518289200, 
    1518292800, 1518296400, 1518300000, 1518303600, 1518307200, 1518310800, 
    1518314400, 1518318000, 1518321600, 1518325200, 1518328800, 1518332400, 
    1518336000, 1518339600, 1518343200, 1518346800, 1518350400, 1518354000, 
    1518357600, 1518361200, 1518364800, 1518368400, 1518372000, 1518375600, 
    1518379200, 1518382800, 1518386400, 1518390000, 1518393600, 1518397200, 
    1518400800, 1518404400, 1518408000, 1518411600, 1518415200, 1518418800, 
    1518422400, 1518426000, 1518429600, 1518433200, 1518436800, 1518440400, 
    1518444000, 1518447600, 1518451200, 1518454800, 1518458400, 1518462000, 
    1518465600, 1518469200, 1518472800, 1518476400, 1518480000, 1518483600, 
    1518487200, 1518490800, 1518494400, 1518498000, 1518501600, 1518505200, 
    1518508800, 1518512400, 1518516000, 1518519600, 1518523200, 1518526800, 
    1518530400, 1518534000, 1518537600, 1518541200, 1518544800, 1518548400, 
    1518552000, 1518555600, 1518559200, 1518562800, 1518566400, 1518570000, 
    1518573600, 1518577200, 1518580800, 1518584400, 1518588000, 1518591600, 
    1518595200, 1518598800, 1518602400, 1518606000, 1518609600, 1518613200, 
    1518616800, 1518620400, 1518624000, 1518627600, 1518631200, 1518634800, 
    1518638400, 1518642000, 1518645600, 1518649200, 1518652800, 1518656400, 
    1518660000, 1518663600, 1518667200, 1518670800, 1518674400, 1518678000, 
    1518681600, 1518685200, 1518688800, 1518692400, 1518696000, 1518699600, 
    1518703200, 1518706800, 1518710400, 1518714000, 1518717600, 1518721200, 
    1518724800, 1518728400, 1518732000, 1518735600, 1518739200, 1518742800, 
    1518746400, 1518750000, 1518753600, 1518757200, 1518760800, 1518764400, 
    1518768000, 1518771600, 1518775200, 1518778800, 1518782400, 1518786000, 
    1518789600, 1518793200, 1518796800, 1518800400, 1518804000, 1518807600, 
    1518811200, 1518814800, 1518818400, 1518822000, 1518825600, 1518829200, 
    1518832800, 1518836400, 1518840000, 1518843600, 1518847200, 1518850800, 
    1518854400, 1518858000, 1518861600, 1518865200, 1518868800, 1518872400, 
    1518876000, 1518879600, 1518883200, 1518886800, 1518890400, 1518894000, 
    1518897600, 1518901200, 1518904800, 1518908400, 1518912000, 1518915600, 
    1518919200, 1518922800, 1518926400, 1518930000, 1518933600, 1518937200, 
    1518940800, 1518944400, 1518948000, 1518951600, 1518955200, 1518958800, 
    1518962400, 1518966000, 1518969600, 1518973200, 1518976800, 1518980400, 
    1518984000, 1518987600, 1518991200, 1518994800, 1518998400, 1519002000, 
    1519005600, 1519009200, 1519012800, 1519016400, 1519020000, 1519023600, 
    1519027200, 1519030800, 1519034400, 1519038000, 1519041600, 1519045200, 
    1519048800, 1519052400, 1519056000, 1519059600, 1519063200, 1519066800, 
    1519070400, 1519074000, 1519077600, 1519081200, 1519084800, 1519088400, 
    1519092000, 1519095600, 1519099200, 1519102800, 1519106400, 1519110000, 
    1519113600, 1519117200, 1519120800, 1519124400, 1519128000, 1519131600, 
    1519135200, 1519138800, 1519142400, 1519146000, 1519149600, 1519153200, 
    1519156800, 1519160400, 1519164000, 1519167600, 1519171200, 1519174800, 
    1519178400, 1519182000, 1519185600, 1519189200, 1519192800, 1519196400, 
    1519200000, 1519203600, 1519207200, 1519210800, 1519214400, 1519218000, 
    1519221600, 1519225200, 1519228800, 1519232400, 1519236000, 1519239600, 
    1519243200, 1519246800, 1519250400, 1519254000, 1519257600, 1519261200, 
    1519264800, 1519268400, 1519272000, 1519275600, 1519279200, 1519282800, 
    1519286400, 1519290000, 1519293600, 1519297200, 1519300800, 1519304400, 
    1519308000, 1519311600, 1519315200, 1519318800, 1519322400, 1519326000, 
    1519329600, 1519333200, 1519336800, 1519340400, 1519344000, 1519347600, 
    1519351200, 1519354800, 1519358400, 1519362000, 1519365600, 1519369200, 
    1519372800, 1519376400, 1519380000, 1519383600, 1519387200, 1519390800, 
    1519394400, 1519398000, 1519401600, 1519405200, 1519408800, 1519412400, 
    1519416000, 1519419600, 1519423200, 1519426800, 1519430400, 1519434000, 
    1519437600, 1519441200, 1519444800, 1519448400, 1519452000, 1519455600, 
    1519459200, 1519462800, 1519466400, 1519470000, 1519473600, 1519477200, 
    1519480800, 1519484400, 1519488000, 1519491600, 1519495200, 1519498800, 
    1519502400, 1519506000, 1519509600, 1519513200, 1519516800, 1519520400, 
    1519524000, 1519527600, 1519531200, 1519534800, 1519538400, 1519542000, 
    1519545600, 1519549200, 1519552800, 1519556400, 1519560000, 1519563600, 
    1519567200, 1519570800, 1519574400, 1519578000, 1519581600, 1519585200, 
    1519588800, 1519592400, 1519596000, 1519599600, 1519603200, 1519606800, 
    1519610400, 1519614000, 1519617600, 1519621200, 1519624800, 1519628400, 
    1519632000, 1519635600, 1519639200, 1519642800, 1519646400, 1519650000, 
    1519653600, 1519657200, 1519660800, 1519664400, 1519668000, 1519671600, 
    1519675200, 1519678800, 1519682400, 1519686000, 1519689600, 1519693200, 
    1519696800, 1519700400, 1519704000, 1519707600, 1519711200, 1519714800, 
    1519718400, 1519722000, 1519725600, 1519729200, 1519732800, 1519736400, 
    1519740000, 1519743600, 1519747200, 1519750800, 1519754400, 1519758000, 
    1519761600, 1519765200, 1519768800, 1519772400, 1519776000, 1519779600, 
    1519783200, 1519786800, 1519790400, 1519794000, 1519797600, 1519801200, 
    1519804800, 1519808400, 1519812000, 1519815600, 1519819200, 1519822800, 
    1519826400, 1519830000, 1519833600, 1519837200, 1519840800, 1519844400, 
    1519848000, 1519851600, 1519855200, 1519858800, 1519862400, 1519866000, 
    1519869600, 1519873200, 1519876800, 1519880400, 1519884000, 1519887600, 
    1519891200, 1519894800, 1519898400, 1519902000, 1519905600, 1519909200, 
    1519912800, 1519916400, 1519920000, 1519923600, 1519927200, 1519930800, 
    1519934400, 1519938000, 1519941600, 1519945200, 1519948800, 1519952400, 
    1519956000, 1519959600, 1519963200, 1519966800, 1519970400, 1519974000, 
    1519977600, 1519981200, 1519984800, 1519988400, 1519992000, 1519995600, 
    1519999200, 1520002800, 1520006400, 1520010000, 1520013600, 1520017200, 
    1520020800, 1520024400, 1520028000, 1520031600, 1520035200, 1520038800, 
    1520042400, 1520046000, 1520049600, 1520053200, 1520056800, 1520060400, 
    1520064000, 1520067600, 1520071200, 1520074800, 1520078400, 1520082000, 
    1520085600, 1520089200, 1520092800, 1520096400, 1520100000, 1520103600, 
    1520107200, 1520110800, 1520114400, 1520118000, 1520121600, 1520125200, 
    1520128800, 1520132400, 1520136000, 1520139600, 1520143200, 1520146800, 
    1520150400, 1520154000, 1520157600, 1520161200, 1520164800, 1520168400, 
    1520172000, 1520175600, 1520179200, 1520182800, 1520186400, 1520190000, 
    1520193600, 1520197200, 1520200800, 1520204400, 1520208000, 1520211600, 
    1520215200, 1520218800, 1520222400, 1520226000, 1520229600, 1520233200, 
    1520236800, 1520240400, 1520244000, 1520247600, 1520251200, 1520254800, 
    1520258400, 1520262000, 1520265600, 1520269200, 1520272800, 1520276400, 
    1520280000, 1520283600, 1520287200, 1520290800, 1520294400, 1520298000, 
    1520301600, 1520305200, 1520308800, 1520312400, 1520316000, 1520319600, 
    1520323200, 1520326800, 1520330400, 1520334000, 1520337600, 1520341200, 
    1520344800, 1520348400, 1520352000, 1520355600, 1520359200, 1520362800, 
    1520366400, 1520370000, 1520373600, 1520377200, 1520380800, 1520384400, 
    1520388000, 1520391600, 1520395200, 1520398800, 1520402400, 1520406000, 
    1520409600, 1520413200, 1520416800, 1520420400, 1520424000, 1520427600, 
    1520431200, 1520434800, 1520438400, 1520442000, 1520445600, 1520449200, 
    1520452800, 1520456400, 1520460000, 1520463600, 1520467200, 1520470800, 
    1520474400, 1520478000, 1520481600, 1520485200, 1520488800, 1520492400, 
    1520496000, 1520499600, 1520503200, 1520506800, 1520510400, 1520514000, 
    1520517600, 1520521200, 1520524800, 1520528400, 1520532000, 1520535600, 
    1520539200, 1520542800, 1520546400, 1520550000, 1520553600, 1520557200, 
    1520560800, 1520564400, 1520568000, 1520571600, 1520575200, 1520578800, 
    1520582400, 1520586000, 1520589600, 1520593200, 1520596800, 1520600400, 
    1520604000, 1520607600, 1520611200, 1520614800, 1520618400, 1520622000, 
    1520625600, 1520629200, 1520632800, 1520636400, 1520640000, 1520643600, 
    1520647200, 1520650800, 1520654400, 1520658000, 1520661600, 1520665200, 
    1520668800, 1520672400, 1520676000, 1520679600, 1520683200, 1520686800, 
    1520690400, 1520694000, 1520697600, 1520701200, 1520704800, 1520708400, 
    1520712000, 1520715600, 1520719200, 1520722800, 1520726400, 1520730000, 
    1520733600, 1520737200, 1520740800, 1520744400, 1520748000, 1520751600, 
    1520755200, 1520758800, 1520762400, 1520766000, 1520769600, 1520773200, 
    1520776800, 1520780400, 1520784000, 1520787600, 1520791200, 1520794800, 
    1520798400, 1520802000, 1520805600, 1520809200, 1520812800, 1520816400, 
    1520820000, 1520823600, 1520827200, 1520830800, 1520834400, 1520838000, 
    1520841600, 1520845200, 1520848800, 1520852400, 1520856000, 1520859600, 
    1520863200, 1520866800, 1520870400, 1520874000, 1520877600, 1520881200, 
    1520884800, 1520888400, 1520892000, 1520895600, 1520899200, 1520902800, 
    1520906400, 1520910000, 1520913600, 1520917200, 1520920800, 1520924400, 
    1520928000, 1520931600, 1520935200, 1520938800, 1520942400, 1520946000, 
    1520949600, 1520953200, 1520956800, 1520960400, 1520964000, 1520967600, 
    1520971200, 1520974800, 1520978400, 1520982000, 1520985600, 1520989200, 
    1520992800, 1520996400, 1521000000, 1521003600, 1521007200, 1521010800, 
    1521014400, 1521018000, 1521021600, 1521025200, 1521028800, 1521032400, 
    1521036000, 1521039600, 1521043200, 1521046800, 1521050400, 1521054000, 
    1521057600, 1521061200, 1521064800, 1521068400, 1521072000, 1521075600, 
    1521079200, 1521082800, 1521086400, 1521090000, 1521093600, 1521097200, 
    1521100800, 1521104400, 1521108000, 1521111600, 1521115200, 1521118800, 
    1521122400, 1521126000, 1521129600, 1521133200, 1521136800, 1521140400, 
    1521144000, 1521147600, 1521151200, 1521154800, 1521158400, 1521162000, 
    1521165600, 1521169200, 1521172800, 1521176400, 1521180000, 1521183600, 
    1521187200, 1521190800, 1521194400, 1521198000, 1521201600, 1521205200, 
    1521208800, 1521212400, 1521216000, 1521219600, 1521223200, 1521226800, 
    1521230400, 1521234000, 1521237600, 1521241200, 1521244800, 1521248400, 
    1521252000, 1521255600, 1521259200, 1521262800, 1521266400, 1521270000, 
    1521273600, 1521277200, 1521280800, 1521284400, 1521288000, 1521291600, 
    1521295200, 1521298800, 1521302400, 1521306000, 1521309600, 1521313200, 
    1521316800, 1521320400, 1521324000, 1521327600, 1521331200, 1521334800, 
    1521338400, 1521342000, 1521345600, 1521349200, 1521352800, 1521356400, 
    1521360000, 1521363600, 1521367200, 1521370800, 1521374400, 1521378000, 
    1521381600, 1521385200, 1521388800, 1521392400, 1521396000, 1521399600, 
    1521403200, 1521406800, 1521410400, 1521414000, 1521417600, 1521421200, 
    1521424800, 1521428400, 1521432000, 1521435600, 1521439200, 1521442800, 
    1521446400, 1521450000, 1521453600, 1521457200, 1521460800, 1521464400, 
    1521468000, 1521471600, 1521475200, 1521478800, 1521482400, 1521486000, 
    1521489600, 1521493200, 1521496800, 1521500400, 1521504000, 1521507600, 
    1521511200, 1521514800, 1521518400, 1521522000, 1521525600, 1521529200, 
    1521532800, 1521536400, 1521540000, 1521543600, 1521547200, 1521550800, 
    1521554400, 1521558000, 1521561600, 1521565200, 1521568800, 1521572400, 
    1521576000, 1521579600, 1521583200, 1521586800, 1521590400, 1521594000, 
    1521597600, 1521601200, 1521604800, 1521608400, 1521612000, 1521615600, 
    1521619200, 1521622800, 1521626400, 1521630000, 1521633600, 1521637200, 
    1521640800, 1521644400, 1521648000, 1521651600, 1521655200, 1521658800, 
    1521662400, 1521666000, 1521669600, 1521673200, 1521676800, 1521680400, 
    1521684000, 1521687600, 1521691200, 1521694800, 1521698400, 1521702000, 
    1521705600, 1521709200, 1521712800, 1521716400, 1521720000, 1521723600, 
    1521727200, 1521730800, 1521734400, 1521738000, 1521741600, 1521745200, 
    1521748800, 1521752400, 1521756000, 1521759600, 1521763200, 1521766800, 
    1521770400, 1521774000, 1521777600, 1521781200, 1521784800, 1521788400, 
    1521792000, 1521795600, 1521799200, 1521802800, 1521806400, 1521810000, 
    1521813600, 1521817200, 1521820800, 1521824400, 1521828000, 1521831600, 
    1521835200, 1521838800, 1521842400, 1521846000, 1521849600, 1521853200, 
    1521856800, 1521860400, 1521864000, 1521867600, 1521871200, 1521874800, 
    1521878400, 1521882000, 1521885600, 1521889200, 1521892800, 1521896400, 
    1521900000, 1521903600, 1521907200, 1521910800, 1521914400, 1521918000, 
    1521921600, 1521925200, 1521928800, 1521932400, 1521936000, 1521939600, 
    1521943200, 1521946800, 1521950400, 1521954000, 1521957600, 1521961200, 
    1521964800, 1521968400, 1521972000, 1521975600, 1521979200, 1521982800, 
    1521986400, 1521990000, 1521993600, 1521997200, 1522000800, 1522004400, 
    1522008000, 1522011600, 1522015200, 1522018800, 1522022400, 1522026000, 
    1522029600, 1522033200, 1522036800, 1522040400, 1522044000, 1522047600, 
    1522051200, 1522054800, 1522058400, 1522062000, 1522065600, 1522069200, 
    1522072800, 1522076400, 1522080000, 1522083600, 1522087200, 1522090800, 
    1522094400, 1522098000, 1522101600, 1522105200, 1522108800, 1522112400, 
    1522116000, 1522119600, 1522123200, 1522126800, 1522130400, 1522134000, 
    1522137600, 1522141200, 1522144800, 1522148400, 1522152000, 1522155600, 
    1522159200, 1522162800, 1522166400, 1522170000, 1522173600, 1522177200, 
    1522180800, 1522184400, 1522188000, 1522191600, 1522195200, 1522198800, 
    1522202400, 1522206000, 1522209600, 1522213200, 1522216800, 1522220400, 
    1522224000, 1522227600, 1522231200, 1522234800, 1522238400, 1522242000, 
    1522245600, 1522249200, 1522252800, 1522256400, 1522260000, 1522263600, 
    1522267200, 1522270800, 1522274400, 1522278000, 1522281600, 1522285200, 
    1522288800, 1522292400, 1522296000, 1522299600, 1522303200, 1522306800, 
    1522310400, 1522314000, 1522317600, 1522321200, 1522324800, 1522328400, 
    1522332000, 1522335600, 1522339200, 1522342800, 1522346400, 1522350000, 
    1522353600, 1522357200, 1522360800, 1522364400, 1522368000, 1522371600, 
    1522375200, 1522378800, 1522382400, 1522386000, 1522389600, 1522393200, 
    1522396800, 1522400400, 1522404000, 1522407600, 1522411200, 1522414800, 
    1522418400, 1522422000, 1522425600, 1522429200, 1522432800, 1522436400, 
    1522440000, 1522443600, 1522447200, 1522450800, 1522454400, 1522458000, 
    1522461600, 1522465200, 1522468800, 1522472400, 1522476000, 1522479600, 
    1522483200, 1522486800, 1522490400, 1522494000, 1522497600, 1522501200, 
    1522504800, 1522508400, 1522512000, 1522515600, 1522519200, 1522522800, 
    1522526400, 1522530000, 1522533600, 1522537200, 1522540800, 1522544400, 
    1522548000, 1522551600, 1522555200, 1522558800, 1522562400, 1522566000, 
    1522569600, 1522573200, 1522576800, 1522580400, 1522584000, 1522587600, 
    1522591200, 1522594800, 1522598400, 1522602000, 1522605600, 1522609200, 
    1522612800, 1522616400, 1522620000, 1522623600, 1522627200, 1522630800, 
    1522634400, 1522638000, 1522641600, 1522645200, 1522648800, 1522652400, 
    1522656000, 1522659600, 1522663200, 1522666800, 1522670400, 1522674000, 
    1522677600, 1522681200, 1522684800, 1522688400, 1522692000, 1522695600, 
    1522699200, 1522702800, 1522706400, 1522710000, 1522713600, 1522717200, 
    1522720800, 1522724400, 1522728000, 1522731600, 1522735200, 1522738800, 
    1522742400, 1522746000, 1522749600, 1522753200, 1522756800, 1522760400, 
    1522764000, 1522767600, 1522771200, 1522774800, 1522778400, 1522782000, 
    1522785600, 1522789200, 1522792800, 1522796400, 1522800000, 1522803600, 
    1522807200, 1522810800, 1522814400, 1522818000, 1522821600, 1522825200, 
    1522828800, 1522832400, 1522836000, 1522839600, 1522843200, 1522846800, 
    1522850400, 1522854000, 1522857600, 1522861200, 1522864800, 1522868400, 
    1522872000, 1522875600, 1522879200, 1522882800, 1522886400, 1522890000, 
    1522893600, 1522897200, 1522900800, 1522904400, 1522908000, 1522911600, 
    1522915200, 1522918800, 1522922400, 1522926000, 1522929600, 1522933200, 
    1522936800, 1522940400, 1522944000, 1522947600, 1522951200, 1522954800, 
    1522958400, 1522962000, 1522965600, 1522969200, 1522972800, 1522976400, 
    1522980000, 1522983600, 1522987200, 1522990800, 1522994400, 1522998000, 
    1523001600, 1523005200, 1523008800, 1523012400, 1523016000, 1523019600, 
    1523023200, 1523026800, 1523030400, 1523034000, 1523037600, 1523041200, 
    1523044800, 1523048400, 1523052000, 1523055600, 1523059200, 1523062800, 
    1523066400, 1523070000, 1523073600, 1523077200, 1523080800, 1523084400, 
    1523088000, 1523091600, 1523095200, 1523098800, 1523102400, 1523106000, 
    1523109600, 1523113200, 1523116800, 1523120400, 1523124000, 1523127600, 
    1523131200, 1523134800, 1523138400, 1523142000, 1523145600, 1523149200, 
    1523152800, 1523156400, 1523160000, 1523163600, 1523167200, 1523170800, 
    1523174400, 1523178000, 1523181600, 1523185200, 1523188800, 1523192400, 
    1523196000, 1523199600, 1523203200, 1523206800, 1523210400, 1523214000, 
    1523217600, 1523221200, 1523224800, 1523228400, 1523232000, 1523235600, 
    1523239200, 1523242800, 1523246400, 1523250000, 1523253600, 1523257200, 
    1523260800, 1523264400, 1523268000, 1523271600, 1523275200, 1523278800, 
    1523282400, 1523286000, 1523289600, 1523293200, 1523296800, 1523300400, 
    1523304000, 1523307600, 1523311200, 1523314800, 1523318400, 1523322000, 
    1523325600, 1523329200, 1523332800, 1523336400, 1523340000, 1523343600, 
    1523347200, 1523350800, 1523354400, 1523358000, 1523361600, 1523365200, 
    1523368800, 1523372400, 1523376000, 1523379600, 1523383200, 1523386800, 
    1523390400, 1523394000, 1523397600, 1523401200, 1523404800, 1523408400, 
    1523412000, 1523415600, 1523419200, 1523422800, 1523426400, 1523430000, 
    1523433600, 1523437200, 1523440800, 1523444400, 1523448000, 1523451600, 
    1523455200, 1523458800, 1523462400, 1523466000, 1523469600, 1523473200, 
    1523476800, 1523480400, 1523484000, 1523487600, 1523491200, 1523494800, 
    1523498400, 1523502000, 1523505600, 1523509200, 1523512800, 1523516400, 
    1523520000, 1523523600, 1523527200, 1523530800, 1523534400, 1523538000, 
    1523541600, 1523545200, 1523548800, 1523552400, 1523556000, 1523559600, 
    1523563200, 1523566800, 1523570400, 1523574000, 1523577600, 1523581200, 
    1523584800, 1523588400, 1523592000, 1523595600, 1523599200, 1523602800, 
    1523606400, 1523610000, 1523613600, 1523617200, 1523620800, 1523624400, 
    1523628000, 1523631600, 1523635200, 1523638800, 1523642400, 1523646000, 
    1523649600, 1523653200, 1523656800, 1523660400, 1523664000, 1523667600, 
    1523671200, 1523674800, 1523678400, 1523682000, 1523685600, 1523689200, 
    1523692800, 1523696400, 1523700000, 1523703600, 1523707200, 1523710800, 
    1523714400, 1523718000, 1523721600, 1523725200, 1523728800, 1523732400, 
    1523736000, 1523739600, 1523743200, 1523746800, 1523750400, 1523754000, 
    1523757600, 1523761200, 1523764800, 1523768400, 1523772000, 1523775600, 
    1523779200, 1523782800, 1523786400, 1523790000, 1523793600, 1523797200, 
    1523800800, 1523804400, 1523808000, 1523811600, 1523815200, 1523818800, 
    1523822400, 1523826000, 1523829600, 1523833200, 1523836800, 1523840400, 
    1523844000, 1523847600, 1523851200, 1523854800, 1523858400, 1523862000, 
    1523865600, 1523869200, 1523872800, 1523876400, 1523880000, 1523883600, 
    1523887200, 1523890800, 1523894400, 1523898000, 1523901600, 1523905200, 
    1523908800, 1523912400, 1523916000, 1523919600, 1523923200, 1523926800, 
    1523930400, 1523934000, 1523937600, 1523941200, 1523944800, 1523948400, 
    1523952000, 1523955600, 1523959200, 1523962800, 1523966400, 1523970000, 
    1523973600, 1523977200, 1523980800, 1523984400, 1523988000, 1523991600, 
    1523995200, 1523998800, 1524002400, 1524006000, 1524009600, 1524013200, 
    1524016800, 1524020400, 1524024000, 1524027600, 1524031200, 1524034800, 
    1524038400, 1524042000, 1524045600, 1524049200, 1524052800, 1524056400, 
    1524060000, 1524063600, 1524067200, 1524070800, 1524074400, 1524078000, 
    1524081600, 1524085200, 1524088800, 1524092400, 1524096000, 1524099600, 
    1524103200, 1524106800, 1524110400, 1524114000, 1524117600, 1524121200, 
    1524124800, 1524128400, 1524132000, 1524135600, 1524139200, 1524142800, 
    1524146400, 1524150000, 1524153600, 1524157200, 1524160800, 1524164400, 
    1524168000, 1524171600, 1524175200, 1524178800, 1524182400, 1524186000, 
    1524189600, 1524193200, 1524196800, 1524200400, 1524204000, 1524207600, 
    1524211200, 1524214800, 1524218400, 1524222000, 1524225600, 1524229200, 
    1524232800, 1524236400, 1524240000, 1524243600, 1524247200, 1524250800, 
    1524254400, 1524258000, 1524261600, 1524265200, 1524268800, 1524272400, 
    1524276000, 1524279600, 1524283200, 1524286800, 1524290400, 1524294000, 
    1524297600, 1524301200, 1524304800, 1524308400, 1524312000, 1524315600, 
    1524319200, 1524322800, 1524326400, 1524330000, 1524333600, 1524337200, 
    1524340800, 1524344400, 1524348000, 1524351600, 1524355200, 1524358800, 
    1524362400, 1524366000, 1524369600, 1524373200, 1524376800, 1524380400, 
    1524384000, 1524387600, 1524391200, 1524394800, 1524398400, 1524402000, 
    1524405600, 1524409200, 1524412800, 1524416400, 1524420000, 1524423600, 
    1524427200, 1524430800, 1524434400, 1524438000, 1524441600, 1524445200, 
    1524448800, 1524452400, 1524456000, 1524459600, 1524463200, 1524466800, 
    1524470400, 1524474000, 1524477600, 1524481200, 1524484800, 1524488400, 
    1524492000, 1524495600, 1524499200, 1524502800, 1524506400, 1524510000, 
    1524513600, 1524517200, 1524520800, 1524524400, 1524528000, 1524531600, 
    1524535200, 1524538800, 1524542400, 1524546000, 1524549600, 1524553200, 
    1524556800, 1524560400, 1524564000, 1524567600, 1524571200, 1524574800, 
    1524578400, 1524582000, 1524585600, 1524589200, 1524592800, 1524596400, 
    1524600000, 1524603600, 1524607200, 1524610800, 1524614400, 1524618000, 
    1524621600, 1524625200, 1524628800, 1524632400, 1524636000, 1524639600, 
    1524643200, 1524646800, 1524650400, 1524654000, 1524657600, 1524661200, 
    1524664800, 1524668400, 1524672000, 1524675600, 1524679200, 1524682800, 
    1524686400, 1524690000, 1524693600, 1524697200, 1524700800, 1524704400, 
    1524708000, 1524711600, 1524715200, 1524718800, 1524722400, 1524726000, 
    1524729600, 1524733200, 1524736800, 1524740400, 1524744000, 1524747600, 
    1524751200, 1524754800, 1524758400, 1524762000, 1524765600, 1524769200, 
    1524772800, 1524776400, 1524780000, 1524783600, 1524787200, 1524790800, 
    1524794400, 1524798000, 1524801600, 1524805200, 1524808800, 1524812400, 
    1524816000, 1524819600, 1524823200, 1524826800, 1524830400, 1524834000, 
    1524837600, 1524841200, 1524844800, 1524848400, 1524852000, 1524855600, 
    1524859200, 1524862800, 1524866400, 1524870000, 1524873600, 1524877200, 
    1524880800, 1524884400, 1524888000, 1524891600, 1524895200, 1524898800, 
    1524902400, 1524906000, 1524909600, 1524913200, 1524916800, 1524920400, 
    1524924000, 1524927600, 1524931200, 1524934800, 1524938400, 1524942000, 
    1524945600, 1524949200, 1524952800, 1524956400, 1524960000, 1524963600, 
    1524967200, 1524970800, 1524974400, 1524978000, 1524981600, 1524985200, 
    1524988800, 1524992400, 1524996000, 1524999600, 1525003200, 1525006800, 
    1525010400, 1525014000, 1525017600, 1525021200, 1525024800, 1525028400, 
    1525032000, 1525035600, 1525039200, 1525042800, 1525046400, 1525050000, 
    1525053600, 1525057200, 1525060800, 1525064400, 1525068000, 1525071600, 
    1525075200, 1525078800, 1525082400, 1525086000, 1525089600, 1525093200, 
    1525096800, 1525100400, 1525104000, 1525107600, 1525111200, 1525114800, 
    1525118400, 1525122000, 1525125600, 1525129200, 1525132800, 1525136400, 
    1525140000, 1525143600, 1525147200, 1525150800, 1525154400, 1525158000, 
    1525161600, 1525165200, 1525168800, 1525172400, 1525176000, 1525179600, 
    1525183200, 1525186800, 1525190400, 1525194000, 1525197600, 1525201200, 
    1525204800, 1525208400, 1525212000, 1525215600, 1525219200, 1525222800, 
    1525226400, 1525230000, 1525233600, 1525237200, 1525240800, 1525244400, 
    1525248000, 1525251600, 1525255200, 1525258800, 1525262400, 1525266000, 
    1525269600, 1525273200, 1525276800, 1525280400, 1525284000, 1525287600, 
    1525291200, 1525294800, 1525298400, 1525302000, 1525305600, 1525309200, 
    1525312800, 1525316400, 1525320000, 1525323600, 1525327200, 1525330800, 
    1525334400, 1525338000, 1525341600, 1525345200, 1525348800, 1525352400, 
    1525356000, 1525359600, 1525363200, 1525366800, 1525370400, 1525374000, 
    1525377600, 1525381200, 1525384800, 1525388400, 1525392000, 1525395600, 
    1525399200, 1525402800, 1525406400, 1525410000, 1525413600, 1525417200, 
    1525420800, 1525424400, 1525428000, 1525431600, 1525435200, 1525438800, 
    1525442400, 1525446000, 1525449600, 1525453200, 1525456800, 1525460400, 
    1525464000, 1525467600, 1525471200, 1525474800, 1525478400, 1525482000, 
    1525485600, 1525489200, 1525492800, 1525496400, 1525500000, 1525503600, 
    1525507200, 1525510800, 1525514400, 1525518000, 1525521600, 1525525200, 
    1525528800, 1525532400, 1525536000, 1525539600, 1525543200, 1525546800, 
    1525550400, 1525554000, 1525557600, 1525561200, 1525564800, 1525568400, 
    1525572000, 1525575600, 1525579200, 1525582800, 1525586400, 1525590000, 
    1525593600, 1525597200, 1525600800, 1525604400, 1525608000, 1525611600, 
    1525615200, 1525618800, 1525622400, 1525626000, 1525629600, 1525633200, 
    1525636800, 1525640400, 1525644000, 1525647600, 1525651200, 1525654800, 
    1525658400, 1525662000, 1525665600, 1525669200, 1525672800, 1525676400, 
    1525680000, 1525683600, 1525687200, 1525690800, 1525694400, 1525698000, 
    1525701600, 1525705200, 1525708800, 1525712400, 1525716000, 1525719600, 
    1525723200, 1525726800, 1525730400, 1525734000, 1525737600, 1525741200, 
    1525744800, 1525748400, 1525752000, 1525755600, 1525759200, 1525762800, 
    1525766400, 1525770000, 1525773600, 1525777200, 1525780800, 1525784400, 
    1525788000, 1525791600, 1525795200, 1525798800, 1525802400, 1525806000, 
    1525809600, 1525813200, 1525816800, 1525820400, 1525824000, 1525827600, 
    1525831200, 1525834800, 1525838400, 1525842000, 1525845600, 1525849200, 
    1525852800, 1525856400, 1525860000, 1525863600, 1525867200, 1525870800, 
    1525874400, 1525878000, 1525881600, 1525885200, 1525888800, 1525892400, 
    1525896000, 1525899600, 1525903200, 1525906800, 1525910400, 1525914000, 
    1525917600, 1525921200, 1525924800, 1525928400, 1525932000, 1525935600, 
    1525939200, 1525942800, 1525946400, 1525950000, 1525953600, 1525957200, 
    1525960800, 1525964400, 1525968000, 1525971600, 1525975200, 1525978800, 
    1525982400, 1525986000, 1525989600, 1525993200, 1525996800, 1526000400, 
    1526004000, 1526007600, 1526011200, 1526014800, 1526018400, 1526022000, 
    1526025600, 1526029200, 1526032800, 1526036400, 1526040000, 1526043600, 
    1526047200, 1526050800, 1526054400, 1526058000, 1526061600, 1526065200, 
    1526068800, 1526072400, 1526076000, 1526079600, 1526083200, 1526086800, 
    1526090400, 1526094000, 1526097600, 1526101200, 1526104800, 1526108400, 
    1526112000, 1526115600, 1526119200, 1526122800, 1526126400, 1526130000, 
    1526133600, 1526137200, 1526140800, 1526144400, 1526148000, 1526151600, 
    1526155200, 1526158800, 1526162400, 1526166000, 1526169600, 1526173200, 
    1526176800, 1526180400, 1526184000, 1526187600, 1526191200, 1526194800, 
    1526198400, 1526202000, 1526205600, 1526209200, 1526212800, 1526216400, 
    1526220000, 1526223600, 1526227200, 1526230800, 1526234400, 1526238000, 
    1526241600, 1526245200, 1526248800, 1526252400, 1526256000, 1526259600, 
    1526263200, 1526266800, 1526270400, 1526274000, 1526277600, 1526281200, 
    1526284800, 1526288400, 1526292000, 1526295600, 1526299200, 1526302800, 
    1526306400, 1526310000, 1526313600, 1526317200, 1526320800, 1526324400, 
    1526328000, 1526331600, 1526335200, 1526338800, 1526342400, 1526346000, 
    1526349600, 1526353200, 1526356800, 1526360400, 1526364000, 1526367600, 
    1526371200, 1526374800, 1526378400, 1526382000, 1526385600, 1526389200, 
    1526392800, 1526396400, 1526400000, 1526403600, 1526407200, 1526410800, 
    1526414400, 1526418000, 1526421600, 1526425200, 1526428800, 1526432400, 
    1526436000, 1526439600, 1526443200, 1526446800, 1526450400, 1526454000, 
    1526457600, 1526461200, 1526464800, 1526468400, 1526472000, 1526475600, 
    1526479200, 1526482800, 1526486400, 1526490000, 1526493600, 1526497200, 
    1526500800, 1526504400, 1526508000, 1526511600, 1526515200, 1526518800, 
    1526522400, 1526526000, 1526529600, 1526533200, 1526536800, 1526540400, 
    1526544000, 1526547600, 1526551200, 1526554800, 1526558400, 1526562000, 
    1526565600, 1526569200, 1526572800, 1526576400, 1526580000, 1526583600, 
    1526587200, 1526590800, 1526594400, 1526598000, 1526601600, 1526605200, 
    1526608800, 1526612400, 1526616000, 1526619600, 1526623200, 1526626800, 
    1526630400, 1526634000, 1526637600, 1526641200, 1526644800, 1526648400, 
    1526652000, 1526655600, 1526659200, 1526662800, 1526666400, 1526670000, 
    1526673600, 1526677200, 1526680800, 1526684400, 1526688000, 1526691600, 
    1526695200, 1526698800, 1526702400, 1526706000, 1526709600, 1526713200, 
    1526716800, 1526720400, 1526724000, 1526727600, 1526731200, 1526734800, 
    1526738400, 1526742000, 1526745600, 1526749200, 1526752800, 1526756400, 
    1526760000, 1526763600, 1526767200, 1526770800, 1526774400, 1526778000, 
    1526781600, 1526785200, 1526788800, 1526792400, 1526796000, 1526799600, 
    1526803200, 1526806800, 1526810400, 1526814000, 1526817600, 1526821200, 
    1526824800, 1526828400, 1526832000, 1526835600, 1526839200, 1526842800, 
    1526846400, 1526850000, 1526853600, 1526857200, 1526860800, 1526864400, 
    1526868000, 1526871600, 1526875200, 1526878800, 1526882400, 1526886000, 
    1526889600, 1526893200, 1526896800, 1526900400, 1526904000, 1526907600, 
    1526911200, 1526914800, 1526918400, 1526922000, 1526925600, 1526929200, 
    1526932800, 1526936400, 1526940000, 1526943600, 1526947200, 1526950800, 
    1526954400, 1526958000, 1526961600, 1526965200, 1526968800, 1526972400, 
    1526976000, 1526979600, 1526983200, 1526986800, 1526990400, 1526994000, 
    1526997600, 1527001200, 1527004800, 1527008400, 1527012000, 1527015600, 
    1527019200, 1527022800, 1527026400, 1527030000, 1527033600, 1527037200, 
    1527040800, 1527044400, 1527048000, 1527051600, 1527055200, 1527058800, 
    1527062400, 1527066000, 1527069600, 1527073200, 1527076800, 1527080400, 
    1527084000, 1527087600, 1527091200, 1527094800, 1527098400, 1527102000, 
    1527105600, 1527109200, 1527112800, 1527116400, 1527120000, 1527123600, 
    1527127200, 1527130800, 1527134400, 1527138000, 1527141600, 1527145200, 
    1527148800, 1527152400, 1527156000, 1527159600, 1527163200, 1527166800, 
    1527170400, 1527174000, 1527177600, 1527181200, 1527184800, 1527188400, 
    1527192000, 1527195600, 1527199200, 1527202800, 1527206400, 1527210000, 
    1527213600, 1527217200, 1527220800, 1527224400, 1527228000, 1527231600, 
    1527235200, 1527238800, 1527242400, 1527246000, 1527249600, 1527253200, 
    1527256800, 1527260400, 1527264000, 1527267600, 1527271200, 1527274800, 
    1527278400, 1527282000, 1527285600, 1527289200, 1527292800, 1527296400, 
    1527300000, 1527303600, 1527307200, 1527310800, 1527314400, 1527318000, 
    1527321600, 1527325200, 1527328800, 1527332400, 1527336000, 1527339600, 
    1527343200, 1527346800, 1527350400, 1527354000, 1527357600, 1527361200, 
    1527364800, 1527368400, 1527372000, 1527375600, 1527379200, 1527382800, 
    1527386400, 1527390000, 1527393600, 1527397200, 1527400800, 1527404400, 
    1527408000, 1527411600, 1527415200, 1527418800, 1527422400, 1527426000, 
    1527429600, 1527433200, 1527436800, 1527440400, 1527444000, 1527447600, 
    1527451200, 1527454800, 1527458400, 1527462000, 1527465600, 1527469200, 
    1527472800, 1527476400, 1527480000, 1527483600, 1527487200, 1527490800, 
    1527494400, 1527498000, 1527501600, 1527505200, 1527508800, 1527512400, 
    1527516000, 1527519600, 1527523200, 1527526800, 1527530400, 1527534000, 
    1527537600, 1527541200, 1527544800, 1527548400, 1527552000, 1527555600, 
    1527559200, 1527562800, 1527566400, 1527570000, 1527573600, 1527577200, 
    1527580800, 1527584400, 1527588000, 1527591600, 1527595200, 1527598800, 
    1527602400, 1527606000, 1527609600, 1527613200, 1527616800, 1527620400, 
    1527624000, 1527627600, 1527631200, 1527634800, 1527638400, 1527642000, 
    1527645600, 1527649200, 1527652800, 1527656400, 1527660000, 1527663600, 
    1527667200, 1527670800, 1527674400, 1527678000, 1527681600, 1527685200, 
    1527688800, 1527692400, 1527696000, 1527699600, 1527703200, 1527706800, 
    1527710400, 1527714000, 1527717600, 1527721200, 1527724800, 1527728400, 
    1527732000, 1527735600, 1527739200, 1527742800, 1527746400, 1527750000, 
    1527753600, 1527757200, 1527760800, 1527764400, 1527768000, 1527771600, 
    1527775200, 1527778800, 1527782400, 1527786000, 1527789600, 1527793200, 
    1527796800, 1527800400, 1527804000, 1527807600, 1527811200, 1527814800, 
    1527818400, 1527822000, 1527825600, 1527829200, 1527832800, 1527836400, 
    1527840000, 1527843600, 1527847200, 1527850800, 1527854400, 1527858000, 
    1527861600, 1527865200, 1527868800, 1527872400, 1527876000, 1527879600, 
    1527883200, 1527886800, 1527890400, 1527894000, 1527897600, 1527901200, 
    1527904800, 1527908400, 1527912000, 1527915600, 1527919200, 1527922800, 
    1527926400, 1527930000, 1527933600, 1527937200, 1527940800, 1527944400, 
    1527948000, 1527951600, 1527955200, 1527958800, 1527962400, 1527966000, 
    1527969600, 1527973200, 1527976800, 1527980400, 1527984000, 1527987600, 
    1527991200, 1527994800, 1527998400, 1528002000, 1528005600, 1528009200, 
    1528012800, 1528016400, 1528020000, 1528023600, 1528027200, 1528030800, 
    1528034400, 1528038000, 1528041600, 1528045200, 1528048800, 1528052400, 
    1528056000, 1528059600, 1528063200, 1528066800, 1528070400, 1528074000, 
    1528077600, 1528081200, 1528084800, 1528088400, 1528092000, 1528095600, 
    1528099200, 1528102800, 1528106400, 1528110000, 1528113600, 1528117200, 
    1528120800, 1528124400, 1528128000, 1528131600, 1528135200, 1528138800, 
    1528142400, 1528146000, 1528149600, 1528153200, 1528156800, 1528160400, 
    1528164000, 1528167600, 1528171200, 1528174800, 1528178400, 1528182000, 
    1528185600, 1528189200, 1528192800, 1528196400, 1528200000, 1528203600, 
    1528207200, 1528210800, 1528214400, 1528218000, 1528221600, 1528225200, 
    1528228800, 1528232400, 1528236000, 1528239600, 1528243200, 1528246800, 
    1528250400, 1528254000, 1528257600, 1528261200, 1528264800, 1528268400, 
    1528272000, 1528275600, 1528279200, 1528282800, 1528286400, 1528290000, 
    1528293600, 1528297200, 1528300800, 1528304400, 1528308000, 1528311600, 
    1528315200, 1528318800, 1528322400, 1528326000, 1528329600, 1528333200, 
    1528336800, 1528340400, 1528344000, 1528347600, 1528351200, 1528354800, 
    1528358400, 1528362000, 1528365600, 1528369200, 1528372800, 1528376400, 
    1528380000, 1528383600, 1528387200, 1528390800, 1528394400, 1528398000, 
    1528401600, 1528405200, 1528408800, 1528412400, 1528416000, 1528419600, 
    1528423200, 1528426800, 1528430400, 1528434000, 1528437600, 1528441200, 
    1528444800, 1528448400, 1528452000, 1528455600, 1528459200, 1528462800, 
    1528466400, 1528470000, 1528473600, 1528477200, 1528480800, 1528484400, 
    1528488000, 1528491600, 1528495200, 1528498800, 1528502400, 1528506000, 
    1528509600, 1528513200, 1528516800, 1528520400, 1528524000, 1528527600, 
    1528531200, 1528534800, 1528538400, 1528542000, 1528545600, 1528549200, 
    1528552800, 1528556400, 1528560000, 1528563600, 1528567200, 1528570800, 
    1528574400, 1528578000, 1528581600, 1528585200, 1528588800, 1528592400, 
    1528596000, 1528599600, 1528603200, 1528606800, 1528610400, 1528614000, 
    1528617600, 1528621200, 1528624800, 1528628400, 1528632000, 1528635600, 
    1528639200, 1528642800, 1528646400, 1528650000, 1528653600, 1528657200, 
    1528660800, 1528664400, 1528668000, 1528671600, 1528675200, 1528678800, 
    1528682400, 1528686000, 1528689600, 1528693200, 1528696800, 1528700400, 
    1528704000, 1528707600, 1528711200, 1528714800, 1528718400, 1528722000, 
    1528725600, 1528729200, 1528732800, 1528736400, 1528740000, 1528743600, 
    1528747200, 1528750800, 1528754400, 1528758000, 1528761600, 1528765200, 
    1528768800, 1528772400, 1528776000, 1528779600, 1528783200, 1528786800, 
    1528790400, 1528794000, 1528797600, 1528801200, 1528804800, 1528808400, 
    1528812000, 1528815600, 1528819200, 1528822800, 1528826400, 1528830000, 
    1528833600, 1528837200, 1528840800, 1528844400, 1528848000, 1528851600, 
    1528855200, 1528858800, 1528862400, 1528866000, 1528869600, 1528873200, 
    1528876800, 1528880400, 1528884000, 1528887600, 1528891200, 1528894800, 
    1528898400, 1528902000, 1528905600, 1528909200, 1528912800, 1528916400, 
    1528920000, 1528923600, 1528927200, 1528930800, 1528934400, 1528938000, 
    1528941600, 1528945200, 1528948800, 1528952400, 1528956000, 1528959600, 
    1528963200, 1528966800, 1528970400, 1528974000, 1528977600, 1528981200, 
    1528984800, 1528988400, 1528992000, 1528995600, 1528999200, 1529002800, 
    1529006400, 1529010000, 1529013600, 1529017200, 1529020800, 1529024400, 
    1529028000, 1529031600, 1529035200, 1529038800, 1529042400, 1529046000, 
    1529049600, 1529053200, 1529056800, 1529060400, 1529064000, 1529067600, 
    1529071200, 1529074800, 1529078400, 1529082000, 1529085600, 1529089200, 
    1529092800, 1529096400, 1529100000, 1529103600, 1529107200, 1529110800, 
    1529114400, 1529118000, 1529121600, 1529125200, 1529128800, 1529132400, 
    1529136000, 1529139600, 1529143200, 1529146800, 1529150400, 1529154000, 
    1529157600, 1529161200, 1529164800, 1529168400, 1529172000, 1529175600, 
    1529179200, 1529182800, 1529186400, 1529190000, 1529193600, 1529197200, 
    1529200800, 1529204400, 1529208000, 1529211600, 1529215200, 1529218800, 
    1529222400, 1529226000, 1529229600, 1529233200, 1529236800, 1529240400, 
    1529244000, 1529247600, 1529251200, 1529254800, 1529258400, 1529262000, 
    1529265600, 1529269200, 1529272800, 1529276400, 1529280000, 1529283600, 
    1529287200, 1529290800, 1529294400, 1529298000, 1529301600, 1529305200, 
    1529308800, 1529312400, 1529316000, 1529319600, 1529323200, 1529326800, 
    1529330400, 1529334000, 1529337600, 1529341200, 1529344800, 1529348400, 
    1529352000, 1529355600, 1529359200, 1529362800, 1529366400, 1529370000, 
    1529373600, 1529377200, 1529380800, 1529384400, 1529388000, 1529391600, 
    1529395200, 1529398800, 1529402400, 1529406000, 1529409600, 1529413200, 
    1529416800, 1529420400, 1529424000, 1529427600, 1529431200, 1529434800, 
    1529438400, 1529442000, 1529445600, 1529449200, 1529452800, 1529456400, 
    1529460000, 1529463600, 1529467200, 1529470800, 1529474400, 1529478000, 
    1529481600, 1529485200, 1529488800, 1529492400, 1529496000, 1529499600, 
    1529503200, 1529506800, 1529510400, 1529514000, 1529517600, 1529521200, 
    1529524800, 1529528400, 1529532000, 1529535600, 1529539200, 1529542800, 
    1529546400, 1529550000, 1529553600, 1529557200, 1529560800, 1529564400, 
    1529568000, 1529571600, 1529575200, 1529578800, 1529582400, 1529586000, 
    1529589600, 1529593200, 1529596800, 1529600400, 1529604000, 1529607600, 
    1529611200, 1529614800, 1529618400, 1529622000, 1529625600, 1529629200, 
    1529632800, 1529636400, 1529640000, 1529643600, 1529647200, 1529650800, 
    1529654400, 1529658000, 1529661600, 1529665200, 1529668800, 1529672400, 
    1529676000, 1529679600, 1529683200, 1529686800, 1529690400, 1529694000, 
    1529697600, 1529701200, 1529704800, 1529708400, 1529712000, 1529715600, 
    1529719200, 1529722800, 1529726400, 1529730000, 1529733600, 1529737200, 
    1529740800, 1529744400, 1529748000, 1529751600, 1529755200, 1529758800, 
    1529762400, 1529766000, 1529769600, 1529773200, 1529776800, 1529780400, 
    1529784000, 1529787600, 1529791200, 1529794800, 1529798400, 1529802000, 
    1529805600, 1529809200, 1529812800, 1529816400, 1529820000, 1529823600, 
    1529827200, 1529830800, 1529834400, 1529838000, 1529841600, 1529845200, 
    1529848800, 1529852400, 1529856000, 1529859600, 1529863200, 1529866800, 
    1529870400, 1529874000, 1529877600, 1529881200, 1529884800, 1529888400, 
    1529892000, 1529895600, 1529899200, 1529902800, 1529906400, 1529910000, 
    1529913600, 1529917200, 1529920800, 1529924400, 1529928000, 1529931600, 
    1529935200, 1529938800, 1529942400, 1529946000, 1529949600, 1529953200, 
    1529956800, 1529960400, 1529964000, 1529967600, 1529971200, 1529974800, 
    1529978400, 1529982000, 1529985600, 1529989200, 1529992800, 1529996400, 
    1530000000, 1530003600, 1530007200, 1530010800, 1530014400, 1530018000, 
    1530021600, 1530025200, 1530028800, 1530032400, 1530036000, 1530039600, 
    1530043200, 1530046800, 1530050400, 1530054000, 1530057600, 1530061200, 
    1530064800, 1530068400, 1530072000, 1530075600, 1530079200, 1530082800, 
    1530086400, 1530090000, 1530093600, 1530097200, 1530100800, 1530104400, 
    1530108000, 1530111600, 1530115200, 1530118800, 1530122400, 1530126000, 
    1530129600, 1530133200, 1530136800, 1530140400, 1530144000, 1530147600, 
    1530151200, 1530154800, 1530158400, 1530162000, 1530165600, 1530169200, 
    1530172800, 1530176400, 1530180000, 1530183600, 1530187200, 1530190800, 
    1530194400, 1530198000, 1530201600, 1530205200, 1530208800, 1530212400, 
    1530216000, 1530219600, 1530223200, 1530226800, 1530230400, 1530234000, 
    1530237600, 1530241200, 1530244800, 1530248400, 1530252000, 1530255600, 
    1530259200, 1530262800, 1530266400, 1530270000, 1530273600, 1530277200, 
    1530280800, 1530284400, 1530288000, 1530291600, 1530295200, 1530298800, 
    1530302400, 1530306000, 1530309600, 1530313200, 1530316800, 1530320400, 
    1530324000, 1530327600, 1530331200, 1530334800, 1530338400, 1530342000, 
    1530345600, 1530349200, 1530352800, 1530356400, 1530360000, 1530363600, 
    1530367200, 1530370800, 1530374400, 1530378000, 1530381600, 1530385200, 
    1530388800, 1530392400, 1530396000, 1530399600, 1530403200, 1530406800, 
    1530410400, 1530414000, 1530417600, 1530421200, 1530424800, 1530428400, 
    1530432000, 1530435600, 1530439200, 1530442800, 1530446400, 1530450000, 
    1530453600, 1530457200, 1530460800, 1530464400, 1530468000, 1530471600, 
    1530475200, 1530478800, 1530482400, 1530486000, 1530489600, 1530493200, 
    1530496800, 1530500400, 1530504000, 1530507600, 1530511200, 1530514800, 
    1530518400, 1530522000, 1530525600, 1530529200, 1530532800, 1530536400, 
    1530540000, 1530543600, 1530547200, 1530550800, 1530554400, 1530558000, 
    1530561600, 1530565200, 1530568800, 1530572400, 1530576000, 1530579600, 
    1530583200, 1530586800, 1530590400, 1530594000, 1530597600, 1530601200, 
    1530604800, 1530608400, 1530612000, 1530615600, 1530619200, 1530622800, 
    1530626400, 1530630000, 1530633600, 1530637200, 1530640800, 1530644400, 
    1530648000, 1530651600, 1530655200, 1530658800, 1530662400, 1530666000, 
    1530669600, 1530673200, 1530676800, 1530680400, 1530684000, 1530687600, 
    1530691200, 1530694800, 1530698400, 1530702000, 1530705600, 1530709200, 
    1530712800, 1530716400, 1530720000, 1530723600, 1530727200, 1530730800, 
    1530734400, 1530738000, 1530741600, 1530745200, 1530748800, 1530752400, 
    1530756000, 1530759600, 1530763200, 1530766800, 1530770400, 1530774000, 
    1530777600, 1530781200, 1530784800, 1530788400, 1530792000, 1530795600, 
    1530799200, 1530802800, 1530806400, 1530810000, 1530813600, 1530817200, 
    1530820800, 1530824400, 1530828000, 1530831600, 1530835200, 1530838800, 
    1530842400, 1530846000, 1530849600, 1530853200, 1530856800, 1530860400, 
    1530864000, 1530867600, 1530871200, 1530874800, 1530878400, 1530882000, 
    1530885600, 1530889200, 1530892800, 1530896400, 1530900000, 1530903600, 
    1530907200, 1530910800, 1530914400, 1530918000, 1530921600, 1530925200, 
    1530928800, 1530932400, 1530936000, 1530939600, 1530943200, 1530946800, 
    1530950400, 1530954000, 1530957600, 1530961200, 1530964800, 1530968400, 
    1530972000, 1530975600, 1530979200, 1530982800, 1530986400, 1530990000, 
    1530993600, 1530997200, 1531000800, 1531004400, 1531008000, 1531011600, 
    1531015200, 1531018800, 1531022400, 1531026000, 1531029600, 1531033200, 
    1531036800, 1531040400, 1531044000, 1531047600, 1531051200, 1531054800, 
    1531058400, 1531062000, 1531065600, 1531069200, 1531072800, 1531076400, 
    1531080000, 1531083600, 1531087200, 1531090800, 1531094400, 1531098000, 
    1531101600, 1531105200, 1531108800, 1531112400, 1531116000, 1531119600, 
    1531123200, 1531126800, 1531130400, 1531134000, 1531137600, 1531141200, 
    1531144800, 1531148400, 1531152000, 1531155600, 1531159200, 1531162800, 
    1531166400, 1531170000, 1531173600, 1531177200, 1531180800, 1531184400, 
    1531188000, 1531191600, 1531195200, 1531198800, 1531202400, 1531206000, 
    1531209600, 1531213200, 1531216800, 1531220400, 1531224000, 1531227600, 
    1531231200, 1531234800, 1531238400, 1531242000, 1531245600, 1531249200, 
    1531252800, 1531256400, 1531260000, 1531263600, 1531267200, 1531270800, 
    1531274400, 1531278000, 1531281600, 1531285200, 1531288800, 1531292400, 
    1531296000, 1531299600, 1531303200, 1531306800, 1531310400, 1531314000, 
    1531317600, 1531321200, 1531324800, 1531328400, 1531332000, 1531335600, 
    1531339200, 1531342800, 1531346400, 1531350000, 1531353600, 1531357200, 
    1531360800, 1531364400, 1531368000, 1531371600, 1531375200, 1531378800, 
    1531382400, 1531386000, 1531389600, 1531393200, 1531396800, 1531400400, 
    1531404000, 1531407600, 1531411200, 1531414800, 1531418400, 1531422000, 
    1531425600, 1531429200, 1531432800, 1531436400, 1531440000, 1531443600, 
    1531447200, 1531450800, 1531454400, 1531458000, 1531461600, 1531465200, 
    1531468800, 1531472400, 1531476000, 1531479600, 1531483200, 1531486800, 
    1531490400, 1531494000, 1531497600, 1531501200, 1531504800, 1531508400, 
    1531512000, 1531515600, 1531519200, 1531522800, 1531526400, 1531530000, 
    1531533600, 1531537200, 1531540800, 1531544400, 1531548000, 1531551600, 
    1531555200, 1531558800, 1531562400, 1531566000, 1531569600, 1531573200, 
    1531576800, 1531580400, 1531584000, 1531587600, 1531591200, 1531594800, 
    1531598400, 1531602000, 1531605600, 1531609200, 1531612800, 1531616400, 
    1531620000, 1531623600, 1531627200, 1531630800, 1531634400, 1531638000, 
    1531641600, 1531645200, 1531648800, 1531652400, 1531656000, 1531659600, 
    1531663200, 1531666800, 1531670400, 1531674000, 1531677600, 1531681200, 
    1531684800, 1531688400, 1531692000, 1531695600, 1531699200, 1531702800, 
    1531706400, 1531710000, 1531713600, 1531717200, 1531720800, 1531724400, 
    1531728000, 1531731600, 1531735200, 1531738800, 1531742400, 1531746000, 
    1531749600, 1531753200, 1531756800, 1531760400, 1531764000, 1531767600, 
    1531771200, 1531774800, 1531778400, 1531782000, 1531785600, 1531789200, 
    1531792800, 1531796400, 1531800000, 1531803600, 1531807200, 1531810800, 
    1531814400, 1531818000, 1531821600, 1531825200, 1531828800, 1531832400, 
    1531836000, 1531839600, 1531843200, 1531846800, 1531850400, 1531854000, 
    1531857600, 1531861200, 1531864800, 1531868400, 1531872000, 1531875600, 
    1531879200, 1531882800, 1531886400, 1531890000, 1531893600, 1531897200, 
    1531900800, 1531904400, 1531908000, 1531911600, 1531915200, 1531918800, 
    1531922400, 1531926000, 1531929600, 1531933200, 1531936800, 1531940400, 
    1531944000, 1531947600, 1531951200, 1531954800, 1531958400, 1531962000, 
    1531965600, 1531969200, 1531972800, 1531976400, 1531980000, 1531983600, 
    1531987200, 1531990800, 1531994400, 1531998000, 1532001600, 1532005200, 
    1532008800, 1532012400, 1532016000, 1532019600, 1532023200, 1532026800, 
    1532030400, 1532034000, 1532037600, 1532041200, 1532044800, 1532048400, 
    1532052000, 1532055600, 1532059200, 1532062800, 1532066400, 1532070000, 
    1532073600, 1532077200, 1532080800, 1532084400, 1532088000, 1532091600, 
    1532095200, 1532098800, 1532102400, 1532106000, 1532109600, 1532113200, 
    1532116800, 1532120400, 1532124000, 1532127600, 1532131200, 1532134800, 
    1532138400, 1532142000, 1532145600, 1532149200, 1532152800, 1532156400, 
    1532160000, 1532163600, 1532167200, 1532170800, 1532174400, 1532178000, 
    1532181600, 1532185200, 1532188800, 1532192400, 1532196000, 1532199600, 
    1532203200, 1532206800, 1532210400, 1532214000, 1532217600, 1532221200, 
    1532224800, 1532228400, 1532232000, 1532235600, 1532239200, 1532242800, 
    1532246400, 1532250000, 1532253600, 1532257200, 1532260800, 1532264400, 
    1532268000, 1532271600, 1532275200, 1532278800, 1532282400, 1532286000, 
    1532289600, 1532293200, 1532296800, 1532300400, 1532304000, 1532307600, 
    1532311200, 1532314800, 1532318400, 1532322000, 1532325600, 1532329200, 
    1532332800, 1532336400, 1532340000, 1532343600, 1532347200, 1532350800, 
    1532354400, 1532358000, 1532361600, 1532365200, 1532368800, 1532372400, 
    1532376000, 1532379600, 1532383200, 1532386800, 1532390400, 1532394000, 
    1532397600, 1532401200, 1532404800, 1532408400, 1532412000, 1532415600, 
    1532419200, 1532422800, 1532426400, 1532430000, 1532433600, 1532437200, 
    1532440800, 1532444400, 1532448000, 1532451600, 1532455200, 1532458800, 
    1532462400, 1532466000, 1532469600, 1532473200, 1532476800, 1532480400, 
    1532484000, 1532487600, 1532491200, 1532494800, 1532498400, 1532502000, 
    1532505600, 1532509200, 1532512800, 1532516400, 1532520000, 1532523600, 
    1532527200, 1532530800, 1532534400, 1532538000, 1532541600, 1532545200, 
    1532548800, 1532552400, 1532556000, 1532559600, 1532563200, 1532566800, 
    1532570400, 1532574000, 1532577600, 1532581200, 1532584800, 1532588400, 
    1532592000, 1532595600, 1532599200, 1532602800, 1532606400, 1532610000, 
    1532613600, 1532617200, 1532620800, 1532624400, 1532628000, 1532631600, 
    1532635200, 1532638800, 1532642400, 1532646000, 1532649600, 1532653200, 
    1532656800, 1532660400, 1532664000, 1532667600, 1532671200, 1532674800, 
    1532678400, 1532682000, 1532685600, 1532689200, 1532692800, 1532696400, 
    1532700000, 1532703600, 1532707200, 1532710800, 1532714400, 1532718000, 
    1532721600, 1532725200, 1532728800, 1532732400, 1532736000, 1532739600, 
    1532743200, 1532746800, 1532750400, 1532754000, 1532757600, 1532761200, 
    1532764800, 1532768400, 1532772000, 1532775600, 1532779200, 1532782800, 
    1532786400, 1532790000, 1532793600, 1532797200, 1532800800, 1532804400, 
    1532808000, 1532811600, 1532815200, 1532818800, 1532822400, 1532826000, 
    1532829600, 1532833200, 1532836800, 1532840400, 1532844000, 1532847600, 
    1532851200, 1532854800, 1532858400, 1532862000, 1532865600, 1532869200, 
    1532872800, 1532876400, 1532880000, 1532883600, 1532887200, 1532890800, 
    1532894400, 1532898000, 1532901600, 1532905200, 1532908800, 1532912400, 
    1532916000, 1532919600, 1532923200, 1532926800, 1532930400, 1532934000, 
    1532937600, 1532941200, 1532944800, 1532948400, 1532952000, 1532955600, 
    1532959200, 1532962800, 1532966400, 1532970000, 1532973600, 1532977200, 
    1532980800, 1532984400, 1532988000, 1532991600, 1532995200, 1532998800, 
    1533002400, 1533006000, 1533009600, 1533013200, 1533016800, 1533020400, 
    1533024000, 1533027600, 1533031200, 1533034800, 1533038400, 1533042000, 
    1533045600, 1533049200, 1533052800, 1533056400, 1533060000, 1533063600, 
    1533067200, 1533070800, 1533074400, 1533078000, 1533081600, 1533085200, 
    1533088800, 1533092400, 1533096000, 1533099600, 1533103200, 1533106800, 
    1533110400, 1533114000, 1533117600, 1533121200, 1533124800, 1533128400, 
    1533132000, 1533135600, 1533139200, 1533142800, 1533146400, 1533150000, 
    1533153600, 1533157200, 1533160800, 1533164400, 1533168000, 1533171600, 
    1533175200, 1533178800, 1533182400, 1533186000, 1533189600, 1533193200, 
    1533196800, 1533200400, 1533204000, 1533207600, 1533211200, 1533214800, 
    1533218400, 1533222000, 1533225600, 1533229200, 1533232800, 1533236400, 
    1533240000, 1533243600, 1533247200, 1533250800, 1533254400, 1533258000, 
    1533261600, 1533265200, 1533268800, 1533272400, 1533276000, 1533279600, 
    1533283200, 1533286800, 1533290400, 1533294000, 1533297600, 1533301200, 
    1533304800, 1533308400, 1533312000, 1533315600, 1533319200, 1533322800, 
    1533326400, 1533330000, 1533333600, 1533337200, 1533340800, 1533344400, 
    1533348000, 1533351600, 1533355200, 1533358800, 1533362400, 1533366000, 
    1533369600, 1533373200, 1533376800, 1533380400, 1533384000, 1533387600, 
    1533391200, 1533394800, 1533398400, 1533402000, 1533405600, 1533409200, 
    1533412800, 1533416400, 1533420000, 1533423600, 1533427200, 1533430800, 
    1533434400, 1533438000, 1533441600, 1533445200, 1533448800, 1533452400, 
    1533456000, 1533459600, 1533463200, 1533466800, 1533470400, 1533474000, 
    1533477600, 1533481200, 1533484800, 1533488400, 1533492000, 1533495600, 
    1533499200, 1533502800, 1533506400, 1533510000, 1533513600, 1533517200, 
    1533520800, 1533524400, 1533528000, 1533531600, 1533535200, 1533538800, 
    1533542400, 1533546000, 1533549600, 1533553200, 1533556800, 1533560400, 
    1533564000, 1533567600, 1533571200, 1533574800, 1533578400, 1533582000, 
    1533585600, 1533589200, 1533592800, 1533596400, 1533600000, 1533603600, 
    1533607200, 1533610800, 1533614400, 1533618000, 1533621600, 1533625200, 
    1533628800, 1533632400, 1533636000, 1533639600, 1533643200, 1533646800, 
    1533650400, 1533654000, 1533657600, 1533661200, 1533664800, 1533668400, 
    1533672000, 1533675600, 1533679200, 1533682800, 1533686400, 1533690000, 
    1533693600, 1533697200, 1533700800, 1533704400, 1533708000, 1533711600, 
    1533715200, 1533718800, 1533722400, 1533726000, 1533729600, 1533733200, 
    1533736800, 1533740400, 1533744000, 1533747600, 1533751200, 1533754800, 
    1533758400, 1533762000, 1533765600, 1533769200, 1533772800, 1533776400, 
    1533780000, 1533783600, 1533787200, 1533790800, 1533794400, 1533798000, 
    1533801600, 1533805200, 1533808800, 1533812400, 1533816000, 1533819600, 
    1533823200, 1533826800, 1533830400, 1533834000, 1533837600, 1533841200, 
    1533844800, 1533848400, 1533852000, 1533855600, 1533859200, 1533862800, 
    1533866400, 1533870000, 1533873600, 1533877200, 1533880800, 1533884400, 
    1533888000, 1533891600, 1533895200, 1533898800, 1533902400, 1533906000, 
    1533909600, 1533913200, 1533916800, 1533920400, 1533924000, 1533927600, 
    1533931200, 1533934800, 1533938400, 1533942000, 1533945600, 1533949200, 
    1533952800, 1533956400, 1533960000, 1533963600, 1533967200, 1533970800, 
    1533974400, 1533978000, 1533981600, 1533985200, 1533988800, 1533992400, 
    1533996000, 1533999600, 1534003200, 1534006800, 1534010400, 1534014000, 
    1534017600, 1534021200, 1534024800, 1534028400, 1534032000, 1534035600, 
    1534039200, 1534042800, 1534046400, 1534050000, 1534053600, 1534057200, 
    1534060800, 1534064400, 1534068000, 1534071600, 1534075200, 1534078800, 
    1534082400, 1534086000, 1534089600, 1534093200, 1534096800, 1534100400, 
    1534104000, 1534107600, 1534111200, 1534114800, 1534118400, 1534122000, 
    1534125600, 1534129200, 1534132800, 1534136400, 1534140000, 1534143600, 
    1534147200, 1534150800, 1534154400, 1534158000, 1534161600, 1534165200, 
    1534168800, 1534172400, 1534176000, 1534179600, 1534183200, 1534186800, 
    1534190400, 1534194000, 1534197600, 1534201200, 1534204800, 1534208400, 
    1534212000, 1534215600, 1534219200, 1534222800, 1534226400, 1534230000, 
    1534233600, 1534237200, 1534240800, 1534244400, 1534248000, 1534251600, 
    1534255200, 1534258800, 1534262400, 1534266000, 1534269600, 1534273200, 
    1534276800, 1534280400, 1534284000, 1534287600, 1534291200, 1534294800, 
    1534298400, 1534302000, 1534305600, 1534309200, 1534312800, 1534316400, 
    1534320000, 1534323600, 1534327200, 1534330800, 1534334400, 1534338000, 
    1534341600, 1534345200, 1534348800, 1534352400, 1534356000, 1534359600, 
    1534363200, 1534366800, 1534370400, 1534374000, 1534377600, 1534381200, 
    1534384800, 1534388400, 1534392000, 1534395600, 1534399200, 1534402800, 
    1534406400, 1534410000, 1534413600, 1534417200, 1534420800, 1534424400, 
    1534428000, 1534431600, 1534435200, 1534438800, 1534442400, 1534446000, 
    1534449600, 1534453200, 1534456800, 1534460400, 1534464000, 1534467600, 
    1534471200, 1534474800, 1534478400, 1534482000, 1534485600, 1534489200, 
    1534492800, 1534496400, 1534500000, 1534503600, 1534507200, 1534510800, 
    1534514400, 1534518000, 1534521600, 1534525200, 1534528800, 1534532400, 
    1534536000, 1534539600, 1534543200, 1534546800, 1534550400, 1534554000, 
    1534557600, 1534561200, 1534564800, 1534568400, 1534572000, 1534575600, 
    1534579200, 1534582800, 1534586400, 1534590000, 1534593600, 1534597200, 
    1534600800, 1534604400, 1534608000, 1534611600, 1534615200, 1534618800, 
    1534622400, 1534626000, 1534629600, 1534633200, 1534636800, 1534640400, 
    1534644000, 1534647600, 1534651200, 1534654800, 1534658400, 1534662000, 
    1534665600, 1534669200, 1534672800, 1534676400, 1534680000, 1534683600, 
    1534687200, 1534690800, 1534694400, 1534698000, 1534701600, 1534705200, 
    1534708800, 1534712400, 1534716000, 1534719600, 1534723200, 1534726800, 
    1534730400, 1534734000, 1534737600, 1534741200, 1534744800, 1534748400, 
    1534752000, 1534755600, 1534759200, 1534762800, 1534766400, 1534770000, 
    1534773600, 1534777200, 1534780800, 1534784400, 1534788000, 1534791600, 
    1534795200, 1534798800, 1534802400, 1534806000, 1534809600, 1534813200, 
    1534816800, 1534820400, 1534824000, 1534827600, 1534831200, 1534834800, 
    1534838400, 1534842000, 1534845600, 1534849200, 1534852800, 1534856400, 
    1534860000, 1534863600, 1534867200, 1534870800, 1534874400, 1534878000, 
    1534881600, 1534885200, 1534888800, 1534892400, 1534896000, 1534899600, 
    1534903200, 1534906800, 1534910400, 1534914000, 1534917600, 1534921200, 
    1534924800, 1534928400, 1534932000, 1534935600, 1534939200, 1534942800, 
    1534946400, 1534950000, 1534953600, 1534957200, 1534960800, 1534964400, 
    1534968000, 1534971600, 1534975200, 1534978800, 1534982400, 1534986000, 
    1534989600, 1534993200, 1534996800, 1535000400, 1535004000, 1535007600, 
    1535011200, 1535014800, 1535018400, 1535022000, 1535025600, 1535029200, 
    1535032800, 1535036400, 1535040000, 1535043600, 1535047200, 1535050800, 
    1535054400, 1535058000, 1535061600, 1535065200, 1535068800, 1535072400, 
    1535076000, 1535079600, 1535083200, 1535086800, 1535090400, 1535094000, 
    1535097600, 1535101200, 1535104800, 1535108400, 1535112000, 1535115600, 
    1535119200, 1535122800, 1535126400, 1535130000, 1535133600, 1535137200, 
    1535140800, 1535144400, 1535148000, 1535151600, 1535155200, 1535158800, 
    1535162400, 1535166000, 1535169600, 1535173200, 1535176800, 1535180400, 
    1535184000, 1535187600, 1535191200, 1535194800, 1535198400, 1535202000, 
    1535205600, 1535209200, 1535212800, 1535216400, 1535220000, 1535223600, 
    1535227200, 1535230800, 1535234400, 1535238000, 1535241600, 1535245200, 
    1535248800, 1535252400, 1535256000, 1535259600, 1535263200, 1535266800, 
    1535270400, 1535274000, 1535277600, 1535281200, 1535284800, 1535288400, 
    1535292000, 1535295600, 1535299200, 1535302800, 1535306400, 1535310000, 
    1535313600, 1535317200, 1535320800, 1535324400, 1535328000, 1535331600, 
    1535335200, 1535338800, 1535342400, 1535346000, 1535349600, 1535353200, 
    1535356800, 1535360400, 1535364000, 1535367600, 1535371200, 1535374800, 
    1535378400, 1535382000, 1535385600, 1535389200, 1535392800, 1535396400, 
    1535400000, 1535403600, 1535407200, 1535410800, 1535414400, 1535418000, 
    1535421600, 1535425200, 1535428800, 1535432400, 1535436000, 1535439600, 
    1535443200, 1535446800, 1535450400, 1535454000, 1535457600, 1535461200, 
    1535464800, 1535468400, 1535472000, 1535475600, 1535479200, 1535482800, 
    1535486400, 1535490000, 1535493600, 1535497200, 1535500800, 1535504400, 
    1535508000, 1535511600, 1535515200, 1535518800, 1535522400, 1535526000, 
    1535529600, 1535533200, 1535536800, 1535540400, 1535544000, 1535547600, 
    1535551200, 1535554800, 1535558400, 1535562000, 1535565600, 1535569200, 
    1535572800, 1535576400, 1535580000, 1535583600, 1535587200, 1535590800, 
    1535594400, 1535598000, 1535601600, 1535605200, 1535608800, 1535612400, 
    1535616000, 1535619600, 1535623200, 1535626800, 1535630400, 1535634000, 
    1535637600, 1535641200, 1535644800, 1535648400, 1535652000, 1535655600, 
    1535659200, 1535662800, 1535666400, 1535670000, 1535673600, 1535677200, 
    1535680800, 1535684400, 1535688000, 1535691600, 1535695200, 1535698800, 
    1535702400, 1535706000, 1535709600, 1535713200, 1535716800, 1535720400, 
    1535724000, 1535727600, 1535731200, 1535734800, 1535738400, 1535742000, 
    1535745600, 1535749200, 1535752800, 1535756400, 1535760000, 1535763600, 
    1535767200, 1535770800, 1535774400, 1535778000, 1535781600, 1535785200, 
    1535788800, 1535792400, 1535796000, 1535799600, 1535803200, 1535806800, 
    1535810400, 1535814000, 1535817600, 1535821200, 1535824800, 1535828400, 
    1535832000, 1535835600, 1535839200, 1535842800, 1535846400, 1535850000, 
    1535853600, 1535857200, 1535860800, 1535864400, 1535868000, 1535871600, 
    1535875200, 1535878800, 1535882400, 1535886000, 1535889600, 1535893200, 
    1535896800, 1535900400, 1535904000, 1535907600, 1535911200, 1535914800, 
    1535918400, 1535922000, 1535925600, 1535929200, 1535932800, 1535936400, 
    1535940000, 1535943600, 1535947200, 1535950800, 1535954400, 1535958000, 
    1535961600, 1535965200, 1535968800, 1535972400, 1535976000, 1535979600, 
    1535983200, 1535986800, 1535990400, 1535994000, 1535997600, 1536001200, 
    1536004800, 1536008400, 1536012000, 1536015600, 1536019200, 1536022800, 
    1536026400, 1536030000, 1536033600, 1536037200, 1536040800, 1536044400, 
    1536048000, 1536051600, 1536055200, 1536058800, 1536062400, 1536066000, 
    1536069600, 1536073200, 1536076800, 1536080400, 1536084000, 1536087600, 
    1536091200, 1536094800, 1536098400, 1536102000, 1536105600, 1536109200, 
    1536112800, 1536116400, 1536120000, 1536123600, 1536127200, 1536130800, 
    1536134400, 1536138000, 1536141600, 1536145200, 1536148800, 1536152400, 
    1536156000, 1536159600, 1536163200, 1536166800, 1536170400, 1536174000, 
    1536177600, 1536181200, 1536184800, 1536188400, 1536192000, 1536195600, 
    1536199200, 1536202800, 1536206400, 1536210000, 1536213600, 1536217200, 
    1536220800, 1536224400, 1536228000, 1536231600, 1536235200, 1536238800, 
    1536242400, 1536246000, 1536249600, 1536253200, 1536256800, 1536260400, 
    1536264000, 1536267600, 1536271200, 1536274800, 1536278400, 1536282000, 
    1536285600, 1536289200, 1536292800, 1536296400, 1536300000, 1536303600, 
    1536307200, 1536310800, 1536314400, 1536318000, 1536321600, 1536325200, 
    1536328800, 1536332400, 1536336000, 1536339600, 1536343200, 1536346800, 
    1536350400, 1536354000, 1536357600, 1536361200, 1536364800, 1536368400, 
    1536372000, 1536375600, 1536379200, 1536382800, 1536386400, 1536390000, 
    1536393600, 1536397200, 1536400800, 1536404400, 1536408000, 1536411600, 
    1536415200, 1536418800, 1536422400, 1536426000, 1536429600, 1536433200, 
    1536436800, 1536440400, 1536444000, 1536447600, 1536451200, 1536454800, 
    1536458400, 1536462000, 1536465600, 1536469200, 1536472800, 1536476400, 
    1536480000, 1536483600, 1536487200, 1536490800, 1536494400, 1536498000, 
    1536501600, 1536505200, 1536508800, 1536512400, 1536516000, 1536519600, 
    1536523200, 1536526800, 1536530400, 1536534000, 1536537600, 1536541200, 
    1536544800, 1536548400, 1536552000, 1536555600, 1536559200, 1536562800, 
    1536566400, 1536570000, 1536573600, 1536577200, 1536580800, 1536584400, 
    1536588000, 1536591600, 1536595200, 1536598800, 1536602400, 1536606000, 
    1536609600, 1536613200, 1536616800, 1536620400, 1536624000, 1536627600, 
    1536631200, 1536634800, 1536638400, 1536642000, 1536645600, 1536649200, 
    1536652800, 1536656400, 1536660000, 1536663600, 1536667200, 1536670800, 
    1536674400, 1536678000, 1536681600, 1536685200, 1536688800, 1536692400, 
    1536696000, 1536699600, 1536703200, 1536706800, 1536710400, 1536714000, 
    1536717600, 1536721200, 1536724800, 1536728400, 1536732000, 1536735600, 
    1536739200, 1536742800, 1536746400, 1536750000, 1536753600, 1536757200, 
    1536760800, 1536764400, 1536768000, 1536771600, 1536775200, 1536778800, 
    1536782400, 1536786000, 1536789600, 1536793200, 1536796800, 1536800400, 
    1536804000, 1536807600, 1536811200, 1536814800, 1536818400, 1536822000, 
    1536825600, 1536829200, 1536832800, 1536836400, 1536840000, 1536843600, 
    1536847200, 1536850800, 1536854400, 1536858000, 1536861600, 1536865200, 
    1536868800, 1536872400, 1536876000, 1536879600, 1536883200, 1536886800, 
    1536890400, 1536894000, 1536897600, 1536901200, 1536904800, 1536908400, 
    1536912000, 1536915600, 1536919200, 1536922800, 1536926400, 1536930000, 
    1536933600, 1536937200, 1536940800, 1536944400, 1536948000, 1536951600, 
    1536955200, 1536958800, 1536962400, 1536966000, 1536969600, 1536973200, 
    1536976800, 1536980400, 1536984000, 1536987600, 1536991200, 1536994800, 
    1536998400, 1537002000, 1537005600, 1537009200, 1537012800, 1537016400, 
    1537020000, 1537023600, 1537027200, 1537030800, 1537034400, 1537038000, 
    1537041600, 1537045200, 1537048800, 1537052400, 1537056000, 1537059600, 
    1537063200, 1537066800, 1537070400, 1537074000, 1537077600, 1537081200, 
    1537084800, 1537088400, 1537092000, 1537095600, 1537099200, 1537102800, 
    1537106400, 1537110000, 1537113600, 1537117200, 1537120800, 1537124400, 
    1537128000, 1537131600, 1537135200, 1537138800, 1537142400, 1537146000, 
    1537149600, 1537153200, 1537156800, 1537160400, 1537164000, 1537167600, 
    1537171200, 1537174800, 1537178400, 1537182000, 1537185600, 1537189200, 
    1537192800, 1537196400, 1537200000, 1537203600, 1537207200, 1537210800, 
    1537214400, 1537218000, 1537221600, 1537225200, 1537228800, 1537232400, 
    1537236000, 1537239600, 1537243200, 1537246800, 1537250400, 1537254000, 
    1537257600, 1537261200, 1537264800, 1537268400, 1537272000, 1537275600, 
    1537279200, 1537282800, 1537286400, 1537290000, 1537293600, 1537297200, 
    1537300800, 1537304400, 1537308000, 1537311600, 1537315200, 1537318800, 
    1537322400, 1537326000, 1537329600, 1537333200, 1537336800, 1537340400, 
    1537344000, 1537347600, 1537351200, 1537354800, 1537358400, 1537362000, 
    1537365600, 1537369200, 1537372800, 1537376400, 1537380000, 1537383600, 
    1537387200, 1537390800, 1537394400, 1537398000, 1537401600, 1537405200, 
    1537408800, 1537412400, 1537416000, 1537419600, 1537423200, 1537426800, 
    1537430400, 1537434000, 1537437600, 1537441200, 1537444800, 1537448400, 
    1537452000, 1537455600, 1537459200, 1537462800, 1537466400, 1537470000, 
    1537473600, 1537477200, 1537480800, 1537484400, 1537488000, 1537491600, 
    1537495200, 1537498800, 1537502400, 1537506000, 1537509600, 1537513200, 
    1537516800, 1537520400, 1537524000, 1537527600, 1537531200, 1537534800, 
    1537538400, 1537542000, 1537545600, 1537549200, 1537552800, 1537556400, 
    1537560000, 1537563600, 1537567200, 1537570800, 1537574400, 1537578000, 
    1537581600, 1537585200, 1537588800, 1537592400, 1537596000, 1537599600, 
    1537603200, 1537606800, 1537610400, 1537614000, 1537617600, 1537621200, 
    1537624800, 1537628400, 1537632000, 1537635600, 1537639200, 1537642800, 
    1537646400, 1537650000, 1537653600, 1537657200, 1537660800, 1537664400, 
    1537668000, 1537671600, 1537675200, 1537678800, 1537682400, 1537686000, 
    1537689600, 1537693200, 1537696800, 1537700400, 1537704000, 1537707600, 
    1537711200, 1537714800, 1537718400, 1537722000, 1537725600, 1537729200, 
    1537732800, 1537736400, 1537740000, 1537743600, 1537747200, 1537750800, 
    1537754400, 1537758000, 1537761600, 1537765200, 1537768800, 1537772400, 
    1537776000, 1537779600, 1537783200, 1537786800, 1537790400, 1537794000, 
    1537797600, 1537801200, 1537804800, 1537808400, 1537812000, 1537815600, 
    1537819200, 1537822800, 1537826400, 1537830000, 1537833600, 1537837200, 
    1537840800, 1537844400, 1537848000, 1537851600, 1537855200, 1537858800, 
    1537862400, 1537866000, 1537869600, 1537873200, 1537876800, 1537880400, 
    1537884000, 1537887600, 1537891200, 1537894800, 1537898400, 1537902000, 
    1537905600, 1537909200, 1537912800, 1537916400, 1537920000, 1537923600, 
    1537927200, 1537930800, 1537934400, 1537938000, 1537941600, 1537945200, 
    1537948800, 1537952400, 1537956000, 1537959600, 1537963200, 1537966800, 
    1537970400, 1537974000, 1537977600, 1537981200, 1537984800, 1537988400, 
    1537992000, 1537995600, 1537999200, 1538002800, 1538006400, 1538010000, 
    1538013600, 1538017200, 1538020800, 1538024400, 1538028000, 1538031600, 
    1538035200, 1538038800, 1538042400, 1538046000, 1538049600, 1538053200, 
    1538056800, 1538060400, 1538064000, 1538067600, 1538071200, 1538074800, 
    1538078400, 1538082000, 1538085600, 1538089200, 1538092800, 1538096400, 
    1538100000, 1538103600, 1538107200, 1538110800, 1538114400, 1538118000, 
    1538121600, 1538125200, 1538128800, 1538132400, 1538136000, 1538139600, 
    1538143200, 1538146800, 1538150400, 1538154000, 1538157600, 1538161200, 
    1538164800, 1538168400, 1538172000, 1538175600, 1538179200, 1538182800, 
    1538186400, 1538190000, 1538193600, 1538197200, 1538200800, 1538204400, 
    1538208000, 1538211600, 1538215200, 1538218800, 1538222400, 1538226000, 
    1538229600, 1538233200, 1538236800, 1538240400, 1538244000, 1538247600, 
    1538251200, 1538254800, 1538258400, 1538262000, 1538265600, 1538269200, 
    1538272800, 1538276400, 1538280000, 1538283600, 1538287200, 1538290800, 
    1538294400, 1538298000, 1538301600, 1538305200, 1538308800, 1538312400, 
    1538316000, 1538319600, 1538323200, 1538326800, 1538330400, 1538334000, 
    1538337600, 1538341200, 1538344800, 1538348400, 1538352000, 1538355600, 
    1538359200, 1538362800, 1538366400, 1538370000, 1538373600, 1538377200, 
    1538380800, 1538384400, 1538388000, 1538391600, 1538395200, 1538398800, 
    1538402400, 1538406000, 1538409600, 1538413200, 1538416800, 1538420400, 
    1538424000, 1538427600, 1538431200, 1538434800, 1538438400, 1538442000, 
    1538445600, 1538449200, 1538452800, 1538456400, 1538460000, 1538463600, 
    1538467200, 1538470800, 1538474400, 1538478000, 1538481600, 1538485200, 
    1538488800, 1538492400, 1538496000, 1538499600, 1538503200, 1538506800, 
    1538510400, 1538514000, 1538517600, 1538521200, 1538524800, 1538528400, 
    1538532000, 1538535600, 1538539200, 1538542800, 1538546400, 1538550000, 
    1538553600, 1538557200, 1538560800, 1538564400, 1538568000, 1538571600, 
    1538575200, 1538578800, 1538582400, 1538586000, 1538589600, 1538593200, 
    1538596800, 1538600400, 1538604000, 1538607600, 1538611200, 1538614800, 
    1538618400, 1538622000, 1538625600, 1538629200, 1538632800, 1538636400, 
    1538640000, 1538643600, 1538647200, 1538650800, 1538654400, 1538658000, 
    1538661600, 1538665200, 1538668800, 1538672400, 1538676000, 1538679600, 
    1538683200, 1538686800, 1538690400, 1538694000, 1538697600, 1538701200, 
    1538704800, 1538708400, 1538712000, 1538715600, 1538719200, 1538722800, 
    1538726400, 1538730000, 1538733600, 1538737200, 1538740800, 1538744400, 
    1538748000, 1538751600, 1538755200, 1538758800, 1538762400, 1538766000, 
    1538769600, 1538773200, 1538776800, 1538780400, 1538784000, 1538787600, 
    1538791200, 1538794800, 1538798400, 1538802000, 1538805600, 1538809200, 
    1538812800, 1538816400, 1538820000, 1538823600, 1538827200, 1538830800, 
    1538834400, 1538838000, 1538841600, 1538845200, 1538848800, 1538852400, 
    1538856000, 1538859600, 1538863200, 1538866800, 1538870400, 1538874000, 
    1538877600, 1538881200, 1538884800, 1538888400, 1538892000, 1538895600, 
    1538899200, 1538902800, 1538906400, 1538910000, 1538913600, 1538917200, 
    1538920800, 1538924400, 1538928000, 1538931600, 1538935200, 1538938800, 
    1538942400, 1538946000, 1538949600, 1538953200, 1538956800, 1538960400, 
    1538964000, 1538967600, 1538971200, 1538974800, 1538978400, 1538982000, 
    1538985600, 1538989200, 1538992800, 1538996400, 1539000000, 1539003600, 
    1539007200, 1539010800, 1539014400, 1539018000, 1539021600, 1539025200, 
    1539028800, 1539032400, 1539036000, 1539039600, 1539043200, 1539046800, 
    1539050400, 1539054000, 1539057600, 1539061200, 1539064800, 1539068400, 
    1539072000, 1539075600, 1539079200, 1539082800, 1539086400, 1539090000, 
    1539093600, 1539097200, 1539100800, 1539104400, 1539108000, 1539111600, 
    1539115200, 1539118800, 1539122400, 1539126000, 1539129600, 1539133200, 
    1539136800, 1539140400, 1539144000, 1539147600, 1539151200, 1539154800, 
    1539158400, 1539162000, 1539165600, 1539169200, 1539172800, 1539176400, 
    1539180000, 1539183600, 1539187200, 1539190800, 1539194400, 1539198000, 
    1539201600, 1539205200, 1539208800, 1539212400, 1539216000, 1539219600, 
    1539223200, 1539226800, 1539230400, 1539234000, 1539237600, 1539241200, 
    1539244800, 1539248400, 1539252000, 1539255600, 1539259200, 1539262800, 
    1539266400, 1539270000, 1539273600, 1539277200, 1539280800, 1539284400, 
    1539288000, 1539291600, 1539295200, 1539298800, 1539302400, 1539306000, 
    1539309600, 1539313200, 1539316800, 1539320400, 1539324000, 1539327600, 
    1539331200, 1539334800, 1539338400, 1539342000, 1539345600, 1539349200, 
    1539352800, 1539356400, 1539360000, 1539363600, 1539367200, 1539370800, 
    1539374400, 1539378000, 1539381600, 1539385200, 1539388800, 1539392400, 
    1539396000, 1539399600, 1539403200, 1539406800, 1539410400, 1539414000, 
    1539417600, 1539421200, 1539424800, 1539428400, 1539432000, 1539435600, 
    1539439200, 1539442800, 1539446400, 1539450000, 1539453600, 1539457200, 
    1539460800, 1539464400, 1539468000, 1539471600, 1539475200, 1539478800, 
    1539482400, 1539486000, 1539489600, 1539493200, 1539496800, 1539500400, 
    1539504000, 1539507600, 1539511200, 1539514800, 1539518400, 1539522000, 
    1539525600, 1539529200, 1539532800, 1539536400, 1539540000, 1539543600, 
    1539547200, 1539550800, 1539554400, 1539558000, 1539561600, 1539565200, 
    1539568800, 1539572400, 1539576000, 1539579600, 1539583200, 1539586800, 
    1539590400, 1539594000, 1539597600, 1539601200, 1539604800, 1539608400, 
    1539612000, 1539615600, 1539619200, 1539622800, 1539626400, 1539630000, 
    1539633600, 1539637200, 1539640800, 1539644400, 1539648000, 1539651600, 
    1539655200, 1539658800, 1539662400, 1539666000, 1539669600, 1539673200, 
    1539676800, 1539680400, 1539684000, 1539687600, 1539691200, 1539694800, 
    1539698400, 1539702000, 1539705600, 1539709200, 1539712800, 1539716400, 
    1539720000, 1539723600, 1539727200, 1539730800, 1539734400, 1539738000, 
    1539741600, 1539745200, 1539748800, 1539752400, 1539756000, 1539759600, 
    1539763200, 1539766800, 1539770400, 1539774000, 1539777600, 1539781200, 
    1539784800, 1539788400, 1539792000, 1539795600, 1539799200, 1539802800, 
    1539806400, 1539810000, 1539813600, 1539817200, 1539820800, 1539824400, 
    1539828000, 1539831600, 1539835200, 1539838800, 1539842400, 1539846000, 
    1539849600, 1539853200, 1539856800, 1539860400, 1539864000, 1539867600, 
    1539871200, 1539874800, 1539878400, 1539882000, 1539885600, 1539889200, 
    1539892800, 1539896400, 1539900000, 1539903600, 1539907200, 1539910800, 
    1539914400, 1539918000, 1539921600, 1539925200, 1539928800, 1539932400, 
    1539936000, 1539939600, 1539943200, 1539946800, 1539950400, 1539954000, 
    1539957600, 1539961200, 1539964800, 1539968400, 1539972000, 1539975600, 
    1539979200, 1539982800, 1539986400, 1539990000, 1539993600, 1539997200, 
    1540000800, 1540004400, 1540008000, 1540011600, 1540015200, 1540018800, 
    1540022400, 1540026000, 1540029600, 1540033200, 1540036800, 1540040400, 
    1540044000, 1540047600, 1540051200, 1540054800, 1540058400, 1540062000, 
    1540065600, 1540069200, 1540072800, 1540076400, 1540080000, 1540083600, 
    1540087200, 1540090800, 1540094400, 1540098000, 1540101600, 1540105200, 
    1540108800, 1540112400, 1540116000, 1540119600, 1540123200, 1540126800, 
    1540130400, 1540134000, 1540137600, 1540141200, 1540144800, 1540148400, 
    1540152000, 1540155600, 1540159200, 1540162800, 1540166400, 1540170000, 
    1540173600, 1540177200, 1540180800, 1540184400, 1540188000, 1540191600, 
    1540195200, 1540198800, 1540202400, 1540206000, 1540209600, 1540213200, 
    1540216800, 1540220400, 1540224000, 1540227600, 1540231200, 1540234800, 
    1540238400, 1540242000, 1540245600, 1540249200, 1540252800, 1540256400, 
    1540260000, 1540263600, 1540267200, 1540270800, 1540274400, 1540278000, 
    1540281600, 1540285200, 1540288800, 1540292400, 1540296000, 1540299600, 
    1540303200, 1540306800, 1540310400, 1540314000, 1540317600, 1540321200, 
    1540324800, 1540328400, 1540332000, 1540335600, 1540339200, 1540342800, 
    1540346400, 1540350000, 1540353600, 1540357200, 1540360800, 1540364400, 
    1540368000, 1540371600, 1540375200, 1540378800, 1540382400, 1540386000, 
    1540389600, 1540393200, 1540396800, 1540400400, 1540404000, 1540407600, 
    1540411200, 1540414800, 1540418400, 1540422000, 1540425600, 1540429200, 
    1540432800, 1540436400, 1540440000, 1540443600, 1540447200, 1540450800, 
    1540454400, 1540458000, 1540461600, 1540465200, 1540468800, 1540472400, 
    1540476000, 1540479600, 1540483200, 1540486800, 1540490400, 1540494000, 
    1540497600, 1540501200, 1540504800, 1540508400, 1540512000, 1540515600, 
    1540519200, 1540522800, 1540526400, 1540530000, 1540533600, 1540537200, 
    1540540800, 1540544400, 1540548000, 1540551600, 1540555200, 1540558800, 
    1540562400, 1540566000, 1540569600, 1540573200, 1540576800, 1540580400, 
    1540584000, 1540587600, 1540591200, 1540594800, 1540598400, 1540602000, 
    1540605600, 1540609200, 1540612800, 1540616400, 1540620000, 1540623600, 
    1540627200, 1540630800, 1540634400, 1540638000, 1540641600, 1540645200, 
    1540648800, 1540652400, 1540656000, 1540659600, 1540663200, 1540666800, 
    1540670400, 1540674000, 1540677600, 1540681200, 1540684800, 1540688400, 
    1540692000, 1540695600, 1540699200, 1540702800, 1540706400, 1540710000, 
    1540713600, 1540717200, 1540720800, 1540724400, 1540728000, 1540731600, 
    1540735200, 1540738800, 1540742400, 1540746000, 1540749600, 1540753200, 
    1540756800, 1540760400, 1540764000, 1540767600, 1540771200, 1540774800, 
    1540778400, 1540782000, 1540785600, 1540789200, 1540792800, 1540796400, 
    1540800000, 1540803600, 1540807200, 1540810800, 1540814400, 1540818000, 
    1540821600, 1540825200, 1540828800, 1540832400, 1540836000, 1540839600, 
    1540843200, 1540846800, 1540850400, 1540854000, 1540857600, 1540861200, 
    1540864800, 1540868400, 1540872000, 1540875600, 1540879200, 1540882800, 
    1540886400, 1540890000, 1540893600, 1540897200, 1540900800, 1540904400, 
    1540908000, 1540911600, 1540915200, 1540918800, 1540922400, 1540926000, 
    1540929600, 1540933200, 1540936800, 1540940400, 1540944000, 1540947600, 
    1540951200, 1540954800, 1540958400, 1540962000, 1540965600, 1540969200, 
    1540972800, 1540976400, 1540980000, 1540983600, 1540987200, 1540990800, 
    1540994400, 1540998000, 1541001600, 1541005200, 1541008800, 1541012400, 
    1541016000, 1541019600, 1541023200, 1541026800, 1541030400, 1541034000, 
    1541037600, 1541041200, 1541044800, 1541048400, 1541052000, 1541055600, 
    1541059200, 1541062800, 1541066400, 1541070000, 1541073600, 1541077200, 
    1541080800, 1541084400, 1541088000, 1541091600, 1541095200, 1541098800, 
    1541102400, 1541106000, 1541109600, 1541113200, 1541116800, 1541120400, 
    1541124000, 1541127600, 1541131200, 1541134800, 1541138400, 1541142000, 
    1541145600, 1541149200, 1541152800, 1541156400, 1541160000, 1541163600, 
    1541167200, 1541170800, 1541174400, 1541178000, 1541181600, 1541185200, 
    1541188800, 1541192400, 1541196000, 1541199600, 1541203200, 1541206800, 
    1541210400, 1541214000, 1541217600, 1541221200, 1541224800, 1541228400, 
    1541232000, 1541235600, 1541239200, 1541242800, 1541246400, 1541250000, 
    1541253600, 1541257200, 1541260800, 1541264400, 1541268000, 1541271600, 
    1541275200, 1541278800, 1541282400, 1541286000, 1541289600, 1541293200, 
    1541296800, 1541300400, 1541304000, 1541307600, 1541311200, 1541314800, 
    1541318400, 1541322000, 1541325600, 1541329200, 1541332800, 1541336400, 
    1541340000, 1541343600, 1541347200, 1541350800, 1541354400, 1541358000, 
    1541361600, 1541365200, 1541368800, 1541372400, 1541376000, 1541379600, 
    1541383200, 1541386800, 1541390400, 1541394000, 1541397600, 1541401200, 
    1541404800, 1541408400, 1541412000, 1541415600, 1541419200, 1541422800, 
    1541426400, 1541430000, 1541433600, 1541437200, 1541440800, 1541444400, 
    1541448000, 1541451600, 1541455200, 1541458800, 1541462400, 1541466000, 
    1541469600, 1541473200, 1541476800, 1541480400, 1541484000, 1541487600, 
    1541491200, 1541494800, 1541498400, 1541502000, 1541505600, 1541509200, 
    1541512800, 1541516400, 1541520000, 1541523600, 1541527200, 1541530800, 
    1541534400, 1541538000, 1541541600, 1541545200, 1541548800, 1541552400, 
    1541556000, 1541559600, 1541563200, 1541566800, 1541570400, 1541574000, 
    1541577600, 1541581200, 1541584800, 1541588400, 1541592000, 1541595600, 
    1541599200, 1541602800, 1541606400, 1541610000, 1541613600, 1541617200, 
    1541620800, 1541624400, 1541628000, 1541631600, 1541635200, 1541638800, 
    1541642400, 1541646000, 1541649600, 1541653200, 1541656800, 1541660400, 
    1541664000, 1541667600, 1541671200, 1541674800, 1541678400, 1541682000, 
    1541685600, 1541689200, 1541692800, 1541696400, 1541700000, 1541703600, 
    1541707200, 1541710800, 1541714400, 1541718000, 1541721600, 1541725200, 
    1541728800, 1541732400, 1541736000, 1541739600, 1541743200, 1541746800, 
    1541750400, 1541754000, 1541757600, 1541761200, 1541764800, 1541768400, 
    1541772000, 1541775600, 1541779200, 1541782800, 1541786400, 1541790000, 
    1541793600, 1541797200, 1541800800, 1541804400, 1541808000, 1541811600, 
    1541815200, 1541818800, 1541822400, 1541826000, 1541829600, 1541833200, 
    1541836800, 1541840400, 1541844000, 1541847600, 1541851200, 1541854800, 
    1541858400, 1541862000, 1541865600, 1541869200, 1541872800, 1541876400, 
    1541880000, 1541883600, 1541887200, 1541890800, 1541894400, 1541898000, 
    1541901600, 1541905200, 1541908800, 1541912400, 1541916000, 1541919600, 
    1541923200, 1541926800, 1541930400, 1541934000, 1541937600, 1541941200, 
    1541944800, 1541948400, 1541952000, 1541955600, 1541959200, 1541962800, 
    1541966400, 1541970000, 1541973600, 1541977200, 1541980800, 1541984400, 
    1541988000, 1541991600, 1541995200, 1541998800, 1542002400, 1542006000, 
    1542009600, 1542013200, 1542016800, 1542020400, 1542024000, 1542027600, 
    1542031200, 1542034800, 1542038400, 1542042000, 1542045600, 1542049200, 
    1542052800, 1542056400, 1542060000, 1542063600, 1542067200, 1542070800, 
    1542074400, 1542078000, 1542081600, 1542085200, 1542088800, 1542092400, 
    1542096000, 1542099600, 1542103200, 1542106800, 1542110400, 1542114000, 
    1542117600, 1542121200, 1542124800, 1542128400, 1542132000, 1542135600, 
    1542139200, 1542142800, 1542146400, 1542150000, 1542153600, 1542157200, 
    1542160800, 1542164400, 1542168000, 1542171600, 1542175200, 1542178800, 
    1542182400, 1542186000, 1542189600, 1542193200, 1542196800, 1542200400, 
    1542204000, 1542207600, 1542211200, 1542214800, 1542218400, 1542222000, 
    1542225600, 1542229200, 1542232800, 1542236400, 1542240000, 1542243600, 
    1542247200, 1542250800, 1542254400, 1542258000, 1542261600, 1542265200, 
    1542268800, 1542272400, 1542276000, 1542279600, 1542283200, 1542286800, 
    1542290400, 1542294000, 1542297600, 1542301200, 1542304800, 1542308400, 
    1542312000, 1542315600, 1542319200, 1542322800, 1542326400, 1542330000, 
    1542333600, 1542337200, 1542340800, 1542344400, 1542348000, 1542351600, 
    1542355200, 1542358800, 1542362400, 1542366000, 1542369600, 1542373200, 
    1542376800, 1542380400, 1542384000, 1542387600, 1542391200, 1542394800, 
    1542398400, 1542402000, 1542405600, 1542409200, 1542412800, 1542416400, 
    1542420000, 1542423600, 1542427200, 1542430800, 1542434400, 1542438000, 
    1542441600, 1542445200, 1542448800, 1542452400, 1542456000, 1542459600, 
    1542463200, 1542466800, 1542470400, 1542474000, 1542477600, 1542481200, 
    1542484800, 1542488400, 1542492000, 1542495600, 1542499200, 1542502800, 
    1542506400, 1542510000, 1542513600, 1542517200, 1542520800, 1542524400, 
    1542528000, 1542531600, 1542535200, 1542538800, 1542542400, 1542546000, 
    1542549600, 1542553200, 1542556800, 1542560400, 1542564000, 1542567600, 
    1542571200, 1542574800, 1542578400, 1542582000, 1542585600, 1542589200, 
    1542592800, 1542596400, 1542600000, 1542603600, 1542607200, 1542610800, 
    1542614400, 1542618000, 1542621600, 1542625200, 1542628800, 1542632400, 
    1542636000, 1542639600, 1542643200, 1542646800, 1542650400, 1542654000, 
    1542657600, 1542661200, 1542664800, 1542668400, 1542672000, 1542675600, 
    1542679200, 1542682800, 1542686400, 1542690000, 1542693600, 1542697200, 
    1542700800, 1542704400, 1542708000, 1542711600, 1542715200, 1542718800, 
    1542722400, 1542726000, 1542729600, 1542733200, 1542736800, 1542740400, 
    1542744000, 1542747600, 1542751200, 1542754800, 1542758400, 1542762000, 
    1542765600, 1542769200, 1542772800, 1542776400, 1542780000, 1542783600, 
    1542787200, 1542790800, 1542794400, 1542798000, 1542801600, 1542805200, 
    1542808800, 1542812400, 1542816000, 1542819600, 1542823200, 1542826800, 
    1542830400, 1542834000, 1542837600, 1542841200, 1542844800, 1542848400, 
    1542852000, 1542855600, 1542859200, 1542862800, 1542866400, 1542870000, 
    1542873600, 1542877200, 1542880800, 1542884400, 1542888000, 1542891600, 
    1542895200, 1542898800, 1542902400, 1542906000, 1542909600, 1542913200, 
    1542916800, 1542920400, 1542924000, 1542927600, 1542931200, 1542934800, 
    1542938400, 1542942000, 1542945600, 1542949200, 1542952800, 1542956400, 
    1542960000, 1542963600, 1542967200, 1542970800, 1542974400, 1542978000, 
    1542981600, 1542985200, 1542988800, 1542992400, 1542996000, 1542999600, 
    1543003200, 1543006800, 1543010400, 1543014000, 1543017600, 1543021200, 
    1543024800, 1543028400, 1543032000, 1543035600, 1543039200, 1543042800, 
    1543046400, 1543050000, 1543053600, 1543057200, 1543060800, 1543064400, 
    1543068000, 1543071600, 1543075200, 1543078800, 1543082400, 1543086000, 
    1543089600, 1543093200, 1543096800, 1543100400, 1543104000, 1543107600, 
    1543111200, 1543114800, 1543118400, 1543122000, 1543125600, 1543129200, 
    1543132800, 1543136400, 1543140000, 1543143600, 1543147200, 1543150800, 
    1543154400, 1543158000, 1543161600, 1543165200, 1543168800, 1543172400, 
    1543176000, 1543179600, 1543183200, 1543186800, 1543190400, 1543194000, 
    1543197600, 1543201200, 1543204800, 1543208400, 1543212000, 1543215600, 
    1543219200, 1543222800, 1543226400, 1543230000, 1543233600, 1543237200, 
    1543240800, 1543244400, 1543248000, 1543251600, 1543255200, 1543258800, 
    1543262400, 1543266000, 1543269600, 1543273200, 1543276800, 1543280400, 
    1543284000, 1543287600, 1543291200, 1543294800, 1543298400, 1543302000, 
    1543305600, 1543309200, 1543312800, 1543316400, 1543320000, 1543323600, 
    1543327200, 1543330800, 1543334400, 1543338000, 1543341600, 1543345200, 
    1543348800, 1543352400, 1543356000, 1543359600, 1543363200, 1543366800, 
    1543370400, 1543374000, 1543377600, 1543381200, 1543384800, 1543388400, 
    1543392000, 1543395600, 1543399200, 1543402800, 1543406400, 1543410000, 
    1543413600, 1543417200, 1543420800, 1543424400, 1543428000, 1543431600, 
    1543435200, 1543438800, 1543442400, 1543446000, 1543449600, 1543453200, 
    1543456800, 1543460400, 1543464000, 1543467600, 1543471200, 1543474800, 
    1543478400, 1543482000, 1543485600, 1543489200, 1543492800, 1543496400, 
    1543500000, 1543503600, 1543507200, 1543510800, 1543514400, 1543518000, 
    1543521600, 1543525200, 1543528800, 1543532400, 1543536000, 1543539600, 
    1543543200, 1543546800, 1543550400, 1543554000, 1543557600, 1543561200, 
    1543564800, 1543568400, 1543572000, 1543575600, 1543579200, 1543582800, 
    1543586400, 1543590000, 1543593600, 1543597200, 1543600800, 1543604400, 
    1543608000, 1543611600, 1543615200, 1543618800, 1543622400, 1543626000, 
    1543629600, 1543633200, 1543636800, 1543640400, 1543644000, 1543647600, 
    1543651200, 1543654800, 1543658400, 1543662000, 1543665600, 1543669200, 
    1543672800, 1543676400, 1543680000, 1543683600, 1543687200, 1543690800, 
    1543694400, 1543698000, 1543701600, 1543705200, 1543708800, 1543712400, 
    1543716000, 1543719600, 1543723200, 1543726800, 1543730400, 1543734000, 
    1543737600, 1543741200, 1543744800, 1543748400, 1543752000, 1543755600, 
    1543759200, 1543762800, 1543766400, 1543770000, 1543773600, 1543777200, 
    1543780800, 1543784400, 1543788000, 1543791600, 1543795200, 1543798800, 
    1543802400, 1543806000, 1543809600, 1543813200, 1543816800, 1543820400, 
    1543824000, 1543827600, 1543831200, 1543834800, 1543838400, 1543842000, 
    1543845600, 1543849200, 1543852800, 1543856400, 1543860000, 1543863600, 
    1543867200, 1543870800, 1543874400, 1543878000, 1543881600, 1543885200, 
    1543888800, 1543892400, 1543896000, 1543899600, 1543903200, 1543906800, 
    1543910400, 1543914000, 1543917600, 1543921200, 1543924800, 1543928400, 
    1543932000, 1543935600, 1543939200, 1543942800, 1543946400, 1543950000, 
    1543953600, 1543957200, 1543960800, 1543964400, 1543968000, 1543971600, 
    1543975200, 1543978800, 1543982400, 1543986000, 1543989600, 1543993200, 
    1543996800, 1544000400, 1544004000, 1544007600, 1544011200, 1544014800, 
    1544018400, 1544022000, 1544025600, 1544029200, 1544032800, 1544036400, 
    1544040000, 1544043600, 1544047200, 1544050800, 1544054400, 1544058000, 
    1544061600, 1544065200, 1544068800, 1544072400, 1544076000, 1544079600, 
    1544083200, 1544086800, 1544090400, 1544094000, 1544097600, 1544101200, 
    1544104800, 1544108400, 1544112000, 1544115600, 1544119200, 1544122800, 
    1544126400, 1544130000, 1544133600, 1544137200, 1544140800, 1544144400, 
    1544148000, 1544151600, 1544155200, 1544158800, 1544162400, 1544166000, 
    1544169600, 1544173200, 1544176800, 1544180400, 1544184000, 1544187600, 
    1544191200, 1544194800, 1544198400, 1544202000, 1544205600, 1544209200, 
    1544212800, 1544216400, 1544220000, 1544223600, 1544227200, 1544230800, 
    1544234400, 1544238000, 1544241600, 1544245200, 1544248800, 1544252400, 
    1544256000, 1544259600, 1544263200, 1544266800, 1544270400, 1544274000, 
    1544277600, 1544281200, 1544284800, 1544288400, 1544292000, 1544295600, 
    1544299200, 1544302800, 1544306400, 1544310000, 1544313600, 1544317200, 
    1544320800, 1544324400, 1544328000, 1544331600, 1544335200, 1544338800, 
    1544342400, 1544346000, 1544349600, 1544353200, 1544356800, 1544360400, 
    1544364000, 1544367600, 1544371200, 1544374800, 1544378400, 1544382000, 
    1544385600, 1544389200, 1544392800, 1544396400, 1544400000, 1544403600, 
    1544407200, 1544410800, 1544414400, 1544418000, 1544421600, 1544425200, 
    1544428800, 1544432400, 1544436000, 1544439600, 1544443200, 1544446800, 
    1544450400, 1544454000, 1544457600, 1544461200, 1544464800, 1544468400, 
    1544472000, 1544475600, 1544479200, 1544482800, 1544486400, 1544490000, 
    1544493600, 1544497200, 1544500800, 1544504400, 1544508000, 1544511600, 
    1544515200, 1544518800, 1544522400, 1544526000, 1544529600, 1544533200, 
    1544536800, 1544540400, 1544544000, 1544547600, 1544551200, 1544554800, 
    1544558400, 1544562000, 1544565600, 1544569200, 1544572800, 1544576400, 
    1544580000, 1544583600, 1544587200, 1544590800, 1544594400, 1544598000, 
    1544601600, 1544605200, 1544608800, 1544612400, 1544616000, 1544619600, 
    1544623200, 1544626800, 1544630400, 1544634000, 1544637600, 1544641200, 
    1544644800, 1544648400, 1544652000, 1544655600, 1544659200, 1544662800, 
    1544666400, 1544670000, 1544673600, 1544677200, 1544680800, 1544684400, 
    1544688000, 1544691600, 1544695200, 1544698800, 1544702400, 1544706000, 
    1544709600, 1544713200, 1544716800, 1544720400, 1544724000, 1544727600, 
    1544731200, 1544734800, 1544738400, 1544742000, 1544745600, 1544749200, 
    1544752800, 1544756400, 1544760000, 1544763600, 1544767200, 1544770800, 
    1544774400, 1544778000, 1544781600, 1544785200, 1544788800, 1544792400, 
    1544796000, 1544799600, 1544803200, 1544806800, 1544810400, 1544814000, 
    1544817600, 1544821200, 1544824800, 1544828400, 1544832000, 1544835600, 
    1544839200, 1544842800, 1544846400, 1544850000, 1544853600, 1544857200, 
    1544860800, 1544864400, 1544868000, 1544871600, 1544875200, 1544878800, 
    1544882400, 1544886000, 1544889600, 1544893200, 1544896800, 1544900400, 
    1544904000, 1544907600, 1544911200, 1544914800, 1544918400, 1544922000, 
    1544925600, 1544929200, 1544932800, 1544936400, 1544940000, 1544943600, 
    1544947200, 1544950800, 1544954400, 1544958000, 1544961600, 1544965200, 
    1544968800, 1544972400, 1544976000, 1544979600, 1544983200, 1544986800, 
    1544990400, 1544994000, 1544997600, 1545001200, 1545004800, 1545008400, 
    1545012000, 1545015600, 1545019200, 1545022800, 1545026400, 1545030000, 
    1545033600, 1545037200, 1545040800, 1545044400, 1545048000, 1545051600, 
    1545055200, 1545058800, 1545062400, 1545066000, 1545069600, 1545073200, 
    1545076800, 1545080400, 1545084000, 1545087600, 1545091200, 1545094800, 
    1545098400, 1545102000, 1545105600, 1545109200, 1545112800, 1545116400, 
    1545120000, 1545123600, 1545127200, 1545130800, 1545134400, 1545138000, 
    1545141600, 1545145200, 1545148800, 1545152400, 1545156000, 1545159600, 
    1545163200, 1545166800, 1545170400, 1545174000, 1545177600, 1545181200, 
    1545184800, 1545188400, 1545192000, 1545195600, 1545199200, 1545202800, 
    1545206400, 1545210000, 1545213600, 1545217200, 1545220800, 1545224400, 
    1545228000, 1545231600, 1545235200, 1545238800, 1545242400, 1545246000, 
    1545249600, 1545253200, 1545256800, 1545260400, 1545264000, 1545267600, 
    1545271200, 1545274800, 1545278400, 1545282000, 1545285600, 1545289200, 
    1545292800, 1545296400, 1545300000, 1545303600, 1545307200, 1545310800, 
    1545314400, 1545318000, 1545321600, 1545325200, 1545328800, 1545332400, 
    1545336000, 1545339600, 1545343200, 1545346800, 1545350400, 1545354000, 
    1545357600, 1545361200, 1545364800, 1545368400, 1545372000, 1545375600, 
    1545379200, 1545382800, 1545386400, 1545390000, 1545393600, 1545397200, 
    1545400800, 1545404400, 1545408000, 1545411600, 1545415200, 1545418800, 
    1545422400, 1545426000, 1545429600, 1545433200, 1545436800, 1545440400, 
    1545444000, 1545447600, 1545451200, 1545454800, 1545458400, 1545462000, 
    1545465600, 1545469200, 1545472800, 1545476400, 1545480000, 1545483600, 
    1545487200, 1545490800, 1545494400, 1545498000, 1545501600, 1545505200, 
    1545508800, 1545512400, 1545516000, 1545519600, 1545523200, 1545526800, 
    1545530400, 1545534000, 1545537600, 1545541200, 1545544800, 1545548400, 
    1545552000, 1545555600, 1545559200, 1545562800, 1545566400, 1545570000, 
    1545573600, 1545577200, 1545580800, 1545584400, 1545588000, 1545591600, 
    1545595200, 1545598800, 1545602400, 1545606000, 1545609600, 1545613200, 
    1545616800, 1545620400, 1545624000, 1545627600, 1545631200, 1545634800, 
    1545638400, 1545642000, 1545645600, 1545649200, 1545652800, 1545656400, 
    1545660000, 1545663600, 1545667200, 1545670800, 1545674400, 1545678000, 
    1545681600, 1545685200, 1545688800, 1545692400, 1545696000, 1545699600, 
    1545703200, 1545706800, 1545710400, 1545714000, 1545717600, 1545721200, 
    1545724800, 1545728400, 1545732000, 1545735600, 1545739200, 1545742800, 
    1545746400, 1545750000, 1545753600, 1545757200, 1545760800, 1545764400, 
    1545768000, 1545771600, 1545775200, 1545778800, 1545782400, 1545786000, 
    1545789600, 1545793200, 1545796800, 1545800400, 1545804000, 1545807600, 
    1545811200, 1545814800, 1545818400, 1545822000, 1545825600, 1545829200, 
    1545832800, 1545836400, 1545840000, 1545843600, 1545847200, 1545850800, 
    1545854400, 1545858000, 1545861600, 1545865200, 1545868800, 1545872400, 
    1545876000, 1545879600, 1545883200, 1545886800, 1545890400, 1545894000, 
    1545897600, 1545901200, 1545904800, 1545908400, 1545912000, 1545915600, 
    1545919200, 1545922800, 1545926400, 1545930000, 1545933600, 1545937200, 
    1545940800, 1545944400, 1545948000, 1545951600, 1545955200, 1545958800, 
    1545962400, 1545966000, 1545969600, 1545973200, 1545976800, 1545980400, 
    1545984000, 1545987600, 1545991200, 1545994800, 1545998400, 1546002000, 
    1546005600, 1546009200, 1546012800, 1546016400, 1546020000, 1546023600, 
    1546027200, 1546030800, 1546034400, 1546038000, 1546041600, 1546045200, 
    1546048800, 1546052400, 1546056000, 1546059600, 1546063200, 1546066800, 
    1546070400, 1546074000, 1546077600, 1546081200, 1546084800, 1546088400, 
    1546092000, 1546095600, 1546099200, 1546102800, 1546106400, 1546110000, 
    1546113600, 1546117200, 1546120800, 1546124400, 1546128000, 1546131600, 
    1546135200, 1546138800, 1546142400, 1546146000, 1546149600, 1546153200, 
    1546156800, 1546160400, 1546164000, 1546167600, 1546171200, 1546174800, 
    1546178400, 1546182000, 1546185600, 1546189200, 1546192800, 1546196400, 
    1546200000, 1546203600, 1546207200, 1546210800, 1546214400, 1546218000, 
    1546221600, 1546225200, 1546228800, 1546232400, 1546236000, 1546239600, 
    1546243200, 1546246800, 1546250400, 1546254000, 1546257600, 1546261200, 
    1546264800, 1546268400, 1546272000, 1546275600, 1546279200, 1546282800, 
    1546286400, 1546290000, 1546293600, 1546297200, 1546300800, 1546304400, 
    1546308000, 1546311600, 1546315200, 1546318800, 1546322400, 1546326000, 
    1546329600, 1546333200, 1546336800, 1546340400, 1546344000, 1546347600, 
    1546351200, 1546354800, 1546358400, 1546362000, 1546365600, 1546369200, 
    1546372800, 1546376400, 1546380000, 1546383600, 1546387200, 1546390800, 
    1546394400, 1546398000, 1546401600, 1546405200, 1546408800, 1546412400, 
    1546416000, 1546419600, 1546423200, 1546426800, 1546430400, 1546434000, 
    1546437600, 1546441200, 1546444800, 1546448400, 1546452000, 1546455600, 
    1546459200, 1546462800, 1546466400, 1546470000, 1546473600, 1546477200, 
    1546480800, 1546484400, 1546488000, 1546491600, 1546495200, 1546498800, 
    1546502400, 1546506000, 1546509600, 1546513200, 1546516800, 1546520400, 
    1546524000, 1546527600, 1546531200, 1546534800, 1546538400, 1546542000, 
    1546545600, 1546549200, 1546552800, 1546556400, 1546560000, 1546563600, 
    1546567200, 1546570800, 1546574400, 1546578000, 1546581600, 1546585200, 
    1546588800, 1546592400, 1546596000, 1546599600, 1546603200, 1546606800, 
    1546610400, 1546614000, 1546617600, 1546621200, 1546624800, 1546628400, 
    1546632000, 1546635600, 1546639200, 1546642800, 1546646400, 1546650000, 
    1546653600, 1546657200, 1546660800, 1546664400, 1546668000, 1546671600, 
    1546675200, 1546678800, 1546682400, 1546686000, 1546689600, 1546693200, 
    1546696800, 1546700400, 1546704000, 1546707600, 1546711200, 1546714800, 
    1546718400, 1546722000, 1546725600, 1546729200, 1546732800, 1546736400, 
    1546740000, 1546743600, 1546747200, 1546750800, 1546754400, 1546758000, 
    1546761600, 1546765200, 1546768800, 1546772400, 1546776000, 1546779600, 
    1546783200, 1546786800, 1546790400, 1546794000, 1546797600, 1546801200, 
    1546804800, 1546808400, 1546812000, 1546815600, 1546819200, 1546822800, 
    1546826400, 1546830000, 1546833600, 1546837200, 1546840800, 1546844400, 
    1546848000, 1546851600, 1546855200, 1546858800, 1546862400, 1546866000, 
    1546869600, 1546873200, 1546876800, 1546880400, 1546884000, 1546887600, 
    1546891200, 1546894800, 1546898400, 1546902000, 1546905600, 1546909200, 
    1546912800, 1546916400, 1546920000, 1546923600, 1546927200, 1546930800, 
    1546934400, 1546938000, 1546941600, 1546945200, 1546948800, 1546952400, 
    1546956000, 1546959600, 1546963200, 1546966800, 1546970400, 1546974000, 
    1546977600, 1546981200, 1546984800, 1546988400, 1546992000, 1546995600, 
    1546999200, 1547002800, 1547006400, 1547010000, 1547013600, 1547017200, 
    1547020800, 1547024400, 1547028000, 1547031600, 1547035200, 1547038800, 
    1547042400, 1547046000, 1547049600, 1547053200, 1547056800, 1547060400, 
    1547064000, 1547067600, 1547071200, 1547074800, 1547078400, 1547082000, 
    1547085600, 1547089200, 1547092800, 1547096400, 1547100000, 1547103600, 
    1547107200, 1547110800, 1547114400, 1547118000, 1547121600, 1547125200, 
    1547128800, 1547132400, 1547136000, 1547139600, 1547143200, 1547146800, 
    1547150400, 1547154000, 1547157600, 1547161200, 1547164800, 1547168400, 
    1547172000, 1547175600, 1547179200, 1547182800, 1547186400, 1547190000, 
    1547193600, 1547197200, 1547200800, 1547204400, 1547208000, 1547211600, 
    1547215200, 1547218800, 1547222400, 1547226000, 1547229600, 1547233200, 
    1547236800, 1547240400, 1547244000, 1547247600, 1547251200, 1547254800, 
    1547258400, 1547262000, 1547265600, 1547269200, 1547272800, 1547276400, 
    1547280000, 1547283600, 1547287200, 1547290800, 1547294400, 1547298000, 
    1547301600, 1547305200, 1547308800, 1547312400, 1547316000, 1547319600, 
    1547323200, 1547326800, 1547330400, 1547334000, 1547337600, 1547341200, 
    1547344800, 1547348400, 1547352000, 1547355600, 1547359200, 1547362800, 
    1547366400, 1547370000, 1547373600, 1547377200, 1547380800, 1547384400, 
    1547388000, 1547391600, 1547395200, 1547398800, 1547402400, 1547406000, 
    1547409600, 1547413200, 1547416800, 1547420400, 1547424000, 1547427600, 
    1547431200, 1547434800, 1547438400, 1547442000, 1547445600, 1547449200, 
    1547452800, 1547456400, 1547460000, 1547463600, 1547467200, 1547470800, 
    1547474400, 1547478000, 1547481600, 1547485200, 1547488800, 1547492400, 
    1547496000, 1547499600, 1547503200, 1547506800, 1547510400, 1547514000, 
    1547517600, 1547521200, 1547524800, 1547528400, 1547532000, 1547535600, 
    1547539200, 1547542800, 1547546400, 1547550000, 1547553600, 1547557200, 
    1547560800, 1547564400, 1547568000, 1547571600, 1547575200, 1547578800, 
    1547582400, 1547586000, 1547589600, 1547593200, 1547596800, 1547600400, 
    1547604000, 1547607600, 1547611200, 1547614800, 1547618400, 1547622000, 
    1547625600, 1547629200, 1547632800, 1547636400, 1547640000, 1547643600, 
    1547647200, 1547650800, 1547654400, 1547658000, 1547661600, 1547665200, 
    1547668800, 1547672400, 1547676000, 1547679600, 1547683200, 1547686800, 
    1547690400, 1547694000, 1547697600, 1547701200, 1547704800, 1547708400, 
    1547712000, 1547715600, 1547719200, 1547722800, 1547726400, 1547730000, 
    1547733600, 1547737200, 1547740800, 1547744400, 1547748000, 1547751600, 
    1547755200, 1547758800, 1547762400, 1547766000, 1547769600, 1547773200, 
    1547776800, 1547780400, 1547784000, 1547787600, 1547791200, 1547794800, 
    1547798400, 1547802000, 1547805600, 1547809200, 1547812800, 1547816400, 
    1547820000, 1547823600, 1547827200, 1547830800, 1547834400, 1547838000, 
    1547841600, 1547845200, 1547848800, 1547852400, 1547856000, 1547859600, 
    1547863200, 1547866800, 1547870400, 1547874000, 1547877600, 1547881200, 
    1547884800, 1547888400, 1547892000, 1547895600, 1547899200, 1547902800, 
    1547906400, 1547910000, 1547913600, 1547917200, 1547920800, 1547924400, 
    1547928000, 1547931600, 1547935200, 1547938800, 1547942400, 1547946000, 
    1547949600, 1547953200, 1547956800, 1547960400, 1547964000, 1547967600, 
    1547971200, 1547974800, 1547978400, 1547982000, 1547985600, 1547989200, 
    1547992800, 1547996400, 1548000000, 1548003600, 1548007200, 1548010800, 
    1548014400, 1548018000, 1548021600, 1548025200, 1548028800, 1548032400, 
    1548036000, 1548039600, 1548043200, 1548046800, 1548050400, 1548054000, 
    1548057600, 1548061200, 1548064800, 1548068400, 1548072000, 1548075600, 
    1548079200, 1548082800, 1548086400, 1548090000, 1548093600, 1548097200, 
    1548100800, 1548104400, 1548108000, 1548111600, 1548115200, 1548118800, 
    1548122400, 1548126000, 1548129600, 1548133200, 1548136800, 1548140400, 
    1548144000, 1548147600, 1548151200, 1548154800, 1548158400, 1548162000, 
    1548165600, 1548169200, 1548172800, 1548176400, 1548180000, 1548183600, 
    1548187200, 1548190800, 1548194400, 1548198000, 1548201600, 1548205200, 
    1548208800, 1548212400, 1548216000, 1548219600, 1548223200, 1548226800, 
    1548230400, 1548234000, 1548237600, 1548241200, 1548244800, 1548248400, 
    1548252000, 1548255600, 1548259200, 1548262800, 1548266400, 1548270000, 
    1548273600, 1548277200, 1548280800, 1548284400, 1548288000, 1548291600, 
    1548295200, 1548298800, 1548302400, 1548306000, 1548309600, 1548313200, 
    1548316800, 1548320400, 1548324000, 1548327600, 1548331200, 1548334800, 
    1548338400, 1548342000, 1548345600, 1548349200, 1548352800, 1548356400, 
    1548360000, 1548363600, 1548367200, 1548370800, 1548374400, 1548378000, 
    1548381600, 1548385200, 1548388800, 1548392400, 1548396000, 1548399600, 
    1548403200, 1548406800, 1548410400, 1548414000, 1548417600, 1548421200, 
    1548424800, 1548428400, 1548432000, 1548435600, 1548439200, 1548442800, 
    1548446400, 1548450000, 1548453600, 1548457200, 1548460800, 1548464400, 
    1548468000, 1548471600, 1548475200, 1548478800, 1548482400, 1548486000, 
    1548489600, 1548493200, 1548496800, 1548500400, 1548504000, 1548507600, 
    1548511200, 1548514800, 1548518400, 1548522000, 1548525600, 1548529200, 
    1548532800, 1548536400, 1548540000, 1548543600, 1548547200, 1548550800, 
    1548554400, 1548558000, 1548561600, 1548565200, 1548568800, 1548572400, 
    1548576000, 1548579600, 1548583200, 1548586800, 1548590400, 1548594000, 
    1548597600, 1548601200, 1548604800, 1548608400, 1548612000, 1548615600, 
    1548619200, 1548622800, 1548626400, 1548630000, 1548633600, 1548637200, 
    1548640800, 1548644400, 1548648000, 1548651600, 1548655200, 1548658800, 
    1548662400, 1548666000, 1548669600, 1548673200, 1548676800, 1548680400, 
    1548684000, 1548687600, 1548691200, 1548694800, 1548698400, 1548702000, 
    1548705600, 1548709200, 1548712800, 1548716400, 1548720000, 1548723600, 
    1548727200, 1548730800, 1548734400, 1548738000, 1548741600, 1548745200, 
    1548748800, 1548752400, 1548756000, 1548759600, 1548763200, 1548766800, 
    1548770400, 1548774000, 1548777600, 1548781200, 1548784800, 1548788400, 
    1548792000, 1548795600, 1548799200, 1548802800, 1548806400, 1548810000, 
    1548813600, 1548817200, 1548820800, 1548824400, 1548828000, 1548831600, 
    1548835200, 1548838800, 1548842400, 1548846000, 1548849600, 1548853200, 
    1548856800, 1548860400, 1548864000, 1548867600, 1548871200, 1548874800, 
    1548878400, 1548882000, 1548885600, 1548889200, 1548892800, 1548896400, 
    1548900000, 1548903600, 1548907200, 1548910800, 1548914400, 1548918000, 
    1548921600, 1548925200, 1548928800, 1548932400, 1548936000, 1548939600, 
    1548943200, 1548946800, 1548950400, 1548954000, 1548957600, 1548961200, 
    1548964800, 1548968400, 1548972000, 1548975600, 1548979200, 1548982800, 
    1548986400, 1548990000, 1548993600, 1548997200, 1549000800, 1549004400, 
    1549008000, 1549011600, 1549015200, 1549018800, 1549022400, 1549026000, 
    1549029600, 1549033200, 1549036800, 1549040400, 1549044000, 1549047600, 
    1549051200, 1549054800, 1549058400, 1549062000, 1549065600, 1549069200, 
    1549072800, 1549076400, 1549080000, 1549083600, 1549087200, 1549090800, 
    1549094400, 1549098000, 1549101600, 1549105200, 1549108800, 1549112400, 
    1549116000, 1549119600, 1549123200, 1549126800, 1549130400, 1549134000, 
    1549137600, 1549141200, 1549144800, 1549148400, 1549152000, 1549155600, 
    1549159200, 1549162800, 1549166400, 1549170000, 1549173600, 1549177200, 
    1549180800, 1549184400, 1549188000, 1549191600, 1549195200, 1549198800, 
    1549202400, 1549206000, 1549209600, 1549213200, 1549216800, 1549220400, 
    1549224000, 1549227600, 1549231200, 1549234800, 1549238400, 1549242000, 
    1549245600, 1549249200, 1549252800, 1549256400, 1549260000, 1549263600, 
    1549267200, 1549270800, 1549274400, 1549278000, 1549281600, 1549285200, 
    1549288800, 1549292400, 1549296000, 1549299600, 1549303200, 1549306800, 
    1549310400, 1549314000, 1549317600, 1549321200, 1549324800, 1549328400, 
    1549332000, 1549335600, 1549339200, 1549342800, 1549346400, 1549350000, 
    1549353600, 1549357200, 1549360800, 1549364400, 1549368000, 1549371600, 
    1549375200, 1549378800, 1549382400, 1549386000, 1549389600, 1549393200, 
    1549396800, 1549400400, 1549404000, 1549407600, 1549411200, 1549414800, 
    1549418400, 1549422000, 1549425600, 1549429200, 1549432800, 1549436400, 
    1549440000, 1549443600, 1549447200, 1549450800, 1549454400, 1549458000, 
    1549461600, 1549465200, 1549468800, 1549472400, 1549476000, 1549479600, 
    1549483200, 1549486800, 1549490400, 1549494000, 1549497600, 1549501200, 
    1549504800, 1549508400, 1549512000, 1549515600, 1549519200, 1549522800, 
    1549526400, 1549530000, 1549533600, 1549537200, 1549540800, 1549544400, 
    1549548000, 1549551600, 1549555200, 1549558800, 1549562400, 1549566000, 
    1549569600, 1549573200, 1549576800, 1549580400, 1549584000, 1549587600, 
    1549591200, 1549594800, 1549598400, 1549602000, 1549605600, 1549609200, 
    1549612800, 1549616400, 1549620000, 1549623600, 1549627200, 1549630800, 
    1549634400, 1549638000, 1549641600, 1549645200, 1549648800, 1549652400, 
    1549656000, 1549659600, 1549663200, 1549666800, 1549670400, 1549674000, 
    1549677600, 1549681200, 1549684800, 1549688400, 1549692000, 1549695600, 
    1549699200, 1549702800, 1549706400, 1549710000, 1549713600, 1549717200, 
    1549720800, 1549724400, 1549728000, 1549731600, 1549735200, 1549738800, 
    1549742400, 1549746000, 1549749600, 1549753200, 1549756800, 1549760400, 
    1549764000, 1549767600, 1549771200, 1549774800, 1549778400, 1549782000, 
    1549785600, 1549789200, 1549792800, 1549796400, 1549800000, 1549803600, 
    1549807200, 1549810800, 1549814400, 1549818000, 1549821600, 1549825200, 
    1549828800, 1549832400, 1549836000, 1549839600, 1549843200, 1549846800, 
    1549850400, 1549854000, 1549857600, 1549861200, 1549864800, 1549868400, 
    1549872000, 1549875600, 1549879200, 1549882800, 1549886400, 1549890000, 
    1549893600, 1549897200, 1549900800, 1549904400, 1549908000, 1549911600, 
    1549915200, 1549918800, 1549922400, 1549926000, 1549929600, 1549933200, 
    1549936800, 1549940400, 1549944000, 1549947600, 1549951200, 1549954800, 
    1549958400, 1549962000, 1549965600, 1549969200, 1549972800, 1549976400, 
    1549980000, 1549983600, 1549987200, 1549990800, 1549994400, 1549998000, 
    1550001600, 1550005200, 1550008800, 1550012400, 1550016000, 1550019600, 
    1550023200, 1550026800, 1550030400, 1550034000, 1550037600, 1550041200, 
    1550044800, 1550048400, 1550052000, 1550055600, 1550059200, 1550062800, 
    1550066400, 1550070000, 1550073600, 1550077200, 1550080800, 1550084400, 
    1550088000, 1550091600, 1550095200, 1550098800, 1550102400, 1550106000, 
    1550109600, 1550113200, 1550116800, 1550120400, 1550124000, 1550127600, 
    1550131200, 1550134800, 1550138400, 1550142000, 1550145600, 1550149200, 
    1550152800, 1550156400, 1550160000, 1550163600, 1550167200, 1550170800, 
    1550174400, 1550178000, 1550181600, 1550185200, 1550188800, 1550192400, 
    1550196000, 1550199600, 1550203200, 1550206800, 1550210400, 1550214000, 
    1550217600, 1550221200, 1550224800, 1550228400, 1550232000, 1550235600, 
    1550239200, 1550242800, 1550246400, 1550250000, 1550253600, 1550257200, 
    1550260800, 1550264400, 1550268000, 1550271600, 1550275200, 1550278800, 
    1550282400, 1550286000, 1550289600, 1550293200, 1550296800, 1550300400, 
    1550304000, 1550307600, 1550311200, 1550314800, 1550318400, 1550322000, 
    1550325600, 1550329200, 1550332800, 1550336400, 1550340000, 1550343600, 
    1550347200, 1550350800, 1550354400, 1550358000, 1550361600, 1550365200, 
    1550368800, 1550372400, 1550376000, 1550379600, 1550383200, 1550386800, 
    1550390400, 1550394000, 1550397600, 1550401200, 1550404800, 1550408400, 
    1550412000, 1550415600, 1550419200, 1550422800, 1550426400, 1550430000, 
    1550433600, 1550437200, 1550440800, 1550444400, 1550448000, 1550451600, 
    1550455200, 1550458800, 1550462400, 1550466000, 1550469600, 1550473200, 
    1550476800, 1550480400, 1550484000, 1550487600, 1550491200, 1550494800, 
    1550498400, 1550502000, 1550505600, 1550509200, 1550512800, 1550516400, 
    1550520000, 1550523600, 1550527200, 1550530800, 1550534400, 1550538000, 
    1550541600, 1550545200, 1550548800, 1550552400, 1550556000, 1550559600, 
    1550563200, 1550566800, 1550570400, 1550574000, 1550577600, 1550581200, 
    1550584800, 1550588400, 1550592000, 1550595600, 1550599200, 1550602800, 
    1550606400, 1550610000, 1550613600, 1550617200, 1550620800, 1550624400, 
    1550628000, 1550631600, 1550635200, 1550638800, 1550642400, 1550646000, 
    1550649600, 1550653200, 1550656800, 1550660400, 1550664000, 1550667600, 
    1550671200, 1550674800, 1550678400, 1550682000, 1550685600, 1550689200, 
    1550692800, 1550696400, 1550700000, 1550703600, 1550707200, 1550710800, 
    1550714400, 1550718000, 1550721600, 1550725200, 1550728800, 1550732400, 
    1550736000, 1550739600, 1550743200, 1550746800, 1550750400, 1550754000, 
    1550757600, 1550761200, 1550764800, 1550768400, 1550772000, 1550775600, 
    1550779200, 1550782800, 1550786400, 1550790000, 1550793600, 1550797200, 
    1550800800, 1550804400, 1550808000, 1550811600, 1550815200, 1550818800, 
    1550822400, 1550826000, 1550829600, 1550833200, 1550836800, 1550840400, 
    1550844000, 1550847600, 1550851200, 1550854800, 1550858400, 1550862000, 
    1550865600, 1550869200, 1550872800, 1550876400, 1550880000, 1550883600, 
    1550887200, 1550890800, 1550894400, 1550898000, 1550901600, 1550905200, 
    1550908800, 1550912400, 1550916000, 1550919600, 1550923200, 1550926800, 
    1550930400, 1550934000, 1550937600, 1550941200, 1550944800, 1550948400, 
    1550952000, 1550955600, 1550959200, 1550962800, 1550966400, 1550970000, 
    1550973600, 1550977200, 1550980800, 1550984400, 1550988000, 1550991600, 
    1550995200, 1550998800, 1551002400, 1551006000, 1551009600, 1551013200, 
    1551016800, 1551020400, 1551024000, 1551027600, 1551031200, 1551034800, 
    1551038400, 1551042000, 1551045600, 1551049200, 1551052800, 1551056400, 
    1551060000, 1551063600, 1551067200, 1551070800, 1551074400, 1551078000, 
    1551081600, 1551085200, 1551088800, 1551092400, 1551096000, 1551099600, 
    1551103200, 1551106800, 1551110400, 1551114000, 1551117600, 1551121200, 
    1551124800, 1551128400, 1551132000, 1551135600, 1551139200, 1551142800, 
    1551146400, 1551150000, 1551153600, 1551157200, 1551160800, 1551164400, 
    1551168000, 1551171600, 1551175200, 1551178800, 1551182400, 1551186000, 
    1551189600, 1551193200, 1551196800, 1551200400, 1551204000, 1551207600, 
    1551211200, 1551214800, 1551218400, 1551222000, 1551225600, 1551229200, 
    1551232800, 1551236400, 1551240000, 1551243600, 1551247200, 1551250800, 
    1551254400, 1551258000, 1551261600, 1551265200, 1551268800, 1551272400, 
    1551276000, 1551279600, 1551283200, 1551286800, 1551290400, 1551294000, 
    1551297600, 1551301200, 1551304800, 1551308400, 1551312000, 1551315600, 
    1551319200, 1551322800, 1551326400, 1551330000, 1551333600, 1551337200, 
    1551340800, 1551344400, 1551348000, 1551351600, 1551355200, 1551358800, 
    1551362400, 1551366000, 1551369600, 1551373200, 1551376800, 1551380400, 
    1551384000, 1551387600, 1551391200, 1551394800, 1551398400, 1551402000, 
    1551405600, 1551409200, 1551412800, 1551416400, 1551420000, 1551423600, 
    1551427200, 1551430800, 1551434400, 1551438000, 1551441600, 1551445200, 
    1551448800, 1551452400, 1551456000, 1551459600, 1551463200, 1551466800, 
    1551470400, 1551474000, 1551477600, 1551481200, 1551484800, 1551488400, 
    1551492000, 1551495600, 1551499200, 1551502800, 1551506400, 1551510000 ;

 latitude = 80.1058 ;

 longitude = 31.4643 ;

 air_pressure_at_sea_level = 98990, 99400, 100000, 100970, 101550, 101900, 
    102330, 102260, 102190, 101900, 102120, 102210, 102080, 102000, 101820, 
    101890, 102110, 102340, 102070, 101260, 100140, 99300, 99510, 100130, 
    100280, 100340, 99890, 99400, 98990, 99250, 99600, 99880, 100480, 100660, 
    100470, 100260, 100660, 102410, 102730, 102700, 102470, 101710, 100190, 
    99560, 98390, 98240, 98880, 100360, 100810, 100810, 100580, 100280, 
    100410, 101260, 101820, 99560, 99410, 100920, 100400, 99770, 103470, 
    103530, 103290, 102950, 102400, 101640, 100780, 100820, 101020, 101000, 
    100780, 100700, 100840, 100890, 101180, 101440, 101730, 101880, 101580, 
    100700, 99770, 100950, 101640, 101710, 101800, 101960, 101820, 101710, 
    101380, 101280, 101370, 101690, 102000, 102250, 102380, 102450, 102370, 
    102410, 102470, 102450, 102440, 102260, 102100, 101810, 101660, 101490, 
    101300, 101320, 101520, 102070, 102070, 101750, 101030, 101290, 100580, 
    100290, 99950, 100040, 100630, 101100, 104830, 101450, 101540, 101740, 
    101810, 101700, 101690, 101450, 101020, 100860, 100520, 100450, 100510, 
    100360, 100280, 100910, 101150, 101800, 101920, 101230, 100630, 99700, 
    99060, 97570, 98500, 99440, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 103060, 103070, 103080, 103060, 
    103050, 103050, 103050, 103050, 103050, 103020, 103010, 103020, 103020, 
    103020, 103010, 103020, 103000, 102990, 102990, 102990, 102980, 102990, 
    103000, 102990, 102980, 102980, 102980, 102880, 102850, 102840, 102830, 
    102810, 102800, 102780, 102780, 102810, 102800, 102790, 102750, 102760, 
    102750, 102710, 102710, 102700, 102680, 102590, 102650, 102610, 102620, 
    102630, 102620, 102580, 102560, 102550, 102560, 102500, 102480, 102450, 
    102460, 102460, 102440, 102420, 102380, 102350, 102350, 102340, 102330, 
    102310, 102320, 102310, 102300, 102320, 102310, 102300, 102330, 102320, 
    102290, 102250, 102240, 102220, 102170, 102150, 102160, 102100, 102150, 
    102110, 102090, 102120, 102110, 102100, 102070, 102050, 102060, 102040, 
    102060, 102050, 102060, 102030, 102020, 102020, 101980, 101990, 101930, 
    101950, 101970, 101940, 101950, 101950, 101930, 101920, 101930, 101940, 
    101930, 101920, 101930, 101920, 101930, 101910, 101930, 101920, 101910, 
    101910, 101940, 101930, 101920, 101940, 101900, 101910, 101920, 101930, 
    101930, 101920, 101930, 101950, 101950, 101960, 101980, 101990, 102010, 
    102020, 102040, 102060, 102090, 102120, 102160, 102190, 102200, 102220, 
    102230, 102240, 102250, 102270, 102280, 102290, 102300, 102330, 102330, 
    102330, 102350, 102340, 102340, 102330, 102330, 102260, 102330, 102320, 
    102280, 102260, 102250, 102300, 102280, 102300, 102300, 102280, 102260, 
    102260, 102260, 102250, 102250, 102280, 102320, 102320, 102330, 102340, 
    102350, 102350, 102340, 102330, 102300, 102310, 102330, 102330, 102330, 
    102360, 102370, 102380, 102370, 102380, 102360, 102330, 102330, 102320, 
    102320, 102320, 102310, 102290, 102290, 102260, 102270, 102270, 102260, 
    102230, 102210, 102210, 102230, 102220, 102250, 102260, 102280, 102270, 
    102250, 102210, 102170, 102160, 102160, 102130, 102120, 102110, 102100, 
    102090, 102080, 102070, 102050, 102020, 101990, 101980, 101980, 101950, 
    101930, 101910, 101900, 101890, 101870, 101860, 101830, 101820, 101780, 
    101740, 101710, 101670, 101670, 101670, 101630, 101630, 101610, 101580, 
    101580, 101540, 101520, 101490, 101480, 101480, 101470, 101490, 101480, 
    101490, 101480, 101470, 101470, 101460, 101450, 101450, 101440, 101430, 
    101440, 101440, 101420, 101430, 101410, 101400, 101390, 101390, 101380, 
    101360, 101330, 101320, 101330, 101330, 101330, 101330, 101320, 101320, 
    101300, 101320, 101280, 101270, 101260, 101260, 101250, 101240, 101240, 
    101210, 101210, 101200, 101210, 101190, 101200, 101190, 101190, 101210, 
    101230, 101260, 101270, 101280, 101310, 101330, 101340, 101350, 101360, 
    101380, 101390, 101400, 101390, 101400, 101420, 101440, 101450, 101450, 
    101460, 101480, 101480, 101480, 101500, 101500, 101510, 101520, 101540, 
    101520, 101540, 101530, 101530, 101520, 101490, 101460, 101430, 101410, 
    101410, 101400, 101370, 101360, 101350, 101320, 101310, 101270, 101250, 
    101210, 101180, 101140, 101130, 101090, 101070, 101020, 101000, 100950, 
    100910, 100860, 100840, 100810, 100780, 100730, 100700, 100660, 100640, 
    100600, 100590, 100560, 100540, 100480, 100480, 100490, 100490, 100500, 
    100520, 100530, 100570, 100620, 100680, 100720, 100750, 100800, 100850, 
    100900, 100950, 100970, 100990, 101050, 101100, 101150, 101180, 101230, 
    101270, 101310, 101310, 101340, 101340, 101340, 101340, 101330, 101340, 
    101340, 101320, 101310, 101340, 101380, 101410, 101410, 101480, 101530, 
    101550, 101590, 101640, 101690, 101730, 101760, 101760, 101770, 101760, 
    101760, 101730, 101730, 101730, 101680, 101660, 101620, 101580, 101500, 
    101460, 101430, 101360, 101350, 101330, 101260, 101200, 101180, 101140, 
    101110, 101080, 101040, 100990, 100930, 100920, 100880, 100820, 100790, 
    100720, 100680, 100570, 100540, 100460, 100410, 100390, 100320, 100250, 
    100230, 100220, 100220, 100230, 100220, 100240, 100230, 100250, 100260, 
    100230, 100220, 100240, 100230, 100250, 100280, 100280, 100350, 100360, 
    100390, 100400, 100400, 100470, 100540, 100570, 100600, 100620, 100630, 
    100620, 100640, 100680, 100710, 100810, 100790, 100790, 100780, 100770, 
    100750, 100750, 100690, 100740, 100720, 100700, 100580, 100590, 100310, 
    100270, 100220, 100140, 100090, 99930, 99850, 99840, 99720, 99710, 99730, 
    99750, 99770, 99750, 99770, 99760, 99740, 99760, 99820, 99830, 99860, 
    99890, 99930, 100020, 100040, 100090, 100060, 100090, 100120, 100120, 
    100160, 100190, 100220, 100250, 100240, 100270, 100340, 100390, 100430, 
    100480, 100510, 100570, 100650, 100720, 100800, 100810, 100860, 100920, 
    100950, 101000, 101030, 101060, 101120, 101150, 101170, 101190, 101200, 
    101240, 101270, 101280, 101270, 101250, 101250, 101220, 101190, 101160, 
    101080, 101020, 101040, 101030, 101000, 100970, 100890, 100810, 100700, 
    100580, 100610, 100560, 100550, 100500, 100500, 100490, 100470, 100420, 
    100390, 100370, 100370, 100340, 100320, 100330, 100330, 100360, 100380, 
    100380, 100430, 100440, 100490, 100510, 100530, 100540, 100570, 100560, 
    100590, 100590, 100590, 100600, 100570, 100560, 100550, 100520, 100510, 
    100490, 100460, 100440, 100430, 100400, 100390, 100370, 100340, 100320, 
    100280, 100270, 100290, 100290, 100320, 100360, 100450, 100460, 100560, 
    100600, 100650, 100700, 100770, 100810, 100850, 100920, 100940, 100950, 
    100990, 101010, 101000, 101010, 101040, 101030, 101020, 101030, 101020, 
    101000, 100990, 100940, 100930, 100870, 100800, 100720, 100650, 100530, 
    100540, 100540, 100460, 100330, 100360, 100080, 100000, 100050, 100130, 
    100010, 100010, 100020, 100010, 99990, 99980, 100000, 100020, 100040, 
    100050, 100070, 100100, 100130, 100160, 100160, 100160, 100130, 100130, 
    100120, 100150, 100150, 100150, 100120, 100120, 100100, 100140, 100140, 
    100130, 100130, 100130, 100120, 100080, 100070, 100070, 100070, 100080, 
    100080, 100060, 100040, 100030, 100000, 99990, 99990, 99980, 99980, 
    99940, 99940, 99950, 99960, 99950, 99960, 99970, 99950, 99920, 99940, 
    99930, 99900, 99880, 99860, 99840, 99830, 99850, 99830, 99820, 99810, 
    99770, 99740, 99750, 99760, 99750, 99770, 99780, 99790, 99810, 99830, 
    99840, 99880, 99910, 99940, 100000, 100060, 100050, 100120, 100160, 
    100230, 100270, 100310, 100340, 100360, 100390, 100430, 100480, 100460, 
    100490, 100510, 100560, 100610, 100620, 100700, 100720, 100730, 100730, 
    100710, 100710, 100680, 100670, 100640, 100600, 100550, 100550, 100540, 
    100470, 100480, 100490, 100460, 100510, 100540, 100590, 100610, 100630, 
    100670, 100770, 100840, 100880, 100900, 101040, 101140, 101230, 101310, 
    101400, 101470, 101500, 101570, 101640, 101660, 101720, 101750, 101790, 
    101880, 101900, 101950, 101970, 101990, 102030, 102030, 102070, 102090, 
    102120, 102130, 102140, 102140, 102130, 102150, 102170, 102170, 102150, 
    102140, 102120, 102150, 102050, 102080, 102030, 102010, 102060, 102110, 
    102100, 102130, 102150, 102130, 102110, 102130, 102120, 102110, 102100, 
    102120, 102130, 102160, 102150, 102150, 102150, 102150, 102150, 102120, 
    102110, 102080, 102080, 102080, 102080, 102080, 102090, 102090, 102080, 
    102070, 102060, 102050, 102040, 102000, 101990, 101980, 101960, 101910, 
    101890, 101880, 101850, 101830, 101800, 101760, 101720, 101670, 101600, 
    101560, 101540, 101520, 101530, 101530, 101580, 101610, 101610, 101600, 
    101560, 101540, 101510, 101500, 101500, 101500, 101510, 101530, 101520, 
    101510, 101520, 101500, 101530, 101560, 101590, 101620, 101640, 101660, 
    101670, 101710, 101730, 101740, 101750, 101760, 101750, 101750, 101740, 
    101750, 101740, 101730, 101710, 101700, 101720, 101680, 101660, 101640, 
    101610, 101560, 101540, 101510, 101490, 101450, 101400, 101360, 101350, 
    101330, 101340, 101310, 101290, 101260, 101230, 101200, 101180, 101130, 
    101080, 101020, 101000, 100940, 100900, 100880, 100820, 100760, 100720, 
    100680, 100740, 100720, 100720, 100710, 100720, 100740, 100740, 100760, 
    100740, 100750, 100750, 100740, 100740, 100700, 100700, 100670, 100680, 
    100650, 100640, 100590, 100570, 100550, 100470, 100440, 100420, 100420, 
    100460, 100470, 100500, 100510, 100530, 100560, 100580, 100570, 100580, 
    100590, 100600, 100570, 100560, 100540, 100510, 100500, 100500, 100480, 
    100460, 100400, 100370, 100370, 100350, 100310, 100290, 100260, 100230, 
    100240, 100240, 100230, 100190, 100160, 100150, 100110, 100110, 100110, 
    100110, 100080, 100040, 100100, 100090, 100010, 100030, 100030, 100010, 
    100010, 100020, 100000, 99980, 99990, 100000, 100010, 100000, 99990, 
    99990, 99980, 99960, 99930, 99930, 99930, 99940, 99940, 99940, 99970, 
    100030, 100090, 100100, 100140, 100160, 100200, 100240, 100300, 100380, 
    100490, 100560, 100630, 100680, 100760, 100850, 100930, 101000, 101090, 
    101180, 101250, 101290, 101360, 101430, 101460, 101470, 101460, 101460, 
    101470, 101460, 101440, 101420, 101400, 101400, 101410, 101370, 101360, 
    101310, 101240, 101230, 101150, 101050, 100960, 100870, 100730, 100580, 
    100500, 100370, 100260, 100120, 99970, 99840, 99710, 99570, 99450, 99370, 
    99240, 99220, 99180, 99190, 99230, 99220, 99250, 99290, 99360, 99430, 
    99520, 99560, 99590, 99670, 99690, 99780, 99840, 99890, 99950, 100000, 
    100080, 100130, 100160, 100230, 100250, 100290, 100330, 100370, 100420, 
    100440, 100500, 100550, 100560, 100610, 100670, 100680, 100700, 100720, 
    100710, 100730, 100750, 100760, 100760, 100750, 100750, 100740, 100740, 
    100730, 100680, 100680, 100680, 100680, 100700, 100700, 100690, 100680, 
    100670, 100720, 100730, 100700, 100700, 100710, 100690, 100680, 100680, 
    100670, 100670, 100680, 100650, 100650, 100630, 100630, 100630, 100610, 
    100620, 100620, 100620, 100620, 100630, 100630, 100600, 100570, 100550, 
    100530, 100500, 100480, 100450, 100430, 100410, 100380, 100350, 100320, 
    100280, 100250, 100200, 100190, 100190, 100180, 100160, 100170, 100190, 
    100210, 100230, 100250, 100240, 100230, 100250, 100250, 100250, 100250, 
    100220, 100210, 100210, 100210, 100200, 100180, 100170, 100150, 100120, 
    100090, 100070, 100050, 100020, 100000, 99980, 99970, 99940, 99920, 
    99900, 99880, 99890, 99870, 99870, 99880, 99870, 99890, 99870, 99870, 
    99850, 99840, 99830, 99800, 99820, 99800, 99750, 99820, 99790, 99810, 
    99840, 99860, 99860, 99840, 99810, 99820, 99820, 99820, 99820, 99820, 
    99840, 99870, 99890, 99890, 99890, 99910, 99930, 99930, 99910, 99920, 
    99930, 99960, 99980, 100010, 100030, 100070, 100100, 100130, 100150, 
    100130, 100130, 100170, 100190, 100180, 100210, 100260, 100240, 100250, 
    100250, 100250, 100250, 100250, 100240, 100200, 100150, 100180, 100200, 
    100250, 100300, 100290, 100300, 100280, 100280, 100290, 100270, 100290, 
    100260, 100230, 100180, 100200, 100220, 100210, 100180, 100170, 100130, 
    100130, 100110, 100090, 100090, 100070, 100070, 100060, 100050, 100060, 
    100020, 100010, 100000, 99990, 99980, 99990, 99980, 99960, 99960, 99970, 
    99990, 100000, 99990, 99990, 100000, 100010, 100010, 100010, 100020, 
    100050, 100090, 100130, 100160, 100220, 100260, 100290, 100300, 100340, 
    100390, 100440, 100480, 100510, 100520, 100550, 100580, 100620, 100670, 
    100700, 100720, 100760, 100790, 100810, 100810, 100840, 100850, 100920, 
    101030, 101140, 101190, 101230, 101280, 101330, 101360, 101440, 101480, 
    101530, 101580, 101650, 101700, 101770, 101820, 101840, 101840, 101870, 
    101910, 101940, 101930, 101990, 102000, 101970, 101960, 101990, 101940, 
    101890, 101830, 101750, 101650, 101510, 101360, 101220, 101030, 100820, 
    100670, 100440, 100170, 99920, 99710, 99500, 99250, 99040, 98830, 98540, 
    98460, 98550, 98610, 98600, 98580, 98560, 98530, 98530, 98520, 98510, 
    98460, 98440, 98450, 98460, 98460, 98480, 98490, 98520, 98560, 98620, 
    98710, 98750, 98770, 98850, 98940, 99050, 99140, 99220, 99280, 99340, 
    99400, 99420, 99450, 99450, 99440, 99440, 99570, 99640, 99680, 99710, 
    99710, 99740, 99740, 99720, 99720, 99770, 99790, 99880, 99930, 99930, 
    99920, 99940, 100010, 100060, 100110, 100090, 100090, 100070, 100150, 
    100290, 100290, 100340, 100300, 100250, 100300, 100310, 100230, 100210, 
    100240, 100240, 100290, 100290, 100270, 100270, 100250, 100260, 100250, 
    100250, 100300, 100280, 100300, 100390, 100410, 100420, 100450, 100550, 
    100590, 100670, 100700, 100760, 100780, 100810, 100830, 100830, 100830, 
    100850, 100910, 100950, 100930, 100890, 100900, 100910, 100930, 100920, 
    100900, 100890, 100900, 100860, 100820, 100800, 100760, 100740, 100680, 
    100590, 100540, 100510, 100470, 100440, 100410, 100380, 100360, 100370, 
    100360, 100350, 100330, 100320, 100310, 100270, 100270, 100250, 100230, 
    100300, 100330, 100310, 100320, 100360, 100420, 100480, 100540, 100610, 
    100660, 100710, 100750, 100790, 100850, 100910, 100940, 100990, 101040, 
    101060, 101110, 101150, 101190, 101200, 101240, 101280, 101290, 101310, 
    101350, 101370, 101390, 101410, 101460, 101490, 101540, 101580, 101620, 
    101630, 101690, 101740, 101780, 101830, 101860, 101910, 101930, 101970, 
    101990, 102020, 102050, 102080, 102120, 102150, 102170, 102210, 102230, 
    102240, 102240, 102260, 102280, 102300, 102290, 102300, 102330, 102350, 
    102350, 102370, 102350, 102330, 102320, 102310, 102270, 102220, 102160, 
    102130, 102040, 101990, 101940, 101860, 101760, 101640, 101550, 101380, 
    101250, 101130, 101000, 100840, 100650, 100480, 100240, 100060, 99910, 
    99760, 99690, 99610, 99520, 99430, 99360, 99300, 99280, 99240, 99230, 
    99240, 99240, 99250, 99270, 99300, 99370, 99430, 99510, 99590, 99630, 
    99700, 99800, 99880, 100010, 100130, 100260, 100410, 100540, 100710, 
    100780, 100910, 101050, 101120, 101220, 101280, 101360, 101410, 101480, 
    101560, 101580, 101660, 101740, 101780, 101870, 101930, 102000, 102100, 
    102170, 102230, 102260, 102320, 102370, 102400, 102410, 102430, 102420, 
    102400, 102380, 102400, 102380, 102360, 102320, 102290, 102290, 102240, 
    102210, 102200, 102210, 102220, 102220, 102230, 102210, 102230, 102240, 
    102210, 102230, 102220, 102160, 102110, 102080, 102050, 102010, 101950, 
    101850, 101780, 101730, 101640, 101600, 101500, 101370, 101320, 101270, 
    101230, 101170, 101110, 101040, 100950, 100840, 100780, 100690, 100550, 
    100440, 100290, 100190, 100080, 100040, 99980, 99900, 99850, 99780, 
    99730, 99660, 99650, 99630, 99590, 99600, 99660, 99730, 99770, 99800, 
    99810, 99840, 99880, 99820, 99800, 99750, 99690, 99680, 99800, 99760, 
    99760, 99760, 99700, 99690, 99660, 99630, 99620, 99550, 99500, 99510, 
    99440, 99410, 99360, 99290, 99250, 99170, 99090, 99130, 99150, 99120, 
    99100, 99090, 99130, 99140, 99230, 99260, 99290, 99410, 99430, 99580, 
    99630, 99740, 99810, 99850, 99910, 100010, 100060, 100080, 100060, 
    100150, 100150, 100220, 100280, 100300, 100340, 100420, 100480, 100520, 
    100530, 100570, 100530, 100550, 100530, 100470, 100440, 100310, 100310, 
    100330, 100300, 100300, 100290, 100270, 100280, 100190, 100190, 100190, 
    100210, 100260, 100320, 100350, 100370, 100390, 100460, 100510, 100540, 
    100580, 100640, 100680, 100730, 100760, 100820, 100900, 100960, 101020, 
    101050, 101090, 101130, 101210, 101250, 101300, 101330, 101380, 101410, 
    101490, 101530, 101600, 101630, 101700, 101730, 101760, 101810, 101850, 
    101880, 101910, 101950, 101990, 102030, 102070, 102110, 102150, 102190, 
    102220, 102230, 102250, 102270, 102310, 102350, 102370, 102390, 102430, 
    102440, 102490, 102490, 102500, 102490, 102480, 102470, 102460, 102410, 
    102410, 102380, 102360, 102350, 102300, 102270, 102250, 102190, 102190, 
    102130, 102050, 101940, 101860, 101770, 101700, 101650, 101570, 101470, 
    101340, 101220, 101150, 101080, 101010, 100900, 100820, 100710, 100640, 
    100600, 100540, 100450, 100350, 100310, 100250, 100230, 100180, 100140, 
    100100, 100080, 100000, 99980, 99880, 99860, 99760, 99680, 99590, 99560, 
    99480, 99350, 99300, 99210, 99090, 99020, 98960, 98880, 98840, 98850, 
    98910, 98990, 99050, 99110, 99170, 99160, 99210, 99230, 99260, 99260, 
    99170, 99060, 98990, 98870, 98790, 98690, 98590, 98500, 98410, 98310, 
    98170, 98090, 97960, 97850, 97780, 97720, 97690, 97700, 97720, 97740, 
    97790, 97860, 97890, 98010, 98100, 98190, 98290, 98390, 98510, 98640, 
    98790, 98890, 99000, 99190, 99410, 99620, 99760, 99900, 100010, 100070, 
    100030, 100100, 100150, 100250, 100280, 100360, 100410, 100420, 100430, 
    100470, 100470, 100460, 100520, 100480, 100490, 100500, 100510, 100520, 
    100510, 100510, 100470, 100470, 100460, 100430, 100410, 100400, 100390, 
    100380, 100420, 100400, 100410, 100480, 100510, 100490, 100440, 100420, 
    100390, 100390, 100420, 100430, 100420, 100490, 100530, 100610, 100660, 
    100650, 100750, 101250, 101250, 101250, 101220, 101200, 101190, 101190, 
    101160, 101100, 101090, 101060, 100960, 100900, 100860, 100820, 100790, 
    100750, 100670, 100670, 100670, 100670, 100680, 100690, 100680, 100720, 
    100770, 100830, 100850, 100890, 101000, 101070, 101130, 101180, 101240, 
    101280, 101350, 101360, 101400, 101430, 101450, 101480, 101500, 101540, 
    101570, 101590, 101640, 101670, 101690, 101700, 101710, 101730, 101740, 
    101740, 101690, 101680, 101690, 101700, 101700, 101700, 101640, 101640, 
    101630, 101620, 101610, 101610, 101580, 101580, 101590, 101600, 101600, 
    101600, 101640, 101640, 101640, 101630, 101630, 101630, 101630, 101640, 
    101650, 101660, 101660, 101670, 101720, 101730, 101730, 101730, 101730, 
    101730, 101690, 101720, 101710, 101700, 101720, 101730, 101810, 101820, 
    101820, 101820, 101790, 101770, 101700, 101700, 101690, 101700, 101690, 
    101680, 101680, 101650, 101630, 101620, 101590, 101570, 101560, 101550, 
    101560, 101560, 101550, 101540, 101590, 101570, 101570, 101560, 101520, 
    101500, 101430, 101440, 101420, 101400, 101380, 101370, 101360, 101330, 
    101320, 101300, 101260, 101230, 101180, 101160, 101140, 101120, 101100, 
    101060, 100940, 100920, 100880, 100850, 100810, 100770, 100690, 100650, 
    100580, 100510, 100380, 100300, 100190, 100070, 99950, 99830, 99720, 
    99610, 99480, 99460, 99410, 99420, 99410, 99440, 99320, 99320, 99310, 
    99290, 99250, 99230, 99180, 99110, 99070, 98960, 98870, 98830, 98430, 
    98440, 98460, 98470, 98500, 98490, 98510, 98470, 98390, 98310, 98190, 
    97930, 97680, 97500, 97340, 97260, 97210, 97210, 97200, 97200, 97190, 
    97220, 97260, 97310, 97350, 97380, 97410, 97420, 97440, 97450, 97460, 
    97480, 97490, 97550, 97590, 97750, 97780, 97830, 97830, 97820, 97850, 
    97900, 97950, 97980, 98010, 98070, 98070, 98150, 98160, 98180, 98190, 
    98190, 98210, 98130, 98150, 98190, 98200, 98220, 98230, 98220, 98250, 
    98270, 98280, 98280, 98290, 98270, 98310, 98320, 98340, 98370, 98400, 
    98430, 98450, 98480, 98500, 98480, 98490, 98460, 98460, 98480, 98510, 
    98500, 98510, 98520, 98530, 98520, 98520, 98530, 98550, 98550, 98570, 
    98580, 98590, 98600, 98630, 98620, 98630, 98640, 98660, 98660, 98680, 
    98580, 98610, 98640, 98650, 98670, 98680, 98690, 98690, 98690, 98710, 
    98760, 98780, 98740, 98780, 98820, 98860, 98920, 98980, 99110, 99150, 
    99190, 99240, 99260, 99300, 99330, 99390, 99440, 99480, 99520, 99560, 
    99630, 99670, 99720, 99780, 99820, 99850, 99890, 99920, 99950, 99990, 
    100040, 100070, 100150, 100160, 100190, 100180, 100170, 100220, 100240, 
    100250, 100260, 100270, 100230, 100220, 100070, 100040, 100010, 99990, 
    99960, 99880, 99840, 99800, 99730, 99660, 99590, 99550, 99460, 99330, 
    99230, 99130, 99010, 98840, 98730, 98550, 98380, 98210, 98050, 97860, 
    97670, 97490, 97330, 97170, 97010, 96840, 96710, 96580, 96470, 96360, 
    96250, 96150, 96050, 95980, 95930, 95900, 95870, 95900, 96070, 96110, 
    96130, 96100, 96080, 96060, 96000, 95930, 95860, 95820, 95760, 95690, 
    95690, 95680, 95690, 95720, 95750, 95800, 95810, 95870, 95940, 95990, 
    96040, 96100, 96160, 96210, 96250, 96280, 96310, 96350, 96320, 96350, 
    96390, 96430, 96460, 96510, 96500, 96580, 96650, 96720, 96780, 96830, 
    96870, 96940, 97000, 97010, 97010, 97090, 97150, 97220, 97280, 97320, 
    97360, 97410, 97470, 97540, 97610, 97680, 97730, 97780, 97920, 97980, 
    98050, 98110, 98160, 98210, 98290, 98360, 98420, 98440, 98440, 98480, 
    98560, 98590, 98600, 98620, 98660, 98690, 98660, 98680, 98720, 98780, 
    98820, 98860, 98940, 98990, 99040, 99080, 99130, 99190, 99180, 99210, 
    99240, 99270, 99260, 99310, 99300, 99320, 99340, 99360, 99340, 99370, 
    99300, 99280, 99260, 99240, 99240, 99220, 99190, 99190, 99170, 99120, 
    99080, 99060, 99090, 99060, 99030, 99030, 99010, 98980, 98970, 98930, 
    98910, 98880, 98860, 98850, 99610, 99620, 99630, 99640, 99660, 99670, 
    99700, 99720, 99740, 99740, 99760, 99690, 99690, 99710, 99720, 99740, 
    99760, 99720, 99740, 99740, 99750, 99790, 99820, 99860, 99890, 99920, 
    99940, 99980, 100050, 99930, 99980, 100030, 100090, 100130, 100180, 
    100260, 100310, 100380, 100410, 100410, 100440, 100470, 100500, 100560, 
    100570, 100610, 100620, 100620, 100620, 100610, 100600, 100570, 100570, 
    100510, 100490, 100460, 100420, 100380, 100360, 100370, 100360, 100340, 
    100330, 100300, 100260, 100250, 100250, 100250, 100260, 100270, 100250, 
    100240, 100260, 100260, 100230, 100250, 100240, 100240, 100250, 100260, 
    100280, 100300, 100280, 100290, 100300, 100270, 100280, 100320, 100290, 
    100330, 100350, 100380, 100420, 100410, 100390, 100430, 100440, 100420, 
    100420, 100430, 100340, 100360, 100390, 100410, 100420, 100420, 100360, 
    100390, 100430, 100460, 100480, 100510, 100530, 100570, 100590, 100620, 
    100670, 100710, 100700, 100730, 100770, 100760, 100770, 100810, 100850, 
    100880, 100950, 100990, 101010, 101030, 101050, 101100, 101100, 101120, 
    101120, 101140, 101160, 101150, 101160, 101170, 101200, 101190, 101160, 
    101140, 101100, 101110, 101030, 100990, 100460, 100480, 100490, 100520, 
    101070, 101100, 101130, 101160, 101190, 101220, 101260, 101260, 101280, 
    101280, 101300, 101310, 101250, 101280, 101310, 101350, 101360, 101350, 
    101410, 101410, 101430, 101420, 101420, 101420, 101360, 101360, 101360, 
    101380, 101380, 101360, 101350, 101330, 101300, 101280, 101240, 101220, 
    101170, 101170, 101150, 101140, 101130, 101110, 101090, 101060, 101010, 
    100990, 100940, 100900, 100800, 100750, 100680, 100610, 100560, 100510, 
    100480, 100410, 100350, 100300, 100220, 100150, 100060, 100010, 99950, 
    99870, 99790, 99700, 99600, 99510, 99430, 99350, 99240, 99140, 98990, 
    98880, 98760, 98640, 98540, 98410, 98320, 98240, 98150, 98030, 97930, 
    97840, 97730, 97620, 97510, 97410, 97310, 97220, 97310, 97220, 97110, 
    97030, 96960, 96930, 96900, 96950, 97020, 97060, 97110, 97150, 97190, 
    97220, 97220, 97200, 97220, 97240, 97100, 97120, 97150, 97200, 97250, 
    97310, 97330, 97360, 97390, 97410, 97420, 97450, 97420, 97440, 97460, 
    97480, 97490, 97490, 97480, 97490, 97490, 97490, 97470, 97490, 97520, 
    97560, 97590, 97600, 97620, 97620, 97660, 97650, 97660, 97650, 97620, 
    97610, 97540, 97530, 97500, 97480, 97480, 97480, 97410, 97400, 97390, 
    97400, 97420, 97460, 97430, 97460, 97480, 97500, 97560, 97600, 97600, 
    97640, 97690, 97720, 97780, 97840, 97830, 97890, 97950, 98010, 98070, 
    98130, 98280, 98340, 98400, 98440, 98490, 98550, 98650, 98670, 98710, 
    98730, 98780, 98820, 99060, 99110, 99160, 99200, 99230, 99310, 99380, 
    99400, 99440, 99460, 99490, 99530, 99570, 99590, 99610, 99640, 99680, 
    99710, 99740, 99760, 99790, 99820, 99870, 99900, 99950, 99970, 100000, 
    100040, 100070, 100120, 100180, 100220, 100270, 100290, 100320, 100360, 
    100420, 100420, 100440, 100460, 100490, 100520, 100590, 100610, 100640, 
    100680, 100730, 100750, 100790, 100800, 100840, 100860, 100860, 100880, 
    100840, 100870, 100900, 100910, 100930, 100950, 100920, 100890, 100890, 
    100920, 100950, 100960, 101000, 101010, 101030, 101040, 101060, 101040, 
    100940, 100930, 100920, 100930, 100910, 100890, 100880, 100880, 100880, 
    100890, 100880, 100890, 100820, 100780, 100750, 100740, 100750, 100750, 
    100770, 100810, 100840, 100890, 100920, 100970, 101050, 101060, 101090, 
    101120, 101120, 101110, 101130, 101140, 101150, 101130, 101100, 101070, 
    101050, 101020, 100980, 100940, 100910, 100890, 100960, 100950, 100950, 
    100970, 101040, 100990, 100990, 101020, 101020, 101020, 101000, 101020, 
    101000, 101010, 101020, 101040, 101040, 101020, 101000, 101000, 101030, 
    101030, 101030, 101080, 101090, 101110, 101110, 101120, 101110, 101070, 
    101060, 101060, 101060, 101060, 101090, 101150, 101170, 101200, 101210, 
    101230, 101260, 101320, 101330, 101370, 101380, 101390, 101420, 101410, 
    101430, 101420, 101450, 101480, 101490, 101560, 101560, 101570, 101580, 
    101570, 101580, 101590, 101600, 101620, 101640, 101660, 101700, 101700, 
    101690, 101700, 101700, 101690, 101720, 101690, 101700, 101720, 101720, 
    101750, 101760, 101860, 101880, 101900, 101900, 101900, 101910, 101930, 
    101970, 102000, 102020, 102050, 102060, 102010, 102020, 102020, 102020, 
    102020, 102020, 102010, 102020, 102010, 101990, 101980, 101980, 102000, 
    101980, 101970, 101960, 101930, 101930, 101910, 101880, 101860, 101840, 
    101820, 101800, 101840, 101800, 101770, 101770, 101760, 101750, 101690, 
    101690, 101690, 101700, 101710, 101710, 101690, 101670, 101660, 101660, 
    101650, 101650, 101640, 101620, 101610, 101600, 101590, 101580, 101590, 
    101550, 101530, 101510, 101500, 101490, 101490, 101480, 101460, 101440, 
    101440, 101440, 101490, 101490, 101480, 101470, 101470, 101450, 101490, 
    101490, 101490, 101500, 101490, 101490, 101530, 101510, 101490, 101460, 
    101470, 101500, 101520, 101510, 101530, 101540, 101560, 101580, 101570, 
    101580, 101590, 101610, 101600, 101600, 101620, 101640, 101640, 101650, 
    101660, 101660, 101630, 101630, 101600, 101570, 101540, 101520, 101490, 
    101470, 101010, 101030, 101040, 101050, 101050, 101060, 101130, 101140, 
    101130, 101120, 101130, 101120, 101080, 101070, 101070, 101090, 101090, 
    101080, 101070, 101060, 101050, 101050, 101070, 101090, 101040, 101010, 
    100980, 100910, 100840, 100740, 100690, 100570, 100450, 100300, 100160, 
    100020, 99940, 99770, 99610, 99480, 99370, 99270, 99120, 99080, 99050, 
    99030, 98990, 98950, 98910, 98830, 98730, 98630, 98510, 98400, 98450, 
    98390, 98340, 98310, 98360, 98440, 98580, 98660, 98710, 98760, 98830, 
    98910, 99040, 99130, 99260, 99390, 99520, 99630, 99740, 99870, 99980, 
    100100, 100170, 100210, 100170, 100190, 100260, 100310, 100340, 100340, 
    100380, 100360, 100310, 100270, 100210, 100140, 100110, 100060, 100020, 
    99970, 99940, 99900, 99970, 99930, 99890, 99850, 99840, 99860, 99970, 
    99990, 100030, 100080, 100150, 100230, 100360, 100390, 100420, 100440, 
    100440, 100460, 100500, 100500, 100500, 100510, 100540, 100560, 100570, 
    100570, 100600, 100590, 100570, 100580, 100630, 100640, 100650, 100660, 
    100660, 100680, 100730, 100710, 100700, 100710, 100720, 100720, 100730, 
    100730, 100730, 100730, 100740, 100730, 100640, 100630, 100640, 100640, 
    100620, 100630, 100610, 100580, 100580, 100580, 100590, 100590, 100520, 
    100520, 100530, 100530, 100520, 100530, 100550, 100580, 100590, 100610, 
    100640, 100670, 100680, 100720, 100760, 100800, 100800, 100820, 100920, 
    100960, 100990, 101030, 101080, 101130, 101230, 101270, 101300, 101310, 
    101320, 101360, 101390, 101430, 101480, 101530, 101590, 101630, 101670, 
    101710, 101760, 101790, 101820, 101840, 101840, 101860, 101870, 101890, 
    101900, 101920, 101980, 102000, 102030, 102050, 102080, 102090, 102130, 
    102160, 102220, 102290, 102370, 102450, 102500, 102550, 102590, 102660, 
    102680, 102720, 102770, 102810, 102840, 102880, 102910, 102940, 102970, 
    103000, 103020, 103040, 103050, 103050, 102980, 102980, 102990, 103020, 
    103030, 103010, 103000, 103000, 102980, 102940, 102890, 102830, 102780, 
    102760, 102720, 102680, 102640, 102580, 102510, 102460, 102400, 102320, 
    102230, 102140, 102060, 101980, 101910, 101840, 101770, 101710, 101640, 
    101570, 101510, 101450, 101360, 101300, 101200, 101160, 101120, 101100, 
    101080, 101060, 101040, 101050, 101060, 101090, 101120, 101140, 101210, 
    101260, 101330, 101390, 101480, 101580, 101700, 101780, 101850, 101930, 
    101990, 102070, 102140, 102230, 102300, 102350, 102400, 102440, 102520, 
    102580, 102650, 102650, 102700, 102750, 102780, 102770, 102780, 102790, 
    102820, 102820, 102790, 102750, 102700, 102640, 102550, 102480, 102550, 
    102480, 102430, 102400, 102370, 102340, 102360, 102300, 102260, 102230, 
    102190, 102160, 102240, 102200, 102150, 102110, 102120, 102080, 102100, 
    102090, 102050, 102010, 101980, 101950, 101860, 101820, 101760, 101710, 
    101670, 101600, 101570, 101490, 101410, 101320, 101270, 101240, 101320, 
    101400, 101530, 101690, 101860, 102020, 102040, 102150, 102240, 102310, 
    102360, 102420, 102530, 102600, 102670, 102710, 102740, 102740, 102790, 
    102790, 102780, 102750, 102740, 102710, 102740, 102720, 102670, 102620, 
    102610, 102570, 102510, 102450, 102360, 102310, 102270, 102190, 102090, 
    102000, 101910, 101850, 101720, 101580, 101540, 101460, 101380, 101320, 
    101270, 101240, 101230, 101270, 101340, 101430, 101520, 101620, 101710, 
    101760, 101850, 101950, 102010, 102070, 102140, 102180, 102190, 102200, 
    102170, 102130, 102260, 102290, 102290, 102260, 102270, 102250, 102240, 
    102230, 102210, 102180, 102170, 102110, 101980, 101920, 101830, 101770, 
    101680, 101640, 101540, 101530, 101520, 101540, 101550, 101590, 101730, 
    101650, 101610, 101530, 101420, 101310, 101170, 101080, 100940, 100790, 
    100640, 100530, 100350, 100290, 100230, 100300, 100450, 100630, 100660, 
    100830, 101020, 101230, 101390, 101560, 101800, 101910, 102030, 102100, 
    102160, 102240, 102330, 102370, 102390, 102420, 102440, 102480, 102510, 
    102480, 102410, 102380, 102270, 102170, 102050, 101910, 101740, 101590, 
    101500, 101410, 101240, 101180, 101110, 101030, 100960, 100880, 100910, 
    100840, 100750, 100680, 100400, 100290, 100250, 100200, 100190, 100230, 
    100350, 100380, 100470, 100670, 100810, 100930, 101050, 101090, 101200, 
    101320, 101430, 101480, 101510, 101520, 101540, 101520, 101490, 101420, 
    101310, 101180, 101080, 100990, 100920, 100870, 100780, 100750, 100810, 
    100850, 100920, 100950, 101030, 101130, 101190, 101300, 101420, 101510, 
    101630, 101790, 101890, 101970, 102050, 102100, 102120, 102200, 102170, 
    102170, 102150, 102100, 102080, 102130, 102090, 102090, 102090, 102080, 
    102090, 102090, 102080, 102060, 102040, 102020, 102000, 101930, 101940, 
    101930, 101900, 101870, 101840, 101800, 101780, 101690, 101640, 101600, 
    101590, 101670, 101640, 101570, 101550, 101560, 101550, 101590, 101590, 
    101560, 101530, 101540, 101530, 101540, 101530, 101510, 101500, 101510, 
    101450, 101410, 101390, 101350, 101320, 101250, 101190, 101190, 101170, 
    101060, 101000, 100980, 100930, 100880, 100810, 100760, 100690, 100660, 
    100670, 100740, 100740, 100710, 100680, 100640, 100600, 100390, 100270, 
    100150, 100040, 99910, 99810, 99790, 99690, 99580, 99490, 99420, 99380, 
    99370, 99450, 99560, 99670, 99740, 99820, 99820, 99820, 99810, 99810, 
    99810, 99900, 99940, 99980, 100010, 100050, 100100, 100130, 100160, 
    100190, 100220, 100250, 100260, 100270, 100280, 100290, 100290, 100260, 
    100220, 100210, 100180, 100130, 100090, 100060, 100030, 99980, 99910, 
    99850, 99800, 99760, 99730, 99680, 99640, 99610, 99580, 99570, 99560, 
    99540, 99520, 99500, 99500, 99480, 99480, 99530, 99570, 99600, 99630, 
    99690, 99720, 99720, 99750, 99780, 99810, 99830, 99850, 99860, 99890, 
    99900, 99910, 99940, 99940, 99920, 99920, 99910, 99900, 99900, 99890, 
    99850, 99860, 99870, 99870, 99870, 99880, 99890, 99910, 99930, 99930, 
    99930, 99930, 99900, 99880, 99880, 99870, 99870, 99880, 99900, 99910, 
    99900, 99890, 99880, 99880, 99880, 99890, 99900, 99930, 99950, 99960, 
    99830, 99860, 99870, 99890, 99890, 99920, 100030, 100050, 100060, 100070, 
    100080, 100100, 100160, 100170, 100170, 100160, 100150, 100150, 100160, 
    100180, 100190, 100210, 100230, 100220, 100230, 100220, 100200, 100130, 
    100060, 99990, 99930, 99840, 99750, 99650, 99560, 99430, 99250, 99190, 
    99080, 99000, 98960, 98910, 98960, 98950, 98900, 98880, 98860, 98830, 
    98790, 98740, 98690, 98640, 98610, 98590, 98440, 98460, 98540, 98720, 
    98910, 99050, 99120, 99180, 99210, 99250, 99270, 99280, 99290, 99310, 
    99330, 99340, 99350, 99380, 99400, 99410, 99430, 99450, 99440, 99440, 
    99420, 99410, 99400, 99380, 99370, 99370, 99380, 99370, 99380, 99380, 
    99390, 99410, 99370, 99370, 99400, 99400, 99420, 99390, 99450, 99450, 
    99410, 99410, 99370, 99360, 99420, 99430, 99430, 99420, 99410, 99400, 
    99380, 99380, 99370, 99360, 99330, 99310, 99260, 99240, 99240, 99220, 
    99200, 99170, 99250, 99230, 99200, 99190, 99160, 99150, 99150, 99140, 
    99140, 99150, 99160, 99150, 99160, 99190, 99210, 99200, 99190, 99190, 
    99140, 99180, 99220, 99250, 99280, 99290, 99340, 99360, 99370, 99390, 
    99390, 99370, 99330, 99350, 99340, 99320, 99310, 99280, 99310, 99300, 
    99270, 99230, 99180, 99110, 99180, 99110, 99050, 99000, 98940, 98880, 
    98850, 98790, 98750, 98700, 98660, 98630, 98660, 98650, 98610, 98610, 
    98580, 98560, 98520, 98520, 98520, 98500, 98450, 98390, 98310, 98260, 
    98170, 98100, 98070, 98030, 98090, 98070, 98070, 98070, 98060, 98050, 
    97920, 97950, 97990, 98060, 98140, 98200, 98300, 98320, 98330, 98330, 
    98280, 98250, 98280, 98260, 98240, 98210, 98200, 98160, 97930, 97880, 
    97840, 97800, 97770, 97740, 97880, 97940, 98020, 98090, 98160, 98230, 
    98340, 98370, 98400, 98450, 98470, 98480, 98500, 98520, 98540, 98550, 
    98570, 98590, 98670, 98680, 98680, 98670, 98640, 98610, 98610, 98620, 
    98610, 98620, 98630, 98630, 98910, 98920, 98940, 98980, 98990, 99000, 
    99020, 99020, 99040, 99050, 99060, 99080, 99170, 99180, 99190, 99210, 
    99210, 99210, 99250, 99250, 99250, 99260, 99290, 99330, 99320, 99360, 
    99430, 99480, 99500, 99540, 99610, 99640, 99660, 99690, 99710, 99710, 
    99860, 99880, 99900, 99910, 99920, 99940, 100000, 100030, 100070, 100120, 
    100170, 100190, 100230, 100270, 100310, 100320, 100320, 100330, 100460, 
    100460, 100470, 100480, 100500, 100520, 100550, 100540, 100550, 100530, 
    100510, 100510, 100490, 100470, 100460, 100440, 100420, 100410, 100470, 
    100440, 100400, 100340, 100290, 100260, 100210, 100160, 100140, 100100, 
    100090, 100080, 100040, 100060, 100060, 100030, 100020, 100020, 100010, 
    100010, 100020, 100050, 100080, 100070, 100090, 100090, 100110, 100110, 
    100100, 100080, 100100, 100090, 100090, 100080, 100060, 100030, 100000, 
    100000, 100010, 100000, 99970, 99940, 99880, 99850, 99830, 99810, 99800, 
    99770, 99800, 99760, 99740, 99700, 99650, 99590, 99430, 99370, 99280, 
    99190, 99110, 99040, 98920, 98840, 98770, 98700, 98620, 98560, 98530, 
    98530, 98520, 98520, 98530, 98530, 98500, 98490, 98470, 98460, 98450, 
    98470, 98440, 98490, 98540, 98610, 98690, 98760, 98780, 98880, 98970, 
    99050, 99110, 99180, 99210, 99300, 99370, 99450, 99550, 99640, 99790, 
    99900, 100000, 100080, 100150, 100220, 100340, 100410, 100470, 100550, 
    100650, 100770, 100830, 100920, 100990, 101070, 101150, 101200, 101280, 
    101360, 101390, 101460, 101550, 101620, 101720, 101770, 101790, 101830, 
    101840, 101840, 101810, 101820, 101830, 101840, 101800, 101740, 101690, 
    101620, 101540, 101440, 101360, 101310, 101320, 101290, 101250, 101250, 
    101280, 101280, 101280, 101280, 101310, 101310, 101310, 101330, 101400, 
    101420, 101430, 101460, 101500, 101530, 101510, 101520, 101560, 101580, 
    101590, 101610, 101560, 101550, 101450, 101450, 101460, 101430, 101420, 
    101460, 101420, 101390, 101400, 101350, 101300, 101260, 101320, 101300, 
    101250, 101260, 101220, 101180, 101170, 101180, 101140, 101120, 101190, 
    101220, 101260, 101310, 101360, 101370, 101410, 101430, 101420, 101440, 
    101430, 101420, 101420, 101430, 101460, 101490, 101550, 101580, 101610, 
    101630, 101670, 101690, 101710, 101740, 101770, 101800, 101800, 101830, 
    101860, 101880, 101880, 101860, 101860, 101860, 101870, 101900, 101920, 
    101930, 101940, 101980, 102030, 102050, 102030, 101960, 101940, 101910, 
    101870, 101830, 101790, 101730, 101720, 101750, 101790, 101780, 101720, 
    101700, 101680, 101630, 101600, 101550, 101500, 101500, 101430, 101360, 
    101330, 101280, 101150, 101070, 101050, 101030, 100970, 100940, 100900, 
    100860, 100790, 100750, 100680, 100610, 100530, 100420, 100370, 100310, 
    100240, 100180, 100130, 100090, 100050, 100010, 99930, 99860, 99830, 
    99740, 99680, 99680, 99610, 99510, 99430, 99350, 99260, 99180, 99100, 
    99050, 98970, 98900, 98780, 98710, 98660, 98650, 98600, 98500, 98360, 
    98330, 98300, 98280, 98180, 98140, 98110, 98070, 98060, 97980, 97960, 
    97960, 97940, 97930, 97920, 97930, 97960, 97970, 97960, 97990, 98020, 
    98050, 98090, 98120, 98160, 98210, 98280, 98340, 98390, 98460, 98520, 
    98600, 98650, 98700, 98750, 98790, 98840, 98900, 98960, 99040, 99080, 
    99120, 99160, 99220, 99260, 99290, 99330, 99370, 99390, 99420, 99470, 
    99510, 99550, 99600, 99650, 99700, 99730, 99810, 99830, 99920, 100000, 
    100090, 100160, 100230, 100290, 100340, 100400, 100450, 100490, 100550, 
    100580, 100610, 100640, 100710, 100790, 100830, 100860, 100890, 100940, 
    100970, 101050, 101120, 101140, 101160, 101230, 101250, 101270, 101360, 
    101400, 101420, 101430, 101470, 101470, 101480, 101490, 101480, 101490, 
    101510, 101480, 101490, 101490, 101470, 101460, 101430, 101400, 101340, 
    101290, 101240, 101210, 101160, 101140, 101090, 101040, 101000, 100910, 
    100820, 100760, 100660, 100570, 100470, 100380, 100310, 100260, 100200, 
    100120, 100050, 100010, 99950, 99840, 99810, 99840, 99870, 99870, 99820, 
    99820, 99830, 99840, 99820, 99840, 99870, 99910, 99920, 99950, 99960, 
    100000, 100050, 100070, 100100, 100120, 100140, 100150, 100170, 100200, 
    100220, 100240, 100270, 100290, 100290, 100310, 100320, 100330, 100400, 
    100410, 100380, 100340, 100350, 100310, 100310, 100390, 100470, 100480, 
    100490, 100470, 100460, 100440, 100450, 100460, 100470, 100460, 100430, 
    100490, 100520, 100520, 100550, 100530, 100500, 100520, 100530, 100550, 
    100500, 100530, 100610, 100650, 100700, 100710, 100730, 100730, 100740, 
    100730, 100760, 100760, 100760, 100780, 100790, 100770, 100770, 100810, 
    100890, 100900, 100970, 100950, 101010, 101010, 101060, 101080, 101060, 
    101070, 101090, 101110, 101140, 101210, 101210, 101120, 101090, 101090, 
    101110, 101120, 101120, 101150, 101170, 101180, 101200, 101190, 101170, 
    101180, 101170, 101150, 101150, 101110, 101110, 101120, 101100, 101110, 
    101150, 101140, 101170, 101180, 101170, 101140, 101130, 101130, 101170, 
    101240, 101250, 101260, 101270, 101270, 101280, 101320, 101310, 101320, 
    101310, 101320, 101320, 101310, 101350, 101360, 101370, 101350, 101370, 
    101390, 101380, 101370, 101360, 101390, 101390, 101410, 101420, 101480, 
    101530, 101530, 101520, 101530, 101550, 101610, 101660, 101650, 101680, 
    101730, 101780, 101810, 101840, 101850, 101880, 101910, 101920, 101910, 
    101940, 101950, 101970, 101950, 101970, 101980, 101990, 101970, 101910, 
    101890, 101860, 101760, 101740, 101690, 101650, 101620, 101580, 101540, 
    101560, 101500, 101420, 101410, 101380, 101360, 101330, 101320, 101300, 
    101340, 101430, 101470, 101410, 101390, 101400, 101470, 101510, 101510, 
    101550, 101550, 101560, 101590, 101620, 101660, 101660, 101720, 101780, 
    101810, 101870, 101840, 101860, 101900, 101930, 101950, 101970, 101980, 
    101960, 101990, 102030, 102020, 102020, 102020, 102020, 102000, 102020, 
    101990, 101960, 101960, 101930, 101930, 101930, 101910, 101880, 101820, 
    101800, 101790, 101740, 101740, 101680, 101650, 101620, 101620, 101610, 
    101600, 101550, 101510, 101510, 101490, 101490, 101480, 101500, 101520, 
    101530, 101490, 101480, 101450, 101430, 101410, 101370, 101340, 101340, 
    101330, 101340, 101310, 101280, 101240, 101180, 101170, 101160, 101160, 
    101140, 101120, 101090, 101120, 101160, 101190, 101190, 101210, 101240, 
    101270, 101250, 101280, 101300, 101280, 101310, 101330, 101350, 101320, 
    101350, 101310, 101290, 101270, 101240, 101260, 101260, 101260, 101240, 
    101210, 101180, 101160, 101170, 101180, 101180, 101150, 101120, 101150, 
    101120, 101100, 101090, 101050, 101010, 101000, 100920, 100810, 100820, 
    100770, 100640, 100620, 100600, 100520, 100430, 100430, 100390, 100300, 
    100220, 100200, 100170, 100210, 100210, 100170, 100160, 100130, 100130, 
    100030, 100030, 100180, 100190, 100160, 100140, 100090, 100030, 100040, 
    100000, 99930, 99840, 99820, 99810, 99770, 99730, 99660, 99570, 99510, 
    99450, 99390, 99390, 99370, 99250, 99310, 99290, 99280, 99180, 99100, 
    99080, 99050, 98970, 99010, 99050, 98990, 98990, 98940, 98990, 98980, 
    98970, 98960, 98990, 98940, 98940, 98930, 99000, 99060, 99100, 99170, 
    99230, 99290, 99310, 99410, 99470, 99510, 99540, 99610, 99660, 99720, 
    99770, 99830, 99890, 99940, 99990, 100020, 100050, 100070, 100110, 
    100120, 100120, 100150, 100160, 100210, 100240, 100290, 100310, 100310, 
    100310, 100310, 100290, 100280, 100310, 100290, 100310, 100330, 100340, 
    100350, 100320, 100310, 100300, 100310, 100310, 100310, 100330, 100330, 
    100340, 100340, 100350, 100350, 100320, 100280, 100250, 100250, 100230, 
    100220, 100190, 100180, 100110, 100070, 100070, 100040, 100020, 99970, 
    99920, 99860, 99790, 99740, 99700, 99640, 99560, 99490, 99410, 99400, 
    99370, 99330, 99340, 99330, 99270, 99260, 99260, 99230, 99220, 99220, 
    99210, 99250, 99260, 99240, 99260, 99270, 99260, 99290, 99310, 99350, 
    99400, 99430, 99460, 99500, 99520, 99540, 99560, 99570, 99600, 99630, 
    99650, 99650, 99660, 99680, 99690, 99690, 99720, 99750, 99740, 99740, 
    99740, 99760, 99790, 99810, 99850, 99900, 99950, 100010, 100070, 100120, 
    100140, 100180, 100230, 100260, 100290, 100310, 100370, 100400, 100400, 
    100410, 100500, 100540, 100540, 100550, 100590, 100630, 100680, 100710, 
    100700, 100720, 100750, 100780, 100830, 100840, 100850, 100870, 100880, 
    100870, 100860, 100880, 100890, 100880, 100860, 100870, 100820, 100750, 
    100760, 100800, 100790, 100780, 100770, 100740, 100750, 100710, 100700, 
    100690, 100700, 100700, 100700, 100700, 100710, 100720, 100720, 100690, 
    100660, 100670, 100680, 100720, 100730, 100730, 100760, 100770, 100770, 
    100790, 100790, 100790, 100820, 100840, 100850, 100880, 100910, 100870, 
    100890, 100940, 101000, 100990, 101020, 101020, 101060, 101070, 101080, 
    101090, 101130, 101110, 101070, 101130, 101140, 101180, 101190, 101220, 
    101260, 101300, 101280, 101320, 101360, 101400, 101460, 101490, 101450, 
    101450, 101480, 101490, 101530, 101550, 101550, 101550, 101570, 101570, 
    101570, 101570, 101590, 101610, 101590, 101580, 101620, 101650, 101670, 
    101690, 101720, 101730, 101700, 101730, 101740, 101750, 101720, 101740, 
    101740, 101780, 101780, 101750, 101750, 101720, 101710, 101660, 101650, 
    101620, 101560, 101520, 101510, 101530, 101510, 101510, 101560, 101510, 
    101540, 101540, 101540, 101520, 101550, 101530, 101550, 101540, 101540, 
    101550, 101530, 101510, 101490, 101490, 101480, 101480, 101470, 101450, 
    101440, 101460, 101460, 101460, 101440, 101440, 101440, 101430, 101420, 
    101420, 101410, 101400, 101400, 101410, 101410, 101420, 101420, 101410, 
    101420, 101420, 101420, 101430, 101430, 101450, 101450, 101480, 101500, 
    101510, 101520, 101530, 101530, 101540, 101530, 101530, 101530, 101520, 
    101530, 101540, 101550, 101580, 101590, 101580, 101590, 101590, 101600, 
    101590, 101600, 101610, 101610, 101630, 101670, 101670, 101640, 101660, 
    101670, 101640, 101620, 101600, 101560, 101520, 101500, 101500, 101480, 
    101440, 101420, 101380, 101370, 101350, 101310, 101290, 101270, 101250, 
    101220, 101200, 101160, 101120, 101110, 101090, 101070, 101050, 101030, 
    100980, 100950, 100930, 100910, 100900, 100900, 100890, 100870, 100860, 
    100840, 100850, 100840, 100840, 100820, 100820, 100830, 100830, 100850, 
    100890, 100890, 100850, 100890, 100910, 100910, 100870, 100870, 100880, 
    100890, 100890, 100930, 100960, 100980, 100990, 100980, 100980, 100980, 
    100970, 100990, 100980, 101000, 101000, 101030, 101060, 101090, 101110, 
    101130, 101100, 101140, 101140, 101130, 101100, 101110, 101120, 101110, 
    101090, 101060, 101040, 101060, 101060, 101080, 101060, 101040, 101030, 
    101050, 101050, 101050, 101030, 101030, 101050, 101050, 101060, 101040, 
    101010, 101010, 101030, 101070, 101090, 101140, 101170, 101200, 101250, 
    101270, 101310, 101340, 101360, 101350, 101370, 101430, 101460, 101490, 
    101500, 101570, 101590, 101640, 101680, 101710, 101730, 101740, 101730, 
    101740, 101780, 101830, 101840, 101880, 101930, 101970, 101970, 102000, 
    102010, 102050, 102050, 102060, 102060, 102120, 102180, 102250, 102250, 
    102280, 102290, 102310, 102320, 102320, 102350, 102370, 102390, 102390, 
    102410, 102410, 102410, 102410, 102420, 102420, 102420, 102430, 102450, 
    102480, 102500, 102510, 102510, 102500, 102480, 102500, 102490, 102490, 
    102480, 102480, 102480, 102480, 102480, 102480, 102480, 102470, 102470, 
    102440, 102420, 102430, 102420, 102420, 102410, 102410, 102420, 102430, 
    102430, 102420, 102420, 102410, 102420, 102400, 102360, 102340, 102310, 
    102310, 102320, 102330, 102330, 102330, 102320, 102310, 102300, 102300, 
    102290, 102260, 102250, 102250, 102280, 102290, 102300, 102270, 102270, 
    102260, 102240, 102210, 102190, 102180, 102200, 102220, 102230, 102260, 
    102290, 102290, 102290, 102320, 102350, 102370, 102370, 102380, 102420, 
    102450, 102480, 102510, 102520, 102540, 102540, 102490, 102550, 102560, 
    102570, 102550, 102590, 102640, 102640, 102670, 102650, 102640, 102620, 
    102640, 102570, 102540, 102430, 102450, 102360, 102180, 102210, 102100, 
    102120, 102040, 101960, 101790, 101540, 101470, 101340, 101180, 101130, 
    101010, 100960, 100860, 100680, 100550, 100490, 100440, 100410, 100390, 
    100370, 100340, 100370, 100360, 100350, 100380, 100450, 100490, 100530, 
    100560, 100580, 100620, 100640, 100660, 100670, 100690, 100710, 100740, 
    100760, 100760, 100770, 100770, 100750, 100750, 100720, 100720, 100710, 
    100660, 100660, 100620, 100620, 100570, 100530, 100490, 100460, 100460, 
    100430, 100420, 100410, 100430, 100420, 100460, 100440, 100500, 100530, 
    100580, 100630, 100720, 100800, 100880, 100980, 101060, 101190, 101310, 
    101390, 101460, 101490, 101520, 101570, 101620, 101630, 101650, 101650, 
    101640, 101650, 101640, 101610, 101590, 101550, 101520, 101480, 101400, 
    101360, 101310, 101250, 101160, 101120, 101080, 101040, 101000, 100990, 
    100980, 100970, 100950, 100950, 100950, 100940, 100970, 100970, 100970, 
    100920, 100930, 100900, 100950, 100960, 100950, 100930, 100940, 100940, 
    100940, 100930, 100900, 100860, 100830, 100780, 100760, 100730, 100700, 
    100680, 100690, 100660, 100610, 100600, 100570, 100520, 100470, 100440, 
    100470, 100440, 100420, 100360, 100320, 100310, 100350, 100410, 100480, 
    100530, 100540, 100600, 100640, 100670, 100720, 100720, 100780, 100820, 
    100860, 100930, 100970, 100940, 101090, 101100, 101150, 101190, 101260, 
    101300, 101320, 101340, 101400, 101460, 101500, 101560, 101570, 101630, 
    101690, 101730, 101780, 101820, 101850, 101870, 101900, 101940, 101960, 
    102010, 102020, 102040, 102040, 102050, 102090, 102100, 102120, 102140, 
    102150, 102190, 102190, 102200, 102200, 102220, 102230, 102240, 102270, 
    102260, 102270, 102280, 102270, 102270, 102270, 102260, 102270, 102280, 
    102280, 102250, 102240, 102230, 102240, 102250, 102240, 102250, 102250, 
    102260, 102280, 102310, 102330, 102350, 102360, 102370, 102380, 102380, 
    102420, 102460, 102500, 102480, 102500, 102480, 102500, 102510, 102500, 
    102490, 102500, 102520, 102530, 102560, 102550, 102550, 102570, 102590, 
    102580, 102590, 102580, 102570, 102550, 102560, 102570, 102560, 102550, 
    102550, 102550, 102540, 102530, 102520, 102500, 102490, 102480, 102460, 
    102460, 102460, 102460, 102430, 102410, 102390, 102370, 102370, 102340, 
    102320, 102290, 102260, 102260, 102250, 102220, 102200, 102170, 102130, 
    102120, 102080, 102050, 102020, 101990, 101980, 101950, 101940, 101910, 
    101860, 101810, 101790, 101750, 101710, 101660, 101620, 101580, 101540, 
    101510, 101460, 101450, 101430, 101400, 101350, 101320, 101280, 101250, 
    101210, 101210, 101200, 101180, 101170, 101170, 101190, 101200, 101200, 
    101210, 101220, 101220, 101210, 101210, 101210, 101220, 101240, 101280, 
    101270, 101290, 101330, 101340, 101350, 101340, 101350, 101370, 101380, 
    101400, 101420, 101440, 101460, 101480, 101490, 101510, 101510, 101510, 
    101490, 101500, 101500, 101500, 101510, 101520, 101500, 101490, 101480, 
    101460, 101480, 101460, 101430, 101460, 101440, 101430, 101430, 101420, 
    101410, 101390, 101370, 101370, 101380, 101370, 101350, 101330, 101310, 
    101280, 101260, 101260, 101270, 101280, 101290, 101300, 101260, 101240, 
    101230, 101230, 101250, 101280, 101310, 101340, 101380, 101400, 101470, 
    101510, 101550, 101600, 101610, 101670, 101700, 101710, 101740, 101780, 
    101800, 101780, 101770, 101770, 101770, 101780, 101920, 101950, 102000, 
    102040, 102090, 102110, 102160, 102220, 102280, 102310, 102340, 102330, 
    102350, 102370, 102380, 102400, 102430, 102440, 102460, 102450, 102470, 
    102460, 102500, 102500, 102500, 102520, 102530, 102550, 102510, 102530, 
    102550, 102550, 102580, 102580, 102600, 102590, 102590, 102540, 102550, 
    102590, 102590, 102580, 102540, 102540, 102530, 102550, 102570, 102540, 
    102550, 102540, 102560, 102550, 102580, 102580, 102600, 102630, 102640, 
    102650, 102630, 102640, 102650, 102650, 102670, 102690, 102700, 102710, 
    102720, 102750, 102750, 102760, 102770, 102770, 102770, 102780, 102790, 
    102810, 102840, 102850, 102850, 102860, 102860, 102860, 102850, 102850, 
    102850, 102830, 102840, 102840, 102870, 102880, 102870, 102860, 102870, 
    102860, 102870, 102860, 102840, 102830, 102840, 102860, 102860, 102850, 
    102860, 102850, 102830, 102830, 102810, 102770, 102750, 102730, 102710, 
    102700, 102700, 102710, 102680, 102650, 102610, 102590, 102570, 102540, 
    102510, 102460, 102430, 102410, 102410, 102400, 102390, 102340, 102290, 
    102260, 102230, 102190, 102150, 102110, 102090, 102040, 102030, 102000, 
    101960, 101890, 101830, 101780, 101690, 101620, 101530, 101480, 101440, 
    101380, 101270, 101210, 101100, 101110, 101100, 101060, 101000, 100940, 
    100890, 100830, 100780, 100730, 100690, 100680, 100640, 100600, 100570, 
    100540, 100520, 100540, 100500, 100560, 100590, 100600, 100610, 100660, 
    100720, 100760, 100770, 100800, 100850, 100900, 100940, 100950, 101000, 
    101050, 101090, 101130, 101190, 101230, 101240, 101280, 101300, 101330, 
    101350, 101410, 101460, 101480, 101530, 101550, 101620, 101670, 101700, 
    101740, 101780, 101830, 101860, 101890, 101910, 101920, 101950, 101990, 
    102010, 102030, 102060, 102080, 102100, 102110, 102140, 102110, 102140, 
    102170, 102190, 102220, 102200, 102250, 102260, 102260, 102280, 102280, 
    102300, 102290, 102290, 102280, 102270, 102260, 102280, 102310, 102300, 
    102290, 102260, 102260, 102250, 102230, 102190, 102150, 102090, 102060, 
    102000, 101950, 101890, 101810, 101720, 101640, 101570, 101450, 101380, 
    101330, 101270, 101250, 101230, 101200, 101200, 101180, 101140, 101120, 
    101120, 101070, 101020, 100990, 100990, 100990, 100970, 100950, 100910, 
    100910, 100890, 100870, 100880, 100870, 100840, 100860, 100880, 100920, 
    100930, 100920, 100900, 100920, 100920, 100900, 100880, 100890, 100880, 
    100870, 100880, 100880, 100880, 100890, 100870, 100870, 100870, 100880, 
    100880, 100870, 100870, 100870, 100840, 100850, 100840, 100830, 100810, 
    100800, 100780, 100750, 100700, 100680, 100670, 100680, 100640, 100620, 
    100580, 100510, 100470, 100390, 100310, 100220, 100120, 99990, 99910, 
    99790, 99670, 99580, 99460, 99340, 99260, 99140, 99020, 98920, 98830, 
    98730, 98640, 98590, 98530, 98470, 98390, 98300, 98230, 98130, 98030, 
    97920, 97820, 97680, 97550, 97430, 97310, 97150, 97090, 97020, 97000, 
    97000, 96990, 96990, 97000, 97000, 97050, 97120, 97200, 97280, 97330, 
    97450, 97500, 97590, 97720, 97890, 97910, 98050, 98100, 98130, 98280, 
    98350, 98420, 98520, 98590, 98660, 98770, 98830, 98890, 98930, 98980, 
    99060, 99130, 99220, 99320, 99400, 99450, 99490, 99510, 99550, 99610, 
    99640, 99650, 99650, 99660, 99660, 99670, 99710, 99740, 99730, 99700, 
    99670, 99710, 99690, 99680, 99720, 99750, 99790, 99810, 99830, 99840, 
    99920, 99930, 99930, 99900, 99890, 99870, 99850, 99950, 99990, 100030, 
    100040, 100070, 100140, 100180, 100260, 100310, 100360, 100390, 100420, 
    100420, 100500, 100550, 100620, 100650, 100700, 100750, 100790, 100830, 
    100880, 100950, 101020, 101080, 101090, 101120, 101170, 101230, 101270, 
    101280, 101290, 101330, 101370, 101380, 101440, 101490, 101520, 101550, 
    101560, 101590, 101620, 101640, 101640, 101650, 101670, 101680, 101700, 
    101720, 101720, 101730, 101730, 101750, 101770, 101780, 101770, 101750, 
    101760, 101760, 101780, 101810, 101830, 101830, 101810, 101820, 101800, 
    101790, 101800, 101780, 101760, 101780, 101790, 101810, 101800, 101810, 
    101800, 101800, 101790, 101810, 101830, 101850, 101860, 101910, 101930, 
    101930, 102010, 102020, 102030, 102050, 102060, 102060, 102070, 102060, 
    102050, 102030, 102020, 102070, 102090, 102120, 102140, 102130, 102180, 
    102190, 102180, 102170, 102150, 102120, 102150, 102140, 102130, 102130, 
    102110, 102100, 102120, 102150, 102140, 102160, 102120, 102150, 102130, 
    102060, 102010, 101960, 101910, 101870, 101840, 101780, 101720, 101700, 
    101640, 101600, 101600, 101620, 101630, 101670, 101680, 101690, 101700, 
    101710, 101730, 101770, 101750, 101770, 101830, 101880, 101880, 101930, 
    101880, 101890, 101910, 101920, 101910, 101960, 101960, 101940, 101990, 
    102010, 102030, 102010, 102030, 102040, 102060, 102070, 102070, 102100, 
    102060, 102070, 102100, 102110, 102150, 102170, 102170, 102180, 102180, 
    102190, 102190, 102180, 102190, 102210, 102200, 102210, 102170, 102130, 
    102060, 102030, 102050, 102030, 102010, 101970, 101930, 101910, 101910, 
    101910, 101850, 101800, 101820, 101830, 101830, 101800, 101780, 101760, 
    101740, 101680, 101640, 101660, 101650, 101690, 101600, 101680, 101720, 
    101730, 101710, 101730, 101720, 101710, 101740, 101740, 101740, 101780, 
    101780, 101790, 101790, 101830, 101820, 101810, 101810, 101820, 101870, 
    101880, 101910, 101930, 101930, 101960, 101970, 101990, 101990, 102010, 
    101990, 101990, 102000, 102030, 102020, 102020, 102010, 101980, 101970, 
    101950, 101950, 101930, 101890, 101890, 101900, 101890, 101890, 101880, 
    101870, 101870, 101860, 101840, 101820, 101770, 101740, 101710, 101700, 
    101710, 101700, 101680, 101650, 101640, 101650, 101630, 101620, 101590, 
    101580, 101540, 101510, 101540, 101540, 101550, 101580, 101570, 101580, 
    101550, 101550, 101550, 101530, 101520, 101540, 101520, 101540, 101540, 
    101540, 101520, 101520, 101520, 101520, 101520, 101530, 101550, 101560, 
    101590, 101580, 101580, 101590, 101590, 101610, 101620, 101630, 101640, 
    101640, 101660, 101680, 101700, 101730, 101710, 101730, 101750, 101790, 
    101810, 101820, 101840, 101850, 101870, 101910, 101950, 101990, 102020, 
    102030, 102060, 102020, 102050, 102020, 102050, 102050, 102100, 102100, 
    102140, 102170, 102180, 102210, 102210, 102220, 102230, 102260, 102300, 
    102290, 102240, 102250, 102320, 102280, 102310, 102310, 102310, 102300, 
    102270, 102270, 102250, 102200, 102220, 102220, 102180, 102210, 102150, 
    102090, 102040, 102010, 101950, 101940, 101880, 101830, 101780, 101730, 
    101700, 101720, 101670, 101630, 101570, 101540, 101530, 101520, 101560, 
    101580, 101600, 101580, 101590, 101600, 101610, 101620, 101640, 101660, 
    101650, 101690, 101700, 101760, 101730, 101770, 101830, 101830, 101860, 
    101850, 101860, 101860, 101860, 101850, 101850, 101830, 101810, 101800, 
    101800, 101790, 101770, 101770, 101770, 101750, 101740, 101710, 101690, 
    101670, 101640, 101650, 101680, 101670, 101650, 101660, 101650, 101670, 
    101680, 101670, 101680, 101700, 101710, 101740, 101750, 101790, 101820, 
    101860, 101860, 101860, 101880, 101890, 101920, 101930, 101940, 101960, 
    102000, 102020, 102040, 102060, 102090, 102080, 102090, 102100, 102100, 
    102090, 102070, 102090, 102100, 102100, 102090, 102050, 102050, 102020, 
    101970, 101940, 101930, 101910, 101870, 101870, 101870, 101860, 101870, 
    101870, 101850, 101830, 101810, 101810, 101770, 101730, 101720, 101680, 
    101630, 101600, 101550, 101520, 101510, 101490, 101500, 101470, 101450, 
    101450, 101420, 101400, 101390, 101360, 101340, 101310, 101310, 101310, 
    101280, 101240, 101190, 101210, 101210, 101210, 101190, 101160, 101110, 
    101120, 101120, 101110, 101110, 101100, 101080, 101100, 101100, 101090, 
    101090, 101070, 101060, 101050, 101040, 101010, 100980, 100960, 100930, 
    100920, 100880, 100870, 100850, 100820, 100780, 100710, 100650, 100620, 
    100580, 100530, 100510, 100490, 100480, 100480, 100470, 100460, 100450, 
    100460, 100450, 100440, 100420, 100430, 100410, 100400, 100390, 100410, 
    100410, 100400, 100390, 100360, 100350, 100350, 100350, 100340, 100330, 
    100330, 100350, 100350, 100360, 100380, 100410, 100440, 100440, 100470, 
    100470, 100480, 100480, 100480, 100470, 100480, 100490, 100500, 100500, 
    100500, 100470, 100460, 100460, 100440, 100430, 100420, 100410, 100370, 
    100360, 100360, 100340, 100310, 100270, 100250, 100240, 100210, 100210, 
    100190, 100200, 100200, 100180, 100180, 100190, 100210, 100240, 100250, 
    100260, 100270, 100300, 100320, 100350, 100380, 100410, 100460, 100480, 
    100520, 100530, 100580, 100610, 100630, 100650, 100680, 100750, 100760, 
    100800, 100850, 100880, 100890, 100920, 100960, 100980, 101020, 101040, 
    101080, 101090, 101110, 101170, 101170, 101180, 101200, 101210, 101220, 
    101220, 101200, 101210, 101200, 101190, 101160, 101160, 101130, 101090, 
    101090, 101080, 101060, 101010, 100960, 100930, 100910, 100900, 100870, 
    100860, 100820, 100770, 100740, 100700, 100680, 100660, 100630, 100620, 
    100600, 100600, 100610, 100610, 100630, 100640, 100650, 100660, 100670, 
    100680, 100690, 100690, 100740, 100770, 100810, 100850, 100870, 100890, 
    100910, 100960, 100970, 100990, 100990, 101040, 101080, 101100, 101110, 
    101150, 101140, 101170, 101200, 101220, 101240, 101290, 101310, 101290, 
    101310, 101340, 101360, 101370, 101390, 101390, 101390, 101410, 101400, 
    101390, 101370, 101310, 101280, 101240, 101240, 101190, 101110, 101090, 
    101030, 101020, 101030, 100980, 100860, 100820, 100780, 100780, 100790, 
    100790, 100790, 100820, 100780, 100780, 100810, 100820, 100850, 100850, 
    100840, 100850, 100890, 100880, 100920, 100910, 100910, 100950, 100960, 
    100970, 100980, 100970, 101010, 101020, 101030, 101060, 101070, 101090, 
    101120, 101130, 101120, 101120, 101140, 101170, 101190, 101190, 101200, 
    101190, 101200, 101220, 101210, 101200, 101210, 101190, 101190, 101200, 
    101210, 101170, 101160, 101180, 101200, 101210, 101210, 101200, 101220, 
    101220, 101210, 101220, 101230, 101250, 101270, 101270, 101300, 101330, 
    101330, 101330, 101350, 101370, 101400, 101430, 101430, 101450, 101480, 
    101500, 101530, 101540, 101570, 101580, 101590, 101640, 101660, 101670, 
    101680, 101690, 101700, 101730, 101770, 101770, 101780, 101800, 101820, 
    101820, 101840, 101850, 101870, 101880, 101890, 101910, 101950, 101950, 
    101960, 101980, 102000, 101990, 101980, 102000, 102010, 102030, 102040, 
    102050, 102080, 102080, 102040, 102090, 102100, 102140, 102170, 102170, 
    102200, 102240, 102280, 102310, 102330, 102370, 102420, 102430, 102460, 
    102490, 102510, 102500, 102500, 102500, 102490, 102490, 102510, 102490, 
    102480, 102510, 102470, 102470, 102420, 102400, 102360, 102320, 102290, 
    102250, 102190, 102140, 102090, 102020, 101960, 101860, 101800, 101700, 
    101650, 101530, 101510, 101480, 101380, 101310, 101240, 101210, 101150, 
    101120, 101080, 101030, 101070, 101040, 101060, 101050, 101060, 101090, 
    101080, 101100, 101090, 101090, 101100, 101070, 101090, 101090, 101100, 
    101100, 101090, 101100, 101090, 101090, 101100, 101080, 101080, 101080, 
    101060, 101050, 101050, 101040, 101040, 101010, 101000, 100950, 100900, 
    100800, 100720, 100640, 100540, 100440, 100330, 100280, 100240, 100220, 
    100160, 100170, 100160, 100110, 100080, 100040, 100040, 100040, 100000, 
    99990, 99950, 99890, 99870, 99950, 99950, 99960, 99900, 99880, 99870, 
    99890, 99950, 100010, 100040, 100090, 100140, 100150, 100180, 100210, 
    100220, 100230, 100280, 100310, 100350, 100400, 100420, 100450, 100460, 
    100490, 100510, 100520, 100520, 100540, 100570, 100570, 100590, 100620, 
    100640, 100660, 100670, 100670, 100680, 100680, 100680, 100700, 100720, 
    100730, 100820, 100860, 100880, 100900, 100930, 100940, 100950, 100930, 
    100910, 100960, 100970, 100990, 101010, 101080, 101080, 101070, 101130, 
    101150, 101170, 101170, 101140, 101170, 101160, 101170, 101180, 101200, 
    101190, 101190, 101210, 101220, 101210, 101150, 101100, 101060, 101060, 
    101020, 101020, 101000, 100980, 100950, 100950, 100920, 100900, 100870, 
    100840, 100840, 100850, 100850, 100890, 100920, 100930, 100940, 100960, 
    100990, 101010, 101020, 101030, 101040, 101070, 101100, 101100, 101120, 
    101150, 101140, 101150, 101150, 101160, 101130, 101100, 101110, 101120, 
    101100, 101110, 101090, 101080, 101090, 101070, 101030, 101030, 101010, 
    100980, 100950, 100950, 100970, 100960, 100940, 100920, 100890, 100870, 
    100830, 100840, 100820, 100800, 100770, 100730, 100710, 100680, 100650, 
    100640, 100630, 100630, 100590, 100530, 100500, 100470, 100430, 100390, 
    100420, 100410, 100410, 100430, 100420, 100430, 100420, 100410, 100380, 
    100340, 100330, 100360, 100400, 100400, 100400, 100380, 100390, 100390, 
    100410, 100410, 100400, 100410, 100410, 100420, 100430, 100440, 100460, 
    100470, 100470, 100460, 100470, 100460, 100490, 100500, 100510, 100520, 
    100550, 100560, 100570, 100610, 100640, 100670, 100700, 100700, 100720, 
    100730, 100760, 100770, 100800, 100820, 100820, 100820, 100820, 100820, 
    100820, 100820, 100800, 100790, 100770, 100820, 100810, 100810, 100850, 
    100850, 100840, 100860, 100860, 100920, 100930, 100950, 100970, 100980, 
    101000, 101020, 101040, 101040, 101060, 101080, 101080, 101080, 101100, 
    101140, 101130, 101130, 101170, 101210, 101240, 101280, 101320, 101340, 
    101380, 101420, 101420, 101460, 101460, 101490, 101530, 101530, 101560, 
    101570, 101600, 101590, 101560, 101590, 101580, 101560, 101550, 101590, 
    101620, 101640, 101640, 101610, 101580, 101570, 101590, 101580, 101560, 
    101520, 101510, 101500, 101490, 101430, 101390, 101350, 101300, 101240, 
    101230, 101200, 101080, 101070, 101040, 100980, 101040, 101000, 100910, 
    100880, 100840, 100830, 100760, 100660, 100680, 100650, 100620, 100590, 
    100590, 100520, 100470, 100430, 100410, 100370, 100300, 100250, 100230, 
    100170, 100120, 100010, 99970, 99960, 100030, 99870, 99850, 99830, 99840, 
    99890, 99900, 99910, 99850, 99860, 99790, 99750, 99800, 99720, 99630, 
    99620, 99540, 99640, 99530, 99550, 99470, 99500, 99500, 99460, 99480, 
    99540, 99510, 99570, 99540, 99540, 99580, 99580, 99590, 99580, 99540, 
    99490, 99500, 99500, 99490, 99480, 99510, 99540, 99590, 99620, 99660, 
    99720, 99780, 99830, 99880, 99930, 99980, 100030, 100060, 100080, 100110, 
    100130, 100120, 100120, 100130, 100130, 100120, 100110, 100050, 100050, 
    100010, 100000, 99990, 99920, 99840, 99830, 99830, 99850, 99870, 99890, 
    99900, 99920, 99910, 99940, 99970, 100000, 100020, 100040, 100080, 
    100090, 100110, 100110, 100110, 100140, 100120, 100130, 100140, 100150, 
    100160, 100160, 100160, 100180, 100240, 100250, 100300, 100340, 100360, 
    100350, 100380, 100420, 100410, 100470, 100490, 100540, 100580, 100600, 
    100620, 100620, 100630, 100630, 100650, 100660, 100670, 100680, 100700, 
    100730, 100750, 100760, 100790, 100790, 100810, 100840, 100850, 100840, 
    100860, 100870, 100860, 100880, 100900, 100910, 100910, 100910, 100900, 
    100910, 100920, 100940, 100950, 100940, 100940, 100950, 100940, 100960, 
    100960, 100970, 100970, 100960, 100960, 100960, 100970, 100960, 100980, 
    100980, 100990, 100990, 100980, 101000, 101010, 101000, 101010, 101000, 
    100990, 101020, 100990, 100970, 100970, 100920, 100900, 100910, 100880, 
    100840, 100800, 100770, 100770, 100680, 100600, 100520, 100450, 100410, 
    100320, 100220, 100170, 100120, 100050, 99970, 99940, 99900, 99900, 
    99920, 99930, 99960, 99980, 99990, 100000, 100020, 100080, 100060, 
    100200, 100330, 100410, 100420, 100520, 100550, 100620, 100660, 100690, 
    100700, 100620, 100590, 100650, 100700, 100700, 100700, 100710, 100760, 
    100870, 100920, 100990, 101040, 101090, 101090, 101140, 101170, 101200, 
    101170, 101150, 101140, 101210, 101230, 101270, 101230, 101280, 101310, 
    101320, 101330, 101330, 101370, 101400, 101390, 101410, 101370, 101380, 
    101410, 101410, 101380, 101370, 101360, 101350, 101370, 101320, 101290, 
    101290, 101310, 101270, 101230, 101180, 101160, 101130, 101120, 101080, 
    101050, 101030, 101030, 101010, 100980, 100950, 100920, 100880, 100850, 
    100830, 100790, 100750, 100710, 100670, 100630, 100590, 100550, 100500, 
    100490, 100490, 100470, 100410, 100390, 100380, 100430, 100430, 100420, 
    100410, 100410, 100410, 100400, 100390, 100390, 100350, 100350, 100340, 
    100330, 100330, 100340, 100340, 100320, 100310, 100290, 100290, 100260, 
    100260, 100250, 100270, 100280, 100270, 100270, 100280, 100260, 100260, 
    100260, 100260, 100250, 100250, 100190, 100190, 100160, 100190, 100210, 
    100190, 100240, 100240, 100220, 100220, 100200, 100200, 100190, 100200, 
    100200, 100190, 100180, 100190, 100180, 100160, 100150, 100140, 100110, 
    100110, 100100, 100090, 100100, 100090, 100100, 100110, 100100, 100090, 
    100110, 100100, 100080, 100080, 100090, 100090, 100130, 100140, 100150, 
    100170, 100180, 100190, 100190, 100210, 100190, 100220, 100230, 100240, 
    100270, 100290, 100340, 100360, 100360, 100370, 100370, 100380, 100410, 
    100420, 100470, 100510, 100560, 100570, 100600, 100630, 100660, 100650, 
    100660, 100660, 100650, 100630, 100630, 100600, 100570, 100550, 100520, 
    100500, 100480, 100460, 100440, 100400, 100400, 100350, 100340, 100310, 
    100340, 100370, 100380, 100380, 100400, 100430, 100480, 100540, 100520, 
    100540, 100570, 100500, 100580, 100640, 100600, 100640, 100660, 100680, 
    100700, 100680, 100670, 100680, 100670, 100670, 100660, 100660, 100640, 
    100650, 100640, 100610, 100580, 100590, 100590, 100570, 100540, 100530, 
    100520, 100510, 100510, 100460, 100410, 100360, 100330, 100300, 100250, 
    100200, 100180, 100140, 100090, 100070, 100000, 99950, 99880, 99830, 
    99780, 99730, 99680, 99590, 99540, 99500, 99460, 99420, 99400, 99380, 
    99370, 99340, 99310, 99280, 99270, 99280, 99290, 99310, 99340, 99370, 
    99420, 99460, 99490, 99510, 99550, 99590, 99640, 99700, 99730, 99770, 
    99830, 99910, 99990, 100070, 100140, 100220, 100280, 100320, 100400, 
    100420, 100500, 100560, 100630, 100680, 100670, 100750, 100830, 100860, 
    100910, 100940, 100900, 100940, 100950, 100960, 100990, 100990, 100990, 
    101020, 101020, 101000, 100970, 100990, 100980, 100980, 101000, 100990, 
    101020, 101040, 101050, 101050, 101060, 101040, 101030, 101050, 101060, 
    101070, 101090, 101110, 101120, 101130, 101170, 101200, 101280, 101310, 
    101370, 101420, 101470, 101500, 101490, 101510, 101520, 101580, 101650, 
    101650, 101770, 101810, 101760, 101770, 101730, 101730, 101750, 101740, 
    101730, 101770, 101780, 101780, 101770, 101730, 101710, 101690, 101670, 
    101670, 101660, 101680, 101690, 101720, 101710, 101740, 101710, 101700, 
    101710, 101660, 101780, 101800, 101850, 101850, 101870, 101850, 101810, 
    101800, 101770, 101740, 101720, 101690, 101670, 101640, 101610, 101580, 
    101570, 101550, 101520, 101500, 101490, 101470, 101470, 101450, 101430, 
    101430, 101390, 101380, 101400, 101420, 101420, 101390, 101430, 101420, 
    101400, 101380, 101380, 101380, 101360, 101360, 101360, 101370, 101380, 
    101380, 101370, 101390, 101360, 101340, 101350, 101320, 101300, 101360, 
    101330, 101340, 101340, 101400, 101460, 101490, 101530, 101560, 101590, 
    101610, 101660, 101650, 101700, 101720, 101750, 101790, 101780, 101810, 
    101790, 101780, 101810, 101830, 101840, 101850, 101790, 101800, 101800, 
    101810, 101790, 101750, 101690, 101650, 101590, 101550, 101530, 101490, 
    101400, 101360, 101330, 101290, 101250, 101170, 101100, 101030, 100960, 
    100830, 100730, 100570, 100460, 100290, 100180, 100060, 99990, 99860, 
    99750, 99690, 99670, 99750, 99760, 99750, 99740, 99710, 99700, 99690, 
    99680, 99650, 99640, 99570, 99480, 99450, 99410, 99340, 99300, 99270, 
    99260, 99220, 99230, 99290, 99300, 99330, 99370, 99390, 99450, 99450, 
    99540, 99560, 99550, 99510, 99510, 99420, 99440, 99470, 99470, 99450, 
    99440, 99440, 99440, 99480, 99520, 99520, 99430, 99510, 99540, 99570, 
    99590, 99610, 99640, 99680, 99690, 99720, 99740, 99750, 99740, 99760, 
    99770, 99770, 99730, 99710, 99690, 99670, 99680, 99710, 99730, 99770, 
    99820, 99870, 99930, 99980, 100020, 100040, 100080, 100140, 100170, 
    100200, 100260, 100280, 100280, 100300, 100360, 100400, 100430, 100510, 
    100620, 100660, 100710, 100740, 100880, 100950, 101010, 101070, 101100, 
    101150, 101180, 101210, 101230, 101280, 101310, 101350, 101390, 101420, 
    101430, 101430, 101430, 101440, 101450, 101460, 101480, 101480, 101480, 
    101510, 101520, 101540, 101550, 101560, 101580, 101580, 101560, 101550, 
    101570, 101590, 101600, 101620, 101620, 101620, 101630, 101650, 101640, 
    101640, 101630, 101650, 101660, 101690, 101730, 101770, 101790, 101810, 
    101830, 101860, 101870, 101880, 101890, 101930, 101960, 101980, 101990, 
    102010, 102050, 102060, 102060, 102090, 102090, 102090, 102100, 102120, 
    102130, 102150, 102160, 102190, 102190, 102190, 102170, 102180, 102170, 
    102170, 102170, 102190, 102190, 102190, 102200, 102210, 102230, 102200, 
    102220, 102230, 102230, 102220, 102200, 102190, 102190, 102190, 102150, 
    102150, 102150, 102160, 102110, 102130, 102060, 102030, 101980, 101960, 
    101940, 101910, 101910, 101860, 101840, 101870, 101910, 101960, 101980, 
    102030, 102080, 102090, 102120, 102160, 102180, 102210, 102250, 102260, 
    102250, 102240, 102220, 102240, 102270, 102200, 102180, 102160, 102110, 
    102050, 102000, 101950, 101900, 101810, 101750, 101630, 101580, 101520, 
    101500, 101450, 101420, 101370, 101370, 101330, 101310, 101310, 101320, 
    101310, 101340, 101390, 101420, 101440, 101480, 101490, 101540, 101560, 
    101570, 101590, 101530, 101560, 101520, 101490, 101480, 101500, 101530, 
    101550, 101570, 101600, 101640, 101650, 101670, 101660, 101640, 101610, 
    101570, 101510, 101450, 101390, 101240, 101170, 101090, 100960, 100970, 
    100920, 100820, 100740, 100680, 100590, 100540, 100500, 100470, 100400, 
    100300, 100280, 100260, 100240, 100190, 100190, 100280, 100270, 100310, 
    100320, 100340, 100380, 100390, 100400, 100400, 100410, 100430, 100450, 
    100470, 100490, 100500, 100550, 100580, 100580, 100580, 100600, 100570, 
    100530, 100500, 100470, 100440, 100390, 100350, 100300, 100220, 100100, 
    99970, 99840, 99750, 99670, 99580, 99540, 99560, 99560, 99560, 99570, 
    99590, 99600, 99600, 99620, 99620, 99640, 99670, 99670, 99670, 99690, 
    99740, 99730, 99740, 99740, 99720, 99760, 99740, 99720, 99690, 99650, 
    99610, 99560, 99490, 99500, 99470, 99440, 99450, 99420, 99390, 99370, 
    99350, 99310, 99280, 99250, 99210, 99150, 99150, 99140, 99130, 99120, 
    99090, 99100, 99100, 99080, 99070, 99060, 99040, 99030, 99040, 99010, 
    98980, 98980, 99010, 99020, 99030, 99050, 99070, 99100, 99130, 99170, 
    99200, 99260, 99300, 99340, 99360, 99370, 99390, 99420, 99400, 99420, 
    99420, 99430, 99430, 99410, 99400, 99370, 99350, 99360, 99380, 99400, 
    99440, 99450, 99480, 99530, 99570, 99590, 99610, 99600, 99550, 99570, 
    99550, 99550, 99570, 99530, 99550, 99580, 99540, 99530, 99580, 99580, 
    99600, 99620, 99590, 99580, 99640, 99680, 99710, 99750, 99760, 99740, 
    99730, 99700, 99750, 99700, 99780, 99920, 99930, 99920, 99930, 99900, 
    99930, 99940, 99920, 99910, 99920, 99920, 99910, 99900, 99890, 99900, 
    99900, 99920, 99920, 99920, 99950, 99940, 99940, 99950, 99960, 99950, 
    99960, 99990, 100000, 99980, 100020, 100010, 100030, 100030, 99990, 
    100050, 100060, 100030, 100070, 100140, 100190, 100230, 100260, 100290, 
    100320, 100370, 100390, 100440, 100470, 100490, 100500, 100530, 100570, 
    100590, 100620, 100640, 100680, 100690, 100720, 100750, 100780, 100790, 
    100800, 100810, 100840, 100880, 100910, 100960, 100980, 101010, 101030, 
    101050, 101050, 101080, 101110, 101150, 101170, 101200, 101210, 101270, 
    101290, 101320, 101300, 101340, 101340, 101340, 101360, 101370, 101370, 
    101380, 101370, 101340, 101330, 101290, 101280, 101280, 101270, 101280, 
    101280, 101280, 101300, 101300, 101280, 101260, 101270, 101270, 101250, 
    101310, 101350, 101370, 101390, 101390, 101410, 101420, 101430, 101460, 
    101450, 101450, 101450, 101440, 101420, 101400, 101360, 101340, 101320, 
    101310, 101310, 101360, 101340, 101310, 101290, 101240, 101230, 101210, 
    101210, 101250, 101220, 101220, 101230, 101240, 101220, 101230, 101210, 
    101170, 101190, 101100, 101090, 101010, 101020, 100990, 100930, 100880, 
    100790, 100820, 100730, 100580, 100490, 100500, 100480, 100370, 100230, 
    100160, 100110, 100020, 100010, 100000, 99980, 99930, 99840, 99800, 
    99770, 99750, 99750, 99730, 99660, 99590, 99590, 99630, 99710, 99760, 
    99750, 99810, 99890, 99910, 99950, 100020, 100060, 100100, 100110, 
    100110, 100130, 100080, 100050, 100020, 100040, 100040, 100030, 100010, 
    100010, 100090, 100120, 100130, 100160, 100160, 100210, 100170, 100240, 
    100230, 100240, 100310, 100350, 100390, 100440, 100440, 100440, 100490, 
    100550, 100650, 100720, 100770, 100830, 100880, 100890, 100940, 100970, 
    101040, 101050, 101090, 101110, 101140, 101190, 101190, 101200, 101210, 
    101240, 101260, 101280, 101170, 101080, 101150, 101160, 101340, 101360, 
    101400, 101440, 101470, 101490, 101510, 101550, 101540, 101560, 101530, 
    101440, 101510, 101540, 101630, 101600, 101590, 101630, 101640, 101660, 
    101660, 101850, 101870, 101780, 101750, 101740, 101740, 101780, 101710, 
    101730, 101790, 101790, 101810, 101800, 101770, 101730, 101710, 101680, 
    101660, 101640, 101620, 101570, 101560, 101570, 101560, 101540, 101510, 
    101470, 101430, 101420, 101400, 101380, 101330, 101330, 101280, 101250, 
    101220, 101200, 101170, 101150, 101100, 101080, 101040, 101000, 100940, 
    100890, 100880, 100790, 100770, 100730, 100680, 100530, 100440, 100420, 
    100380, 100330, 100300, 100210, 100140, 100010, 99950, 99900, 99840, 
    99740, 99690, 99760, 99740, 99740, 99720, 99710, 99710, 99700, 99710, 
    99740, 99800, 99780, 99830, 99870, 99930, 99960, 100020, 100080, 100130, 
    100150, 100210, 100270, 100330, 100390, 100440, 100490, 100530, 100590, 
    100670, 100730, 100790, 100810, 100870, 100920, 101010, 101060, 101100, 
    101150, 101210, 101280, 101330, 101380, 101410, 101450, 101480, 101550, 
    101600, 101660, 101710, 101750, 101790, 101840, 101910, 101940, 101980, 
    102010, 102040, 102050, 102090, 102130, 102160, 102160, 102190, 102210, 
    102220, 102220, 102240, 102230, 102210, 102210, 102190, 102180, 102150, 
    102120, 102070, 102060, 102050, 102010, 101970, 101920, 101880, 101830, 
    101770, 101700, 101620, 101550, 101520, 101480, 101480, 101450, 101410, 
    101400, 101400, 101400, 101360, 101330, 101300, 101290, 101260, 101240, 
    101240, 101230, 101200, 101180, 101150, 101130, 101090, 101060, 101020, 
    100980, 100920, 100880, 100830, 100800, 100740, 100700, 100670, 100620, 
    100580, 100540, 100520, 100510, 100510, 100510, 100500, 100510, 100500, 
    100500, 100500, 100480, 100470, 100460, 100460, 100450, 100430, 100410, 
    100410, 100430, 100420, 100420, 100410, 100390, 100390, 100370, 100360, 
    100330, 100320, 100300, 100310, 100330, 100350, 100370, 100410, 100410, 
    100390, 100370, 100390, 100390, 100420, 100450, 100460, 100460, 100480, 
    100490, 100480, 100470, 100490, 100460, 100490, 100500, 100540, 100540, 
    100580, 100600, 100620, 100640, 100660, 100670, 100680, 100670, 100690, 
    100690, 100690, 100700, 100700, 100710, 100700, 100720, 100700, 100700, 
    100680, 100660, 100660, 100650, 100650, 100650, 100650, 100670, 100670, 
    100670, 100690, 100700, 100700, 100700, 100710, 100710, 100720, 100730, 
    100740, 100750, 100760, 100760, 100770, 100790, 100800, 100820, 100820, 
    100840, 100860, 100890, 100930, 100950, 100950, 100960, 100970, 100980, 
    100990, 101000, 101000, 101020, 101030, 101030, 101040, 101070, 101070, 
    101080, 101090, 101110, 101130, 101120, 101160, 101180, 101180, 101200, 
    101230, 101250, 101270, 101280, 101280, 101310, 101300, 101290, 101290, 
    101310, 101290, 101290, 101290, 101270, 101240, 101200, 101190, 101230, 
    101210, 101200, 101140, 101160, 101170, 101180, 101230, 101200, 101270, 
    101280, 101210, 101210, 101190, 101200, 101200, 101210, 101190, 101180, 
    101170, 101180, 101190, 101250, 101290, 101300, 101320, 101330, 101360, 
    101370, 101320, 101350, 101340, 101410, 101440, 101440, 101460, 101440, 
    101430, 101430, 101430, 101400, 101380, 101370, 101370, 101360, 101330, 
    101320, 101310, 101270, 101280, 101250, 101220, 101190, 101160, 101140, 
    101150, 101150, 101140, 101130, 101100, 101080, 101030, 100990, 100960, 
    100950, 100900, 100890, 100850, 100850, 100820, 100790, 100710, 100650, 
    100600, 100590, 100550, 100510, 100450, 100420, 100410, 100370, 100370, 
    100360, 100330, 100300, 100290, 100310, 100320, 100340, 100340, 100330, 
    100360, 100470, 100520, 100560, 100620, 100670, 100710, 100760, 100840, 
    100910, 100980, 101060, 101120, 101150, 101230, 101270, 101310, 101380, 
    101400, 101440, 101480, 101510, 101540, 101580, 101610, 101620, 101640, 
    101650, 101660, 101660, 101680, 101680, 101670, 101680, 101690, 101710, 
    101720, 101740, 101750, 101740, 101740, 101750, 101750, 101760, 101770, 
    101780, 101780, 101810, 101820, 101830, 101830, 101840, 101830, 101830, 
    101830, 101830, 101820, 101810, 101770, 101780, 101770, 101800, 101780, 
    101780, 101780, 101750, 101760, 101750, 101710, 101660, 101630, 101580, 
    101530, 101490, 101460, 101420, 101400, 101400, 101380, 101330, 101280, 
    101290, 101300, 101300, 101320, 101330, 101330, 101280, 101250, 101220, 
    101210, 101190, 101220, 101240, 101240, 101240, 101210, 101230, 101240, 
    101240, 101250, 101280, 101290, 101300, 101340, 101360, 101400, 101440, 
    101470, 101490, 101520, 101550, 101550, 101590, 101600, 101600, 101610, 
    101610, 101630, 101630, 101630, 101630, 101600, 101610, 101630, 101610, 
    101590, 101560, 101530, 101520, 101510, 101490, 101510, 101520, 101540, 
    101570, 101600, 101650, 101770, 101870, 101940, 102010, 102090, 102240, 
    102350, 102390, 102530, 102650, 102740, 102780, 102860, 102960, 103020, 
    103070, 103130, 103210, 103250, 103320, 103340, 103340, 103360, 103380, 
    103390, 103380, 103350, 103330, 103320, 103300, 103270, 103220, 103220, 
    103200, 103140, 103090, 103050, 103020, 102990, 102940, 102900, 102830, 
    102760, 102710, 102660, 102600, 102510, 102460, 102400, 102330, 102280, 
    102260, 102240, 102250, 102290, 102340, 102380, 102420, 102380, 102450, 
    102480, 102500, 102500, 102500, 102530, 102520, 102520, 102430, 102380, 
    102370, 102330, 102280, 102230, 102160, 102140, 102130, 102110, 102100, 
    102080, 102070, 102070, 102050, 102010, 101970, 101990, 101980, 101950, 
    101920, 101910, 101880, 101870, 101870, 101880, 101890, 101840, 101820, 
    101810, 101810, 101820, 101820, 101800, 101800, 101790, 101770, 101780, 
    101770, 101750, 101720, 101730, 101710, 101710, 101700, 101720, 101730, 
    101740, 101760, 101780, 101780, 101780, 101760, 101760, 101730, 101690, 
    101680, 101650, 101640, 101610, 101550, 101510, 101480, 101380, 101290, 
    101270, 101290, 101290, 101270, 101220, 101170, 101200, 101210, 101190, 
    101160, 101120, 101160, 101150, 101140, 101110, 101080, 101060, 101050, 
    100970, 101030, 100990, 100960, 100960, 100940, 100910, 100840, 100780, 
    100740, 100690, 100650, 100600, 100550, 100510, 100500, 100450, 100410, 
    100350, 100290, 100260, 100190, 100120, 100090, 100020, 100000, 99960, 
    99900, 99860, 99830, 99790, 99770, 99750, 99710, 99700, 99790, 99830, 
    99770, 99890, 99950, 99940, 99870, 99910, 99950, 99930, 99960, 100010, 
    100060, 100120, 100140, 100150, 100290, 100350, 100380, 100400, 100430, 
    100450, 100470, 100530, 100610, 100670, 100750, 100810, 100840, 100910, 
    100930, 100980, 101050, 101080, 101100, 101150, 101160, 101180, 101220, 
    101230, 101240, 101240, 101250, 101260, 101280, 101300, 101310, 101330, 
    101360, 101360, 101370, 101380, 101370, 101360, 101370, 101360, 101340, 
    101320, 101320, 101310, 101300, 101300, 101270, 101260, 101230, 101210, 
    101180, 101150, 101130, 101120, 101080, 101090, 101080, 101040, 101010, 
    101000, 100960, 100900, 100850, 100810, 100740, 100660, 100590, 100500, 
    100430, 100350, 100280, 100190, 100090, 100000, 99910, 99840, 99770, 
    99680, 99660, 99660, 99620, 99590, 99560, 99500, 99540, 99530, 99540, 
    99550, 99540, 99560, 99550, 99550, 99580, 99600, 99640, 99590, 99600, 
    99640, 99630, 99600, 99560, 99530, 99540, 99530, 99540, 99540, 99550, 
    99540, 99530, 99560, 99600, 99600, 99630, 99670, 99760, 99890, 99980, 
    100080, 100120, 100230, 100350, 100450, 100540, 100650, 100690, 100750, 
    100810, 100900, 100970, 101030, 101070, 101090, 101080, 101050, 101000, 
    100950, 100880, 100820, 100730, 100690, 100680, 100650, 100670, 100690, 
    100730, 100740, 100770, 100750, 100750, 100760, 100750, 100740, 100750, 
    100750, 100780, 100760, 100750, 100750, 100810, 100780, 100780, 100780, 
    100720, 100740, 100760, 100750, 100830, 100840, 100860, 100870, 100890, 
    100870, 100840, 100810, 100800, 100810, 100850, 100870, 100900, 100910, 
    100920, 100930, 100940, 100950, 100960, 100960, 100940, 100940, 100970, 
    100940, 100940, 100940, 100890, 100820, 100780, 100750, 100720, 100670, 
    100630, 100600, 100630, 100630, 100620, 100610, 100620, 100620, 100580, 
    100580, 100580, 100580, 100580, 100580, 100600, 100610, 100620, 100640, 
    100630, 100660, 100700, 100690, 100710, 100700, 100680, 100700, 100730, 
    100760, 100790, 100800, 100840, 100840, 100870, 100850, 100870, 100900, 
    100940, 100980, 101030, 101070, 101500, 101530, 101560, 101580, 101610, 
    101630, 101640, 101660, 101690, 101710, 101720, 101760, 101790, 101790, 
    101790, 101800, 101810, 101780, 101810, 101810, 101820, 101850, 101850, 
    101890, 101880, 101880, 101860, 101850, 101820, 101800, 101790, 101750, 
    101730, 101700, 101650, 101650, 101600, 101490, 101310, 101240, 101180, 
    101140, 101170, 101200, 101190, 101210, 101270, 101330, 101380, 101410, 
    101430, 101490, 101520, 101580, 101640, 101700, 101780, 101840, 101900, 
    101980, 102020, 102080, 102090, 102160, 102190, 102230, 102280, 102310, 
    102350, 102380, 102410, 102440, 102470, 102480, 102470, 102450, 102440, 
    102430, 102430, 102420, 102380, 102370, 102330, 102310, 102270, 102250, 
    102210, 102160, 102110, 102050, 102010, 102000, 101950, 101890, 101840, 
    101800, 101760, 101700, 101620, 101510, 101400, 101290, 101210, 101120, 
    101020, 100920, 100820, 100700, 100580, 100480, 100360, 100240, 100170, 
    100080, 100040, 99990, 99940, 99920, 99880, 99850, 99840, 99780, 99710, 
    99640, 99580, 99500, 99400, 99320, 99230, 99110, 99020, 98930, 98880, 
    98820, 98770, 98750, 98740, 98730, 98740, 98760, 98730, 98730, 98730, 
    98740, 98750, 98750, 98770, 98770, 98800, 98870, 98950, 99050, 99130, 
    99210, 99260, 99310, 99350, 99330, 99290, 99310, 99330, 99320, 99280, 
    99280, 99210, 99160, 99080, 99020, 98950, 98810, 98680, 98620, 98540, 
    98510, 98390, 98390, 98350, 98360, 98390, 98390, 98430, 98460, 98520, 
    98580, 98640, 98730, 98790, 98890, 98920, 98990, 99050, 99120, 99170, 
    99200, 99210, 99230, 99200, 99220, 99260, 99230, 99190, 99180, 99140, 
    99110, 99080, 99050, 98950, 98880, 98820, 98760, 98690, 98670, 98560, 
    98550, 98500, 98480, 98500, 98480, 98440, 98450, 98440, 98430, 98460, 
    98490, 98530, 98570, 98630, 98700, 98750, 98780, 98800, 98840, 98870, 
    98890, 98940, 98950, 98980, 98990, 99030, 99070, 99080, 99120, 99150, 
    99170, 99200, 99240, 99260, 99270, 99340, 99420, 99440, 99500, 99560, 
    99640, 99720, 99760, 99830, 99880, 99940, 100010, 100090, 100150, 100200, 
    100250, 100300, 100300, 100330, 100340, 100330, 100350, 100340, 100360, 
    100350, 100370, 100340, 100350, 100360, 100360, 100340, 100360, 100380, 
    100420, 100460, 100500, 100540, 100570, 100620, 100660, 100690, 100690, 
    100670, 100660, 100620, 100560, 100540, 100520, 100500, 100480, 100470, 
    100440, 100420, 100390, 100370, 100320, 100310, 100300, 100280, 100250, 
    100250, 100260, 100240, 100210, 100230, 100190, 100190, 100120, 100160, 
    100100, 100150, 100200, 100190, 100170, 100070, 99980, 100020, 100030, 
    100020, 100020, 100000, 99990, 99950, 99980, 100000, 100020, 100050, 
    100040, 100050, 100070, 100100, 100100, 100140, 100180, 100210, 100240, 
    100280, 100310, 100370, 100440, 100500, 100570, 100610, 100600, 100670, 
    100640, 100700, 100700, 100760, 100820, 100780, 100820, 100840, 100830, 
    100830, 100830, 100790, 100760, 100720, 100670, 100640, 100630, 100600, 
    100590, 100550, 100540, 100540, 100530, 100510, 100500, 100480, 100460, 
    100460, 100470, 100480, 100480, 100470, 100470, 100460, 100460, 100460, 
    100480, 100480, 100490, 100490, 100500, 100530, 100540, 100550, 100530, 
    100530, 100540, 100540, 100550, 100530, 100520, 100490, 100540, 100590, 
    100580, 100590, 100600, 100580, 100560, 100640, 100660, 100670, 100680, 
    100650, 100610, 100550, 100490, 100510, 100580, 100550, 100540, 100590, 
    100600, 100640, 100700, 100730, 100760, 100780, 100830, 100850, 100870, 
    100890, 100890, 100900, 100890, 100860, 100850, 100850, 100880, 100890, 
    100880, 100860, 100860, 100840, 100820, 100810, 100800, 100780, 100740, 
    100730, 100720, 100720, 100710, 100680, 100660, 100650, 100620, 100610, 
    100590, 100570, 100550, 100530, 100520, 100510, 100500, 100480, 100470, 
    100440, 100410, 100420, 100420, 100400, 100400, 100390, 100380, 100390, 
    100390, 100390, 100390, 100400, 100430, 100440, 100470, 100490, 100520, 
    100530, 100570, 100600, 100640, 100650, 100680, 100670, 100660, 100670, 
    100720, 100730, 100750, 100780, 100820, 100850, 100870, 100890, 100930, 
    100920, 100890, 100890, 100910, 100900, 100910, 100930, 100940, 100950, 
    100970, 100980, 101020, 101010, 101050, 101080, 101090, 101140, 101160, 
    101170, 101180, 101240, 101270, 101300, 101310, 101310, 101290, 101260, 
    101230, 101200, 101210, 101150, 101100, 101130, 101120, 101110, 101090, 
    101060, 101040, 101020, 101000, 100990, 100980, 100980, 101020, 101040, 
    101110, 101130, 101150, 101140, 101140, 101150, 101150, 101190, 101230, 
    101230, 101230, 101260, 101290, 101380, 101420, 101450, 101490, 101510, 
    101520, 101530, 101540, _, 101510, 101550, 101600, 101640, 101680, 
    101750, 101770, 101770, 101810, 101800, 101830, 101910, 101940, 102010, 
    102110, 102180, 102240, 102300, 102350, 102410, 102430, 102450, 102470, 
    102480, 102490, 102550, 102640, 102680, 102760, 102810, 102880, 102860, 
    102910, 102930, 102930, 102950, 102990, 103020, 103080, 103090, 103110, 
    103120, 103140, 103160, 103140, 103150, 103130, 103160, 103180, 103230, 
    103260, 103290, 103280, 103280, 103280, 103290, 103310, 103310, 103350, 
    103390, 103420, 103460, 103480, 103510, 103500, 103520, 103550, 103600, 
    103640, 103690, 103720, 103750, 103790, 103820, 103880, 103920, 103940, 
    103940, 103950, 103940, 103980, 103960, 103960, 103980, 103980, 103920, 
    103880, 103950, 103970, 103930, 103910, 103870, 103810, 103780, 103610, 
    103630, 103590, 103620, 103630, 103630, 103630, 103610, 103600, 103620, 
    103620, 103630, 103640, 103650, 103650, 103650, 103650, 103670, 103640, 
    103620, 103610, 103630, 103660, 103670, 103660, 103690, 103710, 103720, 
    103750, 103740, 103750, 103790, 103810, 103830, 103820, 103850, 103830, 
    103830, 103780, 103780, 103780, 103780, 103780, 103750, 103730, 103730, 
    103710, 103710, 103710, 103720, 103720, 103740, 103750, 103760, 103750, 
    103740, 103760, 103770, 103790, 103810, 103800, 103810, 103830, 103860, 
    103870, 103920, 103950, 104000, 103990, 103990, 104010, 104000, 104030, 
    104010, 104030, 104050, 104070, 104100, 104120, 104120, 104090, 104080, 
    104070, 104020, 103990, 103950, 103920, 103890, 103860, 103820, 103770, 
    103740, 103700, 103660, 103610, 103570, 103540, 103490, 103430, 103360, 
    103330, 103290, 103270, 103220, 103160, 103110, 103050, 103040, 103010, 
    102980, 102950, 102930, 102940, 102890, 102880, 102840, 102810, 102760, 
    102750, 102720, 102670, 102670, 102650, 102680, 102690, 102670, 102680, 
    102680, 102670, 102640, 102620, 102590, 102580, 102570, 102560, 102550, 
    102580, 102580, 102580, 102550, 102520, 102490, 102450, 102450, 102450, 
    102450, 102450, 102450, 102450, 102460, 102450, 102410, 102420, 102390, 
    102370, 102330, 102320, 102300, 102290, 102270, 102280, 102260, 102210, 
    102190, 102160, 102130, 102100, 102110, 102090, 102040, 102020, 102020, 
    102030, 102010, 102010, 101960, 101910, 101840, 101770, 101710, 101660, 
    101630, 101580, 101530, 101500, 101480, 101470, 101430, 101420, 101390, 
    101360, 101350, 101350, 101350, 101370, 101400, 101380, 101370, 101370, 
    101400, 101390, 101360, 101350, 101320, 101320, 101270, 101260, 101260, 
    101230, 101180, 101160, 101090, 101060, 101010, 100990, 100980, 100960, 
    100980, 100980, 100980, 101040, 101070, 101140, 101140, 101150, 101160, 
    101210, 101240, 101280, 101300, 101310, 101350, 101370, 101400, 101440, 
    101470, 101470, 101500, 101460, 101520, 101540, 101560, 101610, 101660, 
    101730, 101800, 101790, 101820, 101870, 101900, 101950, 101970, 102050, 
    102120, 102200, 102270, 102360, 102360, 102420, 102460, 102530, 102590, 
    102630, 102700, 102770, 102870, 102950, 103020, 103080, 103130, 103170, 
    103200, 103250, 103290, 103350, 103390, 103450, 103480, 103500, 103550, 
    103580, 103580, 103580, 103540, 103470, 103380, 103380, 103310, 103220, 
    103140, 103040, 102900, 102820, 102670, 102490, 102370, 102310, 102280, 
    102280, 102290, 102310, 102330, 102320, 102320, 102300, 102320, 102330, 
    102290, 102280, 102330, 102380, 102370, 102390, 102450, 102500, 102540, 
    102600, 102670, 102700, 102740, 102770, 102760, 102790, 102810, 102860, 
    102850, 102860, 102900, 102940, 102940, 102950, 102980, 102990, 102990, 
    102970, 103010, 102990, 103070, 103110, 103190, 103230, 103290, 103330, 
    103390, 103410, 103420, 103410, 103430, 103460, 103460, 103470, 103480, 
    103480, 103480, 103480, 103450, 103400, 103350, 103360, 103320, 103260, 
    103200, 103170, 103130, 103100, 103070, 103040, 102970, 102900, 102840, 
    102720, 102670, 102640, 102590, 102530, 102480, 102460, 102390, 102340, 
    102290, 102270, 102240, 102200, 102180, 102140, 102120, 102080, 102080, 
    102090, 102070, 102030, 102000, 102000, 101950, 101910, 101880, 101880, 
    101860, 101860, 101880, 101860, 101860, 101850, 101860, 101890, 101900, 
    101930, 101940, 101970, 101970, 102010, 102050, 102090, 102090, 102110, 
    102130, 102130, 102100, 102050, 102030, 101980, 101920, 101880, 101840, 
    101760, 101640, 101530, 101420, 101410, 101370, 101290, 101220, 101180, 
    101120, 101030, 100930, 100850, 100820, 100740, 100620, 100540, 100480, 
    100420, 100350, 100290, 100260, 100250, 100230, 100210, 100210, 100220, 
    100220, 100220, 100190, 100160, 100110, 100130, 100160, 100200, 100270, 
    100290, 100410, 100670, 100780, 100940, 101060, 101220, 101330, 101430, 
    101580, 101680, 101790, 101870, 101960, 102010, 102040, 102080, 102100, 
    102150, 102160, 102190, 102260, 102310, 102370, 102430, 102490, 102540, 
    102610, 102670, 102740, 102820, 102890, 102930, 102980, 103050, 103090, 
    103150, 103180, 103210, 103230, 103220, 103230, 103220, 103200, 103140, 
    103050, 102980, 102900, 102790, 102670, 102560, 102430, 102250, 102060, 
    101830, 101670, 101510, 101340, 101140, 101120, 101090, 101050, 101080, 
    101160, 101220, 101210, 101280, 101390, 101530, 101690, 101820, 102000, 
    102140, 102270, 102410, 102460, 102530, 102650, 102710, 102770, 102820, 
    102870, 102890, 102920, 102940, 102920, 102910, 102920, 102940, 102950, 
    102970, 102990, 103030, 103030, 103050, 103100, 103130, 103150, 103170, 
    103170, 103190, 103220, 103190, 103070, 103050, 102900, 102830, 102720, 
    102550, 102400, 102220, 101900, 101600, 101360, 101160, 100970, 100710, 
    100340, 100160, 100090, 100030, 99970, 99930, 99840, 99780, 99700, 99620, 
    99570, 99540, 99550, 99500, 99460, 99370, 99290, 99240, 99230, 99270, 
    99260, 99280, 99370, 99710, 99990, 100230, 100520, 100720, 100920, 
    101140, 101260, 101310, 101380, 101710, 101890, 101840, 101990, 102130, 
    102230, 102270, 102320, 102320, 102320, 102350, 102340, 102310, 102280, 
    102220, 102170, 102110, 102050, 101980, 101870, 101750, 101620, 101480, 
    101320, 101140, 100990, 100810, 100670, 100580, 100500, 100430, 100380, 
    100260, 100180, 100080, 99990, 99890, 99790, 99680, 99570, 99490, 99420, 
    99390, 99340, 99320, 99290, 99260, 99260, 99250, 99290, 99300, 99310, 
    99310, 99380, 99420, 99450, 99470, 99470, 99470, 99460, 99430, 99450, 
    99420, 99410, 99420, 99460, 99460, 99490, 99540, 99510, 99510, 99540, 
    99510, 99480, 99430, 99360, 99300, 99280, 99300, 99310, 99250, 99190, 
    99110, 99020, 98940, 98720, 98490, 98320, 97810, 97680, 97640, 97560, 
    97450, 97450, 97480, 97720, 97980, 98360, 98550, 98700, 98880, 99000, 
    99100, 99170, 99200, 99210, 99250, 99300, 99320, 99350, 99390, 99430, 
    99430, 99510, 99570, 99620, 99650, 99640, 99660, 99710, 99780, 99850, 
    99890, 99940, 100000, 100060, 100110, 100180, 100240, 100310, 100360, 
    100400, 100500, 100540, 100590, 100660, 100740, 100740, 100780, 100790, 
    100780, 100610, 100580, 100600, 100620, 100610, 100630, 100650, 100690, 
    100700, 100780, 100820, 100830, 100790, 100770, 100790, 100780, 100790, 
    100770, 100810, 100760, 100800, 100780, 100780, 100760, 100750, 100720, 
    100710, 100700, 100640, 100840, 100880, 100910, 100970, 101020, 101070, 
    101100, 101140, 101170, 101160, 101160, 101180, 101170, 101180, 101160, 
    101180, 101170, 101210, 101190, 101200, 101170, 101100, 101080, 101080, 
    101100, 101100, 101140, 101120, 101120, 101110, 101130, 101130, 101140, 
    101170, 101170, 101170, 101190, 101210, 101180, 101150, 101130, 101160, 
    101090, 101100, 101120, 101120, 101070, 101070, 101010, 100980, 100960, 
    100950, 100910, 100940, 100910, 100880, 100880, 100900, 100910, 100890, 
    100860, 100880, 100830, 100800, 100810, 100750, 100720, 100710, 100710, 
    100700, 100680, 100690, 100720, 100700, 100750, 100730, 100730, 100720, 
    100710, 100670, 100680, 100660, 100610, 100560, 100510, 100470, 100430, 
    100480, 100470, 100490, 100450, 100370, 100380, 100370, 100280, 100260, 
    100250, 100180, 100100, 100010, 99950, 99980, 99930, 99900, 99840, 99880, 
    99870, 99870, 99910, 99870, 99920, 99960, 100050, 100040, 100080, 100120, 
    100190, 100260, 100270, 100300, 100320, 100340, 100380, 100450, 100440, 
    100410, 100460, 100480, 100510, 100550, 100590, 100620, 100640, 100670, 
    100720, 100760, 100800, 100820, 100850, 100840, 100880, 100890, 100960, 
    100970, 101030, 101080, 101140, 101190, 101260, 101320, 101350, 101390, 
    101450, 101490, 101550, 101600, 101630, 101660, 101720, 101780, 101840, 
    101890, 101900, 101930, 101960, 101950, 101960, 101950, 101900, 101880, 
    101880, 101850, 101820, 101770, 101730, 101660, 101600, 101540, 101440, 
    101300, 101170, 101080, 100990, 100880, 100780, 100720, 100630, 100500, 
    100360, 100280, 100210, 100130, 100050, 99970, 99900, 99790, 99720, 
    99630, 99550, 99500, 99460, 99380, 99300, 99240, 99190, 99170, 99120, 
    99090, 99080, 99120, 99190, 99250, 99300, 99350, 99370, 99400, 99430, 
    99420, 99440, 99460, 99460, 99460, 99450, 99450, 99490, 99540, 99540, 
    99540, 99520, 99550, 99570, 99600, 99680, 99770, 99820, 99870, 99950, 
    100030, 100100, 100160, 100200, 100260, 100330, 100390, 100450, 100520, 
    100570, 100640, 100680, 100740, 100770, 100800, 100840, 100920, 100990, 
    101030, 101080, 101120, 101130, 101170, 101170, 101180, 101200, 101180, 
    101140, 101100, 101070, 101020, 101040, 101030, 101000, 100970, 100940, 
    100880, 100870, 100810, 100750, 100730, 100670, 100610, 100570, 100550, 
    100420, 100290, 100210, 100090, 100010, 99930, 99840, 99810, 99760, 
    99720, 99670, 99580, 99430, 99310, 99150, 98990, 98860, 98760, 98710, 
    98700, 98760, 98810, 98870, 98950, 99030, 99090, 99130, 99150, 99230, 
    99280, 99340, 99500, 99630, 99800, 99980, 100110, 100200, 100230, 100280, 
    100300, 100360, 100400, 100450, 100480, 100510, 100550, 100570, 100550, 
    100520, 100540, 100570, 100550, 100590, 100610, 100640, 100690, 100670, 
    100700, 100700, 100730, 100580, 100670, 100690, 100750, 100810, 100900, 
    100870, 100860, 100910, 100960, 101010, 101070, 101120, 101110, 101160, 
    101200, 101250, 101300, 101370, 101420, 101460, 101530, 101580, 101620, 
    101690, 101740, 101780, 101830, 101860, 101890, 101920, 101950, 101990, 
    102030, 102100, 102130, 102170, 102180, 102190, 102210, 102240, 102260, 
    102270, 102270, 102270, 102270, 102260, 102270, 102280, 102280, 102300, 
    102280, 102280, 102230, 102220, 102200, 102200, 102200, 102200, 102200, 
    102190, 102180, 102140, 102100, 102080, 102070, 102040, 102020, 101980, 
    101920, 101880, 101840, 101810, 101770, 101720, 101680, 101620, 101540, 
    101450, 101390, 101300, 101320, 101200, 101210, 101170, 101130, 101070, 
    101010, 100980, 100880, 100840, 100820, 100710, 100740, 100700, 100670, 
    100620, 100610, 100580, 100640, 100640, 100670, 100690, 100700, 100690, 
    100590, 100560, 100450, 100460, 100440, 100410, 100400, 100420, 100410, 
    100530, 100470, 100500, 100580, 100630, 100580, 100590, 100630, 100590, 
    100650, 100710, 100700, 100690, 100710, 100660, 100670, 100620, 100520, 
    100530, 100610, 100720, 100760, 100860, 100970, 101100, 101130, 101250, 
    101340, 101460, 101510, 101570, 101640, 101670, 101720, 101730, 101740, 
    101750, 101770, 101790, 101790, 101800, 101820, 101850, 101840, 101820, 
    101830, 101810, 101820, 101800, 101750, 101690, 101710, 101660, 101560, 
    101520, 101430, 101370, 101310, 101190, 101080, 101010, 100910, 100810, 
    100730, 100680, 100560, 100500, 100390, 100300, 100210, 100150, 100050, 
    100030, 100010, 99980, 100090, 100120, 100200, 100270, 100280, 100330, 
    100450, 100510, 100550, 100730, 100730, 100730, 100750, 100800, 100890, 
    100900, 100920, 100940, 101000, 101060, 101070, 101090, 101170, 101160, 
    101190, 101230, 101250, 101240, 101200, 101220, 101210, 101240, 101210, 
    101200, 101200, 101250, 101260, 101230, 101230, 101250, 101250, 101220, 
    101210, 101230, 101230, 101240, 101230, 101270, 101270, 101290, 101370, 
    101490, 101550, 101710, 101720, 101800, 101820, 101980, 101990, 101980, 
    101980, 102170, 102300, 102330, 102380, 102400, 102420, 102410, 102370, 
    102380, 102390, 102390, 102330, 102270, 102320, 102280, 102270, 102240, 
    102170, 102140, 102090, 102090, 102040, 101970, 101900, 101850, 101760, 
    101680, 101620, 101550, 101500, 101500, 101520, 101540, 101550, 101530, 
    101570, 101570, 101560, 101530, 101510, 101470, 101450, 101400, 101370, 
    101320, 101290, 101270, 101250, 101230, 101210, 101150, 101120, 101120, 
    101140, 101140, 101130, 101120, 101130, 101130, 101160, 101140, 101120, 
    101110, 101100, 101080, 101080, 101100, 101080, 101080, 101040, 101030, 
    101020, 101070, 101080, 101070, 101050, 101030, 101010, 100990, 100980, 
    100960, 100920, 100910, 100870, 100860, 100850, 100860, 100860, 100840, 
    100830, 100850, 100850, 100850, 100860, 100840, 100860, 100870, 100880, 
    100870, 100870, 100850, 100840, 100820, 100840, 100810, 100800, 100800, 
    100790, 100790, 100790, 100800, 100770, 100750, 100760, 100740, 100730, 
    100740, 100750, 100770, 100750, 100760, 100780, 100800, 100820, 100830, 
    100850, 100850, 100860, 100900, 100900, 100900, 100920, 100950, 100960, 
    100960, 100960, 100960, 100970, 100960, 100970, 100960, 100940, 100930, 
    100940, 100970, 100990, 101000, 101010, 101000, 101000, 100990, 100970, 
    100960, 100970, 100950, 100930, 100900, 100880, 100860, 100830, 100830, 
    100790, 100780, 100720, 100660, 100620, 100570, 100540, 100490, 100490, 
    100450, 100580, 100400, 100470, 100550, 100520, 100490, 100460, 100430, 
    100410, 100410, 100330, 100290, 100250, 100220, 100260, 100270, 100320, 
    100210, 100240, 100270, 100310, 100430, 100500, 100550, 100550, 100560, 
    100570, 100590, 100610, 100610, 100620, 100660, 100670, 100660, 100660, 
    100650, 100640, 100550, 100570, 100580, 100650, 100600, 100590, 100620, 
    100640, 100630, 100630, 100630, 100620, 100600, 100600, 100590, 100580, 
    100570, 100570, 100560, 100530, 100560, 100550, 100550, 100510, 100500, 
    100490, 100490, 100450, 100440, 100490, 100490, 100520, 100520, 100500, 
    100500, 100590, 100520, 100530, 100540, 100510, 100510, 100480, 100470, 
    100470, 100460, 100400, 100360, 100320, 100220, 100320, 100400, 100380, 
    100350, 100350, 100360, 100290, 100370, 100330, 100260, 100270, 100290, 
    100290, 100240, 100250, 100230, 100240, 100240, 100270, 100300, 100320, 
    100320, 100320, 100320, 100350, 100370, 100380, 100420, 100420, 100420, 
    100460, 100480, 100510, 100460, 100450, 100460, 100490, 100490, 100510, 
    100520, 100550, 100590, 100610, 100630, 100670, 100700, 100690, 100680, 
    100680, 100760, 100830, 100870, 100920, 100960, 101020, 101060, 101120, 
    101160, 101170, 101210, 101250, 101290, 101330, 101370, 101400, 101450, 
    101480, 101500, 101540, 101580, 101610, 101630, 101650, 101680, 101710, 
    101730, 101740, 101750, 101770, 101800, 101810, 101810, 101800, 101800, 
    101790, 101810, 101800, 101780, 101780, 101740, 101730, 101730, 101720, 
    101680, 101660, 101650, 101660, 101630, 101630, 101600, 101590, 101590, 
    101590, 101580, 101590, 101590, 101590, 101590, 101550, 101520, 101550, 
    101520, 101510, 101490, 101490, 101490, 101490, 101480, 101480, 101450, 
    101440, 101430, 101440, 101440, 101420, 101410, 101430, 101460, 101450, 
    101430, 101420, 101390, 101390, 101400, 101390, 101400, 101410, 101370, 
    101390, 101370, 101350, 101350, 101300, 101270, 101290, 101290, 101250, 
    101230, 101220, 101200, 101210, 101180, 101180, 101180, 101170, 101160, 
    101160, 101160, 101130, 101110, 101070, 101070, 101070, 101080, 101110, 
    101120, 101110, 101140, 101120, 101140, 101180, 101170, 101180, 101220, 
    101240, 101260, 101280, 101280, 101240, 101190, 101080, 101030, 100920, 
    100870, 100840, 100750, 100670, 100760, 100800, 100860, 100890, 100910, 
    100990, 101080, 101140, 101230, 101340, 101400, 101520, 101550, 101570, 
    101640, 101650, 101650, 101650, 101680, 101680, 101670, 101630, 101650, 
    101650, 101650, 101650, 101730, 101780, 101860, 101980, 102000, 102040, 
    102100, 102150, 102180, 102210, 102240, 102250, 102280, 102300, 102320, 
    102340, 102370, 102380, 102410, 102420, 102430, 102410, 102410, 102370, 
    102340, 102330, 102280, 102270, 102190, 102150, 102100, 102050, 102030, 
    102070, 102070, 102040, 102050, 102050, 102060, 102040, 102030, 102010, 
    102000, 101980, 101970, 101960, 101950, 101910, 101920, 101890, 101870, 
    101820, 101750, 101720, 101600, 101520, 101440, 101410, 101350, 101310, 
    101240, 101200, 101090, 101030, 100940, 100850, 100760, 100660, 100580, 
    100500, 100470, 100440, 100450, 100410, 100380, 100350, 100350, 100350, 
    100440, 100510, 100580, 100630, 100690, 100730, 100760, 100820, 100850, 
    100900, 100880, 100890, 100960, 101050, 101150, 101220, 101300, 101370, 
    101480, 101550, 101620, 101690, 101760, 101850, 101870, 101930, 101950, 
    101990, 102050, 102070, 102090, 102120, 102140, 102130, 102120, 102120, 
    102100, 102100, 102090, 102080, 102110, 102100, 102050, 102020, 102010, 
    101950, 101950, 101900, 101860, 101860, 101850, 101810, 101780, 101770, 
    101730, 101690, 101640, 101590, 101570, 101520, 101480, 101490, 101520, 
    101580, 101600, 101600, 101740, 101860, 101930, 102010, 102050, 102060, 
    102120, 102210, 102260, 102310, 102320, 102330, 102450, 102520, 102610, 
    102650, 102650, 102740, 102740, 102750, 102750, 102730, 102710, 102660, 
    102600, 102550, 102500, 102360, 102310, 102250, 102180, 102120, 102050, 
    101990, 101980, 101960, 102020, 102060, 102090, 102160, 102240, 102290, 
    102320, 102310, 102330, 102330, 102330, 102300, 102250, 102210, 102170, 
    102120, 102070, 102020, 101960, 101900, 101860, 101790, 101730, 101670, 
    101600, 101550, 101510, 101470, 101450, 101450, 101480, 101530, 101560, 
    101590, 101660, 101620, 101740, 101780, 101790, 101840, 101870, 101900, 
    101910, 101960, 101990, 102010, 102060, 102060, 102130, 102180, 102190, 
    102250, 102260, 102270, 102330, 102410, 102400, 102430, 102520, 102510, 
    102520, 102510, 102510, 102500, 102560, 102560, 102480, 102410, 102430, 
    102460, 102460, 102410, 102390, 102350, 102300, 102270, 102220, 102200, 
    102130, 102100, 102070, 102020, 101990, 101950, 101880, 101800, 101740, 
    101680, 101620, 101530, 101460, 101420, 101400, 101390, 101390, 101340, 
    101380, 101390, 101440, 101430, 101420, 101380, 101380, 101360, 101350, 
    101340, 101330, 101340, 101340, 101360, 101310, 101280, 101230, 101200, 
    101170, 101140, 101180, 101150, 101180, 101280, 101310, 101310, 101370, 
    101440, 101490, 101520, 101530, 101610, 101710, 101750, 101790, 101820, 
    101820, 101820, 101790, 101790, 101780, 101750, 101700, 101680, 101630, 
    101570, 101530, 101510, 101460, 101420, 101370, 101320, 101270, 101250, 
    101220, 101180, 101150, 101160, 101160, 101160, 101190, 101240, 101270, 
    101310, 101360, 101390, 101430, 101470, 101520, 101620, 101700, 101770, 
    101830, 101910, 102000, 102050, 102120, 102180, 102210, 102240, 102290, 
    102330, 102380, 102420, 102460, 102490, 102480, 102500, 102500, 102510, 
    102490, 102480, 102460, 102490, 102500, 102540, 102530, 102540, 102550, 
    102550, 102540, 102520, 102510, 102500, 102480, 102490, 102510, 102520, 
    102500, 102500, 102480, 102460, 102440, 102420, 102380, 102350, 102310, 
    102300, 102300, 102290, 102250, 102280, 102250, 102250, 102230, 102250, 
    102230, 102220, 102230, 102230, 102220, 102200, 102200, 102190, 102120, 
    102150, 102160, 102150, 102140, 102130, 102160, 102150, 102170, 102170, 
    102160, 102150, 102140, 102130, 102120, 102110, 102060, 102040, 102050, 
    102040, 102020, 102000, 101970, 101960, 101930, 101900, 101890, 101860, 
    101830, 101840, 101840, 101840, 101860, 101840, 101830, 101850, 101840, 
    101810, 101790, 101780, 101760, 101750, 101750, 101700, 101700, 101670, 
    101650, 101640, 101620, 101630, 101620, 101600, 101570, 101560, 101600, 
    101660, 101750, 101820, 101880, 101910, 101950, 101910, 101940, 101900, 
    101960, 101920, 101820, 101800, 101800, 101830, 101810, 101790, 101710, 
    101690, 101680, 101640, 101610, 101860, 101550, 101630, 101660, 101740, 
    101670, 101710, 101700, 101670, 101670, 101710, 101630, 101640, 101760, 
    101750, 101680, 101670, 101710, 101790, 101840, 101890, 101970, 102040, 
    102140, 102160, 102180, 102250, 102370, 102480, 102530, 102590, 102690, 
    102750, 102820, 102850, 102880, 102900, 102900, 102950, 102990, 102940, 
    102890, 102840, 102860, 102840, 102780, 102770, 102790, 102790, 102820, 
    102800, 102760, 102790, 102750, 102660, 102640, 102620, 102610, 102550, 
    102560, 102530, 102530, 102580, 102560, 102530, 102530, 102530, 102510, 
    102520, 102510, 102550, 102560, 102570, 102590, 102630, 102650, 102700, 
    102700, 102730, 102750, 102740, 102740, 102740, 102750, 102780, 102790, 
    102820, 102820, 102820, 102830, 102820, 102780, 102720, 102710, 102610, 
    102600, 102580, 102500, 102430, 102340, 102270, 102220, 102120, 102160, 
    102070, 102160, 102110, 102050, 102000, 102020, 102000, 101980, 102000, 
    101930, 101940, 101940, 101960, 102020, 102050, 102040, 102040, 101990, 
    102080, 102160, 102200, 102210, 102200, 102190, 102250, 102210, 102180, 
    102170, 102170, 102160, 102160, 102130, 102080, 102140, 102160, 102130, 
    102220, 102190, 102260, 102320, 102370, 102400, 102450, 102520, 102570, 
    102580, 102610, 102620, 102640, 102660, 102660, 102620, 102680, 102690, 
    102700, 102710, 102720, 102730, 102680, 102680, 102650, 102630, 102580, 
    102600, 102630, 102570, 102470, 102470, 102600, 102500, 102580, 102580, 
    102540, 102540, 102460, 102350, 102360, 102350, 102320, 102380, 102330, 
    102360, 102340, 102300, 102270, 102270, 102290, 102330, 102290, 102290, 
    102280, 102320, 102290, 102280, 102240, 102200, 102190, 102140, 102100, 
    102030, 101980, 101900, 101830, 101760, 101720, 101690, 101640, 101600, 
    101520, 101550, 101540, 101480, 101440, 101440, 101420, 101390, 101330, 
    101320, 101270, 101230, 101190, 101160, 101160, 101130, 101120, 101060, 
    101060, 101040, 100980, 100960, 100920, 100880, 100820, 100750, 100690, 
    100670, 100610, 100570, 100560, 100560, 100530, 100480, 100460, 100450, 
    100450, 100450, 100450, 100470, 100510, 100530, 100570, 100610, 100660, 
    100710, 100770, 100830, 100890, 100940, 101000, 101060, 101110, 101170, 
    101240, 101300, 101350, 101390, 101440, 101470, 101520, 101530, 101530, 
    101510, 101580, 101590, 101620, 101670, 101680, 101750, 101730, 101750, 
    101800, 101850, 101900, 101830, 101830, 101860, 102190, 101930, 101950, 
    101960, 101970, 101990, 102100, 102200, 102280, 102370, 102470, 102530, 
    102650, 102710, 102760, 102820, 102870, 102920, 103010, 103070, 103150, 
    103230, 103290, 103310, 103380, 103470, 103530, 103580, 103600, 103630, 
    103640, 103720, 103800, 103860, 103970, 104070, 104140, 104200, 104230, 
    104310, 104390, 104460, 104530, 104590, 104610, 104660, 104690, 104710, 
    104730, 104830, 104870, 104890, 104880, 104940, 104940, 104960, 105010, 
    105060, 105070, 105130, 105100, 105120, 105120, 105130, 105240, 105010, 
    105030, 105060, 104940, 104980, 105080, 105120, 105180, 105260, 105290, 
    105310, 105310, 105360, 105380, 105380, 105390, 105390, 105410, 105460, 
    105510, 105570, 105640, 105680, 105720, 105760, 105770, 105800, 105860, 
    105870, 105890, 105900, 105900, 105920, 105950, 105980, 105980, 105980, 
    105980, 105980, 105980, 105950, 105900, 105880, 105850, 105810, 105760, 
    105690, 105620, 105580, 105500, 105430, 105350, 105280, 105170, 105110, 
    105050, 105000, 104960, 104940, 104870, 104780, 104660, 104690, 104540, 
    104450, 104310, 104260, 104200, 104150, 104190, 104120, 104110, 104040, 
    103960, 103830, 103770, 103730, 103670, 103570, 103450, 103410, 103380, 
    103350, 103320, 103300, 103300, 103280, 103270, 103260, 103250, 103240, 
    103230, 103260, 103260, 103280, 103250, 103250, 103200, 103210, 103220, 
    103200, 103170, 103150, 103200, 103210, 103170, 103180, 103180, 103200, 
    103200, 103170, 103140, 103120, 103080, 103040, 103010, 102990, 102980, 
    102970, 102960, 102950, 102950, 102920, 102920, 102910, 102920, 102920, 
    102930, 102990, 103010, 103050, 103050, 103050, 103070, 103080, 103100, 
    103110, 103110, 103110, 103120, 103130, 103130, 103110, 103090, 103090, 
    103070, 103050, 103010, 103000, 102900, 102860, 102900, 102830, 102760, 
    102720, 102610, 102550, 102540, 102550, 102600, 102590, 102590, 102530, 
    102550, 102570, 102570, 102580, 102570, 102570, 102430, 102390, 102430, 
    102490, 102520, 102520, 102520, 102590, 102580, 102600, 102590, 102510, 
    102420, 102200, 102150, 102080, 102140, 102100, 102070, 102140, 102180, 
    102160, 102140, 102180, 102170, 102270, 102270, 102170, 102140, 102160, 
    102210, 102280, 102240, 102310, 102290, 102340, 102370, 102360, 102350, 
    102330, 102300, 102220, 102160, 102180, 102220, 102240, 102220, 102230, 
    102180, 102240, 102270, 102290, 102260, 102300, 102330, 102340, 102360, 
    102360, 102350, 102340, 102310, 102290, 102270, 102270, 102260, 102260, 
    102230, 102220, 102210, 102170, 102150, 102150, 102120, 102080, 102050, 
    102050, 102050, 102020, 102010, 101990, 101970, 101960, 101910, 101850, 
    101800, 101780, 101740, 101680, 101610, 101560, 101510, 101470, 101450, 
    101440, 101420, 101400, 101380, 101350, 101330, 101300, 101280, 101240, 
    101200, 101140, 101130, 101100, 101030, 100950, 100920, 100860, 100820, 
    100730, 100630, 100620, 100610, 100600, 100540, 100500, 100470, 100420, 
    100410, 100350, 100310, 100290, 100250, 100210, 100170, 100180, 100170, 
    100120, 100050, 100070, 100070, 100080, 100100, 100130, 100120, 100130, 
    100070, 100100, 100140, 100160, 100170, 100150, 100120, 100160, 100190, 
    100210, 100220, 100200, 100160, 100160, 100190, 100200, 100180, 100200, 
    100170, 100280, 100320, 100410, 100500, 100590, 100680, 100810, 100900, 
    100970, 101050, 101130, 101220, 101270, 101300, 101340, 101390, 101430, 
    101440, 101460, 101560, 101610, 101610, 101650, 101610, 101590, 101800, 
    101810, 101850, 101790, 101830, 101820, 101900, 101900, 101880, 101900, 
    101900, 101860, 101870, 101840, 101800, 101800, 101790, 101640, 101760, 
    101720, 101700, 101680, 101750, 101810, 101760, 101760, 101780, 101850, 
    101950, 101980, 102030, 102090, 102050, 101980, 102010, 102050, 102030, 
    102100, 102110, 102120, 102200, 102220, 102240, 102230, 102290, 102290, 
    102330, 102370, 102420, 102430, 102450, 102430, 102320, 102430, 102480, 
    102530, 102500, 102460, 102380, 102310, 102280, 102310, 102390, 102390, 
    102400, 102400, 102330, 102380, 102420, 102480, 102530, 102560, 102540, 
    102550, 102560, 102530, 102540, 102560, 102490, 102490, 102470, 102410, 
    102400, 102400, 102360, 102320, 102220, 102210, 102170, 102110, 102070, 
    102000, 102000, 101970, 101910, 101830, 101790, 101720, 101730, 101750, 
    101760, 101680, 101680, 101620, 101590, 101600, 101650, 101630, 101610, 
    101570, 101560, 101550, 101480, 101500, 101440, 101560, 101520, 101500, 
    101500, 101480, 101430, 101450, 101430, 101350, 101320, 101290, 101260, 
    101210, 101160, 101120, 101090, 101020, 101030, 101000, 100990, 100960, 
    100980, 100960, 100980, 100950, 100920, 100900, 100910, 100890, 100870, 
    100840, 100830, 100830, 100820, 100820, 100780, 100780, 100770, 100770, 
    100770, 100720, 100720, 100720, 100690, 100710, 100740, 100740, 100700, 
    100700, 100680, 100650, 100630, 100630, 100610, 100600, 100590, 100600, 
    100610, 100550, 100560, 100540, 100520, 100510, 100460, 100490, 100490, 
    100460, 100460, 100440, 100440, 100470, 100470, 100450, 100520, 100540, 
    100530, 100590, 100570, 100570, 100610, 100630, 100700, 100760, 100740, 
    100790, 100870, 100900, 100910, 100930, 100970, 101020, 101050, 101100, 
    101070, 100940, 101270, 101320, 101330, 101320, 101360, 101410, 101400, 
    101450, 101450, 101490, 101550, 101580, 101590, 101610, 101640, 101660, 
    101640, 101650, 101630, 101630, 101650, 101660, 101670, 101670, 101660, 
    101630, 101630, 101620, 101610, 101580, 101560, 101570, 101560, 101560, 
    101540, 101550, 101550, 101540, 101520, 101500, 101500, 101490, 101490, 
    101470, 101460, 101460, 101490, 101490, 101500, 101510, 101500, 101490, 
    101490, 101470, 101460, 101470, 101470, 101460, 101450, 101410, 101400, 
    101360, 101330, 101290, 101250, 101240, 101210, 101170, 101140, 101080, 
    101050, 101000, 100980, 100940, 100910, 100860, 100850, 100840, 100820, 
    100820, 100780, 100790, 100800, 100800, 100790, 100790, 100770, 100770, 
    100760, 100770, 100800, 100800, 100800, 100830, 100840, 100840, 100860, 
    100840, 100830, 100830, 100810, 100800, 100830, 100890, 100920, 100980, 
    101020, 101060, 101090, 101120, 101160, 101190, 101220, 101230, 101250, 
    101260, 101310, 101340, 101360, 101380, 101400, 101410, 101410, 101400, 
    101400, 101370, 101370, 101370, 101360, 101360, 101330, 101280, 101240, 
    101240, 101210, 101160, 101100, 101070, 101040, 100980, 100940, 100910, 
    100870, 100820, 100750, 100770, 100750, 100730, 100640, 100610, 100620, 
    100570, 100570, 100550, 100520, 100490, 100480, 100480, 100440, 100430, 
    100390, 100390, 100440, 100460, 100460, 100450, 100440, 100430, 100410, 
    100440, 100470, 100440, 100470, 100490, 100480, 100480, 100500, 100500, 
    100520, 100530, 100540, 100540, 100560, 100570, 100570, 100560, 100570, 
    100610, 100610, 100630, 100640, 100670, 100690, 100710, 100710, 100730, 
    100780, 100810, 100840, 100870, 100970, 101000, 100960, 100990, 101000, 
    101020, 101030, 101080, 101110, 101130, 101190, 101220, 101240, 101280, 
    101330, 101350, 101400, 101460, 101460, 101500, 101540, 101590, 101570, 
    101610, 101650, 101670, 101680, 101680, 101730, 101730, 101780, 101810, 
    101870, 101860, 101920, 101950, 101980, 102020, 102060, 102090, 102090, 
    102080, 102040, 102020, 102000, 101970, 101930, 101890, 101850, 101800, 
    101730, 101670, 101650, 101570, 101480, 101410, 101290, 101210, 101040, 
    100950, 100900, 100840, 100800, 100730, 100680, 100650, 100570, 100540, 
    100500, 100500, 100470, 100470, 100410, 100320, 100280, 100260, 100170, 
    100070, 100020, 99970, 99930, 99880, 99820, 99780, 99730, 99710, 99670, 
    99630, 99580, 99580, 99520, 99530, 99560, 99580, 99610, 99660, 99730, 
    99790, 99810, 99840, 99850, 99860, 99820, 99830, 99820, 99770, 99750, 
    99740, 99720, 99720, 99690, 99670, 99620, 99570, 99530, 99540, 99500, 
    99520, 99550, 99580, 99620, 99660, 99690, 99720, 99770, 99810, 99840, 
    99840, 99860, 99860, 99900, 99920, 99930, 99930, 99960, 99940, 99960, 
    99980, 100020, 100060, 100070, 100090, 100110, 100130, 100170, 100220, 
    100240, 100270, 100330, 100360, 100430, 100450, 100470, 100490, 100520, 
    100540, 100540, 100550, 100580, 100570, 100570, 100570, 100570, 100570, 
    100550, 100520, 100500, 100470, 100470, 100470, 100460, 100450, 100460, 
    100460, 100470, 100510, 100560, 100580, 100580, 100630, 100670, 100710, 
    100750, 100780, 100840, 100900, 100930, 100980, 101050, 101050, 101060, 
    101130, 101160, 101200, 101230, 101290, 101320, 101370, 101400, 101430, 
    101450, 101440, 101450, 101460, 101400, 101420, 101410, 101410, 101370, 
    101250, 101250, 101260, 101220, 101080, 100970, 100850, 100800, 100850, 
    100860, 100830, 100780, 100750, 100720, 100690, 100670, 100660, 100600, 
    100590, 100560, 100550, 100580, 100610, 100660, 100710, 100780, 100820, 
    100850, 100880, 100890, 100900, 100930, 100940, 100950, 100980, 101070, 
    101110, 101110, 101130, 101150, 101170, 101200, 101230, 101240, 101270, 
    101300, 101330, 101360, 101390, 101410, 101420, 101430, 101420, 101430, 
    101440, 101470, 101490, 101510, 101540, 101550, 101560, 101570, 101590, 
    101570, 101600, 101560, 101570, 101560, 101570, 101570, 101570, 101560, 
    101520, 101500, 101460, 101420, 101370, 101320, 101240, 101220, 101160, 
    101140, 101100, 101070, 101060, 100990, 100950, 100950, 100910, 100890, 
    100870, 100870, 100900, 100890, 100880, 100880, 100870, 100850, 100830, 
    100800, 100760, 100710, 100670, 100620, 100590, 100540, 100480, 100440, 
    100390, 100350, 100310, 100270, 100230, 100200, 100190, 100190, 100180, 
    100210, 100230, 100250, 100270, 100280, 100290, 100310, 100330, 100340, 
    100350, 100360, 100390, 100420, 100450, 100460, 100480, 100520, 100530, 
    100550, 100550, 100590, 100630, 100660, 100690, 100750, 100830, 100870, 
    100930, 100990, 101010, 101020, 101040, 101070, 101100, 101160, 101180, 
    101210, 101240, 101280, 101290, 101320, 101340, 101340, 101350, 101370, 
    101350, 101360, 101390, 101440, 101440, 101500, 101530, 101530, 101530, 
    101540, 101530, 101570, 101610, 101600, 101600, 101600, 101620, 101650, 
    101680, 101670, 101650, 101620, 101620, 101620, 101590, 101590, 101590, 
    101580, 101570, 101590, 101600, 101590, 101580, 101570, 101540, 101510, 
    101490, 101470, 101460, 101440, 101430, 101410, 101390, 101360, 101350, 
    101330, 101310, 101290, 101260, 101240, 101210, 101190, 101180, 101150, 
    101150, 101120, 101100, 101070, 101040, 101000, 101000, 100980, 100970, 
    100950, 100950, 100970, 100990, 101020, 101030, 101050, 101070, 101080, 
    101100, 101130, 101170, 101200, 101240, 101280, 101300, 101330, 101350, 
    101380, 101390, 101400, 101410, 101420, 101440, 101450, 101470, 101500, 
    101510, 101530, 101510, 101540, 101550, 101570, 101590, 101590, 101610, 
    101620, 101650, 101670, 101690, 101700, 101680, 101670, 101670, 101670, 
    101650, 101630, 101630, 101630, 101610, 101600, 101570, 101570, 101550, 
    101530, 101500, 101470, 101440, 101400, 101380, 101310, 101290, 101280, 
    101260, 101230, 101160, 101140, 101090, 101050, 101020, 101010, 100970, 
    100930, 100920, 100920, 100960, 100960, 100960, 100990, 100980, 101000, 
    101040, 101050, 101100, 101150, 101180, 101220, 101280, 101330, 101370, 
    101390, 101430, 101470, 101490, 101570, 101640, 101680, 101740, 101780, 
    101810, 101850, 101870, 101920, 101950, 101990, 102020, 102050, 102080, 
    102120, 102140, 102190, 102230, 102230, 102260, 102280, 102290, 102320, 
    102360, 102390, 102410, 102470, 102510, 102540, 102560, 102590, 102640, 
    102700, 102740, 102760, 102810, 102830, 102870, 102890, 102930, 102960, 
    102960, 102970, 102970, 102970, 102950, 102950, 102960, 102930, 102950, 
    102940, 102950, 102920, 102910, 102900, 102890, 102900, 102880, 102860, 
    102860, 102850, 102840, 102840, 102840, 102830, 102800, 102800, 102810, 
    102810, 102780, 102780, 102780, 102780, 102750, 102740, 102730, 102730, 
    102720, 102720, 102690, 102690, 102690, 102680, 102690, 102670, 102690, 
    102690, 102700, 102710, 102720, 102720, 102720, 102730, 102750, 102770, 
    102770, 102780, 102800, 102830, 102840, 102850, 102880, 102900, 102930, 
    102950, 102990, 103020, 103040, 103070, 103110, 103130, 103160, 103200, 
    103250, 103250, 103260, 103300, 103320, 103330, 103350, 103370, 103370, 
    103390, 103390, 103390, 103400, 103400, 103390, 103380, 103370, 103360, 
    103310, 103240, 103190, 103130, 103090, 103070, 103020, 102970, 102890, 
    102880, 102820, 102760, 102650, 102560, 102500, 102430, 102360, 102250, 
    102140, 102030, 101920, 101850, 101770, 101650, 101540, 101450, 101390, 
    101360, 101250, 101140, 101140, 101090, 101070, 101060, 101160, 101120, 
    101150, 101170, 101200, 101220, 101270, 101330, 101380, 101450, 101480, 
    101520, 101560, 101630, 101680, 101710, 101770, 101830, 101890, 101930, 
    101970, 102050, 102080, 102080, 102120, 102160, 102180, 102210, 102250, 
    102280, 102300, 102340, 102320, 102320, 102370, 102370, 102340, 102330, 
    102320, 102310, 102310, 102290, 102280, 102250, 102250, 102250, 102260, 
    102220, 102200, 102200, 102200, 102190, 102150, 102160, 102140, 102130, 
    102090, 102090, 102060, 102030, 102010, 101980, 101970, 101970, 101980, 
    102000, 102060, 102120, 102160, 102180, 102190, 102220, 102260, 102300, 
    102320, 102350, 102360, 102400, 102430, 102450, 102480, 102480, 102490, 
    102500, 102500, 102500, 102510, 102530, 102530, 102550, 102580, 102610, 
    102630, 102650, 102670, 102680, 102680, 102660, 102650, 102640, 102660, 
    102670, 102690, 102680, 102700, 102670, 102650, 102640, 102620, 102580, 
    102560, 102520, 102480, 102420, 102350, 102280, 102200, 102150, 102020, 
    101950, 101840, 101740, 101660, 101540, 101460, 101400, 101320, 101240, 
    101200, 101130, 101060, 101020, 100950, 100900, 100820, 100710, 100660, 
    100580, 100510, 100420, 100320, 100260, 100150, 100040, 99960, 99880, 
    99880, 99830, 99840, 99810, 99880, 99920, 99960, 100050, 100110, 100240, 
    100380, 100520, 100610, 100710, 100850, 100960, 101040, 101150, 101210, 
    101290, 101350, 101390, 101430, 101460, 101500, 101490, 101510, 101510, 
    101530, 101560, 101570, 101550, 101530, 101530, 101550, 101550, 101550, 
    101580, 101590, 101670, 101730, 101760, 101760, 101780, 101790, 101790, 
    101790, 101800, 101790, 101800, 101820, 101760, 101840, 101860, 101860, 
    101880, 101880, 101870, 101860, 101870, 101890, 101910, 101930, 101950, 
    101960, 101970, 101960, 101970, 101970, 101950, 101930, 101900, 101910, 
    101890, 101900, 101910, 101920, 101920, 101940, 101960, 101990, 102000, 
    102020, 102040, 102070, 102110, 102160, 102200, 102260, 102280, 102300, 
    102320, 102340, 102350, 102340, 102370, 102380, 102370, 102400, 102400, 
    102420, 102400, 102370, 102310, 102270, 102200, 102070, 101960, 101810, 
    101790, 101650, 101650, 101660, 101680, 101740, 101870, 101940, 101960, 
    102010, 102100, 102140, 102210, 102220, 102260, 102290, 102260, 102270, 
    102220, 102190, 102170, 102140, 102070, 102020, 102000, 102000, 101970, 
    101890, 101860, 101830, 101770, 101720, 101650, 101620, 101550, 101530, 
    101510, 101530, 101530, 101560, 101550, 101540, 101560, 101540, 101570, 
    101540, 101560, 101600, 101630, 101650, 101680, 101740, 101780, 101810, 
    101840, 101880, 101880, 101930, 101950, 101990, 101990, 102050, 102100, 
    102140, 102170, 102200, 102210, 102240, 102260, 102300, 102300, 102360, 
    102410, 102460, 102500, 102530, 102610, 102630, 102660, 102710, 102720, 
    102740, 102760, 102790, 102780, 102790, 102830, 102830, 102820, 102830, 
    102830, 102830, 102790, 102800, 102780, 102770, 102740, 102750, 102780, 
    102790, 102770, 102740, 102730, 102690, 102670, 102630, 102600, 102580, 
    102550, 102550, 102550, 102530, 102480, 102440, 102390, 102330, 102260, 
    102240, 102190, 102080, 101990, 101970, 101990, 101930, 101880, 101800, 
    101790, 101730, 101720, 101700, 101640, 101640, 101610, 101580, 101540, 
    101540, 101490, 101380, 101320, 101260, 101170, 101110, 101080, 101140, 
    101140, 101170, 101270, 101330, 101420, 101460, 101470, 101490, 101450, 
    101460, 101430, 101490, 101530, 101590, 101600, 101650, 101710, 101770, 
    101700, 101720, 101640, 101540, 101530, 101450, 101340, 101250, 101160, 
    101040, 101020, 100990, 100960, 100920, 100870, 100830, 100800, 100770, 
    100750, 100700, 100690, 100770, 100760, 100790, 100830, 100860, 100880, 
    100910, 100940, 100960, 100980, 100990, 101030, 101070, 101090, 101110, 
    101130, 101140, 101210, 101170, 101120, 101080, 101100, 101080, 101080, 
    101010, 100980, 100880, 100800, 100690, 100560, 100450, 100330, 100220, 
    100200, 100230, 100240, 100300, 100380, 100480, 100640, 100770, 100890, 
    100980, 101060, 101100, 101160, 101170, 101180, 101240, 101270, 101230, 
    101190, 101180, 101130, 101030, 101050, 101100, 101110, 101180, 101200, 
    101280, 101330, 101350, 101390, 101420, 101410, 101380, 101360, 101310, 
    101260, 101230, 101200, 101140, 101040, 100960, 100910, 100830, 100770, 
    100710, 100660, 100600, 100560, 100520, 100460, 100470, 100490, 100480, 
    100450, 100430, 100440, 100470, 100530, 100590, 100640, 100680, 100740, 
    100720, 100710, 100690, 100670, 100660, 100670, 100620, 100590, 100570, 
    100560, 100540, 100540, 100540, 100500, 100480, 100460, 100430, 100430, 
    100430, 100460, 100470, 100450, 100490, 100550, 100610, 100580, 100550, 
    100570, 100600, 100760, 100770, 100790, 100770, 100750, 100790, 100860, 
    100880, 100910, 100920, 100950, 100950, 100900, 100900, 100850, 100840, 
    100800, 100780, 100750, 100710, 100690, 100660, 100620, 100580, 100540, 
    100520, 100490, 100460, 100450, 100410, 100440, 100410, 100430, 100400, 
    100400, 100420, 100460, 100470, 100490, 100460, 100480, 100490, 100490, 
    100440, 100390, 100360, 100360, 100360, 100330, 100300, 100300, 100310, 
    100270, 100230, 100220, 100200, 100140, 100090, 100050, 100010, 100000, 
    99970, 99930, 99850, 99800, 99740, 99710, 99710, 99700, 99660, 99580, 
    99530, 99500, 99480, 99480, 99490, 99470, 99490, 99480, 99460, 99410, 
    99430, 99470, 99490, 99460, 99430, 99430, 99440, 99440, 99440, 99470, 
    99440, 99500, 99520, 99570, 99600, 99640, 99710, 99730, 99760, 99780, 
    99810, 99840, 99860, 99890, 99950, 99960, 99990, 100020, 100050, 100060, 
    100040, 100050, 100070, 100100, 100130, 100130, 100130, 100130, 100130, 
    100140, 100130, 100160, 100170, 100190, 100200, 100210, 100210, 100210, 
    100210, 100240, 100260, 100270, 100270, 100280, 100280, 100290, 100290, 
    100300, 100290, 100260, 100230, 100220, 100170, 100150, 100120, 100100, 
    100090, 100080, 100090, 100100, 100110, 100130, 100140, 100140, 100130, 
    100140, 100130, 100120, 100140, 100140, 100150, 100190, 100240, 100250, 
    100300, 100320, 100350, 100400, 100440, 100460, 100490, 100530, 100570, 
    100610, 100670, 100700, 100740, 100750, 100790, 100810, 100810, 100820, 
    100830, 100830, 100800, 100790, 100780, 100800, 100790, 100790, 100770, 
    100800, 100810, 100780, 100820, 100850, 100850, 100900, 100940, 100990, 
    101010, 101050, 101060, 101080, 101110, 101140, 101140, 101130, 101130, 
    101100, 101100, 101100, 101050, 101020, 101000, 100980, 100980, 100960, 
    100910, 100920, 100940, 100960, 100960, 100980, 100980, 100980, 101010, 
    101000, 101030, 101020, 101010, 101050, 101060, 101050, 101060, 101080, 
    101090, 101100, 101100, 101110, 101130, 101140, 101150, 101160, 101160, 
    101170, 101180, 101180, 101190, 101190, 101160, 101160, 101150, 101170, 
    101210, 101220, 101210, 101230, 101240, 101240, 101240, 101240, 101240, 
    101240, 101240, 101240, 101240, 101250, 101220, 101270, 101270, 101270, 
    101270, 101270, 101250, 101220, 101170, 101120, 101080, 101010, 100940, 
    100890, 100820, 100650, 100490, 100330, 100250, 100190, 100140, 100060, 
    100020, 99970, 99920, 99920, 99910, 99840, 99800, 99770, 99730, 99710, 
    99680, 99680, 99650, 99640, 99620, 99630, 99650, 99640, 99650, 99660, 
    99660, 99670, 99680, 99650, 99640, 99610, 99650, 99700, 99820, 99960, 
    100090, 100220, 100350, 100450, 100620, 100800, 100930, 100910, 100990, 
    101060, 101250, 101310, 101370, 101400, 101460, 101510, 101550, 101560, 
    101600, 101650, 101650, 101680, 101680, 101670, 101680, 101660, 101630, 
    101550, 101500, 101470, 101410, 101350, 101350, 101320, 101290, 101260, 
    101220, 101210, 101200, 101190, 101170, 101140, 101140, 101110, 101120, 
    101110, 101120, 101110, 101120, 101130, 101130, 101110, 101100, 101080, 
    101080, 101060, 101080, 101060, 101060, 101040, 101030, 101020, 101030, 
    101020, 101000, 101020, 101020, 101020, 101030, 101020, 101050, 101060, 
    101080, 101080, 101090, 101100, 101110, 101100, 101120, 101140, 101200, 
    101200, 101180, 101170, 101180, 101190, 101250, 101280, 101230, 101160, 
    101150, 101160, 101230, 101300, 101340, 101360, 101400, 101450, 101530, 
    101550, 101590, 101600, 101640, 101680, 101690, 101740, 101780, 101740, 
    101730, 101720, 101680, 101670, 101640, 101560, 101520, 101450, 101370, 
    101300, 101220, 101240, 101170, 101130, 101070, 101050, 101030, 100970, 
    100970, 101030, 101090, 101080, 101170, 101160, 101140, 101140, 101220, 
    101200, 101180, 101200, 101210, 101230, 101180, 101190, 101180, 101090, 
    101090, 101000, 100880, 100820, 100720, 100620, 100610, 100590, 100530, 
    100490, 100530, 100580, 100560, 100560, 100590, 100630, 100650, 100690, 
    100700, 100720, 100800, 100830, 100910, 100960, 100950, 100950, 100930, 
    100940, 100960, 100910, 100900, 100860, 100870, 100860, 100840, 100800, 
    100790, 100770, 100760, 100770, 100820, 100880, 100930, 100970, 101040, 
    101130, 101200, 101260, 101270, 101300, 101320, 101360, 101370, 101400, 
    101430, 101440, 101490, 101530, 101530, 101560, 101560, 101560, 101560, 
    101570, 101570, 101570, 101570, 101490, 101530, 101570, 101520, 101520, 
    101500, 101530, 101460, 101440, 101420, 101390, 101340, 101350, 101330, 
    101290, 101270, 101260, 101220, 101150, 101080, 101050, 101000, 100990, 
    100920, 100920, 100890, 100830, 100530, 100440, 100500, 100440, 100460, 
    100460, 100360, 100310, 100280, 100310, 100290, 100270, 100300, 100350, 
    100350, 100380, 100400, 100420, 100460, 100450, 100420, 100450, 100500, 
    100530, 100570, 100610, 100640, 100660, 100680, 100710, 100760, 100760, 
    100780, 100810, 100850, 100880, 100900, 100970, 100970, 100960, 100990, 
    101020, 101030, 101020, 101020, 100990, 101000, 101020, 101040, 101040, 
    101070, 101060, 101050, 101030, 100960, 100990, 101010, 101000, 100970, 
    100970, 100940, 100940, 100950, 100980, 100980, 100990, 100960, 100930, 
    100910, 100910, 100930, 100930, 100940, 100930, 100860, 100780, 100730, 
    100650, 100630, 100590, 100550, 100540, 100520, 100520, 100520, 100500, 
    100520, 100550, 100550, 100550, 100520, 100500, 100490, 100470, 100450, 
    100440, 100440, 100390, 100330, 100290, 100220, 100150, 100140, 100080, 
    100010, 99940, 99910, 99890, 99860, 99820, 99800, 99780, 99740, 99740, 
    99740, 99700, 99660, 99650, 99650, 99670, 99660, 99650, 99660, 99640, 
    99630, 99610, 99600, 99600, 99610, 99600, 99590, 99590, 99570, 99560, 
    99550, 99530, 99550, 99600, 99650, 99660, 99700, 99730, 99770, 99790, 
    99790, 99810, 99860, 99900, 99890, 99910, 99890, 99860, 99850, 99900, 
    99950, 99980, 100010, 100030, 100050, 100030, 100020, 100030, 100040, 
    100030, 100040, 100020, 100040, 100100, 100110, 100120, 100170, 100220, 
    100270, 100360, 100410, 100460, 100510, 100600, 100650, 100700, 100770, 
    100810, 100890, 100970, 101020, 101070, 101100, 101140, 101190, 101250, 
    101280, 101340, 101390, 101440, 101470, 101500, 101530, 101540, 101550, 
    101570, 101580, 101580, 101560, 101540, 101520, 101520, 101550, 101540, 
    101520, 101460, 101470, 101440, 101420, 101410, 101390, 101370, 101340, 
    101340, 101310, 101300, 101290, 101240, 101220, 101170, 101170, 101110, 
    101090, 101100, 101080, 101090, 101120, 101070, 101040, 101000, 100990, 
    100940, 100870, 100740, 100660, 100640, 100550, 100410, 100280, 100240, 
    100220, 100160, 100130, 100100, 100030, 99970, 99920, 99960, 99880, 
    99890, 99940, 99930, 99860, 99810, 99790, 99760, 99730, 99680, 99700, 
    99660, 99660, 99700, 99670, 99640, 99630, 99640, 99620, 99600, 99580, 
    99560, 99550, 99540, 99550, 99570, 99540, 99550, 99570, 99580, 99580, 
    99600, 99600, 99650, 99680, 99710, 99750, 99780, 99830, 99870, 99900, 
    99940, 99990, 100030, 100070, 100120, 100150, 100200, 100240, 100270, 
    100310, 100320, 100340, 100360, 100360, 100360, 100370, 100380, 100420, 
    100430, 100450, 100490, 100540, 100600, 100670, 100730, 100780, 100810, 
    100870, 100930, 100990, 101040, 101060, 101100, 101160, 101200, 101200, 
    101220, 101250, 101290, 101330, 101360, 101400, 101430, 101470, 101520, 
    101570, 101580, 101610, 101660, 101670, 101700, 101750, 101730, 101780, 
    101840, 101870, 101890, 101930, 101980, 101990, 102000, 102030, 102040, 
    102040, 102070, 102110, 102140, 102150, 102170, 102200, 102180, 102190, 
    102150, 102160, 102150, 102120, 102080, 102050, 102010, 101990, 102070, 
    102030, 101790, 101740, 101790, 101720, 101680, 101420, 101400, 101250, 
    101060, 100880, 100860, 100780, 100780, 100700, 100530, 100490, 100390, 
    100420, 100390, 100390, 100340, 100450, 100460, 100460, 100420, 100320, 
    100210, 100090, 99990, 99920, 99870, 99900, 99970, 100120, 100240, 
    100370, 100480, 100560, 100590, 100640, 100660, 100690, 100800, 100870, 
    100910, 100950, 101010, 101050, 101070, 101090, 101110, 101110, 101130, 
    101160, 101140, 101150, 101170, 101200, 101230, 101220, 101200, 101190, 
    101190, 101180, 101190, 101190, 101200, 101200, 101200, 101200, 101220, 
    101220, 101220, 101220, 101260, 101260, 101290, 101320, 101340, 101350, 
    101410, 101470, 101510, 101540, 101580, 101610, 101600, 101630, 101650, 
    101660, 101650, 101660, 101670, 101670, 101670, 101710, 101700, 101710, 
    101710, 101710, 101700, 101730, 101740, 101740, 101780, 101780, 101780, 
    101790, 101810, 101780, 101790, 101770, 101750, 101730, 101740, 101730, 
    101740, 101720, 101700, 101690, 101670, 101670, 101660, 101610, 101580, 
    101560, 101560, 101540, 101520, 101520, 101500, 101500, 101490, 101470, 
    101440, 101430, 101410, 101420, 101420, 101410, 101410, 101410, 101390, 
    101380, 101380, 101380, 101350, 101350, 101340, 101340, 101350, 101350, 
    101340, 101330, 101350, 101350, 101360, 101330, 101320, 101300, 101300, 
    101250, 101220, 101200, 101190, 101180, 101160, 101150, 101140, 101130, 
    101120, 101110, 101100, 101100, 101100, 101090, 101090, 101110, 101110, 
    101110, 101120, 101120, 101130, 101130, 101130, 101130, 101150, 101160, 
    101180, 101170, 101160, 101180, 101200, 101210, 101220, 101240, 101250, 
    101260, 101300, 101320, 101350, 101360, 101370, 101380, 101410, 101430, 
    101420, 101450, 101440, 101440, 101460, 101430, 101450, 101430, 101430, 
    101430, 101430, 101410, 101380, 101340, 101360, 101360, 101350, 101380, 
    101420, 101450, 101480, 101520, 101540, 101530, 101540, 101580, 101580, 
    101600, 101610, 101600, 101620, 101610, 101610, 101600, 101590, 101600, 
    101590, 101580, 101550, 101580, 101570, 101570, 101590, 101600, 101610, 
    101600, 101600, 101630, 101630, 101640, 101640, 101680, 101700, 101710, 
    101740, 101730, 101720, 101730, 101730, 101740, 101710, 101730, 101700, 
    101680, 101640, 101560, 101550, 101530, 101500, 101450, 101450, 101430, 
    101390, 101410, 101390, 101360, 101370, 101360, 101360, 101340, 101370, 
    101370, 101330, 101350, 101300, 101240, 101180, 101120, 101120, 101140, 
    101100, 101100, 101000, 100960, 100950, 100780, 100690, 100590, 100550, 
    100350, 100340, 100380, 100360, 100330, 100450, 100460, 100440, 100420, 
    100440, 100440, 100440, 100500, 100530, 100580, 100630, 100680, 100750, 
    100810, 100850, 100890, 100960, 100980, 101040, 101080, 101140, 101170, 
    101220, 101270, 101320, 101340, 101350, 101390, 101460, 101480, 101510, 
    101550, 101600, 101640, 101660, 101680, 101720, 101730, 101740, 101750, 
    101760, 101750, 101740, 101750, 101760, 101740, 101750, 101740, 101750, 
    101740, 101750, 101740, 101710, 101730, 101730, 101760, 101720, 101730, 
    101790, 101790, 101770, 101740, 101750, 101730, 101730, 101760, 101750, 
    101740, 101740, 101740, 101720, 101710, 101740, 101720, 101720, 101710, 
    101660, 101680, 101660, 101640, 101620, 101620, 101630, 101620, 101610, 
    101640, 101620, 101620, 101630, 101600, 101640, 101680, 101660, 101680, 
    101700, 101730, 101780, 101850, 101860, 101860, 101850, 101870, 101880, 
    101880, 101880, 101900, 101900, 101900, 101870, 101860, 101830, 101830, 
    101800, 101770, 101730, 101710, 101690, 101670, 101640, 101600, 101570, 
    101540, 101510, 101470, 101440, 101410, 101380, 101360, 101330, 101270, 
    101230, 101190, 101150, 101100, 101040, 100960, 100900, 100830, 100770, 
    100670, 100580, 100540, 100540, 100520, 100500, 100500, 100510, 100530, 
    100530, 100550, 100570, 100710, 100730, 100810, 100840, 100890, 100970, 
    101000, 101040, 101070, 101070, 101070, 101030, 101020, 101040, 101010, 
    100980, 100980, 100960, 100930, 100910, 100880, 100860, 100810, 100760, 
    100750, 100740, 100720, 100710, 100700, 100670, 100660, 100660, 100630, 
    100610, 100600, 100570, 100530, 100500, 100460, 100460, 100440, 100410, 
    100330, 100280, 100200, 100090, 100020, 100000, 99950, 99890, 99840, 
    99800, 99780, 99790, 99830, 99840, 99900, 99910, 99930, 99970, 100000, 
    100040, 100070, 100080, 100110, 100100, 100080, 100080, 100050, 100040, 
    100010, 100000, 99990, 99980, 99960, 99980, 100020, 100020, 100020, 
    99980, 99950, 99900, 99830, 99800, 99760, 99730, 99660, 99610, 99550, 
    99520, 99520, 99490, 99460, 99450, 99420, 99420, 99430, 99460, 99520, 
    99540, 99560, 99610, 99610, 99580, 99570, 99600, 99600, 99550, 99570, 
    99530, 99520, 99530, 99510, 99480, 99520, 99550, 99570, 99600, 99660, 
    99690, 99740, 99800, 99840, 99870, 99880, 99930, 99950, 99950, 99970, 
    99980, 99960, 99940, 99960, 99950, 99930, 99900, 99900, 99930, 99940, 
    99970, 100010, 100090, 100160, 100240, 100280, 100360, 100420, 100510, 
    100570, 100630, 100690, 100710, 100710, 100700, 100660, 100560, 100470, 
    100400, 100310, 100190, 100110, 100010, 99970, 99910, 99920, 99940, 
    99940, 99970, 100030, 100070, 100170, 100240, 100320, 100370, 100410, 
    100430, 100480, 100510, 100500, 100530, 100510, 100530, 100520, 100530, 
    100500, 100480, 100450, 100460, 100440, 100420, 100430, 100430, 100450, 
    100440, 100490, 100500, 100510, 100530, 100540, 100550, 100580, 100610, 
    100640, 100630, 100630, 100640, 100650, 100670, 100670, 100660, 100660, 
    100710, 100680, 100700, 100720, 100720, 100750, 100760, 100790, 100830, 
    100830, 100870, 100900, 100950, 100980, 101020, 101040, 101040, 101090, 
    101100, 101110, 101150, 101190, 101200, 101240, 101280, 101300, 101300, 
    101330, 101340, 101340, 101380, 101410, 101430, 101430, 101440, 101440, 
    101430, 101420, 101370, 101360, 101290, 101250, 101170, 101110, 101090, 
    101040, 101010, 100990, 100950, 100930, 100930, 100910, 100900, 100900, 
    100900, 100920, 100950, 100940, 100950, 100940, 100910, 100860, 100810, 
    100800, 100820, 100740, 100730, 100720, 100720, 100690, 100700, 100700, 
    100680, 100630, 100550, 100550, 100480, 100370, 100270, 100240, 100230, 
    100190, 100220, 100210, 100200, 100160, 100130, 100060, 100010, 99910, 
    99760, 99740, 99760, 99840, 99950, 100040, 100070, 100120, 100190, 
    100260, 100320, 100400, 100400, 100420, 100480, 100500, 100570, 100590, 
    100610, 100670, 100660, 100640, 100630, 100640, 100630, 100580, 100540, 
    100550, 100590, 100590, 100580, 100550, 100620, 100610, 100620, 100620, 
    100640, 100640, 100640, 100660, 100700, 100730, 100730, 100760, 100760, 
    100770, 100780, 100780, 100770, 100780, 100760, 100760, 100760, 100770, 
    100780, 100810, 100820, 100840, 100830, 100810, 100820, 100840, 100840, 
    100840, 100860, 100880, 100870, 100830, 100810, 100780, 100750, 100720, 
    100680, 100680, 100700, 100700, 100700, 100710, 100750, 100790, 100830, 
    100900, 100930, 100990, 101070, 101140, 101190, 101260, 101320, 101370, 
    101430, 101460, 101510, 101540, 101600, 101670, 101710, 101740, 101800, 
    101820, 101820, 101870, 101930, 101940, 101980, 102000, 102000, 102000, 
    102010, 102020, 102040, 102040, 102050, 102020, 101990, 101950, 101890, 
    101850, 101800, 101780, 101730, 101710, 101670, 101620, 101570, 101520, 
    101420, 101360, 101290, 101220, 101170, 101130, 101050, 100990, 100950, 
    100910, 100870, 100850, 100790, 100710, 100690, 100610, 100570, 100530, 
    100490, 100400, 100400, 100380, 100350, 100320, 100290, 100270, 100240, 
    100220, 100250, 100230, 100230, 100250, 100250, 100270, 100260, 100240, 
    100280, 100280, 100340, 100330, 100320, 100340, 100340, 100330, 100330, 
    100320, 100300, 100250, 100190, 100160, 100140, 100110, 100080, 100110, 
    100140, 100130, 100120, 100060, 100060, 100100, 100110, 100110, 100100, 
    100080, 100060, 100060, 99990, 99930, 99890, 99860, 99800, 99710, 99660, 
    99600, 99490, 99480, 99470, 99470, 99420, 99270, 99190, 99200, 99140, 
    99120, 99060, 99040, 99020, 98990, 98880, 98810, 98920, 98950, 98970, 
    98980, 99050, 99100, 99170, 99210, 99290, 99310, 99340, 99430, 99500, 
    99550, 99600, 99690, 99810, 99920, 100040, 100080, 100150, 100250, 
    100290, 100350, 100410, 100460, 100480, 100520, 100560, 100590, 100600, 
    100670, 100720, 100740, 100740, 100740, 100800, 100830, 100870, 100900, 
    100900, 100950, 101000, 101010, 100990, 101020, 101040, 101090, 101170, 
    101200, 101180, 101180, 101200, 101230, 101250, 101230, 101220, 101210, 
    101210, 101240, 101280, 101320, 101330, 101340, 101380, 101390, 101390, 
    101380, 101390, 101390, 101370, 101360, 101350, 101370, 101380, 101390, 
    101390, 101400, 101400, 101410, 101380, 101370, 101380, 101390, 101380, 
    101400, 101410, 101420, 101430, 101450, 101470, 101510, 101510, 101520, 
    101520, 101520, 101520, 101510, 101480, 101510, 101510, 101530, 101530, 
    101520, 101500, 101480, 101470, 101490, 101490, 101500, 101510, 101530, 
    101540, 101550, 101550, 101540, 101530, 101530, 101510, 101500, 101450, 
    101440, 101430, 101400, 101380, 101350, 101320, 101290, 101280, 101250, 
    101230, 101230, 101200, 101200, 101160, 101150, 101120, 101110, 101120, 
    101110, 101090, 101050, 101010, 100990, 100960, 100930, 100950, 100910, 
    100890, 100840, 100850, 100780, 100740, 100670, 100660, 100600, 100590, 
    100550, 100520, 100440, 100390, 100330, 100260, 100170, 100150, 100130, 
    100120, 100070, 100070, 100040, 100010, 100000, 99960, 99920, 99880, 
    99870, 99870, 99830, 99820, 99800, 99830, 99850, 99860, 99860, 99860, 
    99880, 99860, 99890, 99890, 99880, 99900, 99920, 99950, 99950, 99950, 
    99980, 99960, 99950, 99890, 99830, 99770, 99740, 99700, 99660, 99610, 
    99630, 99610, 99630, 99680, 99760, 99810, 99890, 99990, 100070, 100160, 
    100240, 100320, 100350, 100370, 100400, 100390, 100380, 100360, 100340, 
    100290, 100280, 100250, 100240, 100210, 100190, 100180, 100190, 100220, 
    100230, 100320, 100340, 100390, 100480, 100530, 100590, 100640, 100670, 
    100720, 100760, 100770, 100790, 100780, 100780, 100730, 100690, 100650, 
    100670, 100660, 100630, 100650, 100660, 100710, 100720, 100810, 100890, 
    100920, 100980, 101060, 101140, 101180, 101250, 101320, 101330, 101350, 
    101390, 101430, 101410, 101390, 101550, 101620, 101660, 101690, 101680, 
    101700, 101770, 101800, 101810, 101820, 101830, 101810, 101770, 101720, 
    101690, 101670, 101600, 101560, 101520, 101450, 101380, 101290, 101220, 
    101110, 101020, 100980, 100920, 100880, 100770, 100730, 100670, 100570, 
    100530, 100270, 100210, 100200, 100210, 100200, 100210, 100180, 100200, 
    100190, 100210, 100230, 100210, 100280, 100280, 100330, 100420, 100430, 
    100490, 100550, 100630, 100670, 100760, 100850, 100910, 100960, 101030, 
    101120, 101120, 101120, 101180, 101230, 101290, 101310, 101340, 101410, 
    101440, 101450, 101460, 101480, 101500, 101540, 101520, 101550, 101580, 
    101610, 101620, 101640, 101660, 101610, 101590, 101620, 101540, 101510, 
    101430, 101400, 101340, 101230, 101170, 101140, 101050, 101010, 100920, 
    100850, 100790, 100690, 100700, 100660, 100660, 100650, 100680, 100670, 
    100670, 100710, 100740, 100720, 100760, 100770, 100810, 100810, 100840, 
    100830, 100820, 100800, 100760, 100730, 100690, 100690, 100670, 100680, 
    100680, 100700, 100730, 100750, 100800, 100810, 100870, 100900, 100930, 
    100930, 100930, 100940, 100960, 100990, 100990, 101010, 101040, 101080, 
    101140, 101180, 101220, 101260, 101310, 101360, 101420, 101500, 101550, 
    101600, 101630, 101690, 101730, 101770, 101800, 101860, 101890, 101910, 
    101920, 101960, 101970, 102000, 102010, 102020, 102010, 102000, 101980, 
    101960, 101920, 101910, 101860, 101800, 101760, 101730, 101710, 101650, 
    101630, 101610, 101530, 101510, 101470, 101450, 101440, 101440, 101470, 
    101490, 101500, 101510, 101520, 101550, 101550, 101550, 101540, 101530, 
    101530, 101540, 101580, 101610, 101610, 101640, 101600, 101580, 101540, 
    101550, 101570, 101580, 101600, 101610, 101660, 101680, 101710, 101740, 
    101750, 101790, 101830, 101880, 101900, 101940, 102000, 102030, 102050, 
    102100, 102130, 102170, 102200, 102210, 102250, 102290, 102300, 102320, 
    102350, 102390, 102420, 102430, 102450, 102440, 102460, 102490, 102510, 
    102510, 102530, 102550, 102540, 102550, 102570, 102590, 102600, 102630, 
    102640, 102670, 102690, 102700, 102730, 102760, 102770, 102760, 102770, 
    102710, 102680, 102740, 102730, 102760, 102740, 102790, 102830, 102850, 
    102860, 102870, 102890, 102910, 102950, 102970, 102990, 103020, 103020, 
    103050, 103050, 103050, 103070, 103070, 103100, 103110, 103120, 103140, 
    103140, 103150, 103160, 103160, 103170, 103160, 103170, 103170, 103180, 
    103170, 103200, 103210, 103230, 103240, 103250, 103260, 103290, 103290, 
    103290, 103320, 103330, 103360, 103360, 103380, 103380, 103380, 103410, 
    103400, 103420, 103420, 103440, 103430, 103450, 103460, 103460, 103490, 
    103490, 103500, 103480, 103470, 103470, 103480, 103480, 103470, 103460, 
    103450, 103450, 103480, 103460, 103460, 103450, 103440, 103450, 103410, 
    103410, 103420, 103440, 103460, 103460, 103450, 103450, 103420, 103400, 
    103400, 103390, 103370, 103380, 103360, 103350, 103330, 103330, 103330, 
    103330, 103310, 103310, 103310, 103300, 103310, 103300, 103270, 103290, 
    103300, 103320, 103330, 103350, 103350, 103320, 103300, 103300, 103290, 
    103300, 103300, 103280, 103280, 103260, 103250, 103240, 103220, 103210, 
    103210, 103240, 103230, 103230, 103210, 103210, 103220, 103240, 103260, 
    103260, 103270, 103260, 103250, 103240, 103260, 103260, 103270, 103250, 
    103260, 103260, 103270, 103260, 103270, 103240, 103240, 103250, 103230, 
    103240, 103230, 103240, 103260, 103250, 103260, 103290, 103290, 103280, 
    103270, 103250, 103220, 103210, 103220, 103200, 103200, 103200, 103220, 
    103200, 103190, 103190, 103190, 103170, 103140, 103130, 103120, 103110, 
    103100, 103090, 103080, 103130, 103100, 103080, 103070, 103040, 103000, 
    102980, 102960, 102950, 102950, 102930, 102910, 102920, 102900, 102880, 
    102860, 102830, 102810, 102790, 102780, 102790, 102800, 102790, 102790, 
    102780, 102760, 102730, 102710, 102680, 102660, 102630, 102610, 102590, 
    102540, 102530, 102540, 102500, 102500, 102480, 102460, 102420, 102390, 
    102370, 102330, 102330, 102340, 102330, 102310, 102290, 102250, 102200, 
    102130, 102060, 102010, 101940, 101880, 101770, 101660, 101590, 101470, 
    101370, 101310, 101190, 101080, 100970, 100860, 100730, 100570, 100490, 
    100380, 100270, 100150, 100050, 99900, 99780, 99700, 99600, 99540, 99490, 
    99430, 99370, 99300, 99220, 99160, 99110, 99060, 99080, 99190, 99290, 
    99390, 99460, 99560, 99660, 99710, 99740, 99740, 99700, 99640, 99570, 
    99480, 99410, 99330, 99230, 99070, 98900, 98650, 98340, 98080, 98030, 
    97960, 98000, 98010, 98200, 98320, 98470, 98610, 98730, 98820, 98840, 
    98840, 98800, 98780, 98790, 98860, 98940, 98980, 99030, 99080, 99120, 
    99150, 99130, 99140, 99150, 99240, 99290, 99330, 99350, 99390, 99430, 
    99480, 99520, 99570, 99600, 99640, 99640, 99730, 99750, 99790, 99850, 
    99870, 99910, 99930, 99970, 100000, 100030, 100060, 100080, 100100, 
    100130, 100220, 100290, 100370, 100400, 100490, 100570, 100630, 100700, 
    100770, 100830, 100880, 100900, 100940, 100940, 100990, 101020, 101040, 
    101080, 101100, 101140, 101190, 101220, 101240, 101290, 101310, 101330, 
    101350, 101370, 101400, 101420, 101460, 101480, 101520, 101520, 101550, 
    101560, 101580, 101600, 101620, 101620, 101650, 101650, 101670, 101700, 
    101720, 101760, 101770, 101780, 101800, 101830, 101840, 101860, 101850, 
    101870, 101890, 101930, 101950, 101980, 101990, 101990, 101990, 101990, 
    101990, 101990, 102000, 102000, 101990, 101980, 101990, 101980, 101950, 
    101940, 101920, 101900, 101900, 101870, 101860, 101860, 101880, 101880, 
    101880, 101860, 101830, 101820, 101790, 101770, 101730, 101700, 101680, 
    101650, 101630, 101590, 101570, 101540, 101520, 101490, 101460, 101440, 
    101410, 101390, 101360, 101360, 101350, 101320, 101300, 101250, 101220, 
    101170, 101150, 101110, 101070, 101060, 101020, 100990, 100950, 100890, 
    100850, 100780, 100720, 100650, 100530, 100420, 100290, 100200, 100180, 
    100130, 100120, 100090, 100080, 100060, 100030, 99990, 99960, 99920, 
    99880, 99820, 99810, 99780, 99730, 99700, 99650, 99570, 99530, 99520, 
    99510, 99470, 99480, 99490, 99550, 99600, 99620, 99630, 99690, 99790, 
    99820, 99820, 99880, 99910, 99960, 99980, 100010, 100040, 100090, 100110, 
    100170, 100200, 100210, 100210, 100290, 100320, 100330, 100330, 100340, 
    100350, 100340, 100360, 100410, 100470, 100520, 100600, 100700, 100810, 
    100910, 101000, 101120, 101260, 101420, 101560, 101690, 101820, 101890, 
    101960, 102020, 102070, 102120, 102140, 102160, 102180, 102200, 102190, 
    102200, 102210, 102190, 102190, 102160, 102140, 102110, 102080, 102070, 
    102040, 102020, 102000, 101980, 101960, 101930, 101910, 101880, 101850, 
    101820, 101810, 101770, 101770, 101790, 101780, 101750, 101710, 101730, 
    101710, 101680, 101680, 101660, 101650, 101630, 101630, 101660, 101680, 
    101700, 101720, 101740, 101730, 101750, 101760, 101790, 101770, 101780, 
    101810, 101840, 101880, 101880, 101900, 101920, 101910, 101930, 101910, 
    101910, 101910, 101900, 101900, 101880, 101870, 101840, 101800, 101770, 
    101730, 101700, 101660, 101620, 101580, 101480, 101460, 101420, 101370, 
    101310, 101260, 101200, 101130, 101060, 100990, 100920, 100880, 100830, 
    100780, 100750, 100710, 100680, 100640, 100650, 100660, 100670, 100670, 
    100680, 100680, 100690, 100720, 100750, 100780, 100820, 100860, 100880, 
    100890, 100890, 100910, 100920, 100940, 100960, 100990, 101040, 101060, 
    101080, 101100, 101140, 101140, 101150, 101180, 101200, 101250, 101300, 
    101310, 101350, 101420, 101480, 101530, 101550, 101590, 101610, 101650, 
    101660, 101670, 101680, 101700, 101720, 101740, 101750, 101740, 101730, 
    101710, 101710, 101700, 101700, 101710, 101710, 101730, 101770, 101780, 
    101800, 101810, 101800, 101790, 101780, 101800, 101800, 101810, 101820, 
    101820, 101830, 101820, 101820, 101810, 101800, 101800, 101780, 101750, 
    101720, 101690, 101670, 101650, 101650, 101630, 101610, 101570, 101520, 
    101490, 101460, 101420, 101380, 101360, 101320, 101270, 101230, 101210, 
    101180, 101110, 101050, 101000, 100940, 100900, 100850, 100770, 100700, 
    100620, 100520, 100410, 100290, 100190, 100090, 100110, 100120, 100160, 
    100140, 100130, 100140, 100130, 100100, 100100, 100090, 100070, 100030, 
    100000, 99980, 99990, 99990, 99960, 99940, 99890, 99840, 99800, 99720, 
    99650, 99610, 99620, 99610, 99610, 99650, 99710, 99750, 99790, 99830, 
    99900, 99940, 99970, 99990, 100000, 100030, 100040, 100040, 100050, 
    100080, 100080, 100110, 100120, 100140, 100140, 100110, 100100, 100060, 
    100040, 100030, 100010, 99990, 99960, 99960, 99920, 99890, 99850, 99800, 
    99770, 99730, 99760, 99760, 99710, 99670, 99680, 99680, 99700, 99720, 
    99740, 99740, 99730, 99710, 99720, 99700, 99660, 99680, 99670, 99700, 
    99690, 99690, 99670, 99660, 99640, 99620, 99600, 99570, 99550, 99540, 
    99550, 99580, 99590, 99600, 99610, 99570, 99560, 99570, 99750, 99620, 
    99630, 99620, 99620, 99600, 99600, 99600, 99610, 99640, 99660, 99650, 
    99650, 99680, 99690, 99700, 99740, 99760, 99790, 99820, 99820, 99820, 
    99830, 99870, 99920, 99950, 99970, 100000, 100030, 100090, 100140, 
    100180, 100200, 100240, 100250, 100260, 100270, 100280, 100300, 100300, 
    100320, 100370, 100410, 100460, 100490, 100500, 100520, 100530, 100540, 
    100530, 100540, 100560, 100560, 100590, 100590, 100590, 100600, 100590, 
    100580, 100600, 100570, 100590, 100570, 100600, 100610, 100620, 100620, 
    100630, 100640, 100660, 100670, 100640, 100640, 100650, 100660, 100670, 
    100680, 100700, 100720, 100730, 100730, 100750, 100760, 100760, 100760, 
    100780, 100780, 100810, 100810, 100850, 100870, 100860, 100880, 100860, 
    100850, 100860, 100860, 100870, 100890, 100870, 100870, 100880, 100890, 
    100880, 100880, 100880, 100860, 100850, 100840, 100810, 100800, 100780, 
    100770, 100780, 100770, 100760, 100750, 100740, 100700, 100700, 100690, 
    100660, 100650, 100650, 100640, 100640, 100640, 100670, 100700, 100720, 
    100730, 100750, 100740, 100740, 100780, 100750, 100790, 100810, 100840, 
    100860, 100880, 100900, 100930, 100950, 100920, 100940, 100960, 100970, 
    101010, 101040, 101080, 101110, 101110, 101130, 101160, 101170, 101180, 
    101180, 101190, 101190, 101200, 101230, 101260, 101290, 101310, 101300, 
    101330, 101300, 101290, 101260, 101250, 101240, 101220, 101230, 101190, 
    101190, 101160, 101130, 101110, 101120, 101090, 101050, 101000, 100950, 
    100930, 100920, 100910, 100860, 100780, 100760, 100710, 100630, 100530, 
    100330, 100310, 100170, 100100, 100070, 100000, 99860, 99710, 99550, 
    99390, 99290, 99210, 99060, 98940, 98820, 98670, 98630, 98620, 98670, 
    98630, 98620, 98600, 98570, 98510, 98490, 98460, 98450, 98440, 98440, 
    98440, 98460, 98490, 98520, 98610, 98670, 98710, 98840, 98950, 99080, 
    99230, 99370, 99440, 99470, 99630, 99640, 99690, 99790, 99860, 99930, 
    99950, 99950, 99940, 99710, 99710, 99690, 99570, 99440, 99500, 99380, 
    99360, 99340, 99200, 99000, 98900, 98830, 98860, 98760, 98780, 98700, 
    98560, 98470, 98380, 98260, 98160, 98060, 98000, 97920, 97890, 97830, 
    97820, 97820, 97790, 97720, 97670, 97590, 97540, 97540, 97590, 97650, 
    97770, 97850, 97890, 97920, 97950, 97990, 98020, 98050, 98050, 98090, 
    98080, 98080, 98080, 98080, 98050, 98030, 98050, 98050, 98050, 98080, 
    98090, 98120, 98110, 98110, 98120, 98100, 98090, 98070, 98060, 98040, 
    98000, 97990, 97960, 97940, 97950, 97970, 97980, 98010, 98050, 98080, 
    98060, 98120, 98190, 98220, 98300, 98320, 98430, 98520, 98610, 98690, 
    98820, 98890, 98990, 99100, 99230, 99300, 99400, 99520, 99620, 99740, 
    99820, 99890, 99940, 100000, 100060, 100120, 100110, 100140, 100170, 
    100190, 100200, 100200, 100170, 100220, 100200, 100170, 100140, 100090, 
    100050, 99990, 99920, 99970, 99910, 99870, 99860, 99840, 99790, 99770, 
    99730, 99700, 99670, 99610, 99610, 99640, 99670, 99690, 99680, 99690, 
    99670, 99650, 99600, 99580, 99560, 99530, 99500, 99460, 99440, 99400, 
    99370, 99310, 99260, 99180, 99110, 98940, 98930, 98830, 98740, 98700, 
    98660, 98660, 98660, 98680, 98710, 98750, 98770, 98810, 98820, 98810, 
    98780, 98830, 98850, 98950, 98990, 99000, 99050, 99050, 99060, 99040, 
    99030, 99010, 99000, 98990, 98990, 99020, 99060, 99060, 99050, 99030, 
    98960, 98920, 98870, 98800, 98750, 98710, 98680, 98640, 98630, 98630, 
    98660, 98650, 98600, 98630, 98720, 98790, 98890, 99000, 99100, 99180, 
    99230, 99330, 99380, 99450, 99480, 99570, 99620, 99720, 99750, 99790, 
    99840, 99890, 99940, 99960, 99980, 100040, 100090, 100110, 100150, 
    100170, 100220, 100220, 100250, 100340, 100360, 100380, 100450, 100490, 
    100540, 100520, 100550, 100530, 100510, 100470, 100420, 100350, 100280, 
    100250, 100120, 100030, 99920, 99790, 99660, 99520, 99380, 99230, 99040, 
    98830, 98620, 98370, 98090, 97810, 97490, 97310, 97130, 96940, 96790, 
    96690, 96610, 96600, 96630, 96670, 96660, 96660, 96650, 96660, 96660, 
    96690, 96700, 96720, 96760, 96880, 96940, 96990, 97040, 97060, 97090, 
    97100, 97110, 97090, 97060, 97020, 96990, 96960, 96840, 96850, 96800, 
    96770, 96740, 96750, 96750, 96750, 96810, 96740, 96700, 96700, 96750, 
    96860, 97020, 97180, 97340, 97500, 97590, 97710, 97810, 97880, 97970, 
    98040, 98090, 98160, 98180, 98200, 98230, 98280, 98300, 98360, 98400, 
    98490, 98530, 98600, 98640, 98690, 98690, 98710, 98710, 98720, 98730, 
    98730, 98760, 98760, 98760, 98760, 98780, 98790, 98770, 98760, 98750, 
    98730, 98700, 98710, 98720, 98730, 98760, 98800, 98820, 98860, 98900, 
    98900, 98910, 98940, 98970, 99010, 99070, 99130, 99180, 99240, 99320, 
    99350, 99370, 99390, 99410, 99440, 99470, 99480, 99480, 99470, 99470, 
    99490, 99480, 99480, 99470, 99480, 99490, 99520, 99540, 99570, 99600, 
    99610, 99620, 99670, 99710, 99750, 99770, 99800, 99840, 99870, 99900, 
    99930, 99950, 99980, 100020, 100080, 100120, 100130, 100160, 100190, 
    100220, 100240, 100260, 100260, 100270, 100270, 100250, 100180, 100180, 
    100180, 100130, 100070, 100040, 100010, 99970, 99940, 99890, 99850, 
    99830, 99860, 99880, 99860, 99860, 99830, 99790, 99720, 99740, 99700, 
    99630, 99560, 99490, 99440, 99380, 99350, 99320, 99290, 99240, 99220, 
    99180, 99060, 98970, 98850, 98730, 98640, 98620, 98570, 98620, 98660, 
    98690, 98760, 98790, 98790, 98720, 98790, 98860, 98970, 99040, 99080, 
    99170, 99200, 99200, 99220, 99270, 99350, 99390, 99440, 99470, 99500, 
    99530, 99590, 99610, 99630, 99640, 99690, 99740, 99810, 99840, 99860, 
    99870, 99900, 99940, 99960, 100020, 100020, 100010, 100020, 100060, 
    100070, 100110, 100110, 100130, 100140, 100140, 100150, 100190, 100220, 
    100220, 100210, 100230, 100260, 100280, 100270, 100280, 100280, 100260, 
    100280, 100280, 100300, 100280, 100250, 100230, 100210, 100180, 100180, 
    100140, 100140, 100140, 100130, 100110, 100100, 100070, 100050, 100030, 
    99990, 99980, 99960, 99970, 99980, 99970, 99990, 99970, 99940, 99910, 
    99880, 99850, 99840, 99800, 99800, 99760, 99770, 99770, 99760, 99780, 
    99770, 99790, 99790, 99790, 99800, 99810, 99830, 99870, 99900, 99920, 
    99940, 99970, 99980, 99990, 100020, 100050, 100060, 100080, 100100, 
    100130, 100200, 100180, 100190, 100170, 100160, 100140, 100120, 100100, 
    100080, 100080, 100070, 100020, 100010, 99980, 99920, 99880, 99830, 
    99780, 99720, 99660, 99590, 99480, 99400, 99360, 99310, 99240, 99170, 
    99090, 99000, 98930, 98890, 98830, 98780, 98750, 98700, 98650, 98600, 
    98590, 98570, 98540, 98530, 98520, 98500, 98480, 98460, 98420, 98430, 
    98450, 98460, 98480, 98500, 98490, 98510, 98510, 98560, 98580, 98600, 
    98610, 98620, 98620, 98600, 98650, 98680, 98680, 98690, 98720, 98780, 
    98840, 98900, 98940, 98980, 99020, 99070, 99080, 99110, 99130, 99130, 
    99120, 99110, 99130, 99140, 99160, 99130, 99140, 99200, 99210, 99210, 
    99240, 99240, 99240, 99260, 99260, 99270, 99270, 99280, 99280, 99270, 
    99310, 99290, 99260, 99260, 99280, 99260, 99270, 99270, 99250, 99220, 
    99220, 99180, 99150, 99090, 99040, 99000, 98980, 98930, 98910, 98880, 
    98860, 98840, 98810, 98790, 98780, 98770, 98790, 98790, 98790, 98790, 
    98840, 98850, 98870, 98890, 98910, 98950, 98980, 99020, 99060, 99070, 
    99100, 99120, 99160, 99190, 99210, 99240, 99260, 99280, 99340, 99350, 
    99370, 99410, 99430, 99460, 99470, 99480, 99510, 99540, 99560, 99560, 
    99580, 99610, 99630, 99620, 99630, 99660, 99700, 99700, 99680, 99690, 
    99720, 99730, 99780, 99830, 99770, 99840, 99870, 99910, 99950, 99980, 
    100060, 100080, 100090, 100120, 100170, 100210, 100240, 100250, 100290, 
    100330, 100310, 100290, 100300, 100330, 100360, 100390, 100400, 100430, 
    100450, 100410, 100390, 100370, 100390, 100360, 100360, 100360, 100360, 
    100350, 100350, 100350, 100350, 100310, 100330, 100310, 100300, 100290, 
    100280, 100310, 100320, 100330, 100300, 100330, 100310, 100300, 100290, 
    100290, 100310, 100280, 100270, 100270, 100300, 100320, 100310, 100340, 
    100310, 100300, 100310, 100300, 100370, 100350, 100370, 100380, 100350, 
    100360, 100290, 100320, 100380, 100380, 100410, 100440, 100460, 100510, 
    100530, 100530, 100550, 100590, 100640, 100670, 100690, 100750, 100800, 
    100840, 100860, 100890, 100900, 100950, 100990, 101040, 101040, 101090, 
    101100, 101150, 101160, 101160, 101190, 101200, 101220, 101180, 101160, 
    101170, 101190, 101160, 101180, 101150, 101170, 101180, 101190, 101210, 
    101170, 101180, 101230, 101250, 101250, 101270, 101290, 101300, 101290, 
    101310, 101330, 101290, 101280, 101270, 101220, 101190, 101210, 101160, 
    101100, 101050, 100970, 100910, 100820, 100730, 100640, 100530, 100390, 
    100300, 100200, 100010, 99900, 99780, 99700, 99580, 99550, 99400, 99340, 
    99290, 99300, 99270, 99240, 99220, 99210, 99190, 99170, 99110, 99150, 
    99190, 99230, 99350, 99410, 99560, 99590, 99590, 99650, 99690, 99730, 
    99770, 99800, 99890, 99990, 100080, 100170, 100230, 100310, 100350, 
    100390, 100460, 100520, 100560, 100600, 100630, 100640, 100670, 100730, 
    100780, 100810, 100810, 100840, 100900, 100920, 100960, 100970, 100940, 
    100930, 100960, 100980, 100980, 101000, 100970, 100920, 100880, 100790, 
    100720, 100640, 100590, 100520, 100430, 100430, 100340, 100280, 100220, 
    100110, 100080, 100040, 100000, 100010, 99990, 100010, 99980, 99990, 
    100010, 100040, 100030, 100060, 100100, 100100, 100090, 100070, 100070, 
    100040, 100040, 100050, 100080, 100100, 100110, 100080, 100040, 100020, 
    99990, 99970, 99920, 99840, 99810, 99730, 99660, 99590, 99540, 99460, 
    99400, 99370, 99290, 99240, 99250, 99200, 99120, 99200, 99250, 99300, 
    99330, 99310, 99260, 99240, 99250, 99250, 99250, 99210, 99160, 99040, 
    98950, 98860, 98800, 98760, 98710, 98690, 98620, 98610, 98650, 98690, 
    98590, 98650, 98650, 98630, 98630, 98590, 98540, 98480, 98470, 98540, 
    98580, 98580, 98580, 98590, 98620, 98720, 98740, 98810, 98850, 98890, 
    98980, 99090, 99180, 99270, 99360, 99480, 99550, 99690, 99810, 99890, 
    99970, 100070, 100150, 100250, 100310, 100340, 100400, 100440, 100490, 
    100540, 100560, 100590, 100580, 100580, 100580, 100580, 100570, 100590, 
    100580, 100590, 100590, 100620, 100590, 100590, 100610, 100590, 100600, 
    100600, 100590, 100590, 100590, 100600, 100590, 100580, 100600, 100590, 
    100590, 100590, 100600, 100610, 100600, 100590, 100590, 100620, 100620, 
    100640, 100630, 100630, 100640, 100620, 100650, 100650, 100630, 100620, 
    100610, 100670, 100650, 100650, 100650, 100650, 100660, 100680, 100690, 
    100660, 100650, 100640, 100670, 100650, 100640, 100660, 100670, 100660, 
    100690, 100690, 100690, 100710, 100730, 100730, 100760, 100780, 100790, 
    100830, 100850, 100880, 100910, 100930, 100940, 100930, 101030, 101120, 
    101150, 101160, 101220, 101190, 101120, 101240, 101360, 101400, 101420, 
    101380, 101370, 101330, 101290, 101400, 101420, 101450, 101500, 101480, 
    101540, 101560, 101530, 101490, 101540, 101550, 101560, 101570, 101610, 
    101600, 101560, 101540, 101550, 101550, 101610, 101600, 101600, 101590, 
    101590, 101590, 101640, 101640, 101600, 101580, 101650, 101620, 101620, 
    101610, 101640, 101650, 101670, 101790, 101820, 101860, 101850, 101920, 
    101890, 101910, 101900, 101840, 101790, 101970, 101990, 101980, 102020, 
    102030, 102010, 102000, 102010, 102000, 101940, 101920, 101820, 101840, 
    101900, 101940, 101930, 101940, 101920, 101920, 101860, 101760, 101770, 
    101780, 101770, 101750, 101730, 101700, 101670, 101670, 101650, 101610, 
    101540, 101500, 101410, 101290, 101260, 101260, 101260, 101300, 101240, 
    101240, 101210, 101200, 101130, 101090, 101050, 101020, 100950, 100960, 
    100930, 100930, 100940, 100950, 100960, 100920, 100900, 100920, 100910, 
    100940, 100960, 100970, 100970, 100980, 101010, 101080, 101100, 101070, 
    101080, 101080, 101060, 101050, 101030, 101030, 101040, 101060, 101080, 
    101060, 101070, 101090, 101100, 101080, 100960, 100970, 100970, 100940, 
    100970, 101010, 101020, 101050, 101030, 101020, 101000, 101000, 101030, 
    101040, 101030, 101050, 101040, 101070, 101080, 101110, 101130, 101150, 
    101170, 101200, 101200, 101230, 101230, 101240, 101260, 101280, 101320, 
    101360, 101390, 101420, 101410, 101440, 101430, 101460, 101510, 101480, 
    101460, 101480, 101500, 101520, 101600, 101610, 101640, 101680, 101720, 
    101760, 101800, 101820, 101850, 101880, 101910, 101960, 102020, 102050, 
    102060, 102050, 102060, 102100, 102080, 102090, 102120, 102140, 102140, 
    102150, 102200, 102170, 102180, 102190, 102160, 102160, 102150, 102190, 
    102170, 102140, 102130, 102170, 102190, 102200, 102200, 102170, 102180, 
    102170, 102160, 102160, 102150, 102150, 102150, 102180, 102180, 102180, 
    102160, 102170, 102130, 102120, 102100, 102090, 102080, 102100, 102100, 
    102090, 102110, 102110, 102090, 102050, 101990, 101950, 101850, 101830, 
    101830, 101820, 101800, 101770, 101760, 101810, 101780, 101800, 101800, 
    101820, 101840, 101860, 101880, 101900, 101930, 101970, 101990, 101990, 
    101990, 101980, 101960, 101960, 101960, 101920, 101900, 101900, 101900, 
    101890, 101870, 101850, 101840, 101780, 101750, 101750, 101750, 101750, 
    101770, 101800, 101850, 101860, 101880, 101890, 101910, 101890, 101900, 
    101900, 101900, 101890, 101900, 101880, 101910, 101920, 101920, 101950, 
    101940, 101940, 101930, 101910, 101910, 101930, 101920, 101930, 101950, 
    101980, 102010, 102040, 102010, 102000, 102020, 102010, 102020, 102030, 
    102030, 102040, 102070, 102070, 102120, 102150, 102140, 102130, 102120, 
    102140, 102150, 102160, 102180, 102190, 102230, 102270, 102300, 102300, 
    102310, 102330, 102340, 102350, 102360, 102370, 102380, 102390, 102400, 
    102440, 102430, 102430, 102430, 102450, 102460, 102460, 102480, 102500, 
    102490, 102520, 102540, 102570, 102590, 102600, 102600, 102620, 102640, 
    102650, 102660, 102670, 102650, 102660, 102690, 102700, 102720, 102720, 
    102740, 102740, 102740, 102730, 102750, 102760, 102760, 102790, 102800, 
    102840, 102870, 102900, 102890, 102880, 102900, 102870, 102850, 102860, 
    102840, 102870, 102780, 102780, 102800, 102820, 102820, 102770, 102730, 
    102750, 102710, 102680, 102910, 102760, 102780, 102770, 102800, 102800, 
    102770, 102730, 102720, 102680, 102610, 102580, 102600, 102580, 102580, 
    102560, 102530, 102500, 102490, 102460, 102410, 102380, 102300, 102300, 
    102290, 102290, 102250, 102200, 102200, 102130, 102100, 102050, 101990, 
    101830, 101800, 101780, 101690, 101530, 101450, 101410, 101370, 101280, 
    101150, 101090, 101030, 100960, 100880, 100840, 100820, 100800, 100810, 
    100800, 100780, 100780, 100780, 100770, 100760, 100770, 100790, 100770, 
    100770, 100800, 100810, 100850, 100870, 100810, 100800, 100860, 100810, 
    100790, 100790, 100780, 100790, 100800, 100790, 100810, 100820, 100810, 
    100780, 100790, 100800, 100790, 100790, 100810, 100810, 100830, 100870, 
    100860, 100880, 100880, 100920, 100930, 100960, 100970, 100970, 100990, 
    101030, 101050, 101120, 101140, 101180, 101210, 101220, 101250, 101290, 
    101320, 101360, 101400, 101430, 101460, 101500, 101560, 101600, 101620, 
    101630, 101660, 101680, 101710, 101720, 101740, 101750, 101750, 101770, 
    101810, 101820, 101810, 101780, 101770, 101750, 101740, 101730, 101700, 
    101690, 101690, 101740, 101780, 101890, 101960, 102010, 102060, 102120, 
    102210, 102300, 102380, 102440, 102460, 102520, 102540, 102570, 102580, 
    102590, 102570, 102550, 102570, 102540, 102510, 102490, 102480, 102440, 
    102430, 102400, 102330, 102260, 102190, 102140, 102080, 102020, 101950, 
    101920, 101920, 101910, 101920, 101940, 101930, 101910, 101920, 101890, 
    101870, 101860, 101870, 101870, 101860, 101840, 101850, 101840, 101850, 
    101840, 101810, 101770, 101720, 101710, 101690, 101660, 101630, 101650, 
    101640, 101660, 101660, 101630, 101600, 101520, 101450, 101390, 101330, 
    101300, 101260, 101200, 101160, 101120, 101100, 101090, 101110, 101080, 
    101080, 101070, 101060, 101040, 101070, 101070, 101090, 101110, 101100, 
    101110, 101090, 101060, 101070, 101060, 101040, 101000, 101010, 100990, 
    100990, 100970, 100990, 101010, 100990, 100970, 100940, 100910, 100870, 
    100830, 100760, 100750, 100740, 100720, 100740, 100720, 100720, 100810, 
    100880, 100960, 101000, 101070, 101120, 101140, 101200, 101240, 101320, 
    101340, 101350, 101370, 101370, 101390, 101440, 101470, 101550, 101580, 
    101590, 101640, 101690, 101680, 101750, 101820, 101860, 101870, 101890, 
    102000, 102030, 102040, 102110, 102150, 102170, 102220, 102230, 102240, 
    102240, 102250, 102250, 102250, 102260, 102260, 102280, 102280, 102250, 
    102220, 102170, 102140, 102070, 101960, 101880, 101790, 101680, 101630, 
    101550, 101450, 101380, 101270, 101220, 101180, 101120, 101070, 101070, 
    101090, 101110, 101090, 101070, 101090, 101110, 101180, 101240, 101310, 
    101420, 101510, 101590, 101650, 101690, 101740, 101770, 101820, 101820, 
    101850, 101840, 101830, 101810, 101740, 101720, 101650, 101610, 101600, 
    101540, 101500, 101460, 101390, 101320, 101260, 101180, 101070, 100980, 
    100930, 100870, 100800, 100730, 100700, 100670, 100630, 100630, 100650, 
    100620, 100620, 100620, 100660, 100680, 100730, 100790, 100840, 100890, 
    100930, 100980, 100990, 101040, 101120, 101170, 101230, 101280, 101350, 
    101380, 101400, 101440, 101480, 101520, 101550, 101580, 101620, 101640, 
    101660, 101680, 101730, 101740, 101750, 101760, 101790, 101800, 101770, 
    101750, 101780, 101730, 101700, 101700, 101720, 101730, 101780, 101800, 
    101810, 101790, 101820, 101840, 101870, 101890, 101920, 101970, 102040, 
    102090, 102160, 102220, 102280, 102350, 102420, 102450, 102540, 102580, 
    102650, 102710, 102730, 102790, 102820, 102940, 103010, 103010, 103020, 
    103050, 103090, 103120, 103120, 103110, 103150, 103200, 103200, 103180, 
    103180, 103180, 103180, 103170, 103230, 103320, 103370, 103410, 103470, 
    103530, 103560, 103570, 103590, 103620, 103630, 103630, 103610, 103570, 
    103600, 103610, 103600, 103600, 103590, 103560, 103530, 103490, 103470, 
    103440, 103410, 103410, 103400, 103390, 103370, 103360, 103330, 103300, 
    103280, 103260, 103210, 103180, 103140, 103100, 103080, 103060, 103050, 
    103060, 103040, 102990, 102960, 102900, 102880, 102810, 102770, 102730, 
    102690, 102640, 102610, 102560, 102510, 102450, 102390, 102320, 102240, 
    102160, 102080, 101990, 101940, 101870, 101820, 101790, 101730, 101650, 
    101590, 101510, 101430, 101380, 101310, 101260, 101200, 101140, 101150, 
    101140, 101140, 101130, 101110, 101100, 101130, 101110, 101120, 101120, 
    101120, 101150, 101210, 101270, 101310, 101360, 101390, 101430, 101470, 
    101480, 101500, 101510, 101560, 101610, 101650, 101710, 101740, 101780, 
    101790, 101850, 101860, 101860, 101840, 101870, 101840, 101870, 101880, 
    101900, 101940, 101950, 101970, 101990, 101990, 102020, 102000, 102040, 
    102050, 102060, 102060, 102090, 102120, 102150, 102160, 102180, 102190, 
    102200, 102200, 102210, 102210, 102220, 102260, 102300, 102300, 102290, 
    102280, 102260, 102280, 102280, 102270, 102280, 102310, 102320, 102350, 
    102350, 102350, 102330, 102310, 102280, 102240, 102220, 102200, 102180, 
    102170, 102170, 102190, 102210, 102210, 102190, 102160, 102060, 102060, 
    102000, 101960, 101950, 101930, 101900, 101870, 101830, 101820, 101780, 
    101730, 101660, 101600, 101540, 101480, 101420, 101360, 101300, 101240, 
    101190, 101140, 101080, 101020, 100960, 100900, 100820, 100740, 100670, 
    100600, 100520, 100510, 100480, 100420, 100360, 100330, 100290, 100270, 
    100260, 100230, 100240, 100230, 100250, 100290, 100330, 100370, 100400, 
    100440, 100460, 100490, 100510, 100530, 100560, 100580, 100620, 100650, 
    100700, 100730, 100740, 100760, 100780, 100810, 100830, 100860, 100860, 
    100870, 100910, 100940, 100960, 101000, 101040, 101070, 101070, 101100, 
    101110, 101120, 101130, 101140, 101160, 101190, 101230, 101250, 101290, 
    101300, 101300, 101300, 101340, 101370, 101370, 101380, 101400, 101430, 
    101450, 101450, 101440, 101450, 101440, 101460, 101450, 101460, 101450, 
    101420, 101390, 101380, 101380, 101370, 101410, 101390, 101360, 101340, 
    101310, 101250, 101220, 101230, 101200, 101180, 101210, 101230, 101220, 
    101210, 101210, 101190, 101170, 101090, 101080, 101070, 101020, 100970, 
    100940, 100920, 100950, 100960, 100960, 100940, 100930, 100910, 100890, 
    100880, 100850, 100830, 100770, 100670, 100730, 100750, 100740, 100720, 
    100680, 100650, 100640, 100610, 100580, 100570, 100550, 100510, 100490, 
    100460, 100410, 100390, 100350, 100310, 100310, 100290, 100290, 100280, 
    100290, 100310, 100290, 100290, 100280, 100290, 100270, 100260, 100210, 
    100200, 100150, 100120, 100140, 100140, 100090, 99950, 99910, 99870, 
    99810, 99720, 99640, 99610, 99570, 99540, 99530, 99520, 99490, 99480, 
    99440, 99380, 99320, 99240, 99180, 99150, 99170, 99200, 99220, 99220, 
    99230, 99210, 99180, 99160, 99160, 99180, 99190, 99220, 99370, 99390, 
    99460, 99580, 99610, 99630, 99720, 99790, 99900, 99950, 100020, 100090, 
    100140, 100210, 100300, 100340, 100420, 100430, 100520, 100570, 100640, 
    100690, 100740, 100800, 100850, 100930, 101000, 101060, 101120, 101180, 
    101190, 101240, 101280, 101250, 101290, 101340, 101420, 101450, 101500, 
    101570, 101590, 101590, 101610, 101630, 101660, 101650, 101650, 101620, 
    101640, 101630, 101670, 101690, 101710, 101710, 101710, 101700, 101630, 
    101620, 101560, 101480, 101550, 101530, 101460, 101530, 101550, 101600, 
    101550, 101530, 101480, 101480, 101490, 101510, 101510, 101510, 101500, 
    101520, 101490, 101440, 101390, 101370, 101300, 101190, 101110, 101070, 
    101120, 101150, 101120, 101090, 101090, 101040, 101030, 101010, 100990, 
    100940, 100860, 100750, 100730, 100740, 100760, 100810, 100830, 100810, 
    100810, 100810, 100800, 100750, 100750, 100720, 100650, 100590, 100560, 
    100580, 100580, 100560, 100530, 100500, 100490, 100460, 100400, 100360, 
    100290, 100260, 100200, 100190, 100230, 100160, 100110, 100100, 100110, 
    100130, 100150, 100170, 100210, 100210, 100250, 100270, 100280, 100330, 
    100390, 100460, 100540, 100650, 100720, 100810, 100900, 100990, 101080, 
    101160, 101250, 101350, 101400, 101450, 101490, 101560, 101590, 101630, 
    101660, 101690, 101720, 101750, 101840, 101880, 101910, 101960, 101990, 
    102010, 102020, 102010, 102040, 102080, 102110, 102150, 102170, 102190, 
    102210, 102210, 102230, 102230, 102240, 102230, 102240, 102230, 102220, 
    102210, 102200, 102180, 102190, 102180, 102170, 102160, 102140, 102110, 
    102080, 102070, 102040, 102030, 102000, 101940, 101900, 101870, 101810, 
    101760, 101690, 101670, 101630, 101600, 101550, 101520, 101460, 101420, 
    101390, 101370, 101320, 101280, 101230, 101170, 101150, 101120, 101110, 
    101080, 101080, 101050, 101000, 100980, 100940, 100910, 100890, 100840, 
    100800, 100760, 100680, 100660, 100610, 100590, 100570, 100540, 100500, 
    100470, 100430, 100430, 100410, 100410, 100430, 100440, 100430, 100410, 
    100370, 100380, 100360, 100360, 100360, 100350, 100360, 100400, 100450, 
    100490, 100490, 100480, 100490, 100490, 100480, 100440, 100420, 100380, 
    100340, 100340, 100360, 100330, 100330, 100320, 100310, 100310, 100290, 
    100260, 100230, 100220, 100210, 100190, 100180, 100150, 100120, 100100, 
    100060, 100030, 99990, 99970, 99950, 99910, 99880, 99870, 99840, 99800, 
    99790, 99770, 99730, 99680, 99620, 99640, 99630, 99580, 99530, 99510, 
    99530, 99540, 99540, 99500, 99540, 99510, 99510, 99510, 99480, 99430, 
    99390, 99380, 99420, 99440, 99460, 99450, 99500, 99540, 99550, 99650, 
    99690, 99700, 99720, 99680, 99690, 99680, 99670, 99710, 99740, 99760, 
    99800, 99800, 99860, 99880, 99890, 99900, 99920, 99930, 99880, 99900, 
    99980, 100020, 100050, 100090, 100100, 100130, 100180, 100210, 100200, 
    100300, 100400, 100490, 100510, 100520, 100520, 100570, 100670, 100770, 
    100840, 100930, 100990, 101020, 101070, 101250, 101260, 101290, 101340, 
    101380, 101390, 101440, 101450, 101450, 101460, 101460, 101460, 101430, 
    101390, 101350, 101290, 101220, 101160, 101120, 101090, 101060, 101050, 
    101020, 101040, 101000, 100980, 100960, 100910, 100870, 100850, 100830, 
    100820, 100810, 100810, 100820, 100860, 100810, 100770, 100770, 100760, 
    100840, 100770, 100820, 100830, 100750, 100700, 100780, 100850, 100820, 
    100800, 100820, 100900, 100960, 100990, 101000, 101040, 101090, 101130, 
    101160, 101190, 101290, 101380, 101390, 101410, 101400, 101430, 101420, 
    101410, 101430, 101470, 101560, 101620, 101630, 101670, 101690, 101700, 
    101740, 101770, 101790, 101780, 101820, 101840, 101820, 101820, 101820, 
    101840, 101860, 101840, 101850, 101840, 101830, 101810, 101770, 101780, 
    101770, 101710, 101660, 101600, 101560, 101490, 101420, 101340, 101250, 
    101150, 101120, 101070, 101010, 100940, 100880, 100800, 100710, 100610, 
    100460, 100340, 100210, 100120, 100010, 99870, 99750, 99630, 99570, 
    99490, 99440, 99530, 99440, 99370, 99330, 99290, 99260, 99240, 99270, 
    99320, 99330, 99420, 99490, 99560, 99620, 99670, 99730, 99800, 99860, 
    99980, 100100, 100210, 100290, 100380, 100450, 100550, 100630, 100660, 
    100650, 100730, 100750, 100810, 100870, 100900, 100910, 100940, 100970, 
    100970, 100970, 100970, 100950, 100930, 100870, 100820, 100790, 100810, 
    100870, 100910, 100920, 101020, 101020, 101010, 101000, 100990, 100990, 
    100990, 101010, 101000, 100980, 100980, 100920, 100870, 100840, 100790, 
    100720, 100650, 100590, 100530, 100440, 100340, 100260, 100170, 100110, 
    100000, 99880, 99720, 99610, 99470, 99380, 99320, 99210, 99100, 99000, 
    98910, 98870, 98890, 98860, 98770, 98720, 98690, 98660, 98630, 98600, 
    98540, 98540, 98540, 98550, 98520, 98510, 98490, 98460, 98460, 98480, 
    98520, 98550, 98600, 98610, 98650, 98660, 98670, 98690, 98780, 98820, 
    98840, 98880, 98950, 98930, 98970, 98960, 99000, 99040, 99050, 99110, 
    99140, 99180, 99180, 99240, 99230, 99250, 99250, 99260, 99280, 99290, 
    99270, 99250, 99240, 99220, 99210, 99230, 99250, 99250, 99230, 99240, 
    99240, 99220, 99220, 99200, 99160, 99120, 99090, 99110, 99100, 99100, 
    99090, 99080, 99060, 99060, 99040, 99030, 99000, 98980, 98980, 99000, 
    99080, 99160, 99210, 99220, 99230, 99250, 99310, 99340, 99410, 99410, 
    99480, 99490, 99490, 99560, 99660, 99670, 99690, 99730, 99770, 99750, 
    99800, 99810, 99830, 99840, 99880, 99880, 99870, 99890, 99900, 99870, 
    99870, 99840, 99790, 99750, 99710, 99740, 99740, 99680, 99670, 99680, 
    99740, 99760, 99760, 99800, 99830, 99860, 99890, 99950, 100010, 100070, 
    100130, 100180, 100220, 100280, 100330, 100370, 100420, 100400, 100400, 
    100460, 100510, 100570, 100580, 100600, 100720, 100790, 100830, 100800, 
    100760, 100790, 100830, 100840, 100870, 100880, 100870, 100850, 100830, 
    100790, 100770, 100750, 100690, 100650, 100610, 100600, 100610, 100600, 
    100570, 100540, 100500, 100470, 100450, 100430, 100420, 100410, 100440, 
    100480, 100520, 100560, 100590, 100600, 100620, 100610, 100620, 100620, 
    100620, 100580, 100560, 100550, 100590, 100550, 100550, 100550, 100560, 
    100530, 100500, 100470, 100480, 100470, 100460, 100420, 100480, 100520, 
    100560, 100560, 100560, 100560, 100570, 100550, 100550, 100550, 100560, 
    100550, 100540, 100540, 100550, 100560, 100560, 100560, 100530, 100530, 
    100510, 100490, 100450, 100430, 100400, 100400, 100460, 100460, 100440, 
    100440, 100430, 100380, 100410, 100290, 100190, 100150, 100130, 99960, 
    99960, 99820, 99870, 99840, 99780, 99650, 99570, 99530, 99530, 99550, 
    99550, 99510, 99380, 99320, 99300, 99340, 99410, 99510, 99550, 99560, 
    99560, 99540, 99540, 99580, 99550, 99530, 99500, 99480, 99480, 99460, 
    99500, 99460, 99480, 99510, 99510, 99530, 99540, 99540, 99570, 99570, 
    99600, 99600, 99600, 99620, 99630, 99640, 99650, 99660, 99680, 99740, 
    99790, 99820, 99810, 99800, 99830, 99870, 99930, 99940, 99980, 100010, 
    100060, 100090, 100100, 100120, 100160, 100200, 100200, 100160, 100190, 
    100230, 100230, 100220, 100220, 100220, 100240, 100220, 100240, 100230, 
    100190, 100200, 100190, 100170, 100180, 100150, 100150, 100130, 100120, 
    100110, 100080, 100070, 100020, 99980, 99940, 99910, 99870, 99820, 99760, 
    99710, 99650, 99610, 99570, 99520, 99450, 99400, 99330, 99270, 99270, 
    99240, 99210, 99170, 99140, 99100, 99070, 99040, 98980, 98950, 98930, 
    98910, 98900, 98900, 98890, 98880, 98860, 98850, 98840, 98810, 98800, 
    98800, 98810, 98820, 98830, 98850, 98860, 98890, 98890, 98910, 98950, 
    98970, 98990, 99000, 99030, 99060, 99080, 99110, 99130, 99180, 99230, 
    99260, 99280, 99300, 99330, 99350, 99400, 99450, 99490, 99520, 99540, 
    99560, 99570, 99550, 99520, 99500, 99460, 99450, 99430, 99410, 99400, 
    99370, 99350, 99320, 99280, 99280, 99250, 99230, 99200, 99190, 99180, 
    99200, 99230, 99250, 99260, 99290, 99320, 99360, 99400, 99460, 99480, 
    99530, 99580, 99620, 99690, 99740, 99770, 99880, 99940, 100000, 100050, 
    100110, 100180, 100280, 100370, 100450, 100520, 100600, 100680, 100720, 
    100810, 100880, 100930, 101000, 101040, 101050, 101070, 101120, 101130, 
    101120, 101120, 101200, 101240, 101240, 101280, 101340, 101350, 101370, 
    101390, 101390, 101420, 101440, 101420, 101400, 101400, 101380, 101410, 
    101410, 101410, 101540, 101590, 101650, 101740, 101830, 101910, 101980, 
    102060, 102100, 102150, 102220, 102280, 102310, 102390, 102400, 102410, 
    102430, 102430, 102370, 102410, 102370, 102270, 102130, 101960, 101830, 
    101780, 101680, 101420, 101260, 101100, 100900, 100710, 100540, 100410, 
    100290, 100180, 100130, 100140, 100130, 100130, 100110, 100050, 99970, 
    99900, 99810, 99660, 99540, 99460, 99440, 99430, 99430, 99360, 99220, 
    99310, 99450, 99510, 99640, 99690, 99750, 99830, 99940, 100040, 100080, 
    100140, 100180, 100310, 100330, 100360, 100390, 100430, 100450, 100500, 
    100520, 100490, 100500, 100490, 100510, 100630, 100730, 100780, 100800, 
    100920, 101010, 100990, 100990, 100930, 100970, 101000, 100950, 100900, 
    100850, 100820, 100830, 100830, 100810, 100770, 100790, 100800, 100850, 
    100890, 100930, 100890, 100920, 100920, 100890, 100870, 100840, 100820, 
    100830, 100790, 100820, 100860, 100870, 100880, 100880, 100880, 100910, 
    100940, 100890, 100840, 100820, 100790, 100810, 100850, 100880, 100870, 
    100870, 100850, 100780, 100750, 100750, 100680, 100640, 100620, 100530, 
    100540, 100500, 100390, 100360, 100310, 100300, 100220, 100140, 100070, 
    100030, 99990, 99970, 99940, 99910, 99880, 99880, 99900, 99910, 99940, 
    99920, 99920, 99900, 99870, 99880, 99920, 99960, 99940, 99940, 99940, 
    99980, 99980, 100000, 100010, 100000, 99990, 100020, 100040, 100070, 
    100080, 100110, 100080, 100100, 100130, 100130, 100130, 100150, 100160, 
    100150, 100140, 100140, 100100, 100070, 100080, 100080, 100050, 100000, 
    100000, 99970, 99930, 99890, 99880, 99860, 99860, 99820, 99790, 99760, 
    99740, 99720, 99680, 99640, 99610, 99590, 99570, 99560, 99530, 99500, 
    99460, 99410, 99400, 99370, 99340, 99300, 99290, 99280, 99270, 99280, 
    99260, 99280, 99310, 99340, 99360, 99360, 99370, 99420, 99460, 99500, 
    99530, 99550, 99600, 99640, 99670, 99680, 99720, 99740, 99740, 99720, 
    99720, 99740, 99740, 99760, 99790, 99810, 99870, 99900, 100030, 100110, 
    100120, 100190, 100260, 100360, 100430, 100520, 100640, 100710, 100800, 
    100860, 100930, 100970, 101010, 101060, 101120, 101170, 101220, 101300, 
    101350, 101380, 101420, 101480, 101570, 101620, 101650, 101670, 101680, 
    101700, 101730, 101770, 101820, 101850, 101890, 101930, 101950, 101960, 
    102020, 102050, 102070, 102090, 102110, 102140, 102170, 102180, 102180, 
    102190, 102210, 102250, 102230, 102220, 102240, 102210, 102230, 102230, 
    102210, 102180, 102150, 102100, 102040, 102000, 101940, 101880, 101810, 
    101740, 101710, 101660, 101580, 101500, 101440, 101390, 101350, 101310, 
    101250, 101210, 101170, 101180, 101220, 101220, 101220, 101220, 101220, 
    101220, 101200, 101140, 101070, 101010, 100940, 100890, 100760, 100710, 
    100610, 100550, 100450, 100370, 100330, 100260, 100210, 100170, 100120, 
    100090, 100030, 99960, 99910, 99830, 99770, 99730, 99660, 99630, 99590, 
    99580, 99600, 99520, 99530, 99520, 99530, 99590, 99620, 99680, 99680, 
    99620, 99640, 99590, 99660, 99680, 99700, 99710, 99690, 99700, 99680, 
    99690, 99690, 99670, 99660, 99630, 99620, 99610, 99590, 99590, 99570, 
    99570, 99550, 99530, 99530, 99540, 99530, 99550, 99560, 99580, 99590, 
    99600, 99640, 99680, 99730, 99770, 99780, 99850, 99880, 99940, 99970, 
    99960, 100030, 100100, 100150, 100180, 100240, 100240, 100220, 100230, 
    100250, 100310, 100310, 100340, 100340, 100350, 100380, 100420, 100420, 
    100400, 100390, 100390, 100400, 100390, 100390, 100390, 100390, 100380, 
    100360, 100350, 100330, 100330, 100320, 100320, 100320, 100330, 100310, 
    100300, 100290, 100270, 100230, 100190, 100130, 100060, 100010, 99930, 
    99920, 99920, 99950, 99950, 99960, 100010, 100060, 100080, 100120, 
    100140, 100190, 100200, 100240, 100310, 100370, 100440, 100520, 100600, 
    100620, 100650, 100670, 100670, 100650, 100640, 100630, 100640, 100630, 
    100660, 100670, 100690, 100710, 100680, 100670, 100660, 100630, 100610, 
    100580, 100540, 100480, 100450, 100420, 100380, 100320, 100240, 100130, 
    99990, 99810, 99580, 99340, 99170, 98970, 98770, 98630, 98450, 98270, 
    98110, 97930, 97740, 97540, 97330, 97110, 96890, 96660, 96430, 96310, 
    96220, 96130, 96120, 96130, 96160, 96210, 96410, 96590, 96800, 96950, 
    97100, 97170, 97330, 97510, 97780, 97980, 98000, 98100, 98240, 98450, 
    98540, 98600, 98690, 98790, 98870, 98960, 99020, 99060, 99040, 99050, 
    99060, 99030, 99020, 98990, 98940, 98930, 98880, 98830, 98820, 98780, 
    98710, 98670, 98620, 98610, 98560, 98580, 98570, 98550, 98550, 98580, 
    98620, 98630, 98670, 98690, 98790, 98800, 98880, 99000, 99030, 99100, 
    99190, 99270, 99380, 99560, 99620, 99670, 99730, 99820, 99940, 100000, 
    100040, 100080, 100180, 100240, 100310, 100380, 100420, 100420, 100450, 
    100480, 100510, 100510, 100560, 100600, 100590, 100550, 100550, 100550, 
    100550, 100500, 100470, 100420, 100400, 100400, 100400, 100390, 100390, 
    100350, 100310, 100330, 100310, 100270, 100250, 100220, 100230, 100220, 
    100210, 100230, 100260, 100300, 100330, 100360, 100420, 100470, 100500, 
    100530, 100590, 100630, 100730, 100830, 100900, 100990, 101080, 101130, 
    101190, 101240, 101270, 101330, 101360, 101410, 101430, 101490, 101530, 
    101570, 101590, 101600, 101660, 101680, 101700, 101690, 101730, 101780, 
    101820, 101830, 101850, 101850, 101880, 101840, 101840, 101850, 101880, 
    101880, 101880, 101860, 101840, 101880, 101910, 101910, 101900, 101920, 
    101890, 101870, 101880, 101920, 101920, 101940, 101960, 101980, 102000, 
    102030, 102050, 102100, 102160, 102180, 102140, 102130, 102130, 102130, 
    102140, 102190, 102210, 102200, 102220, 102230, 102220, 102230, 102230, 
    102210, 102230, 102240, 102240, 102180, 102160, 102160, 102180, 102150, 
    102100, 102100, 102120, 102100, 102050, 102000, 101990, 102000, 101960, 
    101930, 101880, 101810, 101800, 101800, 101790, 101790, 101750, 101810, 
    101830, 101830, 101820, 101800, 101800, 101790, 101780, 101870, 101820, 
    101720, 101700, 101620, 101630, 101610, 101610, 101560, 101510, 101510, 
    101440, 101390, 101380, 101390, 101370, 101390, 101380, 101400, 101390, 
    101420, 101450, 101480, 101510, 101530, 101570, 101610, 101650, 101710, 
    101750, 101840, 101900, 102000, 102060, 102110, 102180, 102210, 102250, 
    102280, 102320, 102370, 102390, 102420, 102450, 102460, 102480, 102480, 
    102440, 102400, 102360, 102290, 102260, 102230, 102170, 102140, 102070, 
    102020, 101930, 101930, 101940, 101860, 101900, 101950, 101980, 101920, 
    101970, 102020, 102050, 102060, 102060, 102060, 102040, 102030, 102020, 
    102000, 102010, 102000, 102020, 102000, 101980, 101970, 101970, 101970, 
    101970, 101970, 101960, 101940, 101920, 101940, 101940, 101940, 101930, 
    101930, 101920, 101910, 101930, 101940, 101950, 101950, 101960, 101980, 
    101990, 101980, 102000, 102010, 102000, 101990, 101990, 101980, 101960, 
    101970, 101980, 101980, 101990, 102010, 102020, 102040, 102040, 102060, 
    102080, 102110, 102150, 102170, 102190, 102220, 102260, 102300, 102330, 
    102340, 102370, 102380, 102400, 102410, 102420, 102430, 102460, 102480, 
    102490, 102510, 102530, 102530, 102500, 102510, 102500, 102480, 102480, 
    102470, 102470, 102460, 102460, 102460, 102470, 102470, 102430, 102390, 
    102370, 102350, 102330, 102350, 102330, 102330, 102320, 102350, 102340, 
    102330, 102300, 102280, 102260, 102250, 102250, 102170, 102170, 102170, 
    102150, 102160, 102150, 102130, 102120, 102090, 102100, 102090, 102070, 
    102050, 102050, 102060, 102070, 102070, 102090, 102090, 102070, 102110, 
    102110, 102130, 102140, 102140, 102150, 102130, 102140, 102140, 102160, 
    102180, 102200, 102200, 102210, 102220, 102220, 102230, 102280, 102260, 
    102300, 102340, 102340, 102340, 102380, 102390, 102410, 102410, 102440, 
    102450, 102470, 102470, 102460, 102430, 102430, 102430, 102440, 102480, 
    102470, 102450, 102520, 102480, 102540, 102540, 102570, 102610, 102620, 
    102630, 102610, 102600, 102600, 102590, 102560, 102560, 102520, 102530, 
    102520, 102490, 102490, 102450, 102440, 102420, 102410, 102390, 102340, 
    102320, 102300, 102260, 102180, 102120, 102100, 102040, 101980, 101930, 
    101890, 101830, 101770, 101730, 101660, 101590, 101510, 101400, 101290, 
    101190, 101100, 100980, 100860, 100780, 100860, 100980, 101040, 101060, 
    101030, 101070, 101160, 101160, 101190, 101200, 101250, 101300, 101290, 
    101300, 101280, 101280, 101270, 101260, 101240, 101240, 101210, 101200, 
    101170, 101150, 101120, 101100, 101070, 101070, 101050, 101020, 101010, 
    100980, 100960, 100930, 100910, 100860, 100840, 100830, 100820, 100810, 
    100790, 100780, 100760, 100740, 100770, 100760, 100760, 100760, 100760, 
    100760, 100780, 100770, 100780, 100800, 100790, 100780, 100820, 100810, 
    100780, 100800, 100800, 100800, 100810, 100800, 100810, 100810, 100800, 
    100800, 100780, 100760, 100750, 100730, 100720, 100720, 100720, 100720, 
    100710, 100710, 100710, 100690, 100690, 100690, 100690, 100680, 100650, 
    100630, 100630, 100630, 100630, 100630, 100630, 100620, 100600, 100560, 
    100530, 100500, 100510, 100520, 100530, 100540, 100540, 100600, 100630, 
    100690, 100760, 100810, 100840, 100840, 100910, 100950, 100990, 101020, 
    101050, 101070, 101080, 101080, 101090, 101110, 101130, 101130, 101140, 
    101150, 101170, 101190, 101220, 101220, 101240, 101270, 101270, 101260, 
    101260, 101240, 101250, 101260, 101250, 101260, 101260, 101270, 101260, 
    101250, 101250, 101240, 101220, 101200, 101180, 101160, 101150, 101140, 
    101110, 101090, 101110, 101110, 101090, 101110, 101130, 101130, 101170, 
    101230, 101260, 101260, 101280, 101280, 101260, 101260, 101270, 101250, 
    101250, 101250, 101230, 101230, 101240, 101240, 101240, 101250, 101260, 
    101280, 101310, 101330, 101350, 101350, 101340, 101320, 101290, 101270, 
    101240, 101220, 101170, 101120, 101100, 101060, 101020, 101000, 100960, 
    100920, 100880, 100830, 100800, 100780, 100720, 100700, 100680, 100660, 
    100630, 100590, 100550, 100530, 100480, 100400, 100300, 100210, 100110, 
    100020, 99930, 99790, 99710, 99630, 99590, 99490, 99370, 99350, 99310, 
    99270, 99230, 99210, 99180, 99210, 99210, 99220, 99250, 99230, 99280, 
    99340, 99390, 99410, 99470, 99530, 99620, 99750, 99880, 99980, 100070, 
    100100, 100190, 100280, 100330, 100400, 100480, 100590, 100670, 100720, 
    100800, 100880, 100940, 100980, 101040, 101120, 101180, 101260, 101320, 
    101340, 101380, 101390, 101400, 101410, 101450, 101470, 101500, 101540, 
    101570, 101590, 101620, 101610, 101610, 101560, 101520, 101460, 101400, 
    101350, 101320, 101290, 101260, 101220, 101190, 101160, 101120, 101100, 
    101100, 101080, 101050, 101060, 101070, 101090, 101100, 101080, 101050, 
    101020, 100980, 100950, 100910, 100870, 100830, 100790, 100740, 100680, 
    100630, 100550, 100530, 100480, 100430, 100360, 100320, 100260, 100190, 
    100120, 100050, 100010, 100030, 100030, 100070, 100100, 100170, 100200, 
    100240, 100270, 100320, 100380, 100460, 100560, 100620, 100660, 100700, 
    100720, 100810, 100870, 100930, 100980, 101060, 101090, 101130, 101170, 
    101230, 101320, 101370, 101440, 101480, 101510, 101550, 101560, 101590, 
    101650, 101710, 101760, 101790, 101840, 101890, 101930, 101990, 102000, 
    102040, 102050, 102020, 102030, 102080, 102130, 102190, 102240, 102280, 
    102330, 102370, 102390, 102420, 102450, 102460, 102490, 102510, 102500, 
    102510, 102490, 102490, 102550, 102650, 102590, 102590, 102590, 102630, 
    102640, 102660, 102650, 102640, 102630, 102620, 102590, 102590, 102580, 
    102620, 102640, 102610, 102590, 102620, 102560, 102640, 102650, 102680, 
    102630, 102590, 102550, 102570, 102580, 102590, 102610, 102610, 102620, 
    102640, 102690, 102750, 102710, 102780, 102820, 102860, 102880, 102910, 
    102920, 102920, 102950, 102980, 103030, 103060, 103080, 103100, 103170, 
    103220, 103230, 103250, 103250, 103250, 103280, 103300, 103300, 103300, 
    103290, 103310, 103290, 103280, 103270, 103270, 103260, 103230, 103200, 
    103220, 103200, 103190, 103190, 103170, 103170, 103160, 103140, 103080, 
    103070, 103070, 103060, 103030, 103020, 102990, 102940, 102910, 102850, 
    102750, 102680, 102620, 102520, 102450, 102400, 102380, 102340, 102300, 
    102290, 102280, 102290, 102300, 102320, 102340, 102330, 102330, 102360, 
    102380, 102360, 102390, 102400, 102390, 102360, 102380, 102330, 102280, 
    102270, 102260, 102230, 102240, 102230, 102230, 102230, 102210, 102210, 
    102190, 102200, 102200, 102200, 102190, 102190, 102200, 102220, 102230, 
    102240, 102240, 102240, 102220, 102200, 102190, 102130, 102110, 102110, 
    102090, 102080, 102030, 101990, 101980, 101930, 101900, 101870, 101840, 
    101800, 101780, 101780, 101790, 101780, 101780, 101780, 101770, 101770, 
    101770, 101750, 101720, 101670, 101650, 101640, 101650, 101610, 101580, 
    101560, 101540, 101510, 101490, 101450, 101430, 101440, 101450, 101450, 
    101470, 101470, 101480, 101470, 101440, 101430, 101430, 101440, 101390, 
    101380, 101370, 101370, 101420, 101440, 101470, 101480, 101500, 101490, 
    101510, 101480, 101480, 101500, 101480, 101490, 101550, 101580, 101610, 
    101610, 101640, 101640, 101650, 101630, 101610, 101630, 101640, 101660, 
    101670, 101690, 101700, 101710, 101730, 101770, 101780, 101780, 101790, 
    101790, 101790, 101790, 101800, 101830, 101850, 101820, 101820, 101790, 
    101760, 101720, 101680, 101640, 101600, 101560, 101530, 101490, 101470, 
    101430, 101390, 101370, 101350, 101320, 101340, 101320, 101320, 101350, 
    101380, 101390, 101410, 101430, 101460, 101500, 101530, 101560, 101600, 
    101660, 101700, 101750, 101820, 101890, 101970, 102030, 102070, 102130, 
    102160, 102190, 102230, 102300, 102370, 102420, 102480, 102520, 102570, 
    102610, 102650, 102680, 102700, 102700, 102700, 102690, 102680, 102680, 
    102700, 102710, 102680, 102670, 102660, 102640, 102650, 102620, 102610, 
    102600, 102600, 102590, 102580, 102570, 102540, 102510, 102480, 102450, 
    102420, 102380, 102350, 102310, 102240, 102200, 102160, 102150, 102110, 
    102070, 102030, 101980, 101950, 101910, 101870, 101860, 101850, 101850, 
    101840, 101840, 101850, 101830, 101830, 101860, 101860, 101870, 101870, 
    101840, 101850, 101840, 101880, 101880, 101900, 101890, 101910, 101920, 
    101920, 101920, 101920, 101920, 101940, 101970, 101980, 101990, 101980, 
    101980, 102000, 101990, 101970, 101940, 101900, 101860, 101820, 101790, 
    101750, 101690, 101670, 101610, 101600, 101560, 101540, 101490, 101450, 
    101400, 101390, 101400, 101400, 101400, 101390, 101370, 101340, 101320, 
    101310, 101300, 101310, 101330, 101360, 101460, 101520, 101580, 101660, 
    101700, 101730, 101750, 101810, 101850, 101910, 101970, 102020, 102090, 
    102160, 102230, 102250, 102310, 102360, 102390, 102410, 102430, 102440, 
    102460, 102470, 102460, 102490, 102490, 102480, 102470, 102450, 102410, 
    102400, 102380, 102330, 102280, 102240, 102200, 102160, 102110, 102040, 
    102010, 101930, 101900, 101810, 101750, 101680, 101620, 101550, 101500, 
    101470, 101440, 101420, 101390, 101390, 101390, 101420, 101450, 101460, 
    101460, 101470, 101500, 101520, 101560, 101570, 101600, 101610, 101620, 
    101610, 101610, 101600, 101560, 101540, 101510, 101510, 101500, 101480, 
    101450, 101420, 101380, 101370, 101340, 101330, 101320, 101310, 101340, 
    101340, 101380, 101410, 101430, 101440, 101460, 101490, 101480, 101460, 
    101460, 101460, 101480, 101480, 101480, 101460, 101410, 101370, 101330, 
    101280, 101240, 101210, 101180, 101140, 101110, 101090, 101110, 101100, 
    101070, 101020, 100960, 100890, 100820, 100750, 100710, 100650, 100580, 
    100540, 100480, 100450, 100410, 100390, 100380, 100370, 100360, 100320, 
    100290, 100260, 100230, 100210, 100160, 100140, 100110, 100060, 100030, 
    99980, 99940, 99890, 99820, 99810, 99800, 99820, 99840, 99870, 99890, 
    99950, 100000, 100030, 100150, 100240, 100310, 100390, 100380, 100330, 
    100350, 100380, 100480, 100540, 100610, 100670, 100780, 100910, 101000, 
    101050, 101160, 101260, 101320, 101340, 101360, 101370, 101460, 101520, 
    101540, 101580, 101600, 101560, 101590, 101580, 101600, 101580, 101600, 
    101540, 101540, 101520, 101500, 101480, 101430, 101410, 101380, 101350, 
    101280, 101280, 101250, 101210, 101160, 101140, 101120, 101130, 101120, 
    101110, 101140, 101150, 101160, 101180, 101220, 101250, 101270, 101280, 
    101270, 101270, 101290, 101350, 101340, 101310, 101320, 101320, 101320, 
    101290, 101250, 101220, 101190, 101140, 101090, 101070, 101040, 101000, 
    100980, 100990, 100960, 100900, 100890, 100850, 100800, 100760, 100770, 
    100750, 100680, 100700, 100700, 100690, 100680, 100670, 100640, 100650, 
    100670, 100670, 100660, 100690, 100710, 100760, 100800, 100890, 100970, 
    101050, 101110, 101160, 101250, 101320, 101370, 101420, 101480, 101480, 
    101560, 101650, 101680, 101730, 101770, 101790, 101780, 101840, 101850, 
    101840, 101850, 101890, 101910, 101940, 101960, 101960, 101940, 101910, 
    101890, 101900, 101900, 101890, 101920, 101940, 101910, 101890, 101860, 
    101820, 101820, 101820, 101800, 101800, 101790, 101760, 101750, 101740, 
    101720, 101710, 101730, 101750, 101780, 101790, 101790, 101780, 101820, 
    101830, 101840, 101860, 101900, 101920, 101960, 102000, 102030, 102060, 
    102060, 102070, 102070, 102090, 102110, 102180, 102200, 102260, 102290, 
    102310, 102340, 102330, 102320, 102340, 102360, 102360, 102390, 102370, 
    102380, 102370, 102370, 102370, 102360, 102320, 102310, 102310, 102300, 
    102280, 102280, 102300, 102310, 102290, 102310, 102300, 102300, 102280, 
    102300, 102280, 102290, 102290, 102300, 102310, 102320, 102330, 102330, 
    102330, 102330, 102340, 102350, 102370, 102360, 102360, 102380, 102400, 
    102410, 102430, 102430, 102440, 102440, 102440, 102410, 102410, 102420, 
    102410, 102390, 102370, 102350, 102330, 102320, 102320, 102300, 102300, 
    102300, 102290, 102280, 102270, 102290, 102290, 102280, 102260, 102270, 
    102270, 102240, 102240, 102250, 102240, 102230, 102220, 102200, 102180, 
    102150, 102140, 102120, 102100, 102090, 102100, 102070, 102060, 102070, 
    102060, 102020, 102020, 102040, 102050, 102050, 102030, 102040, 102050, 
    102070, 102070, 102050, 102050, 102040, 102030, 102020, 102020, 102010, 
    101990, 101990, 102000, 102000, 101990, 101980, 102020, 102020, 102010, 
    102030, 102030, 102030, 102020, 102020, 102020, 102020, 102010, 101990, 
    101970, 101970, 101980, 101970, 101960, 101950, 101920, 101930, 101930, 
    101910, 101910, 101910, 101890, 101880, 101880, 101890, 101880, 101870, 
    101860, 101850, 101850, 101820, 101800, 101780, 101750, 101740, 101720, 
    101710, 101690, 101660, 101630, 101620, 101600, 101570, 101540, 101510, 
    101470, 101450, 101450, 101440, 101430, 101440, 101410, 101390, 101370, 
    101360, 101340, 101340, 101320, 101310, 101310, 101300, 101300, 101290, 
    101270, 101220, 101200, 101180, 101210, 101180, 101150, 101110, 101100, 
    101110, 101130, 101090, 101050, 101040, 101020, 101010, 100990, 100980, 
    101000, 101010, 101010, 101010, 100990, 100990, 101000, 101040, 101060, 
    101080, 101100, 101110, 101120, 101150, 101180, 101210, 101230, 101240, 
    101260, 101280, 101280, 101300, 101340, 101350, 101350, 101370, 101400, 
    101440, 101470, 101500, 101530, 101550, 101550, 101610, 101660, 101700, 
    101730, 101750, 101770, 101830, 101860, 101880, 101920, 101940, 101960, 
    101980, 101990, 101990, 101990, 102000, 102000, 102010, 102000, 101990, 
    102000, 101990, 101980, 101960, 101950, 101920, 101910, 101930, 101920, 
    101920, 101940, 101930, 101920, 101880, 101870, 101870, 101860, 101820, 
    101790, 101760, 101780, 101750, 101730, 101710, 101690, 101670, 101660, 
    101630, 101600, 101590, 101580, 101580, 101590, 101590, 101590, 101600, 
    101600, 101610, 101630, 101630, 101640, 101650, 101680, 101720, 101750, 
    101770, 101800, 101820, 101840, 101850, 101860, 101870, 101900, 101910, 
    101930, 101930, 101970, 102000, 102060, 102100, 102100, 102100, 102130, 
    102130, 102140, 102150, 102150, 102150, 102160, 102160, 102180, 102190, 
    102190, 102150, 102150, 102150, 102140, 102130, 102110, 102110, 102120, 
    102140, 102140, 102130, 102130, 102130, 102110, 102130, 102110, 102110, 
    102080, 102080, 102070, 102110, 102100, 102120, 102140, 102140, 102160, 
    102170, 102190, 102230, 102270, 102320, 102380, 102430, 102490, 102500, 
    102540, 102550, 102570, 102550, 102580, 102570, 102610, 102640, 102620, 
    102650, 102660, 102670, 102670, 102680, 102700, 102700, 102750, 102740, 
    102770, 102800, 102810, 102830, 102880, 102890, 102880, 102940, 102960, 
    102920, 102900, 102930, 102920, 102900, 102930, 102900, 102880, 102820, 
    102800, 102750, 102700, 102600, 102580, 102530, 102430, 102370, 102310, 
    102270, 102220, 102170, 102090, 102000, 101960, 101950, 101930, 101890, 
    101840, 101840, 101780, 101810, 101790, 101790, 101800, 101780, 101760, 
    101780, 101730, 101690, 101700, 101670, 101650, 101630, 101590, 101520, 
    101420, 101310, 101290, 101210, 101040, 100910, 100820, 100740, 100690, 
    100620, 100590, 100580, 100530, 100550, 100510, 100540, 100560, 100620, 
    100710, 100750, 100700, 100760, 100760, 100770, 100740, 100780, 100760, 
    100750, 100720, 100700, 100650, 100630, 100600, 100590, 100560, 100550, 
    100520, 100510, 100530, 100500, 100530, 100560, 100600, 100620, 100620, 
    100670, 100700, 100720, 100760, 100770, 100800, 100850, 100890, 100900, 
    100880, 100890, 100890, 100910, 100930, 100950, 100970, 101000, 101040, 
    101040, 101060, 101060, 101080, 101060, 101070, 101130, 101170, 101150, 
    101210, 101240, 101270, 101280, 101280, 101310, 101320, 101320, 101310, 
    101310, 101340, 101340, 101320, 101350, 101390, 101390, 101370, 101370, 
    101430, 101420, 101480, 101480, 101500, 101550, 101550, 101550, 101540, 
    101570, 101630, 101660, 101690, 101690, 101690, 101720, 101790, 101850, 
    101900, 101960, 102020, 102060, 102090, 102130, 102170, 102180, 102220, 
    102290, 102300, 102350, 102370, 102400, 102420, 102410, 102400, 102400, 
    102380, 102350, 102370, 102330, 102320, 102300, 102280, 102260, 102210, 
    102180, 102140, 102130, 102090, 102090, 102110, 102120, 102150, 102160, 
    102150, 102090, 102060, 102000, 101930, 101920, 101870, 101850, 101790, 
    101760, 101740, 101710, 101670, 101640, 101590, 101540, 101510, 101460, 
    101440, 101400, 101370, 101370, 101360, 101370, 101370, 101380, 101390, 
    101370, 101350, 101340, 101330, 101340, 101340, 101360, 101370, 101360, 
    101330, 101390, 101400, 101430, 101430, 101470, 101520, 101510, 101560, 
    101600, 101620, 101650, 101680, 101720, 101740, 101750, 101750, 101760, 
    101760, 101790, 101790, 101820, 101820, 101820, 101820, 101830, 101810, 
    101820, 101800, 101810, 101800, 101810, 101840, 101850, 101800, 101810, 
    101800, 101780, 101710, 101710, 101700, 101660, 101600, 101530, 101490, 
    101480, 101440, 101370, 101390, 101410, 101430, 101440, 101440, 101470, 
    101430, 101450, 101470, 101520, 101500, 101490, 101480, 101470, 101460, 
    101450, 101440, 101450, 101450, 101440, 101460, 101460, 101450, 101450, 
    101440, 101430, 101390, 101370, 101360, 101350, 101350, 101330, 101310, 
    101300, 101310, 101330, 101370, 101360, 101360, 101370, 101380, 101410, 
    101440, 101510, 101560, 101620, 101670, 101700, 101710, 101750, 101820, 
    101840, 101850, 101890, 101940, 101970, 102020, 102060, 102120, 102140, 
    102140, 102150, 102140, 102120, 102080, 102060, 102040, 102010, 101990, 
    101930, 101880, 101840, 101790, 101700, 101630, 101560, 101480, 101380, 
    101290, 101210, 101160, 101110, 101050, 100960, 100900, 100870, 100840, 
    100790, 100730, 100690, 100670, 100650, 100620, 100580, 100570, 100550, 
    100470, 100420, 100400, 100370, 100330, 100250, 100210, 100220, 100210, 
    100210, 100240, 100260, 100290, 100280, 100260, 100250, 100340, 100360, 
    100380, 100410, 100440, 100480, 100490, 100570, 100590, 100650, 100720, 
    100780, 100820, 100850, 100870, 100890, 100970, 101020, 101040, 101090, 
    101120, 101120, 101170, 101180, 101180, 101170, 101160, 101170, 101170, 
    101180, 101190, 101190, 101220, 101200, 101200, 101200, 101180, 101190, 
    101180, 101180, 101170, 101160, 101170, 101170, 101150, 101130, 101120, 
    101100, 101110, 101070, 101040, 101030, 101040, 101050, 101050, 101070, 
    101060, 101040, 101020, 101030, 101040, 101050, 101070, 101060, 101080, 
    101100, 101110, 101150, 101170, 101200, 101200, 101190, 101190, 101210, 
    101210, 101220, 101250, 101250, 101260, 101260, 101250, 101250, 101250, 
    101250, 101260, 101280, 101280, 101270, 101290, 101320, 101340, 101370, 
    101390, 101400, 101410, 101420, 101420, 101430, 101440, 101430, 101430, 
    101440, 101440, 101450, 101470, 101470, 101460, 101460, 101460, 101460, 
    101460, 101460, 101460, 101460, 101490, 101510, 101510, 101500, 101480, 
    101470, 101450, 101430, 101410, 101380, 101360, 101330, 101320, 101280, 
    101230, 101220, 101210, 101190, 101150, 101130, 101090, 101030, 100980, 
    100940, 100920, 100890, 100850, 100800, 100770, 100720, 100680, 100660, 
    100620, 100560, 100510, 100490, 100470, 100430, 100390, 100360, 100330, 
    100300, 100260, 100210, 100180, 100190, 100170, 100180, 100180, 100170, 
    100150, 100120, 100120, 100110, 100100, 100090, 100090, 100070, 100070, 
    100070, 100060, 100050, 100060, 100050, 100030, 100010, 99990, 100000, 
    100000, 100010, 100000, 100020, 100010, 100020, 100010, 100000, 100000, 
    100000, 100000, 100000, 99990, 99980, 99960, 99940, 99920, 99910, 99900, 
    99900, 99870, 99880, 99880, 99910, 99950, 99990, 100030, 100090, 100170, 
    100170, 100220, 100330, 100410, 100470, 100520, 100570, 100600, 100640, 
    100680, 100730, 100780, 100810, 100860, 100890, 100910, 100930, 100920, 
    100920, 100880, 100890, 100900, 100920, 100950, 100980, 100980, 101000, 
    101030, 101030, 101010, 101010, 101020, 101030, 101020, 101050, 101100, 
    101130, 101170, 101190, 101210, 101230, 101250, 101270, 101320, 101350, 
    101430, 101480, 101430, 101510, 101530, 101490, 101510, 101510, 101520, 
    101520, 101580, 101600, 101620, 101620, 101630, 101650, 101660, 101660, 
    101660, 101660, 101660, 101650, 101600, 101570, 101620, 101580, 101550, 
    101550, 101550, 101540, 101440, 101490, 101470, 101480, 101490, 101480, 
    101500, 101520, 101510, 101520, 101520, 101510, 101520, 101510, 101480, 
    101500, 101510, 101530, 101590, 101640, 101700, 101780, 101820, 101810, 
    101860, 101910, 101910, 101920, 101960, 102060, 102060, 102110, 102150, 
    102180, 102230, 102260, 102270, 102250, 102210, 102210, 102200, 102240, 
    102260, 102280, 102280, 102320, 102310, 102270, 102260, 102210, 102220, 
    102210, 102130, 102130, 102100, 102060, 102020, 101980, 101890, 101850, 
    101810, 101750, 101640, 101590, 101550, 101470, 101410, 101360, 101340, 
    101320, 101350, 101280, 101250, 101180, 101170, 101160, 101150, 101170, 
    101160, 101180, 101180, 101190, 101210, 101250, 101270, 101310, 101350, 
    101390, 101430, 101470, 101620, 101670, 101740, 101790, 101840, 101900, 
    101950, 101990, 102020, 102050, 102020, 102060, 102080, 102110, 102150, 
    102170, 102180, 102180, 102200, 102160, 102150, 102230, 102220, 102230, 
    102170, 102160, 102140, 102140, 102130, 102120, 102070, 102040, 102050, 
    102030, 102020, 102010, 102090, 102080, 102090, 102100, 102100, 102070, 
    101980, 101960, 101940, 101920, 101900, 101890, 101890, 101900, 101900, 
    101890, 101880, 101860, 101840, 101810, 101790, 101760, 101720, 101690, 
    101690, 101660, 101640, 101610, 101570, 101540, 101520, 101490, 101540, 
    101500, 101380, 101350, 101330, 101300, 101280, 101250, 101210, 101200, 
    101200, 101200, 101160, 101130, 101120, 101110, 101130, 101130, 101110, 
    101110, 101110, 101100, 101090, 101070, 101050, 101010, 100980, 100980, 
    100970, 100970, 100990, 100970, 100960, 100930, 100890, 100880, 100890, 
    100890, 100870, 100860, 100870, 100860, 100850, 100840, 100850, 100840, 
    100840, 100830, 100820, 100780, 100770, 100790, 100800, 100800, 100800, 
    100790, 100760, 100750, 100730, 100720, 100720, 100720, 100720, 100710, 
    100710, 100720, 100720, 100700, 100620, 100640, 100640, 100630, 100650, 
    100630, 100660, 100700, 100750, 100750, 100820, 100870, 100900, 100950, 
    100980, 101010, 101030, 101050, 101010, 101010, 101020, 100970, 101020, 
    101060, 101050, 101050, 101040, 101030, 101010, 101000, 100980, 100960, 
    100950, 101020, 101030, 101050, 101020, 101040, 101080, 101080, 101070, 
    101080, 101020, 101040, 101040, 101040, 101030, 101020, 101000, 100950, 
    100880, 100830, 100820, 100770, 100750, 100770, 100750, 100750, 100750, 
    100750, 100750, 100710, 100690, 100670, 100660, 100640, 100600, 100580, 
    100560, 100540, 100550, 100550, 100530, 100500, 100500, 100460, 100490, 
    100510, 100540, 100580, 100600, 100600, 100520, 100500, 100510, 100550, 
    100600, 100630, 100630, 100640, 100710, 100730, 100740, 100740, 100770, 
    100790, 100820, 100810, 100840, 100880, 100910, 100930, 100980, 101020, 
    101080, 101110, 101140, 101170, 101200, 101230, 101250, 101260, 101260, 
    101280, 101320, 101350, 101350, 101340, 101330, 101340, 101340, 101370, 
    101350, 101300, 101300, 101300, 101300, 101280, 101280, 101320, 101320, 
    101300, 101270, 101260, 101250, 101220, 101190, 101170, 101170, 101170, 
    101140, 101100, 101070, 101080, 101080, 101080, 101030, 101000, 100990, 
    100950, 100850, 100900, 100860, 100820, 100800, 100780, 100730, 100700, 
    100650, 100590, 100560, 100510, 100400, 100340, 100290, 100250, 100200, 
    100150, 100090, 100030, 99960, 99740, 99690, 99660, 99650, 99680, 99730, 
    99790, 99840, 99920, 99970, 100000, 100040, 100060, 100150, 100170, 
    100130, 100080, 100100, 100130, 100160, 100210, 100280, 100340, 100360, 
    100390, 100430, 100470, 100510, 100530, 100580, 100620, 100650, 100670, 
    100700, 100730, 100740, 100730, 100740, 100750, 100710, 100730, 100750, 
    100750, 100760, 100770, 100780, 100800, 100830, 100840, 100830, 100850, 
    100840, 100840, 100900, 100990, 101070, 101130, 101160, 101180, 101230, 
    101280, 101280, 101330, 101380, 101450, 101480, 101530, 101610, 101660, 
    101710, 101760, 101790, 101800, 101820, 101840, 101870, 101900, 101940, 
    101960, 101990, 102040, 102050, 102070, 102070, 102070, 102070, 102070, 
    102070, 102090, 102100, 102120, 102110, 102110, 102110, 102110, 102090, 
    102080, 102070, 102070, 102080, 102070, 102070, 102090, 102090, 102120, 
    102130, 102140, 102140, 102120, 102110, 102110, 102130, 102130, 102130, 
    102130, 102160, 102160, 102150, 102060, 102050, 102040, 101950, 101920, 
    101840, 101830, 101810, 101820, 101820, 101780, 101800, 101770, 101740, 
    101710, 101680, 101660, 101640, 101620, 101600, 101530, 101500, 101460, 
    101420, 101370, 101310, 101250, 101200, 101150, 101130, 101100, 101100, 
    101100, 101080, 101040, 101000, 100960, 100900, 100830, 100750, 100650, 
    100580, 100530, 100500, 100440, 100380, 100350, 100310, 100270, 100250, 
    100240, 100230, 100230, 100250, 100270, 100300, 100350, 100400, 100460, 
    100480, 100480, 100500, 100500, 100480, 100490, 100500, 100500, 100500, 
    100530, 100560, 100570, 100580, 100610, 100650, 100680, 100740, 100740, 
    100760, 100800, 100840, 100900, 100960, 100970, 100990, 101010, 101000, 
    101010, 100990, 100970, 100920, 100840, 100830, 100780, 100720, 100670, 
    100650, 100600, 100570, 100550, 100530, 100540, 100570, 100600, 100600, 
    100600, 100600, 100620, 100620, 100610, 100610, 100590, 100570, 100550, 
    100550, 100560, 100540, 100610, 100640, 100600, 100610, 100590, 100590, 
    100600, 100600, 100590, 100570, 100580, 100560, 100560, 100550, 100580, 
    100610, 100640, 100650, 100680, 100720, 100750, 100810, 100840, 100920, 
    101010, 101070, 101080, 101120, 101090, 101200, 101290, 101310, 101360, 
    101430, 101470, 101490, 101520, 101570, 101610, 101660, 101660, 101680, 
    101690, 101690, 101700, 101700, 101670, 101690, 101690, 101700, 101710, 
    101700, 101690, 101660, 101660, 101670, 101660, 101610, 101610, 101600, 
    101600, 101610, 101600, 101590, 101560, 101550, 101520, 101500, 101480, 
    101490, 101480, 101460, 101440, 101440, 101440, 101430, 101410, 101360, 
    101340, 101320, 101310, 101310, 101300, 101320, 101330, 101340, 101340, 
    101340, 101340, 101340, 101320, 101300, 101290, 101310, 101310, 101310, 
    101330, 101340, 101340, 101320, 101320, 101320, 101290, 101280, 101270, 
    101270, 101280, 101270, 101290, 101300, 101290, 101290, 101300, 101290, 
    101310, 101290, 101280, 101250, 101200, 101180, 101170, 101130, 101130, 
    101100, 101070, 101030, 100990, 100950, 100850, 100910, 100870, 100760, 
    100720, 100680, 100630, 100570, 100500, 100430, 100350, 100270, 100250, 
    100220, 100050, 99990, 99950, 99920, 99870, 99840, 99800, 99780, 99770, 
    99750, 99780, 99910, 99940, 100000, 100050, 99980, 100020, 100060, 
    100130, 100180, 100290, 100400, 100420, 100470, 100530, 100550, 100600, 
    100700, 100750, 100770, 100810, 100850, 100850, 100860, 100870, 100900, 
    100930, 100960, 101030, 101030, 101040, 101060, 101070, 101060, 101060, 
    101050, 101030, 101010, 100990, 100960, 100930, 100900, 100860, 100800, 
    100720, 100660, 100600, 100550, 100500, 100440, 100410, 100370, 100320, 
    100260, 100170, 100080, 99990, 99920, 99870, 99850, 99840, 99780, 99780, 
    99760, 99760, 99850, 99860, 99870, 99880, 99800, 99800, 99800, 99830, 
    99860, 99880, 99890, 99910, 99930, 99950, 99960, 99960, 99950, 99900, 
    99890, 99900, 99900, 99890, 99890, 99920, 99930, 99960, 99980, 99970, 
    99960, 99900, 99900, 99880, 99890, 99880, 99870, 99870, 99870, 99860, 
    99820, 99780, 99780, 99750, 99750, 99770, 99810, 99840, 99850, 99900, 
    100030, 100090, 100090, 100160, 100230, 100310, 100420, 100460, 100540, 
    100650, 100720, 100800, 100880, 101000, 101050, 101110, 101170, 101200, 
    101210, 101220, 101210, 101210, 101120, 101070, 101030, 100960, 100880, 
    100780, 100670, 100570, 100450, 100350, 100410, 100160, 100060, 99940, 
    99850, 99760, 99640, 99480, 99330, 99140, 98940, 98760, 98720, 98480, 
    98400, 98370, 98360, 98310, 98320, 98330, 98340, 98370, 98410, 98460, 
    98560, 98600, 98760, 98890, 98970, 99140, 99270, 99350, 99430, 99480, 
    99580, 99630, 99730, 99790, 99870, 100020, 100040, 100130, 100220, 
    100320, 100430, 100540, 100700, 100820, 100940, 101040, 101150, 101290, 
    101430, 101530, 101580, 101660, 101670, 101710, 101720, 101740, 101750, 
    101800, 101790, 101750, 101740, 101710, 101640, 101590, 101520, 101460, 
    101360, 101280, 101200, 101250, 101050, 100980, 100910, 100840, 100750, 
    100660, 100590, 100490, 100470, 100420, 100430, 100300, 100250, 100210, 
    100140, 100140, 100080, 100030, 99950, 99900, 99850, 99790, 99790, 99650, 
    99590, 99550, 99500, 99430, 99370, 99390, 99430, 99430, 99430, 99420, 
    99420, 99410, 99390, 99370, 99330, 99310, 99280, 99250, 99220, 99190, 
    99120, 99180, 99200, 99280, 99320, 99360, 99360, 99350, 99380, 99460, 
    99470, 99550, 99580, 99590, 99580, 99570, 99530, 99400, 99370, 99340, 
    99310, 99280, 99270, 99260, 99240, 99230, 99240, 99260, 99280, 99310, 
    99350, 99390, 99430, 99470, 99530, 99590, 99650, 99740, 99830, 99880, 
    99920, 99980, 100040, 100100, 100160, 100170, 100230, 100300, 100330, 
    100390, 100510, 100540, 100590, 100600, 100580, 100610, 100650, 100680, 
    100710, 100740, 100760, 100780, 100800, 100790, 100840, 100850, 100860, 
    100870, 100870, 100880, 100890, 100900, 100920, 100950, 100990, 101040, 
    101110, 101190, 101270, 101340, 101350, 101430, 101500, 101550, 101590, 
    101650, 101740, 101810, 101860, 101910, 101920, 101980, 102040, 102080, 
    102110, 102130, 102150, 102160, 102180, 102180, 102190, 102260, 102280, 
    102270, 102290, 102290, 102330, 102330, 102330, 102300, 102270, 102260, 
    102220, 102200, 102210, 102180, 102150, 102120, 102110, 102090, 102060, 
    102020, 102020, 101990, 102010, 102020, 102020, 102020, 102010, 102010, 
    102010, 102000, 102000, 101990, 101960, 101920, 101910, 101910, 101900, 
    101830, 101840, 101760, 101700, 101690, 101690, 101620, 101570, 101560, 
    101550, 101540, 101530, 101530, 101510, 101450, 101410, 101380, 101360, 
    101350, 101330, 101330, 101320, 101310, 101300, 101290, 101280, 101280, 
    101260, 101230, 101200, 101190, 101170, 101140, 101120, 101120, 101090, 
    101060, 101020, 100960, 100900, 100830, 100770, 100690, 100670, 100510, 
    100440, 100380, 100320, 100250, 100170, 100050, 99930, 99800, 99670, 
    99560, 99500, 99430, 99390, 99320, 99240, 99160, 99060, 98960, 98830, 
    98780, 98690, 98710, 98660, 98670, 98530, 98480, 98450, 98400, 98360, 
    98320, 98330, 98300, 98310, 98280, 98250, 98270, 98300, 98320, 98330, 
    98350, 98380, 98610, 98660, 98700, 98530, 98570, 98610, 98630, 98660, 
    98700, 98750, 98790, 98830, 98810, 98860, 98910, 98940, 98980, 99000, 
    99020, 99130, 99160, 99190, 99220, 99160, 99180, 99190, 99200, 99210, 
    99240, 99290, 99340, 99400, 99470, 99510, 99570, 99630, 99630, 99710, 
    99750, 99810, 99910, 99970, 100020, 100060, 100090, 100130, 100210, 
    100300, 100350, 100380, 100450, 100500, 100550, 100590, 100620, 100650, 
    100690, 100730, 100770, 100820, 100860, 100900, 100940, 101010, 101000, 
    101040, 101090, 101120, 101160, 101170, 101190, 101220, 101200, 101200, 
    101200, 101200, 101180, 101150, 101150, 101220, 101280, 101300, 101320, 
    101340, 101400, 101410, 101420, 101420, 101440, 101400, 101500, 101530, 
    101590, 101620, 101600, 101580, 101610, 101620, 101620, 101610, 101610, 
    101600, 101580, 101540, 101500, 101500, 101460, 101480, 101420, 101240, 
    101140, 101020, 100920, 100830, 100750, 100660, 100570, 100460, 100370, 
    100280, 100190, 100100, 100050, 100050, 100050, 100030, 100060, 100060, 
    100050, 100050, 100050, 100080, 100140, 100500, 100290, 100400, 100530, 
    100640, 100750, 100830, 100980, 101150, 101310, 101430, 101530, 101630, 
    101730, 101830, 101930, 102030, 102130, 102180, 102330, 102430, 102500, 
    102490, 102490, 102520, 102540, 102500, 102510, 102400, 102340, 102290, 
    102270, 102240, 102190, 102130, 102050, 101970, 101940, 101880, 101990, 
    101730, 101670, 101660, 101720, 101700, 101680, 101710, 101700, 101710, 
    101720, 101890, 101920, 101880, 101900, 101950, 102000, 102010, 102040, 
    101870, 101880, 101860, 101810, 101760, 101690, 101600, 101430, 101230, 
    101080, 100980, 100920, 100900, 100960, 101080, 101200, 101330, 101460, 
    101580, 101680, 101770, 101850, 101920, 101970, 102000, 102010, 102060, 
    102120, 102140, 102140, 102130, 102120, 102100, 102080, 102100, 102130, 
    102060, 102080, 102050, 102030, 101980, 102000, 102260, 102080, 102140, 
    102200, 102530, 102320, 102390, 102490, 102560, 102660, 102800, 102880, 
    102960, 103050, 103070, 103130, 103280, 103330, 103370, 103420, 103440, 
    103470, 103480, 103480, 103510, 103520, 103550, 103570, 103580, 103560, 
    103550, 103520, 103510, 103490, 103470, 103470, 103470, 103450, 103440, 
    103410, 103390, 103360, 103350, 103320, 103270, 103230, 103210, 103170, 
    103120, 103080, 103030, 102980, 102920, 102850, 102800, 102730, 102680, 
    102620, 102580, 102500, 102440, 102420, 102360, 102280, 102230, 102180, 
    102090, 102040, 101970, 101910, 101850, 101800, 101770, 101740, 101720, 
    101700, 101700, 101710, 101730, 101750, 101800, 101820, 101830, 101850, 
    101860, 101880, 101880, 101860, 101830, 101800, 101770, 101740, 101700, 
    101640, 101570, 101490, 101460, 101450, 101450, 101440, 101440, 101460, 
    101460, 101450, 101440, 101440, 101460, 101470, 101480, 101470, 101500, 
    101520, 101530, 101530, 101520, 101510, 101490, 101470, 101480, 101460, 
    101460, 101460, 101470, 101480, 101490, 101530, 101540, 101540, 101540, 
    101520, 101500, 101490, 101490, 101500, 101510, 101530, 101520, 101490, 
    101490, 101500, 101490, 101500, 101510, 101520, 101530, 101520, 101540, 
    101550, 101550, 101520, 101520, 101530, 101510, 101530, 101570, 101580, 
    101550, 101530, 101600, 101620, 101640, 101670, 101680, 101690, 101760, 
    101770, 101710, 101730, 101750, 101770, 101800, 101840, 101840, 101920, 
    101930, 101930, 102020, 101940, 101940, 101920, 101930, 101950, 101990, 
    102030, 102020, 102020, 102040, 102040, 102050, 102050, 102050, 102030, 
    101970, 101940, 101940, 101860, 101860, 101830, 101810, 101800, 101810, 
    101820, 101820, 101770, 101730, 101740, 101750, 101860, 101870, 101860, 
    101800, 101800, 101790, 101780, 101780, 101770, 101770, 101780, 101800, 
    101810, 101830, 101830, 101830, 101830, 101830, 101830, 101830, 101850, 
    101850, 101860, 101970, 101900, 101910, 101900, 101900, 101850, 101830, 
    101770, 101640, 101530, 101410, 101280, 101130, 100810, 100620, 100450, 
    100370, 100390, 100420, 100660, 100900, 101090, 101200, 101280, 101350, 
    101400, 101450, 101470, 101510, 101550, 101560, 101580, 101630, 101660, 
    101640, 101660, 101680, 101700, 101750, 101770, 101770, 101790, 101830, 
    101850, 101870, 101880, 101960, 101970, 101980, 101960, 101970, 101910, 
    101900, 101880, 101850, 101820, 101790, 101790, 101780, 101720, 101720, 
    101720, 101720, 101710, 101690, 101690, 101690, 101680, 101680, 101840, 
    101780, 101780, 101790, 101720, 101720, 101710, 101710, 101700, 101670, 
    101640, 101650, 101650, 101650, 101650, 101650, 101660, 101680, 101680, 
    101710, 101710, 101700, 101730, 101720, 101720, 101710, 101710, 101700, 
    101720, 101720, 101740, 101750, 101770, 101760, 101760, 101790, 101810, 
    101810, 101820, 101880, 101920, 101950, 101980, 102010, 102040, 102030, 
    102030, 102030, 102110, 102140, 102130, 102130, 102060, 102060, 102040, 
    102000, 101970, 101930, 101880, 101830, 101800, 101780, 101880, 101860, 
    101840, 101750, 101730, 101680, 101670, 101620, 101550, 101540, 101530, 
    101490, 101460, 101540, 101490, 101460, 101440, 101430, 101410, 101400, 
    101240, 101220, 101210, 101180, 101170, 101150, 101150, 101140, 101190, 
    101210, 101350, 101240, 101250, 101260, 101290, 101300, 101330, 101340, 
    101340, 101360, 101340, 101370, 101360, 101220, 101170, 101120, 101050, 
    101030, 101000, 101020, 101010, 101010, 101000, 100990, 101000, 101020, 
    101040, 101020, 101070, 101140, 101130, 101140, 101130, 101270, 101250, 
    101080, 101050, 101020, 101000, 100990, 100960, 100990, 101000, 101010, 
    101150, 101040, 101060, 101090, 101100, 101090, 101120, 101160, 101160, 
    101200, 101240, 101350, 101300, 101330, 101340, 101330, 101300, 101270, 
    101250, 101210, 101160, 101120, 101090, 101070, 101050, 101040, 100990, 
    100940, 100880, 100820, 100780, 100740, 100680, 100650, 100610, 100550, 
    100480, 100410, 100380, 100340, 100290, 100270, 100260, 100340, 100320, 
    100240, 100240, 100250, 100330, 100350, 100360, 100340, 100270, 100310, 
    100350, 100440, 100450, 100520, 100500, 100540, 100580, 100620, 100680, 
    100710, 100740, 100760, 100790, 100810, 100860, 100930, 101010, 101070, 
    101120, 101170, 101210, 101240, 101260, 101300, 101320, 101340, 101360, 
    101370, 101380, 101410, 101440, 101450, 101450, 101460, 101460, 101450, 
    101460, 101450, 101450, 101470, 101460, 101470, 101490, 101490, 101490, 
    101470, 101470, 101460, 101440, 101420, 101430, 101420, 101420, 101430, 
    101420, 101410, 101420, 101420, 101400, 101400, 101390, 101390, 101400, 
    101440, 101460, 101490, 101540, 101580, 101610, 101620, 101630, 101650, 
    101660, 101680, 101690, 101710, 101720, 101750, 101760, 101770, 101770, 
    101780, 101800, 101820, 101830, 101810, 101790, 101800, 101820, 101800, 
    101790, 101790, 101770, 101730, 101690, 101660, 101610, 101580, 101530, 
    101480, 101430, 101470, 101470, 101480, 101480, 101490, 101430, 101410, 
    101480, 101460, 101440, 101440, 101450, 101400, 101430, 101450, 101380, 
    101430, 101430, 101420, 101380, 101370, 101310, 101280, 101240, 101180, 
    101170, 101120, 101070, 101000, 100970, 100890, 100860, 100830, 100780, 
    100730, 100690, 100650, 100600, 100550, 100520, 100530, 100470, 100410, 
    100360, 100350, 100320, 100290, 100200, 100260, 100260, 100230, 100160, 
    100130, 100090, 100060, 100000, 99970, 99970, 99950, 99940, 99920, 99970, 
    100000, 99980, 100010, 99980, 100040, 100040, 100060, 100100, 100160, 
    100320, 100350, 100370, 100410, 100390, 100410, 100500, 100420, 100470, 
    100530, 100560, 100540, 100510, 100560, 100570, 100600, 100610, 100590, 
    100610, 100570, 100530, 100510, 100470, 100480, 100440, 100420, 100340, 
    100300, 100260, 100180, 100140, 100100, 100030, 100000, 99950, 99920, 
    99890, 99870, 99870, 99900, 99900, 99900, 99910, 99890, 99900, 99930, 
    99960, 100010, 100100, 100180, 100320, 100370, 100460, 100540, 100610, 
    100650, 100730, 100740, 100810, 100840, 100910, 100950, 101020, 101070, 
    101070, 101070, 101110, 101150, 101180, 101170, 101180, 101220, 101240, 
    101270, 101290, 101310, 101290, 101300, 101320, 101320, 101270, 101320, 
    101290, 101250, 101270, 101250, 101240, 101230, 101200, 101130, 101080, 
    101060, 100970, 100910, 100820, 100670, 100600, 100500, 100340, 100180, 
    99880, 99680, 99590, 99610, 99410, 99320, 99060, 98860, 98790, 98730, 
    98640, 98450, 98400, 98410, 98380, 98450, 98440, 98390, 98340, 98470, 
    98660, 98770, 98910, 98970, 99010, 99060, 99190, 99260, 99330, 99410, 
    99480, 99640, 99720, 99800, 99850, 99880, 100090, 100090, 99970, 100110, 
    100150, 100230, 100270, 100280, 100290, 100270, 100240, 100230, 100240, 
    100270, 100200, 100230, 100260, 100280, 100280, 100310, 100340, 100370, 
    100400, 100430, 100470, 100470, 100500, 100550, 100560, 100570, 100580, 
    100610, 100620, 100650, 100690, 100740, 100740, 100750, 100760, 100740, 
    100760, 100810, 100840, 100850, 100930, 101000, 101100, 101170, 101230, 
    101250, 101270, 101260, 101310, 101360, 101400, 101410, 101470, 101490, 
    101500, 101520, 101570, 101610, 101650, 101650, 101690, 101730, 101770, 
    101790, 101840, 101910, 101970, 101990, 101990, 102030, 101980, 101940, 
    102050, 102080, 102050, 102030, 102100, 102100, 102100, 102120, 102180, 
    102160, 102200, 102280, 102300, 102300, 102250, 102190, 102210, 102230, 
    102270, 102290, 102270, 102270, 102310, 102410, 102390, 102380, 102340, 
    102320, 102320, 102440, 102510, 102560, 102600, 102600, 102610, 102650, 
    102660, 102660, 102630, 102640, 102670, 102670, 102660, 102650, 102710, 
    102780, 102720, 102680, 102640, 102600, 102620, 102580, 102540, 102500, 
    102430, 102340, 102240, 102140, 102010, 101880, 101690, 101520, 101320, 
    101160, 100960, 100840, 100680, 100510, 100340, 100260, 100170, 100140, 
    100220, 100170, 100170, 100180, 100180, 100140, 100150, 100130, 100160, 
    100180, 100180, 100160, 100230, 100320, 100460, 100560, 100700, 100880, 
    101020, 101060, 101060, 101050, 101040, 100990, 101020, 101010, 100980, 
    101020, 101060, 101050, 101080, 101160, 101180, 101250, 101220, 101200, 
    101150, 101150, 101050, 100970, 100920, 100850, 100760, 100720, 100620, 
    100590, 100490, 100400, 100400, 100340, 100340, 100290, 100290, 100210, 
    100220, 100210, 100140, 100150, 100240, 100260, 100200, 100160, 100190, 
    100170, 100140, 100190, 100180, 100160, 100140, 100190, 100220, 100240, 
    100220, 100250, 100220, 100260, 100330, 100480, 100510, 100600, 100640, 
    100700, 100720, 100720, 100760, 100780, 100830, 100820, 100870, 100900, 
    100940, 100970, 101010, 101060, 101130, 101210, 101280, 101340, 101400, 
    101400, 101490, 101560, 101630, 101690, 101700, 101760, 101700, 101710, 
    101730, 101760, 101800, 101860, 101890, 101950, 102020, 102050, 102110, 
    102090, 102140, 102080, 102210, 102180, 102180, 102150, 102120, 102110, 
    102120, 102130, 102110, 102100, 102010, 101940, 101830, 101830, 101730, 
    101680, 101620, 101620, 101550, 101600, 101570, 101610, 101560, 101540, 
    101590, 101540, 101610, 101610, 101640, 101700, 101670, 101630, 101620, 
    101640, 101620, 101590, 101500, 101390, 101390, 101290, 101100, 101070, 
    101080, 101030, 100940, 100910, 100860, 100840, 100800, 100780, 100750, 
    100760, 100740, 100740, 100760, 100760, 100760, 100720, 100640, 100630, 
    100600, 100640, 100600, 100550, 100570, 100560, 100510, 100470, 100400, 
    100370, 100290, 100180, 100060, 99950, 99840, 99720, 99620, 99540, 99430, 
    99380, 99460, 99470, 99610, 99790, 99950, 100060, 100160, 100250, 100310, 
    100340, 100360, 100380, 100430, 100440, 100450, 100520, 100520, 100520, 
    100610, 100630, 100680, 100720, 100750, 100850, 100880, 100910, 100930, 
    100940, 101000, 101070, 101110, 101130, 101140, 101150, 101230, 101310, 
    101320, 101330, 101330, 101310, 101300, 101300, 101340, 101320, 101360, 
    101360, 101360, 101420, 101400, 101370, 101410, 101410, 101360, 101330, 
    101300, 101290, 101300, 101310, 101280, 101270, 101230, 101180, 101120, 
    101090, 100980, 100940, 100870, 100730, 100570, 100480, 100430, 100360, 
    100310, 100210, 100170, 100120, 100060, 99980, 99940, 99920, 99870, 
    99840, 99800, 99740, 99700, 99650, 99600, 99580, 99520, 99470, 99490, 
    99480, 99480, 99470, 99520, 99570, 99610, 99660, 99700, 99720, 99730, 
    99720, 99710, 99710, 99710, 99710, 99740, 99710, 99730, 99770, 99740, 
    99770, 99830, 99910, 100040, 100190, 100340, 100520, 100690, 100860, 
    100990, 101110, 101260, 101390, 101550, 101670, 101780, 101880, 101970, 
    102060, 102120, 102340, 102410, 102480, 102590, 102700, 102820, 102880, 
    102900, 102960, 103020, 103070, 103120, 103150, 103180, 103210, 103220, 
    103280, 103310, 103320, 103320, 103350, 103380, 103390, 103380, 103370, 
    103360, 103330, 103290, 103270, 103280, 103260, 103210, 103190, 103150, 
    103150, 103080, 103020, 102980, 102960, 102920, 102900, 102880, 102870, 
    102860, 102890, 102890, 102920, 102940, 102960, 102980, 103000, 103010, 
    103030, 103040, 103040, 103090, 103090, 103140, 103140, 103130, 103190, 
    103180, 103180, 103140, 103120, 102950, 103000, 103100, 103150, 103140, 
    103130, 103050, 102990, 102890, 102780, 102730, 102710, 102700, 102580, 
    102420, 102260, 102290, 102280, 102470, 102270, 102320, 102240, 102260, 
    102180, 102160, 102070, 101960, 101770, 101810, 101860, 101760, 101860, 
    101840, 101810, 101930, 101940, 101840, 101900, 101930, 101910, 101940, 
    102000, 102060, 102090, 102120, 102150, 102140, 102160, 102150, 102100, 
    102050, 101990, 102000, 101940, 101860, 101840, 101770, 101710, 101650, 
    101620, 101610, 101550, 101510, 101490, 101460, 101480, 101460, 101440, 
    101400, 101320, 101290, 101270, 101280, 101270, 101270, 101250, 101230, 
    101190, 101160, 101140, 101100, 101010, 100950, 100900, 100810, 100730, 
    100700, 100570, 100500, 100410, 100260, 100100, 100140, 100020, 99920, 
    99710, 99560, 99370, 99250, 99160, 99000, 98860, 98710, 98480, 98420, 
    98050, 98180, 98050, 97900, 97760, 97470, 97370, 97340, 97280, 97320, 
    97200, 97090, 97250, 97380, 97430, 97460, 97520, 97570, 97620, 97690, 
    97710, 97760, 97810, 97840, 97770, 97860, 98260, 98400, 98400, 98420, 
    98460, 98530, 98510, 98560, 98660, 98700, 98740, 98790, 98810, 98800, 
    98840, 98900, 98850, 98910, 98990, 98940, 98990, 98960, 98930, 98890, 
    98800, 98750, 98630, 98520, 98500, 98380, 98360, 98320, 98270, 98260, 
    98220, 98190, 98220, 98230, 98300, 98390, 98500, 98580, 98600, 98640, 
    98620, 98670, 98720, 98750, 98770, 98840, 98890, 98910, 98950, 98970, 
    99010, 99050, 99070, 99100, 99110, 99130, 99150, 99180, 99220, 99230, 
    99260, 99270, 99300, 99350, 99380, 99430, 99470, 99480, 99500, 99520, 
    99570, 99590, 99610, 99640, 99660, 99710, 99720, 99730, 99720, 99720, 
    99730, 99700, 99680, 99630, 99570, 99520, 99450, 99350, 99290, 99170, 
    99080, 98990, 98860, 98680, 98490, 98290, 98110, 97960, 97850, 97740, 
    97670, 97540, 97440, 97440, 97390, 97330, 97250, 97240, 97200, 97150, 
    97150, 97140, 97170, 97180, 97190, 97200, 97250, 97270, 97300, 97360, 
    97430, 97510, 97580, 97630, 97670, 97760, 97800, 97820, 97860, 97890, 
    97930, 97950, 98010, 98030, 98050, 98090, 98120, 98130, 98200, 98200, 
    98170, 98190, 98170, 98260, 98320, 98400, 98420, 98500, 98550, 98580, 
    98640, 98640, 98670, 98690, 98710, 98760, 98810, 98870, 98910, 98960, 
    98960, 99000, 99070, 99080, 99130, 99170, 99210, 99210, 99200, 99180, 
    99180, 99050, 99080, 99080, 99090, 99110, 99080, 99100, 99100, 99070, 
    99100, 99070, 99110, 99120, 99120, 99090, 99080, 99060, 99010, 98950, 
    98920, 98900, 98890, 98890, 98920, 98880, 98840, 98800, 98700, 98640, 
    98580, 98490, 98430, 98370, 98320, 98300, 98320, 98320, 98270, 98270, 
    98260, 98220, 98160, 98140, 98160, 98130, 98080, 98050, 97990, 98000, 
    98030, 98050, 98090, 98080, 98080, 98100, 98110, 98150, 98200, 98250, 
    98300, 98350, 98390, 98360, 98320, 98280, 98270, 98360, 98440, 98490, 
    98560, 98640, 98730, 98830, 98890, 98950, 98970, 99010, 99070, 99070, 
    99180, 99200, 99230, 99270, 99300, 99320, 99340, 99340, 99330, 99310, 
    99310, 99250, 99240, 99210, 99210, 99220, 99240, 99220, 99230, 99210, 
    99230, 99240, 99260, 99260, 99280, 99300, 99310, 99320, 99300, 99300, 
    99340, 99330, 99310, 99300, 99290, 99300, 99300, 99280, 99300, 99300, 
    99340, 99340, 99380, 99340, 99390, 99430, 99460, 99510, 99540, 99550, 
    99560, 99640, 99670, 99780, 99790, 99820, 99830, 99870, 99920, 99950, 
    99980, 100050, 100040, 100080, 100120, 100160, 100200, 100200, 100210, 
    100210, 100210, 100250, 100280, 100330, 100360, 100380, 100390, 100380, 
    100390, 100390, 100400, 100440, 100460, 100480, 100490, 100480, 100550, 
    100520, 100540, 100580, 100580, 100530, 100510, 100540, 100520, 100510, 
    100490, 100440, 100400, 100380, 100410, 100440, 100490, 100460, 100380, 
    100420, 100440, 100490, 100460, 100440, 100460, 100440, 100440, 100480, 
    100470, 100450, 100440, 100440, 100430, 100460, 100530, 100540, 100570, 
    100570, 100580, 100660, 100700, 100720, 100720, 100720, 100700, 100730, 
    100740, 100740, 100760, 100780, 100790, 100790, 100840, 100840, 100820, 
    100830, 100820, 100850, 100850, 100880, 100920, 100920, 100900, 100900, 
    100940, 100930, 100940, 100990, 100980, 101000, 101020, 101020, 101040, 
    101070, 101130, 101110, 101160, 101160, 101210, 101190, 101250, 101260, 
    101300, 101300, 101300, 101350, 101380, 101440, 101490, 101500, 101490, 
    101480, 101460, 101500, 101500, 101500, 101500, 101510, 101510, 101510, 
    101520, 101450, 101500, 101470, 101460, 101510, 101550, 101560, 101600, 
    101650, 101710, 101770, 101800, 101870, 101870, 101860, 101880, 101860, 
    101890, 101900, 101890, 101910, 101950, 101980, 101990, 101960, 101950, 
    101940, 101950, 101950, 101950, 101940, 101930, 101940, 101970, 101990, 
    102010, 102020, 101980, 101940, 101930, 101910, 101860, 101880, 101870, 
    101850, 101850, 101880, 101910, 101890, 101920, 101920, 101910, 101860, 
    101850, 101880, 101830, 101840, 101850, 101860, 101840, 101820, 101790, 
    101760, 101730, 101710, 101690, 101660, 101590, 101500, 101480, 101480, 
    101470, 101460, 101360, 101300, 101220, 101180, 101150, 101090, 101080, 
    101070, 101110, 101100, 100930, 101040, 100930, 100680, 100590, 100550, 
    100500, 100500, 100470, 100480, 100410, 100360, 100260, 100250, 100290, 
    100290, 100280, 100260, 100090, 100010, 99830, 99700, 99640, 99530, 
    99530, 99500, 99410, 99290, 99160, 98990, 98900, 98870, 98800, 98760, 
    98770, 98750, 98740, 98730, 98670, 98560, 98450, 98420, 98500, 98500, 
    98540, 98610, 98740, 98800, 98720, 98840, 98900, 98910, 98950, 99000, 
    99050, 99130, 99120, 99150, 99180, 99130, 99130, 99160, 99150, 99120, 
    99110, 99150, 99150, 99120, 99130, 99140, 99180, 99190, 99170, 99150, 
    99130, 99050, 98970, 98940, 98890, 98870, 98860, 98830, 98780, 98790, 
    98740, 98710, 98670, 98670, 98620, 98590, 98600, 98600, 98600, 98570, 
    98580, 98640, 98750, 98820, 98830, 98850, 98880, 98930, 98940, 98980, 
    99020, 99090, 99130, 99150, 99130, 99180, 99240, 99350, 99470, 99570, 
    99640, 99740, 99790, 99900, 100030, 100140, 100240, 100340, 100410, 
    100480, 100540, 100590, 100640, 100730, 100780, 100840, 100900, 100980, 
    101070, 101110, 101190, 101240, 101300, 101350, 101360, 101400, 101410, 
    101460, 101510, 101570, 101590, 101660, 101690, 101720, 101740, 101750, 
    101770, 101780, 101800, 101830, 101850, 101840, 101860, 101880, 101860, 
    101830, 101840, 101820, 101810, 101760, 101750, 101740, 101740, 101760, 
    101740, 101740, 101720, 101720, 101740, 101730, 101750, 101740, 101720, 
    101730, 101720, 101690, 101690, 101690, 101640, 101590, 101560, 101540, 
    101490, 101420, 101410, 101380, 101320, 101290, 101250, 101210, 101190, 
    101130, 101040, 100990, 100950, 100890, 100810, 100770, 100750, 100690, 
    100610, 100560, 100530, 100470, 100400, 100330, 100310, 100280, 100260, 
    100250, 100270, 100250, 100230, 100210, 100180, 100150, 100090, 100050, 
    100030, 99970, 99930, 99910, 99820, 99750, 99700, 99640, 99590, 99540, 
    99450, 99420, 99400, 99450, 99520, 99620, 99730, 99800, 99870, 99930, 
    99980, 100050, 100050, 100070, 100090, 100150, 100190, 100230, 100290, 
    100320, 100350, 100380, 100390, 100410, 100450, 100450, 100490, 100520, 
    100530, 100530, 100540, 100550, 100560, 100610, 100620, 100630, 100630, 
    100660, 100650, 100700, 100720, 100720, 100740, 100730, 100730, 100740, 
    100740, 100720, 100690, 100670, 100660, 100620, 100620, 100610, 100620, 
    100610, 100610, 100590, 100580, 100590, 100630, 100660, 100680, 100690, 
    100730, 100790, 100850, 100910, 100980, 101030, 101060, 101060, 101150, 
    101150, 101150, 101160, 101130, 101180, 101220, 101250, 101260, 101310, 
    101270, 101280, 101270, 101260, 101260, 101260, 101260, 101240, 101240, 
    101220, 101200, 101190, 101160, 101120, 101080, 101050, 101010, 100960, 
    100930, 100900, 100910, 100890, 100830, 100800, 100740, 100660, 100590, 
    100540, 100540, 100500, 100510, 100500, 100520, 100540, 100580, 100520, 
    100600, 100550, 100580, 100620, 100620, 100620, 100660, 100710, 100740, 
    100850, 100780, 100860, 100880, 100860, 100850, 100850, 100890, 100910, 
    100900, 100930, 100980, 101000, 100970, 100990, 100970, 101000, 101000, 
    100920, 100890, 100940, 100980, 101000, 101020, 101000, 101010, 101030, 
    101020, 101010, 101000, 100990, 101020, 101010, 101010, 101020, 101020, 
    101010, 101000, 100980, 100970, 100970, 100940, 100930, 100940, 100910, 
    100910, 100940, 100940, 100990, 101000, 101030, 101060, 101080, 101070, 
    101080, 101080, 101080, 101110, 101130, 101160, 101160, 101200, 101230, 
    101250, 101250, 101270, 101270, 101290, 101310, 101310, 101340, 101380, 
    101380, 101390, 101370, 101370, 101370, 101390, 101420, 101380, 101400, 
    101390, 101370, 101380, 101450, 101440, 101410, 101410, 101450, 101420, 
    101390, 101360, 101340, 101370, 101390, 101430, 101420, 101460, 101470, 
    101460, 101500, 101520, 101530, 101550, 101560, 101560, 101560, 101590, 
    101600, 101600, 101560, 101530, 101480, 101440, 101400, 101290, 101290, 
    101240, 101180, 101150, 101120, 101080, 101040, 100970, 100910, 100880, 
    100840, 100820, 100780, 100760, 100780, 100810, 100910, 101020, 101080, 
    101160, 101250, 101230, 101340, 101360, 101270, 101330, 101250, 101140, 
    101150, 101030, 100950, 100830, 100670, 100530, 100420, 100350, 100260, 
    100110, 100070, 100060, 100070, 100060, 100010, 100120, 100060, 100110, 
    100210, 100220, 100250, 100320, 100460, 100520, 100600, 100750, 100850, 
    100920, 101050, 101150, 101270, 101410, 101460, 101560, 101770, 101920, 
    101990, 102050, 102120, 102200, 102260, 102340, 102300, 102360, 102370, 
    102360, 102400, 102370, 102400, 102350, 102320, 102220, 102150, 102090, 
    102050, 101950, 101890, 101820, 101720, 101600, 101540, 101410, 101290, 
    101130, 100930, 100760, 100520, 100420, 100290, 100230, 100190, 100150, 
    100120, 100050, 100020, 100020, 99970, 100000, 100020, 100030, 100000, 
    100020, 100010, 100030, 100030, 100030, 100010, 99950, 99950, 99920, 
    99910, 99910, 99920, 99930, 99960, 100000, 100070, 100110, 100140, 
    100180, 100210, 100240, 100260, 100250, 100270, 100310, 100320, 100380, 
    100400, 100460, 100470, 100510, 100520, 100540, 100550, 100570, 100590, 
    100600, 100630, 100660, 100700, 100750, 100790, 100820, 100840, 100880, 
    100930, 101000, 101010, 101050, 101080, 101130, 101160, 101210, 101260, 
    101300, 101320, 101360, 101390, 101410, 101450, 101480, 101510, 101550, 
    101600, 101630, 101640, 101650, 101680, 101690, 101590, 101670, 101700, 
    101660, 101610, 101640, 101610, 101620, 101640, 101640, 101620, 101630, 
    101600, 101630, 101590, 101620, 101640, 101680, 101650, 101700, 101730, 
    101710, 101680, 101670, 101720, 101860, 101880, 101880, 101880, 101910, 
    101930, 101940, 101910, 101870, 101870, 101890, 101900, 101890, 101840, 
    101830, 101800, 101750, 101750, 101760, 101720, 101660, 101650, 101650, 
    101690, 101690, 101690, 101660, 101690, 101690, 101680, 101740, 101720, 
    101740, 101750, 101780, 101750, 101730, 101740, 101730, 101680, 101690, 
    101680, 101640, 101540, 101550, 101530, 101460, 101430, 101400, 101370, 
    101370, 101410, 101450, 101480, 101500, 101520, 101550, 101590, 101620, 
    101630, 101690, 101730, 101720, 101750, 101800, 101850, 101900, 101950, 
    101980, 101970, 101980, 102000, 102050, 102060, 102070, 102070, 102100, 
    102120, 102150, 102160, 102140, 102150, 102160, 102190, 102200, 102180, 
    102200, 102210, 102230, 102260, 102270, 102280, 102250, 102240, 102240, 
    102210, 102210, 102230, 102210, 102210, 102220, 102240, 102260, 102280, 
    102290, 102270, 102270, 102310, 102320, 102320, 102330, 102360, 102380, 
    102430, 102470, 102510, 102530, 102550, 102560, 102580, 102600, 102650, 
    102690, 102700, 102730, 102780, 102810, 102820, 102830, 102800, 102810, 
    102820, 102830, 102850, 102810, 102820, 102840, 102900, 102910, 102900, 
    102940, 102900, 102920, 102920, 102920, 102910, 102900, 102940, 102920, 
    102870, 102920, 102920, 102960, 102860, 102840, 102900, 102840, 102850, 
    102830, 102800, 102860, 102990, 103000, 103010, 103010, 102980, 102970, 
    103010, 103020, 103030, 103020, 102920, 102920, 102950, 102940, 102910, 
    102870, 102820, 102800, 102760, 102730, 102710, 102700, 102680, 102660, 
    102620, 102560, 102490, 102490, 102320, 102180, 102050, 101990, 101890, 
    101770, 101670, 101630, 101600, 101570, 101490, 101390, 101320, 101270, 
    101260, 101250, 101220, 101180, 101170, 101170, 101140, 101110, 101040, 
    100970, 100810, 100670, 100520, 100310, 100120, 99930, 99770, 99650, 
    99530, 99410, 99290, 99200, 99090, 98970, 98840, 98690, 98540, 98380, 
    98270, 98090, 97950, 97860, 97780, 97690, 97620, 97550, 97460, 97390, 
    97450, 97460, 97530, 97620, 97710, 97790, 97840, 97870, 97910, 98040, 
    98090, 98120, 98120, 98100, 98110, 98130, 98160, 98180, 98180, 98200, 
    98210, 98190, 98170, 98150, 98130, 98090, 98020, 97960, 97940, 97910, 
    97850, 97760, 97710, 97670, 97610, 97550, 97480, 97450, 97410, 97390, 
    97400, 97410, 97400, 97410, 97420, 97460, 97500, 97520, 97600, 97690, 
    97800, 97920, 97960, 98060, 98140, 98170, 98200, 98240, 98280, 98350, 
    98380, 98400, 98420, 98430, 98440, 98430, 98420, 98410, 98400, 98410, 
    98400, 98430, 98430, 98440, 98450, 98460, 98490, 98470, 98500, 98480, 
    98450, 98440, 98420, 98400, 98380, 98350, 98330, 98320, 98310, 98300, 
    98250, 98200, 98170, 98110, 98090, 98050, 97960, 97930, 97900, 97870, 
    97830, 97830, 97820, 97820, 97810, 97820, 97810, 97810, 97830, 97870, 
    97920, 97980, 98030, 98060, 98090, 98110, 98160, 98190, 98220, 98260, 
    98260, 98280, 98330, 98380, 98430, 98480, 98510, 98540, 98560, 98590, 
    98640, 98640, 98680, 98720, 98760, 98800, 98830, 98870, 98880, 98880, 
    98900, 98920, 98920, 98910, 98920, 98870, 98880, 98880, 98900, 98900, 
    98910, 98860, 98830, 98800, 98810, 98810, 98820, 98780, 98810, 98810, 
    98800, 98830, 98810, 98770, 98770, 98750, 98750, 98830, 98830, 98840, 
    98840, 98850, 98870, 98870, 98850, 98880, 98870, 98860, 98890, 98910, 
    98950, 98980, 99030, 99050, 99080, 99140, 99190, 99230, 99300, 99350, 
    99420, 99490, 99530, 99550, 99600, 99680, 99710, 99770, 99840, 99880, 
    99930, 99990, 100040, 100080, 100120, 100160, 100220, 100300, 100330, 
    100410, 100460, 100490, 100500, 100580, 100630, 100670, 100720, 100760, 
    100810, 100840, 100880, 100950, 101010, 101110, 101200, 101330, 101430, 
    101510, 101620, 101620, 101710, 101820, 101860, 101830, 101800, 101730, 
    101630, 101480, 101430, 101160, 100990, 100740, 100450, 100210, 99910, 
    99690, 99480, 99150, 99000, 98710, 98640, 98470, 98410, 98330, 98300, 
    98310, 98300, 98310, 98340, 98340, 98290, 98250, 98190, 98170, 98120, 
    98090, 98130, 98150, 98220, 98260, 98240, 98240, 98230, 98250, 98290, 
    98320, 98340, 98420, 98510, 98560, 98610, 98580, 98580, 98600, 98550, 
    98480, 98370, 98300, 98240, 98260, 98180, 98140, 98070, 98020, 98010, 
    97960, 97870, 97880, 97940, 98010, 98070, 98080, 98180, 98330, 98410, 
    98540, 98560, 98580, 98600, 98640, 98660, 98670, 98690, 98750, 98750, 
    98790, 98810, 98840, 98880, 98900, 98910, 98910, 98890, 98890, 98880, 
    98880, 98890, 98870, 98890, 98910, 98890, 98890, 98890, 98890, 98890, 
    98850, 98830, 98780, 98810, 98820, 98820, 98790, 98800, 98770, 98770, 
    98770, 98790, 98780, 98780, 98760, 98750, 98750, 98770, 98780, 98780, 
    98780, 98780, 98780, 98750, 98760, 98760, 98760, 98750, 98740, 98740, 
    98720, 98690, 98720, 98680, 98670, 98650, 98620, 98630, 98660, 98670, 
    98710, 98740, 98750, 98760, 98760, 98760, 98770, 98770, 98770, 98760, 
    98760, 98780, 98780, 98800, 98810, 98800, 98800, 98780, 98790, 98770, 
    98710, 98670, 98620, 98550, 98520, 98440, 98360, 98290, 98140, 98090, 
    98080, 98090, 98130, 98220, 98320, 98430, 98540, 98660, 98780, 98870, 
    98960, 99040, 99130, 99220, 99300, 99360, 99450, 99530, 99630, 99710, 
    99800, 99890, 99960, 100020, 100090, 100150, 100200, 100260, 100320, 
    100370, 100430, 100490, 100540, 100580, 100610, 100620, 100670, 100670, 
    100720, 100750, 100710, 100800, 100830, 100850, 100850, 100950, 100940, 
    100960, 100960, 100960, 101010, 101030, 101000, 100970, 100920, 100860, 
    100760, 100690, 100490, 100490, 100470, 100480, 100460, 100400, 100360, 
    100310, 100270, 100260, 100230, 100180, 100190, 100070, 100030, 99990, 
    99970, 99930, 99870, 99800, 99760, 99730, 99710, 99690, 99700, 99730, 
    99770, 99820, 99830, 99810, 99840, 99870, 99890, 99920, 99950, 100020, 
    100080, 100160, 100190, 100260, 100330, 100400, 100450, 100530, 100570, 
    100640, 100750, 100840, 100950, 100950, 100980, 101010, 101040, 101050, 
    101070, 101170, 101200, 101240, 101310, 101320, 101280, 101340, 101350, 
    101400, 101320, 101330, 101330, 101360, 101320, 101290, 101250, 101250, 
    101220, 101190, 101160, 101100, 101070, 100990, 100980, 100960, 100950, 
    100940, 100880, 100870, 100850, 100870, 100800, 100770, 100790, 100760, 
    100740, 100720, 100690, 100680, 100720, 100700, 100670, 100660, 100660, 
    100620, 100550, 100580, 100620, 100550, 100550, 100530, 100470, 100480, 
    100460, 100500, 100570, 100570, 100540, 100500, 100510, 100520, 100570, 
    100570, 100580, 100600, 100590, 100590, 100590, 100620, 100600, 100640, 
    100680, 100680, 100700, 100700, 100730, 100730, 100760, 100660, 100620, 
    100580, 100480, 100530, 100310, 100430, 100400, 100340, 100350, 100390, 
    100160, 100200, 100130, 100190, 100230, 100170, 100120, 100070, 100010, 
    100010, 100050, 100030, 100020, 99960, 100010, 99980, 99980, 99950, 
    99970, 100030, 100060, 100080, 100110, 100150, 100210, 100290, 100320, 
    100320, 100320, 100340, 100420, 100460, 100490, 100500, 100530, 100540, 
    100530, 100530, 100520, 100510, 100470, 100420, 100440, 100400, 100350, 
    100320, 100290, 100260, 100240, 100230, 100220, 100200, 100160, 100120, 
    100200, 100150, 100100, 100050, 100010, 99950, 99860, 99800, 99740, 
    99690, 99650, 99650, 99680, 99700, 99720, 99750, 99780, 99800, 99820, 
    99830, 99850, 99860, 99850, 99850, 99800, 99790, 99750, 99720, 99690, 
    99630, 99570, 99530, 99460, 99390, 99320, 99270, 99230, 99140, 99060, 
    98990, 98880, 98780, 98690, 98600, 98510, 98430, 98380, 98360, 98340, 
    98330, 98330, 98310, 98320, 98280, 98260, 98230, 98170, 98100, 97990, 
    97900, 98010, 97920, 97810, 97720, 97590, 97470, 97330, 97190, 97020, 
    96850, 96680, 96540, 96430, 96290, 96210, 96210, 96230, 96260, 96260, 
    96270, 96260, 96240, 96230, 96200, 96370, 96340, 96290, 96260, 96220, 
    96170, 96130, 96100, 96080, 96050, 96010, 95960, 95990, 95950, 95920, 
    95910, 95930, 95940, 95950, 95980, 96010, 96040, 96090, 96160, 96250, 
    96320, 96380, 96440, 96490, 96560, 96650, 96720, 96760, 96810, 96860, 
    96920, 97030, 97090, 97160, 97290, 97360, 97390, 97450, 97520, 97590, 
    97630, 97680, 97680, 97720, 97770, 97840, 97910, 97970, 98040, 98120, 
    98200, 98270, 98340, 98410, 98480, 98580, 98670, 98790, 98910, 99010, 
    99090, 99200, 99300, 99340, 99400, 99470, 99500, 99540, 99590, 99670, 
    99750, 99780, 99830, 99880, 99920, 99970, 99990, 100000, 100090, 100110, 
    100090, 100150, 100150, 100160, 100130, 100070, 99980, 99930, 99880, 
    99780, 99760, 99690, 99620, 99570, 99550, 99540, 99570, 99650, 99750, 
    99870, 100000, 100140, 100230, 100380, 100470, 100570, 100700, 100740, 
    100770, 100750, 100700, 100670, 100620, 100550, 100530, 100510, 100420, 
    100350, 100310, 100280, 100260, 100310, 100380, 100450, 100540, 100660, 
    100790, 100930, 101040, 101150, 101300, 101440, 101600, 101680, 101700, 
    101780, 101820, 101880, 101870, 101840, 101750, 101630, 101490, 101320, 
    101100, 100840, 100490, 100230, 99930, 99690, 99500, 99250, 99060, 99120, 
    99110, 99090, 98990, 98970, 98870, 98700, 98480, 98220, 97910, 97540, 
    97320, 97210, 97270, 97520, 97700, 97880, 98030, 98200, 98340, 98550, 
    98630, 98720, 98900, 99110, 99350, 99580, 99780, 99960, 100150, 100370, 
    100520, 100640, 100610, 100700, 100780, 100870, 100960, 101000, 101030, 
    101050, 101040, 101050, 101030, 101010, 101010, 101060, 101080, 101100, 
    101160, 101240, 101290, 101350, 101430, 101440, 101480, 101530, 101560, 
    101610, 101650, 101720, 101750, 101790, 101830, 101850, 101870, 101890, 
    101940, 101950, 101980, 102020, 102050, 102090, 102110, 102120, 102100, 
    102080, 102070, 102110, 102050, 102060, 102070, 102070, 102090, 102070, 
    102030, 102040, 102020, 102050, 102010, 101970, 101950, 101960, 101960, 
    102010, 102010, 102070, 102070, 102030, 102070, 102060, 102090, 102060, 
    102060, 102060, 102080, 102090, 102150, 102150, 102100, 102080, 102060, 
    102090, 102080, 102080, 102090, 102070, 102010, 102010, 102050, 102080, 
    102100, 102090, 102090, 102080, 102060, 102000, 101990, 102000, 102000, 
    102000, 102010, 102010, 102010, 102010, 101990, 101990, 101980, 102010, 
    102020, 101990, 101960, 101940, 101910, 101900, 101920, 101920, 101910, 
    101850, 101780, 101770, 101740, 101680, 101680, 101640, 101600, 101540, 
    101540, 101500, 101450, 101410, 101450, 101370, 101410, 101390, 101320, 
    101330, 101360, 101390, 101390, 101400, 101440, 101410, 101400, 101460, 
    101420, 101440, 101540, 101410, 101410, 101500, 101520, 101540, 101550, 
    101450, 101410, 101420, 101430, 101530, 101460, 101440, 101490, 101460, 
    101520, 101510, 101510, 101530, 101520, 101490, 101560, 101570, 101540, 
    101550, 101570, 101590, 101600, 101590, 101590, 101540, 101500, 101540, 
    101500, 101500, 101470, 101430, 101430, 101460, 101480, 101530, 101520, 
    101490, 101450, 101510, 101560, 101560, 101550, 101550, 101560, 101560, 
    101560, 101540, 101540, 101530, 101540, 101520, 101530, 101550, 101580, 
    101570, 101580, 101550, 101480, 101440, 101430, 101400, 101340, 101280, 
    101210, 101140, 101100, 101070, 101000, 100870, 100820, 100780, 100650, 
    100530, 100470, 100410, 100310, 100240, 100220, 100170, 100090, 100010, 
    99890, 99850, 99840, 99800, 99790, 99730, 99740, 99760, 99790, 99830, 
    99880, 99890, 99930, 99940, 99950, 99900, 99950, 99950, 99940, 99920, 
    99920, 99890, 99850, 99910, 99850, 99780, 99600, 99540, 99480, 99420, 
    99370, 99310, 99260, 99230, 99220, 99210, 99180, 99150, 99140, 99120, 
    99090, 99060, 99060, 99100, 99110, 99090, 99080, 99070, 99100, 99100, 
    99070, 99060, 99060, 99070, 99120, 99160, 99210, 99280, 99360, 99490, 
    99680, 99730, 99770, 99850, 99890, 100000, 100090, 100150, 100180, 
    100280, 100410, 100480, 100540, 100590, 100630, 100680, 100720, 100800, 
    100830, 100850, 100890, 100940, 100960, 100980, 101000, 101000, 100980, 
    100940, 100930, 100930, 100960, 100920, 100870, 100860, 100610, 100460, 
    100470, 100510, 100300, 100270, 100120, 100050, 100560, 100030, 99890, 
    99930, 99880, 99720, 100330, 100300, 99690, 99690, 99670, 99720, 99750, 
    99790, 99800, 99810, 100300, 99910, 100010, 100030, 100070, 100340, 
    100140, 100210, 100230, 100280, 100320, 100380, 100380, 100360, 100340, 
    100390, 100410, 100410, 100420, 100440, 100400, 100300, 100290, 100330, 
    100340, 100300, 100280, 100190, 100190, 100180, 100120, 100040, 99970, 
    99890, 99870, 99810, 99770, 99760, 99770, 99730, 99760, 99750, 99760, 
    99770, 99790, 99860, 99910, 99970, 100040, 100100, 100150, 100230, 
    100290, 100390, 100490, 100590, 100650, 100780, 100890, 100970, 101090, 
    101220, 101240, 101310, 101390, 101520, 101600, 101690, 101740, 101820, 
    101880, 101940, 101810, 101920, 101950, 101990, 102040, 102060, 102100, 
    102090, 102090, 102160, 102250, 102260, 102330, 102360, 102380, 102420, 
    102450, 102480, 102510, 102540, 102550, 102570, 102610, 102670, 102700, 
    102720, 102760, 102790, 102820, 102830, 102850, 102890, 102920, 102950, 
    102980, 103000, 103000, 103020, 103030, 103030, 103050, 103030, 103040, 
    103060, 103040, 103030, 103010, 103000, 102990, 102960, 102950, 102920, 
    102910, 102930, 102880, 102780, 102720, 102720, 102650, 102510, 102420, 
    102230, 102240, 102140, 101980, 101880, 101800, 101770, 101710, 101600, 
    101550, 101410, 101290, 101140, 101020, 100940, 100800, 100710, 100620, 
    100540, 100450, 100380, 100300, 100230, 100130, 100080, 100000, 99900, 
    99880, 99950, 99840, 99800, 99740, 99610, 99570, 99550, 99480, 99300, 
    99240, 99130, 99080, 99050, 98960, 98880, 98800, 98780, 98730, 98710, 
    98730, 98740, 98760, 98750, 98750, 98760, 98810, 98850, 98880, 98920, 
    98940, 99010, 99080, 99140, 99190, 99250, 99320, 99360, 99430, 99480, 
    99520, 99550, 99600, 99640, 99680, 99720, 99760, 99790, 99790, 99810, 
    99840, 99850, 99880, 99860, 99830, 99830, 99840, 99850, 99830, 99830, 
    99810, 99750, 99680, 99620, 99590, 99550, 99580, 99560, 99540, 99480, 
    99450, 99450, 99490, 99450, 99450, 99460, 99470, 99460, 99430, 99470, 
    99500, 99550, 99580, 99590, 99590, 99590, 99610, 99610, 99610, 99630, 
    99640, 99650, 99640, 99690, 99720, 99720, 99730, 99750, 99750, 99760, 
    99800, 99870, 99890, 99940, 99990, 100020, 100030, 100060, 100110, 
    100130, 100120, 100140, 100160, 100170, 100190, 100220, 100240, 100260, 
    100270, 100290, 100290, 100300, 100320, 100340, 100380, 100420, 100470, 
    100470, 100500, 100540, 100550, 100540, 100540, 100550, 100560, 100570, 
    100600, 100610, 100620, 100610, 100590, 100620, 100620, 100600, 100560, 
    100580, 100600, 100590, 100600, 100600, 100590, 100590, 100590, 100550, 
    100530, 100470, 100430, 100410, 100380, 100360, 100330, 100270, 100230, 
    100210, 100170, 100140, 100110, 100020, 100000, 99980, 99990, 99990, 
    100040, 100070, 100080, 100110, 100160, 100190, 100220, 100260, 100300, 
    100360, 100410, 100450, 100510, 100570, 100600, 100640, 100670, 100720, 
    100760, 100770, 100780, 100790, 100810, 100910, 100930, 100940, 100960, 
    100940, 100820, 100800, 100760, 100760, 100730, 100680, 100620, 100570, 
    100520, 100440, 100360, 100280, 100230, 100120, 100040, 99940, 99810, 
    99750, 99740, 99720, 99730, 99780, 99920, 100080, 100230, 100310, 100430, 
    100520, 100620, 100650, 100730, 100810, 100890, 100910, 101010, 101040, 
    101000, 100970, 100920, 100800, 100720, 100620, 100520, 100460, 100320, 
    100200, 100070, 99980, 99850, 99760, 99650, 99560, 99470, 99400, 99370, 
    99320, 99290, 99260, 99280, 99290, 99310, 99340, 99370, 99430, 99510, 
    99610, 99680, 99830, 99920, 100000, 100090, 100090, 100180, 100260, 
    100330, 100390, 100480, 100540, 100570, 100630, 100650, 100680, 100720, 
    100750, 100730, 100720, 100700, 100720, 100720, 100730, 100750, 100750, 
    100760, 100790, 100820, 100850, 100880, 100910, 100940, 100960, 100990, 
    101040, 101130, 101180, 101230, 101240, 101270, 101310, 101340, 101350, 
    101360, 101370, 101390, 101410, 101450, 101450, 101470, 101410, 101390, 
    101370, 101330, 101270, 101260, 101220, 101180, 100990, 100980, 100970, 
    100960, 100920, 100890, 100860, 100840, 100820, 100780, 100760, 100720, 
    100700, 100640, 100650, 100650, 100650, 100610, 100500, 100490, 100560, 
    100520, 100490, 100430, 100280, 100270, 100100, 100190, 100310, 100410, 
    100660, 100850, 100930, 101240, 101230, 101680, 101770, 101870, 102000, 
    102030, 102080, 102040, 102220, 102250, 102270, 102250, 102250, 102290, 
    102320, 102240, 102310, 102370, 102350, 102390, 102380, 102340, 102390, 
    102410, 102360, 102160, 101960, 102180, 101990, 101900, 101790, 101690, 
    101610, 101500, 101450, 101420, 101390, 101320, 101290, 101300, 101290, 
    101290, 101230, 101310, 101330, 101460, 101430, 101450, 101470, 101470, 
    101480, 101580, 101580, 101580, 101590, 101530, 101550, 101650, 101580, 
    101610, 101600, 101610, 101620, 101560, 101600, 101600, 101590, 101570, 
    101610, 101600, 101620, 101590, 101600, 101610, 101570, 101450, 101530, 
    101500, 101500, 101510, 101480, 101500, 101500, 101530, 101590, 101600, 
    101640, 101640, 101660, 101690, 101710, 101740, 101750, 101800, 101820, 
    101850, 101870, 101880, 101910, 101930, 101930, 101940, 101920, 101910, 
    101910, 101930, 101940, 101940, 101950, 101950, 101950, 101940, 101950, 
    101940, 101950, 101950, 101950, 101930, 101920, 101900, 101910, 101950, 
    102000, 102020, 102020, 102010, 102010, 102020, 102050, 102060, 102080, 
    102110, 102130, 102150, 102160, 102140, 102140, 102140, 102140, 102120, 
    102090, 102110, 102110, 102090, 102090, 102070, 102070, 102080, 102060, 
    102050, 102000, 101990, 101980, 101970, 101970, 101950, 101960, 101960, 
    101940, 101930, 101920, 101890, 101870, 101850, 101830, 101830, 101450, 
    101430, 101410, 101400, 101380, 101380, 101380, 101370, 101360, 101370, 
    101380, 101370, 101380, 101370, 101400, 101400, 101410, 101420, 101450, 
    101510, 101570, 101600, 101620, 101670, 101700, 101730, 101790, 101820, 
    101870, 101890, 101900, 101920, 101960, 102000, 102020, 102060, 102070, 
    102080, 102110, 102100, 102110, 102120, 102130, 102110, 102110, 102110, 
    102100, 102060, 102080, 102100, 102110, 102110, 102120, 102120, 102090, 
    102090, 102100, 102120, 102110, 102110, 102080, 102080, 102030, 102010, 
    102000, 102000, 102000, 101970, 101930, 101850, 101730, 101680, 101650, 
    101570, 101540, 101560, 101550, 101500, 101460, 101420, 101400, 101410, 
    101380, 101380, 101380, 101400, 101440, 101480, 101520, 101560, 101610, 
    101640, 101680, 101700, 101700, 101710, 101780, 101800, 101870, 101880, 
    101880, 101900, 101950, 101970, 101990, 101990, 101990, 102000, 102020, 
    102020, 102040, 102100, 102180, 102210, 102200, 102210, 102210, 102250, 
    102290, 102300, 102330, 102350, 102340, 102350, 102360, 102360, 102360, 
    102350, 102330, 102330, 102330, 102290, 102240, 102220, 102200, 102150, 
    102110, 102060, 102040, 101980, 101930, 101880, 101850, 101830, 101790, 
    101750, 101740, 101720, 101690, 101530, 101450, 101490, 101490, 101470, 
    101430, 101380, 101330, 101280, 101220, 101200, 101150, 101090, 101020, 
    100980, 100930, 100900, 100870, 100840, 100830, 100810, 100780, 100770, 
    100780, 100760, 100750, 100740, 100710, 100700, 100690, 100720, 100750, 
    100780, 100840, 100850, 100870, 100870, 100850, 100870, 100890, 100940, 
    100970, 101010, 101020, 101050, 101080, 101100, 101130, 101150, 101160, 
    101150, 101170, 101190, 101200, 101220, 101230, 101240, 101260, 101280, 
    101280, 101280, 101270, 101260, 101290, 101310, 101330, 101330, 101310, 
    101320, 101350, 101360, 101370, 101360, 101360, 101390, 101430, 101440, 
    101480, 101510, 101530, 101540, 101570, 101600, 101630, 101650, 101670, 
    101680, 101720, 101760, 101780, 101830, 101850, 101880, 101890, 101900, 
    101920, 101930, 101940, 101940, 101930, 101970, 101980, 101970, 101930, 
    101910, 101900, 101910, 101890, 101880, 101860, 101820, 101830, 101820, 
    101800, 101790, 101780, 101780, 101770, 101750, 101700, 101700, 101680, 
    101660, 101650, 101640, 101590, 101570, 101580, 101560, 101540, 101520, 
    101500, 101490, 101450, 101430, 101400, 101390, 101340, 101290, 101250, 
    101240, 101190, 101120, 101080, 101030, 100970, 100890, 100860, 100820, 
    100780, 100780, 100780, 100780, 100830, 100840, 100830, 100840, 100890, 
    100990, 101060, 101160, 101240, 101290, 101350, 101430, 101440, 101480, 
    101510, 101570, 101590, 101600, 101600, 101640, 101670, 101720, 101720, 
    101770, 101780, 101810, 101810, 101820, 101850, 101870, 101910, 101930, 
    101940, 101960, 101960, 101970, 101960, 101950, 101920, 101900, 101870, 
    101820, 101760, 101700, 101710, 101670, 101670, 101680, 101660, 101630, 
    101630, 101620, 101620, 101620, 101620, 101630, 101630, 101630, 101640, 
    101630, 101620, 101600, 101580, 101530, 101490, 101490, 101500, 101490, 
    101470, 101470, 101470, 101450, 101460, 101400, 101390, 101360, 101370, 
    101360, 101390, 101370, 101360, 101350, 101290, 101270, 101210, 101200, 
    101170, 101110, 101090, 101060, 101060, 101010, 101010, 100950, 100940, 
    100880, 100840, 100810, 100760, 100710, 100650, 100640, 100570, 100560, 
    100510, 100460, 100410, 100360, 100300, 100210, 100130, 100020, 99950, 
    99850, 99710, 99640, 99520, 99460, 99380, 99350, 99330, 99270, 99290, 
    99290, 99270, 99270, 99280, 99280, 99260, 99260, 99260, 99260, 99240, 
    99220, 99250, 99240, 99300, 99360, 99400, 99430, 99470, 99460, 99520, 
    99560, 99560, 99620, 99720, 99730, 99770, 99810, 99870, 99910, 99960, 
    100030, 100080, 100130, 100180, 100250, 100280, 100330, 100380, 100450, 
    100500, 100530, 100570, 100620, 100680, 100740, 100750, 101000, 101020, 
    101080, 101100, 101110, 101120, 101140, 101160, 101170, 101190, 101170, 
    101180, 101200, 101210, 101200, 101190, 101210, 101220, 101230, 101250, 
    101290, 101330, 101350, 101380, 101390, 101400, 101440, 101480, 101490, 
    101520, 101540, 101560, 101570, 101590, 101650, 101700, 101730, 101790, 
    101830, 101860, 101890, 101920, 101930, 101970, 101980, 102010, 102030, 
    102030, 102060, 102070, 102100, 102120, 102130, 102150, 102170, 102170, 
    102190, 102190, 102190, 102190, 102190, 102200, 102230, 102230, 102230, 
    102240, 102250, 102240, 102230, 102220, 102210, 102200, 102190, 102170, 
    102160, 102150, 102130, 102110, 102100, 102090, 102070, 102060, 102040, 
    102020, 102020, 102040, 102030, 102030, 102020, 102010, 101980, 101970, 
    101960, 101960, 101960, 101930, 101950, 101930, 101920, 101920, 101920, 
    101900, 101900, 101910, 101890, 101850, 101840, 101820, 101800, 101780, 
    101790, 101780, 101760, 101750, 101740, 101720, 101680, 101640, 101600, 
    101610, 101570, 101550, 101560, 101530, 101520, 101510, 101490, 101450, 
    101420, 101400, 101370, 101340, 101330, 101300, 101280, 101250, 101210, 
    101220, 101150, 101100, 101060, 101020, 101000, 100970, 100970, 100900, 
    100950, 100970, 100920, 100910, 100900, 100910, 100900, 100920, 100910, 
    100920, 100900, 100940, 100890, 100970, 101020, 101120, 101150, 101200, 
    101240, 101270, 101290, 101320, 101320, 101360, 101420, 101500, 101500, 
    101530, 101550, 101530, 101530, 101550, 101570, 101570, 101570, 101570, 
    101560, 101580, 101580, 101570, 101590, 101600, 101600, 101570, 101570, 
    101550, 101550, 101540, 101500, 101520, 101530, 101500, 101480, 101450, 
    101400, 101370, 101310, 101290, 101270, 101260, 101210, 101210, 101150, 
    101160, 101120, 101100, 101010, 100960, 100900, 100860, 100740, 100710, 
    100650, 100580, 100500, 100420, 100300, 100220, 100100, 100030, 99970, 
    99920, 99870, 99800, 99770, 99750, 99680, 99650, 99630, 99570, 99530, 
    99500, 99490, 99440, 99380, 99360, 99360, 99340, 99320, 99290, 99260, 
    99230, 99170, 99190, 99130, 99120, 99140, 99150, 99140, 99170, 99160, 
    99140, 99190, 99180, 99200, 99220, 99160, 99150, 99160, 99120, 99110, 
    99110, 99120, 99130, 99090, 99160, 99110, 99090, 99130, 99110, 99140, 
    99170, 99210, 99260, 99300, 99340, 99380, 99390, 99430, 99490, 99510, 
    99530, 99580, 99620, 99650, 99670, 99710, 99770, 99850, 99900, 99960, 
    100000, 100030, 100060, 100110, 100160, 100210, 100250, 100280, 100320, 
    100360, 100380, 100410, 100430, 100470, 100480, 100500, 100520, 100520, 
    100530, 100530, 100570, 100580, 100570, 100570, 100550, 100530, 100580, 
    100580, 100600, 100630, 100630, 100630, 100650, 100670, 100660, 100670, 
    100690, 100650, 100660, 100650, 100670, 100660, 100660, 100640, 100630, 
    100620, 100620, 100610, 100590, 100590, 100570, 100570, 100560, 100560, 
    100550, 100520, 100500, 100510, 100490, 100480, 100470, 100430, 100420, 
    100400, 100420, 100410, 100410, 100420, 100420, 100430, 100420, 100440, 
    100440, 100450, 100460, 100470, 100480, 100520, 100540, 100550, 100540, 
    100550, 100540, 100510, 100490, 100480, 100470, 100470, 100470, 100450, 
    100440, 100380, 100370, 100370, 100350, 100330, 100350, 100320, 100350, 
    100410, 100430, 100480, 100510, 100490, 100500, 100430, 100480, 100500, 
    100500, 100450, 100430, 100410, 100400, 100400, 100330, 100350, 100270, 
    100240, 100240, 100190, 100090, 100020, 100000, 99960, 99920, 99790, 
    99710, 99570, 99470, 99370, 99230, 99140, 99060, 99100, 99070, 99090, 
    99190, 99190, 99170, 99280, 99310, 99280, 99240, 99210, 99190, 99270, 
    99260, 99290, 99270, 99310, 99290, 99340, 99360, 99360, 99430, 99410, 
    99530, 99640, 99710, 99750, 99750, 99810, 99830, 99920, 99960, 100010, 
    100030, 100010, 99990, 99960, 99940, 99960, 99950, 99940, 99970, 99990, 
    100000, 100010, 100050, 100080, 100160, 100180, 100180, 100230, 100210, 
    100270, 100220, 100290, 100330, 100350, 100340, 100350, 100350, 100410, 
    100430, 100440, 100520, 100590, 100650, 100710, 100740, 100790, 100840, 
    100860, 100970, 100980, 100920, 100990, 101040, 101050, 101150, 101200, 
    101250, 101200, 101310, 101330, 101330, 101320, 101310, 101300, 101280, 
    101280, 101280, 101250, 101230, 101190, 101150, 101110, 101130, 101130, 
    101120, 101090, 101080, 101010, 100960, 100950, 100890, 100870, 100880, 
    100870, 100860, 100840, 100850, 100820, 100840, 100820, 100810, 100780, 
    100800, 100780, 100750, 100740, 100720, 100660, 100620, 100650, 100630, 
    100600, 100580, 100540, 100480, 100430, 100460, 100460, 100430, 100430, 
    100420, 100420, 100410, 100390, 100400, 100410, 100420, 100430, 100430, 
    100440, 100410, 100410, 100400, 100360, 100350, 100350, 100380, 100370, 
    100360, 100360, 100350, 100360, 100360, 100360, 100370, 100390, 100410, 
    100430, 100460, 100490, 100520, 100550, 100570, 100590, 100620, 100640, 
    100660, 100670, 100690, 100710, 100720, 100740, 100780, 100800, 100820, 
    100840, 100880, 100910, 100950, 100960, 101010, 101040, 101050, 101080, 
    101120, 101120, 101160, 101170, 101190, 101200, 101220, 101240, 101260, 
    101290, 101310, 101310, 101340, 101340, 101370, 101380, 101400, 101400, 
    101410, 101420, 101420, 101440, 101460, 101480, 101480, 101480, 101490, 
    101500, 101500, 101530, 101540, 101540, 101570, 101580, 101580, 101610, 
    101640, 101640, 101650, 101640, 101650, 101670, 101680, 101690, 101730, 
    101760, 101800, 101810, 101860, 101870, 101910, 101930, 101950, 101980, 
    102000, 102020, 102060, 102080, 102110, 102120, 102130, 102150, 102150, 
    102150, 102180, 102180, 102190, 102200, 102220, 102220, 102230, 102240, 
    102260, 102250, 102270, 102250, 102250, 102260, 102250, 102240, 102240, 
    102250, 102260, 102250, 102270, 102270, 102280, 102280, 102260, 102250, 
    102250, 102260, 102250, 102240, 102260, 102260, 102260, 102260, 102250, 
    102240, 102220, 102200, 102190, 102210, 102180, 102200, 102180, 102190, 
    102170, 102170, 102170, 102140, 102140, 102110, 102080, 102080, 102090, 
    102100, 102080, 102060, 102060, 102030, 102010, 101990, 101990, 101970, 
    101970, 101950, 101950, 101940, 101930, 101910, 101900, 101880, 101860, 
    101880, 101850, 101810, 101800, 101790, 101770, 101770, 101760, 101740, 
    101730, 101720, 101710, 101690, 101680, 101660, 101580, 101560, 101580, 
    101580, 101560, 101580, 101590, 101600, 101590, 101590, 101550, 101580, 
    101590, 101590, 101600, 101600, 101600, 101570, 101540, 101530, 101530, 
    101500, 101490, 101480, 101450, 101430, 101410, 101390, 101370, 101350, 
    101340, 101330, 101340, 101340, 101300, 101290, 101280, 101270, 101280, 
    101290, 101320, 101330, 101340, 101360, 101370, 101370, 101390, 101410, 
    101420, 101440, 101480, 101490, 101520, 101540, 101550, 101580, 101600, 
    101600, 101620, 101640, 101650, 101660, 101670, 101710, 101740, 101760, 
    101780, 101770, 101770, 101780, 101790, 101790, 101770, 101750, 101750, 
    101750, 101760, 101730, 101730, 101710, 101680, 101640, 101640, 101620, 
    101610, 101580, 101580, 101560, 101540, 101480, 101450, 101450, 101430, 
    101430, 101410, 101390, 101380, 101370, 101340, 101380, 101390, 101390, 
    101390, 101400, 101380, 101400, 101420, 101430, 101470, 101480, 101540, 
    101610, 101650, 101680, 101690, 101710, 101740, 101770, 101770, 101750, 
    101730, 101720, 101690, 101680, 101710, 101740, 101740, 101720, 101710, 
    101710, 101710, 101700, 101680, 101690, 101710, 101700, 101690, 101700, 
    101720, 101690, 101680, 101680, 101670, 101630, 101630, 101620, 101600, 
    101560, 101580, 101580, 101540, 101520, 101490, 101470, 101450, 101460, 
    101440, 101440, 101430, 101430, 101430, 101420, 101420, 101390, 101350, 
    101340, 101360, 101340, 101330, 101310, 101330, 101330, 101330, 101330, 
    101350, 101350, 101360, 101370, 101380, 101400, 101430, 101450, 101480, 
    101500, 101550, 101590, 101630, 101660, 101680, 101710, 101740, 101750, 
    101760, 101780, 101790, 101820, 101830, 101850, 101870, 101870, 101910, 
    101920, 101940, 101980, 102000, 102040, 102080, 102120, 102170, 102190, 
    102230, 102280, 102310, 102320, 102350, 102360, 102400, 102390, 102400, 
    102410, 102430, 102430, 102450, 102460, 102470, 102460, 102480, 102480, 
    102490, 102510, 102530, 102550, 102580, 102590, 102610, 102630, 102640, 
    102650, 102680, 102680, 102690, 102670, 102650, 102660, 102650, 102640, 
    102630, 102620, 102610, 102590, 102580, 102560, 102550, 102540, 102550, 
    102570, 102550, 102530, 102510, 102480, 102470, 102430, 102420, 102410, 
    102320, 102350, 102400, 102410, 102350, 102260, 102270, 102270, 102260, 
    102230, 102210, 102160, 102100, 102080, 102010, 102070, 102040, 102010, 
    102020, 101990, 102030, 102030, 102010, 101990, 102040, 102050, 102070, 
    102100, 102120, 102140, 102160, 102180, 102200, 102210, 102240, 102190, 
    102260, 102280, 102250, 102320, 102320, 102330, 102380, 102340, 102350, 
    102380, 102400, 102360, 102340, 102360, 102340, 102350, 102350, 102350, 
    102340, 102320, 102300, 102280, 102250, 102230, 102190, 102200, 102220, 
    102200, 102190, 102200, 102230, 102260, 102300, 102320, 102270, 102280, 
    102290, 102300, 102310, 102330, 102320, 102340, 102350, 102320, 102340, 
    102340, 102340, 102360, 102300, 102340, 102370, 102360, 102360, 102370, 
    102390, 102350, 102320, 102340, 102350, 102290, 102310, 102280, 102270, 
    102260, 102370, 102360, 102240, 102240, 102240, 102240, 102240, 102200, 
    102220, 102190, 102230, 102210, 102250, 102290, 102290, 102280, 102290, 
    102310, 102290, 102280, 102270, 102270, 102300, 102330, 102300, 102330, 
    102320, 102370, 102360, 102370, 102360, 102370, 102360, 102360, 102380, 
    102380, 102400, 102360, 102360, 102350, 102360, 102320, 102320, 102330, 
    102320, 102300, 102230, 102190, 102200, 102200, 102160, 102130, 102120, 
    102130, 102070, 102050, 102010, 102000, 102000, 101980, 101950, 101930, 
    101930, 101900, 101860, 101820, 101810, 101790, 101760, 101720, 101680, 
    101640, 101610, 101580, 101550, 101510, 101480, 101460, 101420, 101360, 
    101320, 101290, 101270, 101260, 101240, 101210, 101230, 101220, 101170, 
    101140, 101100, 101090, 101080, 101040, 101020, 101000, 101010, 101030, 
    101040, 101070, 101050, 101030, 101030, 101040, 100990, 100940, 100890, 
    100850, 100770, 100740, 100670, 100690, 100650, 100650, 100640, 100640, 
    100640, 100660, 100700, 100730, 100740, 100760, 100780, 100750, 100710, 
    100690, 100680, 100610, 100630, 100660, 100710, 100820, 100870, 100910, 
    100910, 100950, 100970, 101010, 101030, 101050, 101070, 101080, 101120, 
    101150, 101170, 101210, 101320, 101220, 101260, 101300, 101330, 101320, 
    101350, 101390, 101380, 101410, 101460, 101460, 101430, 101460, 101590, 
    101590, 101610, 101600, 101640, 101620, 101620, 101630, 101600, 101550, 
    101510, 101480, 101510, 101510, 101480, 101490, 101480, 101480, 101490, 
    101520, 101520, 101540, 101550, 101560, 101590, 101610, 101620, 101600, 
    101600, 101610, 101620, 101630, 101650, 101680, 101690, 101690, 101670, 
    101700, 101710, 101740, 101740, 101740, 101740, 101740, 101740, 101760, 
    101770, 101770, 101770, 101770, 101790, 101750, 101750, 101720, 101680, 
    101680, 101750, 101770, 101790, 101810, 101800, 101780, 101770, 101760, 
    101760, 101740, 101740, 101760, 101750, 101740, 101800, 101800, 101800, 
    101820, 101790, 101750, 101740, 101710, 101680, 101640, 101670, 101690, 
    101680, 101670, 101660, 101640, 101630, 101610, 101580, 101540, 101550, 
    101550, 101510, 101510, 101540, 101520, 101540, 101530, 101510, 101480, 
    101480, 101450, 101440, 101410, 101390, 101400, 101370, 101340, 101310, 
    101260, 101330, 101300, 101260, 101210, 101140, 101080, 101050, 101000, 
    100940, 100890, 100810, 100790, 100700, 100630, 100610, 100570, 100520, 
    100470, 100460, 100400, 100430, 100370, 100370, 100340, 100300, 100260, 
    100280, 100290, 100320, 100330, 100350, 100390, 100410, 100410, 100410, 
    100410, 100400, 100340, 100310, 100290, 100260, 100230, 100210, 100180, 
    100170, 100140, 100100, 100060, 100050, 100030, 100000, 99980, 100040, 
    100040, 100100, 100150, 100170, 100210, 100260, 100310, 100350, 100390, 
    100430, 100480, 100560, 100620, 100660, 100690, 100720, 100760, 100800, 
    100850, 100880, 100930, 100930, 100980, 100990, 101010, 101030, 101070, 
    101070, 101090, 101100, 101120, 101120, 101140, 101160, 101190, 101220, 
    101250, 101290, 101340, 101390, 101440, 101490, 101540, 101600, 101650, 
    101700, 101740, 101780, 101820, 101850, 101890, 101920, 101960, 102000, 
    102020, 102030, 102070, 102120, 102140, 102160, 102180, 102230, 102280, 
    102310, 102320, 102340, 102340, 102330, 102340, 102370, 102400, 102400, 
    102450, 102410, 102400, 102480, 102510, 102510, 102510, 102510, 102510, 
    102500, 102480, 102490, 102460, 102480, 102470, 102470, 102470, 102450, 
    102420, 102410, 102410, 102400, 102380, 102350, 102330, 102300, 102300, 
    102280, 102250, 102220, 102170, 102090, 101980, 101970, 101950, 101950, 
    101910, 101840, 101850, 101900, 101890, 101840, 101840, 101810, 101850, 
    101860, 101880, 101850, 101860, 101880, 101920, 101930, 101950, 101940, 
    102010, 102030, 101980, 102000, 102040, 102080, 102130, 102150, 102170, 
    102180, 102200, 102210, 102290, 102290, 102320, 102350, 102370, 102370, 
    102350, 102460, 102440, 102410, 102430, 102470, 102470, 102470, 102460, 
    102440, 102420, 102440, 102420, 102390, 102360, 102330, 102380, 102390, 
    102390, 102390, 102390, 102410, 102400, 102400, 102350, 102350, 102360, 
    102360, 102390, 102370, 102350, 102330, 102350, 102380, 102340, 102350, 
    102340, 102330, 102320, 102410, 102400, 102400, 102390, 102380, 102380, 
    102400, 102390, 102380, 102400, 102410, 102420, 102430, 102420, 102450, 
    102460, 102440, 102440, 102440, 102450, 102450, 102450, 102460, 102460, 
    102450, 102430, 102410, 102470, 102390, 102380, 102380, 102410, 102410, 
    102400, 102390, 102390, 102380, 102390, 102380, 102360, 102340, 102320, 
    102310, 102300, 102300, 102290, 102310, 102300, 102270, 102270, 102270, 
    102240, 102240, 102250, 102250, 102250, 102270, 102270, 102290, 102310, 
    102320, 102310, 102310, 102320, 102320, 102320, 102290, 102250, 102230, 
    102250, 102280, 102300, 102280, 102240, 102240, 102250, 102250, 102250, 
    102250, 102230, 102250, 102280, 102310, 102330, 102330, 102340, 102350, 
    102360, 102360, 102360, 102350, 102340, 102330, 102320, 102340, 102320, 
    102320, 102290, 102300, 102290, 102260, 102230, 102210, 102190, 102160, 
    102130, 102110, 102070, 102050, 102000, 101950, 101910, 101840, 101790, 
    101760, 101700, 101670, 101630, 101630, 101590, 101570, 101510, 101500, 
    101450, 101400, 101370, 101320, 101290, 101280, 101260, 101250, 101230, 
    101220, 101180, 101160, 101140, 101120, 101110, 101090, 101070, 101050, 
    101020, 101030, 101030, 101030, 101010, 101000, 100980, 100980, 100960, 
    100960, 100970, 100980, 101000, 101030, 101050, 101060, 101080, 101090, 
    101110, 101110, 101110, 101110, 101140, 101130, 101160, 101180, 101210, 
    101220, 101250, 101250, 101250, 101260, 101270, 101280, 101310, 101340, 
    101360, 101380, 101410, 101410, 101410, 101410, 101420, 101400, 101400, 
    101390, 101350, 101330, 101340, 101350, 101340, 101350, 101340, 101350, 
    101340, 101350, 101350, 101340, 101340, 101360, 101370, 101380, 101400, 
    101400, 101410, 101410, 101400, 101410, 101430, 101420, 101430, 101450, 
    101450, 101460, 101480, 101480, 101480, 101480, 101490, 101500, 101500, 
    101490, 101500, 101520, 101540, 101560, 101580, 101590, 101610, 101610, 
    101630, 101630, 101640, 101670, 101680, 101680, 101710, 101710, 101730, 
    101760, 101760, 101760, 101770, 101780, 101800, 101820, 101790, 101820, 
    101820, 101830, 101820, 101840, 101850, 101840, 101830, 101830, 101820, 
    101800, 101780, 101780, 101760, 101750, 101720, 101710, 101670, 101630, 
    101600, 101570, 101530, 101500, 101480, 101450, 101460, 101450, 101430, 
    101400, 101390, 101380, 101360, 101330, 101320, 101320, 101300, 101290, 
    101270, 101250, 101240, 101220, 101210, 101200, 101200, 101200, 101200, 
    101210, 101210, 101210, 101230, 101240, 101270, 101310, 101320, 101340, 
    101370, 101390, 101410, 101430, 101450, 101480, 101510, 101560, 101610, 
    101650, 101680, 101730, 101760, 101780, 101800, 101830, 101890, 101980, 
    102020, 102060, 102140, 102210, 102260, 102300, 102340, 102370, 102390, 
    102410, 102460, 102510, 102570, 102600, 102630, 102670, 102690, 102700, 
    102710, 102710, 102710, 102710, 102750, 102770, 102780, 102780, 102810, 
    102830, 102820, 102810, 102810, 102810, 102800, 102770, 102740, 102720, 
    102710, 102690, 102680, 102650, 102620, 102600, 102580, 102540, 102540, 
    102510, 102450, 102450, 102470, 102480, 102490, 102500, 102500, 102480, 
    102500, 102470, 102430, 102450, 102420, 102390, 102380, 102370, 102300, 
    102270, 102260, 102230, 102190, 102130, 102040, 102000, 101910, 101860, 
    101840, 101780, 101720, 101670, 101570, 101520, 101490, 101380, 101320, 
    101220, 101160, 101120, 101050, 101040, 101030, 101020, 101020, 100980, 
    100950, 100920, 100890, 100930, 100920, 100930, 100960, 100980, 101000, 
    101070, 101140, 101220, 101220, 101230, 101200, 101180, 101150, 101120, 
    101130, 101120, 101110, 101150, 101170, 101150, 101120, 101100, 101070, 
    101060, 101060, 101050, 101070, 101030, 101000, 101000, 100980, 100970, 
    100940, 100900, 100910, 100890, 100890, 100910, 100940, 100980, 101010, 
    101010, 101040, 101040, 101050, 101050, 101050, 101070, 101090, 101060, 
    101070, 101090, 101100, 101100, 101100, 101080, 101100, 101120, 101130, 
    101150, 101190, 101220, 101260, 101310, 101400, 101460, 101510, 101550, 
    101580, 101610, 101630, 101650, 101640, 101710, 101770, 101820, 101870, 
    101940, 101950, 101970, 102040, 102110, 102190, 102210, 102230, 102270, 
    102330, 102370, 102410, 102440, 102480, 102530, 102540, 102540, 102560, 
    102600, 102620, 102660, 102700, 102740, 102750, 102760, 102800, 102820, 
    102820, 102850, 102860, 102870, 102860, 102860, 102850, 102830, 102800, 
    102800, 102750, 102700, 102620, 102550, 102510, 102430, 102380, 102350, 
    102320, 102290, 102230, 102170, 102110, 102080, 102020, 101970, 101930, 
    101900, 101870, 101840, 101820, 101800, 101780, 101750, 101770, 101770, 
    101780, 101790, 101790, 101780, 101780, 101820, 101850, 101860, 101890, 
    101920, 101950, 101960, 101970, 102000, 102020, 102020, 102030, 102040, 
    102040, 102040, 102040, 102010, 101990, 101990, 101960, 101940, 101920, 
    101900, 101860, 101850, 101840, 101840, 101820, 101780, 101760, 101730, 
    101690, 101650, 101620, 101600, 101570, 101550, 101550, 101580, 101570, 
    101540, 101490, 101490, 101470, 101440, 101410, 101460, 101440, 101400, 
    101380, 101410, 101410, 101390, 101390, 101350, 101430, 101400, 101390, 
    101420, 101420, 101430, 101460, 101460, 101470, 101500, 101520, 101540, 
    101550, 101560, 101560, 101570, 101570, 101600, 101610, 101630, 101660, 
    101670, 101710, 101740, 101740, 101740, 101750, 101760, 101750, 101740, 
    101750, 101750, 101770, 101780, 101800, 101800, 101820, 101820, 101830, 
    101830, 101820, 101830, 101840, 101860, 101880, 101870, 101890, 101890, 
    101880, 101870, 101850, 101840, 101810, 101800, 101760, 101740, 101740, 
    101700, 101640, 101590, 101530, 101460, 101410, 101370, 101380, 101320, 
    101270, 101260, 101210, 101170, 101140, 101120, 101090, 101080, 101080, 
    101070, 101100, 101100, 101130, 101160, 101190, 101220, 101270, 101290, 
    101320, 101350, 101340, 101350, 101370, 101370, 101380, 101390, 101390, 
    101380, 101370, 101350, 101350, 101360, 101340, 101310, 101280, 101260, 
    101270, 101260, 101230, 101210, 101200, 101190, 101180, 101180, 101150, 
    101160, 101160, 101150, 101150, 101170, 101170, 101190, 101210, 101200, 
    101210, 101210, 101200, 101170, 101180, 101150, 101170, 101210, 101230, 
    101200, 101230, 101300, 101300, 101300, 101320, 101340, 101360, 101410, 
    101450, 101490, 101520, 101520, 101510, 101530, 101570, 101590, 101580, 
    101570, 101550, 101540, 101510, 101520, 101510, 101520, 101490, 101500, 
    101500, 101460, 101440, 101450, 101380, 101320, 101340, 101310, 101340, 
    101340, 101320, 101310, 101300, 101240, 101220, 101200, 101090, 101130, 
    101010, 101020, 100980, 100950, 100960, 100890, 100860, 100880, 100820, 
    100770, 100830, 100850, 100820, 100810, 100820, 100830, 100800, 100780, 
    100820, 100830, 100800, 100760, 100760, 100700, 100670, 100650, 100520, 
    100490, 100470, 100460, 100400, 100410, 100330, 100290, 100270, 100280, 
    100260, 100200, 100190, 100190, 100180, 100180, 100200, 100200, 100190, 
    100180, 100170, 100150, 100180, 100230, 100240, 100280, 100350, 100420, 
    100440, 100450, 100480, 100500, 100510, 100530, 100570, 100630, 100660, 
    100700, 100730, 100760, 100780, 100800, 100820, 100830, 100890, 100920, 
    100960, 100990, 101020, 101050, 101070, 101090, 101100, 101120, 101130, 
    101130, 101170, 101190, 101230, 101260, 101270, 101290, 101320, 101320, 
    101330, 101330, 101320, 101310, 101290, 101280, 101260, 101240, 101220, 
    101170, 101110, 101050, 100990, 100960, 100960, 100940, 100920, 100880, 
    100890, 100870, 100850, 100830, 100800, 100740, 100660, 100550, 100490, 
    100380, 100330, 100290, 100220, 100140, 100060, 99930, 99860, 99810, 
    99760, 99740, 99730, 99730, 99730, 99740, 99710, 99740, 99750, 99760, 
    99760, 99740, 99750, 99760, 99750, 99730, 99740, 99770, 99780, 99760, 
    99760, 99770, 99770, 99770, 99850, 99880, 99880, 99920, 100030, 100080, 
    100130, 100160, 100230, 100270, 100360, 100430, 100440, 100500, 100570, 
    100560, 100610, 100710, 100750, 100800, 100870, 100940, 101000, 101030, 
    101080, 101070, 101030, 101040, 101010, 101010, 100980, 100950, 100940, 
    100910, 100860, 100790, 100750, 100720, 100670, 100660, 100630, 100620, 
    100630, 100630, 100680, 100710, 100720, 100780, 100810, 100880, 100910, 
    100940, 100960, 100950, 100970, 100950, 100960, 100920, 100870, 100780, 
    100720, 100650, 100580, 100540, 100520, 100500, 100520, 100530, 100590, 
    100600, 100680, 100710, 100760, 100810, 100880, 100920, 100990, 101060, 
    101120, 101190, 101250, 101270, 101390, 101440, 101480, 101510, 101540, 
    101560, 101560, 101570, 101550, 101550, 101530, 101480, 101420, 101360, 
    101320, 101260, 101200, 101150, 101120, 101130, 101150, 101170, 101230, 
    101280, 101340, 101390, 101420, 101450, 101480, 101500, 101560, 101600, 
    101640, 101690, 101720, 101730, 101720, 101720, 101730, 101750, 101720, 
    101680, 101650, 101620, 101620, 101590, 101580, 101520, 101510, 101450, 
    101400, 101350, 101350, 101310, 101280, 101220, 101180, 101180, 101160, 
    101110, 101050, 101070, 101050, 101060, 101100, 101160, 101210, 101280, 
    101360, 101410, 101440, 101500, 101570, 101620, 101660, 101660, 101700, 
    101750, 101780, 101790, 101830, 101840, 101850, 101850, 101830, 101830, 
    101820, 101810, 101780, 101790, 101800, 101740, 101740, 101730, 101690, 
    101670, 101660, 101670, 101620, 101580, 101550, 101520, 101500, 101440, 
    101390, 101320, 101290, 101230, 101220, 101130, 101080, 101040, 101020, 
    101030, 101020, 101010, 101000, 101000, 100970, 101000, 101020, 101040, 
    101050, 101060, 101040, 101050, 101130, 101230, 101270, 101290, 101300, 
    101310, 101320, 101350, 101350, 101360, 101400, 101460, 101470, 101460, 
    101440, 101500, 101580, 101660, 101680, 101720, 101740, 101760, 101780, 
    101770, 101780, 101820, 101780, 101790, 101790, 101780, 101790, 101820, 
    101810, 101780, 101800, 101810, 101780, 101770, 101780, 101790, 101790, 
    101790, 101790, 101750, 101720, 101670, 101660, 101610, 101580, 101560, 
    101530, 101500, 101460, 101430, 101390, 101380, 101340, 101300, 101250, 
    101230, 101190, 101170, 101170, 101170, 101170, 101170, 101180, 101170, 
    101170, 101170, 101150, 101140, 101130, 101160, 101160, 101180, 101210, 
    101270, 101280, 101300, 101340, 101360, 101400, 101410, 101430, 101460, 
    101490, 101510, 101580, 101610, 101650, 101710, 101710, 101730, 101750, 
    101780, 101740, 101800, 101810, 101810, 101800, 101780, 101750, 101720, 
    101650, 101640, 101560, 101480, 101440, 101380, 101310, 101310, 101290, 
    101260, 101230, 101190, 101150, 101110, 101050, 101000, 100940, 100960, 
    100930, 100920, 100890, 100880, 100920, 100880, 100900, 100920, 100930, 
    100980, 101000, 101040, 101070, 101110, 101130, 101200, 101220, 101250, 
    101270, 101340, 101360, 101350, 101390, 101430, 101510, 101510, 101540, 
    101550, 101570, 101590, 101590, 101580, 101580, 101590, 101580, 101600, 
    101610, 101620, 101600, 101610, 101600, 101570, 101550, 101520, 101510, 
    101500, 101480, 101480, 101460, 101430, 101430, 101410, 101380, 101370, 
    101360, 101360, 101350, 101360, 101360, 101380, 101390, 101400, 101410, 
    101440, 101440, 101470, 101470, 101490, 101530, 101540, 101560, 101590, 
    101620, 101640, 101680, 101710, 101760, 101770, 101800, 101830, 101880, 
    101920, 101950, 102000, 102050, 102110, 102140, 102170, 102210, 102240, 
    102250, 102290, 102320, 102350, 102380, 102410, 102450, 102490, 102530, 
    102570, 102590, 102610, 102650, 102700, 102740, 102770, 102770, 102820, 
    102870, 102900, 102910, 102940, 102950, 102960, 102960, 102950, 102950, 
    102950, 102910, 102860, 102800, 102770, 102740, 102710, 102660, 102630, 
    102610, 102530, 102490, 102440, 102340, 102280, 102180, 102140, 102060, 
    101990, 101950, 101870, 101820, 101740, 101670, 101560, 101490, 101390, 
    101260, 101100, 100940, 100770, 100730, 100710, 100740, 100740, 100700, 
    100570, 100420, 100300, 100220, 100120, 100010, 99890, 99710, 99390, 
    99130, 98750, 98360, 98180, 97930, 97620, 97400, 97230, 97100, 96930, 
    96800, 96650, 96490, 96360, 96250, 96150, 96040, 96010, 95990, 96040, 
    96090, 96150, 96200, 96350, 96460, 96620, 96840, 97050, 97190, 97350, 
    97450, 97560, 97670, 97730, 97830, 97930, 98000, 98130, 98200, 98250, 
    98340, 98400, 98470, 98550, 98610, 98670, 98710, 98770, 98840, 98880, 
    98910, 99040, 99100, 99130, 99180, 99220, 99250, 99290, 99310, 99330, 
    99350, 99370, 99380, 99410, 99370, 99400, 99430, 99450, 99480, 99500, 
    99530, 99560, 99580, 99590, 99620, 99650, 99680, 99710, 99740, 99770, 
    99810, 99860, 99910, 99960, 100010, 100060, 100080, 100110, 100200, 
    100260, 100320, 100360, 100420, 100480, 100530, 100580, 100630, 100670, 
    100700, 100740, 100800, 100840, 100860, 100880, 100910, 100940, 100970, 
    101000, 101030, 101050, 101080, 101080, 100920, 100950, 100970, 100990, 
    101020, 101070, 101100, 101140, 101190, 101220, 101230, 101270, 101360, 
    101410, 101450, 101480, 101510, 101550, 101600, 101650, 101710, 101760, 
    101810, 101870, 101940, 102010, 102060, 102120, 102170, 102220, 102270, 
    102320, 102380, 102420, 102420, 102440, 102440, 102490, 102530, 102550, 
    102590, 102610, 102650, 102650, 102680, 102700, 102740, 102760, 102770, 
    102780, 102830, 102850, 102890, 102900, 102880, 102920, 102910, 102920, 
    102910, 102890, 102880, 102900, 102900, 102890, 102890, 102900, 102890, 
    102880, 102910, 102920, 102930, 102920, 102970, 103010, 103020, 103050, 
    103060, 103100, 103100, 103120, 103120, 103130, 103140, 103160, 103140, 
    103130, 103150, 103130, 103120, 103100, 103060, 103030, 103030, 102990, 
    102960, 102930, 102890, 102880, 102860, 102870, 102870, 102820, 102790, 
    102760, 102770, 102750, 102720, 102690, 102690, 102670, 102670, 102660, 
    102640, 102580, 102620, 102610, 102570, 102580, 102550, 102600, 102570, 
    102580, 102590, 102590, 102610, 102570, 102550, 102530, 102490, 102500, 
    102470, 102440, 102400, 102380, 102310, 102310, 102300, 102270, 102230, 
    102180, 102120, 102110, 102050, 102010, 102010, 101990, 101970, 101970, 
    101940, 101910, 101880, 101850, 101800, 101750, 101780, 101720, 101650, 
    101610, 101560, 101510, 101450, 101410, 101370, 101340, 101310, 101260, 
    101230, 101160, 101100, 101090, 101090, 101090, 101060, 101030, 101010, 
    100950, 100920, 100870, 100840, 100840, 100820, 100800, 100760, 100740, 
    100730, 100740, 100710, 100700, 100710, 100680, 100680, 100710, 100720, 
    100720, 100710, 100760, 100810, 100820, 100870, 100890, 100920, 100940, 
    100970, 100990, 101010, 101020, 101040, 101050, 101070, 101080, 101110, 
    101090, 101130, 101120, 101140, 101130, 101130, 101110, 101130, 101130, 
    101150, 101150, 101180, 101190, 101220, 101210, 101220, 101240, 101250, 
    101270, 101290, 101310, 101350, 101380, 101380, 101390, 101400, 101400, 
    101410, 101430, 101420, 101420, 101420, 101420, 101370, 101380, 101370, 
    101350, 101330, 101300, 101250, 101240, 101190, 101140, 101130, 101080, 
    101040, 101010, 100950, 100910, 100860, 100800, 100770, 100640, 100590, 
    100490, 100340, 100240, 100140, 100090, 99970, 99780, 99660, 99510, 
    99320, 99160, 98980, 98810, 98590, 98380, 98190, 98090, 98120, 98210, 
    98360, 98490, 98560, 98670, 98730, 98820, 98880, 98950, 99000, 99110, 
    99110, 99120, 99140, 99160, 99220, 99240, 99300, 99320, 99360, 99400, 
    99400, 99430, 99550, 99570, 99650, 99680, 99730, 99790, 99820, 99880, 
    99930, 99990, 100060, 100150, 100160, 100190, 100240, 100250, 100280, 
    100290, 100300, 100310, 100340, 100380, 100420, 100450, 100460, 100490, 
    100510, 100530, 100560, 100570, 100580, 100620, 100630, 100630, 100650, 
    100630, 100610, 100580, 100530, 100480, 100420, 100360, 100290, 100210, 
    100140, 100090, 100010, 99910, 99820, 99720, 99610, 99470, 99370, 99300, 
    99250, 99200, 99180, 99180, 99160, 99150, 99110, 99070, 99070, 99060, 
    99060, 99090, 99130, 99230, 99340, 99420, 99510, 99620, 99710, 99810, 
    99870, 99910, 99970, 100040, 100130, 100180, 100210, 100280, 100340, 
    100410, 100470, 100530, 100570, 100610, 100630, 100670, 100710, 100730, 
    100750, 100770, 100780, 100790, 100810, 100840, 100840, 100830, 100830, 
    100830, 100830, 100820, 100840, 100810, 100770, 100730, 100720, 100700, 
    100660, 100620, 100570, 100550, 100520, 100500, 100460, 100430, 100420, 
    100410, 100380, 100360, 100310, 100310, 100280, 100250, 100250, 100250, 
    100240, 100220, 100210, 100180, 100200, 100210, 100190, 100220, 100190, 
    100200, 100200, 100210, 100170, 100180, 100200, 100200, 100210, 100200, 
    100220, 100210, 100230, 100240, 100270, 100250, 100290, 100330, 100340, 
    100360, 100390, 100430, 100410, 100420, 100410, 100400, 100390, 100390, 
    100330, 100280, 100250, 100210, 100160, 100080, 99950, 99840, 99700, 
    99670, 99560, 99400, 99350, 99260, 99290, 99290, 99250, 99200, 99090, 
    99030, 98990, 98890, 98830, 98720, 98660, 98570, 98500, 98340, 98120, 
    97880, 97820, 97690, 97700, 97650, 97620, 97620, 97590, 97570, 97500, 
    97460, 97420, 97410, 97390, 97390, 97460, 97520, 97580, 97680, 97810, 
    97930, 97980, 98120, 98180, 98180, 98310, 98290, 98390, 98540, 98760, 
    98920, 99010, 99110, 99280, 99430, 99560, 99610, 99670, 99770, 99870, 
    99980, 100020, 100100, 100170, 100220, 100270, 100320, 100360, 100390, 
    100420, 100470, 100480, 100510, 100540, 100560, 100590, 100610, 100630, 
    100660, 100670, 100660, 100630, 100640, 100610, 100600, 100580, 100570, 
    100580, 100590, 100620, 100600, 100630, 100630, 100620, 100630, 100650, 
    100710, 100750, 100780, 100830, 100870, 100890, 100950, 101010, 101060, 
    101120, 101180, 101210, 101260, 101280, 101290, 101340, 101380, 101400, 
    101430, 101440, 101480, 101520, 101560, 101570, 101610, 101640, 101660, 
    101680, 101720, 101730, 101730, 101740, 101780, 101750, 101760, 101770, 
    101770, 101770, 101800, 101780, 101800, 101760, 101770, 101720, 101710, 
    101670, 101580, 101490, 101430, 101390, 101310, 101330, 101310, 101220, 
    101190, 101170, 101160, 101160, 101090, 101100, 101080, 101110, 101100, 
    101110, 101090, 101080, 101040, 101010, 100980, 100920, 100900, 100870, 
    100830, 100780, 100700, 100700, 100690, 100660, 100590, 100540, 100500, 
    100430, 100370, 100280, 100220, 100090, 100100, 100040, 99990, 99890, 
    99850, 99760, 99630, 99560, 99470, 99390, 99300, 99190, 99060, 98990, 
    98970, 98940, 98910, 98880, 98820, 98820, 98780, 98740, 98740, 98740, 
    98720, 98710, 98710, 98710, 98700, 98720, 98690, 98690, 98720, 98720, 
    98720, 98750, 98770, 98770, 98780, 98730, 98760, 98800, 98810, 98860, 
    98860, 98880, 98880, 98900, 98930, 98960, 98980, 99060, 99100, 99160, 
    99220, 99290, 99360, 99400, 99440, 99560, 99590, 99600, 99670, 99720, 
    99750, 99770, 99740, 99750, 99740, 99730, 99710, 99670, 99660, 99650, 
    99570, 99560, 99530, 99520, 99500, 99490, 99450, 99410, 99390, 99390, 
    99410, 99450, 99500, 99520, 99550, 99600, 99650, 99700, 99780, 99840, 
    99870, 99930, 99990, 100040, 100110, 100210, 100300, 100410, 100490, 
    100560, 100620, 100660, 100740, 100800, 100860, 100890, 100930, 100990, 
    101010, 101020, 101020, 101040, 101000, 100950, 100900, 100910, 100990, 
    101100, 101140, 101150, 101160, 101150, 101120, 101110, 101160, 101200, 
    101240, 101300, 101360, 101400, 101400, 101370, 101320, 101320, 101300, 
    101290, 101270, 101260, 101240, 101250, 101220, 101200, 101180, 101140, 
    101130, 101110, 101100, 101090, 101100, 101100, 101070, 101070, 101040, 
    101080, 101050, 101020, 100990, 100940, 100910, 100840, 100770, 100700, 
    100650, 100580, 100550, 100540, 100540, 100570, 100560, 100530, 100510, 
    100490, 100490, 100430, 100390, 100390, 100370, 100290, 100230, 100190, 
    100150, 100090, 100020, 99930, 99860, 99790, 99730, 99670, 99610, 99570, 
    99540, 99460, 99360, 99320, 99330, 99390, 99440, 99450, 99510, 99520, 
    99530, 99600, 99610, 99590, 99600, 99620, 99650, 99630, 99750, 99770, 
    99800, 99860, 99850, 99860, 99880, 99910, 99900, 99950, 99980, 99970, 
    99980, 99980, 99980, 99990, 100040, 100070, 100100, 100120, 100130, 
    100110, 100120, 100140, 100170, 100190, 100200, 100180, 100210, 100260, 
    100270, 100300, 100300, 100320, 100340, 100390, 100410, 100440, 100480, 
    100530, 100540, 100610, 100730, 100820, 100870, 100920, 100990, 101050, 
    101110, 101150, 101180, 101200, 101280, 101330, 101380, 101450, 101500, 
    101530, 101580, 101670, 101730, 101760, 101840, 101890, 101930, 101980, 
    102050, 102100, 102170, 102200, 102240, 102310, 102370, 102410, 102460, 
    102510, 102540, 102600, 102630, 102660, 102710, 102730, 102760, 102810, 
    102830, 102830, 102830, 102850, 102860, 102880, 102890, 102900, 102900, 
    102890, 102870, 102870, 102840, 102830, 102820, 102770, 102750, 102710, 
    102660, 102620, 102580, 102520, 102460, 102390, 102310, 102200, 102130, 
    102050, 102010, 101970, 101940, 101900, 101860, 101820, 101760, 101690, 
    101640, 101570, 101510, 101480, 101430, 101380, 101340, 101260, 101140, 
    101090, 101040, 100970, 100860, 100770, 100630, 100490, 100410, 100330, 
    100220, 100150, 100020, 99980, 99900, 99870, 99810, 99780, 99750, 99740, 
    99730, 99720, 99750, 99780, 99810, 99830, 99820, 99840, 99890, 99920, 
    99900, 99880, 99890, 99880, 99890, 99870, 99850, 99790, 99710, 99650, 
    99590, 99560, 99520, 99520, 99490, 99430, 99400, 99350, 99300, 99260, 
    99190, 99110, 99050, 99080, 99060, 99040, 99060, 99090, 99130, 99150, 
    99180, 99200, 99200, 99200, 99210, 99220, 99230, 99250, 99260, 99290, 
    99320, 99340, 99340, 99330, 99340, 99330, 99330, 99370, 99460, 99510, 
    99550, 99600, 99660, 99680, 99720, 99720, 99750, 99770, 99840, 99890, 
    99920, 99970, 100000, 100010, 100070, 100080, 100080, 100090, 100110, 
    100110, 100090, 100070, 100070, 100030, 100000, 99960, 99950, 99910, 
    99850, 99760, 99660, 99580, 99470, 99360, 99230, 99090, 98990, 98830, 
    98700, 98590, 98530, 98450, 98370, 98300, 98260, 98210, 98150, 98090, 
    98040, 97980, 97960, 97950, 97940, 97890, 97940, 97970, 98050, 98080, 
    98170, 98240, 98310, 98390, 98540, 98680, 98780, 98880, 98970, 99060, 
    99150, 99240, 99310, 99380, 99470, 99530, 99600, 99640, 99680, 99710, 
    99720, 99770, 99790, 99800, 99840, 99870, 99850, 99850, 99840, 99840, 
    99840, 99790, 99740, 99690, 99610, 99450, 99320, 99270, 99200, 99160, 
    99120, 99070, 99030, 99000, 98950, 98890, 98820, 98750, 98680, 98540, 
    98410, 98480, 98470, 98450, 98480, 98500, 98530, 98560, 98600, 98610, 
    98610, 98580, 98590, 98570, 98570, 98520, 98510, 98520, 98540, 98580, 
    98610, 98650, 98740, 98830, 98930, 99030, 99100, 99140, 99180, 99220, 
    99260, 99260, 99260, 99260, 99240, 99250, 99230, 99320, 99330, 99330, 
    99280, 99250, 99350, 99480, 99590, 99670, 99700, 99770, 99810, 99810, 
    99830, 99850, 99850, 99880, 99910, 99920, 99920, 99940, 99940, 99960, 
    99960, 100010, 100050, 100040, 100040, 100050, 100040, 100040, 100050, 
    100010, 100000, 100020, 100030, 100020, 100030, 100010, 99980, 99960, 
    99900, 99870, 99850, 99830, 99780, 99730, 99730, 99720, 99680, 99670, 
    99650, 99620, 99590, 99540, 99480, 99440, 99400, 99330, 99270, 99230, 
    99210, 99180, 99160, 99140, 99110, 99110, 99090, 99060, 99090, 99150, 
    99160, 99200, 99260, 99310, 99340, 99360, 99390, 99420, 99430, 99450, 
    99470, 99460, 99500, 99530, 99560, 99580, 99590, 99600, 99620, 99610, 
    99610, 99600, 99590, 99620, 99640, 99660, 99690, 99710, 99700, 99710, 
    99690, 99720, 99720, 99730, 99730, 99760, 99730, 99700, 99680, 99710, 
    99730, 99720, 99740, 99730, 99700, 99650, 99650, 99610, 99610, 99590, 
    99590, 99580, 99500, 99410, 99380, 99410, 99350, 99300, 99260, 99250, 
    99260, 99260, 99290, 99340, 99340, 99340, 99400, 99430, 99510, 99520, 
    99610, 99670, 99730, 99790, 99870, 99960, 100040, 100080, 100130, 100180, 
    100220, 100260, 100290, 100290, 100340, 100320, 100380, 100450, 100520, 
    100520, 100510, 100530, 100570, 100650, 100720, 100750, 100770, 100790, 
    100820, 100840, 100850, 100870, 100880, 100910, 100910, 100910, 100900, 
    100900, 100910, 100910, 100900, 100900, 100910, 100930, 100940, 100950, 
    100930, 100950, 100930, 100930, 100910, 100910, 100870, 100860, 100820, 
    100810, 100790, 100770, 100760, 100700, 100640, 100570, 100510, 100450, 
    100400, 100350, 100270, 100160, 100080, 99990, 99890, 99780, 99690, 
    99590, 99600, 99380, 99280, 99200, 99110, 98990, 98870, 98820, 98810, 
    98800, 98800, 98780, 98780, 98760, 98740, 98720, 98650, 98580, 98460, 
    98350, 98340, 98400, 98390, 98300, 98250, 98200, 98230, 98250, 98290, 
    98300, 98290, 98330, 98300, 98270, 98240, 98230, 98080, 98080, 98260, 
    98360, 98340, 98370, 98380, 98430, 98420, 98440, 98430, 98470, 98480, 
    98490, 98570, 98540, 98600, 98560, 98550, 98610, 98490, 98580, 98660, 
    98630, 98640, 98640, 98640, 98640, 98740, 98870, 98860, 98830, 98850, 
    98750, 98680, 98670, 98670, 98680, 98690, 98710, 98740, 98750, 98730, 
    98790, 98790, 98770, 98680, 98690, 98780, 98890, 99000, 99070, 99060, 
    99090, 99150, 99210, 99250, 99290, 99350, 99440, 99480, 99520, 99590, 
    99600, 99630, 99670, 99720, 99760, 99830, 99890, 99950, 100000, 100080, 
    100170, 100250, 100290, 100340, 100410, 100490, 100560, 100590, 100650, 
    100690, 100720, 100760, 100800, 100840, 100900, 100920, 100970, 100960, 
    100950, 100970, 100970, 100960, 100940, 100950, 100960, 100960, 100960, 
    100950, 100930, 100900, 100880, 100840, 100810, 100780, 100790, 100780, 
    100760, 100730, 100710, 100700, 100670, 100630, 100590, 100560, 100570, 
    100530, 100490, 100460, 100420, 100410, 100380, 100330, 100290, 100280, 
    100220, 100180, 100110, 100000, 99970, 99920, 99860, 99770, 99670, 99540, 
    99460, 99380, 99250, 99190, 99110, 99070, 99000, 98990, 98940, 98910, 
    98880, 98880, 98900, 98890, 98890, 98910, 98920, 98940, 99010, 99080, 
    99180, 99240, 99300, 99330, 99330, 99330, 99340, 99340, 99340, 99370, 
    99390, 99390, 99410, 99410, 99410, 99410, 99410, 99430, 99440, 99430, 
    99440, 99430, 99420, 99430, 99470, 99490, 99500, 99510, 99510, 99500, 
    99520, 99530, 99540, 99560, 99520, 99540, 99540, 99520, 99500, 99480, 
    99480, 99500, 99450, 99440, 99420, 99380, 99340, 99300, 99310, 99340, 
    99340, 99340, 99290, 99220, 99220, 99190, 99170, 99170, 99140, 99160, 
    99170, 99200, 99230, 99250, 99270, 99280, 99320, 99350, 99380, 99400, 
    99410, 99440, 99480, 99530, 99540, 99520, 99590, 99620, 99630, 99660, 
    99680, 99740, 99750, 99780, 99850, 99900, 99900, 99950, 99900, 99890, 
    99920, 99890, 99810, 99830, 99810, 99820, 99850, 99890, 99950, 100000, 
    100010, 100140, 100180, 100300, 100410, 100460, 100510, 100570, 100610, 
    100660, 100730, 100810, 100850, 100920, 100970, 101060, 101120, 101210, 
    101320, 101420, 101470, 101450, 101460, 101560, 101550, 101590, 101660, 
    101780, 101870, 101920, 101900, 101940, 101970, 102020, 102100, 102110, 
    102130, 102080, 102170, 102180, 102190, 102180, 102170, 102180, 102200, 
    102220, 102180, 102170, 102180, 102170, 102150, 102130, 102110, 102070, 
    101990, 101900, 101930, 101840, 101720, 101760, 101700, 101630, 101480, 
    101390, 101380, 101240, 101200, 101170, 101140, 101080, 101030, 100980, 
    100820, 100720, 100720, 100700, 100560, 100500, 100410, 100440, 100380, 
    100280, 100120, 100030, 100010, 99920, 99830, 99760, 99760, 99710, 99670, 
    99690, 99690, 99570, 99470, 99430, 99320, 99260, 99210, 99170, 99120, 
    98990, 98920, 98860, 98810, 98780, 98750, 98640, 98600, 98430, 98490, 
    98450, 98470, 98390, 98340, 98270, 98100, 98070, 98100, 98080, 98070, 
    98010, 97920, 97820, 97760, 97720, 97670, 97620, 97560, 97510, 97420, 
    97380, 97380, 97330, 97230, 97140, 97230, 97160, 97140, 97070, 97060, 
    97070, 97010, 96990, 96880, 96880, 96910, 96910, 96950, 96930, 96940, 
    96950, 96970, 97080, 97020, 97060, 97110, 97160, 97230, 97310, 97400, 
    97510, 97570, 97680, 97790, 97900, 98010, 98110, 98150, 98250, 98300, 
    98370, 98440, 98500, 98570, 98620, 98680, 98750, 98820, 98890, 99030, 
    99040, 99110, 99140, 99200, 99230, 99260, 99310, 99370, 99420, 99440, 
    99460, 99540, 99550, 99500, 99510, 99460, 99450, 99400, 99350, 99260, 
    99120, 98980, 98800, 98700, 98630, 98560, 98500, 98440, 98390, 98330, 
    98290, 98260, 98270, 98230, 98180, 98140, 98080, 98010, 97940, 97870, 
    97800, 97720, 97660, 97610, 97600, 97600, 97600, 97650, 97650, 97690, 
    97680, 97660, 97670, 97720, 97620, 97630, 97620, 97610, 97560, 97530, 
    97510, 97460, 97410, 97380, 97360, 97350, 97370, 97380, 97410, 97460, 
    97550, 97580, 97620, 97690, 97730, 97750, 97800, 97810, 97910, 97940, 
    98000, 98010, 98070, 98040, 98000, 97980, 97930, 97900, 97890, 97910, 
    97900, 97930, 97960, 97980, 97990, 98040, 98110, 98190, 98280, 98390, 
    98500, 98590, 98650, 98840, 99040, 99220, 99390, 99560, 99710, 99830, 
    99920, 100060, 100200, 100300, 100410, 100520, 100640, 100790, 100840, 
    100880, 100980, 101070, 101060, 101050, 101030, 100990, 100960, 100930, 
    100880, 100870, 100920, 100970, 101020, 101080, 101160, 101250, 101300, 
    101370, 101420, 101480, 101540, 101590, 101630, 101660, 101700, 101750, 
    101730, 101720, 101700, 101660, 101610, 101560, 101510, 101440, 101360, 
    101310, 101280, 101230, 101180, 101150, 101110, 101060, 101020, 100980, 
    100970, 100890, 100810, 100720, 100570, 100520, 100490, 100480, 100480, 
    100420, 100460, 100350, 100240, 100240, 100270, 100300, 100330, 100320, 
    100380, 100470, 100590, 100590, 100630, 100640, 100640, 100650, 100670, 
    100670, 100660, 100650, 100630, 100650, 100440, 100370, 100120, 100090, 
    100110, 100080, 100050, 100460, 100590, 100670, 100750, 100820, 100890, 
    100960, 101000, 101080, 101130, 101120, 101090, 101090, 101040, 100960, 
    100890, 100820, 100810, 100660, 100520, 100560, 100540, 100570, 100610, 
    100630, 100650, 100690, 100760, 100880, 100870, 100860, 100860, 100880, 
    100900, 100880, 100820, 100760, 100700, 100610, 100540, 100470, 100540, 
    100700, 100780, 101070, 101250, 101430, 101620, 101810, 101950, 102040, 
    102110, 102160, 102180, 102170, 102140, 102140, 102100, 102010, 101940, 
    101870, 101780, 101690, 101620, 101560, 101500, 101430, 101370, 101330, 
    101310, 101310, 101310, 101310, 101300, 101300, 101300, 101310, 101300, 
    101270, 101260, 101250, 101240, 101210, 101200, 101180, 101170, 101200, 
    101240, 101280, 101350, 101410, 101510, 101590, 101620, 101710, 101770, 
    101830, 101890, 101950, 102000, 102040, 102090, 102120, 102160, 102200, 
    102220, 102240, 102250, 102240, 102230, 102210, 102190, 102150, 102130, 
    102120, 102160, 102170, 102100, 102090, 102090, 102060, 102050, 102030, 
    102020, 101970, 101960, 101950, 101940, 101920, 101950, 101940, 101930, 
    101920, 101930, 101900, 101930, 101950, 101950, 101980, 102020, 102030, 
    102080, 102070, 102140, 102170, 102220, 102280, 102320, 102320, 102350, 
    102370, 102400, 102430, 102460, 102470, 102460, 102460, 102450, 102420, 
    102420, 102390, 102350, 102330, 102310, 102290, 102270, 102280, 102290, 
    102290, 102290, 102330, 102330, 102320, 102310, 102300, 102310, 102330, 
    102330, 102330, 102350, 102370, 102370, 102360, 102370, 102360, 102350, 
    102380, 102380, 102390, 102400, 102410, 102420, 102430, 102440, 102410, 
    102450, 102460, 102440, 102440, 102460, 102440, 102450, 102450, 102450, 
    102420, 102400, 102400, 102410, 102420, 102430, 102420, 102420, 102420, 
    102410, 102430, 102410, 102390, 102410, 102410, 102390, 102390, 102370, 
    102360, 102370, 102390, 102410, 102460, 102460, 102480, 102490, 102510, 
    102530, 102550, 102550, 102560, 102590, 102630, 102670, 102710, 102740, 
    102770, 102800, 102830, 102850, 102880, 102910, 102920, 102970, 103030, 
    103080, 103110, 103150, 103180, 103230, 103250, 103270, 103310, 103330, 
    103340, 103380, 103420, 103440, 103470, 103490, 103480, 103490, 103500, 
    103510, 103490, 103480, 103480, 103450, 103450, 103420, 103370, 103350, 
    103300, 103230, 103200, 103160, 103090, 102990, 102910, 102760, 102640, 
    102550, 102450, 102330, 102190, 102040, 101940, 101820, 101720, 101640, 
    101580, 101540, 101530, 101530, 101530, 101510, 101480, 101440, 101390, 
    101370, 101310, 101260, 101210, 101130, 101080, 101010, 100970, 100910, 
    100900, 100900, 100900, 100900, 100870, 100870, 100840, 100810, 100810, 
    100850, 100910, 100920, 100900, 100900, 100920, 100940, 100990, 101010, 
    101030, 101060, 101070, 101090, 101140, 101150, 101120, 101030, 101010, 
    101050, 101140, 101230, 101310, 101430, 101530, 101630, 101730, 101810, 
    101850, 101880, 101940, 101990, 102030, 102060, 102080, 102100, 102140, 
    102170, 102180, 102200, 102240, 102240, 102240, 102180, 102230, 102260, 
    102280, 102340, 102370, 102390, 102420, 102460, 102450, 102450, 102490, 
    102500, 102520, 102540, 102540, 102530, 102500, 102490, 102480, 102460, 
    102430, 102400, 102400, 102420, 102420, 102380, 102380, 102340, 102230, 
    102280, 102310, 102250, 102230, 102190, 102180, 102110, 102070, 102080, 
    102080, 102080, 102070, 102050, 102000, 102060, 102040, 102020, 101930, 
    101910, 101900, 101880, 101840, 101810, 101790, 101780, 101810, 101840, 
    101870, 101870, 101850, 101860, 101860, 101870, 101860, 101830, 101830, 
    101840, 101840, 101830, 101790, 101780, 101750, 101720, 101700, 101680, 
    101660, 101640, 101620, 101600, 101570, 101540, 101490, 101440, 101400, 
    101370, 101330, 101290, 101250, 101230, 101180, 101160, 101120, 101090, 
    101050, 101030, 100980, 100950, 100910, 100890, 100870, 100840, 100810, 
    100800, 100810, 100800, 100780, 100750, 100720, 100710, 100690, 100660, 
    100650, 100640, 100640, 100640, 100640, 100640, 100660, 100650, 100670, 
    100680, 100660, 100680, 100670, 100650, 100650, 100660, 100660, 100640, 
    100570, 100480, 100410, 100320, 100320, 100350, 100360, 100370, 100360, 
    100340, 100360, 100350, 100320, 100280, 100250, 100200, 100190, 100150, 
    100110, 100070, 100020, 99990, 99960, 99950, 99950, 99970, 100000, 
    100030, 100070, 100120, 100160, 100190, 100210, 100270, 100310, 100310, 
    100320, 100320, 100280, 100280, 100280, 100290, 100300, 100280, 100360, 
    100420, 100490, 100510, 100560, 100650, 100670, 100720, 100740, 100820, 
    100840, 100840, 100880, 100950, 100990, 101000, 101010, 101030, 101070, 
    101080, 101100, 101130, 101130, 101160, 101200, 101210, 101260, 101270, 
    101300, 101310, 101300, 101340, 101370, 101390, 101400, 101450, 101470, 
    101510, 101560, 101620, 101600, 101570, 101600, 101620, 101580, 101600, 
    101630, 101630, 101620, 101670, 101680, 101680, 101750, 101740, 101740, 
    101780, 101780, 101800, 101840, 101840, 101840, 101870, 101860, 101860, 
    101860, 101820, 101770, 101730, 101680, 101630, 101580, 101500, 101480, 
    101420, 101370, 101320, 101290, 101250, 101190, 101140, 101070, 100980, 
    100890, 100790, 100700, 100640, 100530, 100460, 100390, 100260, 100160, 
    100020, 99900, 99760, 99640, 99620, 99580, 99530, 99490, 99460, 99420, 
    99390, 99340, 99380, 99340, 99290, 99240, 99230, 99190, 99200, 99200, 
    99170, 99150, 99140, 99120, 99130, 99130, 99080, 99030, 98990, 98960, 
    98960, 98980, 98970, 98920, 98880, 98790, 98790, 98760, 98650, 98590, 
    98540, 98520, 98370, 98470, 98290, 98160, 98020, 97980, 97920, 97920, 
    97920, 97900, 97930, 97980, 98010, 98080, 98100, 98110, 98180, 98230, 
    98290, 98330, 98390, 98390, 98410, 98430, 98490, 98600, 98630, 98680, 
    98690, 98680, 98720, 98780, 98820, 98870, 98950, 98990, 99050, 99030, 
    99000, 99000, 99030, 98980, 98970, 99000, 99000, 99090, 99180, 99200, 
    99240, 99280, 99290, 99230, 99170, 99130, 99110, 99050, 99000, 99020, 
    99000, 99000, 99060, 98980, 98960, 99020, 99090, 99140, 99210, 99200, 
    99240, 99240, 99250, 99270, 99300, 99250, 99200, 99320, 99470, 99530, 
    99500, 99430, 99400, 99360, 99390, 99500, 99540, 99640, 99660, 99680, 
    99710, 99730, 99760, 99790, 99800, 99800, 99820, 99750, 99770, 99810, 
    99810, 99790, 99830, 99890, 99880, 99920, 99900, 99940, 99610, 99570, 
    99680, 99870, 100090, 100120, 100140, 100180, 100180, 100200, 100200, 
    100180, 100160, 100180, 100210, 100260, 100330, 100380, 100390, 100410, 
    100380, 100440, 100510, 100580, 100540, 100630, 100680, 100700, 100730, 
    100700, 100560, 100630, 100750, 100760, 100800, 100730, 100700, 100680, 
    101080, 101390, 101430, 101450, 101470, 101470, 101410, 101460, 101390, 
    101530, 101550, 101490, 101470, 101500, 101550, 101510, 101460, 101440, 
    101380, 101350, 101320, 101220, 101240, 101210, 101180, 101170, 101140, 
    101100, 101070, 101020, 100970, 100940, 100870, 100810, 100740, 100760, 
    100760, 100750, 100730, 100720, 100700, 100670, 100690, 100680, 100700, 
    100700, 100690, 100660, 100660, 100650, 100620, 100620, 100610, 100590, 
    100580, 100540, 100500, 100490, 100470, 100470, 100480, 100460, 100480, 
    100500, 100470, 100470, 100450, 100440, 100420, 100420, 100400, 100380, 
    100390, 100400, 100420, 100440, 100460, 100480, 100480, 100490, 100480, 
    100500, 100500, 100510, 100540, 100570, 100590, 100600, 100610, 100620, 
    100620, 100590, 100580, 100590, 100600, 100610, 100630, 100640, 100630, 
    100600, 100580, 100560, 100550, 100500, 100470, 100460, 100420, 100380, 
    100360, 100330, 100290, 100200, 100150, 100030, 99980, 99930, 99850, 
    99750, 99700, 99550, 99470, 99380, 99160, 99070, 99030, 98970, 98810, 
    98840, 98780, 98760, 98700, 98640, 98570, 98470, 98340, 98220, 98190, 
    98110, 97990, 97880, 97790, 97730, 97680, 97680, 97630, 97600, 97560, 
    97530, 97480, 97510, 97490, 97450, 97450, 97400, 97420, 97440, 97470, 
    97500, 97550, 97590, 97610, 97640, 97720, 97800, 97890, 97970, 98050, 
    98160, 98240, 98320, 98390, 98460, 98510, 98570, 98600, 98630, 98650, 
    98670, 98710, 98780, 98840, 98880, 98950, 98980, 99010, 99030, 99070, 
    99100, 99150, 99190, 99240, 99280, 99320, 99370, 99430, 99480, 99520, 
    99560, 99620, 99650, 99680, 99730, 99770, 99830, 99890, 99950, 99970, 
    100000, 100030, 100050, 100080, 100110, 100140, 100140, 100140, 100150, 
    100180, 100200, 100200, 100220, 100220, 100210, 100200, 100190, 100190, 
    100180, 100180, 100200, 100210, 100230, 100230, 100210, 100220, 100240, 
    100300, 100350, 100390, 100480, 100520, 100580, 100630, 100700, 100770, 
    100840, 100900, 100940, 100960, 100990, 101040, 101070, 101110, 101150, 
    101180, 101280, 101290, 101330, 101390, 101450, 101500, 101540, 101570, 
    101620, 101660, 101710, 101750, 101800, 101800, 101800, 101770, 101770, 
    101780, 101780, 101740, 101700, 101680, 101670, 101690, 101690, 101700, 
    101680, 101620, 101610, 101600, 101570, 101540, 101520, 101520, 101530, 
    101550, 101520, 101460, 101460, 101450, 101430, 101400, 101390, 101350, 
    101360, 101340, 101330, 101290, 101260, 101250, 101230, 101210, 101230, 
    101220, 101200, 101160, 101150, 101130, 101150, 101150, 101130, 101130, 
    101080, 101060, 101080, 101080, 101060, 101020, 101020, 100980, 100930, 
    100880, 100870, 100890, 100880, 100810, 100760, 100720, 100680, 100630, 
    100570, 100490, 100430, 100400, 100370, 100360, 100360, 100370, 100410, 
    100430, 100460, 100500, 100530, 100590, 100620, 100660, 100680, 100690, 
    100690, 100700, 100700, 100710, 100690, 100690, 100650, 100680, 100590, 
    100620, 100650, 100600, 100570, 100500, 100460, 100430, 100380, 100330, 
    100290, 100190, 100120, 100080, 100010, 99880, 99770, 99630, 99540, 
    99440, 99390, 99340, 99250, 99200, 99170, 99170, 99220, 99220, 99220, 
    99220, 99240, 99320, 99290, 99290, 99290, 99290, 99290, 99310, 99320, 
    99340, 99380, 99390, 99440, 99440, 99450, 99430, 99460, 99480, 99520, 
    99570, 99630, 99690, 99720, 99730, 99760, 99820, 99890, 99950, 100030, 
    100080, 100170, 100250, 100330, 100410, 100460, 100510, 100540, 100550, 
    100570, 100550, 100520, 100530, 100500, 100480, 100430, 100380, 100310, 
    100270, 100230, 100180, 100120, 100100, 100110, 100140, 100160, 100190, 
    100250, 100300, 100310, 100360, 100370, 100410, 100440, 100490, 100540, 
    100580, 100630, 100680, 100720, 100760, 100780, 100820, 100860, 100900, 
    100930, 100960, 100980, 101000, 101000, 101010, 101070, 101090, 101060, 
    101100, 101100, 101100, 101140, 101140, 101160, 101180, 101250, 101320, 
    101380, 101440, 101470, 101480, 101530, 101560, 101580, 101630, 101640, 
    101650, 101660, 101680, 101700, 101700, 101690, 101680, 101670, 101650, 
    101650, 101650, 101640, 101640, 101620, 101570, 101590, 101620, 101630, 
    101600, 101590, 101580, 101580, 101540, 101530, 101530, 101560, 101550, 
    101570, 101550, 101550, 101530, 101530, 101530, 101530, 101550, 101560, 
    101580, 101560, 101570, 101550, 101560, 101560, 101530, 101530, 101520, 
    101520, 101500, 101520, 101530, 101540, 101540, 101550, 101560, 101560, 
    101540, 101520, 101510, 101490, 101480, 101460, 101450, 101440, 101420, 
    101410, 101390, 101360, 101330, 101290, 101250, 101240, 101210, 101180, 
    101160, 101130, 101120, 101100, 101080, 101050, 101040, 101000, 100980, 
    100950, 100920, 100880, 100880, 100870, 100850, 100840, 100810, 100820, 
    100800, 100770, 100750, 100760, 100760, 100740, 100720, 100730, 100740, 
    100750, 100770, 100770, 100760, 100770, 100780, 100770, 100760, 100760, 
    100740, 100740, 100720, 100730, 100750, 100720, 100720, 100710, 100680, 
    100680, 100690, 100710, 100720, 100720, 100750, 100770, 100760, 100780, 
    100760, 100760, 100750, 100760, 100760, 100730, 100720, 100740, 100690, 
    100680, 100690, 100670, 100660, 100640, 100630, 100620, 100620, 100640, 
    100650, 100660, 100640, 100660, 100640, 100610, 100590, 100550, 100490, 
    100410, 100430, 100440, 100390, 100430, 100470, 100480, 100430, 100450, 
    100510, 100500, 100490, 100470, 100420, 100360, 100230, 100190, 100240, 
    100290, 100290, 100300, 100320, 100320, 100320, 100380, 100440, 100500, 
    100530, 100610, 100670, 100710, 100730, 100770, 100770, 100770, 100740, 
    100770, 100760, 100750, 100730, 100740, 100730, 100730, 100750, 100800, 
    100800, 100780, 100780, 100780, 100770, 100750, 100710, 100710, 100690, 
    100710, 100760, 100780, 100820, 100830, 100830, 100830, 100820, 100820, 
    100810, 100800, 100800, 100770, 100810, 100800, 100770, 100740, 100710, 
    100660, 100640, 100610, 100560, 100500, 100450, 100420, 100370, 100290, 
    100200, 100150, 100070, 100020, 99990, 99980, 99970, 99970, 100030, 
    100100, 100140, 100170, 100180, 100120, 100130, 100090, 100090, 100070, 
    100070, 100090, 100130, 100190, 100240, 100290, 100350, 100390, 100450, 
    100470, 100500, 100550, 100590, 100580, 100610, 100650, 100690, 100690, 
    100700, 100700, 100690, 100700, 100710, 100720, 100740, 100750, 100770, 
    100810, 100850, 100880, 100950, 100990, 101020, 101060, 101100, 101140, 
    101160, 101170, 101210, 101210, 101230, 101230, 101240, 101240, 101230, 
    101230, 101230, 101250, 101250, 101280, 101280, 101290, 101260, 101280, 
    101300, 101270, 101260, 101260, 101300, 101330, 101360, 101370, 101390, 
    101450, 101470, 101510, 101510, 101530, 101540, 101590, 101610, 101640, 
    101690, 101700, 101660, 101660, 101680, 101760, 101800, 101810, 101810, 
    101820, 101830, 101840, 101850, 101870, 101870, 101880, 101860, 101840, 
    101840, 101790, 101710, 101650, 101600, 101570, 101550, 101520, 101480, 
    101430, 101380, 101340, 101310, 101290, 101230, 101180, 101180, 101160, 
    101130, 101100, 101110, 101110, 101100, 101110, 101130, 101160, 101150, 
    101160, 101150, 101170, 101200, 101210, 101230, 101250, 101260, 101250, 
    101280, 101290, 101290, 101330, 101320, 101340, 101350, 101340, 101330, 
    101290, 101280, 101240, 101220, 101190, 101160, 101090, 101040, 101000, 
    100930, 100900, 100840, 100810, 100770, 100720, 100710, 100670, 100650, 
    100580, 100510, 100450, 100400, 100450, 100420, 100430, 100450, 100470, 
    100500, 100480, 100490, 100540, 100520, 100560, 100530, 100540, 100550, 
    100570, 100530, 100500, 100480, 100430, 100360, 100340, 100280, 100220, 
    100150, 100070, 99960, 99880, 99710, 99520, 99370, 99220, 99070, 98980, 
    98930, 98940, 98920, 98940, 98970, 99000, 98990, 99040, 99040, 99140, 
    99180, 99340, 99560, 99630, 99760, 99910, 100050, 100190, 100220, 100250, 
    100340, 100300, 100240, 100190, 100100, 100000, 99890, 99680, 99470, 
    99220, 98990, 98810, 98580, 98450, 98360, 98360, 98360, 98470, 98530, 
    98620, 98780, 98900, 99000, 99140, 99250, 99410, 99550, 99590, 99680, 
    99740, 99800, 99880, 99960, 100000, 100050, 100010, 100070, 100110, 
    100150, 100160, 100120, 100120, 100120, 100120, 100120, 100100, 100120, 
    100100, 100080, 100070, 100070, 100060, 100100, 100120, 100120, 100150, 
    100220, 100260, 100310, 100370, 100420, 100470, 100540, 100600, 100640, 
    100680, 100730, 100790, 100830, 100850, 100900, 100930, 100970, 101010, 
    101060, 101060, 101030, 101020, 101050, 100970, 100910, 100930, 100870, 
    100800, 100780, 100780, 100750, 100830, 100840, 100840, 100830, 100860, 
    100850, 100890, 100900, 100930, 100930, 100900, 100910, 100940, 100910, 
    100850, 100850, 100840, 100890, 100900, 100890, 100840, 100810, 100780, 
    100750, 100710, 100680, 100660, 100610, 100600, 100590, 100620, 100660, 
    100660, 100650, 100650, 100680, 100660, 100680, 100690, 100720, 100740, 
    100750, 100780, 100810, 100830, 100810, 100790, 100800, 100800, 100820, 
    100840, 100830, 100780, 100800, 100800, 100830, 100820, 100820, 100810, 
    100810, 100790, 100800, 100760, 100750, 100730, 100720, 100710, 100620, 
    100540, 100510, 100510, 100520, 100470, 100450, 100410, 100390, 100330, 
    100310, 100330, 100330, 100320, 100320, 100300, 100290, 100310, 100270, 
    100260, 100260, 100250, 100240, 100260, 100260, 100250, 100240, 100240, 
    100230, 100250, 100240, 100250, 100250, 100260, 100280, 100330, 100360, 
    100380, 100370, 100410, 100430, 100470, 100510, 100530, 100560, 100590, 
    100600, 100630, 100650, 100660, 100670, 100670, 100700, 100690, 100720, 
    100730, 100730, 100740, 100740, 100730, 100740, 100760, 100760, 100770, 
    100780, 100800, 100810, 100830, 100830, 100840, 100850, 100850, 100860, 
    100870, 100870, 100860, 100870, 100870, 100880, 100880, 100870, 100870, 
    100880, 100910, 100930, 100930, 100910, 100920, 100910, 100930, 100930, 
    100930, 100910, 100890, 100890, 100880, 100870, 100850, 100830, 100790, 
    100720, 100660, 100550, 100520, 100500, 100500, 100500, 100500, 100480, 
    100490, 100480, 100450, 100430, 100400, 100350, 100330, 100320, 100360, 
    100350, 100390, 100410, 100420, 100420, 100450, 100460, 100490, 100500, 
    100520, 100520, 100510, 100530, 100550, 100580, 100580, 100560, 100530, 
    100530, 100510, 100490, 100470, 100450, 100420, 100410, 100410, 100380, 
    100390, 100370, 100350, 100340, 100340, 100300, 100250, 100210, 100160, 
    100130, 100120, 100060, 99980, 99920, 99870, 99780, 99720, 99650, 99560, 
    99470, 99370, 99290, 99230, 99190, 99060, 98920, 98770, 98560, 98430, 
    98390, 98400, 98350, 98350, 98300, 98250, 98200, 98120, 98090, 98040, 
    98010, 97990, 98030, 98050, 98070, 97950, 97980, 98110, 98280, 98280, 
    98420, 98440, 98390, 98420, 98450, 98510, 98540, 98610, 98610, 98710, 
    98790, 98820, 98840, 98920, 99100, 99170, 99230, 99280, 99330, 99370, 
    99380, 99390, 99440, 99430, 99440, 99440, 99420, 99400, 99400, 99400, 
    99410, 99440, 99440, 99460, 99450, 99470, 99470, 99450, 99460, 99480, 
    99470, 99470, 99490, 99490, 99470, 99480, 99490, 99520, 99530, 99540, 
    99540, 99570, 99590, 99620, 99630, 99670, 99710, 99730, 99760, 99820, 
    99840, 99880, 99930, 99940, 99940, 99990, 100040, 100080, 100110, 100120, 
    100180, 100220, 100290, 100340, 100380, 100410, 100430, 100470, 100530, 
    100580, 100650, 100720, 100780, 100840, 100920, 100960, 101020, 101040, 
    101090, 101120, 101150, 101200, 101240, 101300, 101350, 101390, 101410, 
    101430, 101450, 101470, 101500, 101530, 101560, 101570, 101580, 101600, 
    101600, 101630, 101630, 101620, 101640, 101630, 101630, 101630, 101620, 
    101630, 101630, 101630, 101620, 101640, 101600, 101610, 101590, 101600, 
    101580, 101550, 101540, 101540, 101560, 101590, 101600, 101610, 101610, 
    101610, 101580, 101580, 101560, 101600, 101620, 101630, 101650, 101680, 
    101700, 101700, 101720, 101720, 101730, 101720, 101740, 101760, 101770, 
    101760, 101820, 101860, 101880, 101890, 101880, 101890, 101890, 101890, 
    101900, 101920, 101930, 101960, 101980, 102010, 102020, 102010, 101980, 
    101960, 101950, 101930, 101930, 101920, 101880, 101870, 101870, 101880, 
    101870, 101830, 101820, 101800, 101760, 101730, 101710, 101700, 101660, 
    101640, 101610, 101590, 101580, 101560, 101540, 101500, 101490, 101460, 
    101460, 101460, 101450, 101450, 101460, 101460, 101490, 101490, 101500, 
    101520, 101560, 101550, 101580, 101590, 101630, 101630, 101620, 101620, 
    101620, 101610, 101600, 101630, 101640, 101650, 101670, 101670, 101690, 
    101720, 101740, 101760, 101750, 101760, 101780, 101780, 101770, 101780, 
    101810, 101830, 101860, 101870, 101880, 101910, 101930, 101940, 101940, 
    101930, 101940, 101950, 101940, 101940, 101930, 101920, 101920, 101920, 
    101900, 101880, 101810, 101800, 101770, 101780, 101780, 101760, 101740, 
    101720, 101700, 101680, 101680, 101640, 101580, 101570, 101540, 101510, 
    101480, 101450, 101450, 101420, 101390, 101360, 101350, 101330, 101280, 
    101250, 101220, 101220, 101210, 101180, 101140, 101120, 101140, 101180, 
    101200, 101240, 101260, 101300, 101340, 101400, 101420, 101430, 101460, 
    101470, 101470, 101460, 101420, 101380, 101350, 101330, 101350, 101370, 
    101380, 101370, 101370, 101370, 101390, 101410, 101370, 101350, 101350, 
    101300, 101300, 101220, 101150, 101070, 101030, 101030, 100970, 100990, 
    100940, 100940, 100970, 101020, 101050, 101090, 101090, 101080, 101090, 
    101110, 101120, 101160, 101220, 101210, 101220, 101220, 101230, 101240, 
    101260, 101240, 101270, 101320, 101330, 101370, 101380, 101380, 101400, 
    101430, 101410, 101370, 101320, 101260, 101330, 101320, 101310, 101290, 
    101240, 101250, 101170, 101140, 101120, 101050, 100980, 100940, 100900, 
    100900, 100880, 100880, 100920, 100880, 100900, 100890, 100880, 100850, 
    100800, 100770, 100780, 100740, 100680, 100640, 100700, 100730, 100690, 
    100660, 100680, 100660, 100720, 100730, 100830, 100840, 100860, 100870, 
    100900, 100920, 100920, 100980, 100950, 100980, 100980, 100980, 101070, 
    101100, 101050, 101050, 101090, 101080, 101060, 101110, 101080, 101080, 
    101080, 101080, 101080, 101100, 101110, 101160, 101170, 101130, 101110, 
    101120, 101090, 101080, 101100, 101100, 101220, 101200, 101230, 101220, 
    101210, 101180, 101230, 101290, 101300, 101280, 101290, 101320, 101310, 
    101340, 101350, 101370, 101390, 101400, 101410, 101430, 101450, 101460, 
    101460, 101470, 101490, 101510, 101530, 101530, 101530, 101520, 101510, 
    101500, 101500, 101480, 101470, 101470, 101470, 101450, 101450, 101440, 
    101440, 101430, 101420, 101410, 101390, 101380, 101350, 101340, 101330, 
    101300, 101280, 101260, 101250, 101240, 101230, 101200, 101160, 101150, 
    101120, 101080, 101060, 101020, 100990, 100920, 100840, 100780, 100670, 
    100610, 100540, 100450, 100390, 100330, 100270, 100150, 100090, 100040, 
    99990, 99920, 99870, 99820, 99750, 99650, 99610, 99620, 99600, 99590, 
    99600, 99600, 99620, 99630, 99640, 99650, 99650, 99660, 99680, 99710, 
    99720, 99740, 99760, 99780, 99790, 99810, 99840, 99860, 99890, 99900, 
    99920, 99970, 100020, 100040, 100070, 100100, 100180, 100230, 100270, 
    100380, 100490, 100530, 100610, 100660, 100700, 100740, 100780, 100820, 
    100860, 100910, 100980, 101070, 101110, 101150, 101210, 101240, 101320, 
    101390, 101460, 101530, 101600, 101680, 101750, 101800, 101860, 101890, 
    101920, 101950, 101990, 102020, 102060, 102110, 102130, 102140, 102110, 
    102120, 102130, 102120, 102100, 102080, 102090, 102050, 102050, 102010, 
    101940, 101900, 101870, 101820, 101810, 101810, 101820, 101760, 101750, 
    101740, 101720, 101720, 101720, 101730, 101720, 101700, 101690, 101640, 
    101610, 101570, 101560, 101540, 101500, 101460, 101420, 101390, 101340, 
    101290, 101240, 101240, 101210, 101170, 101110, 101100, 101110, 101090, 
    101070, 101110, 101150, 101160, 101180, 101200, 101220, 101250, 101310, 
    101380, 101450, 101500, 101570, 101630, 101670, 101710, 101760, 101780, 
    101820, 101840, 101870, 101900, 101940, 101970, 101980, 101980, 101940, 
    101960, 102030, 102040, 102000, 102000, 102020, 102060, 102120, 102170, 
    102240, 102300, 102390, 102440, 102490, 102570, 102660, 102750, 102860, 
    103000, 103120, 103220, 103280, 103350, 103440, 103500, 103580, 103660, 
    103730, 103800, 103850, 103910, 103950, 103970, 104000, 104050, 104090, 
    104090, 104070, 104090, 104110, 104130, 104130, 104170, 104150, 104130, 
    104100, 104070, 104020, 104010, 103980, 103920, 103890, 103810, 103850, 
    103740, 103800, 103780, 103750, 103750, 103750, 103720, 103710, 103690, 
    103670, 103670, 103640, 103620, 103600, 103590, 103580, 103550, 103520, 
    103460, 103390, 103350, 103300, 103260, 103230, 103210, 103170, 103120, 
    103080, 103060, 103020, 102980, 102990, 102980, 102970, 102990, 103000, 
    103020, 103040, 103080, 103140, 103160, 103200, 103230, 103240, 103280, 
    103290, 103330, 103370, 103380, 103430, 103450, 103480, 103490, 103490, 
    103490, 103500, 103460, 103450, 103400, 103370, 103340, 103310, 103270, 
    103250, 103250, 103270, 103260, 103240, 103240, 103220, 103230, 103210, 
    103190, 103190, 103180, 103150, 103110, 103100, 103070, 103030, 102970, 
    102920, 102840, 102770, 102700, 102650, 102550, 102450, 102340, 102270, 
    102190, 102140, 102040, 101930, 101890, 101850, 101840, 101760, 101730, 
    101700, 101650, 101620, 101610, 101620, 101630, 101620, 101640, 101650, 
    101650, 101680, 101680, 101720, 101710, 101730, 101800, 101840, 101850, 
    101890, 101890, 101950, 101960, 102020, 102080, 102110, 102130, 102180, 
    102210, 102250, 102270, 102310, 102330, 102360, 102390, 102430, 102480, 
    102510, 102540, 102560, 102590, 102600, 102610, 102620, 102640, 102660, 
    102690, 102730, 102750, 102760, 102790, 102810, 102830, 102830, 102840, 
    102840, 102850, 102850, 102850, 102870, 102890, 102890, 102900, 102910, 
    102890, 102890, 102880, 102890, 102870, 102860, 102870, 102880, 102890, 
    102900, 102900, 102900, 102900, 102900, 102900, 102860, 102870, 102890, 
    102850, 102850, 102860, 102860, 102880, 102860, 102860, 102850, 102850, 
    102850, 102860, 102870, 102880, 102900, 102910, 102920, 102920, 102940, 
    102930, 102920, 102910, 102910, 102900, 102880, 102860, 102860, 102850, 
    102840, 102850, 102850, 102810, 102780, 102750, 102730, 102710, 102690, 
    102680, 102690, 102690, 102690, 102660, 102620, 102610, 102610, 102560, 
    102560, 102550, 102520, 102530, 102480, 102480, 102490, 102470, 102430, 
    102400, 102380, 102380, 102380, 102340, 102300, 102290, 102280, 102300, 
    102340, 102330, 102320, 102310, 102220, 102190, 102180, 102170, 102150, 
    102170, 102130, 102120, 102100, 102060, 102040, 102010, 101990, 101970, 
    101960, 101980, 101980, 102040, 102070, 102100, 102140, 102050, 102070, 
    102090, 102100, 102100, 102100, 102180, 102160, 102100, 102120, 102180, 
    102210, 102190, 102190, 102180, 102180, 102180, 102180, 102200, 102210, 
    102210, 102230, 102200, 102230, 102230, 102240, 102240, 102240, 102230, 
    102220, 102210, 102170, 102160, 102140, 102120, 102110, 102120, 102120, 
    102110, 102100, 102090, 102100, 102100, 102090, 102100, 102110, 102130, 
    102130, 102160, 102150, 102150, 102170, 102150, 102160, 102150, 102140, 
    102150, 102150, 102150, 102160, 102170, 102170, 102170, 102180, 102180, 
    102170, 102180, 102200, 102190, 102190, 102180, 102200, 102210, 102220, 
    102190, 102140, 102140, 102130, 102090, 102030, 102030, 102020, 101970, 
    101930, 101890, 101820, 101810, 101780, 101750, 101690, 101640, 101650, 
    101640, 101670, 101690, 101710, 101720, 101780, 101810, 101840, 101890, 
    101950, 101970, 102000, 102000, 102000, 102030, 102060, 102080, 102110, 
    102110, 102130, 102160, 102170, 102160, 102140, 102170, 102190, 102190, 
    102170, 102170, 102160, 102160, 102150, 102130, 102110, 102110, 102080, 
    102080, 102040, 102030, 101990, 101950, 101930, 101920, 101870, 101860, 
    101820, 101770, 101740, 101690, 101660, 101630, 101620, 101590, 101540, 
    101530, 101460, 101400, 101350, 101290, 101230, 101130, 101060, 100980, 
    100940, 100860, 100740, 100610, 100590, 100550, 100540, 100550, 100530, 
    100540, 100500, 100510, 100540, 100570, 100570, 100570, 100570, 100540, 
    100550, 100520, 100530, 100550, 100540, 100580, 100590, 100570, 100520, 
    100500, 100510, 100450, 100410, 100380, 100360, 100320, 100220, 100190, 
    100260, 100170, 100130, 100090, 100140, 100120, 100150, 100200, 100210, 
    100190, 100170, 100200, 100210, 100210, 100220, 100210, 100230, 100220, 
    100240, 100260, 100280, 100300, 100330, 100330, 100360, 100380, 100360, 
    100350, 100350, 100360, 100360, 100360, 100350, 100340, 100330, 100310, 
    100300, 100280, 100270, 100250, 100210, 100180, 100160, 100120, 100090, 
    100090, 100070, 100060, 100050, 100020, 99990, 99970, 99940, 99920, 
    99900, 99870, 99850, 99830, 99810, 99800, 99780, 99770, 99760, 99750, 
    99740, 99730, 99740, 99730, 99740, 99750, 99760, 99800, 99820, 99840, 
    99860, 99880, 99910, 99930, 99960, 99970, 100010, 100040, 100070, 100100, 
    100150, 100190, 100210, 100230, 100260, 100270, 100280, 100330, 100340, 
    100380, 100410, 100420, 100440, 100470, 100460, 100470, 100490, 100520, 
    100550, 100580, 100570, 100570, 100570, 100560, 100620, 100700, 100730, 
    100780, 100880, 100930, 101020, 101120, 101140, 101220, 101300, 101360, 
    101420, 101490, 101530, 101560, 101590, 101610, 101650, 101640, 101650, 
    101670, 101680, 101700, 101730, 101760, 101800, 101840, 101860, 101880, 
    101900, 101930, 101960, 101990, 102020, 102040, 102080, 102110, 102110, 
    102120, 102130, 102120, 102120, 102110, 102110, 102090, 102100, 102090, 
    102080, 102090, 102060, 102030, 102010, 101970, 101940, 101910, 101910, 
    101900, 101900, 101900, 101900, 101890, 101880, 101920, 101890, 101870, 
    101860, 101850, 101830, 101870, 101900, 101860, 101840, 101790, 101740, 
    101740, 101750, 101750, 101700, 101800, 101810, 101810, 101770, 101750, 
    101720, 101610, 101560, 101470, 101540, 101490, 101480, 101530, 101590, 
    101550, 101560, 101600, 101650, 101620, 101610, 101590, 101620, 101670, 
    101640, 101640, 101640, 101590, 101600, 101580, 101570, 101570, 101560, 
    101570, 101580, 101580, 101610, 101600, 101630, 101640, 101650, 101620, 
    101620, 101620, 101620, 101650, 101660, 101690, 101680, 101690, 101700, 
    101740, 101750, 101750, 101770, 101780, 101800, 101810, 101810, 101830, 
    101810, 101800, 101810, 101790, 101790, 101810, 101800, 101790, 101760, 
    101760, 101760, 101760, 101700, 101730, 101700, 101660, 101590, 101570, 
    101520, 101420, 101390, 101290, 101230, 101120, 101010, 100930, 100830, 
    100760, 100730, 100680, 100720, 100640, 100590, 100550, 100520, 100460, 
    100450, 100380, 100370, 100360, 100400, 100450, 100480, 100530, 100580, 
    100640, 100700, 100780, 100860, 100990, 101100, 101190, 101310, 101430, 
    101600, 101770, 101950, 102080, 102210, 102340, 102440, 102540, 102650, 
    102750, 102860, 102930, 102990, 103090, 103130, 103180, 103250, 103300, 
    103310, 103330, 103360, 103370, 103370, 103380, 103390, 103400, 103370, 
    103370, 103350, 103320, 103300, 103260, 103230, 103210, 103190, 103180, 
    103180, 103140, 103130, 103110, 103060, 103010, 102960, 102910, 102870, 
    102820, 102780, 102730, 102670, 102630, 102600, 102550, 102480, 102420, 
    102360, 102320, 102250, 102190, 102120, 102070, 102020, 101980, 101940, 
    101890, 101840, 101780, 101720, 101700, 101650, 101590, 101580, 101550, 
    101540, 101490, 101470, 101450, 101430, 101420, 101420, 101510, 101560, 
    101650, 101700, 101760, 101880, 101950, 102010, 102070, 102070, 102100, 
    102120, 102130, 102120, 102100, 102100, 102090, 102080, 102050, 102030, 
    102000, 101930, 101860, 101780, 101730, 101660, 101610, 101540, 101490, 
    101420, 101360, 101320, 101260, 101230, 101190, 101120, 101080, 101030, 
    100990, 100930, 100870, 100800, 100790, 100830, 100800, 100820, 100820, 
    100810, 100810, 100860, 100880, 100920, 100930, 100940, 100960, 100970, 
    100990, 100990, 101000, 100970, 100950, 100990, 100960, 100970, 100980, 
    101020, 101030, 101030, 101020, 101050, 101030, 101040, 101030, 100970, 
    100940, 100980, 101090, 101130, 101170, 101260, 101320, 101360, 101390, 
    101440, 101430, 101480, 101530, 101630, 101700, 101710, 101710, 101780, 
    101810, 101820, 101840, 101860, 101890, 101910, 101900, 101920, 101980, 
    102000, 102020, 102050, 102060, 102050, 102050, 102030, 102050, 102040, 
    102010, 102030, 101990, 101980, 101960, 101960, 101890, 101910, 101900, 
    101870, 101830, 101800, 101790, 101740, 101720, 101690, 101650, 101590, 
    101530, 101490, 101460, 101410, 101340, 101290, 101260, 101220, 101200, 
    101140, 101110, 101060, 101020, 100990, 100950, 100920, 100920, 100930, 
    100930, 100940, 100930, 100940, 100940, 100970, 100970, 100950, 100930, 
    100920, 100950, 100970, 101010, 101020, 101040, 101060, 101070, 101060, 
    101070, 101080, 101080, 101070, 101070, 101080, 101100, 101150, 101150, 
    101150, 101140, 101150, 101150, 101170, 101220, 101230, 101240, 101240, 
    101220, 101200, 101160, 101090, 101060, 101030, 101000, 100940, 100910, 
    100860, 100810, 100810, 100780, 100750, 100780, 100790, 100800, 100800, 
    100790, 100790, 100770, 100780, 100780, 100810, 100790, 100800, 100800, 
    100820, 100810, 100790, 100800, 100800, 100790, 100810, 100810, 100730, 
    100690, 100650, 100700, 100540, 100480, 100410, 100380, 100420, 100300, 
    100190, 100150, 100070, 100150, 100070, 100100, 100060, 100160, 100220, 
    100190, 100190, 100200, 100220, 100240, 100310, 100380, 100410, 100430, 
    100480, 100540, 100580, 100620, 100630, 100660, 100670, 100690, 100710, 
    100750, 100770, 100780, 100820, 100820, 100840, 100860, 100890, 100880, 
    100890, 100890, 100910, 100950, 101050, 100990, 100990, 101010, 101010, 
    101080, 100960, 101060, 101060, 101080, 101170, 101130, 101210, 101170, 
    101170, 101240, 101220, 101240, 101290, 101280, 101280, 101310, 101420, 
    101390, 101420, 101510, 101490, 101520, 101560, 101570, 101650, 101640, 
    101670, 101710, 101760, 101820, 101840, 101890, 101840, 101930, 102020, 
    101990, 102000, 102040, 102070, 102090, 102120, 102160, 102190, 102210, 
    102230, 102230, 102260, 102260, 102250, 102280, 102280, 102270, 102240, 
    102220, 102100, 102160, 102030, 102310, 102090, 101990, 101950, 101860, 
    101770, 101700, 101710, 101480, 100990, 101440, 101370, 101540, 101130, 
    100930, 101000, 100910, 100880, 100860, 100720, 101010, 100820, 100870, 
    100950, 100960, 100970, 101000, 101020, 101020, 101040, 101040, 101050, 
    101080, 101110, 101160, 101110, 101110, 101100, 101110, 101210, 101100, 
    101100, 101150, 101230, 101460, 101260, 101270, 101310, 101350, 101330, 
    101320, 101290, 101270, 101210, 101170, 101170, 101160, 101140, 101140, 
    101150, 101160, 101160, 101160, 101180, 101210, 101220, 101240, 101260, 
    101270, 101260, 101310, 101310, 101300, 101300, 101280, 101300, 101420, 
    101300, 101280, 101270, 101270, 101340, 101260, 101220, 101180, 101130, 
    101050, 101020, 100960, 100840, 100760, 100660, 100610, 100560, 100490, 
    100390, 100340, 100280, 100230, 100170, 100120, 100110, 100080, 100070, 
    100080, 100090, 100160, 100110, 100110, 100110, 100110, 100130, 100130, 
    100140, 100150, 100140, 100240, 100140, 100120, 100120, 100090, 100060, 
    100030, 100270, 100010, 100010, 100000, 100010, 100010, 100030, 100060, 
    100100, 100100, 100150, 100190, 100330, 100250, 100240, 100440, 100260, 
    100300, 100280, 100310, 100380, 100300, 100350, 100330, 100350, 100370, 
    100370, 100420, 100430, 100500, 100560, 100600, 100650, 100690, 100740, 
    100820, 100790, 100790, 100840, 100820, 100850, 100800, 100810, 100860, 
    100890, 100940, 100900, 100900, 100900, 100890, 100890, 100870, 100870, 
    100920, 100910, 100950, 100930, 100930, 100940, 100900, 100960, 100910, 
    100890, 100870, 100860, 100830, 100810, 100830, 100790, 100750, 100720, 
    100690, 100640, 100630, 100590, 100580, 100570, 100560, 100560, 100570, 
    100540, 100540, 100530, 100500, 100460, 100420, 100420, 100460, 100470, 
    100510, 100540, 100620, 100630, 100650, 100640, 100680, 100710, 100720, 
    100720, 100710, 100710, 100700, 100730, 100770, 100790, 100790, 100790, 
    100800, 100840, 100860, 100850, 100880, 100910, 100940, 100970, 100990, 
    101040, 101080, 101120, 101150, 101200, 101240, 101270, 101310, 101350, 
    101400, 101450, 101490, 101520, 101570, 101600, 101620, 101630, 101650, 
    101670, 101680, 101710, 101730, 101760, 101760, 101770, 101770, 101770, 
    101780, 101770, 101770, 101780, 101770, 101780, 101780, 101790, 101760, 
    101720, 101730, 101690, 101650, 101580, 101560, 101550, 101470, 101420, 
    101350, 101330, 101290, 101250, 101170, 101140, 101090, 101040, 101010, 
    100950, 100910, 100880, 100860, 100830, 100840, 100830, 100840, 100860, 
    100830, 100870, 100860, 100860, 100880, 100940, 100970, 100980, 100990, 
    101010, 101040, 101030, 101040, 101040, 101060, 101050, 101060, 101120, 
    101140, 101170, 101210, 101240, 101270, 101310, 101340, 101350, 101370, 
    101400, 101400, 101440, 101460, 101480, 101480, 101500, 101500, 101530, 
    101530, 101530, 101550, 101570, 101580, 101590, 101600, 101630, 101620, 
    101660, 101670, 101680, 101690, 101710, 101720, 101730, 101740, 101770, 
    101780, 101790, 101800, 101810, 101790, 101800, 101830, 101800, 101790, 
    101780, 101770, 101760, 101770, 101750, 101730, 101720, 101720, 101710, 
    101690, 101680, 101650, 101640, 101610, 101600, 101580, 101570, 101560, 
    101550, 101530, 101510, 101490, 101450, 101430, 101420, 101410, 101410, 
    101440, 101410, 101410, 101420, 101430, 101460, 101450, 101460, 101470, 
    101480, 101490, 101500, 101510, 101550, 101530, 101520, 101520, 101530, 
    101530, 101520, 101510, 101500, 101500, 101510, 101530, 101540, 101540, 
    101540, 101540, 101540, 101510, 101510, 101490, 101470, 101460, 101440, 
    101420, 101380, 101350, 101330, 101300, 101270, 101220, 101130, 101090, 
    100990, 101060, 101000, 100960, 100910, 100900, 100870, 100850, 100860, 
    100760, 100710, 100650, 100580, 100550, 100450, 100430, 100270, 100160, 
    100030, 99860, 99580, 99450, 99360, 99370, 99430, 99410, 99440, 99430, 
    99410, 99160, 99200, 99320, 99410, 99480, 99610, 99670, 99780, 99860, 
    99950, 100050, 100130, 100260, 100350, 100480, 100550, 100620, 100690, 
    100740, 100780, 100840, 100890, 100960, 101030, 101080, 101130, 101180, 
    101230, 101290, 101330, 101350, 101410, 101460, 101520, 101580, 101630, 
    101720, 101740, 101820, 101860, 101880, 101900, 101970, 102000, 102000, 
    102010, 102070, 102110, 102160, 102160, 102200, 102230, 102230, 102210, 
    102220, 102250, 102270, 102250, 102280, 102290, 102290, 102330, 102320, 
    102340, 102330, 102330, 102300, 102290, 102290, 102310, 102310, 102320, 
    102340, 102350, 102360, 102350, 102340, 102320, 102300, 102280, 102300, 
    102300, 102320, 102320, 102330, 102340, 102330, 102330, 102360, 102360, 
    102370, 102360, 102390, 102420, 102440, 102470, 102500, 102540, 102540, 
    102560, 102560, 102560, 102570, 102590, 102600, 102600, 102620, 102620, 
    102620, 102610, 102610, 102600, 102600, 102570, 102550, 102550, 102500, 
    102500, 102500, 102470, 102420, 102380, 102380, 102390, 102370, 102350, 
    102300, 102260, 102240, 102210, 102250, 102220, 102160, 102150, 102170, 
    102180, 102170, 102110, 102100, 102070, 102070, 102080, 102090, 102100, 
    102110, 102050, 102090, 102090, 102090, 102080, 102060, 102060, 102040, 
    102000, 102010, 102000, 102010, 101960, 101990, 102010, 101990, 101970, 
    101970, 101920, 101940, 101920, 101800, 101840, 101920, 101800, 101770, 
    101740, 101780, 101800, 101800, 101770, 101720, 101710, 101680, 101730, 
    101720, 101720, 101690, 101680, 101760, 101780, 101750, 101700, 101760, 
    101720, 101770, 101780, 101710, 101640, 101690, 101710, 101720, 101730, 
    101740, 101700, 101580, 101670, 101570, 101550, 101540, 101490, 101450, 
    101400, 101360, 101470, 101430, 101400, 101400, 101440, 101460, 101440, 
    101480, 101460, 101480, 101460, 101440, 101430, 101420, 101390, 101390, 
    101360, 101370, 101340, 101320, 101320, 101290, 101250, 101230, 101220, 
    101200, 101170, 101170, 101150, 101150, 101140, 101120, 101110, 101090, 
    101080, 101080, 101080, 101050, 101040, 101040, 101020, 101010, 101030, 
    101050, 101040, 101010, 101000, 100990, 101010, 101020, 100990, 100980, 
    101010, 101020, 100970, 100970, 100970, 100980, 101000, 100970, 100970, 
    100990, 100970, 100940, 100900, 100880, 100850, 100850, 100840, 100820, 
    100860, 100850, 100820, 100780, 100770, 100710, 100700, 100690, 100680, 
    100660, 100640, 100650, 100640, 100620, 100610, 100600, 100630, 100630, 
    100630, 100660, 100670, 100700, 100730, 100780, 100800, 100830, 100850, 
    100860, 100950, 101000, 101020, 101030, 101090, 101150, 101180, 101250, 
    101280, 101280, 101290, 101290, 101300, 101330, 101340, 101360, 101360, 
    101370, 101380, 101360, 101370, 101380, 101360, 101340, 101290, 101270, 
    101260, 101260, 101230, 101260, 101260, 101250, 101240, 101220, 101120, 
    101070, 101030, 101040, 100940, 100920, 100960, 100960, 100830, 100750, 
    100660, 100580, 100510, 100400, 100340, 100290, 100230, 100200, 100240, 
    100260, 100310, 100440, 100400, 100420, 100390, 100400, 100340, 100320, 
    100330, 100300, 100270, 100230, 100210, 100200, 100190, 100170, 100140, 
    100130, 100120, 100070, 100060, 100060, 100060, 100070, 100100, 100120, 
    100080, 100090, 100070, 100050, 100010, 99980, 99950, 99940, 99940, 
    100010, 100020, 100040, 100050, 100090, 100130, 100150, 100180, 100210, 
    100270, 100290, 100320, 100360, 100410, 100470, 100520, 100570, 100600, 
    100620, 100640, 100700, 100780, 100850, 100880, 100910, 100960, 101020, 
    101090, 101130, 101150, 101180, 101200, 101270, 101350, 101410, 101480, 
    101540, 101550, 101580, 101590, 101610, 101630, 101640, 101630, 101670, 
    101670, 101680, 101680, 101680, 101690, 101700, 101700, 101700, 101710, 
    101690, 101680, 101700, 101710, 101720, 101750, 101760, 101760, 101770, 
    101800, 101810, 101820, 101820, 101820, 101810, 101820, 101810, 101810, 
    101800, 101790, 101770, 101750, 101710, 101710, 101680, 101670, 101640, 
    101640, 101610, 101600, 101590, 101550, 101500, 101530, 101460, 101430, 
    101390, 101350, 101340, 101330, 101310, 101310, 101300, 101280, 101250, 
    101250, 101250, 101270, 101270, 101280, 101300, 101310, 101330, 101370, 
    101390, 101410, 101450, 101480, 101520, 101590, 101620, 101640, 101650, 
    101680, 101700, 101720, 101760, 101750, 101700, 101720, 101760, 101800, 
    101830, 101850, 101880, 101920, 101930, 101980, 102040, 102090, 102140, 
    102170, 102190, 102230, 102250, 102280, 102290, 102290, 102310, 102330, 
    102370, 102380, 102370, 102370, 102360, 102380, 102360, 102350, 102360, 
    102360, 102350, 102370, 102360, 102350, 102360, 102350, 102330, 102310, 
    102320, 102300, 102290, 102270, 102240, 102240, 102250, 102220, 102180, 
    102190, 102170, 102160, 102150, 102120, 102100, 102070, 102060, 102060, 
    102050, 102050, 102020, 101990, 101980, 101950, 101940, 101910, 101870, 
    101840, 101830, 101810, 101780, 101740, 101710, 101680, 101650, 101640, 
    101600, 101560, 101510, 101490, 101480, 101450, 101430, 101420, 101380, 
    101360, 101330, 101300, 101280, 101250, 101220, 101210, 101180, 101170, 
    101170, 101150, 101120, 101110, 101090, 101060, 101030, 101020, 101000, 
    100980, 100980, 101000, 101030, 101030, 101010, 100990, 100990, 100970, 
    100950, 100870, 100830, 100810, 100790, 100770, 100740, 100720, 100710, 
    100710, 100700, 100700, 100710, 100720, 100700, 100710, 100720, 100770, 
    100810, 100840, 100860, 100890, 100880, 100910, 100920, 100930, 100950, 
    100970, 100980, 100980, 100990, 101000, 101010, 101010, 100990, 100980, 
    100970, 100950, 100930, 100930, 100920, 100920, 100910, 100920, 100930, 
    100940, 100960, 100990, 101020, 101050, 101090, 101120, 101120, 101160, 
    101190, 101210, 101220, 101250, 101260, 101260, 101250, 101250, 101260, 
    101260, 101250, 101270, 101300, 101330, 101320, 101300, 101290, 101310, 
    101300, 101270, 101240, 101200, 101180, 101150, 101110, 101080, 101070, 
    101050, 101020, 101010, 101000, 101000, 100960, 100930, 100930, 100930, 
    100940, 100940, 100960, 100940, 100930, 100910, 100890, 100880, 100860, 
    100850, 100830, 100840, 100840, 100820, 100830, 100800, 100780, 100780, 
    100770, 100750, 100710, 100710, 100710, 100710, 100730, 100740, 100760, 
    100760, 100760, 100740, 100740, 100710, 100690, 100670, 100660, 100640, 
    100640, 100620, 100600, 100610, 100610, 100620, 100580, 100550, 100520, 
    100510, 100520, 100520, 100530, 100550, 100540, 100540, 100530, 100510, 
    100490, 100480, 100440, 100420, 100420, 100410, 100410, 100400, 100400, 
    100390, 100370, 100350, 100330, 100330, 100320, 100340, 100340, 100380, 
    100390, 100380, 100400, 100400, 100400, 100410, 100420, 100420, 100430, 
    100440, 100450, 100460, 100460, 100470, 100480, 100490, 100480, 100470, 
    100450, 100430, 100390, 100390, 100380, 100360, 100330, 100310, 100250, 
    100160, 100170, 100160, 100130, 100120, 100090, 100080, 100070, 100090, 
    100090, 100080, 100070, 100050, 100050, 100030, 100020, 100010, 100010, 
    100020, 100040, 100050, 100070, 100070, 100090, 100090, 100120, 100130, 
    100150, 100160, 100210, 100240, 100280, 100310, 100340, 100370, 100360, 
    100370, 100380, 100390, 100380, 100380, 100390, 100410, 100380, 100410, 
    100450, 100450, 100450, 100450, 100460, 100450, 100450, 100450, 100440, 
    100450, 100390, 100380, 100390, 100360, 100300, 100280, 100300, 100270, 
    100230, 100210, 100190, 100170, 100170, 100170, 100170, 100150, 100140, 
    100120, 100110, 100100, 100110, 100120, 100110, 100120, 100140, 100150, 
    100150, 100150, 100170, 100190, 100210, 100220, 100240, 100260, 100290, 
    100320, 100340, 100370, 100390, 100430, 100470, 100500, 100530, 100540, 
    100550, 100570, 100590, 100630, 100650, 100670, 100680, 100690, 100710, 
    100740, 100750, 100770, 100770, 100780, 100790, 100790, 100800, 100800, 
    100790, 100780, 100770, 100770, 100750, 100750, 100830, 100730, 100720, 
    100710, 100700, 100690, 100690, 100670, 100700, 100700, 100690, 100700, 
    100680, 100670, 100670, 100690, 100710, 100720, 100710, 100720, 100740, 
    100760, 100780, 100780, 100790, 100800, 100800, 100790, 100780, 100800, 
    100810, 100830, 100820, 100790, 100760, 100730, 100680, 100650, 100640, 
    100620, 100600, 100580, 100530, 100490, 100460, 100430, 100360, 100330, 
    100310, 100270, 100300, 100320, 100370, 100460, 100580, 100700, 100750, 
    100790, 100800, 100870, 100900, 100970, 101010, 101050, 101090, 101130, 
    101180, 101220, 101270, 101310, 101340, 101350, 101380, 101400, 101400, 
    101410, 101410, 101400, 101370, 101350, 101350, 101330, 101310, 101310, 
    101330, 101320, 101340, 101360, 101390, 101430, 101440, 101460, 101500, 
    101520, 101540, 101550, 101570, 101580, 101590, 101590, 101560, 101550, 
    101570, 101590, 101570, 101560, 101520, 101470, 101450, 101410, 101390, 
    101330, 101280, 101220, 101170, 101090, 101010, 100900, 100820, 100730, 
    100610, 100490, 100380, 100320, 100270, 100260, 100260, 100320, 100360, 
    100430, 100490, 100560, 100640, 100730, 100830, 100900, 100980, 101040, 
    101130, 101200, 101280, 101290, 101290, 101210, 101210, 101140, 101120, 
    101100, 100970, 100910, 100860, 100810, 100740, 100700, 100720, 100670, 
    100670, 100700, 100720, 100830, 100920, 100970, 101010, 101070, 101150, 
    101210, 101200, 101170, 101140, 101090, 101070, 101060, 101050, 101040, 
    101010, 101010, 100960, 100920, 100910, 100860, 100830, 100820, 100810, 
    100820, 100790, 100790, 100750, 100750, 100730, 100690, 100620, 100520, 
    100470, 100470, 100400, 100320, 100250, 100200, 100120, 100050, 99990, 
    99920, 99870, 99810, 99740, 99710, 99720, 99730, 99730, 99790, 99810, 
    99830, 99860, 99860, 99870, 99870, 99890, 99920, 99920, 99950, 99980, 
    99960, 100030, 100090, 100140, 100190, 100270, 100310, 100340, 100400, 
    100470, 100530, 100550, 100590, 100610, 100640, 100600, 100570, 100510, 
    100470, 100380, 100330, 100240, 100210, 100130, 100140, 100080, 100220, 
    100400, 100520, 100580, 100650, 100720, 100770, 100790, 100790, 100860, 
    100890, 100950, 101050, 101070, 101070, 101100, 101170, 101220, 101240, 
    101270, 101290, 101330, 101350, 101350, 101350, 101410, 101430, 101420, 
    101400, 101430, 101430, 101400, 101400, 101360, 101310, 101220, 101140, 
    101100, 101070, 101010, 100890, 100810, 100720, 100690, 100650, 100610, 
    100570, 100530, 100500, 100470, 100410, 100390, 100320, 100280, 100240, 
    100170, 100120, 100140, 100110, 100100, 100080, 100070, 100070, 100060, 
    100040, 100020, 100000, 99970, 99980, 99990, 99970, 99960, 99910, 99890, 
    99890, 99850, 99850, 99840, 99840, 99920, 100000, 100130, 100190, 100270, 
    100350, 100400, 100450, 100510, 100530, 100530, 100540, 100540, 100550, 
    100520, 100520, 100480, 100430, 100390, 100340, 100260, 100180, 100090, 
    100070, 100000, 99930, 99890, 99830, 99760, 99700, 99630, 99620, 99590, 
    99570, 99480, 99380, 99290, 99190, 99150, 99050, 98950, 98860, 98810, 
    98820, 98790, 98750, 98750, 98680, 98640, 98610, 98560, 98500, 98450, 
    98410, 98390, 98360, 98280, 98240, 98150, 98120, 98050, 98000, 97940, 
    97880, 97820, 97770, 97720, 97680, 97630, 97590, 97560, 97540, 97550, 
    97530, 97540, 97570, 97620, 97690, 97750, 97800, 97850, 97910, 97960, 
    98040, 98110, 98190, 98270, 98400, 98500, 98590, 98670, 98700, 98760, 
    98800, 98810, 98860, 98930, 99090, 99150, 99200, 99240, 99290, 99350, 
    99400, 99430, 99460, 99420, 99440, 99440, 99460, 99470, 99480, 99490, 
    99280, 99490, 99470, 99470, 99460, 99420, 99410, 99400, 99400, 99380, 
    99380, 99370, 99350, 99330, 99280, 99240, 99220, 99210, 99200, 99170, 
    99160, 99160, 99170, 99170, 99200, 99210, 99220, 99200, 99190, 99190, 
    99180, 99200, 99200, 99180, 99150, 99100, 99050, 99000, 98950, 98890, 
    98850, 98840, 98860, 98870, 98880, 98900, 98910, 98910, 98880, 98820, 
    98750, 98700, 98630, 98570, 98550, 98560, 98600, 98640, 98720, 98830, 
    98950, 99080, 99190, 99270, 99390, 99530, 99670, 99790, 99870, 99970, 
    100050, 100130, 100190, 100220, 100280, 100320, 100380, 100430, 100490, 
    100550, 100620, 100680, 100740, 100790, 100860, 100900, 100960, 101000, 
    101050, 101090, 101110, 101140, 101170, 101190, 101190, 101180, 101180, 
    101170, 101190, 101180, 101180, 101160, 101160, 101180, 101140, 101120, 
    101100, 101090, 101080, 101070, 101060, 101070, 101020, 100990, 100990, 
    100970, 100960, 100980, 100980, 100980, 101000, 101040, 101020, 101100, 
    101130, 101170, 101200, 101230, 101250, 101290, 101320, 101340, 101360, 
    101370, 101410, 101450, 101470, 101500, 101500, 101510, 101490, 101490, 
    101480, 101460, 101460, 101450, 101430, 101410, 101410, 101370, 101350, 
    101320, 101280, 101280, 101230, 101210, 101180, 101150, 101120, 101100, 
    101080, 101030, 101000, 100980, 100950, 100930, 100890, 100870, 100810, 
    100770, 100760, 100730, 100700, 100670, 100630, 100620, 100600, 100570, 
    100550, 100540, 100570, 100600, 100630, 100670, 100700, 100750, 100800, 
    100840, 100880, 100920, 100970, 101030, 101110, 101160, 101230, 101250, 
    101300, 101340, 101410, 101440, 101450, 101500, 101550, 101600, 101640, 
    101660, 101720, 101730, 101760, 101770, 101770, 101790, 101790, 101810, 
    101800, 101850, 101860, 101860, 101870, 101900, 101900, 101920, 101930, 
    101930, 101920, 101950, 101950, 101920, 101990, 101990, 102020, 102050, 
    102050, 102040, 102030, 102020, 102040, 102060, 102040, 102050, 102100, 
    102090, 102110, 102160, 102110, 102110, 102120, 102090, 102070, 102070, 
    102070, 102050, 102050, 102040, 102020, 102010, 102010, 101970, 101950, 
    101960, 101960, 101890, 101860, 101880, 101890, 101880, 101830, 101820, 
    101800, 101780, 101760, 101730, 101730, 101710, 101720, 101700, 101710, 
    101740, 101730, 101730, 101700, 101710, 101710, 101680, 101670, 101660, 
    101680, 101690, 101670, 101660, 101670, 101650, 101610, 101590, 101510, 
    101490, 101440, 101480, 101510, 101500, 101500, 101490, 101500, 101490, 
    101470, 101460, 101510, 101520, 101530, 101480, 101520, 101540, 101530, 
    101520, 101530, 101570, 101510, 101520, 101610, 101630, 101540, 101590, 
    101570, 101560, 101570, 101540, 101530, 101470, 101450, 101360, 101300, 
    101220, 101180, 101140, 100990, 100920, 100870, 100760, 100600, 100530, 
    100450, 100340, 100210, 100090, 100040, 99940, 99810, 99680, 99630, 
    99610, 99530, 99410, 99460, 99390, 99320, 99250, 99280, 99230, 99190, 
    99250, 99230, 99280, 99340, 99380, 99460, 99570, 99670, 99760, 99870, 
    99960, 100080, 100180, 100310, 100440, 100550, 100590, 100700, 100810, 
    100890, 100990, 101070, 101150, 101240, 101300, 101410, 101480, 101530, 
    101610, 101680, 101750, 101810, 101830, 101860, 101940, 102000, 102000, 
    102050, 102050, 102050, 102060, 102060, 102090, 102060, 102040, 102010, 
    101970, 101960, 101940, 101890, 101830, 101800, 101750, 101710, 101670, 
    101650, 101580, 101510, 101480, 101420, 101360, 101310, 101280, 101270, 
    101240, 101240, 101200, 101180, 101150, 101130, 101100, 100980, 100970, 
    100970, 100910, 100860, 100880, 100790, 100750, 100730, 100730, 100680, 
    100690, 100680, 100670, 100690, 100630, 100600, 100550, 100440, 100310, 
    100240, 100120, 99850, 99730, 99590, 99600, 99350, 99230, 99170, 99050, 
    99060, 99150, 99200, 99330, 99450, 99630, 99800, 99960, 100190, 100310, 
    100360, 100470, 100450, 100500, 100560, 100600, 100650, 100660, 100720, 
    100780, 100870, 100950, 101020, 101090, 101140, 101230, 101270, 101350, 
    101370, 101490, 101490, 101580, 101600, 101650, 101660, 101660, 101660, 
    101660, 101680, 101680, 101690, 101720, 101740, 101770, 101780, 101780, 
    101800, 101750, 101740, 101700, 101650, 101610, 101520, 101460, 101350, 
    101160, 100930, 100720, 100670, 100630, 100590, 100570, 100590, 100630, 
    100690, 100730, 100810, 100860, 100910, 101020, 101090, 101170, 101180, 
    101120, 101100, 101170, 101110, 101060, 101010, 101010, 101010, 100980, 
    101010, 101080, 101150, 101240, 101320, 101390, 101440, 101520, 101600, 
    101700, 101780, 101850, 101870, 101890, 101880, 101880, 101930, 101930, 
    101940, 101950, 101920, 101910, 101890, 101860, 101840, 101820, 101800, 
    101780, 101780, 101800, 101800, 101830, 101860, 101870, 101920, 101910, 
    101970, 101980, 102040, 102060, 102090, 102110, 102100, 102110, 102080, 
    102070, 102050, 102030, 102000, 101940, 101850, 101800, 101780, 101740, 
    101710, 101690, 101700, 101680, 101690, 101690, 101690, 101680, 101710, 
    101710, 101700, 101730, 101740, 101760, 101780, 101790, 101790, 101820, 
    101820, 101800, 101790, 101810, 101820, 101840, 101850, 101830, 101810, 
    101770, 101790, 101760, 101750, 101760, 101780, 101740, 101750, 101780, 
    101800, 101810, 101810, 101870, 101900, 101890, 101910, 101930, 101930, 
    101900, 101890, 101920, 101890, 101850, 101820, 101820, 101820, 101760, 
    101680, 101630, 101570, 101450, 101340, 101310, 101230, 101140, 100950, 
    100920, 100830, 100810, 100740, 100760, 100720, 100720, 100720, 100710, 
    100680, 100630, 100600, 100560, 100520, 100510, 100470, 100430, 100400, 
    100370, 100320, 100310, 100280, 100280, 100280, 100310, 100310, 100290, 
    100270, 100270, 100280, 100270, 100280, 100290, 100290, 100330, 100350, 
    100370, 100360, 100410, 100410, 100420, 100450, 100460, 100460, 100500, 
    100600, 100580, 100560, 100550, 100530, 100490, 100440, 100440, 100340, 
    100290, 100250, 100150, 100040, 100050, 99970, 99910, 99860, 99730, 
    99550, 99410, 99220, 99140, 99080, 98970, 98900, 98890, 98910, 98940, 
    98960, 98980, 98990, 99030, 99050, 99040, 99080, 99110, 99160, 99200, 
    99240, 99260, 99290, 99290, 99300, 99280, 99250, 99290, 99250, 99280, 
    99310, 99340, 99350, 99360, 99400, 99420, 99410, 99410, 99410, 99420, 
    99430, 99430, 99450, 99520, 99550, 99520, 99480, 99490, 99510, 99540, 
    99560, 99560, 99570, 99600, 99620, 99640, 99720, 99740, 99770, 99790, 
    99810, 99810, 99880, 99940, 100000, 100040, 100030, 100060, 100090, 
    100100, 100130, 100140, 100160, 100180, 100280, 100370, 100450, 100520, 
    100610, 100680, 100760, 100820, 100890, 100960, 101010, 101020, 101070, 
    101130, 101210, 101280, 101370, 101440, 101520, 101630, 101680, 101780, 
    101870, 101960, 102060, 102140, 102220, 102280, 102300, 102350, 102370, 
    102390, 102400, 102340, 102280, 102210, 102160, 102110, 102080, 102010, 
    101890, 101830, 101750, 101670, 101580, 101510, 101430, 101360, 101320, 
    101250, 101190, 101140, 101050, 100970, 100850, 100760, 100620, 100550, 
    100490, 100440, 100400, 100400, 100440, 100470, 100530, 100590, 100660, 
    100750, 100850, 100960, 101150, 101370, 101560, 101680, 101800, 101930, 
    102080, 102160, 102280, 102370, 102450, 102540, 102650, 102620, 102650, 
    102630, 102630, 102590, 102500, 102500, 102420, 102310, 102200, 102090, 
    101990, 101840, 101710, 101530, 101370, 101180, 101080, 100910, 100780, 
    100650, 100520, 100490, 100390, 100380, 100410, 100430, 100410, 100450, 
    100490, 100530, 100620, 100710, 100810, 100860, 100970, 101070, 101090, 
    101290, 101320, 101460, 101570, 101650, 101790, 101920, 102060, 102160, 
    102290, 102330, 102400, 102450, 102500, 102480, 102540, 102560, 102540, 
    102530, 102520, 102550, 102560, 102600, 102650, 102660, 102660, 102680, 
    102690, 102710, 102700, 102710, 102660, 102630, 102580, 102500, 102430, 
    102340, 102300, 102250, 102200, 102200, 102120, 102080, 102030, 101970, 
    101920, 101830, 101790, 101720, 101660, 101620, 101550, 101540, 101510, 
    101500, 101450, 101450, 101420, 101390, 101360, 101340, 101330, 101350, 
    101370, 101420, 101450, 101530, 101560, 101580, 101520, 101560, 101550, 
    101520, 101490, 101450, 101420, 101410, 101380, 101300, 101230, 101170, 
    101100, 101040, 100990, 100950, 100920, 100920, 100940, 100960, 100980, 
    101010, 101040, 101080, 101130, 101180, 101230, 101240, 101280, 101310, 
    101330, 101360, 101400, 101440, 101490, 101520, 101550, 101580, 101600, 
    101620, 101660, 101680, 101710, 101740, 101790, 101820, 101840, 101850, 
    101890, 101910, 101950, 101980, 102010, 102040, 102050, 102090, 102140, 
    102180, 102190, 102180, 102200, 102190, 102210, 102220, 102190, 102170, 
    102170, 102170, 102160, 102130, 102100, 102080, 102040, 102040, 101950, 
    101920, 101900, 101820, 101810, 101740, 101670, 101600, 101500, 101370, 
    101230, 101110, 100980, 100830, 100690, 100550, 100460, 100380, 100290, 
    100230, 100160, 100130, 100090, 100080, 100060, 100000, 99960, 99880, 
    99800, 99690, 99640, 99550, 99520, 99480, 99510, 99590, 99650, 99600, 
    99550, 99470, 99430, 99420, 99310, 99330, 99320, 99380, 99460, 99590, 
    99730, 99860, 99960, 100150, 100200, 100360, 100410, 100510, 100640, 
    100780, 100880, 100990, 101010, 101050, 101090, 101090, 101160, 101300, 
    101370, 101380, 101430, 101460, 101490, 101520, 101540, 101530, 101550, 
    101550, 101590, 101620, 101650, 101660, 101690, 101710, 101720, 101740, 
    101730, 101720, 101720, 101700, 101680, 101660, 101610, 101600, 101560, 
    101530, 101510, 101470, 101470, 101460, 101450, 101440, 101460, 101460, 
    101500, 101500, 101500, 101520, 101550, 101550, 101560, 101570, 101550, 
    101550, 101570, 101540, 101540, 101560, 101540, 101510, 101460, 101420, 
    101410, 101420, 101420, 101420, 101400, 101440, 101450, 101460, 101440, 
    101440, 101430, 101420, 101410, 101390, 101360, 101330, 101280, 101270, 
    101250, 101230, 101210, 101200, 101190, 101170, 101140, 101150, 101150, 
    101140, 101180, 101200, 101190, 101260, 101290, 101290, 101290, 101290, 
    101310, 101310, 101300, 101280, 101230, 101210, 101150, 101130, 101020, 
    100960, 100930, 100860, 100760, 100730, 100640, 100600, 100540, 100520, 
    100510, 100530, 100580, 100710, 100750, 100770, 100810, 100880, 101010, 
    101040, 101090, 101210, 101300, 101410, 101480, 101560, 101610, 101650, 
    101660, 101720, 101760, 101810, 101890, 101970, 102070, 102140, 102220, 
    102330, 102450, 102530, 102620, 102710, 102810, 102910, 103010, 103070, 
    103140, 103170, 103210, 103220, 103220, 103240, 103250, 103240, 103200, 
    103210, 103150, 103120, 103170, 103120, 103070, 103050, 102980, 102930, 
    102920, 102860, 102830, 102780, 102750, 102670, 102680, 102690, 102690, 
    102690, 102660, 102670, 102690, 102670, 102640, 102680, 102640, 102630, 
    102650, 102620, 102610, 102560, 102510, 102450, 102440, 102440, 102360, 
    102410, 102310, 102280, 102260, 102200, 102160, 102120, 102060, 102010, 
    101960, 101910, 101890, 101860, 101810, 101790, 101750, 101710, 101680, 
    101640, 101600, 101520, 101500, 101460, 101410, 101370, 101340, 101300, 
    101250, 101230, 101180, 101140, 101130, 101090, 101050, 101040, 101010, 
    100910, 100950, 101000, 100990, 101000, 101070, 101130, 101150, 101210, 
    101220, 101230, 101230, 101280, 101300, 101290, 101280, 101320, 101350, 
    101350, 101380, 101380, 101380, 101420, 101430, 101450, 101460, 101490, 
    101530, 101560, 101540, 101540, 101520, 101520, 101520, 101520, 101540, 
    101570, 101580, 101620, 101650, 101680, 101710, 101710, 101700, 101720, 
    101730, 101750, 101750, 101770, 101770, 101770, 101820, 101850, 101850, 
    101860, 101870, 101910, 101920, 101930, 101930, 101970, 102040, 102070, 
    102060, 102070, 102140, 102180, 102180, 102160, 102250, 102380, 102440, 
    102490, 102540, 102580, 102620, 102750, 102790, 102820, 102890, 102970, 
    103020, 103060, 103090, 103130, 103180, 103210, 103250, 103260, 103310, 
    103340, 103360, 103380, 103400, 103400, 103410, 103420, 103430, 103430, 
    103460, 103490, 103500, 103530, 103530, 103550, 103520, 103540, 103540, 
    103540, 103550, 103550, 103560, 103550, 103550, 103550, 103540, 103510, 
    103500, 103490, 103480, 103450, 103440, 103440, 103430, 103450, 103430, 
    103440, 103440, 103430, 103430, 103450, 103430, 103430, 103440, 103440, 
    103440, 103430, 103410, 103410, 103390, 103390, 103370, 103340, 103300, 
    103280, 103270, 103260, 103260, 103240, 103210, 103180, 103140, 103120, 
    103080, 103040, 103020, 103000, 102980, 102940, 102920, 102880, 102870, 
    102840, 102820, 102800, 102790, 102780, 102780, 102790, 102800, 102790, 
    102800, 102810, 102840, 102860, 102830, 102820, 102840, 102860, 102880, 
    102900, 102900, 102910, 102920, 102940, 102950, 102950, 102940, 102930, 
    102960, 102960, 102970, 102970, 102970, 102980, 102970, 103010, 103010, 
    103010, 103000, 102990, 102970, 102970, 102970, 102960, 102950, 102960, 
    102940, 102910, 102890, 102880, 102850, 102820, 102790, 102760, 102740, 
    102720, 102690, 102650, 102650, 102630, 102590, 102560, 102520, 102480, 
    102410, 102380, 102340, 102310, 102260, 102220, 102180, 102120, 102080, 
    102050, 102030, 102010, 102000, 102010, 102030, 102080, 102120, 102140, 
    102170, 102180, 102190, 102210, 102210, 102210, 102210, 102210, 102220, 
    102220, 102190, 102170, 102160, 102130, 102100, 102060, 102020, 101950, 
    101900, 101850, 101750, 101690, 101600, 101530, 101460, 101370, 101300, 
    101240, 101180, 101120, 101050, 100990, 100930, 100860, 100790, 100730, 
    100680, 100620, 100560, 100490, 100450, 100390, 100330, 100260, 100200, 
    100130, 100020, 99970, 99900, 99810, 99740, 99640, 99560, 99480, 99360, 
    99330, 99190, 99070, 99020, 98910, 98800, 98670, 98610, 98510, 98370, 
    98230, 98140, 98080, 98020, 98000, 98030, 98180, 98330, 98440, 98560, 
    98750, 98700, 98950, 98770, 98920, 99040, 99150, 99260, 99540, 99570, 
    99540, 99690, 99820, 99850, 99780, 99870, 99980, 100020, 100060, 100090, 
    100250, 100340, 100410, 100520, 100550, 100710, 100770, 100860, 100870, 
    100940, 101090, 101150, 101250, 101290, 101350, 101430, 101460, 101500, 
    101580, 101610, 101650, 101660, 101690, 101730, 101800, 101840, 101870, 
    101890, 101920, 101970, 101980, 102010, 102060, 102090, 102130, 102150, 
    102170, 102200, 102230, 102240, 102240, 102240, 102250, 102260, 102250, 
    102250, 102220, 102190, 102170, 102160, 102130, 102090, 102080, 102040, 
    102010, 101970, 101930, 101870, 101830, 101820, 101800, 101790, 101800, 
    101810, 101790, 101720, 101660, 101620, 101570, 101530, 101520, 101480, 
    101470, 101470, 101450, 101420, 101380, 101310, 101280, 101250, 101210, 
    101160, 101110, 101070, 101030, 100990, 100960, 100930, 100880, 100840, 
    100800, 100770, 100720, 100670, 100600, 100540, 100490, 100460, 100420, 
    100410, 100400, 100360, 100260, 100230, 100190, 100150, 100130, 100100, 
    100070, 100050, 100040, 100050, 100040, 100020, 99980, 99930, 99870, 
    99830, 99770, 99670, 99600, 99480, 99440, 99370, 99340, 99190, 99000, 
    98900, 98810, 98670, 98560, 98380, 98220, 98060, 97950, 97830, 97730, 
    97710, 97610, 97530, 97550, 97650, 97730, 97870, 97920, 98000, 98050, 
    98130, 98230, 98250, 98290, 98320, 98420, 98510, 98580, 98670, 98760, 
    98850, 98930, 99000, 99080, 99100, 99120, 99150, 99150, 99130, 99080, 
    98990, 98930, 98840, 98800, 98730, 98690, 98690, 98680, 98710, 98750, 
    98780, 98810, 98830, 98830, 98870, 98860, 98910, 98960, 98970, 99000, 
    99160, 99310, 99420, 99550, 99760, 99880, 100080, 100300, 100460, 100610, 
    100730, 100800, 100970, 101100, 101160, 101220, 101320, 101390, 101420, 
    101490, 101530, 101600, 101660, 101680, 101740, 101780, 101820, 101810, 
    101860, 101900, 101930, 101960, 101960, 101980, 101990, 101970, 101950, 
    101950, 101930, 101940, 101920, 101920, 101920, 101870, 101810, 101770, 
    101800, 101750, 101710, 101680, 101630, 101580, 101540, 101480, 101450, 
    101390, 101350, 101350, 101310, 101280, 101240, 101190, 101150, 101110, 
    101030, 100980, 100960, 100910, 100890, 100830, 100800, 100760, 100720, 
    100740, 100670, 100640, 100640, 100680, 100710, 100720, 100750, 100750, 
    100740, 100720, 100710, 100810, 100830, 100840, 100850, 100860, 100870, 
    100900, 100900, 100900, 100890, 100960, 100980, 101010, 101030, 101060, 
    101060, 101110, 101130, 101160, 101200, 101200, 101230, 101240, 101230, 
    101230, 101260, 101270, 101290, 101280, 101300, 101310, 101330, 101340, 
    101350, 101370, 101400, 101400, 101420, 101420, 101430, 101450, 101490, 
    101520, 101570, 101600, 101630, 101660, 101680, 101680, 101700, 101720, 
    101750, 101790, 101800, 101830, 101830, 101850, 101860, 101870, 101870, 
    101860, 101890, 101880, 101890, 101920, 101960, 101980, 101980, 101990, 
    101990, 101980, 102000, 102010, 101980, 101980, 101980, 101980, 101970, 
    101980, 101950, 101940, 101900, 101860, 101810, 101760, 101730, 101740, 
    101750, 101820, 101880, 101900, 101910, 101910, 101900, 101910, 101900, 
    101900, 101880, 101870, 101850, 101850, 101830, 101820, 101820, 101820, 
    101800, 101800, 101760, 101740, 101680, 101640, 101620, 101600, 101570, 
    101570, 101560, 101550, 101500, 101480, 101450, 101390, 101330, 101350, 
    101330, 101300, 101290, 101300, 101290, 101280, 101230, 101230, 101210, 
    101190, 101170, 101150, 101130, 101120, 101090, 101070, 101090, 101070, 
    101080, 101090, 101110, 101140, 101170, 101220, 101250, 101300, 101340, 
    101360, 101410, 101400, 101380, 101490, 101520, 101620, 101700, 101730, 
    101790, 101820, 101840, 101850, 101880, 101910, 101900, 101870, 101880, 
    101870, 101860, 101840, 101810, 101790, 101780, 101780, 101760, 101730, 
    101700, 101670, 101640, 101620, 101580, 101580, 101560, 101540, 101550, 
    101540, 101520, 101490, 101500, 101480, 101470, 101450, 101420, 101420, 
    101360, 101360, 101370, 101400, 101380, 101370, 101350, 101360, 101330, 
    101340, 101300, 101330, 101300, 101270, 101270, 101290, 101300, 101300, 
    101300, 101250, 101260, 101280, 101280, 101260, 101270, 101240, 101230, 
    101180, 101160, 101170, 101160, 101200, 101170, 101230, 101240, 101260, 
    101270, 101290, 101310, 101320, 101360, 101330, 101340, 101330, 101330, 
    101360, 101370, 101380, 101410, 101400, 101430, 101460, 101510, 101520, 
    101510, 101530, 101530, 101560, 101560, 101580, 101610, 101650, 101670, 
    101680, 101690, 101710, 101720, 101730, 101730, 101740, 101730, 101730, 
    101830, 101810, 101780, 101800, 101770, 101720, 101660, 101630, 101590, 
    101550, 101530, 101620, 101620, 101620, 101580, 101540, 101490, 101470, 
    101390, 101340, 101330, 101310, 101350, 101290, 101240, 101200, 101160, 
    101130, 101080, 101040, 101000, 100970, 100950, 100910, 100880, 100850, 
    100810, 100780, 100790, 100760, 100730, 100700, 100660, 100610, 100600, 
    100580, 100560, 100550, 100550, 100560, 100580, 100600, 100630, 100640, 
    100660, 100670, 100680, 100670, 100660, 100740, 100670, 100660, 100680, 
    100680, 100670, 100590, 100530, 100500, 100420, 100300, 100230, 100120, 
    99940, 99850, 99700, 99530, 99380, 99370, 99410, 99550, 99670, 99770, 
    99870, 99980, 100040, 100130, 100200, 100230, 100230, 100280, 100290, 
    100370, 100410, 100590, 100610, 100640, 100600, 100620, 100660, 100700, 
    100700, 100680, 100680, 100690, 100680, 100630, 100590, 100590, 100810, 
    100810, 100800, 100810, 100820, 100810, 100790, 100780, 100770, 100760, 
    100740, 100720, 100810, 100800, 100790, 100770, 100750, 100750, 100740, 
    100730, 100700, 100700, 100660, 100620, 100530, 100480, 100420, 100400, 
    100370, 100320, 100260, 100200, 100130, 100050, 99980, 99910, 99820, 
    99690, 99560, 99440, 99260, 99110, 99140, 99280, 99440, 99480, 99500, 
    99560, 99430, 99520, 99560, 99590, 99610, 99650, 99700, 99740, 99790, 
    99840, 99850, 99900, 99950, 100000, 100050, 100100, 100170, 100220, 
    100270, 100310, 100360, 100400, 100450, 100510, 100720, 100800, 100880, 
    100970, 101040, 101130, 101210, 101270, 101330, 101380, 101420, 101450, 
    101470, 101530, 101570, 101590, 101600, 101620, 101630, 101650, 101640, 
    101640, 101620, 101610, 101560, 101540, 101520, 101500, 101480, 101460, 
    101430, 101400, 101370, 101330, 101260, 101190, 101140, 101070, 101020, 
    100960, 100910, 100860, 100820, 100770, 100700, 100630, 100590, 100530, 
    100480, 100450, 100430, 100440, 100410, 100400, 100380, 100370, 100370, 
    100360, 100350, 100360, 100370, 100400, 100410, 100420, 100450, 100480, 
    100500, 100510, 100510, 100500, 100510, 100500, 100500, 100530, 100560, 
    100580, 100620, 100650, _, 100690, 100710, 100740, 100730, 100740, 
    100840, 100870, 100900, 100910, 100930, 100950, 100980, 100980, 100980, 
    100980, 100970, 100970, 101010, 101030, 101040, 101070, 101090, 101110, 
    101130, 101130, 101150, 101160, 101160, 101170, 101160, 101170, 101160, 
    101140, 101140, 101150, 101140, 101110, 101080, 101040, 101020, 100980, 
    100960, 100970, 100940, 100910, 100900, 100870, 100830, 100730, 100700, 
    100660, 100630, 100570, 100530, 100490, 100430, 100410, 100350, 100290, 
    100230, 100180, 100130, 100080, 100030, 99940, 99900, 99910, 99930, 
    99940, 99970, 99990, 100040, 100100, 100110, 100150, 100160, 100190, 
    100200, 100240, 100230, 100230, 100230, 100200, 100150, 100120, 100100, 
    100070, 99980, 99930, 99870, 99850, 99870, 99880, 99880, 99890, 99900, 
    99920, 99970, 100030, 100060, 100090, 100160, 100150, 100220, 100270, 
    100270, 100280, 100240, 100220, 100200, 100200, 100160, 100070, 100120, 
    100160, 100170, 100190, 100170, 100160, 100150, 100140, 100110, 100110, 
    100120, 100120, 100110, 100080, 100040, 100010, 99970, 99950, 99940, 
    99900, 99860, 99820, 99820, 99730, 99660, 99710, 99690, 99660, 99650, 
    99620, 99590, 99550, 99540, 99500, 99450, 99460, 99450, 99470, 99470, 
    99510, 99570, 99620, 99660, 99710, 99730, 99760, 99760, 99770, 99710, 
    99620, 99540, 99560, 99520, 99430, 99310, 99210, 99100, 98930, 98760, 
    98500, 98230, 97920, 97570, 97190, 96730, 96450, 96240, 96020, 95980, 
    96000, 96120, 96210, 96380, 96630, 96790, 97010, 97170, 97350, 97460, 
    97620, 97740, 97870, 97950, 98050, 98140, 98190, 98290, 98350, 98410, 
    98450, 98420, 98390, 98330, 98260, 98210, 98160, 98040, 97860, 97670, 
    97370, 97060, 96840, 96800, 96790, 96760, 96820, 96850, 96860, 96920, 
    96950, 96900, 96830, 96850, 96890, 96870, 96850, 96900, 96980, 97050, 
    97100, 97160, 97290, 97400, 97470, 97490, 97440, 97400, 97440, 97470, 
    97460, 97470, 97500, 97500, 97480, 97480, 97460, 97390, 97310, 97260, 
    97210, 97170, 97150, 97110, 97120, 97100, 97090, 97130, 97120, 97120, 
    97150, 97140, 97160, 97170, 97150, 97140, 97150, 97170, 97190, 97280, 
    97340, 97390, 97430, 97480, 97530, 97570, 97580, 97640, 97670, 97680, 
    97660, 97730, 97790, 97800, 97830, 97810, 97830, 97860, 97860, 97880, 
    97870, 97900, 97910, 97920, 97910, 97920, 97960, 97990, 97980, 98010, 
    98060, 98090, 98130, 98150, 98170, 98150, 98130, 98130, 98130, 98130, 
    98130, 98140, 98130, 98120, 98130, 98090, 98060, 98040, 98020, 98060, 
    98020, 97970, 97920, 97970, 97960, 97980, 98020, 98090, 98080, 98030, 
    98060, 98180, 98270, 98340, 98400, 98470, 98570, 98640, 98710, 98790, 
    98920, 98950, 99070, 99180, 99220, 99290, 99470, 99670, 99830, 99940, 
    100050, 100160, 100280, 100380, 100480, 100570, 100660, 100730, 100800, 
    100870, 100910, 100960, 100990, 101020, 101060, 101130, 101150, 101190, 
    101240, 101330, 101380, 101460, 101510, 101520, 101490, 101550, 101580, 
    101580, 101510, 101450, 101430, 101370, 101240, 101150, 101080, 100980, 
    100820, 100620, 100540, 100430, 100290, 100200, 100120, 100020, 100030, 
    99950, 99920, 99860, 99810, 99700, 99730, 99850, 99970, 100080, 100120, 
    100210, 100210, 100280, 100420, 100490, 100570, 100640, 100680, 100750, 
    100800, 100850, 100920, 100980, 101000, 101040, 101050, 101070, 101050, 
    101050, 101100, 101160, 101210, 101190, 101170, 101140, 101130, 101170, 
    101130, 101110, 101100, 101060, 101080, 101110, 101120, 101140, 101140, 
    101140, 101180, 101180, 101220, 101280, 101300, 101350, 101420, 101480, 
    101530, 101620, 101720, 101770, 101810, 101900, 101990, 102050, 102100, 
    102120, 102180, 102240, 102280, 102340, 102340, 102350, 102380, 102400, 
    102410, 102420, 102430, 102430, 102480, 102510, 102540, 102570, 102580, 
    102550, 102580, 102570, 102590, 102600, 102630, 102630, 102670, 102620, 
    102620, 102630, 102650, 102610, 102600, 102530, 102500, 102490, 102480, 
    102490, 102450, 102430, 102370, 102370, 102340, 102290, 102260, 102250, 
    102230, 102230, 102200, 102180, 102160, 102140, 102160, 102160, 102150, 
    102130, 102120, 102110, 102110, 102110, 102070, 102080, 102070, 102100, 
    102080, 102060, 102040, 102030, 102020, 102000, 101980, 101960, 101900, 
    101870, 101850, 101790, 101750, 101660, 101640, 101610, 101550, 101510, 
    101480, 101410, 101370, 101350, 101340, 101330, 101300, 101240, 101230, 
    101190, 101180, 101130, 101060, 100990, 100910, 100830, 100780, 100740, 
    100710, 100670, 100670, 100650, 100630, 100600, 100570, 100540, 100480, 
    100430, 100390, 100310, 100180, 99980, 99920, 99790, 99620, 99480, 99270, 
    99100, 98950, 98910, 98800, 98700, 98570, 98480, 98410, 98350, 98330, 
    98310, 98310, 98350, 98400, 98470, 98500, 98580, 98660, 98720, 98800, 
    98890, 98930, 98970, 98960, 98950, 98920, 98900, 98870, 98890, 98850, 
    98770, 98720, 98750, 98770, 98740, 98690, 98680, 98680, 98650, 98660, 
    98690, 98680, 98680, 98720, 98720, 98720, 98750, 98780, 98780, 98770, 
    98780, 98830, 98900, 98910, 98940, 98970, 98990, 99040, 99060, 99090, 
    99110, 99140, 99160, 99190, 99250, 99270, 99290, 99320, 99330, 99340, 
    99340, 99350, 99320, 99340, 99340, 99340, 99360, 99390, 99390, 99380, 
    99370, 99360, 99330, 99350, 99330, 99330, 99300, 99290, 99250, 99270, 
    99230, 99150, 99130, 99080, 99080, 99020, 98990, 98940, 98840, 98770, 
    98740, 98700, 98630, 98520, 98440, 98390, 98300, 98200, 98110, 98090, 
    98090, 98100, 98080, 98180, 98160, 98170, 98150, 98170, 98170, 98160, 
    98180, 98170, 98210, 98230, 98270, 98300, 98330, 98360, 98390, 98400, 
    98440, 98460, 98450, 98480, 98480, 98500, 98490, 98510, 98530, 98560, 
    98560, 98550, 98560, 98540, 98570, 98570, 98610, 98610, 98640, 98650, 
    98670, 98690, 98710, 98730, 98740, 98750, 98770, 98800, 98830, 98870, 
    98920, 98990, 99010, 99070, 99070, 99100, 99130, 99160, 99170, 99190, 
    99200, 99210, 99230, 99220, 99230, 99220, 99210, 99170, 99180, 99150, 
    99140, 99160, 99190, 99240, 99310, 99360, 99410, 99460, 99500, 99510, 
    99560, 99580, 99590, 99640, 99680, 99710, 99740, 99790, 99800, 99840, 
    99870, 99880, 99880, 99850, 99850, 99850, 99850, 99840, 99820, 99820, 
    99790, 99770, 99790, 99760, 99690, 99730, 99680, 99680, 99720, 99630, 
    99630, 99640, 99680, 99690, 99680, 99700, 99740, 99770, 99760, 99790, 
    99830, 99850, 99890, 99900, 99950, 99980, 100010, 100040, 100050, 100070, 
    100090, 100120, 100160, 100180, 100230, 100260, 100330, 100380, 100440, 
    100460, 100460, 100420, 100400, 100370, 100280, 100190, 100070, 99950, 
    99840, 99700, 99540, 99380, 99210, 99040, 98840, 98620, 98380, 98180, 
    98060, 97920, 97730, 97590, 97500, 97470, 97480, 97470, 97480, 97400, 
    97280, 97220, 97150, 97120, 97030, 96990, 96980, 96960, 96840, 96760, 
    96750, 96760, 96790, 96780, 96830, 97010, 97160, 97280, 97370, 97460, 
    97480, 97570, 97630, 97690, 97760, 97780, 97790, 97860, 97890, 97890, 
    97910, 97910, 97850, 97820, 97820, 97760, 97760, 97750, 97760, 97810, 
    97840, 97880, 97910, 97940, 97930, 97900, 97880, 97880, 97850, 97810, 
    97760, 97710, 97650, 97640, 97600, 97540, 97580, 97620, 97610, 97630, 
    97650, 97670, 97700, 97720, 97740, 97740, 97700, 97650, 97640, 97620, 
    97610, 97630, 97650, 97650, 97730, 97840, 97950, 98050, 98090, 98150, 
    98210, 98250, 98280, 98330, 98370, 98460, 98530, 98630, 98680, 98740, 
    98780, 98840, 98860, 98930, 98990, 99010, 99070, 99190, 99380, 99530, 
    99670, 99810, 99940, 100040, 100160, 100270, 100350, 100430, 100500, 
    100620, 100700, 100740, 100790, 100860, 100900, 100940, 100970, 101010, 
    101050, 101020, 101030, 101060, 101050, 101050, 101070, 101090, 101100, 
    101090, 101090, 101080, 101100, 101110, 101110, 101110, 101110, 101120, 
    101120, 101080, 101050, 101020, 100980, 100970, 100950, 100910, 100900, 
    100880, 100880, 100880, 100850, 100820, 100770, 100780, 100740, 100700, 
    100690, 100630, 100590, 100530, 100520, 100480, 100440, 100410, 100360, 
    100300, 100200, 100070, 99940, 99800, 99650, 99560, 99460, 99390, 99280, 
    99110, 98980, 98840, 98680, 98540, 98370, 98220, 98190, 98140, 98100, 
    98090, 98050, 98100, 98130, 98120, 98160, 98180, 98240, 98290, 98350, 
    98230, 98320, 98380, 98430, 98480, 98480, 98460, 98450, 98450, 98450, 
    98460, 98500, 98550, 98630, 98720, 98810, 98910, 98990, 99080, 99200, 
    99320, 99450, 99530, 99680, 99790, 99900, 100020, 100080, 100110, 100200, 
    100240, 100250, 100280, 100310, 100260, 100330, 100420, 100410, 100430, 
    100480, 100460, 100420, 100400, 100330, 100290, 100250, 100210, 100130, 
    100120, 100130, 100110, 100060, 100040, 99970, 99860, 99830, 99750, 
    99710, 99620, 99590, 99620, 99620, 99640, 99690, 99730, 99750, 99790, 
    99850, 99920, 99960, 100060, 100130, 100210, 100220, 100230, 100240, 
    100250, 100220, 100210, 100170, 100150, 100130, 100110, 100090, 100110, 
    100120, 100170, 100170, 100190, 100220, 100210, 100190, 100150, 100200, 
    100150, 100150, 100120, 100110, 100090, 100030, 99980, 99940, 99880, 
    99820, 99770, 99720, 99680, 99650, 99630, 99620, 99590, 99560, 99550, 
    99520, 99520, 99530, 99520, 99550, 99530, 99530, 99540, 99560, 99570, 
    99590, 99600, 99600, 99590, 99640, 99750, 99800, 99840, 99880, 99950, 
    100010, 100030, 100040, 100090, 100060, 100010, 100020, 100110, 100160, 
    100260, 100300, 100320, 100420, 100490, 100560, 100620, 100660, 100720, 
    100780, 100880, 100970, 101030, 101030, 101040, 101070, 101060, 101040, 
    101040, 101010, 101070, 101110, 101200, 101230, 101260, 101310, 101370, 
    101410, 101450, 101490, 101490, 101540, 101660, 101620, 101630, 101600, 
    101630, 101620, 101610, 101590, 101570, 101560, 101520, 101460, 101380, 
    101330, 101300, 101250, 101230, 101200, 101160, 101140, 101130, 101110, 
    101090, 101060, 101050, 101030, 101000, 100980, 100940, 100940, 100920, 
    100890, 100900, 100920, 100940, 100940, 100930, 100930, 100900, 100860, 
    100840, 100870, 100870, 100850, 100860, 100860, 100880, 100880, 100850, 
    100820, 100770, 100740, 100700, 100640, 100590, 100530, 100510, 100470, 
    100430, 100400, 100370, 100360, 100360, 100370, 100400, 100420, 100440, 
    100500, 100510, 100510, 100550, 100540, 100580, 100640, 100700, 100730, 
    100800, 100840, 100820, 100860, 100850, 100840, 100780, 100750, 100680, 
    100620, 100520, 100530, 100500, 100490, 100450, 100440, 100420, 100450, 
    100440, 100430, 100410, 100390, 100400, 100400, 100340, 100300, 100360, 
    100440, 100490, 100560, 100610, 100670, 100750, 100770, 100840, 100900, 
    100910, 100950, 100970, 101030, 101070, 101140, 101120, 101160, 101130, 
    101170, 101230, 101240, 101290, 101310, 101350, 101370, 101400, 101390, 
    101370, 101340, 101300, 101240, 101210, 101200, 101190, 101140, 101130, 
    101170, 101190, 101200, 101200, 101210, 101270, 101330, 101400, 101440, 
    101500, 101590, 101650, 101710, 101830, 101940, 102030, 102110, 102180, 
    102270, 102310, 102380, 102450, 102530, 102590, 102630, 102700, 102790, 
    102850, 102850, 102890, 102870, 102830, 102840, 102820, 102790, 102770, 
    102740, 102730, 102740, 102730, 102730, 102720, 102760, 102760, 102750, 
    102760, 102730, 102750, 102750, 102760, 102800, 102760, 102770, 102750, 
    102750, 102720, 102710, 102730, 102710, 102710, 102830, 102830, 102810, 
    102830, 102820, 102780, 102780, 102760, 102720, 102720, 102680, 102680, 
    102650, 102610, 102550, 102500, 102460, 102370, 102230, 102130, 102020, 
    101920, 101750, 101630, 101510, 101430, 101300, 101210, 101190, 101050, 
    100970, 100930, 100940, 100980, 101010, 101020, 100980, 100980, 100980, 
    100910, 100860, 100780, 100710, 100590, 100470, 100350, 100220, 100090, 
    99990, 99840, 99680, 99550, 99430, 99310, 99160, 99010, 98880, 98760, 
    98620, 98500, 98420, 98360, 98320, 98280, 98210, 98230, 98240, 98350, 
    98440, 98460, 98590, 98670, 98830, 98990, 99140, 99240, 99290, 99420, 
    99480, 99510, 99490, 99450, 99520, 99450, 99560, 99700, 99740, 99800, 
    99870, 99950, 100050, 100140, 100230, 100360, 100470, 100540, 100630, 
    100710, 100820, 100870, 100980, 101170, 101280, 101400, 101530, 101610, 
    101680, 101740, 101790, 101870, 101930, 101970, 102000, 102050, 102030, 
    101990, 101970, 101930, 101910, 101860, 101810, 101780, 101740, 101680, 
    101620, 101570, 101460, 101390, 101300, 101240, 101190, 101140, 101100, 
    101060, 101020, 100970, 100850, 100790, 100760, 100720, 100710, 100720, 
    100720, 100660, 100690, 100680, 100670, 100630, 100660, 100620, 100620, 
    100630, 100660, 100590, 100540, 100590, 100660, 100670, 100670, 100670, 
    100640, 100600, 100610, 100640, 100670, 100660, 100660, 100700, 100750, 
    100740, 100750, 100770, 100760, 100750, 100740, 100750, 100720, 100720, 
    100700, 100690, 100740, 100770, 100800, 100810, 100780, 100750, 100750, 
    100750, 100730, 100750, 100740, 100740, 100790, 100800, 100820, 100820, 
    100800, 100760, 100720, 100690, 100700, 100690, 100660, 100670, 100640, 
    100650, 100630, 100620, 100610, 100600, 100590, 100570, 100550, 100510, 
    100460, 100430, 100390, 100350, 100310, 100290, 100230, 100200, 100120, 
    100090, 100020, 99970, 99930, 99860, 99820, 99780, 99760, 99670, 99550, 
    99460, 99390, 99280, 99180, 99370, 98930, 98780, 98700, 98630, 98530, 
    98440, 98490, 98550, 98610, 98640, 98690, 98760, 98840, 98840, 98850, 
    98980, 99040, 99020, 98980, 99010, 99070, 99080, 99150, 99240, 99260, 
    99290, 99360, 99400, 99380, 99440, 99620, 99650, 99650, 99750, 99850, 
    99810, 99790, 99850, 99950, 100070, 100240, 100340, 100280, 100300, 
    100340, 100280, 100310, 100300, 100280, 100270, 100250, 100220, 100170, 
    100140, 100100, 100080, 100040, 100000, 99960, 99910, 99880, 99850, 
    99830, 99790, 99730, 99710, 99750, 99760, 99760, 99740, 99730, 99720, 
    99670, 99670, 99640, 99640, 99660, 99640, 99620, 99590, 99560, 99520, 
    99460, 99460, 99410, 99400, 99380, 99410, 99480, 99530, 99540, 99470, 
    99480, 99480, 99550, 99690, 99580, 99540, 99590, 99600, 99560, 99540, 
    99470, 99430, 99410, 99380, 99420, 99440, 99480, 99500, 99510, 99550, 
    99570, 99620, 99660, 99710, 99680, 99750, 99810, 99870, 99880, 99940, 
    99980, 99980, 99980, 100090, 100110, 100170, 100200, 100220, 100220, 
    100270, 100300, 100380, 100450, 100500, 100540, 100630, 100700, 100760, 
    100800, 100890, 100950, 100980, 101020, 101070, 101130, 101200, 101240, 
    101300, 101330, 101370, 101410, 101450, 101470, 101480, 101510, 101530, 
    101560, 101590, 101630, 101650, 101660, 101680, 101700, 101710, 101690, 
    101700, 101790, 101860, 101890, 101890, 101860, 101870, 101830, 101770, 
    101750, 101780, 101820, 101820, 101800, 101820, 101850, 101850, 101830, 
    101810, 101770, 101750, 101740, 101690, 101630, 101570, 101550, 101510, 
    101460, 101390, 101290, 101270, 101260, 101200, 101120, 101080, 101010, 
    100980, 100940, 100880, 100840, 100830, 100800, 100730, 100680, 100630, 
    100610, 100680, 100660, 100630, 100580, 100560, 100510, 100490, 100460, 
    100430, 100440, 100430, 100450, 100450, 100460, 100470, 100460, 100480, 
    100500, 100540, 100560, 100560, 100610, 100630, 100630, 100650, 100670, 
    100690, 100700, 100730, 100760, 100770, 100790, 100800, 100770, 100780, 
    100800, 100860, 100860, 100850, 100840, 100850, 100870, 100860, 100930, 
    100960, 100980, 101030, 101060, 101100, 101100, 101130, 101200, 101240, 
    101310, 101350, 101350, 101390, 101410, 101430, 101490, 101520, 101530, 
    101500, 101530, 101550, 101590, 101600, 101610, 101580, 101580, 101570, 
    101570, 101550, 101570, 101570, 101540, 101530, 101510, 101490, 101480, 
    101450, 101430, 101390, 101340, 101340, 101380, 101330, 101290, 101280, 
    101300, 101280, 101240, 101250, 101230, 101210, 101210, 101210, 101200, 
    101190, 101170, 101100, 101070, 101020, 101010, 100910, 100830, 100770, 
    100710, 100620, 100630, 100590, 100460, 100460, 100400, 100370, 100360, 
    100370, 100460, 100480, 100590, 100660, 100730, 100780, 100800, 100870, 
    100940, 101020, 101080, 100970, 100930, 101040, 101100, 101170, 101150, 
    101140, 101160, 101190, 101240, 101260, 101300, 101310, 101330, 101360, 
    101390, 101420, 101400, 101400, 101410, 101440, 101470, 101470, 101490, 
    101530, 101540, 101560, 101570, 101570, 101590, 101610, 101600, 101600, 
    101630, 101670, 101680, 101680, 101660, 101630, 101600, 101560, 101510, 
    101380, 101280, 101220, 101170, 101050, 100890, 100850, 100830, 100840, 
    100780, 100810, 100740, 100730, 100750, 100730, 100770, 100790, 100820, 
    100860, 100910, 100980, 101030, 101060, 101100, 101130, 101190, 101230, 
    101290, 101370, 101420, 101490, 101520, 101560, 101560, 101570, 101570, 
    101580, 101580, 101590, 101600, 101600, 101580, 101570, 101570, 101570, 
    101550, 101530, 101470, 101400, 101350, 101290, 101250, 101200, 101160, 
    101130, 101060, 100970, 100840, 100710, 100600, 100460, 100290, 100100, 
    100000, 99880, 99670, 99460, 99290, 99160, 99000, 98810, 98630, 98330, 
    97920, 97550, 97310, 97380, 97300, 97390, 97480, 97560, 97560, 97460, 
    97480, 97460, 97390, 97340, 97310, 97300, 97370, 97400, 97460, 97520, 
    97610, 97730, 97840, 98010, 98180, 98390, 98580, 98750, 98920, 99060, 
    99180, 99300, 99420, 99520, 99570, 99700, 99830, 99960, 100090, 100180, 
    100280, 100330, 100450, 100530, 100660, 100670, 100720, 100750, 100810, 
    100830, 100820, 100810, 100810, 100750, 100650, 100550, 100440, 100390, 
    100290, 100200, 100000, 99940, 99870, 99810, 99700, 99680, 99640, 99680, 
    99720, 99690, 99690, 99640, 99690, 99660, 99650, 99650, 99640, 99660, 
    99650, 99610, 99570, 99550, 99490, 99430, 99310, 99230, 99130, 99030, 
    98850, 98710, 98570, 98540, 98400, 98350, 98280, 98250, 98180, 98060, 
    98000, 97990, 97970, 97940, 97890, 97830, 97770, 97760, 97760, 97780, 
    97760, 97770, 97790, 97830, 97850, 97890, 97970, 98000, 98020, 98050, 
    98090, 98110, 98110, 98140, 98170, 98160, 98160, 98150, 98160, 98150, 
    98140, 98130, 98110, 98110, 98090, 98080, 98030, 98020, 98020, 97970, 
    97950, 97900, 97870, 97840, 97790, 97740, 97720, 97690, 97650, 97620, 
    97620, 97610, 97580, 97570, 97540, 97520, 97490, 97530, 97520, 97530, 
    97550, 97580, 97600, 97650, 97680, 97710, 97730, 97760, 97790, 97830, 
    97880, 97930, 97980, 98030, 98080, 98130, 98130, 98130, 98150, 98150, 
    98180, 98180, 98180, 98180, 98210, 98200, 98190, 98190, 98190, 98210, 
    98200, 98180, 98180, 98210, 98230, 98230, 98260, 98280, 98300, 98320, 
    98340, 98370, 98380, 98380, 98400, 98420, 98460, 98510, 98530, 98520, 
    98520, 98550, 98580, 98560, 98570, 98570, 98570, 98560, 98570, 98560, 
    98560, 98560, 98580, 98590, 98610, 98620, 98630, 98640, 98670, 98690, 
    98710, 98760, 98790, 98840, 98890, 98950, 99000, 99060, 99100, 99170, 
    99230, 99280, 99370, 99410, 99470, 99530, 99580, 99630, 99710, 99790, 
    99840, 99910, 99960, 100020, 100050, 100130, 100170, 100200, 100260, 
    100340, 100360, 100370, 100420, 100450, 100460, 100490, 100520, 100530, 
    100540, 100550, 100550, 100550, 100520, 100530, 100530, 100530, 100510, 
    100510, 100510, 100520, 100510, 100500, 100510, 100520, 100470, 100420, 
    100390, 100390, 100310, 100230, 100150, 100150, 100060, 100070, 99980, 
    99770, 99750, 99630, 99400, 99380, 99350, 99260, 99160, 99090, 99070, 
    99100, 99050, 99000, 98970, 98960, 98980, 99020, 99050, 99110, 99160, 
    99230, 99300, 99340, 99440, 99480, 99560, 99570, 99630, 99640, 99670, 
    99710, 99740, 99780, 99770, 99770, 99830, 99860, 99840, 99850, 99830, 
    99830, 99780, 99780, 99710, 99730, 99730, 99730, 99720, 99700, 99690, 
    99660, 99710, 99760, 99760, 99730, 99810, 99880, 99870, 99890, 99890, 
    99810, 99770, 99760, 99750, 99710, 99620, 99520, 99480, 99400, 99270, 
    99240, 99120, 99090, 99090, 99050, 99000, 98960, 98900, 98950, 98980, 
    99040, 99010, 99010, 99060, 99130, 99200, 99250, 99320, 99390, 99420, 
    99400, 99470, 99540, 99580, 99620, 99640, 99650, 99660, 99670, 99750, 
    99680, 99640, 99690, 99650, 99730, 99750, 99830, 99880, 99860, 99860, 
    99930, 99990, 100030, 100120, 100200, 100160, 100110, 100130, 100220, 
    100310, 100420, 100480, 100550, 100620, 100660, 100730, 100770, 100800, 
    100820, 100830, 100800, 100820, 100860, 100860, 100860, 100830, 100800, 
    100830, 100830, 100820, 100800, 100780, 100810, 100820, 100860, 100850, 
    100770, 100790, 100750, 100770, 100750, 100720, 100680, 100710, 100710, 
    100730, 100710, 100630, 100590, 100550, 100520, 100530, 100520, 100530, 
    100490, 100480, 100490, 100480, 100470, 100410, 100360, 100340, 100310, 
    100310, 100300, 100300, 100330, 100330, 100340, 100350, 100340, 100360, 
    100370, 100370, 100370, 100380, 100420, 100410, 100400, 100400, 100420, 
    100420, 100440, 100430, 100440, 100470, 100480, 100460, 100500, 100500, 
    100520, 100540, 100580, 100610, 100640, 100650, 100670, 100660, 100670, 
    100680, 100680, 100670, 100670, 100690, 100690, 100690, 100710, 100730, 
    100740, 100760, 100760, 100760, 100770, 100770, 100790, 100820, 100850, 
    100880, 100890, 100890, 100930, 100930, 100960, 100940, 100980, 101000, 
    100990, 100990, 101050, 101090, 101110, 101110, 101110, 101130, 101150, 
    101150, 101130, 101130, 101130, 101150, 101170, 101190, 101220, 101250, 
    101310, 101320, 101300, 101240, 101240, 101210, 101210, 101170, 101160, 
    101140, 101110, 101090, 101060, 101000, 100930, 100920, 100870, 100840, 
    100820, 100810, 100780, 100750, 100690, 100660, 100630, 100570, 100540, 
    100500, 100470, 100460, 100440, 100430, 100440, 100400, 100440, 100470, 
    100480, 100500, 100550, 100550, 100570, 100610, 100650, 100670, 100710, 
    100780, 100780, 100810, 100830, 100880, 100890, 100940, 100970, 100980, 
    100960, 100980, 101010, 101080, 101130, 101090, 101180, 101270, 101300, 
    101310, 101310, 101320, 101370, 101370, 101380, 101400, 101390, 101360, 
    101330, 101340, 101390, 101400, 101410, 101430, 101420, 101380, 101320, 
    101400, 101400, 101380, 101350, 101350, 101380, 101400, 101430, 101460, 
    101470, 101480, 101560, 101600, 101610, 101620, 101600, 101550, 101550, 
    101580, 101620, 101770, 101800, 101820, 101810, 101820, 101840, 101810, 
    101850, 101860, 101890, 101920, 101990, 101990, 102000, 102040, 102030, 
    102070, 102060, 102060, 102070, 102080, 102090, 102090, 102070, 102040, 
    102060, 102070, 102070, 102050, 102020, 101960, 101960, 101950, 101950, 
    101870, 101830, 101800, 101750, 101760, 101790, 101810, 101840, 101830, 
    101800, 101820, 101840, 101850, 101840, 101840, 101830, 101830, 101840, 
    101850, 101810, 101790, 101750, 101740, 101730, 101720, 101710, 101690, 
    101690, 101690, 101680, 101690, 101670, 101670, 101660, 101650, 101620, 
    101640, 101610, 101600, 101580, 101590, 101550, 101550, 101510, 101480, 
    101470, 101480, 101470, 101460, 101440, 101440, 101430, 101450, 101440, 
    101450, 101470, 101490, 101480, 101500, 101520, 101520, 101540, 101540, 
    101550, 101550, 101600, 101620, 101630, 101660, 101670, 101690, 101700, 
    101710, 101720, 101750, 101760, 101800, 101860, 101880, 101900, 101930, 
    101970, 101990, 102020, 102020, 102040, 102040, 102060, 102100, 102110, 
    102140, 102170, 102190, 102220, 102250, 102260, 102290, 102300, 102310, 
    102330, 102350, 102380, 102380, 102380, 102380, 102390, 102400, 102400, 
    102380, 102370, 102360, 102350, 102340, 102330, 102310, 102280, 102280, 
    102270, 102250, 102220, 102200, 102180, 102180, 102160, 102140, 102150, 
    102130, 102130, 102090, 102070, 102040, 101970, 101880, 101830, 101770, 
    101720, 101670, 101650, 101650, 101660, 101740, 101740, 101760, 101790, 
    101810, 101850, 101860, 101790, 101970, 101890, 102090, 102090, 102070, 
    102080, 102030, 101980, 102010, 102040, 102030, 102070, 102100, 102040, 
    102080, 102070, 102060, 102040, 102010, 102020, 101980, 101950, 101980, 
    101970, 101940, 101860, 101860, 101750, 101700, 101700, 101620, 101590, 
    101640, 101610, 101590, 101640, 101650, 101730, 101760, 101770, 101780, 
    101790, 101830, 101860, 101890, 101890, 101890, 101880, 101900, 101920, 
    101950, 101990, 102030, 102040, 102040, 102060, 102060, 102080, 102060, 
    102080, 102090, 102100, 102110, 102120, 102140, 102140, 102140, 102170, 
    102170, 102250, 102190, 102200, 102210, 102230, 102230, 102260, 102260, 
    102270, 102270, 102260, 102250, 102230, 102210, 102170, 102160, 102210, 
    102190, 102170, 102150, 102140, 102130, 102110, 102090, 102080, 102060, 
    102030, 102050, 102030, 102010, 102000, 101990, 101950, 101960, 101930, 
    101920, 101890, 101860, 101850, 101840, 101830, 101850, 101850, 101860, 
    101890, 101900, 101900, 101910, 101920, 101940, 101950, 101960, 101890, 
    101940, 101930, 101920, 101890, 101900, 101830, 101700, 101580, 101580, 
    101590, 101600, 101620, 101620, 101620, 101610, 101640, 101650, 101640, 
    101730, 101760, 101720, 101710, 101750, 101740, 101750, 101710, 101640, 
    101630, 101660, 101640, 101670, 101690, 101740, 101700, 101650, 101610, 
    101610, 101610, 101600, 101600, 101550, 101500, 101480, 101470, 101560, 
    101580, 101590, 101630, 101640, 101670, 101690, 101690, 101710, 101710, 
    101720, 101740, 101780, 101770, 101790, 101840, 101870, 101890, 101870, 
    101870, 101880, 101890, 101860, 101860, 101880, 101920, 101910, 101920, 
    101910, 101880, 101860, 101850, 101790, 101680, 101670, 101710, 101740, 
    101730, 101720, 101710, 101710, 101710, 101680, 101660, 101640, 101610, 
    101590, 101580, 101560, 101550, 101530, 101520, 101540, 101510, 101440, 
    101440, 101420, 101420, 101430, 101400, 101380, 101390, 101400, 101360, 
    101330, 101290, 101290, 101270, 101270, 101270, 101250, 101250, 101210, 
    101220, 101240, 101260, 101310, 101300, 101300, 101310, 101300, 101340, 
    101360, 101360, 101370, 101370, 101360, 101340, 101320, 101340, 101330, 
    101350, 101330, 101300, 101270, 101270, 101240, 101220, 101220, 101220, 
    101230, 101250, 101260, 101300, 101320, 101310, 101340, 101340, 101340, 
    101390, 101430, 101440, 101460, 101490, 101510, 101490, 101520, 101530, 
    101540, 101540, 101560, 101580, 101610, 101620, 101610, 101640, 101630, 
    101620, 101600, 101590, 101560, 101550, 101530, 101500, 101420, 101350, 
    101280, 101200, 101120, 101040, 101000, 100930, 100860, 100820, 100830, 
    100930, 100910, 100940, 100960, 100970, 101030, 101100, 101140, 101140, 
    101180, 101190, 101200, 101210, 101190, 101200, 101150, 101140, 101110, 
    101050, 101040, 100980, 100920, 100900, 100840, 100800, 100770, 100730, 
    100710, 100650, 100690, 100700, 100700, 100720, 100760, 100770, 100800, 
    100790, 100830, 100850, 100830, 100860, 100860, 100890, 100890, 100930, 
    100950, 101020, 101160, 101250, 101390, 101510, 101590, 101680, 101770, 
    101820, 101940, 102010, 102120, 102210, 102260, 102380, 102460, 102570, 
    102640, 102670, 102750, 102790, 102850, 102890, 102920, 102970, 103040, 
    103060, 103070, 103130, 103170, 103180, 103200, 103200, 103190, 103200, 
    103190, 103180, 103150, 103140, 103100, 103090, 103040, 103010, 102960, 
    102910, 102880, 102830, 102790, 102740, 102660, 102620, 102590, 102560, 
    102530, 102480, 102420, 102380, 102320, 102290, 102170, 102150, 102110, 
    102110, 102110, 102120, 102120, 102100, 102090, 102090, 102090, 102100, 
    102150, 102210, 102260, 102280, 102330, 102340, 102370, 102390, 102440, 
    102460, 102470, 102460, 102460, 102470, 102490, 102530, 102550, 102570, 
    102590, 102600, 102630, 102630, 102600, 102570, 102610, 102600, 102600, 
    102570, 102530, 102480, 102450, 102350, 102270, 102190, 102090, 102000, 
    101890, 101780, 101670, 101610, 101520, 101390, 101310, 101320, 101230, 
    101210, 101200, 101170, 101100, 101080, 101070, 101080, 101050, 101080, 
    101100, 101130, 101170, 101180, 101250, 101290, 101330, 101390, 101460, 
    101520, 101550, 101580, 101630, 101640, 101670, 101700, 101760, 101800, 
    101830, 101860, 101890, 101920, 101910, 101960, 102030, 102130, 102190, 
    102210, 102230, 102240, 102250, 102280, 102320, 102320, 102340, 102350, 
    102370, 102380, 102340, 102350, 102340, 102290, 102270, 102240, 102260, 
    102270, 102270, 102290, 102310, 102320, 102290, 102310, 102400, 102310, 
    102310, 102310, 102370, 102350, 102350, 102390, 102320, 102400, 102450, 
    102400, 102430, 102500, 102670, 102610, 102580, 102600, 102640, 102660, 
    102740, 102750, 102750, 102760, 102790, 102840, 102870, 102880, 102900, 
    102930, 102930, 102950, 102960, 102930, 102930, 102900, 102940, 102940, 
    102960, 102970, 102990, 102990, 103010, 103010, 103020, 103040, 103080, 
    103080, 103080, 103080, 103050, 103040, 103030, 103030, 103010, 102990, 
    102990, 102960, 102940, 102920, 102920, 102910, 102900, 102880, 102880, 
    102880, 102910, 102960, 103000, 103040, 103060, 103110, 103140, 103180, 
    103200, 103220, 103250, 103280, 103300, 103300, 103330, 103340, 103350, 
    103350, 103350, 103340, 103340, 103350, 103330, 103350, 103350, 103340, 
    103330, 103310, 103300, 103290, 103280, 103260, 103220, 103220, 103190, 
    103170, 103190, 103180, 101350, 103140, 103140, 103130, 103110, 103100, 
    103080, 103070, 103050, 103080, 103080, 103100, 103100, 103110, 103090, 
    103080, 103060, 103050, 103060, 103060, 103040, 103050, 103080, 103080, 
    103080, 103060, 103070, 103060, 103040, 103040, 103020, 103020, 103040, 
    103050, 103070, 103080, 103090, 103090, 103090, 103070, 103070, 103050, 
    103040, 103020, 103010, 103010, 103010, 102990, 102990, 102970, 102940, 
    102910, 102910, 102900, 102880, 102870, 102880, 102880, 102890, 102890, 
    102910, 102930, 102910, 102920, 102930, 102930, 102930, 102910, 102890, 
    102880, 102900, 102870, 102870, 102850, 102830, 102810, 102790, 102780, 
    102740, 102740, 102730, 102750, 102750, 102740, 102730, 102740, 102710, 
    102690, 102680, 102660, 102610, 102540, 102470, 102410, 102340, 102290, 
    102220, 102160, 102060, 101970, 101900, 101820, 101740, 101640, 101570, 
    101510, 101420, 101360, 101280, 101230, 101200, 101240, 101290, 101340, 
    101380, 101420, 101430, 101430, 101490, 101520, 101560, 101590, 101560, 
    101550, 101570, 101580, 101580, 101560, 101560, 101540, 101530, 101540, 
    101560, 101540, 101510, 101500, 101500, 101520, 101550, 101530, 101510, 
    101550, 101520, 101590, 101620, 101670, 101770, 101780, 101770, 101770, 
    101820, 101830, 101870, 101840, 101900, 102060, 102080, 102080, 102030, 
    102050, 102140, 102170, 102180, 102180, 102190, 102200, 102190, 102190, 
    102230, 102190, 102210, 102210, 102200, 102190, 102190, 102190, 102190, 
    102210, 102220, 102220, 102200, 102220, 102220, 102230, 102230, 102210, 
    102200, 102190, 102150, 102140, 102150, 102150, 102140, 102120, 102120, 
    102110, 102120, 102110, 102090, 102090, 102090, 102100, 102100, 102130, 
    102140, 102130, 102120, 102110, 102110, 102100, 102080, 102080, 102070, 
    102060, 102050, 102050, 102030, 102040, 102010, 102030, 102030, 102030, 
    102010, 101970, 101960, 101970, 101960, 101980, 101980, 101990, 101960, 
    101940, 101920, 101880, 101870, 101840, 101810, 101810, 101770, 101740, 
    101700, 101680, 101640, 101620, 101580, 101540, 101460, 101400, 101350, 
    101310, 101290, 101260, 101220, 101170, 101130, 101100, 101040, 101000, 
    100950, 100880, 100840, 100820, 100780, 100740, 100710, 100680, 100700, 
    100690, 100670, 100640, 100620, 100600, 100570, 100540, 100520, 100510, 
    100500, 100490, 100500, 100460, 100420, 100370, 100330, 100320, 100290, 
    100280, 100280, 100300, 100320, 100350, 100370, 100390, 100390, 100410, 
    100440, 100460, 100480, 100510, 100540, 100580, 100630, 100650, 100680, 
    100700, 100720, 100750, 100760, 100790, 100800, 100820, 100830, 100850, 
    100870, 100890, 100900, 100920, 100930, 100950, 100970, 100970, 100980, 
    100980, 101010, 101010, 101030, 101050, 101060, 101090, 101110, 101120, 
    101160, 101200, 101220, 101220, 101230, 101210, 101220, 101200, 101190, 
    101170, 101130, 101100, 101090, 101050, 101100, 101140, 101160, 101180, 
    101190, 101190, 101220, 101240, 101240, 101240, 101230, 101250, 101250, 
    101240, 101240, 101240, 101230, 101250, 101260, 101260, 101270, 101280, 
    101290, 101310, 101300, 101320, 101350, 101370, 101410, 101430, 101460, 
    101480, 101520, 101530, 101540, 101540, 101550, 101550, 101570, 101600, 
    101640, 101680, 101720, 101750, 101780, 101800, 101830, 101850, 101900, 
    101950, 101990, 102020, 102060, 102110, 102130, 102160, 102190, 102190, 
    102220, 102230, 102250, 102250, 102260, 102270, 102290, 102310, 102310, 
    102320, 102320, 102290, 102260, 102230, 102250, 102240, 102230, 102230, 
    102200, 102230, 102220, 102190, 102170, 102120, 102090, 102070, 102010, 
    101990, 101970, 101930, 101910, 101820, 101720, 101700, 101630, 101590, 
    101510, 101390, 101330, 101320, 101260, 101200, 101220, 101190, 101220, 
    101200, 101170, 101140, 101150, 101180, 101190, 101220, 101260, 101300, 
    101340, 101380, 101390, 101410, 101440, 101430, 101450, 101480, 101460, 
    101490, 101520, 101560, 101520, 101560, 101590, 101640, 101670, 101740, 
    101800, 101800, 101810, 101850, 101930, 101960, 102020, 101990, 101990, 
    102020, 102010, 102080, 102060, 102090, 102130, 102140, 102180, 102190, 
    102210, 102210, 102250, 102320, 102320, 102360, 102390, 102430, 102470, 
    102500, 102530, 102550, 102590, 102610, 102640, 102680, 102700, 102730, 
    102750, 102760, 102780, 102800, 102870, 102880, 102900, 102940, 102970, 
    102990, 103010, 103040, 103040, 103050, 103100, 103110, 103100, 103110, 
    103090, 103080, 103070, 103050, 103070, 103050, 103030, 103030, 103000, 
    102980, 102990, 102980, 102950, 102940, 102930, 102910, 102890, 102860, 
    102830, 102810, 102790, 102760, 102710, 102660, 102620, 102580, 102560, 
    102510, 102480, 102430, 102400, 102370, 102340, 102360, 102320, 102310, 
    102320, 102290, 102290, 102300, 102310, 102300, 102300, 102320, 102310, 
    102320, 102330, 102340, 102350, 102360, 102380, 102390, 102400, 102420, 
    102440, 102450, 102460, 102450, 102460, 102490, 102490, 102490, 102510, 
    102520, 102510, 102540, 102530, 102540, 102540, 102550, 102530, 102520, 
    102480, 102460, 102440, 102430, 102420, 102410, 102410, 102370, 102370, 
    102350, 102370, 102350, 102360, 102350, 102330, 102340, 102360, 102340, 
    102320, 102320, 102300, 102290, 102300, 102290, 102270, 102240, 102250, 
    102240, 102210, 102220, 102220, 102230, 102220, 102220, 102230, 102220, 
    102220, 102210, 102210, 102210, 102220, 102230, 102250, 102220, 102200, 
    102200, 102190, 102160, 102140, 102150, 102150, 102120, 102120, 102120, 
    102140, 102100, 102050, 102060, 102080, 102100, 102090, 102090, 102110, 
    102090, 102090, 102070, 102080, 102080, 102080, 102080, 102100, 102110, 
    102130, 102170, 102200, 102220, 102240, 102290, 102350, 102380, 102420, 
    102470, 102530, 102600, 102650, 102710, 102740, 102760, 102800, 102830, 
    102850, 102880, 102900, 102920, 102920, 102930, 102940, 102930, 102950, 
    102930, 102900, 102910, 102890, 102880, 102870, 102830, 102840, 102820, 
    102810, 102790, 102750, 102730, 102730, 102710, 102650, 102620, 102570, 
    102540, 102580, 102550, 102510, 102520, 102460, 102450, 102420, 102390, 
    102350, 102360, 102360, 102360, 102410, 102460, 102460, 102490, 102500, 
    102500, 102460, 102440, 102410, 102340, 102290, 102230, 102150, 102070, 
    101950, 101830, 101760, 101670, 101620, 101590, 101550, 101530, 101570, 
    101590, 101570, 101570, 101580, 101590, 101620, 101590, 101580, 101590, 
    101580, 101550, 101520, 101480, 101430, 101390, 101380, 101340, 101310, 
    101310, 101270, 101220, 101150, 101120, 101080, 101050, 101010, 101020, 
    101020, 101010, 101010, 101020, 101010, 100990, 100980, 100960, 100960, 
    100920, 100920, 100900, 100850, 100820, 100800, 100830, 100810, 100790, 
    100760, 100700, 100650, 100630, 100660, 100620, 100590, 100530, 100540, 
    100540, 100470, 100430, 100380, 100220, 100220, 100200, 100190, 100160, 
    100130, 100110, 100030, 99960, 99910, 99870, 99830, 99820, 99830, 99880, 
    99930, 99990, 100020, 100040, 100120, 100170, 100220, 100290, 100310, 
    100280, 100340, 100390, 100400, 100430, 100450, 100460, 100470, 100480, 
    100490, 100490, 100490, 100480, 100480, 100500, 100480, 100500, 100510, 
    100510, 100480, 100480, 100480, 100480, 100440, 100430, 100430, 100430, 
    100420, 100430, 100420, 100440, 100450, 100430, 100430, 100440, 100460, 
    100480, 100480, 100510, 100520, 100550, 100580, 100620, 100630, 100640, 
    100650, 100660, 100690, 100690, 100680, 100690, 100700, 100720, 100740, 
    100740, 100720, 100700, 100680, 100690, 100690, 100680, 100690, 100680, 
    100690, 100710, 100710, 100720, 100720, 100720, 100720, 100710, 100730, 
    100720, 100710, 100680, 100680, 100700, 100690, 100720, 100730, 100720, 
    100710, 100700, 100690, 100680, 100670, 100670, 100680, 100700, 100710, 
    100710, 100710, 100720, 100710, 100730, 100720, 100710, 100710, 100700, 
    100690, 100690, 100680, 100670, 100680, 100670, 100640, 100600, 100580, 
    100560, 100530, 100520, 100520, 100530, 100530, 100500, 100480, 100470, 
    100460, 100440, 100440, 100440, 100450, 100460, 100470, 100500, 100500, 
    100520, 100530, 100550, 100570, 100570, 100600, 100630, 100630, 100670, 
    100680, 100730, 100760, 100770, 100770, 100800, 100800, 100810, 100830, 
    100840, 100830, 100830, 100850, 100850, 100850, 100870, 100870, 100870, 
    100880, 100880, 100870, 100870, 100890, 100910, 100910, 100920, 100920, 
    100940, 100940, 100950, 100960, 100970, 100960, 100980, 100990, 100950, 
    100960, 100960, 100970, 100990, 100980, 100970, 100970, 100950, 100960, 
    100960, 100940, 100970, 100970, 100970, 100970, 100990, 101020, 101020, 
    101010, 101000, 101000, 101010, 101010, 101020, 101030, 101020, 101010, 
    101020, 101000, 101010, 101020, 101020, 101030, 101010, 100990, 101000, 
    101010, 101030, 101040, 101040, 101040, 101020, 101010, 101020, 100990, 
    101010, 101010, 101020, 101010, 100990, 101000, 101020, 101030, 101030, 
    101030, 101020, 101020, 101000, 101010, 101020, 101030, 101040, 101040, 
    101040, 101040, 101050, 101070, 101060, 101060, 101050, 101050, 101050, 
    101050, 101070, 101080, 101090, 101080, 101070, 101060, 101060, 101060, 
    101040, 101020, 101040, 101040, 101050, 101070, 101070, 101040, 101020, 
    100980, 100970, 100970, 100960, 100940, 100920, 100890, 100890, 100860, 
    100840, 100820, 100790, 100770, 100740, 100730, 100690, 100680, 100670, 
    100660, 100680, 100680, 100670, 100650, 100640, 100610, 100600, 100570, 
    100560, 100560, 100550, 100550, 100510, 100460, 100440, 100400, 100370, 
    100340, 100340, 100330, 100360, 100320, 100320, 100340, 100360, 100350, 
    100360, 100360, 100360, 100330, 100330, 100330, 100340, 100320, 100330, 
    100340, 100370, 100370, 100390, 100400, 100410, 100440, 100430, 100460, 
    100450, 100460, 100470, 100480, 100470, 100440, 100440, 100460, 100460, 
    100440, 100410, 100380, 100330, 100280, 100240, 100210, 100250, 100160, 
    100140, 100100, 100090, 100070, 100080, 100090, 100090, 100100, 100140, 
    100180, 100210, 100250, 100320, 100360, 100410, 100460, 100510, 100550, 
    100610, 100630, 100650, 100720, 100790, 100850, 100930, 100990, 101040, 
    101060, 101090, 101130, 101140, 101180, 101210, 101260, 101290, 101340, 
    101370, 101390, 101400, 101400, 101400, 101400, 101390, 101360, 101390, 
    101410, 101470, 101500, 101530, 101540, 101540, 101490, 101490, 101480, 
    101490, 101520, 101500, 101500, 101500, 101520, 101570, 101620, 101650, 
    101650, 101590, 101600, 101560, 101580, 101600, 101630, 101660, 101660, 
    101640, 101610, 101600, 101600, 101590, 101590, 101580, 101560, 101550, 
    101580, 101600, 101590, 101590, 101590, 101600, 101590, 101600, 101580, 
    101580, 101590, 101590, 101580, 101600, 101600, 101590, 101590, 101580, 
    101570, 101580, 101560, 101550, 101530, 101510, 101530, 101510, 101530, 
    101520, 101520, 101490, 101460, 101430, 101410, 101360, 101330, 101310, 
    101270, 101250, 101210, 101170, 101110, 101090, 101020, 100940, 100920, 
    100880, 100810, 100780, 100750, 100700, 100660, 100640, 100600, 100550, 
    100490, 100440, 100370, 100310, 100290, 100250, 100200, 100160, 100170, 
    100150, 100130, 100120, 100100, 100090, 100100, 100110, 100100, 100110, 
    100130, 100160, 100180, 100210, 100230, 100250, 100280, 100300, 100290, 
    100290, 100330, 100380, 100420, 100450, 100490, 100500, 100510, 100510, 
    100520, 100550, 100550, 100570, 100590, 100580, 100590, 100660, 100720, 
    100770, 100780, 100780, 100840, 100840, 100830, 100860, 100880, 100870, 
    100890, 100930, 100910, 100910, 100910, 100900, 100890, 100860, 100870, 
    100860, 100880, 100900, 100880, 100900, 100880, 100880, 100840, 100810, 
    100770, 100730, 100700, 100650, 100590, 100530, 100440, 100350, 100300, 
    100180, 100100, 100050, 99970, 99920, 99810, 99750, 99740, 99660, 99630, 
    99620, 99610, 99630, 99640, 99680, 99730, 99750, 99800, 99870, 99890, 
    99900, 99950, 99990, 100020, 100050, 100090, 100120, 100150, 100190, 
    100230, 100270, 100320, 100370, 100420, 100440, 100500, 100560, 100580, 
    100590, 100610, 100640, 100670, 100690, 100720, 100730, 100740, 100750, 
    100790, 100800, 100800, 100790, 100790, 100780, 100790, 100810, 100820, 
    100840, 100860, 100890, 100890, 100920, 100930, 100940, 100950, 100960, 
    100990, 101000, 101010, 101030, 101040, 101060, 101060, 101080, 101090, 
    101090, 101090, 101070, 101080, 101100, 101090, 101110, 101100, 101100, 
    101110, 101140, 101130, 101120, 101120, 101110, 101110, 101080, 101050, 
    101030, 101020, 101020, 101020, 101010, 100990, 100990, 100970, 100970, 
    100970, 100970, 100980, 100990, 100990, 100990, 101010, 101020, 101030, 
    101040, 101040, 101020, 101030, 101050, 101080, 101110, 101090, 101080, 
    101110, 101090, 101080, 101100, 101090, 101020, 101070, 101060, 101030, 
    100990, 100950, 100910, 100870, 100810, 100670, 100540, 100440, 100320, 
    100270, 100120, 99940, 99860, 99650, 99640, 99520, 99490, 99550, 99550, 
    99580, 99590, 99640, 99700, 99750, 99810, 99850, 99870, 99880, 99910, 
    99990, 100050, 100070, 100120, 100170, 100250, 100300, 100340, 100400, 
    100480, 100580, 100640, 100700, 100770, 100860, 100960, 101050, 101100, 
    101170, 101240, 101300, 101370, 101440, 101480, 101490, 101500, 101510, 
    101560, 101590, 101610, 101600, 101600, 101600, 101570, 101540, 101570, 
    101540, 101500, 101460, 101410, 101410, 101340, 101260, 101170, 101070, 
    101010, 100880, 100810, 100700, 100560, 100480, 100300, 100400, 100340, 
    100380, 100350, 100380, 100410, 100430, 100460, 100500, 100560, 100600, 
    100640, 100670, 100710, 100710, 100730, 100790, 100850, 100840, 100840, 
    100840, 100840, 100840, 100860, 100830, 100870, 100890, 100910, 100930, 
    100950, 101040, 101050, 101090, 101170, 101170, 101210, 101260, 101300, 
    101330, 101320, 101380, 101390, 101390, 101430, 101410, 101380, 101410, 
    101410, 101380, 101350, 101330, 101320, 101320, 101330, 101310, 101290, 
    101210, 101140, 101020, 101020, 100940, 100910, 100890, 100810, 100770, 
    100750, 100670, 100660, 100610, 100610, 100650, 100640, 100660, 100660, 
    100650, 100680, 100690, 100710, 100730, 100780, 100850, 100900, 100910, 
    100880, 100890, 100970, 101000, 101020, 101020, 101030, 101030, 100980, 
    100960, 100910, 100820, 100730, 100680, 100670, 100650, 100630, 100630, 
    100610, 100630, 100660, 100670, 100700, 100730, 100750, 100780, 100810, 
    100870, 100910, 100980, 101020, 101060, 101140, 101200, 101260, 101310, 
    101350, 101410, 101470, 101510, 101570, 101640, 101690, 101740, 101780, 
    101840, 101870, 101890, 101910, 101910, 101830, 101890, 101890, 101870, 
    101870, 101850, 101820, 101780, 101730, 101650, 101590, 101560, 101470, 
    101420, 101370, 101290, 101200, 101150, 101090, 101020, 101030, 101030, 
    101060, 101070, 101130, 101200, 101260, 101350, 101410, 101490, 101550, 
    101600, 101600, 101650, 101640, 101740, 101760, 101810, 101820, 101860, 
    101850, 101850, 101830, 101820, 101790, 101770, 101760, 101750, 101700, 
    101680, 101670, 101670, 101650, 101640, 101670, 101630, 101600, 101570, 
    101540, 101510, 101500, 101490, 101460, 101440, 101420, 101410, 101350, 
    101390, 101370, 101380, 101360, 101350, 101330, 101300, 101320, 101330, 
    101380, 101410, 101440, 101460, 101470, 101480, 101510, 101530, 101550, 
    101560, 101590, 101610, 101610, 101620, 101660, 101660, 101670, 101670, 
    101650, 101640, 101630, 101650, 101610, 101590, 101580, 101560, 101550, 
    101510, 101480, 101450, 101420, 101370, 101350, 101310, 101280, 101280, 
    101250, 101200, 101180, 101150, 101110, 101040, 101010, 100990, 100980, 
    100930, 100870, 100870, 100820, 100810, 100800, 100770, 100740, 100690, 
    100680, 100630, 100600, 100570, 100540, 100540, 100530, 100520, 100500, 
    100500, 100500, 100490, 100470, 100490, 100510, 100520, 100530, 100540, 
    100580, 100620, 100610, 100630, 100650, 100670, 100690, 100720, 100710, 
    100730, 100770, 100750, 100780, 100750, 100750, 100870, 100920, 100930, 
    100940, 100910, 100910, 100920, 101040, 101060, 101050, 101070, 101110, 
    101160, 101170, 101140, 101210, 101220, 101270, 101310, 101340, 101360, 
    101390, 101330, 101320, 101320, 101340, 101320, 101320, 101310, 101280, 
    101290, 101280, 101270, 101260, 101250, 101240, 101230, 101190, 101200, 
    101190, 101180, 101170, 101170, 101180, 101150, 101130, 101130, 101140, 
    101130, 101100, 101050, 101010, 100950, 100890, 100870, 100870, 100850, 
    100850, 100830, 100810, 100750, 100740, 100710, 100680, 100660, 100660, 
    100690, 100690, 100730, 100740, 100740, 100740, 100700, 100720, 100750, 
    100800, 100780, 100740, 100770, 100780, 100820, 100850, 100860, 100850, 
    100850, 100830, 100820, 100810, 100780, 100800, 100790, 100780, 100790, 
    100780, 100790, 100790, 100780, 100740, 100740, 100740, 100750, 100750, 
    100750, 100760, 100770, 100800, 100820, 100840, 100830, 100840, 100820, 
    100850, 100860, 100880, 100900, 100930, 100970, 101000, 101020, 101040, 
    101010, 100990, 101000, 101000, 100990, 100970, 100970, 100980, 100980, 
    100950, 100980, 100990, 100980, 100980, 100980, 100980, 100980, 100990, 
    101020, 101030, 101050, 101040, 101060, 101050, 101050, 101040, 101040, 
    101040, 101040, 101060, 101060, 101090, 101120, 101150, 101170, 101200, 
    101200, 101210, 101210, 101220, 101220, 101210, 101210, 101220, 101230, 
    101230, 101220, 101220, 101230, 101200, 101200, 101200, 101190, 101190, 
    101160, 101210, 101220, 101230, 101250, 101280, 101290, 101310, 101330, 
    101340, 101370, 101400, 101430, 101470, 101490, 101520, 101540, 101590, 
    101600, 101610, 101630, 101630, 101640, 101650, 101680, 101710, 101730, 
    101730, 101750, 101770, 101770, 101790, 101780, 101780, 101760, 101750, 
    101730, 101730, 101710, 101710, 101710, 101700, 101690, 101680, 101670, 
    101670, 101640, 101620, 101610, 101610, 101600, 101600, 101610, 101630, 
    101630, 101660, 101660, 101650, 101640, 101640, 101600, 101590, 101590, 
    101600, 101600, 101620, 101610, 101610, 101620, 101600, 101590, 101590, 
    101590, 101610, 101650, 101700, 101760, 101790, 101810, 101860, 101870, 
    101900, 101920, 101930, 101950, 101960, 101980, 102000, 102030, 102060, 
    102080, 102110, 102120, 102140, 102150, 102160, 102160, 102200, 102210, 
    102230, 102260, 102270, 102260, 102240, 102220, 102230, 102200, 102200, 
    102180, 102160, 102190, 102180, 102160, 102160, 102120, 102070, 102050, 
    102010, 101990, 101970, 101950, 101960, 101950, 101960, 101960, 101940, 
    101960, 101950, 101940, 101940, 101940, 101950, 101950, 101940, 101940, 
    101940, 101940, 101930, 101930, 101910, 101870, 101850, 101840, 101820, 
    101830, 101840, 101800, 101830, 101840, 101810, 101790, 101750, 101720, 
    101700, 101680, 101630, 101620, 101590, 101540, 101500, 101470, 101430, 
    101390, 101360, 101330, 101290, 101280, 101260, 101230, 101230, 101210, 
    101210, 101200, 101160, 101120, 101080, 101070, 101070, 101020, 100980, 
    100970, 100970, 100950, 100920, 100880, 100850, 100870, 100790, 100750, 
    100790, 100770, 100740, 100760, 100750, 100670, 100670, 100620, 100610, 
    100600, 100570, 100560, 100520, 100510, 100470, 100400, 100360, 100310, 
    100220, 100150, 100130, 100120, 100090, 100000, 99960, 99910, 99850, 
    99850, 99810, 99710, 99710, 99690, 99680, 99630, 99560, 99530, 99470, 
    99400, 99300, 99380, 99420, 99440, 99400, 99360, 99330, 99310, 99280, 
    99240, 99190, 99180, 99180, 99170, 99140, 99140, 99150, 99150, 99170, 
    99200, 99240, 99210, 99260, 99260, 99240, 99280, 99320, 99350, 99360, 
    99380, 99410, 99430, 99450, 99450, 99430, 99460, 99480, 99510, 99530, 
    99570, 99540, 99610, 99660, 99670, 99700, 99690, 99730, 99770, 99840, 
    99910, 99960, 100000, 100080, 100150, 100240, 100300, 100350, 100380, 
    100380, 100390, 100380, 100380, 100390, 100390, 100390, 100360, 100330, 
    100320, 100320, 100340, 100360, 100360, 100390, 100460, 100510, 100540, 
    100570, 100590, 100570, 100590, 100640, 100660, 100680, 100620, 100710, 
    100770, 100800, 100800, 100800, 100830, 100910, 100900, 100920, 100930, 
    100940, 100960, 100980, 101030, 101040, 101080, 101090, 101080, 101060, 
    101030, 101040, 101010, 100980, 100960, 100950, 100950, 100960, 100970, 
    100960, 100960, 100950, 100950, 100950, 100950, 100900, 100860, 100840, 
    100820, 100780, 100760, 100750, 100750, 100750, 100770, 100790, 100790, 
    100790, 100800, 100820, 100830, 100810, 100840, 100850, 100850, 100850, 
    100850, 100840, 100790, 100750, 100720, 100710, 100660, 100640, 100600, 
    100570, 100530, 100490, 100450, 100460, 100440, 100430, 100400, 100360, 
    100330, 100320, 100330, 100330, 100340, 100350, 100350, 100330, 100300, 
    100290, 100280, 100300, 100280, 100240, 100290, 100310, 100340, 100350, 
    100400, 100490, 100600, 100690, 100760, 100830, 100880, 100940, 101020, 
    101100, 101160, 101220, 101270, 101310, 101340, 101360, 101380, 101400, 
    101440, 101460, 101500, 101530, 101560, 101590, 101620, 101620, 101630, 
    101610, 101620, 101620, 101630, 101630, 101620, 101630, 101670, 101690, 
    101720, 101740, 101750, 101760, 101770, 101770, 101780, 101780, 101790, 
    101780, 101780, 101790, 101780, 101770, 101770, 101750, 101730, 101740, 
    101750, 101770, 101770, 101780, 101770, 101750, 101760, 101720, 101710, 
    101670, 101640, 101610, 101610, 101560, 101530, 101490, 101470, 101460, 
    101460, 101420, 101400, 101360, 101350, 101330, 101330, 101320, 101300, 
    101300, 101270, 101240, 101230, 101240, 101190, 101140, 101120, 101100, 
    101050, 101020, 100970, 100940, 100950, 100940, 100900, 100850, 100810, 
    100790, 100740, 100690, 100670, 100630, 100600, 100540, 100480, 100440, 
    100390, 100320, 100250, 100240, 100260, 100250, 100250, 100270, 100290, 
    100340, 100400, 100430, 100470, 100480, 100510, 100540, 100550, 100580, 
    100590, 100620, 100660, 100700, 100730, 100740, 100730, 100700, 100720, 
    100710, 100690, 100660, 100660, 100630, 100600, 100570, 100540, 100510, 
    100460, 100410, 100340, 100250, 100110, 100030, 99990, 99990, 99960, 
    99990, 99990, 100020, 100030, 100030, 100010, 100000, 99970, 99950, 
    99910, 99890, 99840, 99810, 99760, 99740, 99740, 99740, 99710, 99700, 
    99670, 99650, 99650, 99660, 99650, 99650, 99660, 99660, 99680, 99700, 
    99700, 99680, 99650, 99630, 99610, 99620, 99600, 99590, 99560, 99510, 
    99480, 99420, 99330, 99260, 99210, 99160, 99100, 99030, 98970, 98950, 
    98900, 98900, 98880, 98870, 98870, 98870, 98910, 98910, 98910, 98950, 
    98970, 98980, 99020, 99050, 99060, 99100, 99120, 99150, 99180, 99210, 
    99270, 99320, 99400, 99400, 99460, 99510, 99590, 99660, 99720, 99820, 
    99870, 99880, 99920, 100000, 100060, 100110, 100230, 100330, 100360, 
    100430, 100470, 100470, 100490, 100570, 100600, 100620, 100630, 100690, 
    100710, 100730, 100760, 100770, 100790, 100790, 100810, 100820, 100830, 
    100840, 100840, 100880, 100880, 100910, 100920, 100940, 100950, 100970, 
    100980, 101010, 101030, 101040, 101090, 101100, 101140, 101150, 101150, 
    101150, 101140, 101140, 101130, 101140, 101150, 101140, 101120, 101120, 
    101120, 101100, 101090, 101050, 101010, 100990, 100970, 100900, 100880, 
    100830, 100780, 100750, 100650, 100550, 100420, 100390, 100290, 100210, 
    100080, 99990, 99920, 99810, 99830, 99790, 99790, 99860, 99930, 99990, 
    100070, 100200, 100260, 100340, 100410, 100480, 100570, 100650, 100720, 
    100790, 100840, 100880, 100940, 100990, 101030, 101090, 101160, 101240, 
    101280, 101320, 101420, 101400, 101470, 101520, 101520, 101570, 101670, 
    101750, 101860, 101960, 102050, 102130, 102180, 102210, 102290, 102330, 
    102380, 102420, 102490, 102480, 102530, 102560, 102570, 102610, 102630, 
    102650, 102650, 102650, 102650, 102670, 102660, 102650, 102640, 102670, 
    102680, 102670, 102670, 102670, 102650, 102650, 102640, 102630, 102600, 
    102590, 102550, 102580, 102580, 102580, 102580, 102540, 102510, 102480, 
    102500, 102490, 102460, 102440, 102430, 102440, 102410, 102390, 102360, 
    102330, 102300, 102310, 102300, 102280, 102240, 102220, 102190, 102200, 
    102200, 102180, 102180, 102170, 102160, 102170, 102150, 102100, 102110, 
    102100, 102090, 102080, 102100, 102070, 102090, 102090, 102100, 102100, 
    102110, 102100, 102130, 102130, 102140, 102140, 102180, 102170, 102180, 
    102170, 102160, 102150, 102150, 102150, 102140, 102140, 102130, 102160, 
    102180, 102180, 102190, 102240, 102260, 102230, 102220, 102210, 102210, 
    102210, 102190, 102190, 102150, 102160, 102170, 102180, 102160, 102150, 
    102160, 102150, 102110, 102100, 102110, 102120, 102100, 102110, 102130, 
    102120, 102100, 102080, 102110, 102090, 102080, 102060, 102050, 102040, 
    102050, 102070, 102090, 102090, 102080, 102060, 102050, 102030, 102010, 
    102010, 102020, 102010, 102020, 102020, 102050, 102050, 102040, 102050, 
    102060, 101990, 101970, 101940, 101920, 101940, 101920, 101910, 101930, 
    101980, 101970, 101980, 101990, 101990, 101940, 101940, 101960, 101980, 
    102000, 102020, 102050, 102070, 102070, 102070, 102020, 102030, 102030, 
    102060, 102100, 102120, 102140, 102140, 102150, 102180, 102170, 102180, 
    102190, 102230, 102220, 102260, 102270, 102290, 102320, 102360, 102380, 
    102360, 102370, 102410, 102380, 102420, 102460, 102500, 102540, 102550, 
    102540, 102570, 102580, 102570, 102570, 102540, 102590, 102610, 102620, 
    102630, 102630, 102620, 102610, 102590, 102570, 102570, 102550, 102540, 
    102500, 102470, 102490, 102450, 102450, 102430, 102420, 102400, 102380, 
    102370, 102330, 102310, 102290, 102270, 102240, 102250, 102230, 102190, 
    102180, 102190, 102190, 102130, 102100, 102070, 102060, 102060, 101990, 
    101980, 101950, 101920, 101880, 101850, 101810, 101780, 101770, 101710, 
    101680, 101670, 101650, 101590, 101580, 101540, 101500, 101470, 101480, 
    101410, 101390, 101340, 101280, 101200, 101140, 101090, 101040, 100980, 
    100920, 100900, 100870, 100850, 100830, 100780, 100750, 100740, 100750, 
    100780, 100800, 100830, 100880, 100930, 100980, 101020, 101050, 101130, 
    101170, 101230, 101300, 101370, 101400, 101440, 101490, 101540, 101560, 
    101580, 101600, 101640, 101670, 101640, 101620, 101600, 101520, 101440, 
    101370, 101380, 101280, 101210, 101190, 101140, 101140, 101050, 100990, 
    100890, 100910, 100860, 100850, 100880, 100890, 100920, 100990, 100990, 
    101000, 100990, 101020, 101020, 101030, 101090, 101160, 101260, 101350, 
    101510, 101590, 101730, 101830, 101910, 102010, 102140, 102240, 102310, 
    102380, 102440, 102570, 102650, 102720, 102750, 102820, 102860, 102880, 
    102940, 102980, 102970, 103030, 103080, 103100, 103140, 103170, 103170, 
    103150, 103160, 103170, 103160, 103130, 103120, 103080, 103060, 103050, 
    103020, 102970, 102930, 102900, 102890, 102850, 102850, 102830, 102840, 
    102820, 102820, 102830, 102840, 102850, 102860, 102850, 102840, 102800, 
    102820, 102790, 102770, 102740, 102710, 102650, 102600, 102540, 102470, 
    102390, 102310, 102230, 102150, 102100, 102040, 101990, 101920, 101870, 
    101810, 101780, 101730, 101670, 101640, 101560, 101550, 101520, 101500, 
    101490, 101500, 101520, 101510, 101510, 101530, 101500, 101480, 101430, 
    101420, 101340, 101320, 101260, 101170, 101100, 101050, 100940, 100920, 
    100780, 100760, 100720, 100700, 100700, 100690, 100660, 100670, 100740, 
    100830, 100960, 101080, 101200, 101350, 101510, 101660, 101780, 101900, 
    102050, 102130, 102250, 102370, 102440, 102530, 102600, 102680, 102730, 
    102780, 102860, 102890, 102940, 102960, 102990, 102960, 102930, 102920, 
    102880, 102870, 102800, 102710, 102620, 102580, 102510, 102460, 102380, 
    102280, 102240, 102120, 102070, 101980, 101920, 101820, 101770, 101700, 
    101660, 101630, 101580, 101560, 101540, 101480, 101470, 101470, 101530, 
    101540, 101540, 101590, 101650, 101720, 101720, 101740, 101740, 101830, 
    101880, 101940, 101990, 102020, 102040, 102050, 102060, 102030, 102040, 
    102020, 102010, 101990, 101950, 101980, 101980, 102010, 102040, 102080, 
    102130, 102190, 102210, 102240, 102290, 102330, 102360, 102370, 102370, 
    102420, 102430, 102450, 102450, 102490, 102570, 102450, 102420, 102370, 
    102400, 102310, 102330, 102340, 102340, 102390, 102380, 102390, 102420, 
    102440, 102450, 102470, 102490, 102500, 102520, 102550, 102510, 102530, 
    102510, 102480, 102500, 102510, 102530, 102520, 102520, 102510, 102530, 
    102490, 102500, 102510, 102540, 102520, 102510, 102510, 102480, 102440, 
    102430, 102430, 102400, 102370, 102330, 102300, 102330, 102300, 102300, 
    102310, 102320, 102300, 102310, 102320, 102290, 102260, 102340, 102360, 
    102360, 102420, 102420, 102460, 102470, 102500, 102480, 102500, 102570, 
    102580, 102590, 102630, 102630, 102640, 102660, 102670, 102660, 102690, 
    102690, 102710, 102720, 102710, 102660, 102660, 102630, 102600, 102580, 
    102540, 102500, 102550, 102570, 102480, 102410, 102400, 102370, 102290, 
    102310, 102260, 102220, 102160, 102140, 102140, 102090, 102030, 102010, 
    102020, 102000, 101990, 102000, 101990, 101920, 101860, 101790, 101760, 
    101690, 101650, 101590, 101510, 101430, 101370, 101310, 101250, 101180, 
    101130, 101040, 100940, 100900, 100860, 100790, 100740, 100700, 100680, 
    100630, 100590, 100570, 100510, 100470, 100430, 100390, 100360, 100310, 
    100240, 100200, 100170, 100170, 100140, 100090, 100050, 100020, 100020, 
    100020, 100010, 99990, 99980, 99990, 99980, 99990, 100020, 100040, 
    100050, 100050, 100070, 100080, 100080, 100080, 100070, 100100, 100110, 
    100130, 100160, 100190, 100200, 100230, 100250, 100270, 100260, 100290, 
    100280, 100320, 100360, 100410, 100470, 100520, 100550, 100560, 100580, 
    100610, 100640, 100680, 100700, 100710, 100760, 100790, 100830, 100860, 
    100900, 100910, 100950, 100960, 100970, 101020, 101040, 101060, 101060, 
    101090, 101110, 101140, 101170, 101210, 101240, 101230, 101200, 101220, 
    101250, 101250, 101270, 101300, 101300, 101330, 101350, 101340, 101340, 
    101360, 101400, 101400, 101390, 101400, 101410, 101420, 101420, 101420, 
    101420, 101420, 101440, 101450, 101460, 101470, 101460, 101450, 101450, 
    101470, 101490, 101520, 101520, 101520, 101520, 101530, 101530, 101530, 
    101540, 101540, 101550, 101580, 101600, 101620, 101650, 101680, 101690, 
    101700, 101720, 101720, 101730, 101730, 101720, 101730, 101760, 101760, 
    101750, 101740, 101730, 101740, 101730, 101740, 101740, 101730, 101720, 
    101710, 101710, 101710, 101690, 101670, 101630, 101600, 101580, 101530, 
    101540, 101530, 101530, 101520, 101510, 101540, 101550, 101550, 101570, 
    101590, 101600, 101600, 101590, 101610, 101600, 101590, 101590, 101600, 
    101590, 101570, 101550, 101550, 101560, 101570, 101570, 101560, 101590, 
    101610, 101630, 101660, 101680, 101680, 101700, 101720, 101710, 101720, 
    101740, 101740, 101730, 101720, 101750, 101750, 101740, 101740, 101740, 
    101730, 101690, 101720, 101730, 101710, 101730, 101740, 101760, 101740, 
    101750, 101760, 101750, 101750, 101770, 101790, 101790, 101800, 101830, 
    101850, 101880, 101920, 101920, 101930, 101950, 101950, 101960, 101990, 
    102030, 102020, 102020, 102040, 102040, 102040, 102050, 102060, 102060, 
    102050, 102080, 102090, 102110, 102120, 102150, 102150, 102200, 102170, 
    102160, 102140, 102140, 102130, 102140, 102120, 102110, 102110, 102090, 
    102070, 102090, 102080, 102080, 102070, 102070, 102070, 102050, 102040, 
    102040, 102040, 102050, 102030, 102040, 102050, 102030, 102010, 102030, 
    102000, 101970, 101860, 101880, 101950, 102000, 102030, 102060, 102070, 
    102080, 102080, 102020, 102040, 102020, 102000, 101960, 101960, 101980, 
    102000, 102030, 102050, 102060, 102060, 102030, 102010, 102010, 102000, 
    101980, 101990, 101990, 101960, 101910, 101910, 101850, 101800, 101770, 
    101730, 101700, 101640, 101620, 101590, 101580, 101550, 101560, 101550, 
    101530, 101540, 101550, 101550, 101540, 101540, 101520, 101550, 101570, 
    101590, 101600, 101610, 101630, 101650, 101660, 101660, 101660, 101650, 
    101630, 101620, 101660, 101700, 101740, 101760, 101780, 101810, 101810, 
    101830, 101850, 101870, 101890, 101920, 101940, 101980, 101980, 102010, 
    102020, 102030, 102030, 102050, 102060, 102070, 102100, 102110, 102130, 
    102150, 102160, 102170, 102150, 102180, 102180, 102180, 102160, 102140, 
    102140, 102140, 102150, 102160, 102170, 102160, 102140, 102110, 102110, 
    102120, 102100, 102110, 102070, 102070, 102050, 102040, 102020, 102000, 
    101970, 101950, 101950, 101930, 101920, 101910, 101890, 101860, 101840, 
    101830, 101840, 101840, 101790, 101760, 101720, 101730, 101750, 101740, 
    101710, 101730, 101710, 101750, 101740, 101780, 101790, 101800, 101820, 
    101850, 101830, 101860, 101880, 101890, 101940, 101940, 101940, 101960, 
    101970, 101980, 101990, 101990, 101990, 102010, 101990, 102010, 102020, 
    102050, 102060, 102050, 102050, 102070, 102080, 102060, 102100, 102090, 
    102110, 102090, 102100, 102090, 102070, 102060, 102040, 102000, 101980, 
    101940, 101930, 101880, 101880, 101790, 101760, 101740, 101680, 101570, 
    101450, 101380, 101260, 101200, 101140, 101090, 101020, 100950, 100930, 
    100850, 100780, 100710, 100660, 100610, 100550, 100530, 100540, 100530, 
    100530, 100550, 100550, 100570, 100570, 100530, 100510, 100490, 100440, 
    100460, 100480, 100490, 100540, 100530, 100560, 100560, 100560, 100590, 
    100650, 100660, 100680, 100740, 100780, 100800, 100800, 100840, 100870, 
    100890, 100930, 100950, 100970, 100980, 100970, 100900, 100870, 100860, 
    100850, 100820, 100810, 100830, 100790, 100740, 100740, 100720, 100700, 
    100700, 100710, 100710, 100670, 100680, 100660, 100670, 100670, 100700, 
    100700, 100710, 100690, 100680, 100680, 100660, 100650, 100680, 100680, 
    100670, 100650, 100640, 100630, 100620, 100610, 100580, 100550, 100510, 
    100480, 100430, 100410, 100350, 100350, 100320, 100290, 100250, 100170, 
    100110, 100070, 100010, 99960, 99900, 99830, 99780, 99710, 99660, 99600, 
    99550, 99470, 99420, 99350, 99280, 99240, 99200, 99090, 99110, 99080, 
    99010, 98990, 98950, 98910, 98890, 98860, 98710, 98650, 98680, 98680, 
    98640, 98590, 98520, 98490, 98460, 98410, 98360, 98340, 98290, 98230, 
    98290, 98230, 98280, 98270, 98170, 98150, 98110, 98120, 98090, 98150, 
    98230, 98310, 98360, 98440, 98500, 98530, 98570, 98600, 98620, 98690, 
    98690, 98650, 98700, 98720, 98770, 98760, 98770, 98800, 98800, 98770, 
    98780, 98830, 98850, 98860, 98930, 98960, 98970, 99000, 99010, 99030, 
    99070, 99080, 99070, 99070, 99080, 99110, 99130, 99150, 99180, 99210, 
    99200, 99190, 99150, 99070, 99030, 98960, 98920, 98920, 98890, 98820, 
    98880, 98880, 98940, 98970, 99000, 98970, 98990, 99000, 99020, 99020, 
    99040, 99020, 99010, 99050, 99040, 99050, 99070, 99090, 99100, 99120, 
    99130, 99140, 99160, 99170, 99180, 99210, 99220, 99240, 99240, 99260, 
    99280, 99300, 99310, 99340, 99360, 99390, 99410, 99430, 99470, 99490, 
    99510, 99510, 99530, 99510, 99500, 99500, 99520, 99510, 99500, 99510, 
    99490, 99490, 99490, 99450, 99430, 99420, 99400, 99380, 99350, 99320, 
    99300, 99270, 99250, 99230, 99210, 99180, 99140, 99080, 99020, 98950, 
    98900, 98820, 98810, 98760, 98740, 98690, 98680, 98660, 98660, 98660, 
    98670, 98610, 98620, 98640, 98600, 98620, 98600, 98580, 98510, 98470, 
    98430, 98420, 98440, 98490, 98500, 98530, 98550, 98560, 98610, 98670, 
    98690, 98740, 98820, 98970, 98960, 99060, 99170, 99260, 99350, 99390, 
    99450, 99470, 99490, 99540, 99600, 99600, 99610, 99620, 99630, 99620, 
    99630, 99640, 99730, 99860, 99880, 99910, 99960, 99990, 100050, 100100, 
    100150, 100180, 100220, 100300, 100330, 100410, 100440, 100490, 100540, 
    100560, 100650, 100700, 100760, 100790, 100830, 100870, 100920, 100960, 
    101010, 101040, 101080, 101120, 101160, 101200, 101210, 101240, 101290, 
    101330, 101380, 101410, 101440, 101480, 101500, 101530, 101560, 101580, 
    101590, 101630, 101650, 101670, 101730, 101760, 101780, 101800, 101820, 
    101840, 101880, 101910, 101920, 101950, 101980, 102030, 102080, 102080, 
    102130, 102190, 102220, 102250, 102300, 102320, 102360, 102370, 102410, 
    102440, 102480, 102490, 102510, 102510, 102520, 102510, 102520, 102520, 
    102510, 102530, 102490, 102480, 102480, 102450, 102430, 102400, 102350, 
    102310, 102270, 102240, 102220, 102170, 102120, 102090, 102060, 102010, 
    101920, 101870, 101790, 101730, 101680, 101690, 101660, 101630, 101620, 
    101600, 101580, 101570, 101560, 101540, 101510, 101480, 101420, 101380, 
    101330, 101240, 101170, 101100, 101120, 101140, 101160, 101230, 101290, 
    101190, 101180, 101290, 101330, 101360, 101370, 101340, 101260, 101280, 
    101240, 101270, 101410, 101470, 101430, 101410, 101360, 101320, 101250, 
    101190, 101210, 101250, 101180, 101140, 101120, 101060, 100960, 100900, 
    100840, 100880, 100850, 100860, 100870, 100870, 100870, 100850, 100800, 
    100730, 100680, 100660, 100730, 100660, 100550, 100510, 100390, 100510, 
    100580, 100570, 100550, 100550, 100510, 100440, 100310, 100300, 100330, 
    100360, 100410, 100430, 100430, 100480, 100470, 100460, 100460, 100430, 
    100420, 100400, 100330, 100270, 100250, 100260, 100300, 100320, 100360, 
    100400, 100450, 100480, 100520, 100540, 100560, 100630, 100620, 100650, 
    100670, 100670, 100700, 100710, 100700, 100690, 100650, 100650, 100690, 
    100700, 100720, 100730, 100740, 100730, 100700, 100730, 100740, 100770, 
    100780, 100820, 100860, 100890, 100920, 100920, 100960, 101000, 101020, 
    101040, 101090, 101120, 101160, 101210, 101310, 101310, 101300, 101270, 
    101310, 101310, 101300, 101320, 101380, 101310, 101330, 101400, 101460, 
    101480, 101520, 101590, 101640, 101650, 101700, 101740, 101750, 101730, 
    101700, 101660, 101800, 101820, 101810, 101820, 101840, 101850, 101840, 
    101840, 101830, 101850, 101870, 101890, 101900, 101880, 101940, 101950, 
    101950, 101940, 101980, 101950, 102020, 101970, 101960, 102000, 102020, 
    102020, 102030, 102020, 102000, 101980, 101960, 101950, 101950, 101930, 
    101900, 101880, 101830, 101810, 101870, 101880, 101870, 101870, 101750, 
    101880, 101940, 102020, 102030, 102020, 102050, 102080, 102100, 102140, 
    102160, 102160, 102180, 102180, 102220, 102220, 102210, 102230, 102250, 
    102260, 102330, 102370, 102380, 102380, 102340, 102420, 102440, 102430, 
    102440, 102440, 102360, 102430, 102450, 102490, 102490, 102520, 102520, 
    102540, 102550, 102550, 102560, 102580, 102600, 102620, 102660, 102720, 
    102770, 102780, 102800, 102820, 102850, 102880, 102890, 102890, 102900, 
    102940, 102980, 102980, 103010, 103010, 103020, 103110, 103150, 103130, 
    103150, 103190, 103210, 103250, 103360, 103400, 103430, 103540, 103520, 
    103510, 103580, 103590, 103630, 103660, 103690, 103720, 103770, 103800, 
    103860, 103860, 103890, 103890, 103900, 103900, 103950, 103950, 103960, 
    103950, 103950, 103970, 104010, 104100, 104090, 104050, 104080, 104100, 
    104120, 104090, 104130, 104100, 104140, 104140, 104090, 104090, 104160, 
    104170, 104220, 104250, 104230, 104220, 104200, 104210, 104220, 104250, 
    104270, 104270, 104270, 104230, 104260, 104270, 104280, 104280, 104270, 
    104280, 104310, 104280, 104290, 104310, 104320, 104310, 104300, 104330, 
    104330, 104290, 104270, 104270, 104250, 104250, 104220, 104180, 104150, 
    104100, 104070, 104050, 104010, 103990, 103960, 103910, 103880, 103850, 
    103800, 103790, 103730, 103670, 103600, 103580, 103560, 103520, 103480, 
    103460, 103450, 103430, 103390, 103350, 103310, 103280, 103240, 103200, 
    103180, 103170, 103130, 103050, 102990, 102950, 102920, 102850, 102800, 
    102750, 102720, 102650, 102580, 102530, 102470, 102420, 102370, 102350, 
    102280, 102240, 102180, 102090, 102000, 101940, 101880, 101820, 101760, 
    101690, 101630, 101550, 101480, 101410, 101330, 101270, 101180, 101080, 
    101010, 100940, 100860, 100790, 100730, 100660, 100610, 100550, 100460, 
    100390, 100360, 100360, 100340, 100340, 100340, 100350, 100350, 100350, 
    100340, 100360, 100340, 100320, 100280, 100270, 100270, 100290, 100330, 
    100330, 100330, 100350, 100350, 100290, 100300, 100340, 100360, 100380, 
    100460, 100530, 100560, 100560, 100570, 100570, 100630, 100630, 100610, 
    100650, 100670, 100630, 100670, 100680, 100700, 100790, 101020, 101070, 
    101100, 101140, 101160, 101180, 101230, 101260, 101250, 101280, 101310, 
    101310, 101300, 101270, 101340, 101330, 101320, 101290, 101290, 101260, 
    101230, 101250, 101230, 101220, 101240, 101290, 101280, 101270, 101270, 
    101280, 101290, 101320, 101340, 101350, 101400, 101400, 101420, 101420, 
    101430, 101420, 101420, 101340, 101350, 101360, 101350, 101330, 101310, 
    101300, 101310, 101310, 101310, 101340, 101300, 101270, 101250, 101260, 
    101230, 101220, 101210, 101200, 101190, 101170, 101150, 101080, 101020, 
    100930, 100820, 100760, 100630, 100450, 100270, 100110, 99900, 99700, 
    99490, 99350, 99330, 99370, 99350, 99340, 99330, 99300, 99330, 99350, 
    99390, 99430, 99480, 99520, 99540, 99550, 99570, 99590, 99570, 99560, 
    99530, 99490, 99450, 99410, 99400, 99380, 99330, 99290, 99260, 99250, 
    99250, 99260, 99270, 99290, 99300, 99310, 99300, 99330, 99340, 99400, 
    99420, 99440, 99450, 99410, 99430, 99440, 99470, 99480, 99400, 99430, 
    99420, 99460, 99540, 99600, 99680, 99730, 99790, 99680, 99870, 99920, 
    99960, 99970, 100010, 99990, 99980, 99960, 100040, 100040, 100060, 
    100080, 100150, 100220, 100220, 100320, 100350, 100410, 100450, 100460, 
    100490, 100520, 100550, 100560, 100550, 100570, 100560, 100570, 100540, 
    100540, 100550, 100530, 100530, 100570, 100580, 100650, 100690, 100640, 
    100700, 100700, 100740, 100760, 100720, 100810, 100780, 100790, 100800, 
    100820, 100800, 100690, 100750, 100710, 100840, 100850, 100910, 101020, 
    101040, 101000, 101100, 101150, 101180, 101220, 101240, 101260, 101310, 
    101370, 101390, 101380, 101440, 101460, 101470, 101550, 101550, 101550, 
    101530, 101590, 101550, 101610, 101630, 101610, 101630, 101600, 101600, 
    101640, 101630, 101570, 101540, 101580, 101540, 101690, 101770, 101810, 
    101820, 101810, 101850, 101900, 101920, 101940, 101960, 101980, 102000, 
    102020, 102030, 102050, 102020, 102020, 102010, 102100, 102160, 102170, 
    102230, 102250, 102260, 102250, 102280, 102340, 102340, 102390, 102360, 
    102380, 102390, 102430, 102440, 102460, 102480, 102470, 102470, 102460, 
    102440, 102420, 102420, 102400, 102400, 102430, 102400, 102370, 102330, 
    102270, 102250, 102240, 102230, 102220, 102180, 102120, 102130, 102100, 
    102080, 102050, 102000, 101980, 101980, 101950, 101920, 101900, 101870, 
    101860, 101840, 101840, 101830, 101800, 101740, 101730, 101730, 101720, 
    101730, 101760, 101770, 101770, 101780, 101770, 101760, 101760, 101710, 
    101740, 101680, 101670, 101700, 101710, 101690, 101680, 101710, 101720, 
    101690, 101670, 101690, 101670, 101660, 101640, 101630, 101580, 101550, 
    101490, 101460, 101390, 101390, 101340, 101310, 101230, 101180, 101150, 
    101120, 101080, 101020, 100940, 100910, 100890, 100780, 100670, 100610, 
    100520, 100440, 100350, 100170, 100300, 99990, 99930, 99880, 99670, 
    99660, 99630, 99570, 99510, 99560, 99450, 99420, 99410, 99400, 99450, 
    99470, 99540, 99590, 99630, 99660, 99690, 99700, 99740, 99790, 99850, 
    99870, 99890, 99890, 99760, 99700, 99710, 99710, 99690, 99720, 99750, 
    99710, 99880, 100050, 100060, 100050, 100090, 100080, 100080, 100070, 
    100050, 100030, 100000, 99970, 99940, 99950, 99990, 99990, 99970, 99930, 
    99950, 99970, 100010, 100200, 100230, 100260, 100250, 100270, 100320, 
    100300, 100150, 100140, 100260, 100280, 100310, 100340, 100340, 100120, 
    100060, 100040, 100090, 100150, 100230, 100310, 100280, 100320, 100360, 
    100390, 100390, 100410, 100410, 100420, 100420, 100430, 100460, 100480, 
    100450, 100450, 100440, 100460, 100460, 100440, 100380, 100390, 100350, 
    100350, 100350, 100360, 100340, 100320, 100340, 100330, 100270, 100300, 
    100270, 100260, 100270, 100230, 100210, 100150, 100140, 100090, 100050, 
    99980, 100000, 100020, 100050, 100080, 100110, 100100, 100120, 100150, 
    100150, 100180, 100190, 100190, 100180, 100190, 100190, 100220, 100250, 
    100250, 100270, 100300, 100320, 100350, 100380, 100450, 100480, 100490, 
    100520, 100530, 100560, 100580, 100580, 100600, 100640, 100610, 100600, 
    100580, 100530, 100490, 100450, 100420, 100400, 100350, 100300, 100290, 
    100270, 100170, 100020, 99880, 99730, 99510, 99350, 99160, 98960, 98760, 
    98550, 98350, 98100, 97820, 97570, 97280, 97000, 96730, 96610, 96560, 
    96550, 96510, 96500, 96460, 96380, 96300, 96230, 96220, 96230, 96250, 
    96270, 96270, 96260, 96250, 96250, 96230, 96310, 96400, 96480, 96580, 
    96680, 96750, 96820, 96890, 96950, 97060, 97200, 97320, 97410, 97480, 
    97520, 97570, 97590, 97670, 97700, 97830, 97970, 98040, 98160, 98260, 
    98330, 98420, 98520, 98620, 98710, 98790, 98800, 98890, 98930, 98920, 
    98930, 98790, 98810, 98850, 98880, 98920, 98980, 98950, 98950, 99000, 
    99080, 99110, 99140, 99130, 99210, 99210, 99250, 99230, 99280, 99360, 
    99430, 99520, 99590, 99640, 99690, 99760, 99820, 99870, 99940, 100000, 
    100020, 100040, 100070, 100090, 100110, 100150, 100180, 100230, 100270, 
    100300, 100320, 100320, 100350, 100350, 100340, 100320, 100380, 100390, 
    100430, 100430, 100410, 100350, 100410, 100400, 100410, 100370, 100370, 
    100410, 100420, 100440, 100510, 100660, 100730, 100760, 100780, 100840, 
    100940, 101040, 101090, 101160, 101240, 101290, 101290, 101330, 101360, 
    101450, 101510, 101520, 101480, 101500, 101560, 101550, 101590, 101600, 
    101670, 101620, 101600, 101670, 101650, 101620, 101600, 101540, 101460, 
    101320, 101150, 100920, 100790, 100770, 100590, 100470, 100400, 100300, 
    100240, 100150, 100130, 100070, 100140, 100180, 100160, 100200, 100260, 
    100320, 100360, 100370, 100400, 100380, 100340, 100330, 100310, 100340, 
    100330, 100320, 100220, 100100, 100080, 100030, 99970, 99860, 99700, 
    99510, 99360, 99170, 98950, 98690, 98470, 98240, 98060, 98010, 97940, 
    97900, 97890, 97880, 97920, 97960, 98030, 98080, 98110, 98130, 98180, 
    98250, 98300, 98400, 98430, 98490, 98540, 98610, 98670, 98700, 98710, 
    98770, 98820, 98870, 98910, 98930, 98890, 98870, 98970, 98940, 98900, 
    98880, 98870, 98850, 98950, 99030, 99060, 99100, 99140, 99170, 99240, 
    99370, 99520, 99620, 99630, 99770, 99920, 100050, 100110, 100120, 100200, 
    100380, 100500, 100560, 100630, 100590, 100660, 100690, 100740, 100770, 
    100820, 100840, 100810, 100840, 100890, 100860, 100890, 100860, 100850, 
    100850, 100860, 100890, 100890, 100880, 100870, 100870, 100880, 100890, 
    100880, 100900, 100940, 100930, 100900, 100920, 100960, 100930, 100920, 
    100950, 100940, 100960, 100930, 100960, 100970, 100940, 100950, 100960, 
    100930, 100910, 100900, 100880, 100860, 100860, 100850, 100840, 100810, 
    100750, 100740, 100740, 100710, 100700, 100680, 100640, 100610, 100600, 
    100600, 100590, 100590, 100570, 100540, 100510, 100490, 100460, 100430, 
    100400, 100380, 100350, 100350, 100360, 100340, 100350, 100340, 100310, 
    100320, 100340, 100340, 100330, 100370, 100400, 100400, 100400, 100380, 
    100360, 100320, 100320, 100300, 100320, 100300, 100300, 100330, 100330, 
    100360, 100390, 100400, 100410, 100430, 100420, 100440, 100460, 100510, 
    100550, 100540, 100560, 100580, 100660, 100620, 100650, 100700, 100720, 
    100730, 100720, 100760, 100790, 100790, 100820, 100850, 100860, 100920, 
    100920, 100920, 100900, 100980, 100940, 100990, 101020, 101020, 101040, 
    101050, 101090, 101080, 101110, 101130, 101130, 101120, 101120, 101110, 
    101140, 101210, 101200, 101220, 101210, 101240, 101270, 101220, 101220, 
    101200, 101230, 101200, 101200, 101220, 101230, 101220, 101210, 101150, 
    101130, 101100, 101070, 100970, 100850, 100660, 100610, 100570, 100470, 
    100500, 100470, 100510, 100530, 100560, 100570, 100610, 100620, 100600, 
    100610, 100610, 100600, 100590, 100590, 100610, 100610, 100610, 100590, 
    100560, 100480, 100460, 100440, 100420, 100420, 100340, 100320, 100310, 
    100280, 100290, 100240, 100220, 100190, 100130, 100080, 100050, 100020, 
    100080, 100170, 100180, 100220, 100250, 100320, 100350, 100420, 100480, 
    100540, 100610, 100670, 100720, 100780, 100830, 100880, 100920, 100970, 
    100990, 101040, 101040, 101090, 101150, 101170, 101170, 101180, 101210, 
    101230, 101230, 101260, 101260, 101270, 101280, 101310, 101330, 101370, 
    101420, 101400, 101420, 101410, 101460, 101490, 101480, 101500, 101510, 
    101530, 101530, 101540, 101550, 101550, 101540, 101550, 101580, 101590, 
    101570, 101570, 101570, 101550, 101550, 101550, 101570, 101550, 101550, 
    101510, 101510, 101490, 101440, 101430, 101420, 101400, 101380, 101370, 
    101380, 101370, 101360, 101340, 101290, 101280, 101240, 101220, 101200, 
    101180, 101160, 101170, 101130, 101130, 101160, 101130, 101100, 101090, 
    101060, 101030, 101040, 101020, 100980, 100940, 100890, 100910, 100880, 
    100860, 100840, 100810, 100810, 100760, 100740, 100710, 100690, 100700, 
    100680, 100650, 100560, 100490, 100430, 100440, 100440, 100510, 100490, 
    100540, 100590, 100610, 100640, 100660, 100730, 100690, 100680, 100610, 
    100530, 100460, 100320, 100190, 100070, 99970, 99830, 99710, 99560, 
    99460, 99240, 99090, 98930, 98800, 98710, 98660, 98620, 98490, 98430, 
    98400, 98340, 98300, 98330, 98390, 98390, 98450, 98500, 98640, 98750, 
    98820, 98940, 99060, 99140, 99210, 99260, 99330, 99360, 99350, 99380, 
    99420, 99460, 99500, 99500, 99550, 99580, 99610, 99610, 99610, 99640, 
    99620, 99620, 99580, 99590, 99590, 99600, 99600, 99650, 99690, 99720, 
    99690, 99710, 99720, 99770, 99790, 99810, 99850, 99880, 99920, 99940, 
    99960, 99960, 99970, 99970, 99990, 100030, 100040, 100080, 100120, 
    100150, 100200, 100260, 100300, 100250, 100280, 100330, 100340, 100380, 
    100390, 100390, 100450, 100560, 100640, 100720, 100770, 100870, 100890, 
    100950, 101000, 101080, 101160, 101220, 101280, 101340, 101400, 101460, 
    101480, 101480, 101530, 101570, 101580, 101660, 101690, 101740, 101790, 
    101820, 101790, 101840, 101830, 101820, 101820, 101840, 101880, 101920, 
    101950, 101990, 102020, 102030, 102000, 101970, 101970, 101900, 101880, 
    101830, 101760, 101750, 101730, 101760, 101750, 101820, 101880, 101950, 
    102000, 102020, 102050, 102060, 102090, 102110, 102150, 102190, 102240, 
    102280, 102320, 102360, 102370, 102370, 102390, 102420, 102390, 102350, 
    102330, 102310, 102310, 102330, 102310, 102280, 102190, 102120, 102040, 
    101980, 101900, 101840, 101750, 101670, 101560, 101520, 101580, 101510, 
    101470, 101430, 101400, 101360, 101360, 101310, 101230, 101060, 100960, 
    100940, 100930, 100900, 100980, 101100, 101300, 101460, 101550, 101640, 
    101720, 101780, 101870, 101910, 101940, 101960, 101950, 101930, 101960, 
    101970, 102000, 102040, 102100, 102090, 102090, 102100, 102090, 102090, 
    102090, 102090, 102100, 102090, 102060, 102080, 102070, 102070, 102090, 
    102110, 102140, 102150, 102150, 102150, 102160, 102150, 102160, 102150, 
    102160, 102160, 102180, 102180, 102200, 102200, 102220, 102200, 102230, 
    102250, 102250, 102270, 102270, 102280, 102280, 102280, 102280, 102300, 
    102270, 102290, 102270, 102270, 102250, 102250, 102220, 102200, 102180, 
    102170, 102140, 102100, 102050, 102020, 101960, 101920, 101920, 101890, 
    101840, 101800, 101760, 101740, 101700, 101640, 101600, 101610, 101590, 
    101570, 101540, 101480, 101470, 101470, 101460, 101440, 101410, 101380, 
    101350, 101320, 101350, 101310, 101280, 101270, 101230, 101250, 101240, 
    101220, 101230, 101190, 101180, 101170, 101140, 101140, 101130, 101130, 
    101130, 101120, 101150, 101100, 101090, 101010, 100950, 100960, 100960, 
    100850, 100840, 100780, 100730, 100690, 100650, 100620, 100570, 100550, 
    100500, 100460, 100490, 100510, 100510, 100530, 100460, 100510, 100540, 
    100630, 100660, 100720, 100760, 100790, 100810, 100790, 100820, 100840, 
    100840, 100850, 100870, 100880, 100910, 100950, 100950, 100960, 101060, 
    101110, 101100, 101110, 101130, 101110, 101120, 101120, 101130, 101110, 
    101090, 101060, 101050, 101020, 100990, 100960, 100920, 100950, 100980, 
    101000, 100990, 101020, 101060, 101080, 101120, 101160, 101180, 101180, 
    101200, 101210, 101240, 101290, 101330, 101360, 101380, 101420, 101420, 
    101450, 101460, 101490, 101490, 101530, 101600, 101630, 101660, 101700, 
    101730, 101730, 101760, 101790, 101800, 101800, 101810, 101840, 101860, 
    101900, 101920, 101920, 101940, 101940, 101950, 101960, 101980, 101970, 
    101960, 101970, 102000, 102040, 102060, 102070, 102080, 102090, 102080, 
    102090, 102110, 102090, 102080, 102090, 102110, 102140, 102130, 102170, 
    102140, 102130, 102180, 102180, 102190, 102190, 102190, 102240, 102280, 
    102320, 102350, 102370, 102410, 102440, 102450, 102490, 102500, 102520, 
    102570, 102600, 102640, 102680, 102720, 102740, 102750, 102770, 102810, 
    102830, 102820, 102820, 102840, 102870, 102890, 102910, 102890, 102880, 
    102870, 102860, 102840, 102800, 102750, 102730, 102680, 102640, 102620, 
    102600, 102560, 102510, 102470, 102390, 102340, 102290, 102220, 102150, 
    102110, 102090, 102080, 102040, 101990, 101940, 101900, 101810, 101720, 
    101690, 101670, 101630, 101580, 101580, 101550, 101540, 101560, 101540, 
    101530, 101550, 101540, 101540, 101530, 101550, 101550, 101540, 101560, 
    101580, 101580, 101580, 101590, 101530, 101550, 101540, 101510, 101470, 
    101440, 101410, 101400, 101320, 101290, 101220, 101170, 101130, 101050, 
    100980, 100880, 100780, 100650, 100530, 100480, 100420, 100350, 100210, 
    100100, 100040, 99920, 99800, 99670, 99580, 99510, 99530, 99470, 99310, 
    99120, 98970, 98770, 98430, 98190, 97930, 97490, 97270, 97150, 97140, 
    97150, 97210, 97260, 97310, 97420, 97520, 97560, 97720, 97850, 98010, 
    98170, 98350, 98530, 98650, 98820, 98940, 99060, 99200, 99320, 99420, 
    99530, 99650, 99860, 100010, 100230, 100380, 100540, 100690, 100750, 
    100840, 100870, 100910, 100960, 100960, 100880, 100790, 100810, 100840, 
    100930, 101020, 101030, 101010, 101010, 101020, 100980, 100930, 100880, 
    100710, 100510, 100340, 100180, 100060, 99730, 99500, 99400, 99250, 
    99130, 99000, 98890, 98820, 98810, 98810, 98780, 98760, 98730, 98750, 
    98750, 98710, 98720, 98700, 98690, 98690, 98710, 98740, 98780, 98830, 
    98840, 98870, 98910, 98940, 98940, 98940, 99000, 99080, 99100, 99140, 
    99210, 99270, 99310, 99380, 99440, 99500, 99560, 99590, 99630, 99670, 
    99730, 99780, 99810, 99850, 99840, 99890, 99920, 99940, 99950, 100010, 
    100060, 100090, 100140, 100200, 100240, 100250, 100240, 100260, 100230, 
    100240, 100230, 100190, 100200, 100190, 100220, 100210, 100150, 100080, 
    100020, 99950, 99870, 99760, 99670, 99560, 99480, 99410, 99310, 99230, 
    99090, 99030, 98900, 98930, 99060, 99230, 99340, 99480, 99530, 99630, 
    99700, 99760, 99780, 99830, 99850, 99870, 99880, 99890, 99920, 99980, 
    100050, 100120, 100190, 100290, 100360, 100450, 100520, 100580, 100610, 
    100680, 100720, 100740, 100790, 100830, 100860, 100920, 100970, 101010, 
    101010, 101030, 101050, 101080, 101110, 101130, 101160, 101180, 101220, 
    101250, 101280, 101300, 101320, 101330, 101350, 101370, 101390, 101370, 
    101380, 101390, 101420, 101440, 101430, 101430, 101400, 101400, 101370, 
    101370, 101380, 101400, 101410, 101430, 101450, 101480, 101490, 101510, 
    101520, 101530, 101550, 101550, 101560, 101560, 101580, 101610, 101630, 
    101660, 101680, 101680, 101690, 101680, 101690, 101690, 101690, 101700, 
    101710, 101700, 101690, 101690, 101700, 101710, 101710, 101700, 101700, 
    101700, 101670, 101700, 101720, 101730, 101750, 101780, 101810, 101850, 
    101860, 101870, 101900, 101900, 101950, 101970, 101970, 101990, 102040, 
    102080, 102110, 102110, 102130, 102170, 102170, 102170, 102170, 102160, 
    102170, 102180, 102210, 102240, 102240, 102260, 102280, 102280, 102300, 
    102320, 102310, 102340, 102360, 102400, 102460, 102520, 102550, 102570, 
    102600, 102650, 102740, 102790, 102840, 102850, 102880, 102900, 102960, 
    103010, 103050, 103100, 103120, 103140, 103180, 103230, 103280, 103280, 
    103290, 103310, 103330, 103370, 103370, 103380, 103380, 103390, 103400, 
    103390, 103380, 103350, 103320, 103320, 103310, 103320, 103320, 103310, 
    103320, 103300, 103310, 103320, 103300, 103260, 103260, 103230, 103230, 
    103220, 103220, 103210, 103180, 103160, 103150, 103130, 103110, 103100, 
    103110, 103080, 103080, 103120, 103140, 103150, 103170, 103150, 103170, 
    103170, 103160, 103140, 103170, 103170, 103190, 103190, 103220, 103220, 
    103230, 103250, 103290, 103310, 103290, 103290, 103300, 103370, 103410, 
    103470, 103510, 103540, 103570, 103590, 103590, 103600, 103620, 103640, 
    103630, 103650, 103620, 103620, 103680, 103680, 103630, 103620, 103610, 
    103600, 103600, 103570, 103560, 103530, 103550, 103550, 103570, 103570, 
    103560, 103580, 103600, 103590, 103630, 103630, 103590, 103580, 103600, 
    103640, 103660, 103690, 103700, 103790, 103760, 103780, 103790, 103790, 
    103790, 103810, 103840, 103860, 103920, 103950, 103970, 104010, 104040, 
    104060, 104070, 104110, 104130, 104160, 104170, 104200, 104220, 104250, 
    104250, 104250, 104250, 104270, 104250, 104230, 104180, 104190, 104150, 
    104150, 104150, 104130, 104080, 104060, 104030, 104020, 104020, 103980, 
    103920, 103880, 103880, 103880, 103870, 103900, 103850, 103830, 103850, 
    103880, 103870, 103920, 103970, 103980, 104030, 104090, 104130, 104220, 
    104280, 104350, 104380, 104410, 104430, 104460, 104460, 104460, 104460, 
    104440, 104410, 104410, 104370, 104340, 104300, 104280, 104230, 104210, 
    104170, 104110, 104100, 104050, 104050, 104010, 103860, 103850, 103810, 
    103840, 103810, 103780, 103670, 103710, 103650, 103590, 103510, 103520, 
    103460, 103430, 103380, 103370, 103280, 103270, 103240, 103230, 103270, 
    103270, 103290, 103310, 103270, 103180, 103080, 103140, 103020, 102950, 
    102790, 102700, 102550, 102430, 102300, 102220, 102170, 102080, 102020, 
    101920, 101830, 101760, 101680, 101640, 101600, 101570, 101570, 101490, 
    101400, 101380, 101310, 101300, 101300, 101310, 101290, 101290, 101350, 
    101360, 101400, 101470, 101490, 101550, 101590, 101650, 101710, 101710, 
    101740, 101770, 101830, 101920, 102020, 102110, 102210, 102270, 102370, 
    102440, 102540, 102610, 102660, 102690, 102710, 102760, 102800, 102810, 
    102830, 102830, 102850, 102870, 102890, 102850, 102820, 102780, 102780, 
    102740, 102720, 102730, 102690, 102660, 102590, 102500, 102460, 102430, 
    102420, 102430, 102350, 102300, 102240, 102240, 102220, 102180, 102210, 
    102200, 102170, 102120, 102120, 102100, 102020, 102090, 102060, 102110, 
    102130, 102200, 102210, 102250, 102220, 102240, 102270, 102280, 102330, 
    102370, 102420, 102460, 102520, 102550, 102590, 102620, 102620, 102640, 
    102670, 102690, 102750, 102810, 102830, 102880, 102910, 102910, 102940, 
    102980, 103040, 103070, 103100, 103150, 103190, 103200, 103220, 103240, 
    103230, 103240, 103260, 103260, 103270, 103280, 103290, 103320, 103320, 
    103320, 103390, 103330, 103330, 103250, 103230, 103220, 103290, 103450, 
    103390, 103330, 103320, 103370, 103400, 103410, 103370, 103350, 103310, 
    103290, 103290, 103260, 103250, 103240, 103230, 103220, 103210, 103220, 
    103160, 103160, 103160, 103150, 103140, 103130, 103150, 103150, 103140, 
    103160, 103170, 103200, 103190, 103190, 103190, 103180, 103180, 103170, 
    103180, 103160, 103160, 103190, 103210, 103220, 103220, 103190, 103190, 
    103190, 103190, 103180, 103170, 103180, 103180, 103190, 103200, 103180, 
    103160, 103170, 103140, 103140, 103130, 103140, 103130, 103120, 103120, 
    103130, 103140, 103160, 103140, 103150, 103150, 103170, 103150, 103160, 
    103140, 103150, 103150, 103190, 103190, 103190, 103190, 103180, 103170, 
    103180, 103180, 103170, 103180, 103180, 103190, 103220, 103230, 103230, 
    103240, 103240, 103250, 103270, 103270, 103250, 103250, 103260, 103280, 
    103290, 103310, 103310, 103320, 103320, 103320, 103320, 103320, 103330, 
    103330, 103370, 103370, 103410, 103410, 103410, 103400, 103420, 103440, 
    103440, 103450, 103430, 103420, 103420, 103430, 103420, 103410, 103380, 
    103380, 103350, 103340, 103310, 103310, 103300, 103300, 103280, 103260, 
    103250, 103240, 103220, 103220, 103210, 103210, 103160, 103180, 103170, 
    103180, 103160, 103170, 103170, 103170, 103150, 103100, 103060, 103040, 
    103010, 102970, 102930, 102880, 102860, 102830, 102780, 102760, 102700, 
    102660, 102620, 102590, 102610, 102600, 102600, 102590, 102630, 102630, 
    102640, 102620, 102560, 102540, 102520, 102490, 102460, 102450, 102430, 
    102410, 102390, 102380, 102370, 102340, 102350, 102380, 102390, 102370, 
    102350, 102360, 102380, 102370, 102380, 102390, 102410, 102440, 102430, 
    102420, 102440, 102450, 102420, 102400, 102430, 102410, 102430, 102440, 
    102460, 102470, 102460, 102480, 102480, 102440, 102470, 102480, 102480, 
    102470, 102470, 102480, 102510, 102510, 102520, 102530, 102550, 102560, 
    102530, 102570, 102580, 102550, 102600, 102620, 102640, 102650, 102640, 
    102640, 102660, 102680, 102700, 102720, 102720, 102730, 102730, 102720, 
    102720, 102710, 102680, 102650, 102630, 102640, 102630, 102630, 102650, 
    102650, 102660, 102670, 102670, 102730, 102700, 102700, 102710, 102730, 
    102720, 102720, 102660, 102640, 102650, 102580, 102640, 102640, 102560, 
    102530, 102520, 102460, 102410, 102420, 102380, 102350, 102290, 102260, 
    102230, 102200, 102150, 102090, 102010, 102000, 101920, 101870, 101810, 
    101750, 101680, 101620, 101530, 101400, 101310, 101180, 101070, 101000, 
    100930, 100850, 100760, 100670, 100570, 100510, 100450, 100360, 100320, 
    100280, 100230, 100250, 100260, 100310, 100350, 100250, 100310, 100380, 
    100380, 100530, 100680, 100730, 100780, 100690, 100810, 100930, 101190, 
    101320, 101350, 101400, 101410, 101410, 101480, 101490, 101630, 101690, 
    101750, 101810, 101850, 101940, 102100, 102140, 102180, 102200, 102260, 
    102230, 102140, 102130, 102150, 102220, 102260, 102320, 102310, 102310, 
    102290, 102290, 102290, 102260, 102260, 102270, 102240, 102250, 102220, 
    102190, 102160, 102140, 102110, 102100, 102070, 102010, 101980, 101980, 
    102040, 101930, 101920, 101890, 101860, 101840, 101830, 101820, 101770, 
    101750, 101740, 101690, 101660, 101620, 101590, 101560, 101510, 101440, 
    101410, 101380, 101330, 101320, 101240, 101190, 101150, 101080, 101060, 
    101010, 100950, 100880, 100830, 100800, 100730, 100690, 100640, 100560, 
    100490, 100450, 100400, 100330, 100270, 100240, 100220, 100200, 100130, 
    100080, 100010, 99960, 99930, 99910, 99930, 100010, 100040, 100010, 
    99950, 99950, 99890, 99820, 99810, 99850, 99910, 99960, 100010, 100030, 
    100100, 100160, 100250, 100320, 100350, 100330, 100290, 100240, 100270, 
    100320, 100390, 100450, 100500, 100530, 100590, 100630, 100630, 100660, 
    100710, 100680, 100650, 100770, 100830, 100820, 100880, 100880, 100900, 
    100970, 101000, 101050, 101140, 101180, 101200, 101240, 101230, 101210, 
    101220, 101280, 101310, 101330, 101360, 101410, 101460, 101500, 101540, 
    101620, 101590, 101710, 101710, 101690, 101700, 101690, 101660, 101690, 
    101690, 101750, 101790, 101790, 101800, 101770, 101770, 101750, 101760, 
    101750, 101720, 101690, 101600, 101490, 101460, 101300, 101110, 100940, 
    100830, 100770, 100730, 100740, 100760, 100750, 100800, 100810, 100860, 
    100880, 100880, 100860, 100850, 100830, 100830, 100800, 100750, 100720, 
    100660, 100640, 100670, 100720, 100740, 100750, 100770, 100780, 100840, 
    100850, 100870, 100890, 100890, 100890, 100890, 100880, 100860, 100870, 
    100820, 100820, 100810, 100800, 100780, 100770, 100760, 100730, 100720, 
    100710, 100690, 100640, 100620, 100600, 100570, 100550, 100530, 100520, 
    100520, 100480, 100470, 100490, 100490, 100500, 100490, 100520, 100550, 
    100580, 100620, 100620, 100640, 100670, 100680, 100690, 100700, 100720, 
    100720, 100750, 100790, 100830, 100860, 100870, 100900, 100890, 100880, 
    100920, 100930, 100950, 100960, 101000, 101040, 101070, 101100, 101120, 
    101120, 101130, 101110, 101120, 101120, 101120, 101130, 101110, 101140, 
    101140, 101140, 101130, 101110, 101120, 101100, 101090, 101090, 101080, 
    101060, 101080, 101090, 101110, 101130, 101130, 101100, 101100, 101080, 
    101080, 101080, 101100, 101120, 101150, 101150, 101160, 101190, 101200, 
    101220, 101220, 101250, 101260, 101250, 101230, 101270, 101320, 101370, 
    101390, 101400, 101420, 101460, 101500, 101540, 101570, 101600, 101640, 
    101660, 101680, 101730, 101760, 101780, 101890, 101940, 101980, 102020, 
    102030, 102070, 102100, 102150, 102190, 102230, 102280, 102320, 102330, 
    102340, 102360, 102360, 102370, 102380, 102420, 102440, 102470, 102520, 
    102550, 102600, 102610, 102660, 102700, 102720, 102740, 102790, 102830, 
    102870, 102890, 102930, 102960, 103010, 103050, 103070, 103080, 103080, 
    103100, 103130, 103140, 103160, 103160, 103190, 103210, 103200, 103200, 
    103210, 103200, 103190, 103200, 103180, 103180, 103160, 103160, 103160, 
    103160, 103160, 103170, 103130, 103120, 103100, 103100, 103100, 103100, 
    103080, 103090, 103070, 103080, 103080, 103040, 103010, 102960, 102950, 
    102960, 102960, 102930, 102910, 102890, 102860, 102850, 102840, 102810, 
    102780, 102730, 102710, 102710, 102670, 102640, 102610, 102580, 102560, 
    102530, 102510, 102490, 102460, 102420, 102390, 102360, 102320, 102310, 
    102280, 102270, 102240, 102220, 102200, 102180, 102150, 102120, 102090, 
    102060, 102040, 102030, 102030, 102030, 102010, 101980, 101970, 101970, 
    101960, 101950, 101950, 101930, 101940, 101950, 101970, 101990, 101960, 
    102000, 102010, 102010, 102010, 101990, 101970, 101960, 101970, 102000, 
    101980, 102020, 101990, 102000, 101970, 101950, 102000, 101940, 101940, 
    101940, 101920, 101890, 101870, 101850, 101820, 101790, 101750, 101710, 
    101740, 101660, 101620, 101600, 101580, 101570, 101570, 101550, 101530, 
    101510, 101490, 101470, 101450, 101410, 101370, 101320, 101250, 101210, 
    101100, 101050, 100930, 100870, 100900, 100950, 100940, 100960, 100960, 
    100950, 100970, 100970, 100970, 100940, 100930, 100930, 100940, 100930, 
    100920, 100900, 100880, 100840, 100790, 100750, 100740, 100700, 100680, 
    100650, 100640, 100630, 100620, 100590, 100570, 100520, 100460, 100390, 
    100300, 100240, 100170, 100090, 100040, 99970, 99900, 99820, 99740, 
    99680, 99630, 99630, 99650, 99680, 99760, 99880, 99970, 100160, 100300, 
    100370, 100440, 100500, 100550, 100630, 100650, 100740, 100820, 100860, 
    100860, 100860, 100850, 100840, 100810, 100790, 100740, 100730, 100760, 
    100790, 100820, 100820, 100780, 100800, 100820, 100810, 100810, 100810, 
    100770, 100780, 100800, 100820, 100880, 100890, 100960, 100950, 101000, 
    101040, 101090, 101110, 101120, 101110, 101090, 101090, 101090, 101060, 
    101040, 100990, 100920, 100830, 100740, 100620, 100470, 100400, 100240, 
    100140, 100030, 99980, 99980, 99980, 100000, 100040, 100090, 100130, 
    100140, 100130, 100140, 100170, 100200, 100220, 100230, 100220, 100270, 
    100280, 100380, 100520, 100630, 100740, 100840, 100950, 101000, 101040, 
    101110, 101080, 101110, 101190, 101210, 101260, 101200, 101280, 101340, 
    101360, 101400, 101390, 101420, 101430, 101430, 101460, 101470, 101480, 
    101490, 101470, 101460, 101460, 101470, 101470, 101490, 101530, 101580, 
    101630, 101680, 101730, 101760, 101850, 101890, 101930, 101990, 102030, 
    102050, 102030, 102060, 102070, 102050, 102010, 101970, 101900, 101860, 
    101830, 101800, 101770, 101700, 101650, 101590, 101560, 101520, 101500, 
    101450, 101410, 101400, 101400, 101420, 101420, 101390, 101350, 101320, 
    101290, 101250, 101230, 101170, 101080, 101010, 100920, 100870, 100840, 
    100760, 100730, 100720, 100680, 100650, 100610, 100590, 100580, 100600, 
    100610, 100650, 100680, 100660, 100570, 100460, 100380, 100410, 100560, 
    100820, 100940, 101000, 101160, 101240, 101360, 101390, 101300, 101430, 
    101430, 101550, 101500, 101570, 101590, 101590, 101660, 101670, 101730, 
    101780, 101880, 101820, 101880, 101970, 102030, 102100, 102160, 102190, 
    102240, 102290, 102320, 102360, 102390, 102410, 102410, 102420, 102430, 
    102400, 102400, 102420, 102440, 102440, 102470, 102480, 102480, 102480, 
    102470, 102470, 102440, 102400, 102370, 102370, 102350, 102300, 102280, 
    102280, 102240, 102230, 102200, 102160, 102140, 102090, 102020, 101970, 
    101900, 101860, 101820, 101820, 101780, 101720, 101730, 101680, 101630, 
    101580, 101540, 101500, 101450, 101410, 101370, 101330, 101260, 101200, 
    101170, 101110, 101040, 101010, 100960, 100910, 100880, 100850, 100800, 
    100780, 100700, 100640, 100530, 100520, 100470, 100440, 100380, 100330, 
    100320, 100260, 100280, 100260, 100290, 100310, 100320, 100390, 100460, 
    100520, 100580, 100670, 100720, 100760, 100820, 100840, 100870, 100890, 
    100880, 100880, 100890, 100850, 100840, 100820, 100820, 100820, 100810, 
    100860, 100900, 100910, 100930, 100930, 100940, 100960, 100960, 100980, 
    100990, 101000, 101030, 101050, 101060, 101060, 101040, 101020, 101010, 
    101000, 100990, 100990, 101000, 101000, 100990, 100990, 100960, 100950, 
    100940, 100940, 100920, 100910, 100900, 100900, 100890, 100890, 100880, 
    100870, 100880, 100870, 100850, 100830, 100810, 100820, 100810, 100810, 
    100800, 100800, 100790, 100770, 100770, 100770, 100770, 100760, 100750, 
    100750, 100760, 100790, 100790, 100790, 100810, 100820, 100840, 100840, 
    100850, 100880, 100870, 100880, 100900, 100920, 100940, 100960, 100980, 
    100980, 101000, 101030, 101040, 101040, 101050, 101060, 101070, 101110, 
    101150, 101160, 101180, 101210, 101240, 101280, 101280, 101270, 101310, 
    101340, 101360, 101400, 101420, 101420, 101420, 101430, 101450, 101450, 
    101450, 101460, 101470, 101480, 101500, 101510, 101530, 101550, 101560, 
    101570, 101590, 101590, 101580, 101580, 101590, 101590, 101590, 101600, 
    101600, 101590, 101580, 101570, 101560, 101550, 101520, 101510, 101490, 
    101490, 101470, 101460, 101450, 101430, 101400, 101360, 101330, 101290, 
    101270, 101230, 101200, 101140, 101100, 101070, 101030, 101010, 100970, 
    100940, 100920, 100900, 100900, 100890, 100880, 100870, 100880, 100890, 
    100920, 100930, 100940, 100960, 100970, 101000, 101000, 101020, 101020, 
    101040, 101030, 101030, 101050, 101070, 101080, 101070, 101090, 101120, 
    101130, 101150, 101150, 101170, 101190, 101210, 101230, 101260, 101300, 
    101340, 101350, 101380, 101390, 101430, 101430, 101420, 101450, 101450, 
    101480, 101470, 101480, 101510, 101520, 101560, 101610, 101640, 101640, 
    101630, 101670, 101720, 101760, 101790, 101830, 101880, 101930, 101960, 
    101980, 102020, 102040, 102080, 102080, 102090, 102140, 102170, 102200, 
    102190, 102210, 102190, 102200, 102210, 102190, 102180, 102180, 102200, 
    102170, 102160, 102210, 102210, 102190, 102200, 102230, 102210, 102190, 
    102180, 102180, 102180, 102220, 102210, 102230, 102220, 102200, 102200, 
    102180, 102180, 102180, 102160, 102170, 102150, 102140, 102120, 102150, 
    102130, 102100, 102090, 102080, 102080, 102080, 102080, 102060, 102070, 
    102070, 102050, 102090, 102110, 102100, 102090, 102050, 102000, 101940, 
    101890, 101790, 101770, 101740, 101690, 101680, 101610, 101610, 101600, 
    101590, 101530, 101450, 101400, 101400, 101360, 101340, 101370, 101360, 
    101360, 101370, 101300, 101300, 101280, 101250, 101220, 101160, 101100, 
    101070, 101080, 101030, 100990, 100980, 100910, 100870, 100830, 100780, 
    100730, 100680, 100590, 100520, 100480, 100430, 100380, 100350, 100310, 
    100270, 100260, 100230, 100250, 100290, 100270, 100290, 100280, 100260, 
    100230, 100180, 100120, 100050, 99990, 99910, 99870, 99810, 99750, 99700, 
    99680, 99650, 99600, 99560, 99550, 99540, 99530, 99510, 99520, 99570, 
    99600, 99650, 99720, 99790, 99890, 99970, 100110, 100190, 100300, 100380, 
    100490, 100560, 100630, 100700, 100760, 100790, 100810, 100820, 100840, 
    100840, 100850, 100820, 100850, 100830, 100830, 100830, 100810, 100780, 
    100770, 100740, 100690, 100630, 100530, 100460, 100370, 100350, 100380, 
    100360, 100410, 100400, 100410, 100440, 100510, 100570, 100640, 100690, 
    100760, 100770, 100880, 100910, 100950, 100990, 100990, 100980, 100960, 
    100910, 100790, 100750, 100700, 100550, 100480, 100360, 100250, 100140, 
    100060, 99930, 99830, 99760, 99720, 99620, 99610, 99680, 99790, 99810, 
    99960, 100070, 100170, 100290, 100410, 100560, 100650, 100730, 100810, 
    100900, 100990, 101040, 101120, 101180, 101220, 101290, 101390, 101450, 
    101480, 101510, 101550, 101620, 101670, 101710, 101720, 101740, 101750, 
    101740, 101750, 101730, 101660, 101570, 101510, 101410, 101260, 101070, 
    100900, 100770, 100510, 100360, 100150, 99980, 99930, 99870, 99860, 
    99890, 99960, 100060, 100170, 100300, 100450, 100570, 100670, 100730, 
    100830, 100930, 101000, 101080, 101190, 101290, 101380, 101460, 101560, 
    101640, 101710, 101750, 101860, 101880, 101900, 101890, 101910, 101900, 
    101870, 101850, 101770, 101700, 101640, 101550, 101420, 101340, 101230, 
    101200, 101170, 101250, 101360, 101420, 101560, 101670, 101860, 102170, 
    102270, 102380, 102510, 102560, 102640, 102720, 102800, 102800, 102830, 
    102860, 102890, 102900, 102880, 102820, 102790, 102780, 102740, 102720, 
    102680, 102640, 102610, 102520, 102490, 102450, 102370, 102270, 102220, 
    102130, 102100, 102080, 102060, 102020, 101990, 101950, 101940, 101910, 
    101860, 101810, 101770, 101750, 101730, 101740, 101720, 101710, 101690, 
    101730, 101670, 101670, 101660, 101620, 101600, 101580, 101600, 101600, 
    101590, 101610, 101640, 101660, 101630, 101650, 101690, 101700, 101710, 
    101740, 101720, 101730, 101770, 101770, 101730, 101700, 101710, 101700, 
    101640, 101570, 101590, 101550, 101530, 101430, 101410, 101470, 101470, 
    101430, 101370, 101290, 101230, 101180, 101090, 101000, 101040, 101080, 
    101090, 101060, 101050, 101060, 101060, 101000, 100990, 100970, 100980, 
    100950, 100980, 100980, 100960, 100950, 100920, 100870, 100830, 100800, 
    100810, 100730, 100640, 100620, 100610, 100630, 100650, 100650, 100620, 
    100580, 100560, 100520, 100480, 100450, 100390, 100310, 100320, 100350, 
    100330, 100300, 100310, 100310, 100280, 100270, 100210, 100230, 100180, 
    100120, 100140, 100190, 100250, 100170, 100110, 100150, 100180, 100160, 
    100130, 100080, 100170, 100150, 100200, 100280, 100340, 100370, 100430, 
    100450, 100440, 100440, 100440, 100440, 100400, 100330, 100240, 100200, 
    100200, 100130, 100130, 100140, 100090, 100070, 100050, 100060, 100040, 
    100030, 100040, 100080, 100140, 100190, 100250, 100280, 100320, 100380, 
    100430, 100470, 100520, 100560, 100600, 100650, 100690, 100720, 100760, 
    100780, 100790, 100820, 100840, 100860, 100860, 100860, 100860, 100880, 
    100890, 100900, 100910, 100930, 100940, 100940, 100940, 100930, 100920, 
    100910, 100890, 100910, 100920, 100920, 100920, 100950, 100970, 101000, 
    101010, 101040, 101060, 101140, 101160, 101220, 101270, 101300, 101340, 
    101370, 101390, 101430, 101440, 101430, 101420, 101400, 101400, 101410, 
    101420, 101420, 101420, 101370, 101390, 101340, 101300, 101240, 101210, 
    101150, 101100, 101070, 101050, 101020, 100970, 100950, 100900, 100840, 
    100800, 100790, 100750, 100710, 100740, 100740, 100730, 100740, 100730, 
    100740, 100740, 100750, 100740, 100750, 100780, 100820, 100880, 100920, 
    100940, 100980, 101000, 101010, 101010, 100980, 100950, 100900, 100870, 
    100800, 100760, 100700, 100660, 100610, 100550, 100490, 100410, 100350, 
    100310, 100280, 100250, 100240, 100240, 100270, 100310, 100370, 100420, 
    100480, 100510, 100560, 100590, 100640, 100670, 100710, 100740, 100760, 
    100780, 100800, 100840, 100880, 100930, 101000, 101050, 101080, 101100, 
    101130, 101180, 101240, 101290, 101340, 101340, 101360, 101370, 101360, 
    101320, 101300, 101280, 101250, 101240, 101200, 101200, 101160, 101160, 
    101150, 101150, 101170, 101170, 101190, 101220, 101260, 101310, 101350, 
    101410, 101460, 101540, 101590, 101620, 101660, 101700, 101730, 101770, 
    101790, 101830, 101850, 101900, 101930, 101960, 101980, 101960, 101950, 
    101960, 101960, 101990, 102020, 102020, 102050, 102090, 102100, 102070, 
    102110, 102110, 102130, 102130, 102120, 102120, 102120, 102110, 102120, 
    102120, 102110, 102100, 102110, 102110, 102100, 102120, 102120, 102140, 
    102170, 102220, 102250, 102250, 102270, 102290, 102300, 102290, 102290, 
    102290, 102280, 102260, 102270, 102250, 102220, 102200, 102210, 102180, 
    102150, 102120, 102100, 102070, 102030, 102000, 101990, 101950, 101880, 
    101830, 101780, 101710, 101670, 101630, 101540, 101470, 101410, 101370, 
    101310, 101260, 101190, 101140, 101090, 101040, 101010, 100990, 100980, 
    100970, 100960, 100920, 100940, 100930, 100930, 100930, 100940, 100940, 
    100920, 100900, 100850, 100830, 100790, 100810, 100810, 100810, 100800, 
    100770, 100740, 100700, 100670, 100650, 100630, 100570, 100550, 100520, 
    100510, 100490, 100480, 100460, 100470, 100450, 100470, 100450, 100450, 
    100450, 100410, 100370, 100340, 100280, 100270, 100240, 100220, 100200, 
    100200, 100190, 100180, 100150, 100120, 100130, 100150, 100190, 100210, 
    100240, 100230, 100230, 100230, 100200, 100220, 100160, 100220, 100300, 
    100360, 100420, 100450, 100500, 100570, 100640, 100630, 100740, 100840, 
    100920, 100970, 101080, 101130, 101170, 101200, 101290, 101330, 101390, 
    101430, 101480, 101510, 101500, 101520, 101530, 101550, 101550, 101560, 
    101550, 101530, 101510, 101490, 101480, 101470, 101460, 101380, 101370, 
    101330, 101340, 101350, 101330, 101260, 101270, 101210, 101240, 101260, 
    101120, 101180, 101140, 101040, 101060, 100950, 100900, 100900, 100780, 
    100700, 100690, 100620, 100590, 100590, 100570, 100520, 100580, 100570, 
    100540, 100510, 100500, 100490, 100480, 100460, 100440, 100400, 100390, 
    100370, 100330, 100250, 100160, 99990, 99910, 99850, 99820, 99690, 99580, 
    99560, 99340, 99230, 99120, 98940, 98770, 98690, 98540, 98380, 98260, 
    98130, 98070, 98050, 98060, 98110, 98120, 98090, 98170, 98290, 98390, 
    98460, 98510, 98570, 98630, 98680, 98580, 98750, 98880, 98950, 99010, 
    99100, 99240, 99420, 99430, 99610, 99700, 99830, 99960, 100100, 100210, 
    100330, 100410, 100500, 100590, 100700, 100780, 100810, 100900, 100950, 
    101020, 101050, 101110, 101180, 101240, 101280, 101320, 101370, 101400, 
    101430, 101440, 101450, 101450, 101470, 101480, 101500, 101500, 101520, 
    101520, 101530, 101540, 101560, 101560, 101550, 101560, 101570, 101580, 
    101590, 101600, 101620, 101620, 101630, 101640, 101640, 101640, 101630, 
    101600, 101610, 101580, 101590, 101570, 101540, 101520, 101500, 101460, 
    101410, 101320, 101240, 101250, 101210, 101190, 101190, 101130, 101040, 
    100960, 100930, 100940, 100890, 100830, 100740, 100720, 100680, 100650, 
    100600, 100560, 100510, 100480, 100470, 100480, 100460, 100460, 100460, 
    100440, 100470, 100460, 100460, 100440, 100410, 100370, 100330, 100310, 
    100230, 100180, 100090, 100010, 99950, 99920, 99860, 99830, 99760, 99760, 
    99730, 99710, 99620, 99610, 99660, 99660, 99660, 99650, 99640, 99630, 
    99620, 99620, 99590, 99610, 99590, 99600, 99620, 99620, 99650, 99680, 
    99720, 99760, 99810, 99860, 99920, 99950, 100000, 100060, 100130, 100180, 
    100220, 100280, 100330, 100370, 100430, 100490, 100540, 100610, 100670, 
    100710, 100750, 100780, 100790, 100810, 100810, 100840, 100880, 100950, 
    100990, 101030, 101070, 101130, 101180, 101190, 101250, 101320, 101350, 
    101420, 101430, 101420, 101440, 101480, 101460, 101440, 101440, 101420, 
    101350, 101330, 101320, 101340, 101340, 101340, 101290, 101270, 101240, 
    101180, 101100, 100980, 100910, 100780, 100750, 100730, 100660, 100590, 
    100600, 100550, 100440, 100420, 100400, 100370, 100330, 100320, 100360, 
    100350, 100360, 100340, 100280, 100270, 100270, 100190, 100160, 100130, 
    100080, 100020, 100000, 99980, 99970, 99930, 99910, 99860, 99830, 99810, 
    99810, 99840, 99840, 99870, 99920, 99960, 100010, 100030, 100100, 100160, 
    100210, 100290, 100350, 100380, 100470, 100550, 100670, 100750, 100830, 
    100890, 101000, 101070, 101110, 101150, 101200, 101240, 101260, 101290, 
    101320, 101300, 101310, 101300, 101290, 101280, 101260, 101250, 101220, 
    101190, 101180, 101170, 101120, 101070, 101040, 101010, 100950, 100880, 
    100840, 100810, 100780, 100670, 100500, 100340, 100250, 100190, 100080, 
    99910, 99730, 99710, 99700, 99720, 99650, 99700, 99700, 99720, 99770, 
    99810, 99820, 99830, 99870, 99920, 99980, 100060, 100160, 100260, 100360, 
    100440, 100500, 100560, 100630, 100660, 100710, 100770, 100780, 100810, 
    100830, 100850, 100870, 100920, 100960, 100980, 101010, 101040, 101050, 
    101070, 101080, 101100, 101120, 101120, 101120, 101140, 101150, 101160, 
    101160, 101150, 101150, 101140, 101150, 101170, 101150, 101170, 101190, 
    101200, 101220, 101250, 101280, 101320, 101320, 101340, 101350, 101380, 
    101390, 101390, 101400, 101420, 101430, 101460, 101450, 101430, 101460, 
    101460, 101440, 101440, 101410, 101420, 101410, 101410, 101420, 101430, 
    101440, 101440, 101420, 101380, 101370, 101330, 101270, 101310, 101390, 
    101340, 101270, 101180, 101230, 101170, 100930, 101050, 101020, 100970, 
    100950, 100830, 100720, 100690, 100520, 100490, 100450, 100330, 100290, 
    100170, 100120, 100040, 100040, 100010, 99960, 99940, 99900, 99880, 
    100060, 100030, 100000, 99950, 99960, 99890, 99900, 99840, 99840, 99820, 
    99800, 99790, 99770, 99740, 99730, 99720, 99690, 99650, 99620, 99590, 
    99550, 99560, 99520, 99490, 99480, 99460, 99430, 99400, 99400, 99380, 
    99390, 99350, 99330, 99350, 99350, 99360, 99330, 99340, 99320, 99300, 
    99280, 99250, 99220, 99180, 99150, 99130, 99120, 99100, 99070, 99050, 
    99030, 99010, 98990, 98970, 98960, 98970, 99000, 99020, 99050, 99110, 
    99160, 99210, 99240, 99260, 99310, 99340, 99350, 99380, 99420, 99470, 
    99500, 99540, 99540, 99590, 99620, 99620, 99670, 99680, 99680, 99690, 
    99680, 99710, 99710, 99740, 99740, 99800, 99810, 99810, 99800, 99820, 
    99830, 99840, 99820, 99810, 99840, 99830, 99840, 99830, 99820, 99810, 
    99780, 99760, 99760, 99800, 99830, 99860, 99890, 99920, 99940, 99960, 
    99990, 99990, 100010, 100020, 100040, 100040, 100070, 100070, 100100, 
    100120, 100160, 100200, 100100, 100060, 100110, 100190, 100270, 100300, 
    100300, 100390, 100410, 100420, 100490, 100550, 100510, 100550, 100580, 
    100600, 100620, 100610, 100590, 100560, 100530, 100470, 100450, 100450, 
    100430, 100410, 100360, 100320, 100310, 100290, 100320, 100310, 100290, 
    100290, 100290, 100260, 100270, 100270, 100240, 100260, 100280, 100260, 
    100260, 100240, 100210, 100210, 100230, 100290, 100330, 100390, 100450, 
    100540, 100600, 100670, 100720, 100770, 100820, 100880, 100940, 100980, 
    101010, 101030, 101070, 101080, 101090, 101100, 101100, 101120, 101170, 
    101210, 101210, 101180, 101170, 101200, 101210, 101200, 101210, 101180, 
    101190, 101210, 101270, 101320, 101350, 101370, 101370, 101420, 101440, 
    101460, 101450, 101470, 101470, 101440, 101420, 101440, 101450, 101440, 
    101440, 101410, 101440, 101430, 101430, 101390, 101350, 101300, 101320, 
    101340, 101360, 101350, 101320, 101320, 101320, 101320, 101310, 101260, 
    101250, 101270, 101240, 101240, 101220, 101220, 101220, 101230, 101240, 
    101220, 101220, 101200, 101210, 101220, 101230, 101240, 101260, 101280, 
    101270, 101290, 101300, 101290, 101300, 101270, 101280, 101300, 101310, 
    101300, 101290, 101300, 101310, 101320, 101300, 101320, 101340, 101360, 
    101350, 101370, 101410, 101450, 101500, 101540, 101540, 101570, 101590, 
    101630, 101640, 101630, 101650, 101680, 101690, 101690, 101690, 101700, 
    101710, 101730, 101720, 101690, 101690, 101690, 101700, 101680, 101680, 
    101660, 101650, 101600, 101550, 101520, 101470, 101440, 101390, 101360, 
    101300, 101290, 101240, 101220, 101190, 101190, 101210, 101200, 101150, 
    101110, 101070, 101060, 101030, 101000, 100990, 100970, 100930, 100910, 
    100840, 100810, 100740, 100680, 100690, 100620, 100650, 100620, 100600, 
    100550, 100490, 100480, 100450, 100430, 100420, 100400, 100390, 100390, 
    100380, 100360, 100370, 100360, 100410, 100450, 100530, 100560, 100560, 
    100600, 100630, 100610, 100550, 100530, 100520, 100470, 100420, 100390, 
    100350, 100310, 100290, 100260, 100250, 100230, 100210, 100180, 100170, 
    100130, 100040, 100000, 100020, 99970, 99940, 99880, 99840, 99820, 99790, 
    99780, 99780, 99730, 99720, 99700, 99730, 99740, 99770, 99840, 99910, 
    99980, 100060, 100130, 100210, 100270, 100340, 100400, 100450, 100450, 
    100440, 100460, 100480, 100470, 100490, 100490, 100520, 100550, 100580, 
    100610, 100650, 100710, 100680, 100700, 100760, 100740, 100710, 100690, 
    100670, 100640, 100570, 100580, 100500, 100420, 100350, 100260, 100140, 
    100050, 99970, 99890, 99880, 99860, 99870, 99900, 99960, 100040, 100090, 
    100120, 100170, 100220, 100260, 100300, 100360, 100420, 100490, 100550, 
    100600, 100640, 100710, 100770, 100800, 100850, 100890, 100920, 100920, 
    100900, 100930, 100920, 100890, 100860, 100810, 100720, 100710, 100670, 
    100620, 100560, 100520, 100480, 100420, 100340, 100290, 100240, 100210, 
    100150, 100150, 100150, 100190, 100250, 100300, 100390, 100460, 100570, 
    100650, 100730, 100780, 100810, 100880, 100930, 100960, 101020, 101050, 
    101090, 101120, 101110, 101120, 101120, 101110, 101070, 101080, 101050, 
    101000, 100930, 100920, 100860, 100840, 100750, 100680, 100600, 100550, 
    100490, 100460, 100470, 100420, 100420, 100430, 100440, 100460, 100460, 
    100490, 100520, 100510, 100550, 100590, 100660, 100710, 100740, 100830, 
    100880, 100940, 101000, 101090, 101140, 101170, 101240, 101270, 101310, 
    101350, 101390, 101460, 101480, 101490, 101520, 101550, 101560, 101550, 
    101560, 101560, 101580, 101560, 101570, 101590, 101610, 101630, 101650, 
    101700, 101740, 101760, 101800, 101850, 101880, 101920, 101960, 101990, 
    102010, 102040, 102070, 102090, 102070, 102040, 102060, 102040, 102040, 
    101990, 101960, 101920, 101880, 101880, 101830, 101790, 101750, 101750, 
    101740, 101690, 101700, 101710, 101720, 101710, 101690, 101700, 101690, 
    101640, 101600, 101600, 101550, 101490, 101440, 101360, 101280, 101020, 
    101090, 100960, 100830, 100690, 100580, 100530, 100430, 100330, 100290, 
    100250, 100230, 100230, 100210, 100250, 100270, 100270, 100300, 100300, 
    100250, 100230, 100210, 100210, 100230, 100250, 100270, 100280, 100310, 
    100320, 100320, 100330, 100360, 100410, 100380, 100430, 100470, 100510, 
    100560, 100580, 100590, 100640, 100670, 100690, 100720, 100770, 100800, 
    100940, 100900, 100970, 101010, 101050, 101120, 101150, 101180, 101200, 
    101210, 101200, 101230, 101230, 101220, 101190, 101160, 101130, 101120, 
    101090, 101040, 101010, 101000, 100970, 100900, 100870, 100810, 100780, 
    100780, 100760, 100760, 100740, 100710, 100700, 100650, 100600, 100600, 
    100580, 100590, 100570, 100540, 100530, 100540, 100520, 100500, 100520, 
    100530, 100560, 100510, 100520, 100500, 100510, 100510, 100450, 100440, 
    100420, 100400, 100370, 100350, 100350, 100320, 100310, 100290, 100290, 
    100280, 100270, 100270, 100260, 100250, 100250, 100250, 100240, 100230, 
    100250, 100280, 100290, 100320, 100350, 100390, 100410, 100470, 100490, 
    100510, 100590, 100680, 100740, 100800, 100910, 100970, 101010, 101040, 
    101090, 101130, 101130, 101100, 101090, 101070, 101040, 100980, 100940, 
    100920, 100900, 100860, 100800, 100760, 100700, 100640, 100620, 100580, 
    100580, 100610, 100580, 100540, 100590, 100630, 100650, 100680, 100700, 
    100710, 100750, 100810, 100850, 100880, 100920, 100890, 100910, 100960, 
    100990, 100990, 100980, 101000, 101030, 101060, 101060, 101130, 101160, 
    101210, 101270, 101320, 101390, 101420, 101460, 101500, 101540, 101570, 
    101590, 101600, 101550, 101510, 101500, 101440, 101420, 101350, 101280, 
    101240, 101180, 101170, 101130, 101140, 101140, 101170, 101160, 101170, 
    101200, 101210, 101190, 101190, 101220, 101290, 101290, 101340, 101380, 
    101420, 101420, 101430, 101430, 101470, 101480, 101450, 101450, 101430, 
    101430, 101390, 101420, 101450, 101500, 101530, 101520, 101550, 101570, 
    101600, 101650, 101680, 101710, 101780, 101850, 101870, 101920, 101950, 
    101960, 101970, 101990, 102030, 102070, 102110, 102150, 102190, 102270, 
    102290, 102330, 102300, 102360, 102340, 102380, 102380, 102350, 102340, 
    102350, 102350, 102360, 102340, 102300, 102290, 102310, 102250, 102210, 
    102170, 102160, 102100, 102100, 102080, 102080, 102080, 102060, 102070, 
    102040, 102010, 102020, 102000, 101960, 101960, 101960, 101950, 101950, 
    101940, 101930, 101940, 101930, 101890, 101850, 101820, 101830, 101840, 
    101870, 101860, 101880, 101910, 101920, 101940, 101950, 102000, 101980, 
    101950, 101950, 102030, 102020, 102110, 102130, 102170, 102220, 102200, 
    102240, 102280, 102350, 102440, 102530, 102470, 102490, 102520, 102530, 
    102560, 102600, 102640, 102640, 102620, 102640, 102640, 102640, 102620, 
    102610, 102610, 102610, 102610, 102600, 102560, 102550, 102530, 102510, 
    102480, 102460, 102430, 102430, 102390, 102370, 102370, 102360, 102330, 
    102280, 102240, 102240, 102210, 102170, 102140, 102110, 102060, 102040, 
    102020, 102000, 101970, 101940, 101910, 101870, 101840, 101790, 101770, 
    101750, 101730, 101720, 101710, 101710, 101710, 101660, 101630, 101650, 
    101610, 101590, 101590, 101550, 101560, 101540, 101530, 101540, 101500, 
    101480, 101500, 101530, 101570, 101590, 101610, 101640, 101660, 101660, 
    101670, 101670, 101660, 101610, 101570, 101470, 101400, 101320, 101340, 
    101300, 101310, 101230, 101080, 101020, 101000, 101010, 100960, 100960, 
    100890, 100840, 100810, 100740, 100720, 100650, 100570, 100490, 100420, 
    100400, 100480, 100390, 100340, 100320, 100280, 100280, 100280, 100180, 
    100090, 100010, 99950, 99850, 99760, 99730, 99660, 99650, 99600, 99580, 
    99590, 99530, 99580, 99560, 99540, 99570, 99530, 99530, 99530, 99500, 
    99470, 99520, 99510, 99520, 99640, 99660, 99720, 99770, 99810, 99840, 
    99870, 99940, 99890, 99890, 99880, 99870, 99900, 99920, 99960, 99990, 
    100030, 100060, 100130, 100150, 100150, 100160, 100190, 100220, 100250, 
    100280, 100280, 100280, 100290, 100320, 100340, 100330, 100340, 100360, 
    100390, 100430, 100460, 100480, 100490, 100500, 100530, 100550, 100560, 
    100570, 100580, 100590, 100610, 100630, 100650, 100680, 100700, 100730, 
    100720, 100740, 100750, 100750, 100760, 100780, 100790, 100850, 100890, 
    100920, 100930, 100950, 100970, 101010, 101020, 101040, 101050, 101050, 
    101070, 101130, 101150, 101130, 101140, 101120, 101120, 101110, 101120, 
    101120, 101100, 101080, 101060, 101080, 101080, 101070, 101080, 101020, 
    101020, 101000, 101010, 101010, 101040, 101000, 100970, 100910, 100890, 
    100840, 100820, 100810, 100760, 100710, 100700, 100690, 100690, 100630, 
    100630, 100620, 100640, 100680, 100680, 100680, 100690, 100680, 100680, 
    100690, 100710, 100680, 100620, 100680, 100710, 100670, 100670, 100630, 
    100670, 100700, 100660, 100640, 100620, 100580, 100580, 100580, 100580, 
    100590, 100600, 100630, 100610, 100590, 100560, 100560, 100520, 100480, 
    100460, 100470, 100480, 100480, 100480, 100480, 100460, 100460, 100470, 
    100450, 100430, 100430, 100430, 100400, 100390, 100390, 100410, 100480, 
    100500, 100500, 100550, 100580, 100610, 100600, 100580, 100580, 100630, 
    100680, 100650, 100640, 100660, 100690, 100710, 100740, 100720, 100760, 
    100760, 100800, 100810, 100830, 100870, 100910, 100930, 100900, 100910, 
    100920, 100930, 100930, 100930, 100950, 100960, 100980, 100990, 101000, 
    101030, 101050, 101060, 101060, 101090, 101120, 101130, 101150, 101160, 
    101170, 101180, 101180, 101190, 101200, 101190, 101160, 101180, 101180, 
    101200, 101210, 101210, 101180, 101180, 101190, 101180, 101180, 101160, 
    101130, 101110, 101100, 101100, 101060, 101050, 101020, 100980, 100950, 
    100930, 100880, 100850, 100820, 100760, 100710, 100610, 100580, 100520, 
    100390, 100190, 100030, 99900, 99800, 99640, 99430, 99320, 99220, 99040, 
    98880, 98760, 98760, 98850, 98870, 98950, 99020, 99040, 99050, 99070, 
    99080, 99060, 99080, 99080, 99080, 99090, 99080, 99040, 99020, 98980, 
    98960, 98910, 98920, 98890, 98890, 98870, 98860, 98850, 98850, 98880, 
    98890, 98900, 98910, 98910, 98900, 98880, 98830, 98720, 98730, 98730, 
    98730, 98750, 98780, 98810, 98750, 98800, 98830, 98850, 98780, 98790, 
    98760, 98820, 98880, 98830, 98860, 98950, 98970, 98950, 99010, 98960, 
    98940, 98980, 99010, 99040, 99020, 98980, 98980, 98970, 99010, 99000, 
    99050, 99120, 99110, 99150, 99190, 99180, 99170, 99220, 99260, 99250, 
    99280, 99280, 99280, 99310, 99320, 99410, 99440, 99450, 99460, 99490, 
    99530, 99590, 99640, 99680, 99740, 99770, 99810, 99840, 99910, 100000, 
    100040, 100100, 100140, 100180, 100240, 100290, 100330, 100380, 100440, 
    100470, 100500, 100540, 100590, 100640, 100660, 100690, 100710, 100750, 
    100800, 100810, 100830, 100860, 100880, 100900, 100930, 100970, 100990, 
    100970, 101010, 100960, 100960, 100970, 100920, 100930, 100910, 100970, 
    100950, 100940, 100890, 100880, 100910, 100900, 100890, 100870, 100920, 
    100880, 100880, 100890, 100880, 100870, 100840, 100840, 100820, 100790, 
    100800, 100840, 100860, 100870, 100900, 100890, 100950, 100970, 100950, 
    100960, 100940, 100900, 100890, 100880, 100910, 100940, 100940, 100920, 
    100920, 100870, 100810, 100800, 100760, 100740, 100660, 100620, 100540, 
    100460, 100410, 100330, 100240, 100130, 100070, 99980, 99890, 99840, 
    99790, 99730, 99700, 99660, 99650, 99640, 99650, 99670, 99700, 99730, 
    99770, 99820, 99880, 99950, 100030, 100080, 100150, 100220, 100310, 
    100360, 100410, 100450, 100490, 100570, 100610, 100660, 100700, 100720, 
    100750, 100780, 100800, 100820, 100840, 100860, 100860, 100890, 100890, 
    100880, 100870, 100880, 100860, 100860, 100870, 100880, 100860, 100840, 
    100850, 100910, 100920, 100930, 100950, 100980, 101020, 101040, 101070, 
    101110, 101130, 101150, 101180, 101200, 101250, 101270, 101300, 101320, 
    101360, 101400, 101420, 101450, 101470, 101460, 101450, 101430, 101400, 
    101380, 101360, 101320, 101300, 101300, 101300, 101280, 101280, 101250, 
    101250, 101250, 101250, 101250, 101230, 101220, 101210, 101180, 101150, 
    101100, 101020, 100960, 100830, 100770, 100710, 100610, 100550, 100400, 
    100310, 100210, 100130, 100010, 99860, 99720, 99550, 99380, 99250, 99150, 
    99110, 99080, 99040, 99130, 99120, 99100, 99120, 99100, 98980, 98840, 
    98800, 98810, 98750, 98760, 98790, 98810, 98850, 98860, 98970, 99080, 
    99210, 99360, 99500, 99690, 99830, 99830, 99980, 100190, 100380, 100510, 
    100580, 100670, 100740, 100830, 100910, 100970, 101050, 101120, 101180, 
    101260, 101300, 101320, 101320, 101310, 101310, 101310, 101300, 101270, 
    101220, 101170, 101120, 101080, 101020, 101020, 100980, 100950, 100940, 
    100880, 100860, 100820, 100790, 100750, 100660, 100620, 100550, 100480, 
    100370, 100280, 100240, 100190, 100160, 100100, 100050, 100020, 99980, 
    99940, 99910, 99900, 99860, 99840, 99850, 99830, 99820, 99800, 99800, 
    99830, 99750, 99630, 99590, 99460, 99350, 99240, 99150, 99110, 99050, 
    99050, 99050, 99130, 99220, 99330, 99470, 99600, 99750, 99880, 99980, 
    100080, 100190, 100330, 100450, 100560, 100670, 100770, 100850, 100930, 
    101050, 101120, 101200, 101280, 101360, 101410, 101460, 101500, 101500, 
    101500, 101510, 101520, 101550, 101550, 101570, 101630, 101680, 101710, 
    101740, 101720, 101750, 101730, 101710, 101640, 101580, 101550, 101470, 
    101400, 101330, 101280, 101230, 101170, 101090, 100970, 100930, 100850, 
    100790, 100720, 100670, 100640, 100640, 100660, 100710, 100750, 100800, 
    100850, 100910, 100990, 101080, 101190, 101240, 101290, 101330, 101380, 
    101410, 101480, 101510, 101530, 101570, 101590, 101610, 101630, 101640, 
    101680, 101740, 101760, 101740, 101750, 101730, 101680, 101670, 101630, 
    101600, 101550, 101500, 101480, 101430, 101420, 101420, 101420, 101420, 
    101440, 101460, 101440, 101460, 101470, 101490, 101510, 101510, 101500, 
    101530, 101560, 101530, 101520, 101510, 101480, 101450, 101380, 101340, 
    101350, 101280, 101250, 101180, 101180, 101160, 101130, 101110, 101100, 
    101120, 101130, 101150, 101140, 101160, 101190, 101200, 101230, 101240, 
    101270, 101300, 101330, 101370, 101370, 101420, 101440, 101480, 101490, 
    101510, 101520, 101520, 101540, 101590, 101600, 101620, 101650, 101640, 
    101650, 101640, 101680, 101720, 101730, 101750, 101770, 101780, 101810, 
    101810, 101820, 101830, 101860, 101870, 101890, 101900, 101920, 101910, 
    101930, 101930, 101930, 101910, 101920, 101930, 101940, 101940, 101900, 
    101920, 101940, 101890, 101850, 101880, 101890, 101840, 101780, 101770, 
    101720, 101690, 101670, 101650, 101610, 101560, 101530, 101500, 101490, 
    101480, 101430, 101390, 101360, 101380, 101340, 101320, 101300, 101310, 
    101340, 101350, 101310, 101290, 101250, 101220, 101200, 101170, 101110, 
    101080, 101030, 100960, 100900, 100860, 100810, 100740, 100670, 100570, 
    100500, 100430, 100380, 100340, 100320, 100280, 100240, 100200, 100170, 
    100130, 100100, 100050, 100020, 99990, 99970, 99990, 100020, 100040, 
    100040, 100010, 99990, 99980, 99960, 99940, 99960, 99980, 100020, 100090, 
    100170, 100230, 100290, 100360, 100410, 100500, 100540, 100600, 100640, 
    100700, 100770, 100840, 100890, 100940, 100970, 100980, 101010, 101050, 
    101080, 101100, 101120, 101100, 101140, 101130, 101170, 101210, 101190, 
    101200, 101190, 101160, 101180, 101210, 101200, 101190, 101220, 101230, 
    101260, 101290, 101320, 101360, 101410, 101440, 101510, 101550, 101580, 
    101590, 101620, 101680, 101700, 101730, 101800, 101820, 101820, 101840, 
    101850, 101880, 101900, 101910, 101930, 101930, 101920, 101930, 101920, 
    101910, 101890, 101890, 101890, 101890, 101890, 101880, 101880, 101870, 
    101840, 101820, 101800, 101770, 101750, 101730, 101690, 101660, 101650, 
    101610, 101580, 101570, 101540, 101510, 101480, 101460, 101450, 101440, 
    101430, 101410, 101400, 101400, 101400, 101400, 101400, 101410, 101410, 
    101420, 101440, 101440, 101450, 101460, 101460, 101460, 101450, 101480, 
    101490, 101510, 101510, 101510, 101510, 101510, 101550, 101540, 101550, 
    101540, 101540, 101540, 101550, 101560, 101570, 101560, 101560, 101580, 
    101580, 101570, 101550, 101550, 101550, 101540, 101530, 101490, 101470, 
    101460, 101440, 101420, 101420, 101410, 101390, 101360, 101340, 101320, 
    101300, 101280, 101280, 101260, 101260, 101210, 101210, 101190, 101150, 
    101120, 101030, 101010, 100970, 100930, 100910, 100850, 100840, 100820, 
    100810, 100770, 100750, 100740, 100710, 100700, 100680, 100680, 100670, 
    100650, 100650, 100660, 100670, 100640, 100610, 100600, 100540, 100500, 
    100490, 100490, 100480, 100480, 100480, 100420, 100370, 100380, 100350, 
    100420, 100430, 100440, 100490, 100550, 100550, 100520, 100520, 100570, 
    100500, 100450, 100400, 100400, 100380, 100390, 100380, 100330, 100290, 
    100330, 100280, 100250, 100150, 100080, 99960, 99920, 99820, 99600, 
    99450, 99380, 99300, 99330, 99290, 99010, 99030, 99030, 98930, 98780, 
    98620, 98550, 98340, 98220, 98230, 98220, 98280, 98290, 98250, 98250, 
    98230, 98150, 98160, 98160, 98200, 98160, 98150, 98090, 98040, 97980, 
    98000, 97940, 97930, 97960, 97920, 97960, 97970, 97950, 97930, 97930, 
    97900, 97890, 97860, 97840, 97830, 97850, 97860, 97890, 97890, 97900, 
    97900, 97890, 97900, 97890, 97880, 97870, 97860, 97860, 97870, 97900, 
    97920, 97960, 97950, 97970, 98030, 98090, 98130, 98150, 98170, 98220, 
    98240, 98300, 98330, 98390, 98420, 98450, 98460, 98480, 98500, 98530, 
    98550, 98550, 98560, 98590, 98620, 98630, 98650, 98650, 98670, 98680, 
    98690, 98700, 98700, 98710, 98740, 98780, 98830, 98880, 98910, 98940, 
    98950, 98970, 99010, 99040, 99050, 99070, 99100, 99120, 99150, 99170, 
    99160, 99170, 99190, 99210, 99220, 99230, 99250, 99270, 99280, 99300, 
    99350, 99390, 99440, 99460, 99480, 99480, 99480, 99480, 99460, 99470, 
    99480, 99500, 99520, 99570, 99610, 99620, 99640, 99650, 99690, 99710, 
    99740, 99750, 99800, 99830, 99870, 99920, 99950, 99970, 99990, 100000, 
    100000, 100000, 99990, 100000, 100000, 100010, 100010, 100020, 100000, 
    99980, 99960, 99950, 99950, 99950, 99970, 100000, 100060, 100090, 100120, 
    100170, 100220, 100290, 100310, 100330, 100340, 100370, 100340, 100320, 
    100320, 100300, 100200, 100190, 100190, 100100, 100060, 100030, 99950, 
    99870, 99810, 99800, 99700, 99740, 99710, 99670, 99760, 99700, 99640, 
    99570, 99620, 99660, 99670, 99660, 99690, 99690, 99650, 99640, 99550, 
    99560, 99550, 99550, 99570, 99690, 99700, 99750, 99750, 99770, 99800, 
    99890, 99910, 99940, 99950, 99960, 99950, 99960, 99990, 100020, 100040, 
    100060, 100100, 100110, 100090, 100060, 100080, 100060, 100060, 100010, 
    100050, 100080, 100110, 100070, 100080, 100140, 100210, 100220, 100260, 
    100260, 100280, 100270, 100250, 100200, 100140, 100130, 100080, 100080, 
    100070, 100080, 100100, 100130, 100110, 100130, 100090, 100110, 100100, 
    100110, 100120, 100120, 100130, 100110, 100100, 100080, 100070, 100030, 
    99980, 99930, 99880, 99840, 99800, 99750, 99690, 99630, 99540, 99440, 
    99350, 99240, 99170, 99110, 99050, 99010, 98970, 98930, 98870, 98820, 
    98780, 98720, 98680, 98650, 98610, 98540, 98530, 98520, 98510, 98510, 
    98500, 98520, 98520, 98510, 98500, 98480, 98490, 98520, 98570, 98600, 
    98640, 98660, 98710, 98700, 98750, 98770, 98750, 98680, 98690, 98670, 
    98690, 98710, 98750, 98720, 98710, 98710, 98680, 98650, 98650, 98610, 
    98600, 98590, 98580, 98600, 98600, 98590, 98630, 98630, 98630, 98650, 
    98660, 98670, 98700, 98690, 98700, 98680, 98690, 98680, 98660, 98620, 
    98610, 98550, 98500, 98490, 98460, 98440, 98450, 98470, 98480, 98480, 
    98490, 98510, 98530, 98510, 98530, 98550, 98550, 98570, 98590, 98610, 
    98650, 98670, 98650, 98660, 98660, 98660, 98650, 98640, 98650, 98660, 
    98670, 98690, 98710, 98720, 98730, 98720, 98720, 98700, 98690, 98690, 
    98690, 98690, 98680, 98690, 98700, 98680, 98710, 98720, 98740, 98760, 
    98760, 98790, 98820, 98860, 98870, 98920, 98970, 99040, 99100, 99150, 
    99230, 99270, 99310, 99350, 99360, 99420, 99470, 99520, 99580, 99680, 
    99770, 99830, 99900, 100010, 100080, 100170, 100260, 100320, 100420, 
    100520, 100600, 100690, 100770, 100860, 100950, 100990, 101060, 101130, 
    101210, 101270, 101340, 101400, 101480, 101530, 101550, 101600, 101610, 
    101610, 101610, 101610, 101600, 101610, 101620, 101620, 101600, 101630, 
    101630, 101630, 101630, 101660, 101700, 101710, 101730, 101750, 101790, 
    101830, 101860, 101840, 101860, 101850, 101840, 101820, 101760, 101750, 
    101690, 101620, 101610, 101550, 101500, 101470, 101430, 101400, 101390, 
    101290, 101210, 101160, 101090, 101010, 100900, 100820, 100770, 100650, 
    100620, 100550, 100440, 100350, 100310, 100300, 100240, 100140, 100080, 
    100040, 99960, 99900, 99820, 99780, 99690, 99730, 99730, 99680, 99600, 
    99570, 99590, 99580, 99600, 99620, 99640, 99640, 99570, 99420, 99480, 
    99540, 99470, 99410, 99390, 99360, 99390, 99400, 99350, 99380, 99390, 
    99420, 99430, 99470, 99500, 99510, 99560, 99610, 99620, 99620, 99650, 
    99710, 99710, 99730, 99760, 99780, 99780, 99830, 99860, 99900, 99930, 
    99960, 100000, 100010, 100030, 100050, 100100, 100120, 100170, 100190, 
    100210, 100250, 100280, 100280, 100320, 100360, 100370, 100390, 100410, 
    100420, 100460, 100460, 100470, 100490, 100520, 100520, 100520, 100510, 
    100490, 100480, 100450, 100420, 100390, 100340, 100300, 100280, 100270, 
    100240, 100200, 100180, 100160, 100110, 100060, 100040, 100010, 99990, 
    99980, 99960, 99960, 99980, 99980, 99960, 99950, 99940, 99920, 99920, 
    99930, 99940, 99940, 99960, 99990, 100020, 100040, 100050, 100080, 
    100100, 100130, 100170, 100190, 100220, 100260, 100330, 100380, 100440, 
    100520, 100560, 100630, 100680, 100730, 100800, 100850, 100880, 100920, 
    100960, 101010, 101060, 101100, 101130, 101140, 101170, 101160, 101150, 
    101140, 101160, 101190, 101190, 101170, 101150, 101140, 101100, 101060, 
    101020, 100990, 100940, 100890, 100850, 100760, 100710, 100670, 100610, 
    100540, 100500, 100410, 100360, 100300, 100290, 100240, 100210, 100180, 
    100140, 100110, 100040, 99950, 99880, 99810, 99770, 99740, 99710, 99670, 
    99620, 99560, 99500, 99430, 99400, 99360, 99360, 99340, 99300, 99300, 
    99330, 99350, 99380, 99420, 99460, 99490, 99520, 99500, 99530, 99540, 
    99560, 99610, 99660, 99700, 99730, 99760, 99810, 99870, 99920, 99970, 
    100010, 100050, 100080, 100150, 100240, 100310, 100370, 100440, 100500, 
    100560, 100610, 100660, 100700, 100760, 100800, 100830, 100880, 100930, 
    100990, 101030, 101070, 101110, 101140, 101150, 101180, 101220, 101260, 
    101260, 101310, 101350, 101410, 101470, 101500, 101540, 101560, 101580, 
    101590, 101610, 101600, 101610, 101650, 101680, 101700, 101740, 101750, 
    101770, 101780, 101780, 101810, 101840, 101860, 101870, 101870, 101880, 
    101950, 101960, 102000, 102040, 102080, 102100, 102140, 102160, 102180, 
    102250, 102250, 102300, 102340, 102360, 102430, 102480, 102500, 102520, 
    102550, 102570, 102620, 102660, 102700, 102730, 102770, 102780, 102810, 
    102840, 102850, 102860, 102870, 102870, 102860, 102840, 102810, 102750, 
    102700, 102640, 102550, 102510, 102490, 102470, 102440, 102400, 102390, 
    102380, 102350, 102350, 102340, 102340, 102310, 102280, 102210, 102100, 
    102020, 101980, 101940, 101910, 101860, 101810, 101780, 101750, 101680, 
    101630, 101590, 101510, 101490, 101440, 101470, 101470, 101480, 101450, 
    101410, 101400, 101410, 101400, 101380, 101350, 101360, 101330, 101300, 
    101280, 101240, 101190, 101160, 101100, 101110, 101060, 101000, 100950, 
    100910, 100860, 100830, 100760, 100670, 100600, 100540, 100440, 100390, 
    100320, 100310, 100330, 100340, 100320, 100340, 100320, 100320, 100310, 
    100310, 100300, 100320, 100340, 100350, 100340, 100390, 100420, 100520, 
    100620, 100710, 100770, 100820, 100960, 101120, 101290, 101480, 101540, 
    101690, 101800, 101840, 101980, 102060, 102090, 102120, 102150, 102180, 
    102180, 102170, 102140, 102090, 102000, 101960, 101870, 101790, 101710, 
    101620, 101570, 101500, 101440, 101370, 101320, 101240, 101180, 101120, 
    101060, 101020, 100970, 100950, 100940, 100910, 100880, 100850, 100850, 
    100840, 100860, 100880, 100890, 101020, 101090, 101120, 101160, 101310, 
    101390, 101420, 101480, 101510, 101550, 101580, 101640, 101680, 101710, 
    101720, 101750, 101800, 101820, 101850, 101880, 101870, 101860, 101830, 
    101790, 101730, 101820, 101870, 101920, 101990, 102040, 102020, 102050, 
    102070, 102120, 102170, 102170, 102160, 102180, 102190, 102200, 102200, 
    102200, 102200, 102190, 102180, 102150, 102130, 102110, 102100, 102100, 
    102090, 102100, 102080, 102070, 102030, 102030, 102020, 101970, 101950, 
    101920, 101890, 101880, 101870, 101870, 101850, 101820, 101820, 101770, 
    101730, 101710, 101680, 101640, 101620, 101610, 101560, 101530, 101500, 
    101470, 101460, 101430, 101380, 101330, 101260, 101230, 101180, 101070, 
    101020, 100970, 100920, 100850, 100840, 100790, 100780, 100730, 100700, 
    100690, 100630, 100620, 100590, 100590, 100620, 100750, 100740, 100760, 
    100780, 100830, 100830, 100860, 100890, 100900, 100930, 100990, 101040, 
    101100, 101150, 101220, 101260, 101290, 101330, 101380, 101430, 101490, 
    101530, 101590, 101650, 101730, 101780, 101860, 101890, 101930, 101960, 
    101990, 102020, 102050, 102130, 102200, 102250, 102300, 102360, 102420, 
    102470, 102530, 102550, 102630, 102690, 102730, 102760, 102810, 102860, 
    102940, 102990, 103020, 103050, 103080, 103090, 103110, 103130, 103150, 
    103180, 103200, 103220, 103250, 103250, 103260, 103290, 103280, 103270, 
    103270, 103270, 103260, 103240, 103250, 103270, 103270, 103240, 103230, 
    103210, 103200, 103170, 103110, 103090, 103040, 102980, 102970, 102930, 
    102910, 102880, 102840, 102790, 102780, 102740, 102690, 102620, 102570, 
    102550, 102510, 102510, 102450, 102420, 102360, 102270, 102200, 102150, 
    102100, 102020, 101970, 101910, 101880, 101830, 101790, 101740, 101670, 
    101600, 101520, 101470, 101420, 101340, 101290, 101210, 101160, 101170, 
    101070, 101050, 101000, 100920, 100880, 100810, 100730, 100700, 100600, 
    100550, 100500, 100450, 100430, 100390, 100340, 100260, 100260, 100280, 
    100260, 100230, 100220, 100240, 100270, 100310, 100350, 100370, 100290, 
    100280, 100330, 100330, 100270, 100200, 100180, 100120, 100170, 100150, 
    100160, 100190, 100170, 100140, 100070, 100050, 100020, 99960, 99910, 
    99890, 99840, 99790, 99680, 99670, 99580, 99530, 99420, 99360, 99170, 
    99180, 99260, 99350, 99380, 99450, 99620, 99800, 99950, 100040, 100150, 
    100310, 100390, 100510, 100610, 100700, 100780, 100820, 100890, 100940, 
    100990, 101010, 101060, 101120, 101170, 101200, 101250, 101300, 101370, 
    101400, 101460, 101500, 101520, 101530, 101530, 101560, 101580, 101570, 
    101580, 101510, 101510, 101510, 101480, 101390, 101330, 101270, 101160, 
    101070, 101010, 100960, 100910, 100860, 100770, 100730, 100680, 100600, 
    100540, 100480, 100420, 100400, 100430, 100380, 100410, 100430, 100480, 
    100500, 100560, 100590, 100600, 100620, 100650, 100660, 100680, 100730, 
    100750, 100790, 100810, 100890, 100920, 100960, 101010, 101050, 101080, 
    101150, 101210, 101300, 101350, 101420, 101510, 101590, 101630, 101610, 
    101670, 101690, 101750, 101760, 101810, 101850, 101870, 101880, 101910, 
    101940, 101970, 101990, 102020, 102020, 102040, 102100, 102150, 102190, 
    102200, 102210, 102250, 102330, 102350, 102470, 102550, 102550, 102540, 
    102640, 102630, 102620, 102510, 102510, 102540, 102440, 102430, 102300, 
    102190, 102040, 101930, 101820, 101680, 101540, 101370, 101210, 101070, 
    101010, 100840, 100760, 100660, 100570, 100540, 100480, 100480, 100430, 
    100410, 100300, 100220, 100090, 100030, 99850, 99700, 99490, 99370, 
    99230, 99060, 98980, 98910, 98940, 99960, 98970, 99080, 99040, 99030, 
    99060, 99050, 99010, 98970, 99240, 99660, 99990, 100250, 100450, 100690, 
    100900, 101080, 101190, 101250, 101320, 101390, 101500, 101530, 101540, 
    101580, 101650, 101690, 101780, 101880, 102000, 102020, 101970, 101950, 
    101920, 101870, 101870, 102000, 101940, 101890, 101870, 101800, 101770, 
    101690, 101630, 101570, 101530, 101480, 101450, 101440, 101400, 101350, 
    101360, 101350, 101360, 101310, 101360, 101420, 101490, 101580, 101620, 
    101700, 101760, 101740, 101760, 101770, 101810, 101810, 101800, 101790, 
    101760, 101740, 101730, 101690, 101660, 101610, 101580, 101550, 101460, 
    101400, 101330, 101260, 101190, 101100, 101000, 100950, 100900, 100800, 
    100730, 100650, 100550, 100510, 100460, 100430, 100390, 100400, 100400, 
    100390, 100430, 100470, 100490, 100530, 100570, 100590, 100590, 100640, 
    100650, 100670, 100680, 100690, 100660, 100740, 100750, 100740, 100740, 
    100770, 100780, 100780, 100770, 100800, 100830, 100830, 100840, 100870, 
    100890, 100920, 100930, 100960, 100980, 100980, 101010, 101000, 101020, 
    101040, 101060, 101100, 101130, 101160, 101160, 101170, 101180, 101200, 
    101200, 101200, 101260, 101290, 101320, 101350, 101380, 101360, 101360, 
    101360, 101370, 101370, 101380, 101390, 101390, 101410, 101420, 101430, 
    101440, 101440, 101450, 101480, 101510, 101530, 101530, 101550, 101590, 
    101630, 101650, 101660, 101680, 101660, 101680, 101670, 101660, 101660, 
    101630, 101630, 101610, 101610, 101620, 101630, 101620, 101600, 101560, 
    101520, 101500, 101480, 101430, 101380, 101360, 101330, 101300, 101270, 
    101230, 101180, 101110, 101050, 100970, 100940, 100830, 100800, 100730, 
    100650, 100620, 100530, 100450, 100420, 100330, 100310, 100290, 100280, 
    100270, 100220, 100240, 100330, 100400, 100440, 100330, 100370, 100380, 
    100540, 100520, 100530, 100550, 100540, 100580, 100630, 100680, 100730, 
    100710, 100710, 100750, 100710, 100700, 100720, 100750, 100740, 100730, 
    100690, 100730, 100760, 100790, 100760, 100730, 100700, 100720, 100670, 
    100660, 100640, 100520, 100530, 100710, 100780, 100770, 100800, 100720, 
    100720, 100630, 100690, 100680, 100730, 100780, 100800, 100930, 101030, 
    101110, 101180, 101270, 101200, 101210, 101250, 101200, 101200, 101180, 
    101260, 101270, 101270, 101250, 101270, 101230, 101210, 101190, 101170, 
    101130, 101140, 101160, 101130, 101150, 101140, 101150, 101140, 101100, 
    101090, 101060, 101030, 100980, 100950, 100870, 100810, 100770, 100720, 
    100650, 100510, 100330, 100290, 100220, 100220, 100130, 100070, 99930, 
    99990, 99950, 99920, 99910, 99900, 99880, 99830, 99780, 99710, 99630, 
    99640, 99670, 99690, 99680, 99710, 99770, 99780, 99800, 99810, 99830, 
    99860, 99850, 99860, 99870, 99900, 99900, 99930, 99940, 99930, 99960, 
    99880, 99860, 99830, 99750, 99770, 99730, 99700, 99700, 99660, 99690, 
    99730, 99740, 99670, 99620, 99680, 99660, 99670, 99670, 99660, 99650, 
    99640, 99660, 99630, 99640, 99590, 99640, 99680, 99700, 99730, 99730, 
    99780, 99790, 99820, 99830, 99810, 99790, 99720, 99680, 99660, 99620, 
    99580, 99580, 99570, 99570, 99570, 99550, 99520, 99470, 99460, 99450, 
    99420, 99400, 99380, 99380, 99330, 99330, 99350, 99400, 99430, 99490, 
    99520, 99540, 99560, 99570, 99570, 99590, 99630, 99680, 99700, 99730, 
    99730, 99730, 99720, 99720, 99710, 99690, 99680, 99660, 99600, 99600, 
    99610, 99560, 99620, 99610, 99550, 99540, 99460, 99370, 99360, 99380, 
    99330, 99280, 99310, 99290, 99300, 99280, 99210, 99190, 99150, 99170, 
    99250, 99160, 99130, 99130, 99160, 99130, 99120, 99150, 99120, 99090, 
    99080, 99070, 99050, 99030, 99020, 99010, 99010, 99020, 99030, 99010, 
    99020, 99030, 99050, 99060, 99050, 99070, 99090, 99110, 99140, 99150, 
    99150, 99140, 99140, 99160, 99190, 99210, 99260, 99300, 99330, 99380, 
    99420, 99450, 99500, 99520, 99550, 99600, 99640, 99670, 99710, 99720, 
    99750, 99780, 99830, 99890, 99920, 99940, 99990, 100040, 100090, 100150, 
    100200, 100260, 100340, 100450, 100510, 100570, 100630, 100650, 100640, 
    100620, 100600, 100570, 100540, 100510, 100450, 100390, 100390, 100360, 
    100420, 100420, 100380, 100380, 100400, 100370, 100310, 100240, 100140, 
    100040, 99930, 99840, 99720, 99550, 99430, 99320, 99240, 99250, 99340, 
    99400, 99500, 99660, 99750, 99810, 99940, 100060, 100130, 100140, 100150, 
    100160, 100200, 100260, 100330, 100390, 100450, 100520, 100530, 100530, 
    100540, 100510, 100470, 100400, 100310, 100180, 100100, 100020, 99940, 
    99850, 99760, 99600, 99450, 99310, 99200, 99060, 98980, 98880, 98850, 
    98840, 98910, 98980, 99050, 99100, 99180, 99220, 99260, 99270, 99290, 
    99290, 99310, 99350, 99330, 99320, 99340, 99370, 99420, 99500, 99590, 
    99680, 99750, 99850, 99920, 100000, 100060, 100110, 100160, 100170, 
    100160, 100140, 100120, 100100, 100070, 100070, 100060, 100040, 100030, 
    100020, 99940, 99850, 99740, 99630, 99590, 99500, 99430, 99360, 99340, 
    99290, 99220, 99200, 99210, 99220, 99220, 99230, 99220, 99240, 99200, 
    99160, 99110, 99090, 99010, 98970, 99100, 99190, 99310, 99380, 99480, 
    99550, 99630, 99680, 99750, 99690, 99810, 99850, 99800, 99810, 99770, 
    99670, 99590, 99560, 99520, 99480, 99490, 99490, 99510, 99550, 99570, 
    99670, 99680, 99820, 99930, 100010, 100170, 100230, 100350, 100520, 
    100670, 100760, 100840, 100990, 101120, 101220, 101330, 101470, 101590, 
    101700, 101800, 101910, 102070, 102090, 102150, 102220, 102250, 102300, 
    102310, 102330, 102350, 102350, 102350, 102380, 102370, 102370, 102370, 
    102400, 102370, 102360, 102260, 102170, 102080, 102040, 101920, 101800, 
    101670, 101590, 101490, 101390, 101300, 101240, 101170, 101120, 101070, 
    101040, 100970, 100950, 100950, 100910, 100890, 100880, 100900, 100890, 
    100880, 100890, 100920, 100850, 100850, 100890, 100880, 100910, 100930, 
    100970, 100960, 101020, 101070, 101100, 101130, 101130, 101150, 101180, 
    101210, 101260, 101310, 101280, 101320, 101320, 101340, 101300, 101300, 
    101270, 101260, 101240, 101220, 101160, 101100, 101060, 101020, 100980, 
    100950, 100920, 100870, 100830, 100800, 100750, 100700, 100670, 100630, 
    100570, 100520, 100480, 100430, 100380, 100320, 100280, 100230, 100200, 
    100160, 100110, 100030, 99970, 99900, 99830, 99810, 99780, 99750, 99730, 
    99670, 99610, 99550, 99440, 99310, 99110, 98930, 98680, 98590, 98390, 
    98170, 98150, 98130, 98050, 97990, 97930, 97870, 97870, 97920, 97960, 
    98010, 98110, 98210, 98400, 98550, 98690, 98870, 99030, 99170, 99220, 
    99320, 99420, 99490, 99580, 99670, 99770, 99860, 99890, 99930, 100000, 
    100020, 100090, 100140, 100140, 100150, 100140, 100110, 100070, 100010, 
    100010, 99980, 100000, 100030, 100040, 100010, 100070, 100020, 100020, 
    100040, 100020, 100020, 100040, 100070, 100070, 100130, 100140, 100140, 
    100160, 100160, 100170, 100200, 100210, 100240, 100260, 100290, 100300, 
    100300, 100320, 100330, 100330, 100320, 100320, 100290, 100280, 100220, 
    100230, 100220, 100210, 100160, 100150, 100140, 100100, 100070, 100040, 
    100010, 100000, 99980, 99970, 99940, 99930, 99870, 99860, 99880, 99860, 
    99830, 99780, 99790, 99790, 99770, 99730, 99750, 99760, 99750, 99780, 
    99790, 99840, 99890, 99920, 99900, 99830, 99860, 99870, 99910, 99930, 
    99960, 99980, 99980, 100000, 100060, 100080, 100110, 100130, 100190, 
    100190, 100190, 100210, 100160, 100140, 100100, 100100, 100070, 100040, 
    100010, 99950, 99940, 99880, 99850, 99800, 99760, 99690, 99610, 99540, 
    99480, 99430, 99360, 99300, 99250, 99210, 99170, 99130, 99090, 99060, 
    99020, 99030, 99030, 99060, 99050, 99070, 99080, 99110, 99130, 99170, 
    99200, 99210, 99190, 99130, 99080, 99050, 99070, 99080, 99120, 99120, 
    99150, 99170, 99230, 99270, 99330, 99490, 99600, 99640, 99650, 99700, 
    99730, 99750, 99850, 99950, 99960, 100000, 100040, 100090, 100090, 
    100090, 100070, 100040, 100040, 100070, 100120, 100180, 100190, 100240, 
    100290, 100300, 100310, 100290, 100260, 100240, 100210, 100210, 100180, 
    100140, 100130, 100110, 100080, 100060, 100020, 100000, 99970, 99950, 
    99930, 99920, 99910, 99920, 99920, 99890, 99860, 99860, 99900, 99920, 
    99950, 99950, 100000, 100060, 100110, 100130, 100160, 100200, 100240, 
    100300, 100350, 100360, 100330, 100350, 100400, 100450, 100510, 100610, 
    100690, 100740, 100770, 100810, 100860, 100910, 100950, 100980, 101040, 
    101100, 101170, 101250, 101310, 101340, 101350, 101330, 101330, 101360, 
    101450, 101450, 101440, 101400, 101390, 101350, 101290, 101220, 101160, 
    101090, 101020, 100920, 100880, 100810, 100770, 100740, 100700, 100650, 
    100640, 100620, 100600, 100600, 100610, 100580, 100580, 100580, 100560, 
    100540, 100520, 100500, 100470, 100440, 100440, 100420, 100420, 100410, 
    100430, 100480, 100520, 100550, 100620, 100640, 100690, 100720, 100800, 
    100840, 100830, 100860, 100850, 100840, 100840, 100890, 100910, 100930, 
    100920, 100900, 100940, 100950, 100960, 100970, 100990, 100990, 100990, 
    100980, 100960, 100990, 100990, 100950, 100960, 100920, 100900, 100930, 
    100870, 100850, 100790, 100770, 100740, 100760, 100770, 100740, 100730, 
    100780, 100750, 100800, 100810, 100850, 100790, 100820, 100840, 100860, 
    100850, 100840, 100850, 100840, 100790, 100790, 100790, 100700, 100740, 
    100770, 100760, 100750, 100760, 100750, 100710, 100710, 100660, 100690, 
    100690, 100630, 100710, 100730, 100710, 100740, 100760, 100800, 100830, 
    100890, 100900, 100940, 101100, 101180, 101330, 101340, 101240, 101210, 
    101250, 101480, 101560, 101610, 101670, 101670, 101670, 101670, 101680, 
    101710, 101730, 101740, 101750, 101740, 101740, 101730, 101720, 101710, 
    101700, 101660, 101620, 101580, 101500, 101440, 101400, 101350, 101280, 
    101190, 101100, 101020, 100920, 100850, 100810, 100770, 100730, 100690, 
    100650, 100590, 100520, 100490, 100430, 100430, 100370, 100330, 100280, 
    100250, 100180, 100110, 100080, 100060, 100090, 100010, 99920, 99870, 
    100030, 100010, 99930, 99970, 99980, 99960, 99860, 99710, 99700, 99650, 
    99560, 99340, 99420, 99600, 99750, 100090, 100220, 100300, 100350, 
    100290, 100280, 100250, 100240, 100180, 100250, 100220, 100210, 100170, 
    100260, 100300, 100210, 100180, 100410, 100510, 100520, 100480, 100510, 
    100430, 100410, 100370, 100360, 100380, 100490, 100460, 100400, 100410, 
    100420, 100400, 100350, 100320, 100300, 100260, 100220, 100180, 100160, 
    100100, 100010, 99950, 99900, 99850, 99790, 99690, 99700, 99680, 99670, 
    99680, 99650, 99580, 99580, 99540, 99380, 99330, 99400, 99460, 99440, 
    99470, 99530, 99570, 99560, 99550, 99540, 99540, 99560, 99530, 99540, 
    99540, 99550, 99570, 99580, 99610, 99610, 99620, 99630, 99680, 99720, 
    99750, 99780, 99780, 99830, 99860, 99900, 99920, 99940, 99980, 100000, 
    100050, 100080, 100100, 100120, 100140, 100110, 100160, 100210, 100180, 
    100210, 100220, 100250, 100250, 100260, 100260, 100230, 100210, 100200, 
    100210, 100240, 100270, 100260, 100270, 100250, 100260, 100270, 100300, 
    100290, 100280, 100270, 100270, 100270, 100290, 100290, 100290, 100310, 
    100260, 100270, 100300, 100310, 100310, 100230, 100180, 100170, 100240, 
    100260, 100360, 100350, 100350, 100320, 100240, 100410, 100430, 100380, 
    100400, 100450, 100470, 100480, 100470, 100460, 100440, 100440, 100450, 
    100450, 100450, 100450, 100450, 100480, 100510, 100490, 100470, 100470, 
    100470, 100470, 100520, 100480, 100480, 100490, 100470, 100450, 100440, 
    100420, 100430, 100400, 100390, 100370, 100360, 100350, 100300, 100270, 
    100270, 100260, 100260, 100250, 100290, 100240, 100220, 100030, 100140, 
    100130, 100110, 100120, 100050, 100070, 100100, 100080, 100030, 100090, 
    100050, 100060, 100080, 100080, 100090, 100080, 100120, 100150, 100190, 
    100190, 100210, 100230, 100250, 100280, 100300, 100360, 100390, 100400, 
    100470, 100450, 100520, 100550, 100640, 100670, 100730, 100750, 100740, 
    100790, 100830, 100830, 100890, 100940, 100990, 101010, 101050, 101080, 
    101100, 101140, 101180, 101210, 101210, 101250, 101290, 101330, 101360, 
    101390, 101430, 101470, 101510, 101510, 101540, 101560, 101630, 101670, 
    101730, 101760, 101760, 101780, 101760, 101780, 101810, 101830, 101880, 
    101910, 101910, 101930, 101940, 101930, 102020, 102050, 102090, 102110, 
    102100, 102140, 102150, 102170, 102210, 102230, 102260, 102320, 102370, 
    102370, 102410, 102460, 102480, 102490, 102520, 102540, 102570, 102590, 
    102620, 102650, 102680, 102710, 102700, 102710, 102690, 102710, 102720, 
    102730, 102740, 102750, 102760, 102780, 102760, 102750, 102730, 102710, 
    102680, 102690, 102670, 102650, 102640, 102640, 102600, 102580, 102560, 
    102550, 102530, 102530, 102510, 102490, 102480, 102470, 102450, 102460, 
    102470, 102470, 102440, 102440, 102430, 102430, 102420, 102420, 102410, 
    102390, 102390, 102400, 102410, 102410, 102410, 102390, 102350, 102300, 
    102320, 102300, 102250, 102280, 102240, 102230, 102240, 102230, 102220, 
    102200, 102180, 102150, 102130, 102130, 102130, 102130, 102140, 102120, 
    102130, 102140, 102170, 102140, 102170, 102190, 102210, 102190, 102180, 
    102140, 102160, 102140, 102070, 102050, 102070, 102050, 102010, 101980, 
    101940, 101920, 101890, 101910, 101880, 101850, 101810, 101790, 101760, 
    101730, 101700, 101670, 101650, 101600, 101570, 101540, 101490, 101460, 
    101450, 101490, 101480, 101480, 101480, 101480, 101510, 101500, 101500, 
    101500, 101520, 101540, 101560, 101610, 101640, 101660, 101680, 101680, 
    101700, 101710, 101730, 101730, 101720, 101730, 101750, 101770, 101800, 
    101790, 101810, 101810, 101830, 101870, 101910, 101930, 101960, 101980, 
    102030, 102050, 102070, 102100, 102110, 102090, 102090, 102120, 102120, 
    102130, 102180, 102150, 102180, 102220, 102240, 102230, 102330, 102220, 
    102200, 102190, 102160, 102130, 102090, 102070, 102030, 102040, 102000, 
    101970, 101950, 101930, 101940, 101910, 101910, 101880, 101880, 101880, 
    101890, 101900, 101900, 101910, 101930, 101890, 101850, 101830, 101830, 
    101810, 101790, 101770, 101770, 101760, 101760, 101780, 101730, 101720, 
    101710, 101710, 101720, 101740, 101760, 101810, 101880, 101960, 102040, 
    102100, 102170, 102230, 102270, 102330, 102380, 102420, 102490, 102550, 
    102590, 102650, 102690, 102740, 102760, 102780, 102800, 102830, 102850, 
    102880, 102900, 102950, 102970, 103010, 103050, 103090, 103110, 103110, 
    103120, 103140, 103150, 103150, 103200, 103220, 103230, 103250, 103280, 
    103290, 103280, 103280, 103280, 103290, 103300, 103300, 103290, 103320, 
    103340, 103360, 103370, 103390, 103380, 103360, 103360, 103340, 103330, 
    103300, 103280, 103270, 103250, 103210, 103180, 103150, 103120, 103060, 
    102990, 102960, 102930, 102900, 102830, 102830, 102840, 102850, 102840, 
    102840, 102820, 102800, 102790, 102780, 102750, 102760, 102750, 102750, 
    102740, 102780, 102750, 102740, 102730, 102710, 102690, 102640, 102600, 
    102580, 102530, 102520, 102460, 102510, 102490, 102500, 102520, 102480, 
    102470, 102420, 102400, 102370, 102360, 102320, 102310, 102320, 102310, 
    102290, 102270, 102270, 102250, 102270, 102260, 102260, 102270, 102270, 
    102300, 102320, 102350, 102370, 102380, 102390, 102390, 102410, 102430, 
    102410, 102410, 102440, 102440, 102430, 102420, 102420, 102400, 102390, 
    102380, 102360, 102330, 102310, 102290, 102280, 102280, 102270, 102230, 
    102200, 102140, 102100, 102050, 102020, 101990, 101950, 101900, 101860, 
    101870, 101820, 101780, 101730, 101690, 101640, 101600, 101570, 101550, 
    101520, 101490, 101460, 101440, 101430, 101400, 101370, 101390, 101350, 
    101310, 101290, 101250, 101240, 101210, 101190, 101180, 101140, 101120, 
    101080, 101000, 100990, 100970, 100950, 100940, 100920, 100900, 100910, 
    100910, 100910, 100910, 100850, 100820, 100830, 100780, 100730, 100700, 
    100690, 100760, 100780, 100730, 100720, 100670, 100600, 100620, 100590, 
    100540, 100500, 100420, 100340, 100320, 100280, 100250, 100280, 100270, 
    100230, 100230, 100200, 100220, 100210, 100260, 100250, 100220, 100190, 
    100160, 100150, 100180, 100200, 100240, 100210, 100130, 100120, 100080, 
    100050, 100030, 99980, 99920, 99920, 99960, 99960, 100000, 100040, 
    100070, 100030, 100060, 100100, 100130, 100140, 100130, 100140, 100080, 
    100040, 100020, 100070, 100120, 100170, 100210, 100230, 100280, 100330, 
    100380, 100420, 100460, 100480, 100510, 100530, 100550, 100560, 100590, 
    100610, 100630, 100630, 100660, 100690, 100690, 100700, 100710, 100720, 
    100740, 100750, 100740, 100750, 100720, 100690, 100690, 100650, 100630, 
    100590, 100570, 100580, 100580, 100580, 100570, 100560, 100530, 100530, 
    100500, 100470, 100430, 100410, 100370, 100340, 100340, 100290, 100250, 
    100220, 100190, 100190, 100220, 100210, 100180, 100150, 100120, 100110, 
    100080, 100080, 100050, 100000, 99970, 99940, 99920, 99900, 99880, 99890, 
    99870, 99830, 99820, 99790, 99780, 99750, 99730, 99710, 99720, 99700, 
    99690, 99660, 99620, 99570, 99540, 99550, 99530, 99540, 99510, 99510, 
    99530, 99540, 99570, 99600, 99630, 99670, 99750, 99740, 99780, 99810, 
    99870, 99890, 99930, 100000, 100020, 100060, 100080, 100100, 100150, 
    100110, 100090, 100040, 100020, 100020, 100030, 100170, 100260, 100340, 
    100350, 100340, 100390, 100420, 100380, 100380, 100370, 100340, 100360, 
    100400, 100400, 100410, 100410, 100410, 100400, 100380, 100350, 100350, 
    100330, 100340, 100390, 100440, 100470, 100460, 100500, 100530, 100540, 
    100550, 100540, 100560, 100580, 100610, 100640, 100710, 100750, 100790, 
    100830, 100890, 100890, 100850, 100900, 100930, 100960, 100970, 100980, 
    100990, 101010, 101050, 100960, 100930, 100920, 100970, 100930, 100880, 
    100940, 100980, 100950, 100990, 100960, 100940, 100890, 100860, 100830, 
    100820, 100770, 100790, 100740, 100670, 100620, 100550, 100430, 100440, 
    100430, 100400, 100310, 100240, 100200, 100160, 100090, 100040, 100000, 
    99980, 99950, 99920, 99900, 99880, 99840, 99780, 99730, 99660, 99660, 
    99610, 99570, 99560, 99550, 99570, 99580, 99610, 99630, 99630, 99690, 
    99720, 99730, 99780, 99820, 99910, 99960, 99990, 100010, 100020, 100030, 
    100100, 100110, 100130, 100140, 100160, 100160, 100190, 100210, 100250, 
    100290, 100300, 100320, 100360, 100390, 100420, 100510, 100520, 100530, 
    100590, 100650, 100680, 100630, 100680, 100650, 100610, 100530, 100410, 
    100260, 100140, 99970, 99870, 99980, 99640, 99520, 99400, 99310, 99170, 
    99120, 99050, 99010, 99010, 98980, 98930, 98890, 98810, 98680, 98560, 
    98490, 98390, 98310, 98190, 98180, 98170, 98140, 98170, 98190, 98210, 
    98220, 98280, 98330, 98380, 98470, 98530, 98650, 98710, 98840, 98940, 
    99040, 99120, 99250, 99320, 99410, 99470, 99620, 99630, 99700, 99730, 
    99800, 99790, 99850, 99840, 99860, 99870, 99790, 99790, 99790, 99740, 
    99670, 99630, 99630, 99640, 99650, 99660, 99650, 99650, 99720, 99800, 
    99820, 99960, 100100, 100240, 100320, 100380, 100450, 100530, 100640, 
    100720, 100850, 100940, 100990, 100970, 101010, 101020, 101050, 101050, 
    101100, 101100, 101090, 101120, 101120, 101090, 101080, 101040, 100980, 
    100980, 100970, 100940, 100980, 100980, 100930, 100930, 100940, 100870, 
    100890, 100910, 100900, 100890, 100950, 100970, 100990, 101000, 100930, 
    100980, 100980, 100990, 101000, 100900, 100850, 100780, 100810, 100800, 
    100770, 100780, 100780, 100770, 100750, 100690, 100680, 100720, 100710, 
    100700, 100610, 100560, 100690, 100690, 100650, 100630, 100620, 100650, 
    100640, 100580, 100380, 100320, 100440, 100470, 100500, 100420, 100390, 
    100350, 100370, 100370, 100320, 100320, 100370, 100410, 100540, 100640, 
    100650, 100690, 100740, 100800, 100830, 100850, 100950, 100920, 100950, 
    100940, 100980, 101000, 101070, 101040, 101040, 101020, 101020, 101040, 
    101030, 100950, 100930, 100870, 100730, 100670, 100630, 100590, 100510, 
    100490, 100460, 100390, 100320, 100260, 100160, 100050, 100040, 99960, 
    99990, 99880, 99770, 99750, 99700, 99690, 99650, 99590, 99540, 99550 ;

 surface_air_pressure_2m = 98800, 99210, 99810, 100780, 101360, 101710, 
    102140, 102070, 102000, 101710, 101930, 102020, 101890, 101810, 101630, 
    101700, 101920, 102150, 101880, 101070, 99950, 99110, 99320, 99940, 
    100090, 100150, 99700, 99210, 98800, 99060, 99410, 99690, 100290, 100470, 
    100280, 100070, 100470, 102220, 102540, 102510, 102280, 101520, 100000, 
    99370, 98200, 98050, 98690, 100170, 100620, 100620, 100390, 100090, 
    100220, 101070, 101630, 99370, 99220, 100730, 100210, 99580, 103280, 
    103340, 103100, 102760, 102210, 101450, 100590, 100630, 100830, 100810, 
    100590, 100510, 100650, 100700, 100990, 101250, 101540, 101690, 101390, 
    100510, 99580, 100760, 101450, 101520, 101610, 101770, 101630, 101520, 
    101190, 101090, 101180, 101500, 101810, 102060, 102190, 102260, 102180, 
    102220, 102280, 102260, 102250, 102070, 101910, 101620, 101470, 101300, 
    101110, 101130, 101330, 101880, 101880, 101560, 100840, 101100, 100390, 
    100100, 99760, 99850, 100440, 100910, 104640, 101260, 101350, 101550, 
    101620, 101510, 101500, 101260, 100830, 100670, 100330, 100260, 100320, 
    100170, 100090, 100720, 100960, 101610, 101730, 101040, 100440, 99510, 
    98870, 97380, 98310, 99250, 99700, 99640, 99600, 99600, 100110, 100200, 
    100280, 100280, 100230, 100260, 100310, 100480, 100580, 100830, 100840, 
    100900, 100890, 100780, 100760, 100780, 100740, 100610, 100580, 100740, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 102770, 102740, 102730, 102720, 102700, 102690, 102670, 
    102670, 102700, 102690, 102680, 102640, 102660, 102640, 102610, 102600, 
    102590, 102570, 102480, 102540, 102510, 102510, 102530, 102510, 102480, 
    102450, 102450, 102460, 102390, 102380, 102340, 102350, 102350, 102330, 
    102310, 102270, 102240, 102250, 102230, 102220, 102200, 102210, 102210, 
    102190, 102210, 102200, 102200, 102220, 102210, 102180, 102150, 102130, 
    102110, 102060, 102040, 102050, 101990, 102040, 102000, 101980, 102020, 
    102010, 101990, 101960, 101940, 101950, 101930, 101950, 101950, 101950, 
    101930, 101910, 101920, 101870, 101880, 101830, 101850, 101860, 101830, 
    101850, 101840, 101820, 101820, 101820, 101830, 101820, 101810, 101820, 
    101810, 101830, 101810, 101820, 101810, 101810, 101800, 101830, 101820, 
    101810, 101840, 101790, 101800, 101820, 101820, 101820, 101810, 101820, 
    101840, 101840, 101850, 101870, 101890, 101910, 101910, 101940, 101960, 
    101980, 102020, 102050, 102080, 102090, 102110, 102130, 102130, 102140, 
    102160, 102170, 102180, 102200, 102220, 102220, 102220, 102240, 102230, 
    102230, 102220, 102220, 102150, 102220, 102210, 102170, 102160, 102140, 
    102190, 102170, 102200, 102190, 102180, 102160, 102150, 102150, 102140, 
    102140, 102170, 102210, 102210, 102220, 102240, 102240, 102240, 102230, 
    102220, 102190, 102200, 102220, 102230, 102230, 102250, 102260, 102270, 
    102260, 102270, 102250, 102230, 102220, 102210, 102210, 102210, 102200, 
    102180, 102180, 102150, 102160, 102160, 102150, 102120, 102100, 102100, 
    102120, 102110, 102140, 102150, 102170, 102160, 102140, 102100, 102060, 
    102050, 102050, 102020, 102010, 102000, 101990, 101980, 101970, 101970, 
    101950, 101920, 101890, 101870, 101870, 101850, 101820, 101800, 101790, 
    101790, 101760, 101750, 101720, 101710, 101670, 101640, 101610, 101570, 
    101560, 101560, 101530, 101520, 101500, 101470, 101470, 101440, 101410, 
    101380, 101370, 101370, 101360, 101380, 101370, 101380, 101370, 101370, 
    101360, 101350, 101340, 101340, 101340, 101320, 101330, 101330, 101310, 
    101330, 101300, 101300, 101280, 101290, 101270, 101250, 101220, 101210, 
    101220, 101220, 101220, 101220, 101210, 101210, 101190, 101210, 101180, 
    101160, 101160, 101150, 101140, 101130, 101140, 101110, 101100, 101100, 
    101100, 101080, 101090, 101080, 101080, 101100, 101130, 101150, 101160, 
    101170, 101200, 101220, 101230, 101240, 101260, 101270, 101280, 101290, 
    101290, 101290, 101310, 101330, 101340, 101340, 101350, 101370, 101370, 
    101370, 101390, 101400, 101400, 101410, 101430, 101410, 101430, 101430, 
    101420, 101410, 101380, 101350, 101320, 101300, 101300, 101290, 101260, 
    101250, 101240, 101220, 101210, 101170, 101140, 101100, 101070, 101030, 
    101020, 100990, 100970, 100920, 100900, 100850, 100810, 100760, 100740, 
    100710, 100680, 100630, 100590, 100560, 100530, 100500, 100490, 100460, 
    100440, 100370, 100370, 100380, 100390, 100400, 100420, 100430, 100460, 
    100520, 100570, 100620, 100640, 100700, 100750, 100800, 100840, 100860, 
    100890, 100940, 100990, 101040, 101070, 101120, 101170, 101200, 101200, 
    101230, 101230, 101230, 101240, 101230, 101230, 101230, 101210, 101210, 
    101240, 101270, 101300, 101310, 101370, 101420, 101440, 101480, 101530, 
    101580, 101620, 101650, 101650, 101660, 101650, 101650, 101620, 101620, 
    101620, 101570, 101550, 101520, 101470, 101400, 101350, 101330, 101260, 
    101240, 101220, 101150, 101090, 101070, 101040, 101000, 100980, 100930, 
    100880, 100830, 100810, 100770, 100710, 100680, 100610, 100580, 100470, 
    100430, 100350, 100300, 100280, 100220, 100150, 100120, 100110, 100120, 
    100120, 100110, 100140, 100130, 100140, 100150, 100130, 100110, 100130, 
    100130, 100140, 100170, 100180, 100240, 100250, 100280, 100290, 100300, 
    100370, 100430, 100460, 100490, 100520, 100520, 100510, 100540, 100580, 
    100610, 100700, 100680, 100680, 100670, 100660, 100640, 100640, 100580, 
    100640, 100620, 100590, 100470, 100490, 100200, 100170, 100120, 100040, 
    99990, 99830, 99740, 99730, 99620, 99610, 99620, 99650, 99670, 99640, 
    99670, 99660, 99640, 99650, 99720, 99720, 99760, 99790, 99830, 99920, 
    99940, 99980, 99960, 99980, 100010, 100010, 100060, 100090, 100120, 
    100140, 100140, 100160, 100230, 100280, 100320, 100370, 100410, 100470, 
    100540, 100610, 100700, 100710, 100760, 100810, 100840, 100890, 100920, 
    100950, 101020, 101050, 101060, 101080, 101090, 101130, 101170, 101180, 
    101160, 101150, 101140, 101120, 101080, 101050, 100980, 100920, 100940, 
    100930, 100890, 100860, 100790, 100700, 100590, 100480, 100500, 100460, 
    100440, 100400, 100390, 100380, 100360, 100310, 100290, 100270, 100270, 
    100230, 100220, 100220, 100220, 100250, 100280, 100280, 100320, 100330, 
    100380, 100410, 100420, 100440, 100470, 100460, 100490, 100490, 100490, 
    100490, 100470, 100460, 100440, 100420, 100400, 100390, 100360, 100330, 
    100330, 100290, 100280, 100260, 100230, 100220, 100170, 100170, 100190, 
    100190, 100210, 100260, 100340, 100360, 100450, 100500, 100550, 100590, 
    100660, 100700, 100740, 100820, 100830, 100840, 100880, 100900, 100890, 
    100900, 100940, 100920, 100920, 100920, 100910, 100890, 100880, 100830, 
    100820, 100760, 100690, 100610, 100540, 100420, 100440, 100430, 100360, 
    100230, 100250, 99980, 99890, 99940, 100020, 99900, 99910, 99910, 99910, 
    99880, 99880, 99900, 99910, 99930, 99950, 99960, 99990, 100030, 100050, 
    100050, 100050, 100030, 100020, 100020, 100050, 100040, 100040, 100020, 
    100010, 100000, 100040, 100030, 100020, 100030, 100030, 100010, 99970, 
    99970, 99970, 99970, 99980, 99980, 99950, 99940, 99920, 99890, 99880, 
    99880, 99880, 99870, 99840, 99830, 99850, 99850, 99840, 99850, 99860, 
    99840, 99820, 99830, 99820, 99800, 99770, 99750, 99740, 99730, 99740, 
    99730, 99710, 99700, 99660, 99640, 99650, 99650, 99650, 99660, 99670, 
    99690, 99700, 99720, 99740, 99780, 99810, 99840, 99890, 99960, 99950, 
    100020, 100060, 100120, 100170, 100200, 100240, 100260, 100280, 100330, 
    100370, 100360, 100390, 100410, 100450, 100500, 100520, 100590, 100620, 
    100620, 100620, 100610, 100610, 100580, 100570, 100540, 100490, 100450, 
    100440, 100430, 100360, 100370, 100380, 100360, 100410, 100440, 100480, 
    100510, 100530, 100570, 100660, 100730, 100780, 100800, 100940, 101030, 
    101120, 101200, 101290, 101360, 101400, 101470, 101530, 101550, 101610, 
    101640, 101690, 101770, 101790, 101840, 101860, 101880, 101920, 101930, 
    101970, 101980, 102010, 102020, 102030, 102030, 102020, 102040, 102060, 
    102070, 102040, 102030, 102010, 102040, 101940, 101970, 101920, 101910, 
    101960, 102000, 101990, 102020, 102040, 102020, 102000, 102030, 102010, 
    102000, 102000, 102020, 102020, 102050, 102040, 102040, 102040, 102040, 
    102040, 102010, 102010, 101970, 101980, 101970, 101970, 101970, 101990, 
    101990, 101970, 101960, 101950, 101940, 101930, 101890, 101880, 101870, 
    101850, 101810, 101780, 101770, 101750, 101720, 101690, 101650, 101610, 
    101560, 101500, 101450, 101430, 101410, 101420, 101430, 101470, 101510, 
    101510, 101490, 101450, 101430, 101410, 101400, 101400, 101400, 101410, 
    101420, 101410, 101410, 101410, 101390, 101420, 101450, 101490, 101510, 
    101530, 101550, 101570, 101600, 101620, 101630, 101640, 101650, 101640, 
    101650, 101630, 101650, 101640, 101620, 101610, 101600, 101610, 101570, 
    101560, 101540, 101500, 101450, 101430, 101400, 101390, 101340, 101290, 
    101260, 101240, 101220, 101240, 101210, 101190, 101150, 101120, 101090, 
    101070, 101030, 100980, 100910, 100890, 100840, 100800, 100770, 100710, 
    100660, 100620, 100580, 100640, 100610, 100620, 100610, 100620, 100630, 
    100630, 100650, 100640, 100650, 100640, 100630, 100630, 100600, 100590, 
    100560, 100580, 100540, 100530, 100480, 100460, 100440, 100370, 100340, 
    100320, 100320, 100350, 100370, 100390, 100410, 100430, 100460, 100470, 
    100470, 100470, 100480, 100490, 100470, 100460, 100440, 100410, 100400, 
    100390, 100370, 100360, 100300, 100270, 100270, 100240, 100210, 100180, 
    100160, 100130, 100140, 100140, 100130, 100090, 100060, 100050, 100010, 
    100000, 100000, 100000, 99980, 99930, 100000, 99980, 99910, 99920, 99920, 
    99900, 99900, 99920, 99900, 99880, 99890, 99890, 99910, 99900, 99880, 
    99880, 99880, 99850, 99820, 99830, 99820, 99840, 99830, 99840, 99870, 
    99920, 99980, 99990, 100030, 100050, 100090, 100130, 100190, 100270, 
    100380, 100460, 100520, 100580, 100650, 100740, 100830, 100890, 100980, 
    101070, 101140, 101180, 101250, 101330, 101350, 101360, 101350, 101350, 
    101360, 101350, 101330, 101310, 101290, 101290, 101300, 101260, 101250, 
    101200, 101140, 101120, 101050, 100940, 100850, 100760, 100620, 100470, 
    100390, 100270, 100150, 100020, 99860, 99730, 99610, 99460, 99340, 99270, 
    99130, 99110, 99080, 99080, 99130, 99120, 99150, 99190, 99250, 99320, 
    99420, 99450, 99490, 99560, 99580, 99670, 99740, 99780, 99840, 99890, 
    99970, 100020, 100050, 100120, 100140, 100180, 100220, 100260, 100310, 
    100330, 100390, 100440, 100450, 100500, 100560, 100580, 100590, 100610, 
    100600, 100630, 100640, 100650, 100650, 100640, 100640, 100630, 100630, 
    100620, 100580, 100570, 100570, 100570, 100590, 100590, 100580, 100570, 
    100570, 100610, 100630, 100590, 100590, 100600, 100580, 100570, 100570, 
    100570, 100560, 100570, 100550, 100540, 100520, 100520, 100520, 100500, 
    100510, 100510, 100510, 100510, 100520, 100520, 100490, 100460, 100440, 
    100420, 100400, 100370, 100340, 100320, 100300, 100270, 100240, 100210, 
    100180, 100140, 100090, 100080, 100080, 100070, 100060, 100060, 100080, 
    100100, 100120, 100140, 100130, 100120, 100140, 100140, 100140, 100140, 
    100110, 100110, 100100, 100100, 100090, 100070, 100060, 100040, 100010, 
    99980, 99960, 99940, 99920, 99890, 99870, 99870, 99840, 99810, 99790, 
    99780, 99780, 99770, 99760, 99770, 99760, 99780, 99760, 99760, 99740, 
    99730, 99720, 99690, 99710, 99690, 99640, 99710, 99680, 99700, 99730, 
    99750, 99750, 99730, 99700, 99710, 99710, 99710, 99710, 99710, 99730, 
    99760, 99780, 99780, 99780, 99800, 99820, 99820, 99800, 99810, 99820, 
    99850, 99870, 99900, 99920, 99960, 99990, 100020, 100040, 100020, 100020, 
    100060, 100080, 100070, 100100, 100150, 100130, 100140, 100140, 100140, 
    100140, 100140, 100140, 100100, 100040, 100070, 100090, 100140, 100190, 
    100180, 100190, 100170, 100170, 100180, 100170, 100180, 100150, 100120, 
    100070, 100090, 100110, 100100, 100070, 100070, 100030, 100020, 100000, 
    99980, 99980, 99960, 99960, 99950, 99940, 99950, 99910, 99900, 99890, 
    99880, 99870, 99880, 99880, 99850, 99850, 99860, 99880, 99890, 99880, 
    99880, 99890, 99900, 99900, 99900, 99920, 99950, 99980, 100020, 100050, 
    100120, 100150, 100180, 100200, 100230, 100290, 100330, 100370, 100410, 
    100410, 100440, 100480, 100510, 100560, 100590, 100610, 100650, 100680, 
    100700, 100700, 100730, 100750, 100810, 100920, 101030, 101080, 101120, 
    101170, 101220, 101250, 101330, 101370, 101420, 101480, 101540, 101590, 
    101660, 101710, 101730, 101730, 101760, 101800, 101830, 101820, 101880, 
    101890, 101860, 101850, 101880, 101830, 101780, 101720, 101640, 101540, 
    101400, 101250, 101110, 100920, 100710, 100570, 100330, 100060, 99810, 
    99600, 99400, 99140, 98940, 98720, 98440, 98350, 98440, 98500, 98500, 
    98480, 98460, 98430, 98430, 98420, 98410, 98350, 98330, 98350, 98350, 
    98360, 98370, 98380, 98410, 98450, 98520, 98610, 98650, 98660, 98740, 
    98830, 98940, 99030, 99110, 99170, 99230, 99290, 99310, 99340, 99350, 
    99340, 99330, 99470, 99530, 99580, 99600, 99600, 99630, 99630, 99610, 
    99610, 99660, 99690, 99770, 99830, 99830, 99810, 99840, 99910, 99950, 
    100010, 99990, 99990, 99960, 100040, 100180, 100180, 100230, 100190, 
    100140, 100200, 100200, 100120, 100100, 100130, 100130, 100180, 100190, 
    100160, 100170, 100140, 100150, 100140, 100150, 100190, 100180, 100190, 
    100280, 100300, 100310, 100340, 100450, 100480, 100570, 100590, 100650, 
    100680, 100700, 100720, 100730, 100720, 100740, 100800, 100840, 100820, 
    100780, 100800, 100810, 100820, 100810, 100800, 100780, 100790, 100750, 
    100710, 100690, 100650, 100630, 100570, 100480, 100430, 100400, 100360, 
    100330, 100300, 100270, 100250, 100270, 100250, 100240, 100230, 100220, 
    100200, 100160, 100160, 100150, 100120, 100190, 100220, 100200, 100220, 
    100250, 100310, 100370, 100430, 100500, 100550, 100610, 100640, 100690, 
    100740, 100810, 100830, 100880, 100930, 100950, 101010, 101040, 101080, 
    101090, 101140, 101170, 101180, 101200, 101240, 101260, 101280, 101300, 
    101350, 101380, 101430, 101470, 101510, 101520, 101580, 101630, 101670, 
    101720, 101750, 101800, 101820, 101860, 101880, 101910, 101940, 101970, 
    102010, 102040, 102060, 102100, 102120, 102130, 102130, 102150, 102170, 
    102190, 102180, 102190, 102220, 102240, 102240, 102260, 102240, 102220, 
    102210, 102200, 102160, 102110, 102050, 102020, 101930, 101890, 101830, 
    101750, 101650, 101530, 101440, 101270, 101150, 101020, 100890, 100730, 
    100540, 100370, 100140, 99960, 99810, 99650, 99580, 99510, 99410, 99320, 
    99260, 99200, 99180, 99140, 99130, 99140, 99140, 99150, 99170, 99190, 
    99270, 99330, 99400, 99480, 99520, 99590, 99700, 99780, 99910, 100020, 
    100150, 100310, 100430, 100600, 100670, 100800, 100940, 101010, 101110, 
    101180, 101250, 101300, 101370, 101450, 101470, 101550, 101630, 101670, 
    101760, 101820, 101890, 101990, 102060, 102120, 102150, 102210, 102260, 
    102290, 102290, 102310, 102310, 102290, 102270, 102290, 102270, 102250, 
    102210, 102180, 102180, 102130, 102100, 102090, 102100, 102110, 102120, 
    102120, 102100, 102120, 102130, 102100, 102120, 102110, 102050, 102000, 
    101970, 101940, 101900, 101840, 101740, 101670, 101620, 101530, 101490, 
    101390, 101260, 101210, 101160, 101120, 101060, 101010, 100940, 100840, 
    100730, 100680, 100580, 100450, 100330, 100180, 100090, 99980, 99940, 
    99880, 99800, 99740, 99680, 99620, 99560, 99540, 99520, 99490, 99500, 
    99560, 99630, 99670, 99700, 99700, 99730, 99770, 99720, 99690, 99650, 
    99580, 99580, 99690, 99660, 99660, 99650, 99600, 99590, 99550, 99530, 
    99510, 99440, 99400, 99400, 99330, 99300, 99260, 99180, 99150, 99060, 
    98990, 99020, 99040, 99020, 98990, 98980, 99020, 99030, 99120, 99150, 
    99180, 99300, 99320, 99470, 99520, 99630, 99700, 99740, 99800, 99900, 
    99950, 99970, 99950, 100040, 100040, 100110, 100170, 100190, 100220, 
    100310, 100370, 100410, 100420, 100460, 100420, 100440, 100420, 100360, 
    100330, 100200, 100200, 100220, 100190, 100190, 100180, 100160, 100170, 
    100080, 100080, 100080, 100100, 100150, 100210, 100240, 100260, 100280, 
    100350, 100400, 100430, 100470, 100530, 100570, 100620, 100650, 100710, 
    100790, 100850, 100910, 100940, 100980, 101020, 101100, 101140, 101190, 
    101220, 101270, 101300, 101380, 101420, 101490, 101520, 101590, 101620, 
    101650, 101700, 101740, 101770, 101800, 101840, 101880, 101920, 101960, 
    102000, 102040, 102080, 102110, 102120, 102140, 102160, 102200, 102240, 
    102260, 102280, 102320, 102330, 102380, 102380, 102390, 102380, 102370, 
    102360, 102350, 102300, 102300, 102270, 102250, 102240, 102190, 102160, 
    102140, 102080, 102080, 102030, 101950, 101830, 101750, 101670, 101590, 
    101540, 101470, 101360, 101230, 101110, 101040, 100970, 100900, 100800, 
    100710, 100600, 100530, 100490, 100430, 100340, 100250, 100200, 100150, 
    100120, 100070, 100040, 100000, 99970, 99900, 99870, 99780, 99750, 99660, 
    99570, 99490, 99460, 99380, 99240, 99190, 99110, 98980, 98920, 98860, 
    98770, 98730, 98740, 98800, 98880, 98940, 99000, 99060, 99050, 99100, 
    99130, 99160, 99150, 99060, 98960, 98890, 98760, 98680, 98590, 98490, 
    98390, 98300, 98200, 98070, 97980, 97850, 97750, 97670, 97620, 97590, 
    97600, 97620, 97640, 97690, 97760, 97780, 97910, 98000, 98080, 98180, 
    98290, 98400, 98530, 98680, 98790, 98890, 99090, 99300, 99510, 99650, 
    99790, 99910, 99960, 99920, 99990, 100040, 100140, 100170, 100250, 
    100300, 100310, 100320, 100360, 100360, 100350, 100410, 100370, 100380, 
    100390, 100400, 100410, 100400, 100400, 100360, 100360, 100350, 100320, 
    100300, 100290, 100280, 100270, 100310, 100290, 100300, 100370, 100400, 
    100380, 100330, 100310, 100280, 100280, 100310, 100320, 100310, 100380, 
    100420, 100500, 100550, 100540, 100640, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 101440, 101510, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 101180, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 101340, 101340, 
    101350, 101330, 101310, 101350, 101310, 101280, 101290, 101240, 101200, 
    101150, 101210, 101190, 101150, 101150, 101110, 101080, 101070, 101070, 
    101040, 101020, 101080, 101110, 101150, 101200, 101250, 101260, 101300, 
    101320, 101310, 101330, 101320, 101310, 101320, 101330, 101350, 101390, 
    101440, 101480, 101510, 101520, 101560, 101580, 101600, 101630, 101660, 
    101690, 101690, 101720, 101750, 101780, 101770, 101750, 101750, 101750, 
    101770, 101790, 101810, 101830, 101830, 101880, 101920, 101940, 101920, 
    101850, 101830, 101800, 101760, 101720, 101680, 101620, 101610, 101640, 
    101690, 101670, 101610, 101590, 101580, 101530, 101490, 101440, 101390, 
    101390, 101320, 101250, 101220, 101170, 101040, 100970, 100940, 100920, 
    100860, 100830, 100790, 100750, 100680, 100640, 100570, 100500, 100420, 
    100310, 100260, 100200, 100130, 100070, 100020, 99990, 99940, 99910, 
    99830, 99750, 99720, 99630, 99580, 99570, 99500, 99400, 99330, 99240, 
    99150, 99070, 98990, 98940, 98860, 98790, 98670, 98600, 98550, 98540, 
    98500, 98390, 98260, 98220, 98190, 98170, 98080, 98040, 98000, 97970, 
    97950, 97880, 97860, 97850, 97830, 97820, 97820, 97830, 97860, 97870, 
    97860, 97880, 97910, 97940, 97980, 98010, 98050, 98110, 98170, 98230, 
    98280, 98350, 98410, 98490, 98540, 98590, 98640, 98680, 98740, 98790, 
    98850, 98930, 98980, 99010, 99050, 99110, 99150, 99180, 99220, 99260, 
    99290, 99310, 99360, 99400, 99450, 99490, 99540, 99590, 99630, 99700, 
    99730, 99800, 99890, 99980, 100050, 100130, 100180, 100230, 100290, 
    100340, 100380, 100440, 100470, 100500, 100530, 100600, 100680, 100720, 
    100750, 100780, 100830, 100860, 100940, 101010, 101030, 101050, 101120, 
    101140, 101160, 101250, 101290, 101310, 101320, 101350, 101360, 101370, 
    101380, 101370, 101370, 101400, 101370, 101380, 101380, 101360, 101350, 
    101320, 101280, 101220, 101180, 101130, 101100, 101050, 101030, 100980, 
    100930, 100890, 100800, 100710, 100650, 100550, 100460, 100360, 100270, 
    100200, 100150, 100090, 100010, 99940, 99900, 99840, 99730, 99700, 99730, 
    99760, 99760, 99720, 99710, 99720, 99730, 99710, 99730, 99760, 99800, 
    99820, 99850, 99850, 99890, 99950, 99960, 99990, 100020, 100030, 100040, 
    100060, 100100, 100110, 100140, 100160, 100180, 100180, 100200, 100210, 
    100230, 100290, 100300, 100270, 100230, 100240, 100200, 100210, 100280, 
    100370, 100370, 100380, 100360, 100350, 100330, 100340, 100350, 100360, 
    100350, 100320, 100380, 100410, 100410, 100440, _, 100390, _, 100420, 
    100440, 100390, 100420, 100500, 100540, 100590, 100600, 100620, 100620, 
    100630, 100620, 100650, 100650, 100650, 100660, 100670, 100650, 100660, 
    100700, 100770, 100790, 100860, 100840, 100900, 100890, 100950, 100960, 
    100940, 100960, 100970, 101000, 101030, 101090, 101100, 101010, 100980, 
    100980, 101000, 101010, 101010, 101030, 101060, 101070, 101090, 101080, 
    101050, 101070, 101060, 101040, 101040, 101000, 100990, 101000, 100990, 
    100990, 101040, 101030, 101060, 101070, 101050, 101020, 101010, 101020, 
    101050, 101130, 101140, _, 101160, 101160, 101170, 101210, 101200, 
    101210, 101200, 101210, 101200, 101200, 101230, 101240, 101260, 101240, 
    101250, 101280, 101260, 101260, 101250, 101270, 101280, 101300, 101310, 
    101360, 101410, 101420, 101400, 101420, 101430, 101490, 101550, 101540, 
    101570, 101620, 101670, 101690, 101720, 101740, 101770, 101800, 101810, 
    101800, 101830, 101840, 101860, 101840, 101850, 101870, 101880, 101850, 
    101800, 101780, 101740, 101640, 101620, 101580, 101540, 101510, 101470, 
    101430, 101450, 101380, 101310, 101290, 101270, 101250, 101220, 101200, 
    101190, 101230, 101320, 101360, 101290, 101280, 101290, 101360, 101400, 
    101390, 101440, 101440, 101450, 101480, 101510, 101550, 101550, _, 
    101670, 101700, 101760, 101730, 101750, 101790, _, 101830, 101850, 
    101870, 101840, 101880, 101910, 101910, 101910, 101900, 101900, 101890, 
    101910, 101880, 101840, 101850, 101810, 101820, 101810, 101790, 101770, 
    101710, 101690, 101680, 101630, 101620, 101570, 101530, 101510, 101510, 
    101500, 101480, 101430, 101390, 101400, 101380, 101380, 101360, 101390, 
    101410, 101410, 101380, 101360, 101340, 101310, 101300, 101250, 101230, 
    101220, 101220, 101220, 101200, 101170, 101130, 101070, 101060, 101050, 
    101050, 101030, 101010, 100980, 101010, 101040, 101070, 101080, 101100, 
    101130, 101150, 101130, 101160, 101180, 101160, 101200, 101220, 101240, 
    101210, 101230, 101200, 101180, 101160, 101120, 101140, 101150, 101150, 
    101130, 101090, 101070, 101050, 101050, 101070, 101070, 101040, 101010, 
    101040, 101000, 100990, 100980, 100940, 100900, 100880, 100810, 100700, 
    100710, 100650, 100530, 100510, 100490, 100400, 100320, 100320, 100280, 
    100190, 100110, 100090, 100060, 100090, 100100, 100060, 100050, 100020, 
    100010, 99920, 99920, 100070, 100080, 100050, 100030, 99980, 99920, 
    99930, 99890, 99820, 99730, 99710, 99700, 99660, 99620, 99550, 99460, 
    99400, 99340, 99280, 99280, 99260, 99140, 99200, 99180, 99170, 99070, 
    98990, 98970, 98940, 98860, 98900, 98940, 98880, 98880, 98830, 98880, 
    98870, 98860, 98850, 98880, 98830, 98840, 98830, 98890, 98950, 98990, 
    99060, 99120, 99180, 99200, 99300, 99370, 99400, 99440, 99500, 99560, 
    99610, 99660, 99720, 99780, 99830, 99880, 99910, 99940, 99960, 100000, 
    100010, 100010, 100040, 100060, 100100, 100130, 100180, 100200, 100200, 
    100200, 100200, 100180, 100170, 100200, 100180, 100200, 100220, 100230, 
    100240, 100210, 100200, 100190, 100200, 100200, 100200, 100220, 100220, 
    100230, 100230, 100240, 100240, 100210, 100170, 100140, 100140, 100120, 
    100110, 100080, 100070, 100000, 99960, 99960, 99930, 99910, 99860, 99810, 
    96750, 99680, 99630, 99580, 99530, 99450, 99380, 99300, 99290, 99260, 
    99220, 99230, 99220, 99160, 99150, 99150, 99120, 99110, 99110, 99100, 
    99140, 99150, 99130, 99150, 99160, 99150, 99180, 99200, 99240, 99290, 
    99320, 99350, 99390, 99410, 99430, 99450, 99460, 99490, 99520, 99540, 
    99540, 99550, 99570, 99580, 99580, 99610, 99650, 99640, 99640, 99640, 
    99650, 99680, 99700, 99750, 99790, 99840, 99910, 99960, 100010, 100040, 
    100070, 100120, 100150, 100180, 100200, 100260, 100290, 100300, 100300, 
    100390, 100430, 100430, 100440, 100480, 100520, 100570, 100600, 100590, 
    100610, 100640, 100670, 100720, 100730, 100740, 100760, 100770, 100760, 
    100750, 100770, 100770, 100760, 100750, 100760, 100710, 100630, 100650, 
    100690, 100680, 100670, 100660, 100630, 100640, 100590, 100590, 100580, 
    100590, 100590, 100590, 100590, 100600, 100600, 100610, 100580, 100550, 
    100560, 100560, 100610, 100620, 100620, 100650, 100660, 100660, 100680, 
    100680, 100680, 100710, 100730, 100740, 100770, 100800, 100760, 100780, 
    100820, 100890, 100880, 100910, 100910, 100950, 100960, 100970, 100980, 
    101020, 101000, 100960, 101020, 101030, 101060, 101080, 101110, 101150, 
    101190, 101170, 101210, 101250, 101290, 101350, 101380, 101340, 101340, 
    101360, 101380, 101410, 101440, 101440, 101430, 101450, 101450, 101460, 
    101460, 101480, 101500, 101470, 101470, 101500, 101530, 101560, 101580, 
    101610, 101620, 101590, 101610, 101630, 101630, 101610, 101630, 101630, 
    101670, 101660, 101630, 101640, 101600, 101590, 101550, 101530, 101500, 
    101450, 101410, 101390, 101420, 101390, 101390, 101450, 101400, 101430, 
    101430, 101430, 101400, 101440, 101420, 101430, 101430, 101430, 101430, 
    101420, 101400, 101380, 101370, 101370, 101360, 101360, 101340, 101330, 
    101340, 101350, 101350, 101330, 101320, 101330, 101320, 101310, 101310, 
    101300, 101290, 101280, 101290, 101300, 101300, 101310, 101300, 101300, 
    101310, 101310, 101320, 101310, 101340, 101340, 101370, 101390, 101400, 
    101410, 101410, 101420, 101430, 101410, 101410, 101420, 101410, 101410, 
    101430, 101430, 101470, 101470, 101470, 101480, 101470, 101490, 101480, 
    101480, 101490, 101500, 101510, 101560, 101560, 101530, 101550, 101560, 
    101530, 101510, 101490, 101440, 101410, 101390, 101390, 101370, 101320, 
    101310, 101270, 101250, 101230, 101200, 101180, 101150, 101130, 101110, 
    101080, 101050, 101010, 101000, 100970, 100960, 100940, 100910, 100870, 
    100840, 100810, 100800, 100790, 100790, 100770, 100760, 100750, 100730, 
    100740, 100730, 100720, 100710, 100710, 100710, 100710, 100730, 100770, 
    100770, 100730, 100770, 100800, 100790, 100760, 100760, 100770, 100770, 
    100780, 100810, 100850, 100860, 100880, 100870, 100870, 100860, 100860, 
    100880, 100870, 100890, 100890, 100910, 100950, 100980, 101000, 101020, 
    100990, 101020, 101020, 101010, 100990, 101000, 101010, 100990, 100980, 
    100950, 100930, 100940, 100940, 100970, 100940, 100930, 100920, 100940, 
    100930, 100940, 100920, 100920, 100940, 100930, 100950, 100920, 100900, 
    100900, 100920, 100960, 100970, 101030, 101050, 101090, 101140, 101150, 
    101190, 101230, 101250, 101240, 101260, 101320, 101350, 101370, 101380, 
    101460, 101480, 101530, 101570, 101590, 101610, 101620, 101610, 101620, 
    101670, 101720, 101720, 101760, 101820, 101850, 101850, 101890, 101900, 
    101940, 101930, 101950, 101950, 102010, 102070, 102130, 102140, 102160, 
    102180, 102190, 102210, 102210, 102230, 102250, 102280, 102280, 102300, 
    102300, 102300, 102290, 102300, 102300, 102300, 102320, 102340, 102360, 
    102380, 102400, 102400, 102380, 102370, 102380, 102380, 102380, 102360, 
    102370, 102370, 102360, 102360, 102360, 102370, 102360, 102350, 102320, 
    102310, 102310, 102300, 102310, 102300, 102300, 102310, 102320, 102310, 
    102300, 102310, 102300, 102300, 102280, 102250, 102230, 102190, 102200, 
    102210, 102220, 102220, 102220, 102210, 102200, 102190, 102190, 102170, 
    102150, 102140, 102140, 102170, 102180, 102190, 102160, 102160, 102150, 
    102130, 102100, 102080, 102070, 102090, 102110, 102120, 102150, 102170, 
    102180, 102180, 102210, 102240, 102260, 102260, 102270, 102310, 102340, 
    102370, 102400, 102410, 102430, 102430, 102380, 102440, 102450, 102460, 
    102430, 102480, 102520, 102520, 102560, 102540, 102530, 102510, 102520, 
    102460, 102430, 102320, 102340, 102250, 102070, 102100, 101990, 102010, 
    101930, 101850, 101680, 101430, 101360, 101230, 101080, 101020, 100900, 
    100850, 100750, 100570, 100450, 100390, 100330, 100310, 100290, 100270, 
    100230, 100260, 100250, 100240, 100280, 100340, 100380, 100420, 100450, 
    100480, 100510, _, 100560, 100560, 100580, 100610, 100630, 100650, 
    100650, 100660, 100660, 100640, 100640, 100620, 100620, 100600, 100550, 
    100550, 100520, 100510, 100470, 100420, 100380, 100350, 100350, 100320, 
    100320, 100300, 100320, 100310, 100350, 100330, 100390, 100430, 100480, 
    100520, 100620, 100690, 100770, 100870, 100950, 101080, 101200, 101280, 
    101340, 101380, 101400, 101450, 101500, 101510, 101540, 101540, 101520, 
    101540, 101530, 101500, 101480, 101440, 101400, 101370, 101290, 101250, 
    101200, 101140, 101050, 101010, 100970, 100930, 100890, 100880, 100870, 
    100860, 100840, 100840, 100840, 100830, 100860, 100860, 100860, 100810, 
    100820, 100790, 100840, 100850, 100840, 100820, 100830, 100830, 100830, 
    100820, 100790, 100750, 100720, 100670, 100650, 100620, 100590, 100570, 
    100590, 100550, 100510, 100490, 100460, 100410, 100360, 100330, 100360, 
    100330, 100310, 100260, 100210, 100200, 100240, 100300, 100370, 100430, 
    100440, 100490, 100530, 100560, 100610, 100610, 100670, 100710, 100750, 
    100820, 100860, 100840, 100990, 100990, 101040, 101080, 101150, 101190, 
    101210, 101230, 101290, 101350, 101390, 101450, 101470, 101520, 101580, 
    101620, 101670, 101710, 101740, 101760, 101790, 101830, 101850, 101900, 
    101910, 101930, 101930, 101940, 101980, 101990, 102010, 102030, 102040, 
    102080, 102080, 102090, 102090, 102110, 102120, 102130, 102160, 102150, 
    102160, 102170, 102160, 102160, 102160, 102150, 102160, 102170, 102160, 
    102140, 102130, 102120, 102130, 102140, 102130, 102140, 102140, 102150, 
    102170, 102200, 102210, 102240, 102250, 102260, 102260, 102270, 102310, 
    102350, 102380, 102370, 102380, 102370, 102390, 102390, 102390, 102380, 
    102390, 102410, 102410, 102450, 102440, 102440, 102460, 102480, 102470, 
    102480, 102460, 102450, 102440, 102450, 102460, 102450, 102440, 102430, 
    102430, 102430, 102420, 102410, 102390, 102380, 102370, 102350, 102350, 
    102350, 102350, 102320, 102300, 102280, 102260, 102250, 102230, 102210, 
    102180, 102150, 102150, 102130, 102100, 102090, 102060, 102020, 102000, 
    101970, 101940, 101910, 101880, 101870, 101840, 101820, 101790, 101740, 
    101700, 101680, 101640, 101600, 101550, 101510, 101470, 101430, 101400, 
    101350, 101340, 101320, 101290, 101240, 101210, 101170, 101140, 101100, 
    101100, 101090, 101070, 101060, 101060, 101080, 101090, 101090, 101100, 
    101110, 101110, 101100, 101100, 101110, 101110, 101130, 101170, 101160, 
    101180, 101220, 101230, 101240, 101230, 101240, 101260, 101270, 101290, 
    101320, 101330, 101350, 101370, 101380, 101400, 101400, 101400, 101380, 
    101390, 101390, 101390, 101400, 101410, 101390, 101380, 101370, 101350, 
    101370, 101350, 101320, 101350, 101330, 101320, 101320, 101310, 101310, 
    101280, 101260, 101270, 101270, 101260, 101240, 101220, 101200, 101170, 
    101150, 101150, 101160, 101170, 101180, 101190, 101150, 101130, 101120, 
    101120, 101140, 101170, 101200, 101230, 101270, 101290, 101360, 101410, 
    101440, 101490, 101500, 101560, 101590, 101600, 101630, 101670, 101690, 
    101670, 101660, 101660, 101660, 101670, 101810, 101840, 101890, 101930, 
    101980, 102000, 102050, 102110, 102170, 102200, 102230, 102220, 102240, 
    102260, 102270, 102290, 102320, 102330, 102350, 102340, 102360, 102350, 
    102390, 102390, 102390, 102390, 102410, 102440, 102400, 102420, 102430, 
    102440, 102470, 102470, 102490, 102480, 102470, 102430, 102440, 102470, 
    102470, 102470, 102430, 102420, 102420, 102440, 102460, 102430, 102430, 
    102430, 102440, 102440, 102470, 102470, 102490, 102520, 102520, 102540, 
    102520, 102520, 102530, 102540, 102550, 102570, 102590, 102600, 102610, 
    102630, 102640, 102650, 102660, 102660, 102660, 102660, 102670, 102700, 
    102730, 102740, 102740, 102740, 102750, 102750, 102740, 102740, 102740, 
    102720, 102720, 102730, 102750, 102770, 102750, 102750, 102760, 102750, 
    102760, 102750, 102730, 102720, 102730, 102750, 102750, 102740, 102740, 
    102740, 102710, 102710, 102690, 102650, 102640, 102620, 102600, 102590, 
    102590, 102590, 102570, 102540, 102490, 102480, 102460, 102430, 102390, 
    102350, 102320, 102300, 102300, 102290, 102280, 102230, 102180, 102150, 
    102120, 102080, 102040, 102000, 101980, 101930, 101920, 101890, 101850, 
    101780, 101720, 101670, 101580, 101510, 101420, 101370, 101330, 101270, 
    101160, 101100, 100990, 101010, 100990, 100950, 100890, 100830, 100780, 
    100730, 100670, 100620, 100590, 100570, 100530, 100500, 100460, 100430, 
    100410, 100430, 100390, 100450, 100480, 100490, 100510, 100550, 100610, 
    100650, 100660, 100690, 100740, 100800, 100830, 100840, 100890, 100940, 
    100980, 101020, 101080, 101120, 101130, 101170, 101200, 101220, 101240, 
    101300, 101350, 101370, 101420, 101440, 101510, 101560, 101600, 101630, 
    101670, 101720, 101750, 101780, 101800, 101810, 101840, 101880, 101900, 
    101920, 101950, 101960, 101990, 102000, 102030, 102000, 102030, 102060, 
    102080, 102110, 102090, 102140, 102150, 102150, 102170, 102170, 102190, 
    102180, 102180, 102170, 102160, 102150, 102170, 102200, 102190, 102180, 
    102150, 102150, 102140, 102120, 102080, 102040, 101980, 101950, 101890, 
    101840, 101780, 101700, 101610, 101530, 101460, 101340, 101270, 101220, 
    101160, 101150, 101120, 101090, 101090, 101070, 101030, 101010, 101010, 
    100970, 100910, 100880, 100880, 100880, 100860, 100840, 100800, 100800, 
    100780, 100770, 100770, 100760, 100730, 100750, 100770, 100810, 100820, 
    100810, 100790, 100810, 100810, 100790, 100770, 100780, 100770, 100760, 
    100770, 100770, 100780, 100790, 100770, 100770, 100760, 100770, 100770, 
    100770, 100770, 100760, 100730, 100740, 100740, 100720, 100700, 100690, 
    100670, 100640, 100590, 100570, 100560, 100570, 100530, 100510, 100470, 
    100410, 100370, 100280, 100200, 100110, 100010, 99890, 99810, 99680, 
    99560, 99470, 99350, 99240, 99150, 99040, 98910, 98810, 98720, 98630, 
    98530, 98480, 98430, 98360, 98280, 98200, 98120, 98030, 97930, 97820, 
    97710, 97570, 97440, 97330, 97210, 97050, 96980, 96920, 96890, 96890, 
    96880, 96890, 96890, 96900, 96950, 97020, 97090, 97180, 97220, 97340, 
    97400, 97490, 97610, 97780, 97800, 97940, 97990, 98030, 98180, 98240, 
    98320, 98410, 98480, 98560, 98660, 98720, 98780, 98820, 98870, 98960, 
    99030, 99120, 99210, 99290, 99340, 99390, 99400, 99440, 99500, 99530, 
    99540, 99550, 99550, 99560, 99570, 99600, 99630, 99620, 99590, 99560, 
    99600, 99580, 99580, 99610, 99640, 99680, 99700, 99720, 99730, 99820, 
    99820, 99820, 99790, 99780, 99760, 99750, 99840, 99880, 99920, 99930, 
    99970, 100030, 100080, 100160, 100210, 100250, 100280, 100320, 100310, 
    100400, 100450, 100510, 100540, 100600, 100640, 100680, 100720, 100780, 
    100840, 100910, 100980, 100980, 101010, 101060, 101130, 101160, 101170, 
    101180, 101220, 101260, 101270, 101330, 101380, 101420, 101440, 101450, 
    101480, 101510, 101540, 101540, 101540, 101560, 101570, 101600, 101610, 
    101620, 101620, 101620, 101640, 101660, 101670, 101660, 101640, 101650, 
    101660, 101670, 101700, 101720, 101720, 101700, 101710, 101690, 101680, 
    101690, 101670, 101650, 101670, 101680, 101700, 101700, 101700, 101690, 
    101690, 101690, 101700, 101720, 101740, 101750, 101800, 101830, 101830, 
    101900, 101910, 101920, 101940, 101950, 101950, 101960, 101950, 101940, 
    101930, 101910, 101960, 101990, 102010, 102030, 102030, 102070, 102080, 
    102070, 102060, 102040, 102010, 102040, 102030, 102030, 102020, 102000, 
    101990, 102010, 102040, 102040, 102050, 102010, 102040, 102020, 101950, 
    101900, 101860, 101800, 101760, 101730, 101670, 101610, 101590, 101530, 
    101490, 101490, 101510, 101520, 101560, 101570, 101580, 101590, 101600, 
    101630, 101660, 101640, 101660, 101720, 101770, 101770, 101820, 101770, 
    101790, 101800, 101810, 101800, 101850, 101850, 101830, 101880, 101900, 
    101920, 101900, 101920, 101930, 101950, 101960, 101960, 101990, 101950, 
    101960, 101990, 102000, 102040, 102060, 102070, 102080, 102070, 102090, 
    102080, 102070, 102080, 102100, 102090, 102100, 102060, 102020, 101950, 
    101920, 101940, 101920, 101900, 101860, 101820, 101800, 101800, 101800, 
    101740, 101690, 101720, 101720, 101720, 101700, 101670, 101660, 101630, 
    101570, 101530, 101550, 101540, 101580, 101490, 101580, 101610, 101630, 
    101600, 101620, 101610, 101610, 101630, 101630, 101630, 101670, 101670, 
    101680, 101680, 101720, 101710, 101700, 101700, 101720, 101760, 101770, 
    101810, 101820, 101820, 101850, 101860, 101880, 101880, 101900, 101880, 
    101880, 101890, 101920, 101910, 101910, 101900, 101870, 101860, 101840, 
    101850, 101820, 101790, 101780, 101790, 101780, 101780, 101770, 101760, 
    101760, 101750, 101740, 101710, 101660, 101630, 101600, 101590, 101600, 
    101590, 101570, 101540, 101530, 101540, 101520, 101510, 101480, 101470, 
    101430, 101410, 101430, 101430, 101450, 101470, 101460, 101480, 101450, 
    101440, 101440, 101420, 101410, 101430, 101410, 101430, 101430, 101440, 
    101410, 101410, 101410, 101420, 101410, 101420, 101440, 101450, 101480, 
    101480, 101470, 101490, 101490, 101510, 101520, 101520, 101530, 101540, 
    101560, 101570, 101590, 101620, 101610, 101630, 101640, 101690, 101700, 
    101710, 101730, 101740, 101760, 101800, 101840, 101880, 101910, 101920, 
    101950, 101910, 101940, 101910, 101940, 101940, 102000, 101990, 102030, 
    102060, 102080, 102110, 102100, 102110, 102130, 102150, 102190, 102180, 
    102130, 102140, 102210, 102170, 102200, 102210, 102200, 102190, 102160, 
    102170, 102140, 102090, 102120, 102120, 102080, 102100, 102050, 101980, 
    101940, 101900, 101840, 101830, 101770, 101720, 101670, 101620, 101600, 
    101610, 101560, 101520, 101460, 101440, 101420, 101410, 101460, 101470, 
    101490, 101480, 101480, 101490, 101500, 101510, 101550, 101560, 101540, 
    101580, 101590, 101650, 101620, 101660, 101720, 101720, 101750, 101740, 
    101750, 101750, 101760, 101750, 101750, 101730, 101700, 101690, 101690, 
    101690, 101660, 101660, 101660, 101650, 101630, 101610, 101580, 101560, 
    101540, 101550, 101570, 101570, 101540, 101550, 101540, 101560, 101570, 
    101560, 101570, 101590, 101610, 101630, 101640, 101680, 101720, 101750, 
    101750, 101750, 101770, 101780, 101810, 101820, 101830, 101850, 101890, 
    101910, 101930, 101950, 101980, 101980, 101990, 101990, 101990, 101980, 
    101960, 101980, 101990, 101990, 101990, 101940, 101940, 101920, 101860, 
    101840, 101820, 101800, 101770, 101760, 101770, 101750, 101760, 101760, 
    101740, 101730, 101700, 101710, 101670, 101620, 101610, 101570, 101520, 
    101490, 101450, 101410, 101410, 101380, 101400, 101360, 101340, 101340, 
    101310, 101290, 101280, 101260, 101230, 101200, 101200, 101200, 101170, 
    101130, 101080, 101100, 101100, 101100, 101080, 101050, 101010, 101010, 
    101020, 101000, 101000, 100990, 100980, 101000, 100990, 100980, 100980, 
    100960, 100960, 100950, 100940, 100900, 100880, 100850, 100830, 100820, 
    100780, 100750, 100740, 100710, 100680, 100600, 100540, 100520, 100480, 
    100430, 100410, 100380, 100380, 100380, 100360, 100350, 100340, 100360, 
    100340, 100320, 100310, 100320, 100300, 100290, 100290, 100300, 100310, 
    100300, 100280, 100250, 100250, 100240, 100240, 100230, 100220, 100230, 
    100240, 100250, 100250, 100270, 100310, 100330, 100340, 100360, 100360, 
    100370, 100370, 100380, 100360, 100370, 100380, 100400, 100390, 100390, 
    100370, 100360, 100350, 100330, 100320, 100310, 100310, 100270, 100260, 
    100250, 100240, 100200, 100170, 100150, 100140, 100100, 100100, 100090, 
    100090, 100090, 100070, 100070, 100080, 100100, 100130, 100150, 100150, 
    100160, 100190, 100220, 100250, 100270, 100310, 100350, 100370, 100410, 
    100420, 100470, 100500, 100520, 100540, 100580, 100650, 100660, 100690, 
    100740, 100770, 100790, 100810, 100850, 100880, 100910, 100930, 100970, 
    100980, 101010, 101060, 101070, 101070, 101090, 101100, 101120, 101110, 
    101100, 101100, 101090, 101080, 101060, 101050, 101020, 100990, 100990, 
    100980, 100950, 100900, 100850, 100830, 100810, 100790, 100770, 100750, 
    100710, 100660, 100630, 100600, 100580, 100560, 100530, 100520, 100500, 
    100500, 100500, 100500, 100530, 100540, 100540, 100550, 100560, 100570, 
    100580, 100590, 100640, 100670, 100700, 100740, 100760, 100790, 100810, 
    100860, 100860, 100880, 100890, 100930, 100970, 100990, 101000, 101040, 
    101030, 101060, 101090, 101120, 101140, 101180, 101200, 101190, 101200, 
    101230, 101250, 101270, 101290, 101280, 101280, 101300, 101290, 101280, 
    101260, 101200, 101180, 101140, 101140, 101090, 101010, 100980, 100920, 
    100920, 100920, 100880, 100760, 100710, 100680, 100670, 100690, 100690, 
    100680, 100720, 100670, 100680, 100700, 100710, 100740, 100740, 100740, 
    100750, 100780, 100770, 100810, 100800, 100810, 100840, 100850, 100860, 
    100870, 100860, 100900, 100920, 100920, 100950, 100960, 100990, 101010, 
    101020, 101010, 101010, 101030, 101070, 101080, 101090, 101100, 101080, 
    101100, 101110, 101110, 101090, 101100, 101080, 101080, 101090, 101100, 
    101070, 101060, 101070, 101100, 101100, 101110, 101090, 101110, 101110, 
    101100, 101110, 101120, 101150, 101160, 101170, 101190, 101220, 101220, 
    101220, 101250, 101270, 101290, 101320, 101330, 101340, 101370, 101390, 
    101430, 101440, 101460, 101470, 101480, 101530, 101550, 101560, 101580, 
    101590, 101590, 101620, 101660, 101660, 101670, 101690, 101710, 101720, 
    101730, 101740, 101760, 101770, 101790, 101810, 101840, 101850, 101850, 
    101870, 101890, 101880, 101870, 101900, 101910, 101920, 101930, 101950, 
    101980, 101970, 101930, 101980, 101990, 102030, 102060, 102060, 102090, 
    102140, 102170, 102200, 102220, 102270, 102310, 102320, 102360, 102380, 
    102400, 102400, 102390, 102390, 102380, 102390, 102400, 102380, 102370, 
    102400, 102370, 102360, 102310, 102290, 102250, 102210, 102180, 102140, 
    102080, 102040, 101980, 101910, 101850, 101760, 101690, 101590, 101540, 
    101430, 101410, 101370, 101270, 101200, 101130, 101100, 101050, 101020, 
    100980, 100920, 100960, 100930, 100950, 100950, 100960, 100980, 100980, 
    100990, 100980, 100980, 101000, 100970, 100980, 100980, 100990, 100990, 
    100990, 100990, 100990, 100980, 100990, 100970, 100970, 100970, 100950, 
    100940, 100950, 100940, 100940, 100900, 100890, 100850, 100790, 100690, 
    100610, 100530, 100430, 100340, 100220, 100180, 100130, 100110, 100060, 
    100070, 100050, 100000, 99980, 99930, 99930, 99930, 99890, 99890, 99840, 
    99790, 99770, 99850, 99850, 99850, 99790, 99780, 99760, 99780, 99840, 
    99900, 99940, 99980, 100040, 100050, 100080, 100100, 100110, 100120, 
    100180, 100210, 100240, 100300, 100320, 100350, 100360, 100380, 100400, 
    100410, 100420, 100440, 100460, 100470, 100490, 100510, 100530, 100550, 
    100560, 100560, 100570, 100580, 100580, 100590, 100610, 100630, 100710, 
    100760, 100770, 100790, 100820, 100830, 100840, 100820, 100800, 100850, 
    100860, 100880, 100900, 100970, 100980, 100960, 101020, 101040, 101060, 
    101070, 101040, 101060, 101050, 101060, 101070, 101090, 101090, 101090, 
    101110, 101110, 101110, 101050, 101000, 100960, 100950, 100910, 100910, 
    100890, 100870, 100840, 100840, 100810, 100790, 100760, 100740, 100740, 
    100740, 100750, 100780, 100810, 100820, 100830, 100860, 100890, 100900, 
    100910, 100920, 100940, 100970, 100990, 100990, 101010, 101040, 101040, 
    101050, 101050, 101050, 101020, 101000, 101010, 101010, 101000, 101000, 
    100990, 100970, 100980, 100960, 100930, 100920, 100910, 100870, 100840, 
    100850, 100870, 100850, 100840, 100810, 100790, 100760, 100730, 100730, 
    100710, 100690, 100660, 100620, 100600, 100570, 100550, 100530, 100530, 
    100520, 100480, 100430, 100400, 100370, 100330, 100290, 100310, 100310, 
    100310, 100330, 100310, 100330, 100310, 100300, 100270, 100230, 100230, 
    100260, 100290, 100290, 100300, 100270, 100280, 100280, 100310, 100300, 
    100290, 100300, 100310, 100310, 100320, 100340, 100350, 100370, 100360, 
    100350, 100370, 100350, 100380, 100390, 100400, 100420, 100440, 100450, 
    100470, 100500, 100530, 100560, 100600, 100590, 100610, 100630, 100660, 
    100670, 100700, 100710, 100710, 100710, 100720, 100710, 100710, 100710, 
    100700, 100680, 100660, 100710, 100710, 100710, 100750, 100740, 100740, 
    100750, 100750, 100810, 100820, 100840, 100860, 100870, 100900, 100910, 
    100930, 100940, 100950, 100970, 100970, 100970, 101000, 101030, 101030, 
    101020, 101260, 101100, 101130, 101170, 101210, 101230, 101270, 101320, 
    101310, 101350, 101350, 101390, 101420, 101420, 101460, 101470, 101490, 
    101480, 101450, 101480, 101470, 101450, 101440, 101490, 101510, 101540, 
    101540, 101500, 101480, 101460, 101480, 101470, 101460, 101420, 101400, 
    101390, 101390, 101320, 101280, 101240, 101190, 101130, 101120, 101090, 
    100980, 100960, 100930, 100880, 100940, 100900, 100800, _, 100730, 
    100730, 100660, 100550, 100580, _, 100520, 100480, 100490, 100420, 
    100360, 100320, 100300, 100260, 100190, 100150, 100120, 100060, 100020, 
    99910, 99870, 99850, 99920, 99770, 99750, 99730, 99740, 99780, 99790, 
    99810, 99750, 99760, 99690, 99650, 99690, 99620, 99530, 99520, 99430, 
    99530, 99430, 99450, 99360, 99400, 99400, 99360, 99380, 99430, 99400, 
    99470, 99440, 99440, 99480, 99470, 99490, 99480, 99430, 99380, 99400, 
    99400, 99380, 99370, _, 99430, 99480, 99510, 99560, 99620, 99680, 99720, 
    99780, _, 99870, 99920, 99960, 99970, 100010, 100020, 100020, 100020, 
    100030, 100030, 100020, 100010, 99940, 99940, 99910, 99890, 99880, 99820, 
    99740, 99730, 99720, 99740, 99760, 99780, 99790, 99810, 99800, 99840, 
    99870, 99900, 99910, 99940, 99970, 99990, 100010, 100000, 100000, 100040, 
    100010, 100030, 100040, 100040, 100050, 100050, 100060, 100080, 100140, 
    100140, 100200, 100240, 100250, 100250, 100270, 100310, 100300, 100360, 
    100390, 100440, 100480, 100500, 100520, 100510, 100530, 100530, 100550, 
    100550, 100570, 100580, 100590, 100620, 100650, 100660, 100680, 100680, 
    100700, 100730, 100740, 100740, 100750, 100770, 100750, 100780, 100800, 
    100800, 100800, 100810, 100800, 100800, 100810, 100830, 100840, 100830, 
    100830, 100840, 100840, 100860, 100850, 100860, 100860, 100850, 100850, 
    100850, 100860, 100860, 100880, 100870, _, 100890, 100870, 100890, 
    100910, 100900, 100900, 100890, 100880, 100910, 100880, 100860, 100860, 
    100810, 100800, 100800, 100770, 100740, 100700, 100670, 100660, 100570, 
    100490, 100410, 100340, 100300, 100210, 100110, _, 100010, 99940, 99870, 
    99840, 99800, 99800, _, 99820, 99860, 99880, 99890, 99900, 99910, 99980, 
    99950, 100100, 100220, 100310, 100310, 100410, 100450, 100520, 100550, 
    100590, 100600, 100510, 100480, 100550, 100600, 100590, 100600, 100600, 
    100660, 100760, 100820, 100890, 100930, 100980, 100980, 101040, 101060, 
    101100, 101060, 101040, 101030, 101100, 101130, 101160, 101130, 101170, 
    101200, 101210, 101220, 101220, _, 101290, 101280, 101310, 101270, 
    101270, 101300, 101300, 101270, 101260, _, 101250, 101260, 101210, 
    101190, 101180, 101200, 101170, 101120, 101070, 101050, 101030, 101020, 
    100980, 100950, 100930, 100920, _, 100880, 100850, 100820, 100770, 
    100740, 100730, 100680, 100650, 100610, 100560, 100520, 100490, 100450, 
    100400, 100390, 100390, 100360, 100300, 100290, 100280, 100320, 100320, 
    100310, 100310, 100310, 100310, 100300, 100290, 100280, 100250, 100250, 
    100240, 100230, 100220, 100240, 100240, 100210, 100210, 100190, 100180, 
    100160, 100150, 100140, 100170, 100180, 100170, 100170, 100170, 100150, 
    100160, 100160, 100160, 100150, 100150, 100080, 100080, 100050, 100090, 
    100100, 100080, 100130, 100130, 100110, 100110, 100100, 100090, 100090, 
    100090, 100090, 100080, 100080, 100090, 100070, 100060, 100050, 100030, 
    100000, 100010, 99990, 99990, 100000, 99990, 99990, 100000, 100000, 
    99990, 100000, 99990, 99970, 99970, 99980, 99990, 100020, 100030, 100050, 
    100070, 100070, 100080, 100080, 100100, 100080, 100110, 100120, 100140, 
    100160, 100190, 100230, 100250, 100250, 100260, 100270, 100280, 100300, 
    100320, _, 100410, 100450, 100460, 100500, 100520, 100550, 100540, 
    100550, 100550, _, 100530, 100530, 100490, 100460, 100440, 100420, 
    100390, 100370, 100360, 100330, 100300, 100300, 100250, 100230, 100200, 
    100230, 100260, 100270, 100270, 100290, 100330, 100370, 100430, 100420, 
    100440, 100470, 100400, 100470, 100540, 100500, 100540, _, 100570, 
    100600, 100580, 100570, 100580, 100570, 100570, 100550, 100550, 100530, 
    100540, 100530, 100510, 100480, 100490, 100480, 100460, 100430, 100420, 
    100410, 100400, 100400, 100360, 100310, 100260, 100230, 100200, 100140, 
    100090, 100070, 100030, 99990, 99960, 99900, 99850, 99780, 99730, 99680, 
    99620, 99580, 99480, 99440, 99400, 99360, 99320, 99300, 99280, 99270, 
    99230, 99210, 99180, 99170, 99180, 99180, 99210, 99240, 99270, 99320, 
    99360, 99390, 99400, 99440, 99490, 99530, 99590, 99630, 99660, 99720, 
    99810, 99890, 99960, 100040, 100120, 100170, 100210, 100290, 100310, 
    100400, 100450, 100530, 100570, 100560, 100640, 100720, 100760, 100800, 
    100830, 100790, 100830, 100850, 100850, 100890, 100880, 100890, 100920, 
    100920, 100900, 100870, 100880, 100870, 100870, 100890, 100880, 100910, 
    100930, 100950, 100940, 100950, 100930, 100930, 100950, 100950, 100960, 
    100980, 101010, 101020, 101030, 101060, 101100, 101170, 101210, 101260, 
    101310, 101360, 101390, 101380, 101400, 101420, 101470, 101540, 101550, 
    101660, 101700, 101650, 101660, 101630, 101630, 101640, 101630, 101620, 
    101660, 101680, 101670, 101660, 101620, 101600, 101590, 101570, 101560, 
    101560, 101570, 101590, 101610, 101610, 101630, 101600, 101590, 101600, 
    101560, 101670, 101690, 101740, 101740, 101760, 101740, 101710, 101700, 
    101660, 101630, 101610, 101590, 101560, 101530, 101500, 101470, 101460, 
    101440, 101410, 101400, 101380, 101360, 101360, 101340, 101330, 101320, 
    101280, 101280, 101290, 101310, 101310, 101280, 101320, 101320, 101290, 
    101270, 101270, 101270, 101260, 101250, 101250, 101260, 101280, 101280, 
    101270, 101280, 101260, 101230, 101250, 101210, 101190, 101260, 101220, 
    101230, 101240, 101300, 101350, 101380, 101410, 101450, 101480, 101510, 
    101560, 101540, 101590, 101620, 101650, 101680, 101670, 101700, 101680, 
    101670, 101700, 101720, 101730, 101740, 101690, 101700, 101690, 101700, 
    101680, 101640, 101580, 101540, 101480, 101440, 101420, 101380, 101290, 
    101250, 101220, 101180, 101150, 101060, 100990, 100920, 100860, 100720, 
    100620, 100460, 100350, 100180, 100070, 99960, 99890, 99760, 99650, 
    99580, 99570, 99640, 99660, 99640, 99630, 99610, 99600, 99580, 99570, 
    99550, 99530, 99460, 99380, 99350, 99310, 99240, 99200, 99170, 99150, 
    99110, 99120, 99180, 99200, 99220, 99270, 99290, 99340, 99340, 99430, 
    99450, 99440, 99390, 99390, 99310, 99340, 99370, 99360, 99350, 99330, 
    99340, 99330, 99380, 99410, 99420, 99320, 99400, 99440, 99460, 99480, 
    99510, 99540, 99570, 99590, 99620, 99630, 99640, 99630, 99660, 99670, 
    99660, 99630, 99600, 99590, 99570, 99580, 99600, 99620, 99670, 99710, 
    99760, 99830, 99870, 99910, 99940, 99980, 100040, 100060, 100090, 100160, 
    100180, 100180, 100200, 100260, 100290, 100320, 100400, 100510, 100560, 
    100600, 100630, 100770, 100840, 100900, 100960, 100990, 101040, 101070, 
    101100, 101130, 101170, 101210, 101240, 101280, 101310, 101320, 101330, 
    101320, 101330, 101340, 101360, 101370, 101380, 101380, 101400, 101410, 
    101430, 101450, 101460, 101470, 101470, 101450, 101440, 101460, 101480, 
    101490, 101510, 101510, 101520, 101520, 101540, 101530, 101530, 101520, 
    101540, 101560, 101580, 101630, 101660, 101680, 101700, 101730, 101750, 
    101770, 101770, 101790, 101830, 101850, 101870, 101890, 101910, 101940, 
    101950, 101960, 101980, 101980, 101980, 101990, 102010, 102020, 102040, 
    102050, 102080, 102080, 102080, 102070, 102070, 102060, 102070, 102070, 
    102080, 102090, 102080, 102090, 102110, 102120, 102100, 102110, 102120, 
    102120, 102110, 102090, 102080, 102080, 102080, 102050, 102040, 102040, 
    102050, 102010, 102020, 101960, 101920, 101870, 101860, 101840, 101800, 
    101810, 101760, 101740, 101760, 101800, 101860, 101870, 101930, 101970, 
    101980, 102020, 102050, 102070, 102110, 102140, 102150, 102140, 102130, 
    102110, 102130, 102160, 102090, 102070, 102050, 102000, 101940, 101900, 
    101840, 101800, 101700, 101650, 101520, 101480, 101410, 101390, 101350, 
    101310, 101270, 101260, 101230, 101200, 101200, 101210, 101210, 101240, 
    101280, 101320, 101340, 101370, 101380, 101430, 101450, 101460, 101490, 
    101420, 101450, 101410, 101380, 101430, 101390, 101420, 101450, 101460, 
    101490, 101540, 101540, 101570, 101550, 101530, 101500, 101470, 101400, 
    101350, 101290, 101130, 101070, 100990, 100860, 100870, 100810, 100720, 
    100630, 100570, 100490, 100430, 100400, 100370, 100300, 100200, 100180, 
    100150, 100140, 100090, 100080, 100180, 100160, 100200, 100220, 100230, 
    100270, 100290, 100300, 100290, 100300, 100320, 100340, 100370, 100380, 
    100400, 100440, 100470, 100470, 100480, 100490, 100460, 100420, 100400, 
    100370, 100340, 100290, 100250, 100190, 100110, 99990, 99860, 99740, 
    99650, 99570, 99470, 99440, 99460, 99460, 99460, 99460, 99490, 99500, 
    99500, 99510, 99520, 99530, 99560, 99570, 99570, 99580, 99630, 99620, 
    99640, 99640, 99610, 99660, 99640, 99620, 99590, 99550, 99510, 99460, 
    99390, 99400, 99360, 99340, 99340, 99310, 99280, 99260, 99240, 99200, 
    99170, 99140, 99110, 99050, 99040, 99030, 99030, 99020, 98990, 98990, 
    99000, 98970, 98970, 98950, 98930, 98930, 98930, 98910, 98880, 98880, 
    98910, 98920, 98920, 98940, 98960, 99000, 99030, 99060, 99100, 99160, 
    99200, 99240, 99250, 99270, 99290, 99310, 99300, 99320, 99310, 99320, 
    99330, 99310, 99300, 99270, 99240, 99250, 99280, 99300, 99340, 99350, 
    99380, 99430, 99460, 99490, 99510, 99500, 99440, 99470, 99440, 99440, 
    99460, 99420, 99450, 99480, 99440, 99430, 99470, 99470, 99490, 99520, 
    99480, 99510, 99540, 99580, 99610, 99640, 99650, 99630, 99630, 99600, 
    99650, 99590, 99670, 99810, 99830, 99810, 99830, 99800, 99830, 99830, 
    99810, 99810, 99820, 99810, 99810, 99800, 99790, 99790, 99800, 99810, 
    99820, 99810, 99840, 99840, 99830, 99840, 99860, 99840, 99850, 99890, 
    99900, 99870, 99910, 99910, 99930, 99930, 99880, 99940, 99950, 99920, 
    99970, 100030, 100090, 100130, 100150, 100180, 100220, 100260, 100280, 
    100330, 100370, 100380, 100390, 100420, 100460, 100490, 100520, 100530, 
    100570, 100590, 100620, 100650, 100670, 100690, 100700, 100710, 100730, 
    100770, 100800, 100850, 100880, 100900, 100920, 100940, 100950, 100980, 
    101010, 101040, 101060, 101090, 101110, 101160, 101180, 101210, 101190, 
    101240, 101230, 101230, 101250, 101250, 101260, 101270, 101260, 101230, 
    101220, 101190, 101180, 101170, 101160, 101170, 101170, 101170, 101200, 
    101190, 101170, 101150, 101160, 101160, 101140, 101210, 101240, 101260, 
    101290, 101290, 101310, 101310, 101330, 101350, 101350, 101340, 101340, 
    101330, 101320, 101290, 101250, 101230, 101210, 101210, 101210, 101260, 
    101240, 101210, 101180, 101130, 101130, 101100, 101100, 101150, 101110, 
    101120, 101120, 101130, 101120, 101120, 101100, 101060, 101080, 100990, 
    100990, 100900, 100910, 100880, 100820, 100780, 100690, 100710, 100620, 
    100480, 100380, 100390, 100370, 100260, 100120, 100050, 100010, 99920, 
    99910, 99900, 99880, 99820, 99740, 99690, 99660, 99640, 99640, 99620, 
    99560, 99490, 99480, 99520, 99600, 99650, 99650, 99710, 99780, 99800, 
    99840, 99910, 99960, 100000, 100010, 100010, 100020, 99980, 99940, 99910, 
    99930, 99940, 99930, 99910, 99910, 99980, 100020, 100030, 100050, 100050, 
    100100, 100140, 100140, 100120, 100130, 100200, 100250, 100290, 100340, 
    100330, 100330, 100380, 100440, 100540, 100610, 100660, 100720, 100780, 
    100790, 100840, 100870, 100930, 100940, 100990, 101010, 101040, 101080, 
    101080, 101090, 101100, 101130, 101160, 101170, 101060, 100970, 101050, 
    101060, 101240, 101260, 101300, 101340, 101360, 101380, 101400, 101440, 
    101430, 101450, 101430, 101330, 101400, 101440, 101520, 101490, 101490, 
    101520, 101530, 101550, 101560, 101740, 101760, 101670, 101640, 101630, 
    101630, 101670, 101600, 101630, 101680, 101680, 101700, 101690, 101670, 
    101620, 101600, 101570, 101550, 101530, 101510, 101460, 101460, 101460, 
    101450, 101430, 101400, 101360, 101330, 101310, 101290, 101280, 101230, 
    101220, 101180, 101140, 101110, 101090, 101070, 101040, 101000, 100970, 
    100940, 100890, 100830, 100790, 100780, 100690, 100660, 100620, 100580, 
    100430, 100340, 100320, 100270, 100220, 100190, 100100, 100030, 99900, 
    99850, 99790, 99740, 99630, 99590, 99650, 99640, 99630, 99610, 99610, 
    99600, 99590, 99600, 99630, 99700, 99670, 99730, 99760, 99820, 99850, 
    99910, 99970, 100020, 100040, 100100, 100160, 100230, 100290, 100330, 
    100380, 100430, 100480, 100560, 100620, 100680, 100710, 100760, 100820, 
    100900, 100950, 100990, 101040, 101100, 101170, 101220, 101280, 101300, 
    101340, 101380, 101450, 101500, 101550, 101600, 101640, 101690, 101740, 
    101800, 101830, 101870, 101900, 101930, 101940, 101980, 102020, 102050, 
    102060, 102080, 102100, 102110, 102110, 102130, 102120, 102100, 102100, 
    102090, 102070, 102040, 102010, 101960, 101950, 101950, 101910, 101860, 
    101820, 101770, 101720, 101660, 101590, 101510, 101440, 101420, 101380, 
    101380, 101340, 101310, 101290, 101290, 101290, 101250, 101220, 101190, 
    101180, 101150, 101130, 101130, 101120, 101090, 101070, 101050, 101020, 
    100980, 100950, 100910, 100870, 100810, 100770, 100730, 100690, 100630, 
    100590, 100560, 100520, 100470, 100440, 100420, 100400, 100400, 100400, 
    100400, 100400, 100400, 100390, 100390, 100370, 100360, 100360, 100360, 
    100340, 100330, 100310, 100300, 100320, 100310, 100310, 100300, 100290, 
    100280, 100260, 100250, 100220, 100210, 100190, 100200, 100230, 100240, 
    100260, 100300, 100300, 100280, 100260, 100290, 100280, 100310, 100340, 
    100360, 100350, 100370, 100390, 100370, 100360, 100380, 100350, 100380, 
    100390, 100430, 100430, 100470, 100490, 100510, 100530, 100550, 100570, 
    100570, 100560, 100590, 100580, 100590, 100590, 100590, 100600, 100590, 
    100610, 100590, 100590, 100580, 100560, 100550, 100550, 100550, 100540, 
    100550, 100560, 100560, 100560, 100580, 100590, 100590, 100590, 100600, 
    100600, 100610, 100620, 100630, 100650, 100650, 100660, 100670, 100680, 
    100690, 100710, 100720, 100730, 100760, 100780, 100820, 100840, 100850, 
    100850, 100860, 100870, 100880, 100890, 100890, 100910, 100920, 100920, 
    100940, 100960, 100960, 100970, 100980, 101000, 101020, 101020, 101050, 
    101070, 101070, 101090, 101120, 101150, 101160, 101170, 101180, 101200, 
    101190, 101190, 101180, 101200, 101190, 101180, 101180, 101160, 101130, 
    101090, 101080, 101120, 101100, 101090, 101030, 101060, 101060, 101080, 
    101120, 101090, 101160, 101180, 101110, 101100, 101090, 101090, 101100, 
    101100, 101090, 101070, 101070, 101070, 101090, 101140, 101190, 101190, 
    101220, 101220, 101260, 101270, 101220, 101240, 101230, 101300, 101330, 
    101340, 101350, 101340, 101320, 101320, 101320, 101290, 101270, 101260, 
    101260, 101250, 101220, 101210, 101200, 101160, 101170, 101140, 101110, 
    101080, 101050, 101030, 101040, 101050, 101030, 101020, 100990, 100970, 
    100920, 100880, 100850, 100840, 100790, 100780, 100740, 100750, 100710, 
    100680, 100600, 100540, 100490, 100480, 100440, 100410, 100350, 100310, 
    100300, 100260, 100270, 100250, 100230, 100200, 100190, 100200, 100210, 
    100240, 100230, 100220, 100260, 100360, 100410, 100450, 100510, 100560, 
    100600, 100650, 100730, 100800, 100870, 100950, 101010, 101040, 101120, 
    101160, 101200, 101270, 101290, 101330, 101370, 101410, 101430, 101470, 
    101500, 101510, 101530, 101540, 101550, 101550, 101570, 101570, 101560, 
    101570, 101580, 101600, 101610, 101630, 101640, 101630, 101630, 101640, 
    101640, 101660, 101660, 101670, 101680, 101700, 101710, 101720, 101720, 
    101730, 101720, 101720, 101720, 101720, 101710, 101700, 101670, 101680, 
    101670, 101690, 101670, 101680, 101670, 101640, 101650, 101640, 101610, 
    101550, 101530, 101470, 101420, 101380, 101350, 101320, 101300, 101290, 
    101270, 101220, 101170, 101180, 101190, 101190, 101210, 101220, 101220, 
    101170, 101140, 101110, 101100, 101090, 101110, 101130, 101140, 101130, 
    101100, 101120, 101140, 101140, 101150, 101180, 101180, 101190, 101230, 
    101250, 101300, 101330, 101360, 101390, 101420, 101440, 101440, 101480, 
    101490, 101500, 101500, 101500, 101530, 101530, 101530, 101530, 101490, 
    101500, 101520, 101500, 101480, 101450, 101420, 101410, 101400, 101390, 
    101400, 101410, 101430, 101460, 101490, 101540, 101670, 101760, 101830, 
    101900, 101980, 102130, 102240, 102280, 102420, 102540, 102630, 102670, 
    102750, 102850, 102900, 102960, 103020, 103090, 103140, 103200, 103230, 
    103220, 103250, 103270, 103280, 103270, 103240, 103220, 103210, 103190, 
    103160, 103110, 103110, 103090, 103030, 102980, 102940, 102910, 102880, 
    102830, 102790, 102730, 102650, 102600, 102550, 102490, 102400, 102350, 
    102290, 102220, 102180, 102150, 102130, 102150, 102190, 102230, 102240, 
    102310, 102270, 102340, 102370, 102400, 102390, 102390, 102420, 102410, 
    102410, 102320, 102280, 102260, 102230, 102180, 102120, 102050, 102030, 
    102020, 102000, 101990, 101970, 101960, 101960, 101940, 101910, 101860, 
    101880, 101870, 101840, 101810, 101800, 101770, 101760, 101760, 101780, 
    101780, 101730, 101710, 101710, 101710, 101710, 101710, 101690, 101690, 
    101680, 101670, 101680, 101660, 101640, 101610, 101620, 101600, 101600, 
    101590, 101610, 101620, 101630, 101650, 101680, 101670, 101670, 101660, 
    101650, 101620, 101580, 101570, 101540, 101530, 101500, 101440, 101400, 
    101370, 101280, 101190, 101170, 101190, 101180, 101170, 101120, 101070, 
    101090, 101100, 101080, 101050, 101010, 101050, 101040, 101030, 101000, 
    100970, 100950, 100940, 100870, 100920, 100880, 100850, 100860, 100830, 
    100800, 100730, 100670, 100630, 100590, 100550, 100490, 100440, 100410, 
    100390, 100350, 100310, 100250, 100180, 100150, 100080, 100020, 99980, 
    99910, 99890, 99850, 99800, 99750, 99720, 99690, 99670, 99650, 99600, 
    99590, 99680, 99730, 99670, 99790, 99840, 99830, 99770, 99810, 99850, 
    99830, 99850, 99900, 99950, 100010, 100030, 100040, 100180, 100240, 
    100270, 100290, 100330, 100340, 100370, 100420, 100500, 100570, 100640, 
    100710, 100740, 100800, 100830, 100880, 100950, 100970, 101000, 101040, 
    101050, 101070, 101110, 101120, 101130, 101140, 101140, 101150, 101180, 
    101190, 101200, 101220, 101250, 101250, 101270, 101270, 101260, 101250, 
    101270, 101250, 101230, 101220, 101210, 101200, 101190, 101190, 101160, 
    101150, 101120, 101100, 101080, 101040, 101020, 101010, 100970, 100980, 
    100970, 100930, 100910, 100890, 100850, 100800, 100740, 100700, 100630, 
    100550, 100480, 100400, 100320, 100240, 100170, 100080, 99980, 99900, 
    99810, 99730, 99670, 99570, 99560, 99550, 99510, 99490, 99450, 99390, 
    99430, 99420, 99430, 99450, 99440, 99450, 99450, 99450, 99470, 99490, 
    99530, 99480, 99490, 99530, 99520, 99500, 99450, 99420, 99430, 99420, 
    99440, 99430, 99440, 99430, 99420, 99450, 99490, 99490, 99530, 99560, 
    99650, 99780, 99870, 99970, 100010, 100120, 100240, 100340, 100430, 
    100540, 100580, 100640, 100710, 100790, 100860, 100920, 100960, 100980, 
    100970, 100950, 100900, 100840, 100780, 100720, 100620, 100590, 100570, 
    100550, 100570, 100580, 100620, 100630, 100660, 100650, 100650, 100660, 
    100640, 100640, 100640, 100640, 100670, 100660, 100650, 100650, 100700, 
    100670, 100670, 100670, 100610, 100630, 100650, 100650, 100720, 100730, 
    100760, 100760, 100780, 100760, 100730, 100700, 100690, 100700, 100740, 
    100770, 100790, 100800, 100810, 100820, 100830, 100840, 100850, 100850, 
    100830, 100830, 100860, 100830, 100830, 100830, 100780, 100720, 100670, 
    100650, 100610, 100560, 100520, 100490, 100530, 100520, 100510, 100500, 
    100510, 100510, 100470, 100470, 100470, 100480, 100470, 100480, 100490, 
    100500, 100520, 100530, 100530, 100550, 100600, 100580, 100600, 100600, 
    100570, 100590, 100630, 100650, 100680, 100690, 100730, 100730, 100760, 
    100740, 100760, 100790, 100830, 100870, 100920, _, 101400, 101430, 
    101450, 101470, 101500, 101520, 101530, 101550, 101580, 101600, 101610, 
    101650, 101690, 101680, 101680, 101690, 101700, 101670, 101700, 101700, 
    101710, 101740, 101740, 101780, 101770, 101770, 101750, 101740, 101710, 
    101690, 101680, 101640, 101620, 101590, 101540, 101540, 101490, 101390, 
    101200, 101130, 101070, 101030, 101060, 101090, 101090, 101100, 101160, 
    101220, 101270, 101310, 101330, 101380, 101410, 101470, 101530, 101590, 
    101670, 101730, 101790, 101870, 101910, 101970, 101990, 102060, 102080, 
    102120, 102170, 102200, 102240, 102270, 102300, 102330, 102360, 102370, 
    102360, 102340, 102330, 102320, 102320, 102310, 102270, 102260, 102220, 
    102200, 102160, 102140, 102100, 102050, 102000, 101950, 101900, 101890, 
    101840, 101780, 101730, 101690, 101650, 101590, 101520, 101400, 101290, 
    101190, 101100, 101010, 100920, 100810, 100710, 100590, 100480, 100380, 
    100250, 100140, 100070, 99980, 99930, 99890, 99840, 99810, 99770, 99750, 
    99730, 99680, 99610, 99540, 99480, 99400, 99300, 99210, 99120, 99000, 
    98910, 98830, 98770, 98710, 98670, 98650, 98630, 98630, 98640, 98650, 
    98630, 98630, 98630, 98640, 98650, 98650, 98670, 98660, 98700, 98770, 
    98850, 98940, 99030, 99100, 99150, 99200, 99240, 99220, 99180, 99200, 
    99220, 99220, 99170, 99170, 99100, 99060, 98970, 98910, 98840, 98700, 
    98570, 98510, 98440, 98400, 98290, 98290, 98250, 98250, 98280, 98280, 
    98320, 98360, 98420, 98470, 98540, 98620, 98680, 98790, 98820, 98880, 
    98940, 99010, 99060, 99090, 99110, 99120, 99090, 99110, 99150, 99120, 
    99080, 99070, 99030, 99010, 98980, 98940, 98840, 98780, 98720, 98650, 
    98590, 98560, 98450, 98440, 98400, 98370, 98390, 98370, 98340, 98350, 
    98330, 98320, 98350, 98380, 98420, 98470, 98530, 98590, 98650, 98670, 
    98690, 98730, 98760, 98780, 98830, 98840, 98870, 98880, 98920, 98960, 
    98970, 99010, 99040, 99060, 99090, 99130, 99150, 99160, 99230, 99310, 
    99330, 99390, 99450, 99530, 99610, 99650, 99720, 99770, 99830, 99900, 
    99980, 100040, 100090, 100140, 100190, 100190, 100220, 100230, 100220, 
    100240, 100230, 100250, 100240, 100260, 100230, 100240, 100250, 100250, 
    100230, 100250, 100270, 100310, 100350, 100390, 100430, 100460, 100510, 
    100550, 100580, 100580, 100560, 100550, 100510, 100450, 100430, 100410, 
    100390, 100370, 100370, 100330, 100310, 100280, 100260, 100210, 100200, 
    100190, 100170, 100140, 100140, 100150, 100130, 100100, 100120, 100080, 
    100080, 100010, 100050, 100000, 100040, 100090, 100080, 100060, 99970, 
    99870, 99910, 99920, 99910, 99910, 99890, 99880, 99840, 99880, 99890, 
    99910, 99940, 99940, 99940, 99960, 99990, 99990, 100040, 100070, 100110, 
    100130, 100170, 100200, 100260, 100330, 100390, 100460, 100500, 100490, 
    100560, 100530, 100590, 100590, 100650, 100710, 100680, 100710, 100730, 
    100710, 100710, 100720, 100680, 100650, 100610, 100560, 100530, 100520, 
    100490, 100480, 100440, 100430, 100430, 100420, 100400, 100390, 100370, 
    100350, 100350, 100360, 100350, 100370, 100360, 100360, 100350, 100350, 
    100350, 100370, 100370, 100380, 100380, 100400, 100420, 100430, 100450, 
    100430, 100420, 100440, 100430, 100440, 100420, 100410, 100380, 100430, 
    100480, 100470, 100480, 100500, 100470, 100460, 100530, 100550, 100560, 
    100570, 100540, 100510, 100440, 100380, 100400, 100470, 100440, 100430, 
    100480, 100500, 100540, 100590, 100620, 100650, 100670, 100720, 100740, 
    100760, 100780, 100780, 100790, 100780, 100760, 100740, 100740, 100770, 
    100780, 100770, 100760, 100750, 100730, 100710, 100700, 100690, 100670, 
    100630, 100620, 100610, 100610, 100600, 100570, 100550, 100540, 100510, 
    100500, 100480, 100460, 100440, 100420, 100410, 100400, 100390, 100370, 
    100360, 100330, 100300, 100310, 100310, 100290, 100290, 100280, 100270, 
    100280, 100280, 100280, 100280, 100290, 100320, 100330, 100360, 100380, 
    100410, 100420, 100460, 100490, 100520, 100540, 100570, 100560, 100550, 
    100560, 100610, 100620, 100640, 100670, 100710, 100740, 100760, 100780, 
    100820, 100810, 100780, 100780, 100800, 100790, 100800, 100820, 100830, 
    100840, 100860, 100870, 100910, 100890, 100940, 100970, 100980, 101020, 
    101050, 101060, 101070, 101130, 101160, 101190, 101190, 101190, 101180, 
    101150, 101120, 101080, 101090, 101040, 100990, 101020, 101000, 101000, 
    100980, 100950, 100930, 100910, 100890, 100880, 100870, 100870, 100900, 
    100930, 101000, 101020, 101040, 101030, 101030, 101030, 101040, 101080, 
    101120, 101120, 101120, 101150, 101180, 101270, _, _, _, _, _, _, _, _, 
    _, 101440, 101480, 101520, 101570, 101630, 101650, 101660, 101700, 
    101680, 101720, 101800, 101830, 101900, 101990, 102070, 102120, 102190, 
    102230, 102290, 102320, 102340, 102350, 102360, 102380, _, 102530, 
    102570, 102650, 102690, 102760, 102740, 102790, 102820, 102820, 102830, 
    102880, 102910, 102970, 102970, 103000, 103010, 103030, 103050, 103030, 
    103040, 103020, 103050, 103070, 103120, 103150, 103170, 103170, 103160, 
    103170, 103180, 103190, 103200, 103240, 103280, 103310, 103350, 103360, 
    103390, 103390, 103410, 103440, 103490, 103530, 103580, 103610, 103640, 
    103680, 103710, 103770, 103810, 103830, 103830, 103830, 103830, 103860, 
    103850, 103850, 103860, 103860, 103800, 103770, 103840, 103850, 103810, 
    103790, 103750, 103690, 103660, 103500, 103520, 103480, 103500, 103510, 
    103520, 103510, 103490, 103490, 103500, 103510, 103520, 103530, 103540, 
    103540, 103540, 103530, 103560, 103530, 103510, 103500, 103520, 103550, 
    103560, 103550, 103580, 103600, 103610, 103640, 103630, 103640, 103680, 
    103690, 103720, 103710, 103730, 103720, 103710, 103660, 103660, 103660, 
    103670, 103660, 103640, 103620, 103620, 103600, 103590, 103600, 103610, 
    103610, 103630, 103630, 103640, 103630, 103630, 103650, 103660, 103680, 
    103700, 103690, 103690, 103720, 103750, 103760, 103810, 103830, 103880, 
    103880, 103870, 103900, 103890, 103910, 103900, 103910, _, 103960, 
    103980, 104010, 104000, 103980, 103970, 103950, 103910, 103870, 103840, 
    103810, 103780, 103750, 103710, 103660, 103630, 103590, 103540, 103500, 
    103460, 103430, 103380, 103320, 103250, 103220, 103180, 103160, 103100, 
    103050, 103000, 102940, 102930, 102900, 102870, 102840, 102820, 102830, 
    102780, 102770, 102730, 102700, 102650, 102640, 102610, 102570, 102560, 
    102540, 102580, 102580, 102560, 102570, 102570, 102560, 102530, 102510, 
    102480, 102470, 102460, 102450, 102440, 102470, 102470, 102470, 102440, 
    102410, 102380, 102340, 102340, 102340, 102340, 102340, 102340, 102340, 
    102350, 102340, 102300, 102310, 102280, 102260, 102220, 102210, 102190, 
    102180, 102160, 102170, 102150, 102100, 102080, 102050, 102020, 101990, 
    101990, 101980, 101930, 101910, 101910, 101910, 101900, 101900, 101850, 
    101800, 101730, 101660, 101600, 101550, 101520, 101470, 101420, 101390, 
    101370, 101360, 101320, 101310, 101280, 101250, 101230, 101240, 101240, 
    101260, 101290, 101270, 101250, 101260, 101290, 101270, 101250, 101240, 
    101210, 101200, 101160, 101150, 101150, 101120, 101070, 101050, 100980, 
    100940, 100900, 100880, 100870, 100850, 100870, 100860, 100870, 100930, 
    100960, 101030, 101020, 101040, 101040, 101090, 101120, 101160, 101180, 
    101200, 101240, 101260, 101290, 101320, 101350, 101350, 101390, 101340, 
    101410, 101430, 101440, 101500, 101550, 101620, 101680, 101680, 101710, 
    101750, 101790, 101830, 101860, 101940, 102010, 102090, 102160, 102250, 
    102250, 102310, 102350, 102420, 102470, 102520, 102590, 102660, 102760, 
    102840, 102900, 102970, 103020, 103060, 103090, 103130, 103180, 103240, 
    103280, 103340, 103370, 103390, 103440, 103470, 103470, 103470, 103430, 
    103360, 103270, 103260, 103200, 103110, 103030, 102930, 102790, 102710, 
    102560, 102380, 102260, 102200, 102170, 102170, 102180, 102200, 102220, 
    102210, 102220, 102200, 102210, 102220, 102190, 102170, 102220, 102270, 
    102260, 102280, 102340, 102390, 102430, 102490, 102560, 102590, 102630, 
    102670, 102650, 102680, 102700, 102750, 102740, 102750, 102790, 102830, 
    102830, 102840, 102880, 102880, 102880, 102860, 102900, 102880, 102960, 
    103000, 103080, 103120, 103180, 103220, 103280, 103300, 103310, 103300, 
    103320, 103350, 103350, 103360, 103370, 103370, 103370, 103370, 103340, 
    103290, 103240, 103250, 103210, 103150, 103090, 103060, 103020, 102990, 
    102960, 102930, 102860, 102790, 102730, 102610, 102560, 102540, 102480, 
    102420, 102370, 102350, 102280, 102240, 102180, 102160, 102130, 102100, 
    102070, 102030, 102010, 101970, 101980, 101980, 101960, 101920, 101890, 
    101890, 101840, 101800, 101770, 101770, 101750, 101750, 101770, 101750, 
    101750, 101740, 101750, 101780, 101790, 101820, 101830, 101860, 101860, 
    101900, 101940, 101980, 101980, 102000, 102020, 102020, 101990, 101940, 
    101920, 101870, 101810, 101770, 101730, 101650, 101530, 101420, 101310, 
    101300, 101260, 101180, 101110, 101070, 101010, 100920, 100820, 100740, 
    100710, 100630, 100510, 100440, 100380, 100310, 100240, 100180, 100150, 
    100140, 100120, 100110, 100100, 100110, 100110, 100110, 100080, 100050, 
    100000, 100020, 100050, 100090, 100160, 100180, 100300, 100550, 100670, 
    100830, 100950, 101110, 101220, 101310, 101470, 101560, 101670, 101750, 
    101850, 101900, 101930, 101970, 101990, 102030, 102040, 102080, 102140, 
    102190, 102250, 102320, 102370, 102420, 102500, 102550, 102630, 102700, 
    102770, 102820, 102870, 102930, 102970, 103030, 103070, 103090, 103110, 
    103100, 103120, 103100, 103090, 103030, 102930, 102860, 102780, 102680, 
    102560, 102450, 102310, 102140, 101950, 101720, 101570, 101400, 101230, 
    101030, 101020, 100980, 100940, 100970, 101050, 101110, 101100, _, 
    101280, 101420, 101580, 101710, 101890, 102030, 102160, 102290, 102350, 
    102410, 102540, 102590, 102650, 102710, 102760, 102780, 102810, 102830, 
    102810, 102800, 102800, 102830, 102840, 102850, 102870, 102910, 102910, 
    102930, 102980, 103010, 103030, 103060, 103050, 103080, 103110, 103070, 
    102950, 102940, 102790, 102710, 102600, 102440, 102290, 102110, 101790, 
    101490, 101250, 101050, 100860, 100610, 100230, 100050, 99980, 99920, 
    99870, 99820, 99730, 99670, 99600, 99510, 99460, 99430, 99450, 99400, 
    99350, 99260, 99180, 99140, 99130, 99160, 99160, 99180, 99260, 99600, 
    99880, 100120, 100410, 100610, 100810, 101030, 101150, 101200, 101260, 
    101590, 101780, 101720, 101880, 102020, 102120, 102160, 102210, 102210, 
    102200, 102240, 102220, 102200, 102170, 102110, 102050, 102000, 101930, 
    101860, 101760, 101630, 101510, 101360, 101210, 101030, 100880, 100700, 
    100560, 100470, 100390, 100320, 100270, 100150, 100070, 99970, 99870, 
    99780, 99680, 99570, 99460, 99380, 99310, 99270, 99230, 99210, 99180, 
    99150, 99150, 99130, 99180, 99190, 99200, 99200, 99260, 99310, 99340, 
    99360, 99360, 99360, 99350, 99320, 99330, 99310, 99300, 99310, 99350, 
    99350, 99380, 99430, 99400, 99400, 99430, 99390, 99360, 99320, 99250, 
    99190, 99170, 99190, 99190, 99140, 99070, 99000, 98910, 98830, 98610, 
    98380, 98210, 97700, 97580, 97530, 97450, 97340, 97350, 97380, 97610, 
    97870, 98250, 98440, 98590, 98770, 98890, 98990, 99060, 99090, 99100, 
    99140, 99190, 99210, 99240, 99280, 99320, 99320, 99400, 99460, 99510, 
    99540, 99530, 99560, 99600, 99670, 99740, 99780, 99830, 99890, 99950, 
    100000, 100070, 100130, 100200, 100250, 100290, 100390, 100430, 100480, 
    100550, 100630, 100630, 100670, 100680, 100670, 100500, 100470, 100490, 
    100510, 100500, 100520, 100540, 100580, 100600, 100670, 100710, 100720, 
    100690, 100660, 100680, 100670, 100680, 100660, 100700, 100650, 100690, 
    100670, 100670, 100650, 100650, 100610, 100600, 100590, 100540, 100730, 
    100770, 100800, 100860, 100910, 100960, 100990, 101030, 101060, 101050, 
    101050, 101070, 101060, 101070, 101050, 101070, 101060, 101100, 101090, 
    101090, 101060, 100990, 100970, 100980, 100990, 100990, 101030, 101010, 
    101010, 101010, 101020, 101020, 101030, 101060, 101060, 101060, 101080, 
    101100, 101070, 101040, 101020, 101050, 100980, 100990, 101010, 101010, 
    100960, 100960, 100900, 100870, 100850, 100850, 100810, 100830, 100810, 
    100770, 100770, 100790, 100800, 100780, 100750, 100770, 100720, 100690, 
    100700, 100650, 100620, 100610, 100600, 100590, 100570, 100580, 100620, 
    100600, 100640, 100620, 100620, 100620, 100600, 100560, 100570, 100550, 
    100500, 100460, 100410, 100370, 100330, 100370, 100360, 100380, 100340, 
    100260, 100270, 100260, 100180, 100150, 100140, 100080, 99990, 99900, 
    99840, 99880, 99820, 99790, 99730, 99770, 99760, 99770, 99800, 99770, 
    99810, 99850, 99940, 99940, 99970, 100010, 100090, 100150, 100160, 
    100200, 100210, 100240, 100280, 100340, 100330, 100310, 100350, 100370, 
    100410, _, 100480, 100510, 100530, 100560, 100610, 100650, 100690, 
    100720, 100740, 100730, 100770, 100780, 100850, 100860, 100920, 100970, 
    101030, 101080, 101150, 101210, 101240, 101280, 101340, 101380, 101440, 
    101490, 101520, 101550, 101610, 101670, 101730, 101780, 101790, 101820, 
    101850, 101840, 101850, 101840, 101790, 101770, 101770, 101740, 101710, 
    101660, 101620, 101550, 101490, 101430, 101330, 101190, 101060, 100970, 
    100880, 100780, 100670, 100610, 100520, 100390, 100250, 100180, 100100, 
    100030, 99950, 99860, 99800, 99680, 99610, 99520, 99450, 99400, 99350, 
    99270, 99190, 99130, 99080, 99070, 99010, 98980, 98970, 99010, 99080, 
    99140, 99190, 99240, 99260, 99300, 99320, 99320, 99340, 99360, 99360, 
    99350, 99340, 99340, 99390, 99430, 99430, 99440, 99420, 99440, 99460, 
    99500, 99570, 99660, 99710, 99760, 99840, 99930, 99990, 100050, 100090, 
    100150, 100220, 100280, 100350, 100410, 100460, 100530, 100570, 100630, 
    100660, 100700, 100730, 100810, 100880, 100920, 100970, 101010, 101020, 
    101060, 101060, 101070, 101090, 101070, 101030, 100990, 100960, 100910, 
    100930, 100920, 100890, 100860, 100830, 100770, 100760, 100700, 100650, 
    100630, 100560, 100500, 100460, 100440, 100310, 100180, 100100, 99980, 
    99900, 99820, 99740, 99700, 99650, 99620, 99570, 99470, 99320, 99200, 
    99040, 98890, 98810, 98650, 98600, 98590, 98650, 98700, 98770, 98840, 
    98920, 98980, 99020, 99040, 99120, 99170, 99230, 99390, 99520, 99690, 
    99870, 100000, 100090, 100110, 100170, 100190, 100250, 100290, 100340, 
    100370, 100400, 100440, 100460, 100440, 100410, 100430, 100460, 100440, 
    100480, 100500, 100530, 100570, 100560, 100590, 100590, 100610, 100470, 
    100560, 100580, _, 100700, 100790, 100760, 100750, 100800, 100850, 
    100900, 100960, 101010, 101000, 101050, 101090, 101140, 101190, 101260, 
    101300, 101350, 101420, 101460, 101510, 101580, 101630, 101670, 101710, 
    101740, 101780, 101810, 101840, 101870, 101920, 101990, 102020, 102050, 
    102070, 102080, 102100, 102120, 102140, 102160, 102160, 102160, 102150, 
    102150, 102160, 102160, 102170, 102180, 102170, 102160, 102110, 102110, 
    102080, 102090, 102090, 102090, 102090, 102080, 102070, 102030, 101980, 
    101960, 101950, 101930, 101900, 101870, 101810, 101770, 101730, 101700, 
    101660, 101610, 101560, 101510, 101430, 101340, 101280, 101190, 101200, 
    101090, 101090, 101060, 101020, 100960, 100900, 100870, 100770, 100730, 
    100710, 100600, 100630, 100590, 100560, 100510, 100500, 100460, 100530, 
    100530, 100560, 100580, 100590, 100570, 100470, 100450, 100340, 100350, 
    100330, 100300, 100290, 100310, 100300, 100410, 100360, 100390, 100460, 
    100510, 100470, 100480, 100520, 100480, 100540, 100600, 100590, 100580, 
    100600, 100540, 100560, 100510, 100410, 100420, 100500, 100610, 100650, 
    100750, 100850, 100990, 101010, 101140, 101220, 101350, 101400, 101460, 
    101530, 101560, 101610, 101620, 101630, 101640, 101660, 101680, 101680, 
    101690, 101710, 101740, 101720, 101710, 101710, 101690, 101700, 101680, 
    101630, 101580, 101590, 101550, 101440, 101410, 101320, 101260, 101190, 
    101080, 100970, 100900, 100790, 100690, 100610, 100570, 100450, 100380, 
    100270, 100180, 100090, 100040, 99940, 99920, 99900, 99870, 99980, 
    100000, 100090, 100150, 100170, 100210, 100340, 100400, 100440, 100620, 
    100610, 100620, 100640, 100690, 100770, 100790, 100810, 100830, 100890, 
    100940, 100950, 100980, 101050, 101050, 101070, 101120, 101130, 101130, 
    101080, 101100, 101090, 101120, 101090, 101080, 101090, 101140, 101140, 
    101110, 101110, 101140, 101130, 101110, 101090, 101120, 101120, 101130, 
    101120, 101160, 101150, 101180, 101260, 101380, 101440, 101590, 101600, 
    101690, 101710, 101860, 101880, 101870, 101870, 102060, 102190, 102210, 
    102270, 102290, 102300, 102290, 102260, 102270, 102280, 102270, 102220, 
    102160, 102200, 102170, 102150, 102130, 102050, 102030, 101980, 101970, 
    101920, 101860, 101790, 101730, 101650, 101570, 101500, 101430, 101380, 
    101380, 101400, 101430, 101440, 101410, 101460, 101460, 101440, 101420, 
    101390, 101360, 101330, 101280, 101250, 101210, 101180, 101160, 101140, 
    101120, 101100, 101040, 101010, 101010, 101030, 101030, 101020, 101010, 
    101010, 101010, 101040, 101030, 101010, 101000, 100990, 100970, 100960, 
    100980, 100970, 100970, 100920, 100910, 100900, 100960, 100970, 100950, 
    100940, 100910, 100900, 100880, 100870, 100850, 100810, 100790, 100750, 
    100750, 100740, 100750, 100750, 100730, 100720, 100740, 100740, 100740, 
    100740, 100730, 100740, 100760, 100770, 100760, 100760, 100740, 100730, 
    100710, 100730, 100690, 100690, 100680, 100680, 100680, 100680, 100690, 
    100660, 100640, 100650, 100630, 100620, 100630, 100640, 100660, 100640, 
    100650, 100670, 100690, 100710, 100720, 100740, 100740, 100750, 100780, 
    100790, 100790, 100800, 100840, 100840, 100850, 100850, 100850, 100860, 
    100840, 100860, 100840, 100830, 100820, 100830, 100850, 100880, 100890, 
    100890, 100880, 100890, 100880, 100860, 100850, 100850, 100840, 100820, 
    100790, 100770, 100750, 100720, 100720, 100670, 100660, 100610, 100550, 
    100510, 100460, 100430, 100380, 100380, 100340, 100470, 100290, 100360, 
    100430, 100410, 100380, 100350, 100320, 100300, 100300, 100220, 100180, 
    100140, 100110, 100150, 100160, 100210, 100100, 100130, 100160, 100200, 
    100320, 100390, 100440, 100440, 100450, 100450, 100480, 100490, 100500, 
    100510, 100550, 100560, 100550, 100550, 100540, 100530, 100440, 100460, 
    100470, 100530, 100490, 100480, 100510, 100530, 100520, 100520, 100520, 
    100510, 100490, 100480, 100470, 100470, 100460, 100460, 100450, 100420, 
    100440, 100440, 100440, 100400, 100390, 100380, 100380, 100340, 100330, 
    100380, 100380, 100400, 100410, 100390, 100380, 100480, 100410, 100420, 
    100420, 100400, 100400, 100370, 100360, 100360, 100340, 100290, 100240, 
    100210, 100110, 100200, 100280, 100260, 100240, 100230, 100250, 100180, 
    100260, 100220, 100150, 100160, 100190, 100180, 100140, 100140, 100120, 
    100130, 100130, 100160, 100190, 100210, 100210, 100210, 100220, 100240, 
    100260, 100270, 100320, 100320, 100320, 100360, 100370, 100400, 100350, 
    100340, 100350, 100380, 100380, 100400, 100410, 100440, 100480, 100500, 
    100520, 100560, 100590, 100580, 100580, 100570, 100650, 100720, 100760, 
    100810, 100850, 100910, 100950, 101010, 101050, 101060, 101100, 101140, 
    101180, 101220, 101260, 101290, 101340, 101370, 101390, 101430, 101470, 
    101500, 101520, 101540, 101570, 101600, 101620, 101630, 101640, 101660, 
    101690, 101700, 101700, 101690, 101690, 101680, 101700, 101690, 101670, 
    101670, 101630, 101620, 101620, 101610, 101570, 101550, 101540, 101550, 
    101520, 101520, 101490, 101480, 101480, 101480, 101470, 101470, 101480, 
    101480, 101480, 101440, 101410, 101440, 101410, 101400, 101380, 101370, 
    101370, 101380, 101370, 101370, 101340, 101330, 101320, 101330, 101330, 
    101310, 101300, 101310, 101340, 101330, 101320, 101310, 101280, 101280, 
    101290, 101280, 101290, 101300, 101260, 101280, 101260, 101240, 101240, 
    101190, 101160, 101180, 101180, 101140, 101120, 101110, 101090, 101100, 
    101070, 101070, 101070, 101060, 101050, 101050, 101050, 101030, 101010, 
    100960, 100960, 100970, 100980, 101010, 101010, 101010, 101030, 101020, 
    101030, 101070, 101060, 101070, 101110, 101130, 101150, 101170, 101170, 
    101140, 101080, 100970, 100920, 100810, 100760, 100730, 100640, 100560, 
    100650, 100690, 100750, 100780, 100800, 100880, 100970, 101030, 101120, 
    101230, 101290, 101410, 101440, 101460, 101530, 101540, 101540, 101540, 
    101570, 101570, 101560, 101520, 101540, 101540, 101540, 101540, 101620, 
    101660, 101750, 101870, 101890, 101930, 101990, 102030, 102070, 102100, 
    102130, 102140, 102170, 102190, 102210, 102230, 102260, 102270, 102300, 
    102310, 102320, 102300, 102290, 102250, 102230, 102220, 102170, 102160, 
    102080, 102040, 101990, 101940, 101920, 101960, 101960, 101920, 101940, 
    101940, 101950, 101930, 101920, 101900, 101890, 101870, 101860, 101850, 
    101840, 101810, 101810, 101780, 101760, 101710, 101640, 101610, 101490, 
    101410, 101330, 101300, 101240, 101200, 101140, 101090, 100980, 100920, 
    100830, 100750, 100650, 100550, 100480, 100400, 100360, 100330, 100350, 
    100300, 100270, 100240, 100240, 100250, 100330, 100400, 100470, 100520, 
    100580, 100620, 100650, 100710, 100730, 100790, 100760, 100770, 100850, 
    100940, 101040, 101110, 101190, 101250, 101370, 101440, 101510, 101580, 
    101640, 101730, 101760, 101810, 101830, 101880, 101930, 101960, 101980, 
    102010, 102030, 102010, 102010, 102000, 101990, 101990, 101970, 101960, 
    101990, 101990, 101940, 101910, 101900, 101840, 101830, 101790, 101740, 
    101750, 101740, 101700, 101670, 101660, 101620, 101580, 101530, 101480, 
    101460, 101410, 101370, 101380, 101410, 101460, 101490, 101490, 101630, 
    101740, 101820, 101900, 101930, 101940, 102000, 102090, 102150, 102190, 
    102200, 102210, 102330, 102400, 102490, 102530, 102530, 102620, 102620, 
    102630, 102630, 102610, 102590, 102540, 102480, 102430, 102380, 102240, 
    102190, 102130, 102060, 102000, 101930, 101880, 101860, 101850, 101910, 
    101940, 101980, 102040, 102120, 102170, 102200, 102190, 102210, 102210, 
    102210, 102180, 102130, 102100, 102050, 102000, 101960, 101900, 101840, 
    101790, 101740, 101670, 101610, 101560, 101480, 101430, 101390, 101350, 
    101330, 101330, 101360, 101410, 101440, 101470, 101540, 101500, 101610, 
    101650, 101670, 101720, 101750, 101780, 101790, 101840, 101870, 101890, 
    101930, 101940, 102010, 102060, 102060, 102130, 102140, 102140, 102210, 
    102280, 102280, 102310, 102400, 102390, 102400, 102390, 102390, 102380, 
    102440, 102430, 102360, 102290, 102310, 102340, 102340, 102280, 102270, 
    102230, 102180, 102150, 102090, 102080, 102000, 101970, 101950, 101900, 
    101870, 101830, 101760, 101680, 101620, 101560, 101500, 101410, 101340, 
    101300, 101280, 101270, 101270, 101230, 101270, 101280, 101330, 101310, 
    101300, 101260, 101260, 101240, 101230, 101220, 101210, 101220, 101220, 
    101240, 101190, 101160, 101110, 101090, 101050, 101020, 101060, 101030, 
    101060, 101160, 101190, 101190, 101250, 101320, 101380, 101400, 101410, 
    101490, 101590, 101630, 101670, 101700, 101700, 101700, 101670, 101680, 
    101670, 101630, 101580, 101570, 101510, 101450, 101420, 101400, 101350, 
    101300, 101250, 101200, 101150, 101130, 101100, 101070, 101040, 101040, 
    101040, 101040, 101070, 101120, 101150, 101190, 101240, 101270, 101310, 
    101350, 101400, 101500, 101580, 101650, 101710, 101790, 101880, 101930, 
    102000, 102060, 102090, 102130, 102180, 102220, 102270, 102300, 102340, 
    102370, 102360, 102380, 102380, 102390, 102370, 102360, 102340, 102370, 
    102380, 102420, 102410, 102420, 102430, 102430, 102430, 102400, 102390, 
    102380, 102360, 102370, 102390, 102400, 102380, 102380, 102360, 102340, 
    102320, 102300, 102260, 102230, 102190, 102190, 102180, 102170, 102140, 
    102160, 102130, 102130, 102120, 102130, 102110, 102100, 102110, 102110, 
    102100, 102080, 102080, 102070, 102000, 102030, 102040, 102030, 102020, 
    102010, 102040, 102040, 102060, 102050, _, 102040, 102020, 102010, 
    102000, 101990, 101950, 101930, 101930, 101930, _, 101890, 101850, 
    101840, 101810, 101790, 101770, 101750, 101720, 101720, 101730, 101720, 
    101740, 101720, 101710, 101730, 101720, 101700, 101670, 101670, 101650, 
    101640, 101630, 101580, 101580, _, 101530, 101530, 101510, 101510, 
    101510, 101490, 101450, 101450, 101480, 101540, 101630, 101700, 101760, 
    101790, 101830, 101790, 101820, 101770, 101830, 101800, 101700, 101680, 
    101680, 101700, 101690, 101670, 101590, 101570, 101560, 101520, 101490, 
    _, 101430, 101510, 101540, 101620, 101560, 101590, 101580, 101550, 
    101550, 101600, 101510, 101520, 101640, 101630, 101560, _, 101590, 
    101670, 101720, 101770, 101850, 101920, 102020, 102040, 102060, 102130, 
    102250, 102360, 102410, 102470, 102570, 102630, 102700, 102730, 102760, 
    102780, 102780, 102830, 102870, 102820, 102760, 102720, 102740, 102720, 
    102660, 102650, 102670, 102670, 102700, 102680, 102640, 102670, 102620, 
    102540, 102520, 102500, 102490, 102430, 102440, 102410, 102410, 102460, 
    102440, 102410, 102410, 102410, 102390, 102400, 102390, 102430, 102440, 
    102450, 102470, 102510, 102530, 102580, 102580, 102610, 102630, 102620, 
    102620, 102620, 102630, 102660, 102670, 102700, 102700, 102690, 102710, 
    102700, 102660, 102600, 102590, 102490, 102480, 102460, 102380, 102310, 
    102230, 102150, 102100, 102010, 102040, 101950, 102040, 101990, 101940, 
    101890, 101910, 101890, 101870, 101880, 101810, 101820, 101820, 101850, 
    101900, 101940, 101920, 101920, 101880, 101970, 102040, 102090, 102090, 
    102080, 102070, 102130, 102100, 102060, 102060, 102060, 102040, 102050, 
    102010, 101960, 102030, 102040, 102010, 102100, 102070, 102140, 102200, 
    102250, 102280, 102330, 102400, 102450, 102460, 102490, 102500, 102520, 
    102540, 102540, 102510, 102560, 102570, 102580, 102600, 102600, 102610, 
    102560, 102560, 102530, 102510, 102460, 102480, 102510, 102450, 102350, 
    102350, 102480, 102380, 102460, 102460, 102420, 102420, 102340, 102230, 
    102240, 102230, 102200, 102260, 102210, 102240, 102220, 102180, 102150, 
    102150, 102170, 102210, 102170, 102170, 102160, 102200, 102170, 102170, 
    102120, 102080, 102070, 102030, 101980, 101910, 101870, 101780, 101710, 
    101650, 101600, 101570, 101530, 101480, 101410, 101430, 101420, 101370, 
    101320, 101320, 101310, 101270, 101210, 101200, 101150, 101120, 101080, 
    101050, 101040, 101020, 101010, 100940, 100940, 100930, 100860, 100840, 
    100800, 100760, 100700, 100630, 100570, 100560, 100500, 100450, 100440, 
    100440, 100410, 100370, 100350, 100330, 100330, 100330, 100340, 100360, 
    100390, 100410, 100460, 100500, 100550, 100590, 100660, 100720, 100770, 
    100820, 100890, 100950, 101000, 101060, 101130, 101180, 101230, 101270, 
    101330, 101360, 101400, 101410, 101410, 101400, 101460, 101470, 101510, 
    101550, 101560, 101630, 101610, 101640, 101690, 101730, 101790, 101710, 
    101710, 101740, 101800, 101830, 101840, 101850, 101860, 101880, 101990, 
    102080, 102170, 102250, 102360, 102420, 102540, 102590, 102640, 102700, 
    102760, 102810, 102900, 102960, 103030, 103120, 103180, 103200, 103270, 
    103360, 103410, 103460, 103490, 103510, 103530, 103610, 103680, 103750, 
    103850, 103960, 104020, 104090, 104110, 104200, 104280, 104350, 104410, 
    104470, 104490, 104540, 104570, 104590, 104620, 104710, 104750, 104780, 
    104760, 104820, 104820, 104850, 104890, 104940, 104960, 105010, 104980, 
    105010, 105010, 105010, 105120, 104890, 104920, 104950, 104820, 104860, 
    104970, 105000, 105060, 105140, 105170, 105190, 105200, 105240, 105270, 
    105260, 105280, 105270, 105290, 105340, 105390, 105450, 105520, 105560, 
    105610, 105640, 105650, 105690, 105740, 105750, 105770, 105790, 105780, 
    105810, 105830, 105870, 105870, 105860, 105870, 105860, 105860, 105830, 
    105790, 105760, 105730, 105690, 105640, 105580, 105510, 105460, 105390, 
    105320, 105240, 105160, 105060, 104990, 104930, 104890, 104840, 104830, 
    104750, 104660, 104550, 104580, 104420, 104330, 104190, 104140, 104090, 
    104040, 104080, 104000, 103990, 103930, 103850, 103720, 103660, 103620, 
    103560, 103460, 103330, 103300, 103270, 103230, 103200, 103190, 103190, 
    103170, 103150, 103150, 103140, 103130, 103110, 103140, 103140, 103160, 
    103130, 103140, 103090, 103090, 103110, 103080, 103050, 103030, 103080, 
    103100, 103060, 103070, 103060, 103080, 103080, 103050, 103020, 103000, 
    102960, 102920, 102890, 102880, 102870, 102860, 102840, 102830, 102830, 
    102800, 102800, 102790, 102800, 102800, 102810, 102870, 102890, 102930, 
    102930, 102930, 102950, 102960, 102980, 102990, 102990, 102990, 103000, 
    103010, 103010, 102990, 102970, 102970, 102950, 102930, 102890, 102880, 
    102790, 102740, 102790, 102720, 102640, 102610, 102490, 102440, 102420, 
    102440, 102480, 102470, 102470, 102420, 102430, 102450, 102460, 102460, 
    102450, 102450, 102310, 102270, 102310, 102370, 102410, 102410, 102400, 
    102470, 102460, 102480, 102470, 102400, 102310, 102090, 102040, 101970, 
    102030, 101990, 101960, 102030, 102070, 102040, 102030, 102070, 102060, 
    102160, 102160, 102050, 102030, 102050, 102100, 102160, 102130, 102190, 
    102180, 102230, 102260, 102250, 102230, 102220, 102190, 102110, 102050, 
    102070, 102100, 102130, 102100, 102120, 102060, 102120, 102160, 102170, 
    102150, 102180, 102210, 102230, 102250, 102240, 102230, 102220, 102200, 
    102180, 102160, 102150, 102140, 102140, 102110, 102110, 102090, 102060, 
    102030, 102030, 102000, 101960, 101940, 101930, 101930, 101910, 101890, 
    101880, 101850, 101850, 101790, 101740, 101690, 101660, 101630, 101560, 
    101500, 101440, 101400, 101360, 101330, 101330, 101310, 101280, 101270, 
    101240, 101220, 101190, 101170, 101130, 101090, 101030, 101020, 100990, 
    100920, 100840, 100810, 100750, 100710, 100620, 100520, 100510, 100500, 
    100490, 100430, 100390, 100360, 100310, 100290, 100240, 100200, 100180, 
    100140, 100100, 100060, 100070, 100060, 100010, 99940, 99960, 99960, 
    99970, 99990, 100020, 100020, 100020, 99960, 99990, 100030, 100050, 
    100060, 100040, 100010, 100050, 100080, 100110, 100110, 100090, 100050, 
    100050, 100080, 100090, 100070, 100090, 100060, 100170, 100210, 100300, 
    100390, 100480, 100570, 100700, 100790, 100860, 100940, 101010, 101110, 
    101160, 101190, 101230, 101280, 101320, 101330, 101350, 101450, 101500, 
    101500, 101540, 101500, 101480, 101680, 101700, 101740, 101680, 101720, 
    101710, 101790, 101790, 101770, 101780, 101790, 101750, 101760, 101720, 
    101690, 101690, 101670, 101530, 101640, 101610, 101590, 101570, 101640, 
    101690, 101640, 101650, 101670, 101730, 101840, 101870, 101920, 101970, 
    101940, 101870, 101900, 101940, 101920, 101990, 102000, 102010, 102080, 
    102110, 102130, 102120, 102170, 102170, 102220, 102260, 102310, 102320, 
    102340, 102320, 102200, 102320, 102360, 102410, 102380, 102350, 102270, 
    102190, 102160, 102190, 102270, 102270, 102280, 102280, 102220, 102260, 
    102300, 102370, 102410, 102440, 102420, 102430, 102440, 102410, 102420, 
    102440, 102370, 102380, 102350, 102290, 102280, 102280, 102250, 102200, 
    102110, 102090, 102050, 101990, 101950, 101880, 101890, 101860, 101800, 
    101710, 101670, 101600, 101610, 101630, 101650, 101560, 101560, 101500, 
    101470, 101490, 101540, 101510, 101490, 101450, 101440, 101430, 101360, 
    101380, 101320, 101440, 101400, 101380, 101380, 101360, 101310, 101330, 
    101310, 101230, 101200, 101170, 101140, 101100, 101040, 101000, 100970, 
    100900, 100910, 100880, 100870, 100850, 100870, 100840, 100860, 100840, 
    100800, 100790, 100790, 100780, 100750, 100720, 100710, 100710, 100700, 
    100710, 100660, 100660, 100650, 100650, 100660, 100600, 100600, 100600, 
    100570, 100590, 100620, 100620, 100590, 100590, 100570, 100530, 100510, 
    100520, 100500, 100480, 100470, 100480, 100490, 100440, 100440, 100420, 
    100400, 100390, 100350, 100370, 100380, 100340, 100340, 100330, 100330, 
    100350, 100360, 100340, 100410, 100420, 100410, 100480, 100460, 100460, 
    100500, 100520, 100590, 100640, 100620, 100670, 100750, 100790, 100800, 
    100810, 100850, 100910, 100940, 100990, 100960, 100820, 101150, 101210, 
    101210, 101200, _, 101290, 101280, 101330, 101330, 101380, 101430, 
    101470, 101480, 101490, 101520, 101540, 101520, 101530, 101520, 101520, 
    101530, 101550, 101550, 101560, 101540, 101510, 101510, 101500, 101500, 
    101470, 101450, 101450, 101440, 101440, 101420, 101440, 101440, 101430, 
    101400, 101380, 101390, 101380, 101380, 101360, 101350, 101350, 101370, 
    101380, 101390, 101390, 101380, 101370, 101380, 101350, 101340, 101360, 
    101350, 101340, 101340, 101300, 101280, 101250, 101210, 101180, 101140, 
    101130, 101090, 101060, 101030, 100960, 100940, 100890, 100870, 100830, 
    100800, 100750, 100740, 100730, 100700, 100710, 100670, 100680, 100690, 
    100690, 100670, 100680, 100660, 100650, 100650, 100650, 100680, 100690, 
    100680, 100720, 100730, 100730, 100750, 100730, 100720, 100720, 100690, 
    100690, 100720, 100780, 100810, 100860, 100900, 100940, 100970, 101010, 
    101050, 101080, 101100, 101110, 101130, 101150, 101200, 101220, 101250, 
    101260, 101290, 101290, 101290, 101290, 101290, 101260, 101250, 101250, 
    101240, 101240, 101210, 101160, 101120, 101120, 101090, 101050, 100980, 
    100950, 100920, 100860, 100820, 100800, 100750, 100710, 100640, 100650, 
    100630, 100610, 100530, 100490, 100500, 100450, 100460, 100440, 100400, 
    100370, 100360, 100360, 100320, 100320, 100270, 100280, 100320, 100340, 
    100340, 100330, 100330, 100320, 100300, 100320, 100350, 100330, 100360, 
    100380, 100370, 100360, 100390, 100390, 100400, 100420, 100420, 100420, 
    100440, 100450, 100460, 100440, 100460, 100490, 100490, 100520, 100520, 
    100550, 100570, 100590, 100600, 100610, 100670, 100690, 100720, 100750, 
    100850, 100880, 100840, 100880, 100890, 100910, 100920, 100960, 101000, 
    101010, 101080, 101100, 101130, 101170, 101210, 101230, 101290, 101340, 
    101350, 101390, 101420, 101480, 101460, 101500, 101540, 101550, 101560, 
    101560, 101620, 101620, 101670, 101700, 101750, 101750, 101810, 101840, 
    101870, 101900, 101940, 101980, 101970, 101960, 101930, 101910, 101880, 
    101850, 101810, 101770, 101740, 101690, 101620, 101560, 101530, 101460, 
    101370, 101300, 101180, 101100, 100930, 100840, 100790, 100730, 100690, 
    100620, 100570, 100540, 100460, 100430, 100400, 100390, 100360, 100360, 
    100310, 100220, 100180, 100160, 100060, 99960, 99920, 99870, 99820, 
    99770, 99720, 99670, 99620, 99600, 99560, 99530, 99480, 99480, 99420, 
    99430, 99450, 99470, 99500, 99560, 99630, 99690, 99710, 99730, 99750, 
    99760, 99720, 99720, 99710, 99670, 99640, 99630, 99620, 99620, 99580, 
    99560, 99510, 99460, 99430, 99430, 99400, 99420, 99450, 99480, 99520, 
    99550, 99590, 99610, 99660, 99710, 99740, 99730, 99760, 99750, 99790, 
    99810, 99830, 99830, 99860, 99840, 99850, 99870, 99910, 99950, 99960, 
    99990, 100000, 100030, 100060, 100110, 100130, 100170, 100230, 100260, 
    100320, 100350, 100360, 100390, 100410, 100440, 100430, 100440, 100470, 
    100470, 100460, 100460, 100460, 100460, 100440, 100410, 100390, 100370, 
    100370, 100360, 100360, 100340, 100350, 100350, 100360, 100410, 100450, 
    100470, 100470, 100520, 100560, 100600, 100650, 100670, 100730, 100790, 
    100820, 100880, 100940, 100940, 100950, 101020, 101050, 101100, 101120, 
    101180, 101210, 101260, 101290, 101320, 101340, 101330, 101340, 101350, 
    101290, 101310, 101300, 101300, 101260, 101140, 101140, 101150, 101110, 
    100970, 100870, 100740, 100690, 100740, 100750, 100720, 100670, 100650, 
    100610, 100580, 100570, 100550, 100490, 100490, 100460, 100440, 100470, 
    100500, 100560, 100610, 100670, 100710, 100740, 100770, 100780, 100800, 
    100820, 100840, 100840, 100870, 100960, 101000, 101000, 101020, 101050, 
    101060, 101090, 101120, 101130, 101160, 101190, 101220, 101250, 101280, 
    101300, 101310, 101320, 101310, 101320, 101330, 101360, _, 101400, 
    101430, 101440, 101450, 101460, 101480, 101460, 101490, 101450, 101460, 
    101460, 101460, 101460, 101460, 101460, 101420, 101390, 101350, 101310, 
    101260, 101210, 101130, 101110, 101060, 101030, 100990, 100960, 100950, 
    100880, 100840, 100840, 100800, 100780, 100760, 100760, 100790, 100780, 
    100770, 100770, 100760, 100740, 100720, 100690, 100650, 100600, 100560, 
    100510, 100480, 100430, 100370, 100330, 100280, 100240, 100200, 100160, 
    100120, 100090, 100080, 100080, 100070, 100100, 100120, 100140, 100160, 
    100170, 100180, 100210, 100220, 100230, 100240, 100250, 100280, 100310, 
    100340, 100350, 100370, 100410, 100420, 100440, 100440, 100480, 100520, 
    100560, 100590, 100640, 100720, 100770, 100820, 100880, 100900, 100910, 
    100930, 100960, 100990, 101050, 101070, 101100, 101130, 101170, 101180, 
    101210, 101230, 101230, 101240, 101260, 101240, 101250, 101280, 101330, 
    101330, 101390, 101410, 101420, 101420, 101420, 101410, 101450, 101490, 
    101490, 101490, 101490, 101510, 101540, 101570, 101560, 101540, 101510, 
    101510, 101500, 101480, 101480, 101480, 101470, 101460, 101480, 101490, 
    101480, 101470, 101460, 101430, 101400, 101380, 101360, 101350, 101330, 
    101310, 101300, 101270, 101250, 101240, 101220, 101200, 101180, 101150, 
    101130, 101100, 101080, 101070, 101040, 101040, 101010, 100990, 100960, 
    100930, 100890, 100890, 100870, 100860, 100840, 100840, 100860, 100880, 
    100910, 100920, 100940, 100960, 100970, 101000, 101020, 101060, 101090, 
    101130, 101170, 101190, 101220, 101240, 101270, 101280, 101290, 101300, 
    101320, 101330, 101340, 101360, 101390, 101400, 101420, 101400, 101430, 
    101440, 101460, 101480, 101480, 101500, 101510, 101540, 101560, 101580, 
    101590, 101570, 101560, 101560, 101560, 101540, 101520, 101520, 101520, 
    101500, 101490, 101460, 101460, 101440, 101420, 101390, 101360, 101330, 
    101290, 101270, 101210, 101180, 101170, 101150, 101120, 101050, 101030, 
    100980, 100940, 100920, 100900, 100860, 100820, 100810, 100820, 100860, 
    100850, 100850, 100880, 100870, 100900, 100930, 100940, 100990, 101040, 
    101070, 101120, 101170, 101220, 101260, 101280, 101320, 101360, 101380, 
    101470, 101530, 101580, 101630, 101670, 101700, 101740, 101760, 101810, 
    101850, 101880, 101910, 101940, 101970, 102010, 102030, 102080, 102120, 
    102120, 102150, 102170, 102180, 102210, 102250, 102270, 102300, 102360, 
    102390, 102420, 102450, 102480, 102530, 102590, 102630, 102650, 102690, 
    102720, 102760, 102780, 102820, 102850, 102850, 102860, 102860, 102860, 
    102840, 102840, 102840, 102820, 102840, 102830, 102840, 102810, 102790, 
    102790, 102780, 102790, 102770, 102750, 102750, 102740, 102730, 102730, 
    102730, 102720, 102680, 102690, 102700, 102690, 102670, 102670, 102670, 
    102660, 102640, 102630, 102620, 102620, 102610, 102610, 102580, 102570, 
    102580, 102570, 102580, 102560, 102570, 102580, 102590, 102590, 102610, 
    102610, 102610, 102620, 102630, 102660, 102660, 102670, 102690, 102710, 
    102730, 102740, 102770, 102790, 102820, 102840, 102880, 102910, 102920, 
    102960, 102990, 103020, 103050, 103090, 103140, 103140, 103150, 103180, 
    103200, 103220, 103240, 103260, 103250, 103280, 103280, 103280, 103290, 
    103280, 103280, 103270, 103260, 103250, 103200, 103130, 103080, 103010, 
    102980, 102960, 102910, 102860, 102780, 102770, 102710, 102650, 102540, 
    102450, 102390, 102320, 102250, 102140, 102040, 101920, 101810, 101740, 
    101660, 101540, 101430, 101340, 101280, 101250, 101140, 101040, 101030, 
    100980, 100960, 100960, 101050, 101010, 101040, 101070, 101100, 101110, 
    101160, 101230, 101270, 101340, 101370, 101410, 101450, 101520, 101570, 
    101600, 101660, 101720, 101780, 101820, 101860, 101940, 101970, 101970, 
    102020, 102050, 102070, 102110, 102140, 102170, 102190, 102230, 102210, 
    102220, 102260, 102260, 102230, 102220, 102220, 102200, 102200, 102180, 
    102170, 102140, 102140, 102150, 102160, 102120, 102090, 102090, 102090, 
    102080, 102040, 102050, 102030, 102020, 101980, 101980, 101950, 101920, 
    101900, 101870, 101870, 101860, 101870, 101890, 101950, 102010, 102050, 
    102060, 102080, 102110, 102150, 102190, 102210, 102240, 102240, 102290, 
    102320, 102340, 102370, 102370, 102380, 102380, 102390, 102390, 102400, 
    102420, 102420, 102440, 102470, 102500, 102520, 102540, 102560, 102570, 
    102570, 102550, 102540, 102530, 102550, 102560, 102570, 102570, 102580, 
    102560, 102540, 102530, 102510, 102470, 102450, 102410, 102370, 102310, 
    102240, 102170, 102090, 102030, 101910, 101840, 101730, 101630, 101550, 
    101430, 101350, 101290, 101210, 101130, 101090, 101020, 100950, 100910, 
    100840, 100790, 100710, 100610, 100550, 100470, 100400, 100310, 100210, 
    100160, 100050, 99940, 99850, 99770, 99770, 99720, 99740, 99700, 99780, 
    99820, 99850, 99950, 100000, 100130, 100270, 100410, 100500, 100610, 
    100740, 100850, 100930, 101040, 101100, 101180, 101240, 101290, 101320, 
    101350, 101390, 101380, 101400, 101400, 101420, 101450, 101460, 101440, 
    101420, 101420, 101440, 101440, 101440, 101470, 101480, 101560, 101620, 
    101650, 101650, 101670, 101680, 101680, 101680, 101690, 101680, 101690, 
    101710, 101650, 101730, 101750, 101750, 101770, 101770, 101760, 101760, 
    101770, 101780, 101800, 101820, 101840, 101850, 101860, 101850, 101860, 
    101860, 101840, 101820, 101790, 101800, 101780, 101790, 101800, 101810, 
    101810, 101830, 101850, 101880, 101890, 101910, 101930, 101960, 102000, 
    102050, 102090, 102150, 102170, 102190, 102210, 102230, 102240, 102230, 
    102260, 102270, 102260, 102290, 102290, 102310, 102290, 102260, 102200, 
    102160, 102090, 101960, 101850, 101700, 101680, 101540, 101540, 101550, 
    101570, 101630, 101760, 101830, 101860, 101900, 101990, 102030, 102100, 
    102110, 102150, 102180, 102150, 102160, 102110, 102080, 102060, 102030, 
    101960, 101910, 101890, 101900, 101860, 101790, 101750, 101720, 101660, 
    101610, 101540, 101510, 101450, 101420, 101400, 101420, 101430, 101450, 
    101440, 101440, 101450, 101430, 101460, 101440, 101460, 101490, 101520, 
    101550, 101580, 101630, 101670, 101700, 101730, 101780, 101770, 101830, 
    101850, 101880, 101880, 101940, 101990, 102030, 102070, 102090, 102110, 
    102130, 102150, 102190, 102190, 102250, 102300, 102350, 102390, 102420, 
    102500, 102520, 102550, 102600, 102610, 102630, 102650, 102680, 102670, 
    102680, 102720, 102720, 102710, 102720, 102720, 102720, 102680, 102700, 
    102670, 102660, 102640, 102650, 102670, 102690, 102670, 102630, 102620, 
    102580, 102560, 102520, 102490, 102470, 102450, 102450, 102440, 102420, 
    102370, 102330, 102290, 102220, 102150, 102130, 102080, 101970, 101880, 
    101860, 101880, 101830, 101770, 101700, 101680, 101620, 101620, 101590, 
    101540, 101540, 101510, 101470, 101430, 101440, 101390, 101270, 101210, 
    101150, 101060, 101040, 100980, 101030, 101040, 101060, 101170, 101230, 
    101290, 101350, 101370, 101380, 101340, 101350, 101330, 101380, 101420, 
    101500, 101510, 101540, 101610, 101660, 101590, 101610, 101530, 101430, 
    101420, 101340, 101230, 101150, 101050, 100940, 100910, 100880, 100850, 
    100810, 100760, 100740, 100710, 100660, 100640, 100600, 100580, 100670, 
    100660, 100690, 100730, 100760, 100780, 100800, 100830, 100850, 100870, 
    100890, 100920, 100960, 100980, 101000, 101030, 101030, 101100, 101060, 
    101010, 100970, 100990, 100970, 100970, 100900, 100880, 100770, 100690, 
    100580, 100460, 100350, 100220, 100110, 100090, 100120, 100140, 100200, 
    100280, 100380, 100530, 100660, 100780, 100870, 100950, 100990, 101050, 
    101060, 101070, 101130, 101160, 101120, 101090, 101070, 101020, 100930, 
    100950, 100990, 101000, 101070, 101090, 101180, 101220, 101240, 101280, 
    101310, 101300, 101280, 101250, 101200, 101150, 101120, 101090, 101030, 
    100940, 100850, 100800, 100720, 100660, 100600, 100550, 100490, 100450, 
    100410, 100360, 100360, 100380, 100380, 100350, 100330, 100340, 100360, 
    100420, 100480, 100540, 100580, 100630, 100620, 100610, 100580, 100570, 
    100550, 100560, 100520, 100480, 100470, 100450, 100430, 100430, 100440, 
    100400, 100370, 100350, 100320, 100320, 100330, 100350, 100370, 100340, 
    100380, 100450, 100510, 100470, 100450, 100470, 100490, 100650, 100660, 
    100680, 100670, 100640, 100680, 100750, 100780, 100800, 100810, 100840, 
    100840, 100790, 100790, 100750, 100730, 100690, 100670, 100640, 100600, 
    100580, 100550, 100510, 100480, 100430, 100410, 100380, 100350, 100340, 
    100300, 100330, 100310, 100320, 100290, 100290, 100310, 100360, 100360, 
    100380, 100350, 100370, 100390, 100380, 100330, 100280, 100260, 100250, 
    100260, 100220, 100200, 100200, 100200, 100170, 100130, 100110, 100090, 
    100030, 99990, 99940, 99900, 99890, 99870, 99820, 99740, 99690, 99630, 
    99610, 99600, 99590, 99550, 99480, 99430, 99390, 99370, 99370, 99380, 
    99370, 99380, 99380, 99350, 99300, 99330, 99360, 99380, 99350, 99330, 
    99330, 99330, 99340, 99330, 99370, 99330, 99400, 99410, 99470, 99490, 
    99540, 99600, 99620, 99660, 99670, 99700, 99730, 99750, 99780, 99840, 
    99850, 99880, 99920, 99940, 99950, 99930, 99940, 99960, 99990, 100020, 
    100020, 100020, 100020, 100020, 100030, 100020, 100050, 100070, 100080, 
    100090, 100100, 100110, 100110, 100110, 100130, 100150, 100160, 100170, 
    100170, 100180, 100180, 100190, 100200, 100190, 100160, 100130, 100110, 
    100070, 100040, 100010, 100000, 99980, 99980, 99980, 99990, 100010, 
    100020, 100030, 100030, 100030, 100030, 100020, 100020, 100030, 100030, 
    100050, 100080, 100130, 100140, 100190, 100220, 100250, 100290, 100330, 
    100350, 100380, 100430, 100460, 100510, 100560, 100590, 100630, 100650, 
    100680, 100700, 100700, 100720, 100720, 100720, 100690, 100680, 100680, 
    100690, 100690, 100680, 100660, 100690, 100700, 100680, 100710, 100740, 
    100750, 100800, 100830, 100870, 100900, 100940, 100950, 100980, 101000, 
    101030, 101030, 101020, 101020, 100990, 100990, 100990, 100940, 100910, 
    100900, 100880, 100870, 100860, 100810, 100820, 100830, 100860, 100860, 
    100880, 100880, 100870, 100900, 100900, 100920, 100910, 100910, 100950, 
    100950, 100950, 100950, 100970, 100980, 100990, 101000, 101010, 101030, 
    101030, _, 101060, 101050, 101070, 101070, 101070, 101080, 101080, 
    101060, 101060, 101050, 101070, 101110, 101110, 101110, 101120, _, 
    101130, 101130, 101140, 101140, 101140, 101130, 101130, 101130, 101140, 
    101120, 101160, 101160, 101170, _, 101160, 101150, 101120, 101060, 
    101020, 100980, 100910, 100830, 100790, 100720, 100550, 100380, 100230, 
    100150, 100080, 100030, 99960, 99910, 99870, 99810, 99820, 99800, 99730, 
    99700, 99670, 99630, 99610, 99570, 99580, 99550, 99540, 99510, 99520, 
    99550, 99540, 99540, 99550, 99550, 99560, 99580, 99540, 99530, 99500, 
    99540, 99590, 99720, 99860, 99990, 100110, 100240, 100350, 100520, 
    100700, _, _, _, _, _, 101210, 101270, 101300, 101350, 101400, 101440, 
    101450, 101490, 101540, 101550, 101570, 101580, 101570, 101570, 101560, 
    101520, 101450, 101400, 101360, 101310, 101240, 101240, 101210, 101180, 
    101150, 101120, 101100, 101100, 101080, 101060, 101030, 101030, 101000, 
    101010, 101010, 101010, 101000, 101010, _, 101020, 101000, 101000, 
    100970, 100980, 100950, 100970, 100960, 100960, 100940, 100920, 100910, 
    100930, 100910, 100900, 100910, 100910, 100910, 100920, 100910, 100950, 
    100950, 100970, 100970, 100980, 100990, 101010, 100990, 101010, 101040, 
    101090, 101090, 101070, 101070, 101080, 101080, 101150, 101170, 101120, 
    101050, 101040, 101050, 101120, 101190, 101230, 101250, _, 101340, 
    101430, 101450, 101480, 101490, 101540, 101570, 101580, 101630, 101670, 
    101640, 101620, 101610, 101580, 101570, 101530, 101460, 101420, 101340, 
    101270, 101190, 101110, 101130, 101070, 101020, 100960, 100940, 100920, 
    100870, 100870, 100930, 100990, 100970, 101060, 101050, 101030, 101030, 
    101120, 101100, 101070, 101090, 101100, 101130, 101080, 101080, 101070, 
    100980, 100980, 100890, 100770, 100710, 100610, 100510, 100510, 100480, 
    100430, 100390, 100430, 100470, 100460, 100460, 100480, 100530, 100540, 
    100580, 100600, 100610, 100700, 100730, 100810, 100850, 100840, 100840, 
    100820, 100840, 100860, 100810, 100790, 100750, 100770, 100750, 100740, 
    100690, 100680, 100660, 100650, 100670, 100720, 100770, 100820, 100860, 
    100940, 101020, 101100, 101150, 101170, 101190, 101220, 101250, 101270, 
    101290, 101330, 101340, 101380, 101420, 101430, 101450, 101450, 101450, 
    101450, 101460, 101460, 101470, 101460, 101380, 101420, 101460, 101420, 
    101410, 101390, 101430, 101350, 101330, 101310, 101290, 101240, 101240, 
    101230, 101190, 101160, 101160, 101120, 101050, 100970, 100940, 100890, 
    100880, 100810, 100810, 100790, 100720, 100430, 100330, 100390, 100340, 
    100360, 100350, 100260, 100210, 100180, 100210, 100180, 100160, 100190, 
    100250, 100250, 100280, 100300, 100310, 100350, 100350, 100320, 100350, 
    100400, 100430, 100470, 100510, 100530, 100560, 100580, 100610, 100650, 
    100660, _, 100710, 100740, 100770, 100790, 100860, 100860, 100850, 
    100890, 100920, 100930, 100910, 100920, 100880, 100890, 100910, 100930, 
    100930, 100960, 100960, 100940, 100920, 100860, 100880, 100910, 100900, 
    100870, 100870, 100840, _, 100850, 100880, 100880, 100890, 100860, 
    100830, 100800, 100810, 100820, 100820, 100830, 100820, 100750, 100680, 
    100620, 100550, 100520, 100490, 100450, 100430, 100410, 100410, 100410, 
    100400, 100410, 100450, 100440, 100450, 100410, 100400, 100380, 100370, 
    100350, 100330, 100330, 100280, 100220, 100190, 100110, 100050, 100030, 
    99980, 99910, 99840, 99810, 99780, 99760, 99720, 99690, 99670, 99640, 
    99630, 99630, 99590, 99560, 99540, 99540, 99560, 99550, 99540, 99550, 
    99540, 99520, 99510, 99500, 99500, 99500, 99500, 99480, 99480, 99460, 
    99460, 99440, 99420, 99450, 99490, 99540, 99560, 99590, 99620, 99660, 
    99690, 99680, 99710, _, 99790, 99790, 99810, 99790, 99760, 99740, 99800, 
    99840, 99870, 99910, 99930, 99950, 99930, 99920, 99920, 99930, 99930, 
    99940, 99920, 99930, 99990, 100000, 100010, 100060, 100120, 100170, 
    100250, 100310, 100350, 100400, 100490, 100540, 100590, 100660, 100700, 
    100780, 100860, 100910, 100960, 100990, 101030, 101080, 101140, 101170, 
    101230, 101280, 101330, 101360, 101390, 101420, 101430, 101440, 101460, 
    101470, 101470, 101450, 101430, 101420, 101420, 101440, 101430, 101410, 
    101360, 101360, 101330, 101310, 101300, 101280, 101260, 101230, 101230, 
    101200, 101200, 101180, 101140, 101110, 101060, 101060, 101000, 100990, 
    100990, 100980, 100980, 101010, 100960, 100930, 100900, 100880, 100830, 
    100760, 100630, 100550, 100530, 100450, 100300, 100180, _, 100110, 
    100050, _, 100000, 99930, 99860, 99810, 99850, 99780, 99780, 99840, 
    99820, 99750, 99710, 99680, 99650, 99620, 99580, 99590, 99550, 99550, 
    99590, 99560, 99530, 99520, 99530, 99510, 99490, 99480, 99450, 99440, 
    99440, 99440, 99460, 99440, 99450, 99470, 99470, 99470, 99490, 99490, 
    99540, 99570, 99600, 99650, 99680, 99730, 99760, 99800, 99840, 99880, 
    99930, 99960, 100020, 100040, 100090, 100130, 100170, 100200, 100220, 
    100240, 100250, 100260, 100260, 100260, 100280, 100310, 100330, 100340, 
    100390, 100430, 100500, 100560, 100620, 100670, 100700, 100760, 100830, 
    100880, 100940, 100950, 101000, 101050, 101090, 101100, 101120, 101140, 
    101190, 101230, 101250, 101300, 101330, _, 101410, 101460, 101480, 
    101510, 101550, 101560, 101600, 101640, 101620, 101670, 101730, 101770, 
    101780, 101820, 101880, 101890, 101890, 101920, 101930, 101930, _, _, 
    102030, 102050, 102060, 102090, 102070, 102080, 102040, 102050, 102050, 
    102010, 101980, 101950, 101900, 101880, 101960, 101920, 101680, 101640, 
    101680, 101610, 101580, 101320, 101300, 101150, 100950, 100780, 100750, 
    100680, 100680, 100600, 100430, 100380, 100290, 100320, 100280, 100280, 
    100230, 100350, 100350, 100360, 100320, 100210, 100100, 99980, 99880, 
    99810, 99770, 99790, 99860, 100010, 100140, 100260, 100370, 100460, 
    100480, 100530, 100560, 100580, 100690, 100760, 100800, 100840, _, 
    100940, 100970, 100980, 101000, 101000, 101020, 101050, 101040, _, 
    101070, 101090, 101120, 101110, 101100, 101090, 101080, 101070, 101080, 
    101080, 101100, 101090, 101090, 101090, 101110, 101110, 101120, 101110, 
    101150, 101150, 101180, 101200, 101230, 101240, 101300, 101360, 101400, 
    101440, 101470, 101500, 101500, 101530, 101550, 101550, 101550, 101560, 
    101570, 101560, 101560, 101600, 101590, 101600, 101600, 101610, 101600, 
    101620, 101630, 101630, 101670, 101680, 101670, 101690, 101700, 101680, 
    101680, 101660, 101650, 101620, 101630, 101630, 101640, 101610, 101590, 
    101590, 101570, 101560, 101550, 101510, 101470, 101450, 101450, 101430, 
    101420, 101420, 101390, 101390, 101390, 101360, 101340, 101320, 101300, 
    101310, 101310, 101310, 101300, 101300, 101280, 101280, 101280, 101270, 
    101250, 101240, 101230, 101230, 101240, 101240, 101230, 101220, 101240, 
    101250, 101250, 101220, 101220, 101200, 101190, 101140, 101110, 101090, 
    101080, 101080, 101050, 101040, 101040, 101020, 101020, 101000, 100990, 
    100990, 101000, 100980, 100980, 101010, 101010, 101000, 101020, 101010, 
    101020, 101020, 101020, 101020, 101040, 101050, 101080, 101070, 101060, 
    101070, 101100, 101100, 101120, 101140, 101140, 101150, 101190, 101210, 
    101240, 101250, 101270, 101280, 101300, 101320, 101320, 101350, 101340, 
    101340, 101350, 101330, 101350, 101330, 101330, 101330, 101330, 101300, 
    101280, 101240, 101250, 101260, 101240, 101280, 101310, 101350, 101380, 
    101410, 101440, 101420, 101440, 101470, 101480, 101490, 101500, 101490, 
    101510, 101510, 101510, 101500, 101480, 101490, 101490, 101470, 101440, 
    101480, 101470, 101460, 101480, 101490, 101500, 101500, 101490, 101520, 
    101520, 101540, 101530, 101570, 101600, 101610, 101640, 101630, 101620, 
    101620, 101620, 101630, 101610, 101620, 101600, 101570, 101530, 101460, 
    101440, 101420, 101390, 101350, 101350, 101320, 101280, 101310, 101280, 
    101260, 101260, 101260, 101250, 101230, 101260, 101260, 101220, 101240, 
    101190, 101130, 101080, 101010, 101020, 101030, 100990, 101000, 100890, 
    100850, 100840, 100670, 100590, 100480, 100450, 100240, 100230, 100280, 
    100250, 100230, 100340, 100350, 100340, 100310, 100330, 100330, 100340, 
    100400, 100420, 100480, 100530, 100570, 100640, 100710, 100740, 100790, 
    100850, 100870, 100930, 100980, 101030, 101070, 101120, 101170, 101210, 
    101230, 101250, 101280, 101350, 101380, 101400, 101440, 101490, 101530, 
    101550, 101570, 101620, 101620, 101640, 101650, 101650, 101640, 101630, 
    101650, 101650, 101630, 101640, 101630, 101650, 101630, 101640, 101640, 
    101600, 101620, 101620, 101630, 101630, 101620, 101680, 101680, 101660, 
    101630, 101640, 101630, 101630, 101650, 101640, 101630, 101630, 101630, 
    101620, 101630, 101640, 101630, 101620, 101600, 101550, 101570, 101550, 
    101530, 101510, 101510, 101520, 101510, 101500, 101530, 101510, 101520, 
    101530, 101500, 101530, 101580, 101560, 101580, 101590, 101620, 101670, 
    101750, 101750, 101750, 101750, 101760, 101770, 101770, 101770, 101790, 
    101800, 101790, 101770, 101760, 101720, 101720, 101690, 101670, 101620, 
    101610, 101580, 101560, 101530, 101490, 101460, 101430, 101400, 101360, 
    101340, 101300, 101270, 101260, 101220, 101160, 101130, 101080, 101040, 
    101000, 100940, 100850, 100790, 100720, 100660, 100570, 100480, 100430, 
    100430, 100420, 100400, 100400, 100410, 100420, 100420, 100440, 100470, 
    100600, 100620, 100700, 100740, 100780, 100860, 100900, 100930, 100970, 
    100960, 100970, 100920, 100910, 100930, 100910, 100870, 100870, 100850, 
    100820, 100800, 100780, 100760, 100710, 100660, 100650, 100630, 100610, 
    100600, 100590, 100560, 100550, 100550, 100530, 100510, 100490, 100470, 
    100430, 100390, 100360, 100350, 100340, 100300, 100230, 100170, 100100, 
    99990, 99920, 99900, 99840, 99780, 99740, 99700, 99680, 99690, 99730, 
    99740, 99790, 99810, 99820, 99870, 99890, 99940, 99960, 99970, 100010, 
    99990, 99970, 99970, 99950, 99930, 99900, 99890, 99880, 99880, 99860, 
    99870, 99910, 99910, 99910, 99870, 99850, 99800, 99730, 99690, 99660, 
    99620, 99550, 99500, 99450, 99420, 99410, 99390, 99360, 99340, 99310, 
    99310, 99330, 99350, 99420, 99430, 99450, 99500, 99500, 99470, 99470, 
    99500, 99490, 99450, 99460, 99420, 99410, 99420, 99410, 99380, 99420, 
    99440, 99460, 99500, 99550, 99580, 99630, 99700, 99730, 99760, 99780, 
    99830, 99840, 99850, 99860, 99870, 99850, 99840, 99850, 99850, 99820, 
    99800, 99790, 99820, 99830, 99860, 99900, 99980, 100050, 100130, 100180, 
    100260, 100310, 100400, 100470, 100520, 100580, 100600, 100600, 100590, 
    100550, 100450, 100360, 100300, 100200, 100090, 100010, 99900, 99870, 
    99800, 99820, 99830, 99840, 99860, 99930, 99960, 100070, 100130, 100210, 
    100270, 100310, 100330, 100370, 100400, 100400, 100420, 100410, 100430, 
    100410, 100430, 100400, 100370, 100340, 100350, 100340, 100310, 100330, 
    100330, 100340, 100340, 100390, 100400, 100410, 100430, 100440, 100450, 
    100480, 100500, 100530, 100530, 100530, 100530, 100540, 100560, 100560, 
    100550, 100560, 100600, 100580, 100590, 100610, 100620, 100640, 100660, 
    100690, 100730, 100730, 100770, 100790, 100850, 100880, 100910, 100940, 
    100930, 100990, 101000, 101000, 101040, 101080, 101090, 101130, 101170, 
    101190, 101200, 101230, 101230, 101230, 101280, 101310, 101320, 101330, 
    101330, 101340, 101320, 101320, 101270, 101250, 101190, 101150, 101070, 
    101010, 100980, 100940, 100900, 100880, 100840, 100830, 100830, 100810, 
    100790, 100790, 100800, 100820, 100840, 100830, 100840, 100840, 100800, 
    100760, 100710, 100690, 100710, 100630, 100630, 100610, 100620, 100580, 
    100590, 100590, 100580, 100520, 100450, 100440, 100370, 100270, 100170, 
    100140, 100120, 100090, 100120, 100110, 100090, 100060, 100020, 99950, 
    99900, 99800, 99660, 99630, 99660, 99730, 99840, 99930, 99970, 100020, 
    100090, 100160, 100210, 100290, 100300, 100320, 100380, 100400, 100460, 
    100480, 100510, 100570, 100550, 100540, 100530, 100540, 100520, 100470, 
    100440, 100450, 100480, 100490, 100470, 100450, 100520, 100510, 100520, 
    100520, 100530, 100540, 100530, 100560, 100600, 100620, 100630, 100660, 
    100660, 100670, 100670, 100670, 100660, 100680, 100660, 100650, 100650, 
    100670, 100670, 100710, 100710, 100730, 100730, 100710, 100720, 100730, 
    100730, 100740, 100750, 100770, 100760, 100720, 100700, 100680, 100620, 
    100610, 100570, 100570, 100600, 100590, 100600, 100610, 100650, 100680, 
    100730, 100800, 100830, 100890, 100960, 101030, 101090, 101160, 101220, 
    101270, 101320, 101350, 101400, 101440, 101490, 101570, 101600, 101640, 
    101690, 101710, 101710, 101760, 101820, 101840, 101870, 101900, 101900, 
    101890, 101900, 101910, 101930, 101940, 101940, 101910, 101880, 101840, 
    101780, 101740, 101690, 101670, 101630, 101600, 101560, 101510, 101470, 
    101420, 101310, 101250, 101190, 101110, 101060, 101020, 100950, 100880, 
    100830, 100810, 100760, 100740, 100690, 100610, 100590, 100500, 100460, 
    100390, 100390, 100290, 100300, 100280, 100250, 100210, 100180, 100160, 
    100130, 100120, 100140, 100130, 100120, 100150, 100150, 100160, 100150, 
    100140, 100170, 100170, 100230, 100230, 100210, 100230, 100230, 100230, 
    100230, 100210, 100200, 100150, 100090, 100050, 100030, 100010, 99970, 
    100000, 100030, 100020, 100010, 99960, 99960, 99990, 100000, 100010, 
    99990, 99980, 99950, 99950, 99890, 99830, 99790, 99750, 99690, 99610, 
    99550, 99490, 99380, 99380, 99370, 99370, 99310, 99170, 99090, 99100, 
    99040, 99010, 98960, 98940, 98920, 98890, 98780, 98810, 98820, 98850, 
    98870, 98870, 98950, 98990, 99070, 99100, 99190, 99210, 99240, 99330, 
    99400, 99450, 99490, 99580, 99700, 99810, 99930, 99980, 100050, 100140, 
    100190, 100240, 100310, 100350, 100370, 100410, 100450, 100480, 100490, 
    100560, 100610, 100640, 100630, 100630, 100690, 100720, 100770, 100790, 
    100800, 100850, 100890, 100910, 100890, 100910, 100930, 100980, 101060, 
    101090, 101070, 101080, 101090, 101120, 101140, 101120, 101120, 101110, 
    101110, 101130, 101180, 101210, 101230, 101230, 101270, 101280, 101280, 
    101270, 101280, 101290, 101270, 101260, 101250, 101270, 101280, 101280, 
    101280, 101290, 101290, 101300, 101270, 101260, 101270, 101280, 101270, 
    101290, 101300, 101320, 101320, 101340, 101370, 101400, 101400, 101410, 
    101410, 101410, 101410, 101400, 101380, 101400, 101400, 101420, 101420, 
    101410, 101390, 101370, 101360, 101380, 101380, 101400, 101410, 101420, 
    101430, 101440, 101440, 101430, 101420, 101420, 101410, 101400, 101340, 
    101340, 101320, 101290, 101270, 101240, 101210, 101190, 101170, 101140, 
    101130, 101130, 101090, 101090, 101060, 101040, 101010, 101010, 101020, 
    101000, 100990, 100940, 100910, 100880, 100850, 100820, 100840, 100810, 
    100780, 100730, 100740, 100670, 100630, 100560, 100560, 100490, 100490, 
    100440, 100410, 100340, 100280, 100220, 100150, 100060, 100050, 100020, 
    100010, 99960, 99960, 99940, 99910, 99890, 99860, 99810, 99770, 99760, 
    99760, 99730, 99710, 99700, 99720, 99740, 99750, 99760, 99750, 99770, 
    99760, 99780, 99790, 99780, 99800, 99820, 99840, 99840, 99850, 99870, 
    99860, 99840, 99790, 99720, 99670, 99640, 99590, 99560, 99500, 99530, 
    99510, 99520, 99570, 99650, 99710, 99790, 99880, 99960, 100060, 100130, 
    100210, 100250, 100260, 100300, 100280, 100270, 100250, 100240, 100180, 
    100170, 100150, 100140, 100110, 100070, 100070, 100090, 100120, 100130, 
    100210, 100230, 100280, 100380, 100430, 100490, 100540, 100560, 100610, 
    100650, 100660, 100680, 100670, 100670, 100620, 100590, 100550, 100560, 
    100550, 100520, 100540, 100550, 100600, 100620, 100700, 100780, 100810, 
    100870, 100950, 101040, 101080, 101150, 101210, 101230, 101240, 101280, 
    101320, 101300, 101290, 101440, 101520, 101550, 101580, 101580, 101590, 
    101660, 101690, 101700, 101710, 101730, 101700, 101670, 101610, 101580, 
    101560, 101490, 101450, 101410, 101340, 101280, 101180, 101120, 101010, 
    100910, 100880, 100810, 100780, 100660, 100620, 100560, 100460, 100420, 
    100170, 100110, 100100, 100100, 100100, 100100, 100080, 100100, 100090, 
    100100, 100130, 100100, 100170, 100170, 100220, 100320, 100320, 100390, 
    100450, 100530, 100560, 100650, 100750, 100800, 100860, 100920, 101010, 
    101010, 101010, 101070, 101130, 101180, 101210, 101230, 101300, 101330, 
    101340, 101360, 101380, 101390, 101430, 101420, 101450, 101480, 101500, 
    101510, 101530, 101560, 101500, 101490, 101510, 101440, 101400, 101330, 
    101290, 101240, 101130, 101070, 101040, 100940, 100900, 100810, 100740, 
    100680, 100580, 100590, 100550, 100560, 100540, 100570, 100570, 100570, 
    100610, 100630, 100620, 100660, 100660, 100700, 100710, 100730, 100720, 
    100710, 100690, 100650, 100620, 100580, 100580, 100560, 100570, 100580, 
    100600, 100630, 100640, 100690, 100700, 100770, 100790, 100820, 100820, 
    100820, 100830, 100850, 100890, 100890, 100900, 100930, 100970, 101030, 
    101070, 101110, 101160, 101200, 101250, 101310, 101390, 101440, 101490, 
    101520, 101580, 101630, 101660, 101690, 101760, 101790, 101810, 101810, 
    101850, 101860, 101890, 101900, 101910, 101900, 101890, 101870, 101860, 
    101820, 101800, 101760, 101700, 101650, 101630, 101600, 101540, 101520, 
    101500, 101430, 101400, 101370, 101340, 101340, 101330, 101360, 101390, 
    101400, 101410, 101410, 101440, 101440, 101450, 101440, 101420, 101430, 
    101430, 101480, 101500, 101500, 101530, 101500, 101470, 101440, 101440, 
    101470, 101470, 101500, 101510, 101550, 101570, 101590, 101640, 101640, 
    101680, 101720, 101770, 101800, 101840, 101890, 101920, 101950, 102000, 
    102020, 102060, 102090, 102110, 102140, 102180, 102190, 102220, 102240, 
    102280, 102310, 102320, 102340, 102330, 102350, 102380, 102400, 102400, 
    102420, 102440, 102430, 102450, 102460, 102480, 102490, 102520, 102530, 
    102560, 102590, 102590, 102620, 102650, 102660, 102650, 102660, 102600, 
    102570, 102630, 102620, 102650, 102640, 102690, 102720, 102740, 102750, 
    102770, 102780, 102800, 102840, _, 102880, 102910, 102910, 102940, 
    102940, 102940, 102960, 102960, 102990, 103000, 103010, 103030, 103030, 
    103040, 103050, 103050, 103060, 103050, 103060, 103060, 103070, 103060, 
    103090, 103100, 103120, 103130, 103140, 103150, 103180, 103190, 103190, 
    103210, 103220, 103250, 103260, 103270, _, 103270, 103300, 103300, 
    103310, 103310, 103330, 103320, 103340, 103350, 103360, 103380, 103380, 
    103390, 103370, 103360, _, 103370, 103370, 103360, 103350, 103340, 
    103340, 103370, 103350, 103350, 103340, 103340, 103340, 103300, 103300, 
    103320, _, 103350, _, 103340, 103340, 103310, 103290, 103290, 103280, 
    103260, 103270, 103250, 103240, 103220, _, 103230, 103220, 103200, 
    103200, 103200, 103200, 103200, 103190, 103170, 103180, 103190, 103210, 
    103220, 103240, 103240, 103210, 103190, 103190, 103180, 103190, 103190, 
    103170, 103170, 103150, 103140, 103130, 103110, 103100, 103100, 103130, 
    103120, 103120, 103100, 103100, 103110, 103130, 103150, 103150, 103160, 
    103150, 103140, 103130, 103150, 103150, 103160, 103140, 103150, 103150, 
    103160, 103150, 103140, 103130, 103130, 103140, 103120, 103130, 103120, 
    103130, 103150, 103140, 103150, 103180, 103180, 103170, 103160, 103140, 
    103110, 103100, 103110, 103100, 103090, 103100, 103110, 103100, 103080, 
    103080, 103080, 103060, 103030, 103020, 103010, 103000, 102990, 102980, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 102650, 102620, 102600, 102570, 102550, 102520, 102510, 102490, 
    102440, 102420, 102430, 102390, 102390, 102370, 102350, 102310, 102280, 
    102260, 102230, 102220, 102230, 102220, 102200, 102190, 102150, 102100, 
    102020, 101950, 101900, 101830, 101770, 101660, 101550, 101490, 101360, 
    101260, 101200, 101080, 100970, 100870, 100750, 100620, 100470, 100380, 
    100280, 100160, 100050, 99940, 99800, 99670, 99590, 99500, 99430, 99380, 
    99320, 99270, 99200, 99120, 99060, 99010, _, 98980, 99080, 99180, 99290, 
    99360, 99460, 99550, 99610, 99630, 99640, 99590, 99530, 99460, 99370, 
    99310, 99230, 99120, 98960, 98790, 98540, 98240, 97970, 97930, 97860, 
    97900, 97900, 98090, 98220, 98370, 98510, 98630, 98720, 98740, 98740, 
    98690, 98680, 98690, 98760, 98830, 98870, 98930, 98970, 99020, 99050, 
    99030, 99030, 99050, 99130, 99180, 99230, 99240, 99290, 99330, 99370, 
    99410, 99460, 99490, 99530, 99540, 99620, 99640, 99680, 99750, 99770, 
    99800, 99830, 99860, 99900, 99930, 99950, 99980, _, 100020, 100110, 
    100180, 100270, 100290, 100380, 100460, 100530, 100600, 100660, 100720, 
    100770, 100800, 100830, 100840, 100880, 100910, 100940, 100970, 100990, 
    101030, 101080, 101120, 101130, 101190, _, 101220, 101240, 101260, 
    101290, 101310, 101350, 101370, 101410, 101410, 101440, 101450, 101470, 
    101490, 101510, 101510, 101540, 101540, 101560, 101590, 101610, 101650, 
    101660, 101670, 101690, 101720, 101730, 101750, 101740, 101760, 101790, 
    101820, 101840, 101870, 101880, 101880, 101880, 101880, 101880, 101880, 
    101890, 101890, 101880, 101870, 101880, 101870, 101840, 101830, 101810, 
    101790, 101790, 101760, 101750, 101750, 101770, 101770, 101770, 101750, 
    101720, 101710, 101680, 101660, 101620, 101590, 101570, 101550, 101520, 
    101480, 101460, 101430, 101410, 101380, 101360, 101330, 101310, 101280, 
    101260, 101260, 101240, 101210, 101190, 101150, 101110, 101060, 101040, 
    101000, 100970, 100950, 100910, 100880, 100840, 100790, 100740, 100680, 
    _, 100550, 100420, 100310, 100180, 100090, 100070, 100020, 100020, 99990, 
    99980, 99950, 99920, 99890, 99860, 99810, 99780, 99710, 99710, 99680, 
    99630, 99600, 99550, 99470, 99420, 99410, 99400, 99360, 99370, 99390, 
    99450, 99490, 99520, 99530, 99580, 99690, 99720, 99710, 99770, 99800, 
    99850, 99870, 99900, 99930, 99980, 100000, 100060, 100100, 100100, 
    100110, 100190, 100220, 100220, 100220, 100230, 100240, 100240, 100260, 
    100310, 100360, 100410, 100490, 100600, 100700, 100810, 100900, 101010, 
    101150, 101310, 101450, 101580, 101710, 101780, 101850, 101910, 101960, 
    102010, 102030, 102050, 102070, 102080, 102080, 102090, 102100, 102080, 
    102080, 102050, 102030, 102000, 101970, 101960, 101930, 101910, 101890, 
    _, 101850, 101820, _, 101770, 101740, 101710, 101690, 101660, 101650, 
    101680, 101670, 101640, 101600, 101620, 101600, 101570, 101570, 101550, 
    101540, 101520, 101520, 101550, 101570, 101590, 101610, 101630, 101620, 
    101640, 101650, 101670, 101660, 101670, 101700, 101730, 101770, 101770, 
    101790, 101810, 101800, 101820, 101800, 101800, 101800, 101790, 101790, 
    101770, 101760, 101730, 101690, 101660, 101620, 101590, 101550, 101510, 
    101470, 101370, 101350, 101310, 101260, 101200, 101150, 101090, 101020, 
    100950, 100880, 100810, 100770, 100720, 100670, 100640, 100600, 100570, 
    100530, 100540, _, 100560, 100560, 100570, 100570, 100580, 100610, 
    100640, 100670, 100710, 100750, 100770, 100780, 100780, 100800, 100810, 
    100830, 100850, 100880, 100930, 100950, 100970, 100990, 101030, 101030, 
    101040, 101070, 101090, 101140, 101190, 101200, 101240, 101310, 101370, 
    101410, 101440, 101480, 101500, 101540, 101550, 101560, 101570, 101590, 
    101610, 101630, 101640, 101630, 101620, 101600, 101600, 101590, 101590, 
    101600, 101600, 101620, 101660, 101670, 101690, _, 101690, 101670, 
    101670, 101690, 101690, 101690, 101700, 101710, 101710, 101710, 101710, 
    101700, 101690, _, 101670, 101640, 101610, 101580, 101560, 101540, 
    101540, 101520, 101500, 101460, 101410, 101380, 101350, 101310, 101270, 
    101250, 101210, 101160, 101120, 101100, 101060, 101000, 100940, 100890, 
    100830, 100790, 100740, 100660, 100590, 100510, 100420, 100310, 100180, 
    100080, 99980, 100000, 100010, 100050, 100030, 100020, 100030, 100030, 
    99990, 100000, 99980, 99960, 99920, 99890, 99870, _, 99880, 99850, 99830, 
    99780, 99730, 99690, 99620, _, 99500, 99510, 99500, 99500, 99540, 99600, 
    99640, 99680, 99720, 99790, 99830, 99860, 99880, 99890, 99920, 99930, 
    99930, 99940, 99970, 99970, 100000, 100010, 100030, 100030, 100000, 
    99990, 99950, 99930, _, 99900, 99880, 99850, 99850, 99810, 99780, 99740, 
    99690, 99660, 99620, 99650, 99650, 99600, 99570, 99570, 99570, 99590, 
    99610, 99630, 99630, 99620, 99600, 99610, 99590, 99550, 99570, 99560, 
    99590, 99580, 99580, 99560, 99550, 99530, 99510, 99490, 99460, 99450, 
    99430, 99440, 99470, 99480, 99490, 99500, 99460, 99450, _, _, _, 99520, 
    99510, 99510, 99490, 99490, 99490, 99500, 99530, 99550, 99540, 99540, 
    99570, 99580, 99590, 99630, 99650, 99680, 99710, 99710, 99710, 99720, 
    99760, 99810, 99840, 99870, 99890, 99920, 99980, 100030, 100070, 100090, 
    100130, 100140, 100150, 100160, 100170, 100190, 100190, 100210, 100260, 
    100300, 100350, 100380, 100390, 100410, 100420, 100430, 100420, 100430, 
    100450, 100450, 100470, 100480, 100480, 100490, 100480, 100460, 100480, 
    100460, 100480, 100460, 100490, 100490, 100510, 100510, 100510, 100530, 
    100540, 100560, 100530, 100530, 100540, 100540, 100560, 100570, 100590, 
    100610, 100620, 100620, 100640, 100650, 100650, 100650, 100660, 100660, 
    100690, 100700, 100730, 100750, 100750, 100770, 100750, 100740, 100750, 
    100750, 100760, 100780, 100760, 100760, 100770, 100780, 100770, 100770, 
    100770, 100750, 100730, 100730, 100700, 100690, 100670, 100660, 100670, 
    100660, 100650, 100640, 100630, 100590, 100590, 100580, 100550, 100540, 
    100540, 100530, 100530, 100530, 100560, 100590, 100610, 100620, 100640, 
    100630, 100630, 100670, 100640, 100680, 100700, 100730, 100750, 100770, 
    100790, 100820, 100830, 100810, 100830, 100850, 100850, 100900, 100930, 
    _, 100990, 101000, 101020, 101040, 101060, 101070, 101070, 101080, 
    101070, 101090, 101120, 101150, 101170, 101190, 101190, 101210, 101190, 
    101180, 101150, 101130, 101130, 101110, 101120, 101080, 101080, 101050, 
    101020, 101000, 101010, 100980, 100940, _, 100840, 100820, 100810, 
    100800, 100750, 100670, 100650, 100600, 100520, 100420, 100220, 100210, 
    100060, 99990, 99960, 99890, 99750, _, 99450, 99280, 99180, 99100, 98950, 
    98830, 98710, 98560, 98520, 98520, 98560, 98530, 98510, 98490, 98470, 
    98410, 98390, 98360, 98350, 98330, 98330, _, 98350, 98380, 98420, 98510, 
    98560, 98600, 98730, 98850, 98970, 99120, 99260, 99330, 99360, 99520, 
    99530, 99590, 99680, 99750, 99820, 99840, 99840, 99830, 99600, 99600, 
    99580, 99460, 99330, 99390, 99270, 99250, 99230, 99090, 98890, 98790, 
    98720, 98750, 98650, 98670, 98590, 98460, 98360, 98270, 98160, 98060, 
    97960, 97900, 97820, 97790, 97730, _, 97720, 97680, 97610, 97560, 97490, 
    97440, 97440, 97490, 97550, 97660, 97740, 97780, 97810, 97840, 97880, 
    97910, 97940, 97940, 97980, 97980, 97980, _, 97970, 97940, 97930, 97940, 
    97940, 97940, 97970, 97990, 98010, 98010, 98010, 98020, 97990, 97980, 
    97960, 97950, 97930, 97900, 97880, 97850, 97830, 97850, 97860, 97870, 
    97900, 97940, 97970, 97950, 98020, 98090, 98120, 98190, 98210, 98320, 
    98410, 98500, 98580, 98710, 98780, 98880, 98990, 99120, 99190, 99290, 
    99410, 99510, 99630, 99710, 99780, 99820, 99880, 99930, 99970, 99980, 
    100030, 100060, 100080, 100090, 100090, 100060, 100110, 100090, 100060, 
    100030, 99980, 99940, 99880, 99810, 99860, 99800, 99760, 99750, 99740, 
    99680, 99660, 99620, 99590, 99560, 99510, 99510, 99540, 99570, 99580, 
    99580, 99580, 99560, 99540, 99500, 99480, 99450, 99420, 99390, 99350, 
    99340, 99300, 99260, 99200, 99150, 99080, 99000, 98840, 98820, 98720, 
    98640, 98590, 98550, 98560, 98550, 98570, 98610, 98650, 98670, 98700, 
    98710, 98710, 98670, 98720, 98740, 98840, 98880, 98890, 98940, 98940, 
    98950, 98930, 98920, 98900, 98890, 98880, 98890, 98910, 98950, 98950, 
    98950, 98930, 98850, 98810, 98760, 98690, 98640, 98600, 98570, 98530, 
    98520, 98530, 98560, 98540, 98490, 98520, 98620, 98680, 98780, 98890, 
    98990, 99070, 99120, 99220, 99270, 99340, 99370, 99460, 99510, 99610, 
    99640, 99680, 99730, 99780, 99830, 99850, 99870, 99930, 99980, 100000, 
    100040, 100060, 100110, 100110, 100140, 100230, 100240, 100270, 100340, 
    100380, 100430, 100410, 100440, 100420, 100400, 100360, 100310, 100240, 
    100170, 100140, 100010, 99920, 99810, 99680, 99550, 99410, 99270, 99120, 
    98930, 98720, 98520, 98260, 97980, 97710, 97390, 97210, 97030, 96830, 
    96690, 96590, 96510, 96500, 96530, 96560, 96560, 96560, 96550, 96560, 
    96560, 96590, 96600, 96620, 96660, 96770, 96840, 96890, 96930, 96960, 
    96990, 96990, 97000, 96990, 96960, 96910, 96890, 96860, 96740, 96750, 
    96700, 96670, 96640, 96650, 96650, 96650, 96710, 96640, 96590, 96600, 
    96640, 96760, 96920, 97080, 97230, 97390, 97480, 97600, 97710, 97770, 
    97860, 97940, 97990, 98060, 98080, 98090, 98120, 98170, 98190, 98250, 
    98300, 98380, 98430, 98490, 98530, 98590, 98580, 98610, 98600, 98620, 
    98620, 98620, 98650, 98650, 98650, 98660, 98670, 98680, 98660, 98650, 
    98640, 98620, 98600, 98600, 98610, 98620, 98650, 98690, 98710, 98750, 
    98790, 98790, 98810, 98840, 98860, 98900, 98970, 99020, 99070, 99130, 
    99210, 99240, 99260, 99280, 99300, 99330, 99360, 99370, 99370, 99360, 
    99370, 99380, 99370, 99370, 99360, 99370, 99380, 99420, 99440, 99460, 
    99490, 99500, 99510, 99560, 99610, 99640, 99660, 99690, 99730, 99760, 
    99790, 99820, 99840, 99870, 99910, 99970, 100010, 100020, 100050, 100080, 
    100110, 100120, 100150, 100150, 100160, 100160, 100140, 100070, 100080, 
    100070, 100020, 99960, 99940, 99900, 99860, 99830, 99790, 99750, 99730, 
    99750, 99770, 99750, 99750, 99720, 99690, 99620, 99630, 99600, 99530, 
    99450, 99380, 99330, 99270, 99250, 99220, 99180, 99130, 99110, 99070, 
    98960, 98870, 98750, 98630, 98540, 98510, 98470, 98520, 98550, 98590, 
    98650, 98680, 98680, 98620, 98690, 98760, 98860, 98930, 98980, 99060, 
    99100, 99090, 99110, 99170, 99240, 99280, 99330, 99360, 99390, 99430, 
    99480, 99510, 99530, 99540, 99590, 99640, 99700, 99730, 99750, 99760, 
    99800, 99830, 99850, 99910, 99920, 99900, 99910, 99950, 99960, 100000, 
    100000, 100020, 100030, 100030, 100040, 100080, 100110, 100110, 100100, 
    100120, 100140, 100170, 100160, 100170, 100170, 100150, 100170, 100170, 
    100190, 100170, 100130, 100110, 100100, 100070, 100070, 100030, 100030, 
    100030, 100020, 100000, 99990, 99960, 99940, 99920, 99880, 99860, 99850, 
    99860, 99870, 99860, 99870, 99860, 99830, 99800, 99770, 99740, 99730, 
    99690, 99690, 99650, 99660, 99660, 99650, 99670, 99660, 99670, 99680, 
    99680, 99690, 99700, 99720, 99760, 99790, 99810, 99830, 99860, 99870, 
    99880, 99900, 99940, 99950, 99970, 99990, 100020, 100090, 100070, 100080, 
    100060, 100050, 100030, 100000, 99990, 99970, 99970, 99960, 99910, 99900, 
    99870, 99810, 99770, 99720, 99670, 99610, 99550, 99480, 99370, 99290, 
    99250, 99200, 99130, 99060, 98980, 98890, 98820, 98780, 98720, 98670, 
    98640, 98590, 98540, 98490, 98480, 98460, 98430, 98420, 98410, 98390, 
    98370, 98350, 98300, 98320, 98340, 98350, 98370, 98390, 98380, 98400, 
    98400, 98440, 98470, 98490, 98500, 98510, 98510, 98490, 98540, 98560, 
    98570, 98580, 98600, 98660, 98730, 98790, 98820, 98870, 98910, 98950, 
    98960, 98990, 99020, 99020, 99010, 99000, 99020, 99030, 99050, 99020, 
    99020, 99090, 99100, 99100, 99130, 99130, 99130, 99150, 99150, 99160, 
    99160, 99170, 99170, 99160, 99200, 99180, 99150, 99150, 99170, 99150, 
    99160, 99160, 99140, 99110, 99110, 99070, 99040, 98980, 98940, 98900, 
    98870, 98820, 98800, 98770, 98750, 98730, 98700, 98680, 98670, 98660, 
    98680, 98680, 98690, 98680, 98730, 98740, 98760, 98780, 98800, 98840, 
    98870, 98910, 98950, 98960, 98980, 99010, 99050, 99070, 99090, 99130, 
    99140, 99170, 99230, 99240, 99260, 99290, 99320, 99340, 99350, 99360, 
    99400, 99420, 99450, 99440, 99470, 99490, 99520, 99510, 99520, 99540, 
    99590, 99580, 99570, 99580, 99610, 99620, 99670, 99720, 99650, 99730, 
    99760, 99800, 99830, 99860, 99950, 99960, 99980, 100010, 100060, 100100, 
    100120, 100140, 100180, 100220, 100200, 100180, 100190, 100210, 100260, 
    100270, 100280, 100320, 100340, 100300, 100270, 100250, 100280, 100250, 
    100250, 100250, 100250, 100230, 100230, 100240, 100230, 100200, 100210, 
    100200, 100190, 100180, 100170, 100200, 100200, 100210, 100190, 100210, 
    100190, 100190, 100180, 100170, 100190, 100160, 100160, 100160, 100190, 
    100210, 100190, 100230, 100200, 100190, 100200, 100190, 100260, 100240, 
    100250, 100270, 100240, 100240, 100180, 100210, 100270, 100270, 100300, 
    100330, 100350, 100390, 100410, 100410, 100440, 100480, 100520, 100560, 
    100580, 100630, 100690, 100730, 100740, 100770, 100790, 100840, 100880, 
    100930, 100930, 100970, 100990, 101040, 101050, 101040, 101080, 101080, 
    101110, 101070, 101040, 101060, 101080, 101050, 101070, 101040, 101060, 
    101070, 101080, 101100, 101060, 101070, 101120, 101130, 101140, 101150, 
    101180, 101180, 101170, 101200, 101220, 101180, 101170, 101150, 101100, 
    101080, 101100, 101040, 100990, 100940, 100860, 100790, 100700, 100610, 
    100530, 100410, 100280, 100190, 100090, 99900, 99790, 99670, 99590, 
    99470, 99440, 99290, 99230, 99180, 99190, 99160, 99130, 99120, 99100, 
    99070, 99060, 99000, 99040, 99090, 99120, 99240, 99300, 99450, 99480, 
    99480, 99540, 99590, 99610, 99660, 99690, 99780, 99880, 99970, 100060, 
    100130, 100190, 100220, 100280, 100340, 100410, 100450, 100480, 100520, 
    100530, 100550, 100620, 100670, 100700, 100700, 100730, 100790, 100800, 
    100840, 100860, 100830, 100820, 100850, 100860, 100870, 100880, 100850, 
    100810, 100760, 100670, 100600, 100530, 100480, 100410, 100320, 100320, 
    100230, 100170, 100110, 100000, 99970, 99940, 99890, 99900, 99880, 99910, 
    99870, 99880, 99900, 99930, 99930, 99950, 99990, 100000, 99980, 99960, 
    99960, 99940, 99930, 99950, 99970, 99990, 100000, 99970, 99940, 99920, 
    99880, 99860, 99820, 99730, 99710, 99620, 99550, 99480, 99440, 99360, 
    99300, 99260, 99180, 99140, 99140, 99090, 99020, 99090, 99140, 99190, 
    99230, 99210, 99160, 99140, 99140, 99140, 99150, 99110, 99060, 98940, 
    98850, 98760, 98700, 98650, 98610, 98590, 98510, 98510, 98550, 98590, 
    98490, 98540, 98550, 98530, 98520, 98480, 98430, 98380, 98370, 98440, 
    98480, 98480, 98480, 98490, 98510, 98610, 98640, 98700, 98750, 98790, 
    98870, 98990, 99080, 99160, 99260, 99370, 99450, 99590, 99700, 99780, 
    99860, 99960, 100040, 100140, 100200, 100230, 100290, 100330, 100380, 
    100430, 100450, 100480, 100470, 100470, 100470, 100470, 100460, 100480, 
    100470, 100480, 100480, 100510, 100480, 100490, 100500, 100480, 100490, 
    100490, 100480, 100480, 100490, 100490, 100480, 100470, 100490, 100480, 
    100480, 100480, 100490, 100500, 100490, 100480, 100480, 100510, 100510, 
    100530, 100520, 100520, 100530, 100520, 100540, 100540, 100530, 100510, 
    100500, 100560, 100540, 100540, 100540, 100540, 100550, 100570, 100580, 
    100550, 100540, 100530, 100560, 100540, 100530, 100550, 100560, 100550, 
    100580, 100580, 100580, 100600, 100630, 100620, 100650, 100670, 100680, 
    100720, 100740, 100770, 100800, 100820, 100830, 100820, 100920, 101010, 
    101040, 101050, 101110, 101080, 101010, 101130, 101250, 101290, 101300, 
    101270, 101250, 101220, 101180, 101280, 101310, 101330, 101380, 101360, 
    101420, 101440, 101420, 101380, 101420, 101440, 101450, 101460, 101500, 
    101490, 101450, 101420, 101440, 101440, 101490, 101490, 101480, 101480, 
    101480, 101480, 101530, 101520, 101480, 101470, 101530, 101510, 101500, 
    101490, 101520, 101540, 101550, 101680, 101710, 101750, 101740, 101800, 
    101780, 101800, 101780, 101720, 101670, 101860, 101870, 101860, 101910, 
    101910, 101890, 101880, 101890, 101890, 101830, 101800, 101710, 101730, 
    101780, 101820, 101820, 101830, 101810, 101800, 101740, 101650, 101650, 
    101670, 101660, 101640, 101610, 101590, 101560, 101560, 101540, 101490, 
    101430, 101380, 101300, 101180, 101150, 101150, 101140, 101190, 101130, 
    101120, 101100, 101090, 101020, 100980, 100940, 100910, 100840, 100840, 
    100810, 100820, 100830, 100840, 100850, 100810, 100790, 100800, 100800, 
    100820, 100840, 100850, 100860, 100870, 100900, 100960, 100990, 100950, 
    100970, 100970, 100940, 100940, 100920, 100920, 100930, 100950, 100970, 
    100950, 100960, 100970, 100990, 100960, 100840, 100860, 100860, 100830, 
    100860, 100900, 100910, 100940, 100910, 100910, 100890, 100880, 100920, 
    100920, 100910, 100940, 100920, 100950, 100960, 101000, 101020, 101030, 
    101050, 101080, 101090, 101110, 101110, 101130, 101150, 101160, 101200, 
    101240, 101280, 101300, 101300, 101320, 101320, 101340, 101390, 101360, 
    101340, 101360, 101390, 101410, 101490, 101490, 101520, 101560, 101610, 
    101650, 101680, 101700, 101740, 101770, 101800, 101840, 101910, 101940, 
    101940, 101940, 101950, 101990, 101970, 101970, 102010, 102020, 102020, 
    102030, 102080, 102050, 102060, 102070, 102040, 102040, 102030, 102070, 
    102050, 102030, 102020, 102050, 102070, 102090, 102090, 102050, 102060, 
    102050, 102050, 102040, 102030, 102040, 102040, 102060, 102060, 102060, 
    102040, 102060, 102020, 102010, 101990, 101970, 101970, 101990, 101980, 
    101970, 101990, 102000, 101980, 101940, 101880, 101840, 101740, 101720, 
    101720, 101710, 101690, 101660, 101650, 101700, 101670, 101690, 101690, 
    101710, 101730, 101750, 101770, 101790, 101820, 101860, 101880, 101880, 
    101880, 101870, 101850, 101850, 101840, 101810, 101790, 101790, 101790, 
    101780, 101760, 101730, 101730, 101670, 101640, 101640, 101640, 101640, 
    101660, 101690, 101730, 101740, 101770, 101770, 101800, 101780, 101790, 
    101790, 101790, 101780, 101780, 101770, 101800, 101800, 101800, 101840, 
    101830, 101820, 101810, 101800, 101800, 101810, 101810, 101810, 101840, 
    101860, 101890, 101930, 101900, 101880, 101900, 101900, 101910, 101910, 
    101920, 101930, 101950, 101960, 102010, 102030, 102030, 102010, 102010, 
    102020, 102040, 102050, 102060, 102070, 102110, 102150, 102190, 102190, 
    102200, 102220, 102230, 102230, 102240, 102250, 102260, 102280, 102290, 
    102320, 102320, 102320, 102310, 102330, 102340, 102340, 102360, 102390, 
    102370, 102400, 102420, 102460, 102470, 102490, 102480, 102500, 102520, 
    102530, 102540, 102550, 102540, 102540, 102580, 102590, 102610, 102600, 
    102620, 102620, 102630, 102610, 102630, 102640, 102640, 102680, 102680, 
    102720, 102750, 102780, 102780, 102770, 102780, 102750, 102730, 102740, 
    102720, 102750, 102660, 102660, 102680, 102710, 102710, 102650, 102620, 
    102640, 102590, 102570, 102790, 102640, 102670, 102660, 102680, 102680, 
    102660, 102620, 102600, 102560, 102500, 102460, 102480, 102470, 102460, 
    102440, 102410, 102380, 102370, 102340, 102300, 102270, 102190, 102180, 
    102170, 102170, 102140, 102080, 102090, 102020, 101990, 101940, 101880, 
    101710, 101690, 101670, 101570, 101410, 101330, 101290, 101260, 101170, 
    101040, 100980, 100920, 100850, 100770, 100730, 100710, 100690, 100710, 
    100690, 100670, 100670, 100670, 100660, 100650, 100660, 100680, 100660, 
    100670, 100690, 100700, 100740, 100760, 100700, 100690, 100750, 100700, 
    100680, 100680, 100670, 100680, 100690, 100680, 100700, 100710, 100700, 
    100670, 100680, 100690, 100680, 100680, 100700, 100700, 100720, 100760, 
    100750, 100770, 100770, 100810, 100820, 100850, 100860, 100870, 100880, 
    100920, 100940, 101010, 101030, 101070, 101100, 101120, 101140, 101190, 
    101210, 101260, 101290, 101320, 101350, 101390, 101450, 101490, 101510, 
    101520, 101550, 101570, 101600, 101610, 101630, 101640, 101640, 101660, 
    101700, 101710, 101700, 101670, 101660, 101640, 101630, 101620, 101590, 
    101580, 101580, 101630, 101670, 101780, 101850, 101890, 101950, 102010, 
    102100, 102190, 102270, 102330, 102340, 102400, 102420, 102460, 102470, 
    102480, 102460, 102440, 102460, 102430, 102400, 102370, 102370, 102330, 
    102320, 102290, 102220, 102140, 102080, 102030, 101970, 101910, 101840, 
    101810, 101810, 101800, 101810, 101830, 101810, 101800, 101810, 101780, 
    101760, 101750, 101760, 101760, 101740, 101730, 101740, 101730, 101730, 
    101730, 101700, 101660, 101610, 101600, 101580, 101550, 101520, 101540, 
    101530, 101550, 101550, 101520, 101490, 101410, 101340, 101290, 101220, 
    101190, 101150, 101100, 101050, 101010, 100990, 100980, 101000, 100970, 
    100970, 100960, 100950, 100930, 100960, 100960, 100980, 101000, 100990, 
    101000, 100980, 100950, 100960, 100960, 100930, 100890, 100900, 100880, 
    100880, 100860, 100880, 100900, 100880, 100860, 100830, 100800, 100760, 
    100720, 100660, 100650, 100630, 100610, 100630, 100620, 100610, 100700, 
    100770, 100850, 100890, 100960, 101010, 101020, 101090, 101130, 101210, 
    101230, 101240, 101260, 101260, 101280, 101330, 101360, 101440, 101470, 
    101480, 101530, 101580, 101560, 101640, 101710, 101740, 101760, 101780, 
    101890, 101920, 101930, 102000, 102040, 102060, 102110, 102120, 102130, 
    102130, 102140, 102140, 102140, 102140, 102150, 102160, 102170, 102140, 
    102100, 102060, 102030, 101960, 101850, 101770, 101680, 101570, 101520, 
    101440, 101340, 101260, 101160, 101110, 101070, 101010, 100960, 100960, 
    100980, 101000, 100980, 100960, 100980, 101000, 101070, 101130, 101200, 
    101310, 101400, 101480, 101540, 101580, 101620, 101660, 101700, 101710, 
    101730, 101730, 101720, 101700, 101630, 101600, 101540, 101500, 101490, 
    101430, 101390, 101350, 101280, 101210, 101150, 101070, 100970, 100880, 
    100820, 100760, 100690, 100620, 100590, 100560, 100520, 100520, 100540, 
    100510, 100510, 100510, 100550, 100580, 100620, 100680, 100730, 100790, 
    100820, 100870, 100880, 100930, 101020, 101060, 101120, 101170, 101240, 
    101270, 101290, 101330, 101370, 101410, 101440, 101470, 101510, 101530, 
    101550, 101570, 101620, 101630, 101640, 101650, 101680, 101690, 101660, 
    101640, 101670, 101620, 101590, 101590, 101610, 101620, 101660, 101690, 
    101700, 101680, 101710, 101730, 101760, 101780, 101810, 101860, 101930, 
    101980, 102050, 102110, 102170, 102240, 102310, 102340, 102430, 102470, 
    102530, 102590, 102620, 102680, 102710, 102820, 102890, 102900, 102910, 
    102940, 102970, 103010, 103010, 103000, 103040, 103090, 103090, 103070, 
    103070, 103070, 103070, 103060, 103120, 103210, 103260, 103300, 103360, 
    103410, 103450, 103460, 103480, 103500, 103520, 103520, 103500, 103460, 
    103490, 103500, 103490, 103480, 103480, 103440, 103410, 103380, 103360, 
    103330, 103300, 103290, 103290, 103270, 103260, 103250, 103210, 103180, 
    103170, 103140, 103100, 103070, 103020, 102990, 102970, 102950, 102940, 
    102950, 102930, 102880, 102850, 102790, 102760, 102690, 102660, 102620, 
    102570, 102530, 102500, 102450, 102400, 102340, 102280, 102210, 102130, 
    102050, 101970, 101880, 101830, 101760, 101710, 101680, 101620, 101540, 
    101480, 101400, 101320, 101270, 101200, 101150, 101090, 101030, 101040, 
    101030, 101030, 101020, 101000, 100990, 101020, 101000, 101020, 101010, 
    101020, 101040, 101100, 101160, 101200, 101250, 101280, 101320, 101360, 
    101370, 101390, 101400, 101450, 101500, 101540, 101600, 101630, 101670, 
    101680, 101740, 101750, 101750, 101730, 101760, 101730, 101760, 101770, 
    101790, 101830, 101840, 101860, 101880, 101880, 101910, 101890, 101930, 
    101940, 101950, 101950, 101980, 102010, 102040, 102050, 102070, 102080, 
    102090, 102090, 102100, 102100, 102110, 102150, 102180, 102190, 102180, 
    102170, 102150, 102160, 102170, 102160, 102170, 102200, 102210, 102240, 
    102240, 102240, 102220, 102200, 102170, 102130, 102110, 102090, 102070, 
    102060, 102060, 102080, 102100, 102100, 102080, 102050, 101950, 101950, 
    101890, 101850, 101840, 101820, 101800, 101760, 101720, 101710, 101670, 
    101620, 101560, 101490, 101440, 101370, 101310, 101250, 101190, 101130, 
    101080, 101040, 100970, 100910, 100850, 100790, 100710, 100630, 100560, 
    100490, 100410, 100400, 100370, 100310, 100260, 100230, 100190, 100170, 
    100150, 100120, 100130, 100130, 100140, 100180, 100220, 100260, 100290, 
    100330, 100350, 100380, 100400, 100420, 100450, 100470, 100520, 100540, 
    100590, 100620, 100630, 100650, 100680, 100700, 100730, 100750, 100750, 
    100760, 100800, 100830, 100850, 100900, 100930, 100960, 100960, 100990, 
    101000, 101020, 101020, 101030, 101050, 101080, 101120, 101140, 101180, 
    101190, 101190, 101190, 101230, 101260, 101260, 101270, 101290, 101320, 
    101340, 101340, 101330, 101340, 101330, 101350, 101340, 101350, 101340, 
    101310, 101280, 101270, 101270, 101260, 101300, 101280, 101250, 101230, 
    101200, 101150, 101110, 101120, 101090, 101070, 101100, 101120, 101110, 
    101110, 101100, 101080, 101060, 100980, 100970, 100970, 100910, 100870, 
    100830, 100820, 100850, 100850, 100850, 100830, 100820, 100810, 100790, 
    100770, 100740, 100720, 100660, 100560, 100630, 100640, 100630, 100610, 
    100570, 100540, 100530, 100500, 100470, 100460, 100440, 100410, 100380, 
    100350, 100310, 100280, 100240, 100210, 100200, 100180, 100180, 100170, 
    100180, 100200, 100180, 100190, 100180, 100180, 100160, 100150, 100100, 
    100090, 100040, 100010, 100030, 100030, 99980, 99850, 99800, 99760, 
    99700, 99610, 99530, 99510, 99460, 99430, 99420, 99410, 99390, 99370, 
    99330, 99270, 99220, 99140, 99080, 99040, 99060, 99090, 99110, 99120, 
    99120, 99100, 99080, 99060, 99050, 99070, 99080, 99120, 99260, 99280, 
    99360, 99470, 99500, 99520, 99610, 99690, 99800, 99840, 99910, 99990, 
    100040, 100110, 100200, 100240, 100310, 100330, 100410, 100470, 100530, 
    100590, 100640, 100700, 100740, 100820, 100890, 100950, 101010, 101070, 
    101080, 101130, 101170, 101140, 101180, 101230, 101310, 101340, 101390, 
    101460, 101480, 101490, 101510, 101530, 101550, 101550, 101540, 101510, 
    101530, 101520, 101560, 101580, 101600, 101600, 101600, 101590, 101530, 
    101510, 101450, 101380, 101440, 101420, 101350, 101420, 101440, 101490, 
    101440, 101420, 101370, 101370, 101390, 101400, 101400, 101400, 101390, 
    101410, 101380, 101330, 101280, 101260, 101200, 101080, 101010, 100960, 
    101010, 101040, 101010, 100980, 100990, 100930, 100920, 100910, 100890, 
    100830, 100760, 100640, 100620, 100630, 100650, 100700, 100730, 100700, 
    100710, 100700, 100690, 100640, 100640, 100620, 100550, 100480, 100450, 
    100470, 100470, 100450, 100430, 100390, 100390, 100350, 100290, 100250, 
    100190, 100160, 100100, 100080, 100120, 100060, 100000, 100000, 100010, 
    100020, 100040, 100070, 100100, 100100, 100150, 100160, 100170, 100230, 
    100290, 100360, 100440, 100540, 100610, 100710, 100790, 100880, 100970, 
    101050, 101150, 101240, 101300, 101340, 101380, 101450, 101480, 101520, 
    101550, 101580, 101610, 101640, 101730, 101770, 101800, 101850, 101880, 
    101900, 101910, 101900, 101930, 101970, 102000, 102040, 102060, 102080, 
    102100, 102100, 102120, 102120, 102130, 102120, 102130, 102120, 102100, 
    102100, 102090, 102070, 102080, 102070, 102060, 102050, 102030, 102000, 
    101970, 101960, 101930, 101920, 101890, 101830, 101790, 101760, 101700, 
    101650, 101580, 101560, 101520, 101490, 101440, 101420, 101350, 101310, 
    101280, 101260, 101220, 101170, 101120, 101060, 101040, 101010, 101000, 
    100970, 100970, 100940, 100900, 100870, 100830, 100800, 100780, 100730, 
    100700, 100650, 100570, 100550, 100500, 100480, 100460, 100440, 100390, 
    100370, 100320, 100320, 100300, 100300, 100320, 100330, 100320, 100300, 
    100270, 100270, 100250, 100260, 100250, 100240, 100250, 100290, 100340, 
    100380, 100380, 100380, 100380, 100380, 100370, 100340, 100310, 100270, 
    100230, 100230, 100250, 100230, 100230, 100210, 100210, 100200, 100190, 
    100150, 100120, 100110, 100100, 100090, 100070, 100050, 100010, 99990, 
    99950, 99920, 99880, 99860, 99840, 99800, 99770, 99760, 99730, 99690, 
    99690, 99660, 99620, 99570, 99510, 99530, 99520, 99480, 99420, 99400, 
    99430, 99440, 99440, 99390, 99430, 99400, 99400, 99400, 99380, 99320, 
    99280, 99280, 99310, 99330, 99360, 99350, 99400, 99430, 99450, 99540, 
    99580, 99590, 99610, 99570, 99580, 99570, 99560, 99610, 99630, 99660, 
    99690, 99700, 99760, 99770, 99780, 99770, 99810, 99830, 99770, 99790, 
    99870, 99910, 99940, 99990, 100000, 100030, 100070, 100100, 100090, 
    100190, 100290, 100390, 100400, 100420, 100410, 100460, 100560, 100660, 
    100740, 100820, 100880, 100910, 100960, 101140, 101150, 101180, 101230, 
    101270, 101280, 101330, 101340, 101340, 101340, 101350, 101350, 101320, 
    101280, 101240, 101180, 101110, 101050, 101010, 100980, 100950, 100940, 
    100910, 100930, 100900, 100870, 100850, 100800, 100760, 100740, 100720, 
    100710, 100690, 100700, 100710, 100740, 100700, 100660, 100660, 100650, 
    100720, 100660, 100710, 100710, 100630, 100580, 100670, 100730, 100700, 
    100680, 100710, 100790, 100850, 100880, 100890, 100930, 100980, 101020, 
    101050, 101080, 101180, 101260, 101270, 101300, 101290, 101320, 101300, 
    101290, 101320, 101350, 101450, 101500, 101520, 101550, 101580, 101580, 
    101620, 101660, 101670, 101660, 101710, 101720, 101710, 101710, 101700, 
    101730, 101740, 101720, 101730, 101730, 101720, 101690, 101660, 101670, 
    101660, 101590, 101540, 101490, 101450, 101370, 101310, 101220, 101140, 
    101030, 101010, 100960, 100900, 100830, 100770, 100690, 100600, 100500, 
    100350, 100230, 100110, 100010, 99900, 99760, 99640, 99520, 99460, 99380, 
    99330, 99420, 99330, 99270, 99230, 99190, 99150, 99130, 99160, 99210, 
    99220, 99310, 99380, 99450, 99510, 99560, 99610, 99690, 99740, 99870, 
    99990, 100100, 100170, 100270, 100340, 100440, 100520, 100540, 100540, 
    100620, 100640, 100700, 100750, 100790, 100800, 100830, 100860, 100860, 
    100860, 100860, 100840, 100820, 100760, 100710, 100690, 100700, 100760, 
    100800, 100810, 100910, 100910, 100900, 100890, 100880, 100880, 100880, 
    100900, 100890, 100880, 100840, 100810, 100760, 100730, 100680, 100610, 
    100540, 100480, 100420, 100330, 100230, 100160, 100060, 100010, 99890, 
    99770, 99610, 99500, 99370, 99280, 99220, 99110, 98990, 98890, 98810, 
    98770, 98780, 98750, 98670, 98610, 98580, 98560, 98530, 98490, 98430, 
    98440, 98430, 98440, 98420, 98400, 98380, 98350, 98360, 98380, 98420, 
    98450, 98500, 98510, 98540, 98550, 98560, 98580, 98680, 98720, 98730, 
    98780, 98840, 98820, 98860, 98860, 98890, 98940, 98940, 99000, 99040, 
    99080, 99080, 99130, 99120, 99140, 99140, 99150, 99170, 99180, 99170, 
    99150, 99130, 99110, 99110, 99130, 99140, 99140, 99130, 99140, 99130, 
    99110, 99110, 99090, 99050, 99010, 98980, 99000, 98990, 98990, 98980, 
    98970, 98950, 98950, 98930, 98930, 98890, 98870, 98870, 98890, 98970, 
    99050, 99100, 99110, 99120, 99140, 99200, 99230, 99300, 99300, 99370, 
    99380, 99380, 99450, 99550, 99560, 99580, 99620, 99660, 99640, 99690, 
    99700, 99720, 99730, 99770, 99770, 99760, 99780, 99790, 99760, 99760, 
    99720, 99670, 99630, 99600, 99630, 99630, 99570, 99560, 99570, 99620, 
    99650, 99650, 99690, 99720, 99750, 99770, 99830, 99900, 99960, 100010, 
    100070, 100110, 100160, 100220, 100260, 100310, 100280, 100280, 100340, 
    100390, 100450, 100460, 100490, 100610, 100680, 100720, 100680, 100650, 
    100670, 100710, 100720, 100750, 100760, 100760, 100730, 100720, 100680, 
    100650, 100630, 100580, 100540, 100500, 100490, 100500, 100490, 100460, 
    100430, 100390, 100360, 100340, 100310, 100310, 100300, 100330, 100370, 
    100410, 100450, 100470, 100490, 100500, 100500, 100500, 100510, 100510, 
    100460, 100450, 100440, 100470, 100440, 100440, 100440, 100440, 100410, 
    100390, 100360, 100360, 100350, 100340, 100310, 100370, 100400, 100440, 
    100440, 100440, 100450, 100450, 100430, 100430, 100440, 100440, 100440, 
    100420, 100430, 100440, 100450, 100450, 100450, 100410, 100420, 100400, 
    100370, 100330, 100310, 100290, 100280, 100350, 100340, 100330, 100320, 
    100320, 100260, 100290, 100170, 100080, 100040, 100020, 99850, 99850, 
    99710, 99750, 99720, 99670, 99540, 99460, 99420, 99420, 99430, 99440, 
    99400, 99270, 99210, 99190, 99230, 99300, 99400, 99440, 99440, 99440, 
    99430, 99430, 99470, 99440, 99420, 99390, 99370, 99370, 99350, 99380, 
    99350, 99370, 99400, 99400, 99420, 99430, 99420, 99460, 99460, 99490, 
    99490, 99490, 99510, 99520, 99530, 99540, 99550, 99570, 99630, 99680, 
    99710, 99700, 99690, 99710, 99760, 99810, 99830, 99860, 99900, 99950, 
    99970, 99990, 100010, 100050, 100090, 100080, 100050, 100080, 100120, 
    100120, 100110, 100110, 100110, 100120, 100110, 100120, 100120, 100080, 
    100090, 100080, 100060, 100060, 100040, 100030, 100010, 100010, 100000, 
    99960, 99950, 99910, 99870, 99830, 99790, 99760, 99710, 99640, 99600, 
    99540, 99500, 99450, 99410, 99330, 99290, 99220, 99160, 99160, 99130, 
    99090, 99060, 99030, 98990, 98960, 98930, 98860, 98840, 98820, 98800, 
    98780, 98790, 98780, 98770, 98740, 98730, 98730, 98700, 98690, 98680, 
    98690, 98710, 98720, 98740, 98750, 98780, 98780, 98800, 98840, 98850, 
    98870, 98890, 98920, 98940, 98960, 99000, 99020, 99070, 99120, 99150, 
    99170, 99190, 99210, 99240, 99290, 99340, 99370, 99410, 99430, 99440, 
    99460, 99440, 99410, 99390, 99350, 99330, 99320, 99300, 99290, 99260, 
    99240, 99210, 99170, 99170, 99140, 99120, 99090, 99070, 99070, 99090, 
    99120, 99140, 99150, 99180, 99210, 99250, 99290, 99350, 99370, 99420, 
    99470, 99510, 99580, 99630, 99660, 99770, 99830, 99890, 99940, 100000, 
    100060, 100170, 100260, 100330, 100410, 100490, 100570, 100600, 100700, 
    100770, 100820, 100880, 100920, 100940, 100960, 101010, 101010, 101000, 
    101010, 101090, 101130, 101130, 101170, 101220, 101240, 101260, 101280, 
    101270, 101310, 101330, 101310, 101280, 101290, 101260, 101290, 101290, 
    101290, 101420, 101470, 101540, 101620, 101720, 101790, 101870, 101950, 
    101980, 102030, 102100, 102160, 102190, 102280, 102290, 102290, 102320, 
    102320, 102260, 102300, 102260, 102150, 102020, 101850, 101720, 101660, 
    101570, 101310, 101150, 100990, 100790, 100610, 100430, 100300, 100180, 
    100070, 100020, 100040, 100020, 100020, 100000, 99940, 99860, 99790, 
    99700, 99550, 99430, 99350, 99330, 99320, 99320, 99250, 99110, 99200, 
    99340, 99400, 99530, 99580, 99640, 99720, 99830, 99930, 99970, 100030, 
    100060, 100190, 100220, 100250, 100280, 100310, 100330, 100390, 100410, 
    100380, 100390, 100380, 100390, 100520, 100610, 100670, 100690, 100810, 
    100890, 100880, 100870, 100820, 100860, 100890, 100840, 100790, 100740, 
    100710, 100710, 100710, 100690, 100660, 100680, 100690, 100730, 100780, 
    100810, 100780, 100810, 100800, 100770, 100760, 100730, 100710, 100710, 
    100680, 100710, 100750, 100750, 100760, 100760, 100760, 100790, 100820, 
    100770, 100730, 100700, 100680, 100700, 100740, 100760, 100750, 100750, 
    100740, 100660, 100630, 100630, 100560, 100540, 100510, 100420, 100430, 
    100380, 100280, 100240, 100200, 100180, 100110, 100030, 99960, 99920, 
    99880, 99860, 99830, 99800, 99770, 99760, 99780, 99800, 99820, 99810, 
    99800, 99780, 99750, 99760, 99810, 99850, 99830, 99830, 99820, 99870, 
    99860, 99890, 99890, 99890, 99870, 99900, 99930, 99950, 99970, 100000, 
    99970, 99990, 100020, 100020, 100010, 100030, 100050, 100040, 100030, 
    100030, 99990, 99960, 99970, 99970, 99930, 99890, 99890, 99850, 99820, 
    99780, 99770, 99750, 99750, 99710, 99680, 99650, 99620, 99600, 99570, 
    99530, 99500, 99470, 99460, 99440, 99420, 99390, 99350, 99300, 99290, 
    99260, 99230, 99190, 99180, 99170, 99160, 99160, 99150, 99170, 99200, 
    99220, 99250, 99250, 99260, 99310, 99350, 99380, 99420, 99440, 99480, 
    99530, 99560, 99570, 99610, 99630, 99630, 99610, 99610, 99630, 99630, 
    99650, 99680, 99690, 99750, 99790, 99920, 100000, 100000, 100080, 100150, 
    100240, 100320, 100400, 100520, 100600, 100690, 100740, 100810, 100860, 
    100900, 100950, 101000, 101060, 101110, 101190, 101230, 101260, 101310, 
    101360, 101450, 101500, 101530, 101560, 101560, 101580, 101610, 101650, 
    101710, 101730, 101770, 101810, 101830, 101840, 101910, 101930, 101950, 
    101970, 101990, 102020, 102050, 102060, 102070, 102070, 102090, 102130, 
    102110, 102100, 102120, 102090, 102110, 102110, 102090, 102070, 102030, 
    101990, 101920, 101890, 101820, 101770, 101700, 101630, 101600, 101550, 
    101470, 101380, 101330, 101280, 101240, 101200, 101140, 101100, 101060, 
    101070, 101110, 101110, 101110, 101100, 101100, 101100, 101090, 101030, 
    100960, 100900, 100830, 100770, 100650, 100600, 100500, 100440, 100340, 
    100260, 100220, 100140, 100100, 100060, 100010, 99980, 99920, 99850, 
    99800, 99720, 99660, 99620, 99550, 99520, 99480, 99470, 99490, 99410, 
    99410, 99400, 99420, 99480, 99500, 99570, 99560, 99500, 99530, 99480, 
    99550, 99570, 99580, 99590, 99570, 99580, 99560, 99570, 99580, 99560, 
    99550, 99520, 99510, 99490, 99470, 99480, 99460, 99460, 99430, 99420, 
    99420, 99420, 99420, 99430, 99450, 99470, 99470, 99490, 99530, 99560, 
    99620, 99650, 99670, 99730, 99760, 99820, 99860, 99840, 99910, 99990, 
    100030, 100060, 100120, 100120, 100100, 100120, 100140, 100190, 100190, 
    100220, 100230, 100240, 100260, 100300, 100310, 100290, 100280, 100270, 
    100280, 100270, 100280, 100270, 100280, 100260, 100250, 100230, 100210, 
    100210, 100200, 100210, 100210, 100210, 100200, 100190, 100180, 100150, 
    100110, 100070, 100020, 99950, 99890, 99820, 99810, 99810, 99840, 99840, 
    99850, 99890, 99940, 99970, 100000, 100030, 100070, 100080, 100130, 
    100200, 100260, 100330, 100410, 100480, 100510, 100540, 100560, 100560, 
    100540, 100530, 100520, 100530, 100520, 100550, 100560, 100580, 100600, 
    100570, 100560, 100550, 100520, 100500, 100470, 100430, 100370, 100340, 
    100310, 100270, 100210, 100130, 100020, 99890, 99700, 99470, 99240, 
    99070, 98860, 98670, 98530, 98340, 98160, 98010, 97830, 97630, 97430, 
    97230, 97000, 96790, 96560, 96330, 96210, 96120, 96030, 96020, 96020, 
    96060, 96110, 96310, 96480, 96690, 96840, 96990, 97060, 97220, 97400, 
    97670, 97870, 97890, 97990, 98130, 98340, 98430, 98490, 98570, 98680, 
    98760, 98850, 98900, 98950, 98930, 98940, 98940, 98920, 98910, 98880, 
    98830, 98810, 98770, 98720, 98710, 98670, 98590, 98560, 98500, 98500, 
    98450, 98470, 98450, 98440, 98440, 98470, 98510, 98510, 98560, 98580, 
    98680, 98690, 98770, 98880, 98920, 98990, 99070, 99160, 99270, 99450, 
    99510, 99560, 99620, 99700, 99830, 99890, 99930, 99960, 100060, 100130, 
    100200, 100260, 100310, 100310, 100340, 100370, 100390, 100400, 100450, 
    100490, 100480, 100430, 100440, 100430, 100430, 100390, 100360, 100300, 
    100290, 100290, 100280, 100270, 100280, 100240, 100200, 100220, 100200, 
    100160, 100140, 100110, 100120, 100100, 100100, 100120, 100150, 100190, 
    100220, 100240, 100310, 100360, 100390, 100420, 100480, 100520, 100620, 
    100720, 100780, 100880, 100970, 101020, 101070, 101130, 101160, 101210, 
    101250, 101290, 101320, 101370, 101410, 101450, 101480, 101490, 101540, 
    101560, 101580, 101580, 101620, 101670, 101700, 101710, 101740, 101740, 
    101770, 101730, 101730, 101730, 101760, 101770, 101760, 101750, 101730, 
    101760, 101800, 101800, 101790, 101810, 101780, 101760, 101770, 101800, 
    101810, 101820, 101840, 101870, 101890, 101910, 101940, 101990, 102050, 
    102070, 102030, 102020, 102010, 102020, 102030, 102070, 102100, 102090, 
    102110, 102110, 102100, 102110, 102110, 102100, 102110, 102120, 102130, 
    102070, 102050, 102050, 102060, 102030, 101990, 101990, 102010, 101990, 
    101940, 101880, 101880, 101890, 101850, 101820, 101760, 101690, 101690, 
    101680, 101670, 101670, 101640, 101690, 101720, 101720, 101700, 101690, 
    101680, 101680, 101670, 101780, 101710, 101610, 101590, 101500, 101520, 
    101490, 101490, 101450, 101400, 101400, 101320, 101280, 101270, 101280, 
    101260, 101280, 101270, 101290, 101280, 101310, 101340, 101370, 101400, 
    101420, 101450, 101500, 101540, 101590, 101640, 101730, 101790, 101880, 
    101950, 102000, 102060, 102100, 102140, 102170, 102210, 102250, 102280, 
    102310, 102330, 102350, 102370, 102360, 102330, 102290, 102240, 102170, 
    102150, 102110, 102050, 102030, 101960, 101910, 101820, 101810, 101830, 
    101750, 101790, 101840, 101860, 101810, 101860, 101910, 101940, 101950, 
    101950, 101950, 101930, 101920, 101910, 101890, 101900, 101890, 101900, 
    101880, 101870, 101850, 101860, 101850, 101860, 101860, 101850, 101830, 
    101810, 101830, 101830, 101830, 101820, 101820, 101810, 101800, 101820, 
    101830, 101840, 101840, 101850, 101860, 101880, 101870, 101890, 101900, 
    101890, 101880, 101880, 101860, 101850, 101850, 101870, 101870, 101880, 
    101900, 101910, 101930, 101920, 101950, 101970, 101990, 102040, 102060, 
    102080, 102110, 102150, 102190, 102220, 102230, 102260, 102270, 102280, 
    102300, 102300, 102310, 102350, 102360, 102380, 102400, 102410, 102420, 
    102390, 102390, 102390, 102370, 102370, 102360, 102360, 102350, 102340, 
    102350, 102350, 102350, 102320, 102280, 102260, 102240, 102220, 102240, 
    102220, 102210, 102210, 102240, 102230, 102220, 102190, 102160, 102150, 
    102140, 102130, 102060, 102050, 102060, 102040, 102050, 102030, 102010, 
    102000, 101980, 101990, 101970, 101960, 101940, 101940, 101950, 101950, 
    101950, 101970, 101970, 101960, 102000, 102000, 102010, 102030, 102020, 
    102030, 102020, 102030, 102020, 102050, 102070, 102090, 102090, 102100, 
    102100, 102110, 102120, 102170, 102140, 102180, 102220, 102230, 102230, 
    102270, 102280, 102300, 102300, 102330, 102330, 102360, 102350, 102350, 
    102320, 102320, 102320, 102330, 102370, 102360, 102340, 102410, 102370, 
    102430, 102430, 102450, 102500, 102510, 102520, 102500, 102490, 102490, 
    102480, 102450, 102450, 102410, 102420, 102410, 102380, 102380, 102340, 
    102330, 102310, 102300, 102280, 102230, 102210, 102190, 102160, 102070, 
    102020, 101990, 101940, 101870, 101820, 101780, 101720, 101660, 101620, 
    101550, 101480, 101400, 101290, 101180, 101090, 100990, 100870, 100750, 
    100670, 100750, 100870, 100930, 100950, 100920, 100960, 101050, 101050, 
    101080, 101090, 101140, 101190, 101180, 101190, 101170, 101170, 101160, 
    101150, 101130, 101130, 101100, 101080, 101060, 101040, 101010, 100990, 
    100960, 100960, 100940, 100910, 100900, 100870, 100850, 100820, 100800, 
    100750, 100730, 100720, 100710, 100700, 100680, 100670, 100650, 100630, 
    100660, 100650, 100650, 100650, 100650, 100650, 100670, 100660, 100670, 
    100690, 100680, 100670, 100710, 100700, 100670, 100690, 100690, 100690, 
    100700, 100690, 100690, 100700, 100680, 100690, 100670, 100650, 100640, 
    100620, 100610, 100610, 100610, 100610, 100600, 100600, 100600, 100580, 
    100580, 100580, 100580, 100560, 100540, 100520, 100520, 100520, 100520, 
    100520, 100520, 100510, 100490, 100450, 100420, 100390, 100400, 100410, 
    100420, 100430, 100430, 100490, 100520, 100580, 100650, 100700, 100730, 
    100730, 100800, 100840, 100880, 100910, 100940, 100960, 100960, 100970, 
    100980, 101000, 101020, 101020, 101030, 101040, 101060, 101080, 101110, 
    101110, 101130, 101160, 101160, 101150, 101150, 101130, 101140, 101150, 
    101140, 101140, 101150, 101160, 101140, 101140, 101140, 101130, 101110, 
    101090, 101060, 101040, 101040, 101030, 101000, 100980, 101000, 101000, 
    100980, 100990, 101020, 101020, 101060, 101120, 101150, 101150, 101160, 
    101170, 101150, 101150, 101160, 101140, 101140, 101140, 101120, 101120, 
    101130, 101130, 101130, 101140, 101140, 101170, 101190, 101220, 101240, 
    101240, 101230, 101210, 101180, 101160, 101130, 101100, 101060, 101010, 
    100990, 100950, 100910, 100890, 100850, 100810, 100770, 100720, 100690, 
    100670, 100610, 100590, 100570, 100550, 100520, 100490, 100450, 100420, 
    100370, 100300, 100200, 100100, 100000, 99920, 99820, 99690, 99610, 
    99520, 99480, 99390, 99270, 99250, 99200, 99160, 99120, 99110, 99080, 
    99100, 99100, 99110, 99140, 99120, 99180, 99230, 99280, 99300, 99360, 
    99420, 99510, 99640, 99770, 99870, 99960, 99990, 100080, 100170, 100220, 
    100290, 100370, 100480, 100560, 100610, 100690, 100770, 100830, 100870, 
    100930, 101010, 101070, 101150, 101210, 101230, 101260, 101280, 101290, 
    101300, 101340, 101360, 101390, 101430, 101460, 101480, 101510, 101500, 
    101500, 101450, 101410, 101350, 101290, 101240, 101210, 101180, 101150, 
    101110, 101080, 101050, 101010, 100990, 100990, 100970, 100940, 100950, 
    100960, 100980, 100990, 100970, 100940, 100910, 100870, 100840, 100800, 
    100760, 100720, 100680, 100630, 100570, 100520, 100440, 100420, 100370, 
    100320, 100250, 100210, 100160, 100080, 100010, 99940, 99900, 99920, 
    99920, 99960, 99990, 100060, 100090, 100130, 100160, 100210, 100270, 
    100350, 100450, 100510, 100550, 100590, 100610, 100700, 100760, 100820, 
    100870, 100950, 100980, 101020, 101060, 101120, 101210, 101260, 101330, 
    101370, 101400, 101440, 101450, 101480, 101540, 101600, 101650, 101680, 
    101730, 101780, 101820, 101880, 101890, 101930, 101940, 101910, 101920, 
    101970, 102020, 102080, 102130, 102170, 102220, 102260, 102280, 102310, 
    102340, 102340, 102380, 102400, 102390, 102400, 102380, 102380, 102440, 
    102540, 102470, 102480, 102480, 102520, 102530, 102550, 102530, 102530, 
    102520, 102510, 102480, 102480, 102470, 102510, 102530, 102490, 102480, 
    102500, 102450, 102530, 102540, 102560, 102520, 102480, 102440, 102450, 
    102460, 102480, 102500, 102500, 102510, 102530, 102580, 102640, 102600, 
    102670, 102710, 102750, 102770, 102800, 102810, 102810, 102840, 102870, 
    102910, 102950, 102970, 102990, 103050, 103100, 103120, 103140, 103140, 
    103140, 103170, 103180, 103180, 103180, 103180, 103200, 103180, 103170, 
    103160, 103160, 103150, 103120, 103090, 103110, 103080, 103080, 103080, 
    103060, 103060, 103050, 103030, 102970, 102960, 102960, 102950, 102920, 
    102910, 102880, 102830, 102800, 102740, 102640, 102570, 102510, 102420, 
    102350, 102290, 102270, 102230, 102190, 102180, 102170, 102180, 102190, 
    102210, 102230, 102220, 102220, 102250, 102280, 102250, 102280, 102290, 
    102280, 102250, 102270, 102230, 102180, 102160, 102150, 102120, 102130, 
    102120, 102120, 102120, 102100, 102100, 102080, 102090, 102090, 102090, 
    102080, 102080, 102090, 102110, 102130, 102130, 102130, 102130, 102110, 
    102090, 102080, 102020, 102000, 102000, 101980, 101970, 101920, 101880, 
    101870, 101820, 101800, 101760, 101740, 101690, 101670, 101680, 101680, 
    101670, 101670, 101670, 101660, 101660, 101660, 101640, 101610, 101570, 
    101540, 101540, 101540, 101510, 101470, 101450, 101430, 101410, 101380, 
    101340, 101320, 101330, 101340, 101340, 101360, 101360, 101370, 101360, 
    101330, 101320, 101320, 101330, 101280, 101270, 101260, 101270, 101310, 
    101330, 101370, 101370, 101390, 101380, 101400, 101380, 101370, 101390, 
    101380, 101390, 101440, 101480, 101500, 101500, 101530, 101530, 101540, 
    101520, 101500, 101520, 101540, 101550, 101560, 101580, 101590, 101600, 
    101620, 101660, 101670, 101670, 101680, 101680, 101680, 101680, 101690, 
    101720, 101740, 101720, 101710, 101680, 101650, 101610, 101570, 101540, 
    101500, 101450, 101420, 101380, 101370, 101320, 101280, 101260, 101240, 
    101220, 101230, 101210, 101220, 101250, 101280, 101290, 101300, 101320, 
    101360, 101390, 101430, 101450, 101490, 101550, 101590, 101640, 101710, 
    101780, 101860, 101920, 101960, 102020, 102050, 102080, 102120, 102190, 
    102260, 102310, 102370, 102410, 102460, 102500, 102540, 102570, 102590, 
    102590, 102590, 102580, 102570, 102570, 102590, 102600, 102570, 102560, 
    102550, 102530, 102540, 102510, 102500, 102490, 102490, 102480, 102470, 
    102460, 102440, 102410, 102370, 102340, 102310, 102270, 102240, 102200, 
    102130, 102090, 102050, 102040, 102000, 101960, 101920, 101880, 101840, 
    101800, 101760, 101750, 101740, 101740, 101730, 101730, 101740, 101730, 
    101720, 101750, 101750, 101760, 101760, 101740, 101740, 101740, 101770, 
    101780, 101790, 101780, 101800, 101810, 101810, 101810, 101810, 101810, 
    101830, 101870, 101880, 101880, 101870, 101870, 101890, 101880, 101860, 
    101830, 101790, 101750, 101710, 101680, 101640, 101580, 101560, 101510, 
    101500, 101460, 101430, 101380, 101340, 101300, 101280, 101300, 101300, 
    101300, 101280, 101260, 101230, 101210, 101210, 101190, 101200, 101220, 
    101260, 101350, 101410, 101470, 101550, 101590, 101620, 101640, 101700, 
    101740, 101800, 101860, 101910, 101980, 102050, 102120, 102140, 102200, 
    102250, 102280, 102300, 102320, 102330, 102350, 102360, 102350, 102380, 
    102380, 102370, 102360, 102340, 102300, 102290, 102270, 102220, 102170, 
    102130, 102090, 102050, 102000, 101930, 101900, 101830, 101790, 101710, 
    101650, 101570, 101510, 101440, 101390, 101360, 101330, 101310, 101280, 
    101280, 101280, 101310, 101340, 101350, 101350, 101360, 101390, 101410, 
    101450, 101460, 101490, 101500, 101510, 101500, 101500, 101490, 101450, 
    101430, 101400, 101400, 101390, 101370, 101340, 101310, 101270, 101260, 
    101230, 101220, 101210, 101200, 101230, 101230, 101270, 101300, 101320, 
    101330, 101350, 101380, 101370, 101360, 101350, 101350, 101370, 101370, 
    101370, 101350, 101300, 101260, 101220, 101170, 101140, 101100, 101070, 
    101040, 101010, 100980, 101000, 100990, 100960, 100910, 100860, 100790, 
    100720, 100650, 100600, 100540, 100480, 100440, 100380, 100350, 100300, 
    100290, 100270, 100270, 100250, 100210, 100180, 100150, 100120, 100100, 
    100060, 100030, 100000, 99960, 99920, 99880, 99830, 99780, 99720, 99700, 
    99700, 99720, 99730, 99760, 99780, 99840, 99890, 99920, 100040, 100130, 
    100200, 100280, 100270, 100220, 100240, 100270, 100370, 100430, 100500, 
    100570, 100680, 100810, 100890, 100940, 101050, 101150, 101210, 101230, 
    101250, 101260, 101350, 101410, 101430, 101470, 101490, 101450, 101480, 
    101470, 101490, 101470, 101490, 101430, 101430, 101410, 101390, 101370, 
    101320, 101310, 101270, 101240, 101170, 101180, 101140, 101100, 101050, 
    101030, 101010, 101020, 101010, 101010, 101030, 101040, 101050, 101070, 
    101120, 101140, 101160, 101170, 101160, 101160, 101180, 101240, 101230, 
    101200, 101210, 101210, 101210, 101180, 101140, 101110, 101080, 101030, 
    100980, 100960, 100930, 100890, 100870, 100880, 100850, 100800, 100780, 
    100740, 100690, 100660, 100670, 100640, 100570, 100590, 100590, 100590, 
    100580, 100560, 100540, 100550, 100560, 100560, 100550, 100580, 100600, 
    100650, 100690, 100780, 100860, 100940, 101000, 101060, 101140, 101220, 
    101270, 101310, 101370, 101370, 101460, 101540, 101580, 101620, 101660, 
    101680, 101670, 101730, 101740, 101730, 101750, 101780, 101800, 101830, 
    101850, 101850, 101830, 101800, 101780, 101800, 101800, 101780, 101810, 
    101830, 101810, 101780, 101760, 101710, 101710, 101710, 101690, 101690, 
    101680, 101650, 101640, 101630, 101610, 101610, 101620, 101640, 101670, 
    101680, 101680, 101670, 101710, 101720, 101730, 101750, 101790, 101820, 
    101860, 101890, 101920, 101950, 101950, 101960, 101960, 101980, 102000, 
    102070, 102090, 102150, 102180, 102200, 102230, 102220, 102210, 102230, 
    102250, 102250, 102280, 102270, 102270, 102260, 102260, 102260, 102250, 
    102210, 102200, 102200, 102190, 102170, 102170, 102190, 102200, 102180, 
    102210, 102190, 102190, 102170, 102190, 102180, 102180, 102180, 102190, 
    102200, 102210, 102220, 102220, 102220, 102220, 102230, 102240, 102260, 
    102250, 102250, 102270, 102290, 102300, 102320, 102320, 102330, 102330, 
    102330, 102310, 102300, 102310, 102300, 102280, 102260, 102240, 102230, 
    102210, 102210, 102190, 102200, 102190, 102180, 102170, 102170, 102180, 
    102180, 102170, 102150, 102160, 102160, 102140, 102140, 102140, 102130, 
    102120, 102120, 102090, 102070, 102040, 102030, 102010, 101990, 101980, 
    101990, 101970, 101950, 101960, 101950, 101910, 101910, 101940, 101940, 
    101940, 101930, 101930, 101950, 101960, 101960, 101950, 101940, 101930, 
    101920, 101910, 101910, 101910, 101880, 101880, 101890, 101890, 101880, 
    101880, 101910, 101910, 101900, 101920, 101920, 101920, 101910, 101910, 
    101910, 101920, 101900, 101880, 101860, 101860, 101870, 101860, 101850, 
    101840, 101810, 101820, 101820, 101800, 101800, 101800, 101780, 101770, 
    101770, 101780, 101770, 101760, 101750, 101740, 101740, 101710, 101690, 
    101680, 101640, 101630, 101610, 101610, 101590, 101550, 101530, 101510, 
    101490, 101460, 101430, 101400, 101370, 101350, 101350, 101340, 101330, 
    101330, 101300, 101290, 101270, 101260, 101240, 101230, 101210, 101200, 
    101200, 101200, 101190, 101180, 101160, 101110, 101090, 101070, 101110, 
    101070, 101040, 101010, 101000, 101000, 101020, 100990, 100940, 100930, 
    100920, 100910, 100890, 100870, 100890, 100900, 100900, 100900, 100880, 
    100880, 100890, 100930, 100950, 100970, 100990, 101000, 101020, 101040, 
    101070, 101110, 101120, 101130, 101160, 101180, 101170, 101200, 101230, 
    101240, 101250, 101270, 101300, 101340, 101360, 101390, 101420, 101440, 
    101440, 101500, 101560, 101590, 101620, 101640, 101670, 101730, 101750, 
    101770, 101820, 101830, 101860, 101880, 101880, 101880, 101880, 101890, 
    101890, 101910, 101890, 101890, 101890, 101880, 101870, 101850, 101840, 
    101810, 101800, 101820, 101810, 101810, 101830, 101820, 101810, 101780, 
    101760, 101760, 101760, 101720, 101680, 101660, 101670, 101640, 101620, 
    101610, 101590, 101570, 101550, 101520, 101490, 101490, 101470, 101480, 
    101490, 101480, 101490, 101490, 101490, 101500, 101520, 101520, 101540, 
    101540, 101580, 101610, 101640, 101670, 101700, 101710, 101730, 101740, 
    101750, 101770, 101790, 101800, 101820, 101830, 101860, 101900, 101950, 
    101990, 101990, 101990, 102020, 102030, 102030, 102040, 102040, 102040, 
    102050, 102050, 102070, 102080, 102080, 102040, 102040, 102040, 102030, 
    102020, 102000, 102010, 102020, 102030, 102040, 102020, 102030, 102030, 
    102000, 102020, 102010, 102000, 101970, 101970, 101960, 102000, 102000, 
    102010, 102030, 102040, 102060, 102060, 102080, 102120, 102160, 102210, 
    102270, 102320, 102380, 102390, 102430, 102440, 102460, 102440, 102470, 
    102460, 102500, 102530, 102510, 102540, 102550, 102570, 102560, 102570, 
    102590, 102590, 102640, 102630, 102660, 102690, 102700, 102720, 102770, 
    102780, 102770, 102830, 102850, 102810, 102790, 102820, 102820, 102790, 
    102820, 102790, 102770, 102710, 102690, 102640, 102590, 102490, 102470, 
    102420, 102320, 102260, 102200, 102160, 102110, 102060, 101990, 101900, 
    101850, 101840, 101820, 101790, 101730, 101740, 101680, 101700, 101690, 
    101680, 101690, 101680, 101660, 101670, 101630, 101590, 101590, 101570, 
    101550, 101520, 101480, 101410, 101310, 101210, 101190, 101100, 100930, 
    100800, 100720, 100640, 100580, 100510, 100490, 100470, 100430, 100440, 
    100400, 100430, 100460, 100520, 100600, 100640, 100590, 100650, 100650, 
    100660, 100630, 100670, 100660, 100640, 100620, 100590, 100550, 100530, 
    100490, 100490, 100450, 100440, 100410, 100410, 100420, 100390, 100420, 
    100450, 100500, 100510, 100520, 100560, 100590, 100610, 100650, 100670, 
    100700, 100740, 100780, 100790, 100770, 100790, 100790, 100810, 100820, 
    100840, 100860, 100900, 100930, 100930, 100950, 100960, 100970, 100960, 
    100960, 101020, 101060, 101040, 101100, 101130, 101170, 101180, 101170, 
    101200, 101210, 101210, 101200, 101200, 101230, 101230, 101220, 101240, 
    101280, 101280, 101270, 101260, 101320, 101320, 101370, 101370, 101390, 
    101440, 101450, 101440, 101430, 101460, 101530, 101550, 101580, 101580, 
    101580, 101610, 101690, 101740, 101790, 101850, 101910, 101960, 101980, 
    102020, 102060, 102070, 102110, 102180, 102190, 102240, 102260, 102290, 
    102310, 102300, 102290, 102290, 102270, 102250, 102260, 102220, 102220, 
    102190, 102170, 102150, 102100, 102080, 102040, 102030, 101980, 101980, 
    102000, 102010, 102040, 102050, 102040, 101980, 101950, 101890, 101830, 
    101810, 101760, 101740, 101690, 101660, 101630, 101610, 101560, 101530, 
    101480, 101440, 101400, 101350, 101330, 101290, 101260, 101260, 101260, 
    101270, 101260, 101270, 101290, 101260, 101250, 101230, 101230, 101230, 
    101230, 101250, 101260, 101250, 101230, 101280, 101290, 101320, 101320, 
    101360, 101410, 101400, 101450, 101490, 101510, 101540, 101570, 101610, 
    101630, 101640, 101640, 101650, 101650, 101680, 101680, 101710, 101720, 
    101720, 101710, 101720, 101710, 101720, 101700, 101710, 101700, 101700, 
    101730, 101740, 101700, 101710, 101690, 101670, 101600, 101610, 101600, 
    101560, 101490, 101430, 101380, 101380, 101340, 101270, 101290, 101310, 
    101320, 101330, 101330, 101360, 101320, 101350, 101370, 101410, 101390, 
    101390, 101380, 101360, 101350, 101340, 101340, 101340, 101340, 101340, 
    101350, 101360, 101350, 101340, 101330, 101320, 101280, 101260, 101250, 
    101240, 101240, 101220, 101200, 101200, 101210, 101220, 101260, 101250, 
    101260, 101270, 101270, 101300, 101340, 101410, 101450, 101510, 101560, 
    101600, 101600, 101640, 101710, 101740, 101740, 101780, 101830, 101860, 
    101920, 101960, 102010, 102030, 102030, 102040, 102030, 102010, 101970, 
    101960, 101930, 101900, 101880, 101820, 101770, 101730, 101680, 101590, 
    101530, 101450, 101380, 101270, 101180, 101100, 101050, 101000, 100940, 
    100850, 100800, 100760, 100730, 100680, 100630, 100590, 100570, 100540, 
    100510, 100480, 100470, 100440, 100370, 100320, 100290, 100260, 100220, 
    100140, 100100, 100120, 100100, 100110, 100130, 100160, 100190, 100170, 
    100160, 100140, 100230, 100260, 100270, 100300, 100340, 100370, 100390, 
    100470, 100480, 100540, 100620, 100670, 100720, 100740, 100770, 100780, 
    100860, 100920, 100940, 100990, 101010, 101010, 101060, 101070, 101080, 
    101060, 101050, 101060, 101060, 101080, 101080, 101090, 101120, 101090, 
    101090, 101090, 101070, 101080, 101070, 101070, 101070, 101050, 101070, 
    101060, 101040, 101020, 101010, 100990, 101000, 100960, 100930, 100930, 
    100940, 100940, 100950, 100960, 100950, 100940, 100920, 100930, 100930, 
    100950, 100960, 100960, 100970, 100990, 101000, 101040, 101060, 101090, 
    101090, 101080, 101080, 101100, 101100, 101110, 101140, 101140, 101150, 
    101150, 101140, 101140, 101140, 101150, 101150, 101170, 101170, 101170, 
    101180, 101210, 101240, 101260, 101280, 101290, 101310, 101310, 101310, 
    101330, 101330, 101330, 101320, 101340, 101340, 101350, 101360, 101360, 
    101350, 101350, 101360, 101350, 101350, 101350, 101350, 101360, 101380, 
    101400, 101400, 101390, 101380, 101360, 101350, 101330, 101300, 101270, 
    101260, 101230, 101210, 101170, 101130, 101110, 101100, 101080, 101040, 
    101020, 100980, 100920, 100880, 100840, 100810, 100780, 100740, 100700, 
    100660, 100620, 100570, 100550, 100510, 100460, 100400, 100380, 100370, 
    100320, 100290, 100260, 100230, 100200, 100150, 100110, 100080, 100080, 
    100070, 100070, 100070, 100070, 100040, 100020, 100020, 100000, 100000, 
    99990, 99980, 99960, 99970, 99960, 99960, 99950, 99950, 99950, 99930, 
    99900, 99890, 99900, 99900, 99900, 99890, 99910, 99910, 99910, 99900, 
    99890, 99890, 99900, 99900, 99890, 99880, 99870, 99850, 99840, 99810, 
    99800, 99790, 99790, 99770, 99770, 99780, 99800, 99850, 99880, 99920, _, 
    _, 100060, 100120, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 101330, 101370, _, 101400, 101420, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 101510, 101480, 101450, 101440, 101440, _, _, _, 
    101370, _, 101380, 101370, 101400, 101420, 101400, 101410, _, _, _, 
    101400, 101370, 101390, 101400, 101430, 101480, 101530, 101590, 101670, 
    101710, 101700, 101750, 101800, 101800, 101810, 101850, 101950, 101950, 
    102000, 102040, 102070, 102120, 102150, 102160, 102140, 102110, _, _, _, 
    102150, 102170, 102170, 102210, 102200, 102170, 102160, 102100, 102110, 
    102100, 102020, 102020, 101990, 101950, 101910, _, _, _, _, 101640, 
    101530, 101480, 101440, 101360, 101300, 101250, 101230, 101220, 101240, 
    101170, 101140, 101070, 101060, 101050, _, _, _, _, _, _, 101110, 101140, 
    101160, _, 101240, _, 101320, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 102040, 102070, _, 102080, 102090, 102060, _, _, _, _, _, 102050, 
    102030, 102030, 102020, 102010, 101960, 101930, 101940, 101920, 101910, 
    _, _, _, _, _, _, _, _, 101860, 101840, _, 101790, 101780, _, 101790, 
    101790, 101780, 101770, _, _, 101710, 101680, _, _, 101590, 101580, 
    101560, 101530, 101500, _, 101430, 101410, _, _, _, _, 101240, 101230, 
    101190, 101170, 101140, 101110, 101090, 101090, 101100, 101060, _, _, 
    101000, 101020, 101020, 101000, _, 101000, _, _, _, _, _, _, _, 100870, 
    100860, 100880, 100870, 100850, 100820, 100780, 100780, 100790, 100790, 
    100760, 100750, 100760, 100750, 100740, 100730, 100740, 100730, 100730, 
    100720, 100720, 100680, 100660, 100690, 100700, 100690, 100690, 100680, 
    100650, 100640, 100620, 100620, 100620, 100610, 100610, 100600, 100600, 
    100620, 100620, 100590, 100520, 100530, 100530, 100530, 100540, 100520, 
    100550, 100590, 100640, 100640, 100720, 100760, 100790, 100840, 100870, 
    100900, 100920, 100950, 100900, 100900, 100910, 100860, 100910, 100950, 
    100940, 100940, 100930, 100920, 100900, 100890, 100870, 100850, 100840, 
    100910, 100930, 100940, 100910, 100930, 100970, 100970, 100960, 100980, 
    100920, 100930, 100930, 100930, 100920, 100910, 100890, 100840, 100780, 
    100720, 100710, 100660, 100650, 100660, 100640, 100640, 100640, 100650, 
    100640, 100600, 100580, 100570, 100550, 100530, 100500, 100470, 100460, 
    100430, 100440, 100440, 100420, 100390, 100390, 100360, 100380, 100410, 
    100440, 100470, 100490, 100490, 100410, 100390, 100400, _, _, 100520, 
    100520, _, _, _, _, _, _, _, _, _, 100740, 100770, 100800, 100830, 
    100880, 100910, 100970, 101000, 101030, 101070, 101090, 101120, 101140, 
    101160, 101150, 101170, 101210, _, _, _, _, _, _, _, 101240, 101190, _, 
    _, 101190, 101170, 101170, 101220, _, 101190, 101160, 101150, 101140, _, 
    101080, 101060, 101060, 101060, _, _, 100960, 100970, 100970, 100970, 
    100920, 100890, 100880, 100840, _, 100790, 100760, 100710, 100700, _, 
    100630, 100590, 100550, _, _, _, _, _, _, _, _, _, _, _, _, _, 99580, 
    99550, 99550, 99570, 99620, 99680, 99730, 99820, 99860, 99890, 99930, _, 
    _, _, _, _, 99990, 100020, _, 100110, 100170, 100230, 100250, 100280, _, 
    _, 100410, 100420, 100470, 100510, 100540, 100560, _, 100620, _, _, _, _, 
    _, _, _, _, 100660, 100660, 100670, _, 100730, 100730, 100730, 100740, _, 
    100730, _, _, 100960, 101020, 101050, 101070, 101130, 101170, 101180, 
    101220, _, _, _, 101420, 101510, 101550, 101600, 101660, 101680, 101690, 
    _, _, _, 101790, 101830, 101850, 101880, 101930, 101940, 101960, 101970, 
    101960, _, _, 101970, 101980, 102000, 102010, 102000, 102000, 102010, 
    102000, 101980, _, 101960, 101960, 101970, 101960, 101960, 101980, 
    101990, 102010, _, 102030, 102030, 102010, 102000, 102000, 102020, 
    102020, 102020, _, _, _, _, _, 101940, 101930, 101840, 101810, 101730, 
    101730, 101700, 101720, 101710, 101680, 101700, _, _, 101600, _, 101560, 
    101540, 101510, 101490, 101430, 101390, 101350, _, 101260, 101210, 
    101140, 101100, 101040, 101020, 100990, 100990, _, 100970, 100940, 
    100900, 100860, 100790, 100720, 100640, 100550, _, 100430, 100390, _, 
    100280, 100240, _, _, 100140, 100130, 100120, _, 100140, 100170, 100190, 
    100240, 100290, 100360, 100370, 100380, 100400, 100390, 100370, 100380, 
    100390, 100400, 100390, 100420, 100460, 100460, 100480, 100500, 100540, 
    100570, 100630, 100630, 100650, 100690, 100730, 100800, 100850, 100860, 
    100880, 100910, 100890, 100900, 100890, 100870, 100820, 100730, 100720, 
    100670, 100620, 100570, 100540, 100500, 100470, 100440, 100420, 100440, 
    100470, 100490, 100490, 100490, 100490, 100510, 100520, 100500, 100500, 
    100480, 100470, 100440, 100450, 100450, 100440, 100500, 100530, 100490, 
    100510, 100490, 100480, 100490, 100490, _, 100470, 100470, 100450, 
    100450, 100450, 100470, 100500, 100530, 100540, 100580, 100610, 100650, 
    100700, 100740, 100820, 100900, 100960, 100970, 101010, 100980, 101090, 
    101190, 101200, 101250, 101320, 101360, _, 101410, 101460, 101500, 
    101550, 101550, 101570, 101580, 101580, 101590, _, _, _, 101580, 101590, 
    101600, 101590, 101580, 101560, 101550, 101560, _, _, _, 101490, 101490, 
    101500, 101490, 101480, 101450, 101440, 101410, 101390, _, _, _, _, _, _, 
    _, _, _, _, 101230, 101210, _, 101200, 101190, 101210, 101220, 101240, 
    101230, _, _, _, _, _, _, _, _, 101200, 101220, 101230, 101230, 101210, 
    101210, 101210, 101180, _, _, 101160, 101170, 101160, 101180, 101190, 
    101180, 101190, 101190, _, _, _, _, _, _, 101070, 101060, 101020, 101020, 
    100990, 100960, 100920, 100880, _, _, _, _, _, 100610, 100580, 100520, 
    100460, 100390, 100320, 100240, _, _, _, _, 99890, 99850, 99810, 99770, 
    99730, 99700, 99680, 99660, 99650, _, _, _, _, _, _, 99910, 99950, 
    100020, 100070, 100180, 100290, 100310, 100360, _, _, _, _, 100640, 
    100660, 100700, 100740, 100740, 100760, 100760, 100790, _, 100850, 
    100920, 100920, 100930, 100950, 100960, 100950, 100950, _, _, 100900, 
    100880, 100850, 100830, 100800, 100760, 100700, 100610, _, _, 100440, 
    100390, 100330, 100310, 100260, 100220, 100150, 100070, _, 99890, 99820, 
    99760, 99750, 99730, 99680, 99680, 99650, _, _, _, _, _, _, 99690, 99700, 
    _, 99750, 99770, _, 99800, 99830, 99840, 99850, 99850, 99840, 99800, 
    99790, 99800, 99790, 99780, _, _, _, _, _, _, _, _, 99790, 99780, 99780, 
    99780, 99770, 99760, 99760, 99750, _, 99670, 99680, 99640, 99650, 99670, 
    99700, 99730, 99740, _, _, _, _, 100050, 100120, 100210, 100310, 100350, 
    100430, 100540, 100610, _, 100770, 100900, 100950, 101010, 101060, 
    101090, 101100, 101110, _, _, _, 100960, 100920, 100860, 100770, 100670, 
    100560, 100460, 100340, _, _, _, 99950, 99830, 99750, 99660, 99540, 
    99370, 99230, 99040, 98840, _, _, _, 98300, 98260, 98260, 98200, 98210, 
    98230, 98230, 98270, _, 98360, 98450, 98500, 98650, 98790, 98870, 99030, 
    99160, 99250, 99320, 99370, 99470, 99520, 99620, 99680, _, _, _, 100030, 
    100120, 100210, 100320, 100430, 100590, 100710, 100830, _, 101040, 
    101180, 101320, 101420, 101470, 101550, 101570, 101600, 101610, 101630, 
    _, _, _, _, 101630, 101600, 101530, 101480, 101420, 101350, 101250, 
    101170, _, _, _, 100870, 100800, 100730, 100650, 100550, 100490, 100380, 
    100360, _, _, _, 100140, 100110, 100040, 100030, 99980, 99920, 99850, 
    99790, 99750, _, _, _, 99480, 99450, 99390, 99330, 99260, 99280, 99320, 
    99320, _, _, _, 99300, 99280, 99270, 99230, 99210, 99170, 99140, 99110, 
    _, _, _, 99100, 99170, 99210, 99250, 99260, 99240, 99270, 99350, _, _, _, 
    _, _, _, _, _, 99260, 99240, 99200, 99170, 99160, 99150, 99130, 99130, _, 
    _, 99170, 99210, 99240, 99290, 99320, 99370, 99420, 99480, _, _, _, _, _, 
    _, _, _, _, _, 100120, 100190, 100230, _, _, _, 100480, 100500, 100470, 
    _, 100540, _, _, 100630, _, 100670, _, _, _, 100740, 100750, 100760, 
    100760, _, _, 100800, _, _, 100880, 100930, _, 101080, 101160, _, _, _, 
    _, _, _, _, _, _, 101750, _, _, _, _, _, _, _, 102050, 102050, 102070, 
    102080, 102090, 102150, _, _, _, _, _, 102220, 102220, _, 102160, 102150, 
    102110, 102090, 102100, _, _, 102010, 102000, 101980, _, 101910, 101910, 
    101880, 101900, _, _, 101910, 101900, 101900, 101900, 101890, 101900, 
    101880, _, 101810, 101800, 101800, 101800, 101720, 101730, 101650, 
    101590, _, 101580, _, 101460, 101460, 101450, 101430, 101430, 101420, 
    101400, 101350, 101300, 101280, 101250, 101240, 101220, 101220, _, _, 
    101190, 101180, _, _, 101160, 101120, 101090, 101080, _, _, 101010, 
    101010, 100990, 100950, 100910, 100850, 100800, 100720, 100660, _, _, _, 
    100330, 100270, 100210, _, _, _, 99830, 99690, 99560, 99450, 99390, 
    99330, 99280, _, 99130, 99050, 98950, 98850, 98730, 98680, 98580, 98610, 
    _, _, _, 98370, 98350, 98300, _, 98210, 98230, 98200, 98200, 98170, 
    98140, 98160, _, 98220, _, 98250, _, _, _, _, _, 98470, 98500, _, 98560, 
    _, 98640, _, 98720, 98700, _, 98810, 98830, 98870, 98900, _, _, _, _, _, 
    _, 99070, _, 99090, _, 99130, _, 99230, _, _, _, 99460, 99520, 99520, 
    99600, 99650, 99700, 99800, 99860, _, 99950, 99980, 100020, _, 100190, 
    100240, 100270, 100340, _, _, 100490, 100510, 100540, 100580, 100620, 
    100660, 100710, _, 100790, _, _, _, 100930, 100980, 101010, 101050, 
    101060, 101080, 101110, 101090, _, _, 101090, _, _, 101040, 101110, 
    101170, _, 101210, _, _, _, _, _, _, _, _, 101420, 101480, 101510, 
    101490, 101470, 101500, 101510, _, 101510, 101500, 101490, 101470, 
    101430, 101390, 101390, _, _, _, _, 101030, 100910, _, 100720, 100640, _, 
    100470, 100360, 100260, 100170, _, 99990, _, 99950, 99940, 99930, 99960, 
    _, _, 99950, 99950, 99970, _, _, _, 100290, 100420, 100530, 100640, 
    100730, 100870, 101040, 101200, _, 101420, _, 101620, _, _, 101920, _, _, 
    _, 102320, 102380, 102380, 102380, 102410, 102420, 102390, 102400, 
    102290, _, 102180, _, 102130, _, 102020, 101940, 101860, 101830, _, _, _, 
    101560, 101560, 101610, 101590, 101570, 101610, 101590, 101610, _, _, _, 
    _, _, _, _, _, _, _, 101770, 101750, 101700, 101660, 101580, 101500, 
    101320, 101120, _, _, 100810, _, 100860, 100970, _, 101230, 101360, _, _, 
    _, _, 101810, _, 101890, 101900, 101950, 102010, _, _, 102020, _, _, 
    101970, _, 102020, 101950, 101970, 101940, 101920, 101880, _, _, _, 
    102030, _, _, _, 102290, 102380, 102450, 102550, 102690, 102770, 102850, 
    102930, 102960, _, _, _, _, 103310, 103330, 103360, 103370, 103370, 
    103400, 103400, 103430, _, 103470, 103450, 103440, 103410, 103400, 
    103380, 103360, 103360, 103360, 103340, 103330, 103300, 103280, 103250, 
    103230, 103200, 103160, _, _, _, _, 102970, 102920, _, 102810, 102740, 
    102690, 102620, 102570, 102510, 102470, 102390, _, _, _, _, 102120, 
    102070, 101980, 101930, 101860, 101810, 101740, 101700, _, _, 101610, 
    101590, 101590, 101600, 101620, 101640, 101690, 101710, _, _, 101740, 
    101770, 101760, 101750, 101720, 101680, 101660, 101630, _, _, 101460, 
    101380, 101350, 101340, 101330, 101330, 101330, 101350, _, _, 101330, 
    101330, 101350, 101360, 101370, 101360, 101390, 101410, 101410, 101410, 
    101410, 101400, 101380, 101360, 101370, 101350, 101340, 101350, _, _, _, 
    _, 101430, 101430, 101420, 101410, 101380, 101380, _, _, 101400, 101420, 
    101410, 101380, 101380, 101390, 101380, 101390, _, _, 101410, 101400, 
    101420, 101440, 101430, 101410, _, 101420, 101390, _, _, 101460, 101440, 
    101420, 101490, 101510, 101530, 101560, 101570, _, _, _, _, 101610, 
    101640, 101650, 101690, 101720, 101730, 101810, 101820, _, _, _, 101820, 
    101810, 101810, 101840, 101870, 101920, 101910, 101910, 101930, _, _, 
    101940, 101930, 101920, 101850, 101830, 101820, 101750, 101750, _, 
    101700, 101690, 101700, 101710, 101710, 101660, 101620, 101620, _, _, _, 
    _, _, 101690, 101670, 101660, 101670, 101660, 101650, 101670, 101690, _, 
    _, 101720, 101720, _, 101720, 101720, 101720, 101740, 101740, _, _, _, 
    101800, 101790, 101780, 101740, 101720, 101660, 101530, 101420, _, _, 
    101020, 100700, 100520, 100340, 100260, 100280, 100310, 100550, 100790, 
    _, _, 101170, 101240, 101290, 101340, 101360, 101400, 101440, 101450, _, 
    _, _, _, 101550, 101570, 101590, 101630, 101660, 101660, 101680, 101720, 
    _, _, _, _, _, _, _, _, _, 101790, 101770, 101740, 101710, 101680, 
    101680, 101670, 101610, 101610, 101610, 101610, 101600, 101570, 101580, 
    101580, 101570, _, _, _, _, _, _, 101600, 101590, 101600, 101580, 101560, 
    101530, 101530, 101530, _, _, 101530, 101550, 101570, 101570, 101600, 
    101600, 101590, 101620, _, _, 101600, 101600, 101590, 101600, 101610, 
    101630, 101640, 101660, 101650, 101650, 101680, 101700, 101700, 101720, 
    101770, _, 101840, 101870, 101900, 101920, 101920, 101920, _, _, _, _, _, 
    _, 101950, 101930, 101890, 101860, 101820, 101770, 101720, 101690, _, _, 
    _, _, _, 101620, 101570, 101560, 101510, 101440, 101430, 101420, 101380, 
    _, _, _, _, _, _, _, _, _, 101120, 101100, 101070, 101060, 101040, 
    101040, 101040, 101080, _, _, _, 101140, 101150, 101180, 101190, 101220, 
    101240, 101230, 101250, _, _, _, _, 101060, 101010, 100950, 100920, 
    100890, 100920, 100910, 100900, _, _, 100900, 100910, 100940, 100920, 
    100960, 101030, 101030, 101040, _, _, _, _, 100940, 100910, 100900, 
    100880, 100860, 100880, 100890, _, _, _, 100950, 100990, 100990, 100980, 
    101010, 101050, 101050, 101100, _, _, _, 101220, 101240, 101230, 101200, 
    101160, 101140, 101100, 101050, _, _, 100960, 100940, 100930, 100880, 
    100830, 100770, 100720, 100670, _, _, _, 100500, 100440, 100380, 100300, 
    100270, 100230, 100180, 100170, _, _, _, _, 100130, 100140, 100220, 
    100240, 100250, 100230, 100160, 100200, _, _, _, _, _, 100430, 100480, 
    100510, 100570, _, 100630, 100650, 100680, 100700, 100750, 100820, 
    100900, 100960, 101020, 101060, _, 101130, 101150, 101190, 101210, 
    101230, 101250, 101260, _, _, _, _, _, _, _, _, 101350, 101340, 101340, 
    101360, 101350, 101360, 101380, 101380, 101380, 101360, 101360, 101350, 
    101330, 101310, 101320, 101310, 101310, 101320, 101310, 101300, 101310, 
    101310, 101290, 101290, 101280, 101280, 101290, 101330, 101350, 101380, 
    101430, 101460, 101500, 101510, 101520, 101540, 101550, 101570, 101580, 
    101600, 101610, 101640, 101650, 101660, 101660, 101670, 101690, 101710, 
    101710, 101690, 101680, 101690, 101700, 101690, 101680, 101680, 101660, 
    101620, 101580, 101550, 101500, 101470, 101420, 101370, 101320, 101360, 
    101360, 101370, 101370, 101380, 101320, 101300, 101360, 101350, 101330, 
    101330, 101340, 101290, 101320, 101340, 101260, 101310, 101310, 101300, 
    101270, 101250, 101190, 101170, 101130, 101060, 101050, 101010, 100950, 
    100890, 100860, 100770, 100750, 100710, 100670, 100620, 100580, 100540, 
    100490, 100430, 100410, 100420, 100350, 100300, 100250, 100240, 100200, 
    100170, 100090, 100140, 100150, 100120, 100050, 100020, 99980, 99940, 
    99890, 99860, 99860, 99830, 99830, 99810, 99860, 99890, 99860, 99890, 
    99870, 99930, 99930, 99940, 99980, 100040, 100210, 100240, 100250, 
    100300, 100280, 100290, 100390, 100300, 100350, 100410, 100440, 100430, 
    100390, 100440, 100460, 100480, 100490, 100470, 100490, 100450, 100420, 
    100400, 100360, 100360, 100320, 100300, 100230, 100190, 100150, 100070, 
    100030, 99990, 99920, 99890, 99840, 99810, 99780, 99760, 99760, 99790, 
    99790, 99790, 99800, 99780, 99790, 99810, 99840, 99900, 99980, 100070, 
    100200, 100260, 100350, 100430, 100500, 100530, 100610, 100620, 100690, 
    100730, 100790, 100840, 100900, 100950, 100960, 100950, 100990, 101030, 
    101060, 101050, 101060, 101100, 101120, 101150, 101170, 101190, 101180, 
    101180, 101200, 101200, 101150, 101200, 101170, 101130, 101150, 101130, 
    101120, 101110, 101090, 101010, 100970, 100950, 100860, 100800, 100700, 
    100560, 100480, 100380, 100230, 100060, 99770, 99570, 99480, 99490, 
    99300, 99200, 98950, 98750, 98680, 98620, 98530, 98340, 98300, 98300, 
    98270, 98340, 98330, 98290, 98230, 98360, 98550, 98660, 98800, 98860, 
    98900, 98950, 99080, 99150, 99220, 99300, 99370, 99520, 99610, 99690, 
    99730, 99770, 99980, 99970, 99860, 99990, 100040, 100110, 100150, 100170, 
    100170, 100150, 100130, 100110, 100130, 100160, 100080, 100110, 100150, 
    100160, 100160, 100190, 100220, 100260, 100280, 100320, 100360, 100360, 
    100390, 100440, 100440, 100450, 100460, 100500, 100500, 100540, 100580, 
    100630, 100620, 100630, 100650, 100630, 100640, 100700, 100730, 100730, 
    100810, 100880, 100990, 101050, 101110, 101130, 101160, 101150, 101190, 
    101250, 101280, 101290, 101350, 101370, 101380, 101400, 101450, 101500, 
    101530, 101540, 101580, 101620, 101650, 101670, 101720, 101800, 101850, 
    101880, 101880, 101910, 101860, 101820, 101940, 101970, 101930, 101910, 
    101980, 101990, 101990, 102000, 102060, 102050, 102090, 102160, 102190, 
    102180, 102130, 102080, 102100, 102120, 102160, 102180, 102160, 102160, 
    102190, 102290, 102280, 102270, 102230, 102200, 102210, 102330, 102390, 
    102450, 102480, 102480, 102500, 102540, 102550, 102550, 102510, 102520, 
    102560, 102550, 102540, 102530, 102590, 102670, 102600, 102560, 102530, 
    102480, 102510, 102460, 102430, 102380, 102320, 102230, 102120, 102030, 
    101890, 101770, 101580, 101400, 101210, 101050, 100840, 100730, 100570, 
    100400, 100230, 100150, 100060, 100030, 100110, 100050, 100060, 100070, 
    100060, 100030, 100040, 100020, 100050, 100070, 100070, 100040, 100120, 
    100210, 100350, 100450, 100580, 100770, 100910, 100940, 100940, 100930, 
    100920, 100870, 100910, 100890, 100870, 100910, 100940, 100940, 100970, 
    101040, 101060, 101130, 101110, 101080, 101040, 101030, 100930, 100860, 
    100810, 100740, 100650, 100610, 100500, 100470, 100380, 100290, 100290, 
    100230, 100230, 100170, 100170, 100100, 100110, 100090, 100030, 100030, 
    100130, 100150, 100090, 100040, 100080, 100050, 100030, 100080, 100070, 
    100040, 100030, 100080, 100110, 100130, 100110, 100130, 100110, 100140, 
    100220, 100370, 100390, 100490, 100530, 100590, 100610, 100610, 100650, 
    100670, 100710, 100710, 100760, 100790, 100820, 100850, 100890, 100950, 
    101020, 101090, 101160, 101230, 101290, 101280, 101370, 101440, 101510, 
    101570, 101580, 101640, 101580, 101590, 101610, 101640, 101680, 101740, 
    101770, 101830, 101900, 101930, 101990, 101970, 102020, 101960, 102090, 
    102060, 102060, 102030, 102000, 102000, 102010, 102010, 101990, 101980, 
    101890, 101820, 101710, 101710, 101620, 101560, 101510, 101500, 101440, 
    101480, 101450, 101500, 101440, 101430, 101470, 101420, 101500, 101500, 
    101530, 101580, 101550, 101520, 101500, 101530, 101510, 101480, 101390, 
    101280, 101280, 101170, 100990, 100960, 100970, 100920, 100830, 100800, 
    100750, 100730, 100690, 100680, 100640, 100650, 100630, 100630, 100650, 
    100650, 100650, 100610, 100540, 100520, 100500, 100530, 100490, 100440, 
    100470, 100450, 100410, 100360, 100300, 100260, 100180, 100070, 99950, 
    99840, 99730, 99610, 99510, 99440, 99320, 99280, 99370, 99360, 99500, 
    99670, 99840, 99950, 100050, 100130, 100200, 100230, 100240, 100270, 
    100310, 100330, 100330, 100410, 100410, 100410, 100490, 100510, 100570, 
    100610, 100630, 100730, 100760, 100800, 100810, 100820, 100890, 100950, 
    101000, 101010, 101020, 101040, 101110, 101190, 101200, 101220, 101210, 
    101200, 101190, 101190, 101230, 101210, 101250, 101240, 101240, 101300, 
    101290, 101260, 101300, 101290, 101250, 101220, 101200, 101170, 101190, 
    101200, 101160, 101160, 101120, 101070, 101010, 100980, 100870, 100830, 
    100760, 100620, 100460, 100370, 100320, 100250, 100210, 100100, 100060, 
    100010, 99950, 99870, 99840, 99820, 99760, 99740, 99690, 99630, 99600, 
    99550, 99490, 99480, 99410, 99370, 99390, 99380, 99380, 99370, 99410, 
    99460, 99510, 99550, 99580, 99610, 99620, 99610, 99610, 99600, 99600, 
    99600, 99630, 99600, 99620, 99660, 99630, 99660, 99720, 99800, 99930, 
    100080, 100220, 100410, 100580, 100750, 100880, 101000, 101150, 101280, 
    101430, 101560, 101670, 101770, 101850, 101940, 102010, 102220, 102300, 
    102360, 102470, 102580, 102710, 102770, 102790, 102840, 102900, 102950, 
    103010, 103040, 103060, 103090, 103110, 103160, 103200, 103200, 103200, 
    103240, 103280, 103270, 103270, 103260, 103250, 103220, 103180, 103160, 
    103160, 103150, 103090, 103070, 103030, 103040, 102970, 102910, 102870, 
    102850, 102810, 102780, 102770, 102760, 102750, 102780, 102780, 102810, 
    102830, 102850, 102870, 102890, 102900, 102910, 102930, 102930, 102980, 
    102980, 103030, 103030, 103010, 103080, 103060, 103070, 103020, 103000, 
    102840, 102890, 102980, 103030, 103020, 103010, 102930, 102870, 102770, 
    102670, 102620, 102600, 102590, 102470, 102300, 102140, 102180, 102160, 
    102350, 102160, 102200, 102130, 102140, 102070, 102050, 101960, 101850, 
    101650, 101690, 101750, 101650, 101740, 101720, 101700, 101810, 101820, 
    101730, 101780, 101810, 101800, 101820, 101890, 101940, 101970, 102010, 
    102030, 102020, 102040, 102030, 101980, 101940, 101880, 101880, 101820, 
    101750, 101720, 101660, 101600, 101530, 101510, 101500, 101440, 101390, 
    101380, 101350, 101370, 101340, 101330, 101290, 101200, 101180, 101160, 
    101170, 101150, 101150, 101130, 101120, 101070, 101050, 101030, 100980, 
    100900, 100830, 100790, 100700, 100620, 100580, 100460, 100380, 100300, 
    100140, 99980, 100020, 99900, 99800, 99600, 99450, 99260, 99140, 99050, 
    98890, 98750, 98590, 98370, 98310, 97940, 98070, 97950, 97790, 97660, 
    97360, 97260, 97230, 97180, 97220, 97100, 96990, 97150, 97280, 97320, 
    97360, 97410, 97470, 97520, 97590, 97600, 97660, 97700, 97740, 97660, 
    97760, 98150, 98290, 98290, 98310, 98350, 98420, 98400, 98450, 98550, 
    98590, 98640, 98680, 98700, 98690, 98730, 98790, 98740, 98800, 98890, 
    98830, 98880, 98850, 98820, 98780, 98690, 98640, 98520, 98410, 98400, 
    98270, 98260, 98210, 98170, 98150, 98110, 98080, 98110, 98120, 98190, 
    98290, 98400, 98470, 98490, 98530, 98510, 98560, 98610, 98640, 98660, 
    98730, 98780, 98800, 98840, 98860, 98900, 98940, 98960, 98990, 99000, 
    99020, 99040, 99070, 99110, 99120, 99150, 99160, 99190, 99240, 99280, 
    99320, 99360, 99370, 99390, 99410, 99450, 99480, 99500, 99530, 99550, 
    99600, 99610, 99620, 99610, 99610, 99620, 99580, 99570, 99520, 99460, 
    99410, 99340, 99240, 99190, 99060, 98970, 98880, 98760, 98570, 98380, 
    98180, 98010, 97860, 97740, 97630, 97570, 97430, 97340, 97340, 97280, 
    97220, 97140, 97130, 97100, 97050, 97050, 97040, 97060, 97070, 97080, 
    97100, 97150, 97160, 97190, 97260, 97320, 97400, 97470, 97530, 97570, 
    97650, 97690, 97720, 97750, 97780, 97820, 97840, 97910, 97920, 97940, 
    97990, 98020, 98020, 98090, 98090, 98070, 98080, 98070, 98150, 98210, 
    98290, 98310, 98390, 98440, 98470, 98530, 98530, 98560, 98580, 98600, 
    98650, 98690, 98760, 98800, 98850, 98850, 98890, 98960, 98970, 99020, 
    99060, 99100, 99100, 99090, 99070, 99080, 98950, 98970, 98980, 98990, 
    99000, 98980, 98990, 99000, 98970, 99000, 98960, 99000, 99010, 99010, 
    98990, 98980, 98950, 98900, 98840, 98820, 98790, 98790, 98780, 98810, 
    98770, 98730, 98700, 98590, 98530, 98470, 98380, 98330, 98270, 98210, 
    98200, 98220, 98210, 98160, 98160, 98150, 98110, 98050, 98030, 98050, 
    98020, 97980, 97940, 97880, 97900, 97920, 97940, 97980, 97970, 97970, 
    97990, 98000, 98040, 98080, 98140, 98190, 98240, 98280, 98250, 98210, 
    98170, 98170, 98250, 98330, 98390, 98450, 98530, 98620, 98730, 98780, 
    98840, 98860, 98900, 98960, 98970, 99070, 99090, 99120, 99160, 99190, 
    99220, 99230, 99230, 99220, 99200, 99200, 99140, 99130, 99100, 99100, 
    99110, 99130, 99110, 99120, 99100, 99120, 99130, 99150, 99150, 99160, 
    99190, 99200, 99200, 99190, 99190, 99230, 99210, 99200, 99190, 99180, 
    99190, 99190, 99170, 99190, 99190, 99230, 99230, 99270, 99230, 99280, 
    99320, 99350, 99400, 99430, 99440, 99440, 99530, 99560, 99660, 99680, 
    99710, 99720, 99760, 99810, 99840, 99870, 99940, 99920, 99970, 100000, 
    100050, 100090, 100090, 100100, 100090, 100090, 100130, 100160, 100220, 
    100250, 100260, 100270, 100270, 100270, 100270, 100290, 100320, 100350, 
    100360, 100380, 100360, 100430, 100410, 100420, 100470, 100470, 100410, 
    100400, 100420, 100410, 100390, 100370, 100320, 100290, 100260, 100300, 
    100330, 100370, 100340, 100270, 100300, 100320, 100380, 100350, 100330, 
    100340, 100320, 100320, 100360, 100350, 100340, 100330, 100320, 100310, 
    100340, 100410, 100430, 100460, 100460, 100470, 100550, 100580, 100600, 
    100610, 100600, 100580, 100610, 100630, 100620, 100640, 100660, 100670, 
    100670, 100720, 100720, 100710, 100720, 100700, 100730, 100730, 100760, 
    100800, 100800, 100780, 100780, 100820, 100810, 100820, 100870, 100860, 
    100880, 100900, 100910, 100920, 100950, 101010, 100990, 101040, 101040, 
    101090, 101070, 101130, 101140, 101180, 101180, 101180, 101230, 101260, 
    101320, 101370, 101380, 101370, 101360, 101340, 101380, 101380, 101380, 
    101380, 101400, 101390, 101400, 101400, 101330, 101390, 101370, 101350, 
    101400, 101430, 101440, 101500, 101530, 101600, 101650, 101680, 101750, 
    101750, 101740, 101760, 101740, 101770, 101780, 101770, 101790, 101830, 
    101860, 101870, 101840, 101830, 101820, 101830, 101830, 101840, 101820, 
    101810, 101820, 101850, 101870, 101890, 101900, 101860, 101820, 101810, 
    101790, 101740, 101760, 101750, 101730, 101730, 101760, 101790, 101770, 
    101800, 101800, 101790, 101740, 101730, 101760, 101710, 101720, 101730, 
    101740, 101720, 101700, 101670, 101640, 101610, 101590, 101570, 101550, 
    101480, 101380, 101360, 101360, 101360, 101340, 101240, 101190, 101100, 
    101060, 101040, 100980, 100970, 100950, 100990, 100980, 100810, 100930, 
    100810, 100570, 100480, 100440, 100380, 100390, 100350, 100370, 100300, 
    100240, 100140, 100130, 100180, 100180, 100170, 100150, 99980, 99890, 
    99720, 99590, 99530, 99420, 99420, 99390, 99300, 99170, 99050, 98880, 
    98790, 98760, 98700, 98650, 98660, 98640, 98630, 98620, 98590, 98480, 
    98340, 98320, 98400, 98390, 98440, 98510, 98630, 98700, 98620, 98730, 
    98790, 98800, 98840, 98890, 98950, 99030, 99010, 99050, 99070, 99030, 
    99020, 99050, 99040, 99020, 99000, 99050, 99040, 99010, 99020, 99040, 
    99080, 99090, 99060, 99040, 99030, 98950, 98870, 98830, 98780, 98760, 
    98750, 98720, 98680, 98680, 98630, 98600, 98570, 98560, 98510, 98480, 
    98490, 98500, 98500, 98470, 98480, 98530, 98640, 98710, 98720, 98740, 
    98770, 98820, 98840, 98880, 98910, 98990, 99020, 99050, 99020, 99080, 
    99130, 99240, 99360, 99460, 99530, 99640, 99680, 99790, 99930, 100030, 
    100130, 100230, 100300, 100370, 100430, 100480, 100530, 100620, 100670, 
    100740, 100800, 100870, 100960, 101000, 101080, 101130, 101190, 101240, 
    101250, 101280, 101300, 101350, 101400, 101460, 101480, 101550, 101580, 
    101610, 101630, 101640, 101660, 101670, 101690, 101720, 101740, 101730, 
    101750, 101770, 101750, 101720, 101730, 101710, 101700, 101650, 101640, 
    101630, 101630, 101650, 101630, 101630, 101610, 101610, 101630, 101620, 
    101640, 101630, 101610, 101620, 101600, 101570, 101580, 101570, 101530, 
    101480, 101460, 101420, 101380, 101310, 101290, 101260, 101210, 101180, 
    101140, 101090, 101070, 101020, 100930, 100880, 100840, 100780, 100700, 
    100660, 100640, 100580, 100500, 100450, 100420, 100360, 100290, 100220, 
    100200, 100170, 100150, 100150, 100160, 100140, 100130, 100110, 100080, 
    100040, 99980, 99940, 99920, 99860, 99830, 99810, 99710, 99640, 99600, 
    99530, 99480, 99430, 99350, 99310, 99290, 99350, 99410, 99520, 99620, 
    99700, 99770, 99820, 99880, 99940, 99940, 99960, 99980, 100040, 100080, 
    100120, 100180, 100210, 100240, 100270, 100280, 100300, 100340, 100340, 
    100380, 100410, 100420, 100430, 100440, 100450, 100450, 100500, 100510, 
    100520, 100520, 100550, 100540, 100590, 100610, 100610, 100640, 100620, 
    100630, 100630, 100630, 100620, 100590, 100560, 100550, 100520, 100510, 
    100500, 100510, 100500, 100500, 100480, 100470, 100490, 100520, 100550, 
    100570, 100580, 100620, 100680, 100740, 100790, 100870, 100920, 100950, 
    100950, 101040, 101040, 101030, 101040, 101010, 101060, 101100, 101140, 
    101150, 101200, 101160, 101170, 101160, 101150, 101150, 101150, 101150, 
    101130, 101130, 101110, 101090, 101080, 101050, 101010, 100970, 100940, 
    100890, 100850, 100820, 100790, 100800, 100780, 100720, 100680, 100630, 
    100550, 100480, 100430, 100430, 100390, 100400, 100390, 100400, 100430, 
    100470, 100410, 100490, 100440, 100470, 100510, 100510, 100510, 100550, 
    100600, 100630, 100740, 100660, 100750, 100770, 100750, 100740, 100740, 
    100780, 100790, 100790, 100820, 100870, 100880, 100860, 100870, 100860, 
    100880, 100890, 100810, 100780, 100820, 100860, 100880, 100910, 100880, 
    100900, 100920, 100900, 100890, 100890, 100880, 100900, 100900, 100900, 
    100910, 100910, 100890, 100880, 100860, 100860, 100850, 100830, 100810, 
    100830, 100800, 100800, 100820, 100820, 100870, 100890, 100910, 100940, 
    100970, 100960, 100970, 100960, 100970, 101000, 101010, 101050, 101050, 
    101080, 101120, 101130, 101140, 101160, 101150, 101180, 101190, 101190, 
    101220, 101260, 101260, 101270, 101250, 101250, 101250, 101270, 101300, 
    101260, 101280, 101270, 101250, 101260, 101330, 101320, 101290, 101290, 
    101330, 101300, 101270, 101240, 101220, 101250, 101270, 101310, 101300, 
    101340, 101350, 101340, 101380, 101410, 101410, 101430, 101440, 101440, 
    101440, 101470, 101490, 101480, 101440, 101410, 101360, 101320, 101280, 
    101170, 101170, 101130, 101060, 101030, 101010, 100960, 100930, 100860, 
    100790, 100760, 100730, 100700, 100670, 100650, 100660, 100700, 100790, 
    100900, 100970, 101040, 101130, 101110, 101230, 101240, 101150, 101210, 
    101140, 101020, 101040, 100920, 100830, 100710, 100560, 100420, 100310, 
    100240, 100150, 100000, 99960, 99940, 99950, 99950, 99900, 100010, 99950, 
    100000, 100100, 100110, 100140, 100210, 100350, 100410, 100480, 100640, 
    100730, 100810, 100940, 101040, 101150, 101300, 101350, 101440, 101650, 
    101800, 101880, 101930, 102000, 102080, 102140, 102230, 102180, 102240, 
    102260, 102250, 102280, 102250, 102280, 102240, 102210, 102100, 102030, 
    101980, 101930, 101840, 101770, 101700, 101600, 101490, 101430, 101300, 
    101180, 101020, 100810, 100650, 100410, 100310, 100180, 100120, 100080, 
    100050, 100020, 99940, 99920, 99910, 99860, 99890, 99910, 99930, 99890, 
    99910, 99900, 99920, 99920, 99920, 99900, 99850, 99840, 99810, 99800, 
    99800, 99810, 99830, 99850, 99900, 99960, 100000, 100040, 100080, 100110, 
    100130, 100160, 100140, 100160, 100200, 100210, 100280, 100290, 100350, 
    100360, 100400, 100410, 100430, 100440, 100460, 100480, 100490, 100520, 
    100550, 100590, 100640, 100680, 100700, 100720, 100770, 100820, 100890, 
    100900, 100940, 100970, 101020, 101050, 101100, 101150, 101190, 101210, 
    101240, 101270, 101300, 101340, 101360, 101400, 101430, 101480, 101510, 
    101530, 101530, 101560, 101580, 101470, 101550, 101580, 101540, 101490, 
    101520, 101490, 101500, 101520, 101530, 101510, 101510, 101480, 101520, 
    101470, 101500, 101520, 101570, 101530, 101580, 101620, 101590, 101560, 
    101550, 101610, 101740, 101760, 101770, 101760, 101790, 101810, 101820, 
    101790, 101750, 101750, 101780, 101780, 101770, 101720, 101710, 101680, 
    101640, 101630, 101640, 101600, 101550, 101540, 101530, 101570, 101570, 
    101570, 101540, 101570, 101570, 101560, 101620, 101600, 101620, 101630, 
    101660, 101630, 101610, 101620, 101610, 101560, 101570, 101560, 101520, 
    101420, 101430, 101410, 101350, 101310, 101290, 101250, 101250, 101300, 
    101330, 101360, 101400, 101400, 101430, 101470, 101500, 101510, 101570, 
    101600, 101600, 101630, 101680, 101730, 101780, 101830, 101860, 101850, 
    101860, 101880, 101930, 101940, 101950, 101950, 101980, 102000, 102020, 
    102040, 102020, 102030, 102040, 102070, 102080, 102060, 102080, 102090, 
    102110, 102140, 102150, 102160, 102130, 102120, 102120, 102090, 102090, 
    102110, 102090, 102090, 102100, 102130, 102150, 102150, 102170, 102150, 
    102150, 102190, 102200, 102200, 102210, 102240, 102260, 102310, 102350, 
    102390, 102410, 102430, 102440, 102460, 102480, 102530, 102570, 102580, 
    102610, 102660, 102690, 102700, 102710, 102680, 102690, 102700, 102710, 
    102720, 102690, 102700, 102720, 102780, 102790, 102770, 102820, 102780, 
    102800, 102800, 102800, 102790, 102780, 102820, 102800, 102750, 102800, 
    102800, 102840, 102740, 102720, 102780, 102720, 102730, 102710, 102680, 
    102740, 102870, 102880, 102890, 102890, 102860, 102850, 102890, 102900, 
    102910, 102900, 102800, 102800, 102830, 102830, 102800, 102750, 102700, 
    102690, 102640, 102610, _, 102580, _, _, 102500, 102440, 102370, 102370, 
    102210, 102060, 101930, 101870, 101780, 101650, 101560, 101510, 101480, 
    101460, 101370, 101270, 101210, 101160, 101150, 101140, 101110, 101070, 
    101060, 101060, 101030, 101000, 100930, 100860, 100700, 100560, 100410, 
    100200, 100010, 99830, 99660, 99540, 99420, 99300, 99180, 99100, 98980, 
    98870, 98740, 98580, 98440, 98280, 98160, 97990, 97840, 97760, 97680, 
    97590, 97520, 97440, 97350, 97290, 97350, 97360, 97420, 97510, 97600, 
    97680, 97730, 97770, 97800, 97930, 97980, 98010, 98010, 97990, 98010, 
    98020, 98050, 98070, 98080, 98090, 98100, 98080, _, 98040, 98020, _, _, 
    97850, _, 97800, 97740, 97650, _, 97560, _, 97440, 97370, 97340, 97300, 
    97280, _, 97300, 97290, 97310, 97310, 97350, 97390, 97420, 97490, 97580, 
    97690, 97810, 97850, _, 98030, _, 98090, 98130, 98170, 98240, 98270, 
    98290, 98310, 98320, 98330, 98300, 98310, 98300, 98290, 98290, 98290, 
    98320, 98320, 98340, 98340, 98350, 98380, 98360, 98380, 98370, 98340, 
    98330, 98310, 98290, 98270, 98240, 98240, 98210, 98200, 98190, 98140, 
    98090, 98060, 98000, 97990, 97940, 97850, 97820, 97790, 97750, 97720, 
    97720, 97710, 97700, 97700, 97710, 97700, 97700, 97720, 97760, 97810, 
    97870, 97920, 97950, 97970, 98000, 98050, 98080, 98110, 98150, 98150, 
    98170, 98210, 98270, 98320, 98370, 98400, 98430, 98450, 98480, 98520, 
    98530, 98570, 98610, 98640, 98680, 98720, 98750, 98770, 98770, 98780, 
    98810, 98810, 98800, 98810, 98760, 98770, 98770, 98790, 98790, 98790, 
    98750, 98710, 98690, 98690, 98690, 98700, 98670, 98700, 98700, 98690, 
    98720, 98700, 98660, 98660, 98630, 98640, 98720, 98720, 98720, 98730, 
    98740, 98760, 98760, 98740, 98760, 98750, 98740, 98770, 98790, 98840, 
    98870, 98910, 98940, 98970, 99030, 99070, 99110, 99180, 99240, 99310, 
    99380, 99410, 99430, 99480, 99560, 99590, 99660, 99730, 99770, 99810, 
    99870, 99920, 99970, 100000, 100040, 100100, 100180, 100220, 100290, 
    100340, 100370, 100390, 100470, 100520, 100550, 100600, 100640, 100690, 
    100720, 100770, 100830, 100890, 100990, 101080, 101220, 101310, 101390, 
    101500, 101500, 101590, 101700, 101740, 101710, 101680, 101610, 101510, 
    101370, 101260, 101040, 100870, 100620, 100340, 100090, 99800, 99580, 
    99370, 99040, 98890, 98600, 98530, 98360, 98300, 98220, 98190, 98200, 
    98200, 98200, 98240, 98240, 98190, 98150, 98080, 98070, 98020, 97980, 
    98020, 98050, 98110, 98150, 98140, 98140, 98120, 98140, 98190, 98220, 
    98240, 98320, 98410, 98460, 98510, 98470, 98470, 98500, 98450, 98370, 
    98270, 98190, 98140, 98160, 98070, 98030, 97960, 97910, 97900, 97850, 
    97770, 97770, 97830, 97900, 97960, 97970, 98080, 98220, 98300, 98430, 
    98450, 98470, 98490, 98530, 98540, 98560, 98580, 98640, 98640, 98680, 
    98700, 98730, 98770, 98780, 98790, 98790, 98780, 98770, 98770, 98770, 
    98780, 98760, 98780, 98800, 98780, 98780, 98780, 98780, 98780, 98740, 
    98710, 98670, 98690, 98710, 98700, 98680, 98690, 98660, 98660, 98660, 
    98680, 98670, 98660, 98650, 98630, 98630, 98650, 98670, 98670, 98670, 
    98660, 98670, 98640, 98650, 98650, 98650, 98640, 98630, 98630, 98610, 
    98580, 98600, 98560, 98560, 98540, 98500, 98520, 98550, 98560, 98600, 
    98620, 98640, 98650, 98640, 98640, 98650, 98660, 98650, 98640, 98650, 
    98660, 98660, 98680, 98700, 98690, 98690, 98670, 98680, 98660, 98600, 
    98560, 98510, 98440, 98400, 98330, 98240, 98180, 98020, 97980, 97980, 
    97980, 98020, 98110, 98210, 98320, 98430, 98540, 98660, 98760, 98850, 
    98930, 99010, 99110, 99190, 99250, 99330, 99420, 99510, 99590, 99680, 
    99770, 99840, 99900, 99980, 100040, 100090, 100140, 100210, 100250, 
    100320, 100370, 100430, 100470, 100500, 100500, 100560, 100550, 100610, 
    100630, 100600, 100690, 100710, 100740, 100730, 100830, 100820, 100840, 
    100840, 100840, 100890, 100910, 100880, 100850, 100810, 100750, 100650, 
    100580, 100370, 100380, 100360, 100370, 100350, 100290, 100250, 100200, 
    100160, 100150, 100120, 100070, 100080, 99960, 99920, 99880, 99860, 
    99820, 99760, 99690, 99660, 99620, 99600, 99580, 99590, 99620, 99660, 
    99710, 99720, 99700, 99730, 99760, 99780, 99810, 99840, 99910, 99970, 
    100050, 100080, 100150, 100220, 100290, 100340, 100420, 100450, 100530, 
    100640, 100730, 100840, 100840, 100870, 100890, 100920, 100940, 100960, 
    101050, 101080, 101120, 101200, 101200, 101170, 101230, 101230, 101290, 
    101210, 101220, 101220, 101240, 101210, 101180, 101140, 101140, 101100, 
    101080, 101040, 100990, 100950, 100880, 100870, 100850, 100840, 100820, 
    100770, 100750, 100730, 100750, 100690, 100650, 100670, 100650, 100620, 
    100600, 100580, 100560, 100600, 100580, 100560, 100540, 100550, 100500, 
    100430, 100460, 100510, 100440, 100430, 100420, 100350, 100370, 100350, 
    100390, 100450, 100460, 100430, 100390, 100390, 100410, 100460, 100460, 
    100470, 100480, 100480, 100470, 100480, 100510, 100490, 100530, 100570, 
    100570, 100590, 100590, 100620, 100620, 100650, 100550, 100510, 100460, 
    100370, 100420, 100200, 100320, 100290, 100220, 100230, 100280, 100050, 
    100090, 100020, 100080, 100120, 100060, 100010, 99960, 99900, 99900, 
    99940, 99930, 99910, 99860, 99900, 99880, 99880, 99850, 99860, 99930, 
    99960, 99980, 100010, 100040, 100100, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 101770, 101760, 101720, 101640, 101520, 101380, 101200, 100990, 
    100730, 100380, 100120, 99820, 99590, 99400, 99140, 98960, 99020, 99000, 
    98980, 98890, 98870, 98760, 98600, 98370, 98110, 97810, 97430, 97210, 
    97100, 97170, 97420, 97600, 97780, 97920, 98090, 98230, 98440, 98520, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 101320, 101330, 101370, 101410, 101450, 101490, 101530, 
    101610, 101640, 101680, 101710, 101740, 101760, 101770, 101820, 101840, 
    101860, 101900, 101930, 101970, 102000, 102000, 101990, 101960, 101950, 
    102000, 101930, 101940, 101960, 101950, 101970, 101950, 101920, 101920, 
    101910, 101930, 101890, 101850, 101830, 101840, 101840, 101890, 101890, 
    101950, 101950, 101910, 101950, 101950, 101970, 101940, 101940, 101940, 
    101960, 101980, 102030, 102030, 101980, 101960, 101940, 101970, 101960, 
    101960, 101970, 101950, 101890, 101900, 101930, 101960, 101980, 101970, 
    101970, 101970, 101940, 101890, 101870, 101880, 101880, 101880, 101900, 
    101890, 101890, 101890, 101870, 101870, 101860, 101890, 101900, 101870, 
    101850, 101820, 101790, 101790, 101810, 101800, 101790, 101740, 101670, 
    101660, 101630, 101560, 101560, 101530, 101480, 101430, 101430, 101390, 
    101330, 101290, _, 101250, _, _, 101200, 101220, 101250, 101270, 101270, 
    101290, _, 101290, 101280, _, 101300, 101320, _, 101290, 101300, _, _, _, 
    _, 101330, 101290, 101300, 101310, _, 101340, 101330, 101370, 101350, 
    101410, 101390, 101390, 101420, 101400, 101370, 101440, 101450, 101420, 
    101440, 101450, 101470, 101480, 101470, 101470, 101420, 101380, 101420, 
    101380, 101380, 101350, 101310, 101310, 101340, 101360, 101420, 101400, 
    101370, 101330, 101390, 101440, 101440, 101430, 101430, 101450, 101440, 
    101440, 101420, 101430, 101410, 101420, 101410, 101410, 101430, 101470, 
    101450, 101470, 101440, 101360, 101330, 101320, 101290, 101220, 101160, 
    101090, 101030, 100990, 100950, 100880, 100750, 100710, 100670, 100540, 
    100420, 100360, 100300, 100200, 100140, 100110, 100060, 99980, 99900, 
    99780, 99750, 99730, 99690, 99680, 99630, 99630, 99660, 99690, 99720, 
    99770, 99790, 99820, 99840, 99850, 99800, 99840, 99850, 99840, 99810, 
    99810, 99780, 99740, _, _, _, 99500, 99440, 99370, 99320, 99270, 99200, 
    99150, 99120, 99120, 99100, 99070, 99040, 99030, 99010, 98980, 98950, 
    98950, 98990, 99000, 98980, 98970, 98970, 98990, 98990, 98960, 98950, 
    98950, 98960, 99010, 99050, 99110, 99170, 99250, 99380, 99570, 99620, 
    99660, 99740, 99780, 99890, 99970, 100040, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 100500, 100350, 100360, 
    100390, 100190, 100160, 100000, 99940, _, 99920, 99780, 99820, 99760, 
    99610, _, _, 99580, 99580, 99560, 99610, 99630, 99680, 99690, 99700, _, 
    99800, 99900, 99920, 99960, _, 100030, 100100, 100120, 100170, 100210, 
    100270, 100270, 100250, 100230, 100280, 100300, 100300, 100310, 100330, 
    100290, 100190, 100180, 100220, 100230, 100190, 100170, 100070, 100080, 
    100060, 100010, 99930, 99850, 99780, 99760, 99700, 99660, 99640, 99660, 
    99620, 99650, 99640, 99650, 99660, 99680, 99750, 99800, 99850, 99920, 
    99980, 100030, 100110, 100180, 100270, 100380, 100480, 100540, 100660, 
    100770, 100860, 100980, 101100, 101120, 101200, 101280, 101410, 101480, 
    101570, 101620, 101700, 101760, 101820, _, 101810, 101830, 101870, 
    101920, 101940, 101980, 101980, 101970, 102040, 102130, 102140, 102210, 
    102240, 102260, 102300, 102340, 102360, 102390, 102430, 102430, 102450, 
    102500, 102560, 102580, 102600, 102640, 102670, 102710, 102710, 102740, 
    102770, 102810, 102830, 102870, 102880, 102880, 102900, 102920, 102910, 
    102930, 102920, 102920, 102950, 102920, 102920, 102900, 102880, 102870, 
    102840, 102830, 102810, 102800, 102810, 102760, 102660, 102600, 102610, 
    102540, 102400, 102310, 102120, 102130, 102030, 101860, 101760, 101680, 
    101660, 101600, 101490, 101430, 101300, 101180, 101030, 100910, 100830, 
    100690, 100600, 100520, 100430, 100340, 100270, 100200, 100120, 100020, 
    99980, 99890, 99800, 99770, _, 99730, 99690, 99630, 99500, 99460, 99450, 
    99370, 99190, 99140, 99030, 98980, 98950, 98860, 98780, 98690, 98670, 
    98620, 98610, 98630, 98630, 98650, 98650, 98650, 98650, 98700, 98740, 
    98770, 98820, 98830, 98910, 98970, 99030, 99080, 99140, 99210, 99250, 
    99330, 99380, 99410, 99440, 99490, 99530, 99570, 99610, 99660, 99680, 
    99690, 99700, 99730, 99740, 99770, 99760, 99730, 99720, 99730, 99740, 
    99720, 99720, 99710, 99640, 99570, 99510, 99480, 99440, 99470, 99450, 
    99430, 99380, 99340, 99340, 99380, 99350, 99340, 99350, 99360, 99350, 
    99330, 99360, 99400, 99450, 99470, 99480, 99480, 99490, 99500, 99500, 
    99510, 99520, 99530, 99550, 99540, 99580, 99610, 99610, 99620, 99640, 
    99640, 99650, 99690, 99760, 99780, 99830, 99880, 99910, 99930, 99960, 
    100000, 100020, 100010, 100030, 100050, 100060, 100080, 100110, 100130, 
    100150, 100160, 100180, 100180, 100190, 100210, 100230, 100270, 100310, 
    100360, 100360, 100390, 100430, 100440, 100430, 100430, 100450, 100450, 
    100460, 100490, 100500, 100510, 100500, 100480, 100510, 100510, 100490, 
    100450, 100470, 100490, 100480, 100490, 100500, 100480, 100490, 100480, 
    100440, 100420, 100360, 100320, 100300, 100270, 100250, 100220, 100160, 
    100130, 100100, 100070, 100040, 100000, 99910, 99890, 99870, 99880, 
    99880, 99930, 99960, 99970, 100000, 100050, 100090, 100110, 100150, 
    100200, 100260, 100300, 100350, 100410, 100460, 100490, 100530, 100570, 
    100610, 100650, 100660, 100670, 100680, 100700, 100800, 100820, 100830, 
    100850, 100830, 100710, 100690, 100650, 100650, 100630, 100570, 100520, 
    100470, 100410, 100330, 100260, 100180, 100130, 100020, 99930, 99840, 
    99710, 99640, 99630, 99620, 99630, 99680, 99820, 99980, 100120, 100200, 
    100320, 100410, 100510, 100540, 100620, 100700, 100780, 100800, 100900, 
    100930, 100890, 100860, 100810, 100690, 100610, 100510, 100410, 100350, 
    100210, 100090, 99960, 99870, 99740, 99650, 99540, 99450, 99360, 99300, 
    99260, 99210, 99180, 99160, 99180, 99180, 99210, 99230, 99260, 99330, 
    99410, 99500, 99570, 99720, 99810, 99890, 99980, 99980, 100060, 100150, 
    100220, 100280, 100360, 100430, 100460, 100520, 100540, 100570, 100610, 
    100640, 100620, 100610, 100590, 100610, 100610, 100610, 100640, 100640, 
    100650, 100680, 100710, 100730, 100760, 100800, 100830, 100850, 100880, 
    100930, 101020, 101070, 101110, 101120, 101160, 101200, 101220, 101240, 
    101240, 101260, 101280, 101300, 101340, 101330, 101350, 101300, 101280, 
    101260, 101220, 101160, 101150, 101110, 101070, 100880, 100870, 100860, 
    100850, 100810, 100770, 100750, 100730, 100710, 100660, 100650, 100610, 
    100590, 100530, 100540, 100540, 100540, 100500, 100390, 100380, 100450, 
    100410, 100380, 100320, 100170, 100160, 99990, 100080, 100200, 100300, 
    100550, 100740, 100820, 101130, 101120, 101570, 101660, 101750, 101890, 
    101910, 101970, 101930, 102110, 102130, 102150, 102140, 102140, 102180, 
    102200, 102130, 102200, 102250, 102240, 102280, 102260, 102220, 102270, 
    102300, 102240, 102050, 101850, 102070, 101880, 101790, 101680, 101580, 
    101500, 101390, 101340, 101310, 101280, 101200, 101180, 101190, 101180, 
    101170, 101120, 101190, 101210, 101340, 101320, 101340, 101350, 101360, 
    101370, 101470, 101470, 101470, 101480, 101410, 101440, 101530, 101460, 
    101500, 101490, 101500, 101510, 101450, 101490, 101480, 101480, 101460, 
    101500, 101480, 101500, 101480, 101480, 101490, 101460, 101340, 101410, 
    101390, 101390, 101400, 101370, 101390, 101390, 101420, 101480, 101490, 
    101530, 101530, 101550, 101580, 101600, 101630, 101640, 101690, 101710, 
    101740, 101760, 101760, 101790, 101820, 101810, 101830, 101800, 101800, 
    101800, 101810, 101820, 101830, 101840, 101840, 101840, 101830, 101830, 
    101830, 101840, 101830, 101840, 101820, 101810, 101790, 101800, 101840, 
    101890, 101910, 101900, 101900, 101890, 101910, 101940, 101950, 101970, 
    102000, 102020, 102040, 102050, 102030, 102030, 102030, 102030, 102010, 
    101980, 101990, 101990, 101970, 101970, 101960, 101950, 101960, 101950, 
    101940, 101880, 101870, 101870, 101860, 101860, 101830, 101850, 101850, 
    101830, 101820, 101810, 101780, 101760, 101730, 101710, 101710, 101340, 
    101320, 101300, 101290, 101270, 101270, 101270, 101260, 101250, 101260, 
    101270, 101260, 101260, 101260, 101290, 101290, 101300, 101310, 101330, 
    101400, 101450, 101480, 101510, 101550, 101590, 101620, 101670, 101710, 
    101760, 101780, 101790, 101810, 101840, 101880, 101900, 101940, 101960, 
    101970, 102000, 101990, 101990, 102010, 102020, 102000, 101990, 102000, 
    101990, 101950, 101960, 101990, 102000, 102000, 102010, 102000, 101980, 
    101980, 101990, 102010, 101990, 101990, 101970, 101960, 101920, 101900, 
    101890, 101890, 101890, 101860, 101820, 101740, 101620, 101570, 101540, 
    101460, 101440, 101450, 101440, 101390, 101350, 101310, 101290, 101300, 
    101270, 101270, 101270, 101290, 101330, 101370, 101410, 101450, 101500, 
    101530, 101570, 101580, 101590, 101600, 101670, 101690, 101760, 101760, 
    101770, 101790, 101830, 101860, 101870, 101880, 101880, 101890, 101900, 
    101910, 101920, 101990, 102060, 102100, 102090, 102100, 102090, 102140, 
    102180, 102180, 102220, 102240, 102230, 102240, 102250, 102250, 102250, 
    102230, 102220, 102220, 102210, 102170, 102130, 102100, 102080, 102040, 
    102000, 101950, 101930, 101870, 101820, 101760, 101740, 101720, 101680, 
    101640, 101630, 101610, 101580, 101420, 101340, 101370, 101380, 101360, 
    101320, 101270, 101220, 101170, 101110, 101080, 101030, 100980, 100910, 
    100860, 100820, 100780, 100760, 100730, 100720, 100700, 100670, 100660, 
    100670, 100650, 100640, 100630, 100600, 100580, 100580, 100610, 100630, 
    100670, 100720, 100740, 100760, 100760, 100740, 100760, 100780, 100830, 
    100860, 100900, 100910, 100940, 100970, 100990, 101020, 101040, 101050, 
    101040, 101060, 101080, 101090, 101110, 101110, 101130, 101150, 101170, 
    101170, 101170, 101150, 101150, 101180, 101200, 101210, 101210, 101200, 
    101210, 101230, 101250, 101250, 101240, 101250, 101280, 101310, 101320, 
    101360, 101400, 101420, 101430, 101450, 101490, 101520, 101530, 101560, 
    101570, 101610, 101650, 101670, 101710, 101740, 101760, 101780, 101790, 
    101800, 101820, 101830, 101830, 101820, 101860, 101860, 101850, 101820, 
    101790, 101790, 101800, 101780, 101770, 101740, 101710, 101720, 101710, 
    101690, 101680, 101670, 101670, 101660, 101630, 101590, 101590, 101570, 
    101550, 101540, 101530, 101480, 101460, 101470, 101450, 101430, 101410, 
    101390, 101380, 101340, 101320, 101290, 101270, 101230, 101180, 101140, 
    101130, 101080, 101010, 100970, 100920, 100860, 100780, 100750, 100710, 
    100670, 100670, 100670, 100670, 100730, 100730, 100730, 100740, 100780, 
    100880, 100950, 101050, 101130, 101180, 101240, 101310, 101330, 101370, 
    101400, 101460, 101480, 101490, 101490, 101530, 101560, 101610, 101610, 
    101660, 101670, 101690, 101700, 101710, 101730, 101760, 101800, 101820, 
    101830, 101850, 101850, 101860, 101840, 101840, 101810, 101790, 101760, 
    101710, 101650, 101590, 101600, 101560, 101560, 101570, 101550, 101520, 
    101520, 101510, 101510, 101510, 101510, 101520, 101520, 101520, 101530, 
    101520, 101510, 101490, 101470, 101420, 101380, 101380, 101390, 101380, 
    101360, 101360, 101360, 101340, 101350, 101300, 101290, 101260, 101260, 
    101260, 101280, 101270, 101250, 101240, 101190, 101170, 101100, 101090, 
    101060, 101000, 100980, 100960, 100950, 100900, 100900, 100840, 100830, 
    100780, 100740, 100700, 100650, 100610, 100550, 100530, 100460, 100460, 
    100410, 100360, 100300, 100260, 100190, 100100, 100020, 99920, 99850, 
    99740, 99610, 99540, 99420, 99350, 99280, 99250, 99230, 99160, 99190, 
    99190, 99160, 99170, 99170, 99170, 99150, 99160, 99160, 99150, 99140, 
    99110, 99150, 99140, 99190, 99250, 99290, 99330, 99360, 99350, 99420, 
    99450, 99450, 99510, 99610, 99620, 99660, 99700, 99770, 99800, 99850, 
    99920, 99970, 100020, 100070, 100140, 100170, 100220, 100270, 100340, 
    100390, 100420, 100460, 100510, 100570, 100630, 100640, 100890, 100910, 
    100970, 100990, 101000, 101010, 101030, 101050, 101060, 101080, 101060, 
    101070, 101090, 101100, 101090, 101080, 101100, 101110, 101120, 101140, 
    101190, 101220, 101240, 101270, 101290, 101300, 101340, 101370, 101380, 
    101410, 101430, 101450, 101470, 101480, 101550, 101590, 101620, 101680, 
    101720, 101750, 101780, 101810, 101820, 101860, 101880, 101900, 101920, 
    101920, 101950, 101960, 101990, 102010, 102020, 102040, 102060, 102060, 
    102080, 102080, 102080, 102080, 102080, 102090, 102120, 102120, 102120, 
    102130, 102140, 102130, 102120, 102110, 102100, 102090, 102080, 102060, 
    102050, 102040, 102020, 102010, 102000, 101980, 101960, 101950, 101930, 
    101910, 101910, 101930, 101920, 101920, 101910, 101900, 101870, 101860, 
    101850, 101850, 101850, 101820, 101850, 101820, 101810, 101810, 101810, 
    101800, 101790, 101800, 101780, 101740, _, 101710, 101690, 101670, 
    101690, _, 101650, _, _, 101610, 101570, 101530, 101490, 101500, 101460, 
    101440, 101450, 101420, 101410, _, 101380, 101340, 101310, 101290, _, 
    101240, 101220, 101190, 101170, _, 101100, 101110, 101040, _, _, 100910, 
    100870, 100860, 100860, 100800, 100840, 100860, 100810, 100800, 100790, 
    100800, 100790, 100820, 100800, 100810, 100790, 100830, 100780, 100860, 
    100910, 101010, 101040, 101100, 101140, 101160, 101190, 101210, 101220, 
    101250, 101310, 101390, 101390, 101430, 101440, 101420, 101420, 101440, 
    101460, 101460, 101460, 101460, 101450, 101470, 101470, 101460, 101480, 
    101490, 101490, 101460, 101460, 101440, 101440, 101430, 101400, 101410, 
    101420, 101390, 101370, 101340, 101290, 101260, 101200, 101190, 101170, 
    101160, 101100, 101100, 101050, 101060, 101010, 100980, 100910, 100850, 
    100790, 100750, 100630, 100600, 100550, 100470, 100390, 100310, 100190, 
    100110, 99990, 99920, 99860, 99810, 99760, 99690, 99660, 99640, 99570, 
    99540, 99520, 99470, 99430, 99390, 99390, 99330, 99270, 99260, 99250, 
    99230, 99220, 99180, 99150, 99130, 99070, 99090, 99020, 99020, 99030, 
    99050, 99040, 99070, 99060, 99030, 99080, 99080, 99100, 99110, 99050, 
    99050, 99060, 99010, 99000, 99010, 99020, 99020, 98980, 99050, 99000, 
    98990, 99020, 99000, 99030, 99060, 99110, 99150, 99190, 99240, 99280, 
    99290, 99320, 99380, 99400, 99420, 99470, 99520, 99540, 99570, 99600, 
    99670, 99740, 99800, 99850, 99900, 99920, 99950, 100010, 100060, 100100, 
    100140, 100180, 100210, 100250, 100270, 100300, 100330, 100360, 100370, 
    100400, 100410, 100410, 100430, 100420, 100460, 100470, 100460, 100460, 
    100440, 100430, 100470, 100480, 100490, 100520, 100520, 100530, 100550, 
    100560, 100560, 100560, 100580, 100550, 100550, 100540, 100560, 100550, 
    100550, 100530, 100520, 100520, 100510, 100500, 100490, 100480, 100460, 
    100470, 100460, 100450, 100440, 100410, 100390, 100400, 100390, 100370, 
    100360, 100330, 100310, 100300, 100310, 100300, 100310, 100310, 100310, 
    100320, 100310, 100330, 100330, 100340, 100360, 100360, 100370, 100410, 
    100430, 100440, 100440, 100450, 100430, 100400, 100390, 100370, 100360, 
    100360, 100370, 100350, 100330, 100280, 100260, 100260, 100240, 100230, 
    100250, 100210, 100250, 100310, 100330, 100380, 100400, 100390, 100390, 
    100330, 100370, 100390, 100390, 100340, 100320, 100300, 100290, 100290, 
    100230, 100240, 100160, 100130, 100140, 100090, 99980, 99920, 99890, 
    99850, 99810, 99690, 99600, 99470, 99360, 99260, 99130, 99040, 98950, 
    98990, 98970, 98990, 99080, 99080, 99070, 99180, 99200, 99180, 99130, 
    99110, 99090, 99170, 99160, 99180, 99170, 99200, 99180, 99230, 99250, 
    99250, 99320, 99300, 99420, 99530, 99600, 99650, 99650, 99710, 99720, 
    99820, 99850, 99900, 99920, 99910, 99880, 99850, 99830, 99860, 99840, 
    99830, 99870, 99880, 99890, 99910, 99950, 99970, 100050, 100070, 100070, 
    100120, 100110, 100160, 100120, 100190, 100220, 100240, 100240, 100240, 
    100240, 100310, 100320, 100340, 100410, 100480, 100550, 100610, 100630, 
    100680, 100730, 100750, 100860, 100870, 100810, 100880, 100930, 100940, 
    101040, 101100, 101140, 101100, 101200, 101220, 101220, 101210, 101200, 
    101190, 101180, 101170, 101170, 101150, 101130, 101090, 101040, 101000, 
    101020, 101020, 101010, 100980, 100970, 100900, 100860, 100840, 100780, 
    100770, 100770, 100760, 100750, 100730, 100740, 100710, 100730, 100710, 
    100700, 100680, 100690, 100670, 100650, 100630, 100610, 100550, 100510, 
    100540, 100530, 100500, 100470, 100430, 100370, 100330, 100360, 100350, 
    100330, 100320, 100320, 100310, 100300, 100280, 100290, 100310, 100310, 
    100330, 100320, 100330, 100310, 100300, 100290, 100250, 100240, 100250, 
    100270, 100260, 100250, 100250, 100240, 100250, 100260, 100250, 100260, 
    100280, 100310, 100330, 100350, 100390, 100410, 100440, 100460, 100490, 
    100510, 100530, 100550, 100560, 100590, 100600, 100620, 100630, 100670, 
    100700, 100710, 100730, 100770, 100800, 100850, 100860, 100900, 100930, 
    100940, 100980, 101010, 101010, 101050, 101060, 101080, 101100, 101110, 
    101130, 101150, 101180, 101200, 101210, 101230, 101240, 101270, 101270, 
    101290, 101290, 101300, 101310, 101310, 101330, 101360, 101380, 101370, 
    101370, 101390, 101400, 101390, 101420, 101430, 101430, 101460, 101470, 
    101480, 101500, 101530, 101530, 101540, 101530, 101550, 101570, 101570, 
    101580, 101620, 101650, 101690, 101710, 101750, 101760, 101800, 101820, 
    101840, 101870, 101890, 101910, 101950, 101970, 102000, 102010, 102020, 
    102040, 102040, 102040, 102070, 102070, 102080, 102100, 102110, 102110, 
    102120, 102130, 102150, 102140, 102170, 102140, 102140, 102150, 102140, 
    102130, 102130, 102140, 102150, 102140, 102160, 102160, 102160, 102170, 
    102150, 102140, 102140, 102150, 102140, 102130, 102150, 102160, 102150, 
    102150, 102140, 102130, 102100, 102090, 102080, 102100, 102070, 102090, 
    102080, 102080, 102070, 102060, 102060, 102030, 102030, 102000, 101970, 
    101970, 101980, 101990, 101970, 101950, 101950, 101920, 101910, 101880, 
    101880, 101860, 101860, 101850, 101840, 101830, 101820, 101800, 101790, 
    101770, 101750, 101770, 101750, 101710, 101690, 101680, 101660, 101660, 
    101650, 101640, 101620, 101610, 101600, 101580, 101580, 101550, 101470, 
    101450, 101470, 101470, 101450, 101480, 101490, 101500, 101480, 101480, 
    101450, 101480, 101480, 101480, 101500, 101490, 101490, 101460, 101430, 
    101420, 101420, 101390, 101380, 101370, 101350, 101320, 101310, 101280, 
    101260, 101240, 101230, 101220, 101230, 101230, 101200, 101180, 101180, 
    101160, 101170, 101180, 101210, 101230, 101240, 101250, 101270, 101270, 
    101280, 101310, 101310, 101330, 101370, 101390, 101410, 101430, 101440, 
    101470, 101490, 101490, 101510, 101530, 101540, 101560, 101560, 101600, 
    101630, 101650, 101670, 101660, 101660, 101690, 101680, 101680, 101660, 
    101640, 101640, 101640, 101650, 101620, 101620, 101600, 101570, 101530, 
    101540, 101510, 101500, 101480, 101470, 101450, 101430, 101380, 101340, 
    101340, 101320, 101320, 101300, 101290, 101280, 101260, 101230, 101270, 
    101280, 101280, 101290, 101290, 101270, 101290, 101320, 101320, 101360, 
    101370, 101430, 101500, 101540, 101570, 101580, 101600, 101640, 101660, 
    101660, 101640, 101630, 101610, 101590, 101570, 101600, 101630, 101630, 
    101620, 101600, 101600, 101610, 101590, 101570, 101580, 101600, 101590, 
    101590, 101600, 101610, 101580, 101570, 101570, 101560, 101530, 101520, 
    101520, 101490, 101450, 101470, 101480, 101440, 101410, 101380, 101360, 
    101340, 101350, 101340, 101330, 101320, 101320, 101320, 101310, 101310, 
    101270, 101250, 101230, 101250, 101230, 101220, 101200, 101220, 101230, 
    101220, 101220, 101240, 101240, 101250, 101260, 101270, 101300, 101320, 
    101350, 101370, 101400, 101450, 101490, 101520, 101550, 101570, 101600, 
    101630, 101640, 101650, 101680, 101680, 101720, 101720, 101740, 101760, 
    101760, 101800, 101810, 101830, 101880, 101900, 101930, 101970, 102010, 
    102070, 102090, 102120, 102180, 102210, 102220, 102240, 102260, 102300, 
    102290, 102300, 102300, 102320, 102320, 102350, 102360, 102370, 102350, 
    102380, 102370, 102380, 102400, 102420, 102440, 102470, 102490, 102510, 
    102540, 102540, 102540, 102570, 102570, 102580, 102570, 102540, 102550, 
    102540, 102530, 102520, 102510, 102500, 102480, 102470, 102450, 102440, 
    102430, 102440, 102460, 102440, 102420, 102400, 102380, 102360, 102330, 
    102310, 102300, 102210, 102240, 102300, 102300, 102250, 102150, 102160, 
    102170, 102150, 102120, 102100, 102050, 101990, 101970, 101900, 101960, 
    101930, 101910, 101910, 101880, 101930, 101930, 101900, 101880, 101940, 
    _, 101960, 101990, 102010, 102040, 102050, 102070, 102080, 102100, 
    102130, 102080, 102150, 102170, 102140, 102220, 102220, _, _, _, 102240, 
    _, 102290, 102250, 102230, 102260, 102230, 102240, _, _, 102230, _, 
    102190, 102170, 102150, 102120, 102080, _, 102110, _, 102080, _, _, 
    102150, 102200, 102210, 102170, _, 102180, _, 102210, 102230, 102220, _, 
    102250, 102220, 102240, _, 102240, 102250, 102190, _, 102260, 102250, _, 
    102260, 102280, 102240, 102210, 102230, 102240, 102180, 102200, 102170, 
    102170, _, _, _, _, 102130, 102130, _, 102130, 102090, 102110, 102090, 
    102120, 102100, 102140, 102180, 102180, 102170, 102190, 102210, 102180, 
    _, _, 102160, _, 102220, 102190, 102220, 102210, 102260, 102260, 102260, 
    102250, 102260, 102250, 102250, 102270, 102270, 102290, 102250, 102250, 
    102240, 102250, 102210, 102220, 102230, 102220, 102190, 102120, 102090, 
    102090, 102090, 102050, 102020, 102010, 102020, 101970, 101940, 101910, 
    101890, 101900, 101880, 101850, 101820, 101830, 101790, _, 101710, 
    101700, 101690, 101650, 101620, _, 101530, 101510, _, 101440, 101410, 
    101370, 101360, 101320, 101250, _, 101180, 101160, 101160, 101130, 
    101110, 101120, 101110, 101060, 101030, 101000, 100980, 100970, 100930, 
    100910, 100890, 100910, 100930, 100930, 100960, 100940, 100920, 100920, 
    100940, 100890, 100830, 100780, 100740, 100670, 100630, 100560, 100580, 
    100540, 100540, 100530, 100540, 100540, 100550, 100590, 100620, 100630, 
    100650, 100670, 100650, 100610, 100580, 100580, 100510, 100520, 100550, 
    100610, 100710, 100760, 100810, 100810, 100850, 100860, 100900, 100930, 
    100940, 100970, 100970, 101020, 101050, 101070, 101100, 101210, 101110, 
    _, 101190, 101220, 101220, 101250, 101290, 101270, 101300, 101350, 
    101360, 101320, 101360, 101480, 101480, 101500, 101500, 101540, 101510, 
    101520, 101520, 101490, 101440, 101400, 101370, 101400, 101400, 101380, 
    101390, 101370, 101370, 101380, 101420, 101410, 101440, 101450, 101450, 
    101480, 101510, 101510, 101490, 101500, 101500, 101510, 101530, 101540, 
    101580, 101580, 101580, 101560, 101590, 101610, 101630, 101630, 101630, 
    101630, 101630, 101630, 101650, 101660, 101660, 101660, 101670, 101680, 
    101650, 101640, 101610, 101580, 101570, 101640, 101660, 101680, 101700, 
    101690, 101680, 101660, 101650, 101650, 101630, 101630, 101650, 101640, 
    101630, 101690, 101690, 101700, 101710, 101680, 101650, 101630, 101600, 
    101570, 101540, 101560, 101590, 101570, 101560, 101550, 101530, 101520, 
    101500, 101470, 101440, 101440, 101440, 101400, 101400, 101440, 101410, 
    101430, 101420, 101400, 101380, 101380, 101350, 101330, 101300, 101280, 
    101290, 101260, 101230, 101200, 101150, 101230, 101200, 101150, 101100, 
    101040, 100970, 100940, 100900, 100840, 100780, 100700, 100680, 100590, 
    100530, 100510, 100460, 100410, 100370, 100350, 100290, 100320, 100270, 
    100260, 100230, 100190, 100160, 100170, 100180, 100210, 100220, 100250, 
    100280, 100300, 100310, 100300, _, 100290, 100230, _, _, 100150, _, _, 
    100080, 100070, _, 99990, 99950, 99950, _, _, 99880, 99930, 99940, 99990, 
    100040, 100060, 100110, 100160, _, 100250, 100290, 100330, 100380, 
    100450, _, 100560, 100580, _, 100650, 100700, 100740, 100770, 100820, 
    100820, 100870, 100890, 100900, 100920, 100960, 100960, 100990, 100990, 
    101020, 101010, 101040, _, 101080, 101120, 101140, 101180, _, 101280, 
    101330, 101380, 101430, 101490, 101540, _, 101640, 101670, _, 101750, _, 
    _, 101850, 101890, _, 101930, 101960, 102010, 102030, 102050, 102080, 
    102120, 102170, 102200, 102220, 102230, _, 102220, 102230, _, 102290, 
    102290, 102340, 102300, 102290, 102370, 102400, 102400, _, _, 102400, _, 
    102370, 102380, 102360, 102370, 102360, _, 102360, 102350, 102320, _, _, 
    102290, _, 102240, 102220, 102200, 102200, 102170, 102150, 102120, 
    102070, 101990, 101880, 101870, 101840, 101840, 101810, 101740, 101750, 
    101800, 101780, 101740, 101730, 101710, 101750, 101750, 101780, 101750, 
    _, 101770, 101810, 101830, 101850, 101840, 101900, 101930, 101870, 
    101890, 101930, 101970, 102030, 102040, 102060, 102070, 102090, 102110, 
    102190, 102180, 102210, 102240, 102260, 102260, 102240, 102350, 102330, 
    102300, _, 102370, _, _, 102360, _, 102320, 102340, _, 102280, _, 102220, 
    102270, _, 102290, _, 102280, 102310, 102300, _, _, _, _, _, _, 102270, 
    102240, 102220, _, 102270, 102230, 102250, _, 102220, 102220, 102310, _, 
    _, 102280, _, 102280, 102300, 102280, 102280, 102290, 102310, 102310, 
    102330, 102310, 102340, 102350, 102340, _, 102330, _, 102350, 102350, 
    102360, _, 102340, 102320, _, _, _, 102280, _, _, _, _, _, 102280, 
    102280, 102280, 102280, 102250, 102240, 102220, 102200, _, 102190, 
    102190, 102200, 102190, 102160, _, 102160, 102130, 102130, _, 102140, 
    102140, 102160, 102170, 102190, _, 102210, 102200, _, _, _, 102210, _, _, 
    102120, 102140, 102180, 102190, 102170, 102130, _, 102140, _, _, 102140, 
    102130, 102140, _, 102200, 102220, 102220, _, _, 102250, _, 102250, 
    102240, 102230, _, 102220, 102230, 102220, 102220, 102190, 102190, 
    102180, _, 102130, 102100, _, 102050, 102030, 102010, 101970, 101940, 
    101890, 101840, 101800, 101740, 101690, 101650, 101600, 101560, 101530, 
    101520, 101480, 101470, 101410, 101390, 101350, 101290, 101260, 101210, 
    101180, 101170, 101160, 101140, 101130, 101110, 101070, 101060, 101040, 
    101010, 101000, 100990, 100960, 100950, 100920, 100920, 100930, 100920, 
    100910, 100890, 100880, 100870, 100850, 100860, 100860, 100870, 100900, 
    _, 100940, 100950, 100970, 100990, 101000, 101000, 101010, 101010, 
    101030, 101030, 101060, 101070, 101100, 101120, 101140, 101140, _, 
    101160, 101160, 101170, 101200, 101240, 101260, 101280, 101300, 101310, 
    101300, 101310, 101320, 101300, 101290, 101290, 101240, 101220, 101230, 
    101250, 101240, 101250, 101230, 101240, 101230, 101240, 101240, 101240, 
    101230, 101250, 101260, 101270, 101290, 101290, 101310, 101310, 101300, 
    101300, 101330, 101310, 101320, 101340, 101350, 101350, 101380, 101380, 
    101380, 101380, 101390, 101390, 101390, 101380, 101390, 101420, 101440, 
    101460, 101470, 101480, 101500, 101510, 101520, 101530, 101530, 101560, 
    101570, 101580, 101610, 101610, 101630, 101650, 101660, 101650, 101660, 
    101670, 101690, 101710, 101690, 101710, 101720, 101720, 101720, 101730, 
    101750, 101730, 101730, 101720, 101710, 101690, 101670, 101670, 101650, 
    101640, 101620, 101600, 101570, 101530, 101490, 101460, 101430, 101400, 
    101370, 101350, 101350, 101340, 101330, 101290, 101290, 101280, 101260, 
    101230, 101210, 101220, 101200, 101180, 101160, 101140, 101130, 101110, 
    101110, 101100, 101100, 101090, 101090, 101100, 101100, 101110, 101130, 
    101140, 101170, 101200, 101220, 101240, 101260, 101280, 101310, 101330, 
    101350, 101370, 101400, 101450, 101500, 101550, 101580, 101620, 101650, 
    101670, 101690, 101720, 101780, 101870, 101910, 101950, 102030, 102100, 
    102150, 102190, 102240, 102260, 102280, 102300, 102350, 102400, 102460, 
    102490, 102520, 102560, 102580, 102590, 102600, 102610, 102600, 102610, 
    102650, 102670, 102680, 102670, 102700, 102730, 102720, 102700, 102700, 
    102710, 102690, 102660, 102630, 102610, 102600, 102580, 102570, 102540, 
    102510, 102490, 102480, 102440, 102430, 102400, 102340, 102350, 102360, 
    102370, 102380, 102400, 102390, 102370, 102390, 102360, 102320, 102340, 
    102310, 102280, 102270, 102260, 102200, 102170, 102150, 102120, 102080, 
    102020, 101930, 101900, 101810, 101750, 101730, 101670, 101610, 101560, 
    101470, 101420, 101390, 101280, 101210, 101110, 101050, 101010, 100950, 
    100930, 100930, 100910, 100910, 100870, 100840, 100820, 100790, 100820, 
    100810, 100820, 100850, 100880, 100890, 100960, 101030, 101110, 101110, 
    101120, 101090, 101070, 101040, 101010, 101020, 101020, 101010, 101040, 
    101060, 101050, 101020, 101000, 100970, 100960, 100950, 100950, 100960, 
    100930, 100900, 100900, 100880, 100860, 100830, 100800, 100800, 100790, 
    100780, 100800, 100840, 100870, 100900, 100900, 100930, 100940, 100940, 
    100950, 100950, 100960, 100980, 100950, 100970, 100990, 100990, 100990, 
    100990, 100980, 100990, 101010, 101020, 101040, 101080, 101110, 101160, 
    101200, 101290, 101360, 101410, 101440, 101480, 101500, 101520, 101550, 
    101530, 101600, 101660, 101720, 101770, 101830, 101840, 101860, 101930, 
    102000, 102080, 102100, 102120, 102170, 102220, 102260, 102300, 102330, 
    102370, 102420, 102430, 102430, 102460, 102490, 102510, 102550, 102590, 
    102630, 102640, 102650, 102700, 102710, 102720, 102740, 102750, 102770, 
    102750, 102750, 102740, 102720, 102690, 102690, 102640, 102590, 102510, 
    102440, 102400, 102320, 102270, 102240, 102210, 102180, 102120, 102060, 
    102010, 101970, 101910, 101860, 101820, 101790, 101760, 101730, 101710, 
    101690, 101670, 101650, 101670, 101660, 101670, 101680, 101680, 101680, 
    101670, 101710, 101740, 101750, 101780, 101810, 101840, 101850, 101870, 
    101890, 101910, 101910, 101920, 101930, 101930, 101930, 101930, 101900, 
    101880, 101880, 101850, 101830, 101810, 101790, 101750, 101750, 101740, 
    101740, 101710, 101680, 101650, 101620, 101580, 101540, 101510, 101490, 
    101460, 101450, 101450, 101480, 101460, 101430, 101380, 101380, 101360, 
    101330, 101300, 101350, 101330, 101300, 101270, 101300, 101300, 101280, 
    101280, 101240, 101320, 101300, 101280, 101320, 101310, 101330, 101360, 
    101350, 101360, 101390, 101410, 101430, 101440, 101450, 101450, 101460, 
    101460, 101490, 101510, 101530, 101550, 101570, 101600, 101630, 101630, 
    101630, 101640, 101650, 101640, 101640, 101640, 101640, 101660, 101670, 
    101690, 101690, 101710, 101720, 101720, 101720, 101720, 101720, 101740, 
    101760, 101770, 101770, 101780, 101780, 101770, 101760, 101740, 101730, 
    101700, 101700, 101650, 101640, 101630, 101590, 101540, 101480, 101420, 
    101360, 101310, 101260, 101280, 101210, 101160, 101150, 101100, 101060, 
    101040, 101020, 100980, 100970, 100970, 100960, 101000, 101000, 101020, 
    101050, 101080, 101110, 101160, 101180, 101210, 101240, 101230, 101240, 
    101260, 101260, 101270, 101280, 101280, 101270, 101260, 101240, 101250, 
    101250, 101240, 101200, 101170, 101150, 101160, 101150, 101130, 101100, 
    101100, 101090, 101070, 101070, 101050, 101050, 101050, 101040, 101050, 
    101060, 101060, 101080, 101100, 101100, 101110, 101100, 101100, 101060, 
    101070, 101040, 101060, 101100, 101120, 101100, 101120, 101190, 101190, 
    101200, 101220, 101240, 101250, 101300, 101340, 101380, 101410, 101410, 
    101400, 101420, 101460, 101480, 101470, 101460, 101440, 101430, 101410, 
    101410, 101410, 101410, 101380, 101390, 101390, 101350, 101330, 101340, 
    101270, 101220, 101230, 101200, 101230, 101230, 101210, 101200, 101190, 
    101130, 101110, 101090, 100990, 101020, 100910, 100920, 100870, 100840, 
    100850, 100790, 100750, 100770, 100710, 100660, 100720, 100740, 100710, 
    100700, 100710, 100730, 100700, 100670, 100720, 100720, 100690, 100660, 
    100650, 100590, 100560, 100540, 100410, 100370, 100370, 100350, 100290, 
    100300, 100220, 100180, 100160, 100180, 100160, 100090, 100090, 100090, 
    100070, 100070, 100090, 100090, 100090, 100070, 100060, 100050, _, 
    100120, 100140, 100170, 100240, 100320, 100330, 100340, 100370, 100390, 
    100400, 100420, 100460, 100520, 100560, 100590, 100620, 100650, 100680, 
    100690, 100710, 100720, 100780, 100810, 100850, 100880, 100910, 100950, 
    100970, _, 100990, 101010, 101020, 101030, 101060, 101080, 101120, 
    101150, 101160, 101180, 101210, 101220, 101220, 101220, 101210, 101200, 
    101190, 101180, 101160, 101130, 101110, _, 101000, 100950, 100890, 
    100850, 100850, 100840, 100810, 100780, 100780, 100770, 100740, 100720, 
    100700, 100630, 100550, 100450, 100380, 100270, 100220, 100180, 100110, 
    100040, 99960, 99830, 99750, 99700, 99650, 99640, 99620, 99630, 99620, 
    99630, 99600, 99640, 99640, 99660, 99660, 99640, 99640, 99650, 99640, 
    99630, 99640, 99670, 99670, 99650, 99660, 99660, 99670, 99660, 99740, 
    99780, 99780, 99810, 99920, 99980, 100020, 100050, 100120, 100170, 
    100250, 100320, 100340, 100390, 100460, 100450, 100510, 100610, 100650, 
    100690, 100760, 100830, 100890, 100920, 100970, 100960, 100920, 100930, 
    100900, 100910, 100870, 100840, 100830, 100800, 100750, 100680, 100640, 
    100610, 100560, 100550, 100530, 100510, 100530, 100530, 100570, 100600, 
    100620, 100670, 100700, 100770, 100810, 100830, 100850, 100850, 100860, 
    100840, 100850, 100820, 100760, 100680, 100610, 100540, 100470, 100440, 
    100410, 100390, 100410, 100430, 100480, 100490, 100570, 100610, 100650, 
    100700, 100780, 100810, 100880, 100950, 101010, 101080, 101140, 101160, 
    101280, 101340, 101370, 101400, 101430, 101460, 101460, 101460, 101440, 
    101430, 101430, 101390, 101310, 101260, 101220, 101150, 101090, 101050, 
    101020, 101020, 101040, 101060, 101130, 101170, 101230, 101290, 101310, 
    101340, 101370, 101400, 101460, 101490, 101540, 101580, 101610, 101620, 
    101610, 101620, 101620, 101640, 101610, 101580, 101540, 101520, 101510, 
    101480, 101470, 101420, 101400, 101340, 101300, 101240, 101240, 101210, 
    101180, 101120, 101080, 101080, 101050, 101010, 100950, 100970, 100940, 
    100950, 100990, 101050, 101110, 101160, 101250, 101300, 101340, 101390, 
    101460, 101510, 101560, 101550, 101590, 101640, 101670, 101680, 101720, 
    _, 101740, 101740, 101720, 101720, 101710, 101700, 101670, 101690, 
    101690, 101640, 101630, 101620, 101580, 101560, 101560, 101560, 101510, 
    101480, 101440, 101420, 101390, 101330, 101280, 101210, 101180, 101120, 
    101110, 101020, 100970, 100940, 100910, 100920, 100910, 100900, 100900, 
    100900, 100870, 100890, 100920, 100930, 100950, 100960, 100930, 100940, 
    101020, 101120, 101160, 101180, 101190, 101200, 101210, 101240, 101240, 
    101250, 101290, 101350, 101360, 101360, 101330, 101390, 101470, 101550, 
    101570, 101610, 101630, 101650, 101670, 101660, 101670, 101710, 101680, 
    101680, 101680, 101670, 101680, 101710, 101700, 101670, 101690, 101700, 
    101680, 101660, 101670, 101680, 101680, 101690, 101680, 101640, 101620, 
    101570, 101550, 101500, 101480, 101460, 101420, 101350, 101350, 101330, 
    101280, 101270, 101230, 101190, 101150, 101120, 101080, 101070, 101060, 
    101060, 101070, 101060, 101070, 101060, 101060, 101060, 101040, 101030, 
    101030, 101050, 101050, 101070, 101100, 101160, 101170, 101190, 101230, 
    101250, 101290, 101300, 101320, 101340, 101380, 101410, 101470, 101510, 
    101540, 101600, 101610, 101620, 101640, 101670, 101640, 101690, 101700, 
    101710, 101700, 101670, 101640, 101610, 101540, 101530, 101450, 101370, 
    101340, 101280, 101200, 101200, 101180, 101150, 101120, 101090, 101040, 
    101000, 100940, 100890, 100830, 100860, 100830, 100810, 100790, 100770, 
    100810, 100780, 100790, 100810, 100820, 100870, 100900, 100930, 100960, 
    101010, 101020, 101090, 101110, 101150, 101170, 101240, 101250, 101240, 
    101290, 101320, 101400, 101400, 101430, 101450, 101460, 101480, 101480, 
    101470, 101480, 101480, 101470, 101500, 101500, 101510, 101490, 101500, 
    101490, 101460, 101440, 101420, 101400, 101390, 101370, 101370, _, 
    101320, 101320, _, 101270, 101270, 101250, 101250, 101240, 101250, 
    101250, 101270, 101280, 101290, 101310, 101330, 101340, 101360, 101360, 
    101380, 101420, 101430, 101450, _, _, _, _, _, _, _, 101690, 101720, 
    101780, 101810, 101840, 101890, 101940, 102000, 102030, 102060, 102100, 
    102130, 102140, 102180, 102210, 102240, 102270, 102300, 102340, 102380, 
    102410, 102460, 102480, 102500, 102540, 102590, 102630, 102660, 102660, 
    102710, 102760, 102780, 102800, 102830, 102840, 102850, 102850, 102840, 
    102840, 102840, 102800, 102750, 102690, 102660, 102630, 102600, 102550, 
    102520, 102500, 102430, 102380, 102330, 102230, 102170, 102070, 102030, 
    101950, 101880, 101840, 101760, 101720, 101630, 101560, 101450, 101380, 
    101280, 101150, 101000, 100830, 100670, 100620, 100610, 100630, 100630, 
    100600, 100460, 100310, 100190, 100120, 100020, 99900, 99790, 99610, 
    99290, 99020, 98640, 98260, 98070, 97820, 97520, 97300, 97120, 96990, 
    96830, 96690, 96550, 96390, 96260, 96150, 96050, 95940, 95910, 95890, 
    95940, 95990, 96040, 96100, 96250, 96360, 96520, 96740, 96950, 97080, 
    97250, 97350, 97460, 97560, 97630, 97720, 97830, 97890, 98020, 98100, 
    98150, 98230, 98300, 98360, 98450, 98500, 98570, 98610, 98670, 98740, 
    98780, 98810, 98930, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 102010, 
    102060, 102110, 102160, 102210, 102270, 102310, 102310, 102330, 102330, 
    102380, 102420, 102440, 102480, 102500, 102540, 102540, 102570, 102590, 
    102630, 102650, 102660, 102670, 102720, 102740, 102780, 102790, 102770, 
    102810, 102800, 102810, _, 102780, 102770, 102790, 102790, 102780, 
    102780, 102790, 102780, 102770, 102800, 102810, 102820, 102810, 102860, 
    102900, 102910, 102940, 102950, 102990, 102990, 103010, 103010, 103020, 
    103030, 103050, 103030, 103020, 103040, 103020, 103010, 102990, 102950, 
    102920, 102920, 102880, 102850, 102820, 102790, 102770, 102750, 102760, 
    102760, 102710, 102680, 102650, 102660, 102640, 102620, 102580, 102580, 
    102560, 102560, 102550, 102530, 102470, 102510, 102500, 102460, 102470, 
    102450, 102490, 102470, 102480, 102480, 102480, 102500, 102460, 102450, 
    102420, 102380, 102390, _, 102340, 102300, 102270, 102200, _, 102190, 
    102160, 102120, 102070, 102010, 102000, 101940, 101900, 101900, 101890, 
    101860, 101860, 101840, 101810, 101770, 101740, 101700, 101640, 101670, 
    101610, 101540, 101510, 101450, 101410, 101340, 101300, 101270, 101240, 
    101200, 101160, 101120, 101050, 100990, 100980, 100980, 100980, 100960, 
    100930, 100900, 100850, 100820, 100770, 100740, 100730, 100710, 100690, 
    100660, 100630, 100630, 100630, 100610, 100600, 100600, 100580, 100580, 
    100600, 100610, 100610, 100610, 100650, 100700, 100710, 100760, 100780, 
    100810, 100840, _, 100890, 100900, 100910, 100930, 100950, 100960, 
    100980, 101000, 100990, 101020, 101010, 101030, 101020, 101020, 101000, 
    101020, 101030, 101040, 101050, 101070, 101080, 101110, 101110, 101120, 
    101130, 101150, 101160, 101180, 101200, 101240, 101280, 101270, 101280, 
    101290, 101300, 101310, 101330, 101310, 101320, 101320, 101310, 101260, 
    101270, 101270, 101250, 101230, 101190, 101140, 101130, 101080, 101030, 
    101020, 100980, 100930, 100910, 100850, 100800, 100750, 100690, 100660, 
    100540, 100480, 100380, 100240, 100140, 100030, 99980, 99870, 99670, 
    99550, 99410, 99220, 99050, 98870, 98700, 98490, 98280, 98080, 97990, 
    98010, 98110, 98250, 98380, 98460, 98570, 98630, 98720, 98780, 98850, 
    98890, 99010, 99000, 99010, 99040, 99060, 99110, 99140, 99190, 99210, 
    99260, 99300, 99290, 99330, 99440, 99470, 99540, 99580, 99620, 99680, 
    99710, 99770, 99830, 99880, 99960, 100050, 100050, 100080, 100140, 
    100140, 100170, 100190, 100190, 100200, 100240, 100280, 100310, 100350, 
    100350, 100380, 100400, 100430, 100450, 100460, 100480, 100510, 100530, 
    100520, 100540, 100520, 100500, 100470, 100420, 100370, 100310, 100250, 
    _, _, 100040, 99990, 99910, 99810, 99710, _, 99500, 99370, _, 99190, 
    99140, 99100, 99080, 99070, 99060, 99050, 99000, 98960, 98960, 98960, 
    98960, 98980, 99030, 99130, 99230, 99320, 99400, 99510, 99600, 99700, 
    99760, 99810, 99870, 99930, 100020, 100070, 100100, 100170, 100230, 
    100300, 100360, 100420, 100460, 100500, 100520, 100560, 100600, 100620, 
    100640, 100660, 100670, 100690, 100700, 100730, 100730, 100720, 100720, 
    100720, 100720, 100710, 100730, 100700, 100660, 100620, 100610, 100590, 
    100550, 100510, 100460, 100440, 100410, 100390, 100350, 100330, 100310, 
    100300, 100270, 100250, 100200, 100200, 100170, 100140, 100140, 100140, 
    100130, 100120, 100100, 100070, 100090, 100100, 100090, 100110, 100080, 
    100090, 100100, 100100, 100060, 100070, 100090, 100090, 100100, 100090, 
    100110, 100110, 100120, 100130, 100160, 100150, 100180, 100220, 100230, 
    100260, 100280, 100320, 100300, 100310, 100300, _, 100280, 100280, 
    100220, 100170, 100140, 100100, 100050, 99980, 99840, 99730, 99590, 
    99570, 99450, 99300, 99240, 99150, 99180, 99180, 99150, 99090, 98980, 
    98920, 98880, 98790, 98720, 98620, 98560, 98470, 98390, 98230, 98020, 
    97780, 97720, 97590, 97600, 97550, 97510, 97520, 97490, 97470, 97400, 
    97360, 97320, 97310, 97290, 97290, 97350, 97410, 97480, 97580, 97700, 
    97820, 97880, 98020, 98080, 98070, 98200, 98180, 98290, 98440, 98650, 
    98820, 98900, 99000, 99170, 99320, 99450, 99510, 99570, 99660, 99760, 
    99870, 99910, 99990, 100060, 100110, 100150, 100210, 100250, 100280, 
    100310, 100360, 100370, 100400, 100430, 100450, 100480, 100500, 100520, 
    100550, 100560, 100540, 100520, 100530, 100500, 100490, 100470, 100460, 
    100470, 100480, 100510, 100490, 100520, 100520, 100510, 100520, 100540, 
    100600, 100640, 100670, 100720, 100760, 100780, 100840, 100900, 100950, 
    101010, 101060, 101100, 101150, 101170, 101180, 101220, 101270, 101290, 
    101320, 101330, 101370, 101410, 101450, 101460, 101490, 101530, 101550, 
    101570, 101600, 101620, 101610, 101630, 101670, 101640, 101650, 101650, 
    101660, 101660, 101690, 101670, 101690, 101650, 101650, 101610, 101600, 
    101560, 101470, 101380, 101310, 101280, 101200, 101220, 101200, 101110, 
    101080, 101060, 101050, 101050, 100980, 100990, 100970, 101000, 100990, 
    101000, 100980, 100970, 100930, 100900, 100870, 100810, 100790, 100760, 
    100720, 100680, 100600, 100590, 100580, 100550, 100480, 100430, 100400, 
    100320, 100270, 100180, 100110, 99990, 100000, 99930, 99880, 99780, 
    99740, 99650, 99530, 99450, 99370, 99280, 99200, 99080, 98950, 98890, 
    98860, 98840, 98810, 98780, 98720, 98720, 98670, 98640, 98640, 98630, 
    98620, _, 98610, 98600, 98590, 98620, 98580, 98580, 98610, 98620, 98610, 
    98640, 98670, 98670, 98670, 98630, 98660, 98690, 98710, 98750, 98750, 
    98770, 98780, 98810, 98830, 98860, 98880, 98950, 99000, 99050, 99120, 
    99190, 99250, 99290, 99330, 99450, 99480, 99500, 99560, 99610, 99650, 
    99660, 99640, 99640, 99630, 99620, 99600, 99560, 99550, 99540, 99460, 
    99450, 99420, 99410, 99400, 99380, 99340, 99300, 99280, 99290, _, 99340, 
    99390, 99410, 99440, 99490, 99540, 99600, 99670, 99730, 99760, 99820, 
    99880, 99930, 100000, 100100, 100190, 100300, 100370, 100450, 100510, 
    100550, 100620, 100690, 100750, 100780, 100810, 100870, 100890, 100900, 
    100910, 100930, 100890, 100840, 100790, 100800, 100880, 100990, 101030, 
    101040, 101050, 101040, 101010, 101000, 101040, 101090, 101130, 101190, 
    101250, 101290, 101290, 101260, 101210, 101210, 101190, 101180, 101160, 
    101150, 101130, 101140, 101110, 101090, 101070, 101030, 101020, 101000, 
    100990, 100980, 100990, 100990, 100970, 100960, 100930, 100970, 100940, 
    100910, 100880, 100830, 100800, 100740, 100660, 100590, 100540, 100470, 
    100440, 100430, 100430, 100460, 100460, 100420, 100400, 100380, 100380, 
    100320, 100280, 100290, 100270, 100190, 100120, 100090, 100040, 99990, 
    99910, 99820, 99750, 99680, 99630, 99570, 99510, 99460, 99430, 99350, 
    99250, 99210, 99220, 99280, 99330, 99340, 99400, 99410, 99420, 99500, 
    99500, 99490, 99490, 99510, 99540, 99520, 99650, 99670, 99700, 99750, 
    99740, 99760, 99770, 99800, 99800, 99850, 99880, 99860, 99870, 99870, 
    99870, 99890, 99930, 99960, 99990, 100010, 100020, 100000, 100010, 
    100040, 100060, 100080, 100090, 100080, 100110, 100160, 100170, 100200, 
    100190, 100220, 100230, 100280, 100300, 100340, 100380, 100430, 100440, 
    100510, 100620, 100710, 100760, 100820, 100880, 100940, 101000, _, 
    101080, 101090, 101180, 101220, 101270, 101340, 101390, 101420, 101480, 
    101560, 101620, 101660, 101730, 101780, 101820, 101870, 101940, 102000, 
    102060, 102090, 102130, 102200, 102270, 102300, 102360, 102400, 102430, 
    102490, 102520, 102560, 102600, 102620, 102650, 102700, 102720, 102730, 
    102720, 102740, 102750, 102770, 102780, 102790, 102790, _, 102760, 
    102760, 102730, 102720, 102710, 102660, 102640, 102600, 102550, 102510, 
    102470, 102410, 102350, 102280, 102200, 102100, 102030, 101940, 101900, 
    101860, 101830, 101790, 101750, 101710, 101660, 101580, 101530, _, 
    101400, 101370, 101320, 101270, 101230, 101150, 101030, 100980, 100940, 
    100860, 100750, 100660, 100530, 100390, 100310, 100220, 100110, 100040, 
    99910, 99870, 99790, 99760, 99710, 99670, 99640, 99630, 99630, 99610, 
    99640, 99680, 99700, 99720, 99720, 99730, 99790, 99820, 99800, 99770, 
    99780, 99770, 99790, 99770, 99740, _, 99600, _, 99490, 99450, 99420, 
    99410, 99380, 99320, 99300, 99240, 99200, 99150, 99080, 99000, 98950, 
    98980, 98960, 98940, 98950, 98990, 99030, 99040, 99080, 99090, 99090, 
    99100, 99110, _, 99120, 99140, 99150, 99190, 99210, 99240, 99240, 99230, 
    99230, 99220, 99220, 99270, 99350, 99400, 99450, 99490, 99550, 99580, 
    99610, 99620, 99640, 99660, 99730, 99780, 99820, 99860, 99890, 99900, 
    99960, 99970, 99970, 99990, 100000, 100000, 99980, 99960, 99960, 99920, 
    99890, 99850, 99840, 99800, 99740, _, 99550, 99470, 99360, 99250, 99120, 
    98980, 98880, 98720, 98590, 98480, 98420, 98340, 98270, 98200, 98150, 
    98100, 98050, 97980, 97930, 97880, 97860, 97850, 97840, 97780, 97830, 
    97870, 97950, 97980, 98060, 98130, 98210, 98280, 98430, 98580, 98680, 
    98770, 98870, 98950, 99050, 99130, 99200, 99270, 99360, 99430, 99500, 
    99530, 99570, 99600, 99620, 99660, 99680, 99700, 99730, 99760, 99740, 
    99740, 99730, 99730, 99730, 99680, 99630, 99580, 99510, 99340, 99210, 
    99160, 99090, 99050, 99010, 98960, 98930, 98900, 98840, 98790, _, 98650, 
    98580, 98440, 98300, 98370, 98360, 98350, 98370, 98390, 98420, 98450, 
    98490, 98500, 98500, 98470, 98480, 98460, 98460, 98410, _, 98410, 98430, 
    98470, 98500, 98540, 98630, 98720, 98820, 98920, 98990, 99030, 99070, 
    99110, 99150, 99150, 99160, 99150, 99130, 99150, 99120, 99220, 99230, 
    99220, 99170, 99150, 99240, 99370, 99480, 99570, 99590, 99660, 99700, 
    99710, 99720, 99740, 99740, 99770, 99810, 99810, 99820, 99830, 99830, 
    99850, 99860, 99900, 99940, 99930, 99930, 99940, 99940, 99930, 99940, 
    99900, 99890, 99910, 99920, 99910, 99920, 99900, 99870, 99850, 99800, 
    99770, 99740, 99720, 99670, 99630, 99630, 99610, 99570, 99570, _, 99510, 
    99480, 99430, 99370, _, 99290, 99220, 99160, 99130, 99100, 99080, _, 
    99030, 99000, 99000, 98980, 98950, 98980, 99050, 99050, 99090, 99150, 
    99210, 99230, 99250, 99290, 99320, 99320, 99340, 99360, 99350, 99390, 
    99430, 99450, 99480, 99480, 99490, 99510, 99500, 99500, 99490, 99480, 
    99510, 99530, 99560, 99580, 99600, 99600, 99600, 99580, 99610, 99610, 
    99620, 99620, 99650, 99620, 99600, 99570, 99600, 99620, 99620, 99630, 
    99620, 99590, 99540, 99540, 99500, 99500, 99480, 99480, 99470, _, 99300, 
    99270, 99300, 99240, 99190, 99160, 99140, 99150, 99150, 99190, 99230, _, 
    99240, 99300, 99320, 99410, 99420, 99500, 99570, 99620, 99680, 99760, 
    99850, 99930, 99970, 100020, 100080, _, 100150, 100180, 100190, 100230, 
    100210, _, 100340, 100410, 100410, 100400, _, 100460, _, 100610, 100640, 
    100660, _, _, 100730, 100740, 100760, 100770, 100800, 100800, _, _, 
    100790, _, 100810, 100790, 100790, 100810, 100820, _, 100850, 100830, 
    100840, 100820, 100820, 100800, 100800, 100770, 100750, 100710, _, 
    100680, 100660, 100660, _, 100530, _, _, 100340, 100290, 100240, 100160, 
    100050, _, 99880, 99780, 99670, 99580, _, _, _, 99170, 99090, 99010, 
    98890, 98770, 98720, 98710, 98690, 98690, 98670, 98680, 98660, 98640, 
    98610, 98540, 98480, 98350, 98240, 98240, 98300, 98280, 98190, 98140, 
    98100, 98120, 98150, 98190, 98190, 98190, 98220, 98200, 98160, 98140, 
    98130, 97970, 97970, 98160, 98260, 98230, 98270, 98280, 98330, 98320, 
    98330, 98330, 98370, 98370, 98380, 98460, 98430, 98490, 98450, 98440, 
    98500, 98390, _, 98550, 98520, 98530, 98530, 98530, 98530, 98630, 98760, 
    98750, 98730, 98750, 98640, 98570, 98560, 98560, 98570, 98580, 98600, 
    98630, 98650, 98620, 98680, 98690, 98660, 98580, 98590, 98680, _, 98890, 
    98970, 98960, 98990, 99040, 99100, 99150, 99190, 99240, 99330, 99380, 
    99420, 99480, 99490, 99520, 99560, 99610, 99650, 99720, 99790, 99840, 
    99890, 99970, 100060, 100140, 100180, 100240, 100300, 100380, 100450, 
    100480, 100540, 100580, 100610, 100650, 100690, 100730, 100790, 100800, 
    100860, 100840, 100840, 100860, _, 100850, 100830, 100840, 100840, 
    100850, 100840, _, 100810, 100790, 100770, 100730, 100700, 100670, 
    100680, 100670, 100650, 100620, 100590, 100590, 100550, 100520, 100480, 
    100450, 100460, 100420, 100380, 100340, 100310, 100300, 100270, 100220, 
    100170, 100160, 100110, 100070, 100000, 99890, 99860, 99810, 99740, 
    99660, 99560, 99430, 99350, 99270, 99140, 99080, 99010, 98960, 98890, 
    98880, 98840, 98800, 98770, 98780, 98790, 98780, 98780, 98800, 98810, 
    98830, 98900, 98970, 99070, 99130, 99190, 99220, 99220, 99220, 99230, 
    99230, 99230, 99260, 99270, 99280, 99300, 99300, 99300, _, 99300, 99320, 
    99330, 99320, 99330, 99310, 99310, 99320, 99360, 99380, 99390, 99400, 
    99400, 99390, 99410, 99420, 99430, 99450, 99410, 99430, 99430, 99410, 
    99390, 99370, 99370, 99380, 99340, 99320, 99310, 99270, 99230, 99190, 
    99200, 99230, 99230, 99230, 99180, 99110, 99110, 99080, 99060, 99060, 
    99030, 99050, 99060, 99090, 99120, 99140, 99160, 99170, 99210, 99240, 
    99270, 99290, 99300, 99330, 99370, 99420, 99430, 99410, 99480, 99510, 
    99520, 99550, 99570, 99630, 99640, 99670, 99730, 99780, 99780, 99840, 
    99790, 99780, 99810, 99780, 99700, 99720, 99700, 99710, 99740, 99770, 
    99840, 99890, 99900, 100030, 100070, 100190, 100300, 100340, 100400, 
    100460, 100500, 100550, 100620, 100690, 100740, 100810, 100860, 100950, 
    101010, 101100, 101210, 101320, 101360, 101340, 101350, 101440, 101440, 
    101470, 101540, 101660, 101750, 101800, 101780, 101820, 101850, 101900, 
    101990, 101990, 102010, 101970, 102050, 102070, 102080, 102060, 102060, 
    102060, 102080, 102100, 102070, 102060, 102070, 102050, 102040, 102010, 
    101990, 101960, 101870, 101790, 101820, 101730, 101610, 101640, 101590, 
    101520, 101370, 101270, 101260, 101130, 101080, 101050, 101020, 100970, 
    100920, 100870, 100700, 100610, 100610, 100590, 100450, 100390, 100300, 
    100330, 100260, 100170, 100010, 99920, 99900, 99810, 99720, 99650, 99650, 
    99600, 99560, 99580, 99580, 99460, 99360, 99320, 99210, 99150, 99100, 
    99060, 99020, 98880, 98810, 98750, 98710, 98680, 98650, 98530, 98490, 
    98320, 98390, 98350, 98360, 98290, 98240, 98160, 98000, 97970, 98000, 
    97980, 97970, 97910, 97810, 97710, 97660, 97620, 97570, 97520, 97450, 
    97400, 97320, 97270, 97280, 97230, 97130, 97030, 97130, 97060, 97030, 
    96970, 96960, 96970, 96910, 96890, 96780, 96770, 96800, 96800, 96840, 
    96830, _, 96840, _, _, _, 96950, _, _, 97130, _, 97300, 97400, 97470, 
    97580, 97680, _, _, 98000, 98040, 98140, 98190, 98260, _, _, 98460, 
    98510, _, _, 98710, _, _, _, 99000, 99030, 99090, _, 99150, _, 99260, 
    99310, 99330, _, _, _, _, 99400, 99350, 99340, 99290, _, 99150, 99010, 
    98870, 98690, _, 98520, _, _, 98330, 98280, 98230, 98190, 98160, 98160, 
    _, 98080, _, 97970, 97900, _, _, 97700, 97610, 97550, 97500, 97490, 
    97490, 97490, 97540, 97540, 97580, _, 97550, 97560, 97610, 97510, 97520, 
    97510, 97500, 97450, 97430, 97400, 97350, 97300, 97270, 97250, 97240, 
    97270, 97270, _, 97350, 97440, 97470, 97510, 97580, 97620, 97640, 97700, 
    97700, 97800, 97830, 97890, 97900, 97960, _, 97890, 97870, 97820, _, 
    97780, 97800, 97790, 97820, _, 97870, 97870, 97930, _, _, 98170, _, 
    98390, 98480, 98540, 98730, 98930, 99110, _, _, 99600, 99710, 99810, _, 
    100090, 100180, _, _, 100530, 100670, _, 100770, 100860, 100950, 100950, 
    _, 100910, 100880, _, 100820, _, 100760, _, 100860, 100910, 100970, 
    101040, 101140, 101190, 101260, 101310, 101370, 101420, 101480, _, 
    101550, 101590, 101640, 101620, 101610, _, 101550, 101500, 101450, 
    101400, _, 101260, 101200, 101180, 101120, 101080, 101040, 101000, 
    100950, 100920, 100870, 100870, 100780, _, 100610, 100470, _, 100380, 
    100370, 100370, 100310, 100350, 100250, 100130, 100140, _, _, 100220, 
    100210, _, 100370, 100480, 100480, 100520, _, _, 100540, 100560, 100560, 
    _, 100540, 100520, 100550, 100330, 100260, 100010, 99980, 100010, 99980, 
    99950, 100350, 100480, _, 100650, _, _, 100860, 100900, 100970, 101020, 
    101010, 100980, 100980, _, _, _, 100720, 100710, _, 100410, 100460, 
    100430, _, 100500, _, 100550, _, 100650, 100770, 100760, 100750, 100760, 
    _, _, 100780, 100720, _, 100600, _, _, _, 100430, _, _, _, 101140, 
    101330, _, 101700, _, _, 102000, 102060, 102070, 102060, 102030, 102030, 
    101990, 101900, _, 101760, 101680, 101580, _, _, 101390, 101320, _, _, 
    101210, _, 101200, _, _, 101190, _, 101200, 101190, 101160, _, _, 101130, 
    101110, 101090, 101070, 101060, 101090, 101130, 101170, 101240, 101310, 
    101400, 101480, 101510, 101600, _, 101720, _, 101840, _, 101930, 101980, 
    102010, _, 102090, 102110, 102130, _, 102130, 102120, 102100, _, _, _, _, 
    _, _, _, 101980, 101980, 101950, 101940, 101920, 101910, 101860, 101850, 
    101840, 101830, 101810, 101840, 101830, 101820, 101810, 101820, 101790, 
    101810, 101840, 101830, 101870, 101910, 101920, 101960, 101960, 102030, 
    102050, 102110, 102170, 102200, 102200, 102230, 102260, 102280, 102310, 
    102350, 102360, 102340, 102340, 102330, 102310, 102300, 102270, 102240, 
    102220, 102200, 102180, 102150, 102170, 102180, 102180, 102180, 102210, 
    102210, 102200, 102200, 102190, 102190, 102210, 102220, 102220, 102240, 
    102260, 102250, 102240, 102260, 102250, 102240, 102260, 102270, 102270, 
    102290, 102300, 102310, 102320, 102330, 102330, 102340, 102340, 102330, 
    102320, 102340, 102330, 102340, 102340, 102330, 102310, 102290, 102290, 
    102290, 102300, 102310, 102300, 102300, 102300, 102300, 102310, 102300, 
    102280, 102300, 102290, 102280, 102270, 102260, 102260, 102260, 102280, 
    102300, 102350, 102350, 102370, 102380, 102400, 102420, 102430, 102440, 
    102460, 102480, 102520, 102550, 102600, 102630, 102650, 102690, 102720, 
    102740, 102770, 102800, 102810, 102860, 102920, 102970, 102990, 103030, 
    103060, 103120, 103140, 103160, 103200, 103220, 103230, 103260, 103300, 
    103330, 103360, 103370, 103370, 103380, 103390, 103390, 103380, 103370, 
    103370, 103340, 103330, 103310, 103260, 103240, 103190, 103110, 103080, 
    103040, 102980, 102880, 102790, 102650, 102530, 102440, 102330, 102210, 
    102080, 101930, 101830, 101710, 101610, 101530, 101470, 101430, 101420, 
    101420, 101420, 101390, 101380, 101330, 101280, 101250, 101200, 101150, 
    101100, 101020, 100970, 100900, 100860, 100800, 100790, 100790, 100790, 
    100780, 100760, 100760, 100730, 100700, 100700, 100740, 100800, 100810, 
    100790, 100790, 100800, 100830, 100880, 100900, 100920, 100950, 100960, 
    100980, 101020, 101040, 101010, 100920, 100900, 100940, 101030, 101120, 
    101200, 101320, 101420, 101520, 101620, 101690, 101730, 101760, 101820, 
    101880, 101910, 101950, 101960, 101980, 102020, 102060, 102070, 102090, 
    102130, 102130, 102120, 102070, 102120, 102150, 102170, 102230, 102260, 
    102280, 102310, 102350, 102340, 102340, 102380, 102390, 102410, 102430, 
    102430, 102410, 102390, 102380, 102370, 102350, 102320, 102290, 102290, 
    102310, 102310, 102270, 102270, 102230, 102120, 102170, 102200, 102140, 
    102120, 102080, 102070, 102000, 101960, 101970, 101970, 101970, 101960, 
    101940, 101890, 101960, 101930, 101910, 101820, 101800, 101790, 101770, 
    101730, 101700, 101680, 101670, 101700, 101730, 101760, 101760, 101740, 
    101750, 101750, 101760, 101750, 101720, 101720, 101730, 101730, 101720, 
    101680, 101670, 101640, 101610, 101590, 101570, 101550, 101540, 101520, 
    101490, 101460, 101430, 101380, 101330, 101290, 101260, 101220, 101180, 
    101140, 101120, 101070, 101050, 101010, 100980, 100940, 100920, 100870, 
    100840, 100800, 100780, 100760, 100730, 100700, 100690, 100700, 100690, 
    100670, 100640, 100610, 100600, 100580, 100550, 100540, 100530, 100530, 
    100530, 100530, 100530, 100550, 100540, 100560, 100570, 100550, 100570, 
    100560, 100540, 100550, 100550, 100550, 100530, 100460, 100370, 100300, 
    100210, 100210, 100250, 100250, 100260, 100250, 100230, 100250, 100240, 
    100210, 100170, 100140, 100100, 100080, 100040, 100010, 99960, 99910, 
    99890, 99850, 99840, 99840, 99860, 99890, 99920, 99960, 100010, 100050, 
    100090, 100100, 100160, 100200, 100200, 100210, 100210, 100170, 100170, 
    100170, 100180, 100190, 100170, 100250, 100310, 100380, 100400, 100450, 
    100540, 100560, 100610, 100630, 100710, 100730, 100730, 100770, 100840, 
    100880, 100890, 100900, 100920, 100960, 100970, 101000, 101020, 101020, 
    101050, 101090, 101100, 101150, 101170, 101200, 101200, 101200, 101240, 
    101260, 101280, 101290, 101350, 101360, 101390, 101450, 101510, 101490, 
    101460, 101490, 101510, 101470, 101500, 101530, 101530, 101520, 101560, 
    101570, 101580, 101640, 101630, 101630, 101670, 101670, 101690, 101730, 
    101730, 101730, 101760, 101750, 101750, 101750, 101710, 101660, 101620, 
    101570, 101530, 101480, 101390, 101370, 101310, 101260, 101210, 101180, 
    101140, 101080, 101030, 100960, 100870, 100780, 100690, 100590, 100530, 
    100420, 100350, 100280, 100160, 100050, 99920, 99790, 99650, 99530, 
    99510, 99470, 99430, 99390, 99350, 99310, 99280, 99230, 99270, 99240, 
    99190, 99130, 99120, 99090, 99080, 99090, 99060, 99040, 99030, 99010, 
    99030, 99020, 98970, 98920, 98880, 98850, 98850, 98870, 98860, 98810, 
    98770, 98690, 98680, 98650, 98540, 98490, 98430, 98420, 98260, 98370, 
    98180, 98050, 97910, 97870, 97810, 97810, 97810, 97790, 97830, 97870, 
    97910, 97970, 98000, 98010, 98070, 98130, 98190, 98230, 98280, 98280, 
    98300, 98320, 98380, 98490, 98520, 98570, 98590, 98580, 98620, 98670, 
    98710, 98760, 98840, 98890, 98940, 98900, 98890, 98890, 98920, 98880, 
    98860, 98890, 98890, 98980, 99070, 99100, 99140, 99170, 99180, 99130, 
    99060, 99020, 99000, 98950, 98890, 98910, 98890, 98900, 98950, 98870, 
    98860, 98910, 98990, 99030, 99100, 99090, 99130, 99130, 99140, 99170, 
    99190, 99150, 99100, 99210, 99360, 99430, 99390, 99320, 99300, 99250, 
    99280, 99390, 99440, 99530, 99550, 99570, 99600, 99620, 99650, 99680, 
    99700, 99690, 99710, 99640, 99660, 99700, 99700, 99690, 99730, 99780, 
    99770, 99810, 99790, 99830, 99500, 99460, 99570, 99760, 99980, 100010, 
    100030, 100070, 100070, 100090, 100090, 100070, 100050, 100070, 100100, 
    100150, 100220, 100270, 100280, 100300, 100270, 100330, 100400, 100470, 
    100430, 100520, 100570, 100590, 100620, 100590, 100450, 100520, 100640, 
    100650, 100690, 100620, 100590, 100570, 100970, 101280, 101310, 101340, 
    101360, 101360, 101300, 101350, 101270, 101410, 101440, 101380, 101360, 
    101390, 101440, 101400, 101350, 101330, 101270, 101240, 101210, 101110, 
    101130, 101100, 101070, 101050, 101030, 100990, 100960, 100910, 100860, 
    100830, 100760, 100690, 100630, 100650, 100650, _, 100620, 100610, 
    100590, 100560, 100580, 100570, 100590, 100590, 100580, 100550, 100550, 
    100530, 100510, 100500, 100500, 100480, 100470, 100430, 100390, 100380, 
    100360, 100350, 100370, 100350, 100370, 100380, 100360, 100350, 100340, 
    100320, 100310, 100310, _, 100270, 100280, 100290, 100310, 100330, 
    100350, 100360, 100370, 100380, 100370, 100380, 100390, 100400, 100420, 
    100460, 100480, 100490, 100500, _, 100500, 100480, 100470, 100480, 
    100490, 100500, 100520, 100530, 100510, 100490, 100470, 100440, 100430, 
    100390, 100360, 100340, 100310, 100270, 100250, 100220, 100170, 100090, 
    100040, 99920, 99870, 99820, 99740, 99640, 99590, 99440, _, 99270, 99050, 
    98970, 98920, 98860, 98700, 98740, 98680, 98650, _, 98530, 98460, 98360, 
    98230, 98110, 98080, 98000, 97880, 97780, 97690, 97620, 97570, 97580, 
    97520, 97500, 97450, 97420, 97370, 97400, 97390, 97350, 97350, 97290, 
    97310, 97340, 97360, 97400, 97450, 97490, 97510, 97530, 97610, 97690, 
    97780, 97860, 97950, 98060, 98130, 98220, 98280, 98350, 98400, 98470, 
    98500, 98520, 98540, 98570, 98610, 98680, 98740, 98780, 98840, 98870, 
    98900, 98930, 98960, 98990, 99040, 99080, 99130, 99180, 99220, 99270, 
    99320, 99370, 99410, 99450, 99510, 99540, 99570, 99620, 99660, 99720, 
    99780, 99840, 99860, 99890, 99920, 99940, 99970, 100000, 100030, 100030, 
    100040, 100040, 100070, 100090, 100100, 100110, 100110, 100100, 100090, 
    100080, 100080, 100070, 100080, 100090, 100110, 100120, 100120, 100100, 
    100110, 100130, 100190, 100240, 100280, 100370, 100410, 100470, 100520, 
    100590, 100660, 100730, 100790, 100820, 100850, 100880, 100920, 100960, 
    101000, 101040, 101070, 101170, 101180, 101220, 101280, 101340, 101390, 
    101430, 101460, 101510, 101550, 101600, 101640, 101690, 101690, 101690, 
    101660, 101660, 101670, 101670, 101630, 101590, 101570, 101560, 101580, 
    101580, 101590, 101570, 101520, 101500, 101490, 101460, 101430, 101410, 
    101410, 101430, 101440, 101410, 101350, 101350, 101340, 101320, 101290, 
    101280, 101240, 101260, 101230, 101220, 101180, 101150, 101140, 101120, 
    101110, 101120, 101110, 101090, 101050, 101050, 101020, 101040, 101040, 
    101020, 101020, 100970, 100950, 100970, 100960, 100950, 100910, 100910, 
    100870, 100820, 100770, 100760, 100780, 100780, 100700, 100650, 100620, 
    100570, 100520, 100470, 100390, 100330, 100290, 100260, 100250, 100250, 
    100260, 100310, 100330, 100350, 100400, 100430, 100480, 100510, 100550, 
    100570, 100580, 100580, 100600, 100590, 100600, 100580, 100580, 100540, 
    100570, 100480, 100510, 100540, 100490, 100460, 100400, 100360, 100320, 
    100270, 100230, 100180, 100080, 100010, 99970, 99900, 99770, 99670, 
    99530, 99440, 99340, 99280, 99230, 99150, 99090, 99060, 99070, 99110, 
    99110, 99110, 99110, 99140, _, 99180, 99190, 99180, 99180, 99190, 99200, 
    99220, 99240, 99270, 99290, 99330, 99340, 99350, 99330, 99350, 99370, 
    99420, 99460, 99520, 99580, 99610, 99620, 99660, 99710, 99780, 99840, 
    99930, 99970, 100060, 100140, 100220, 100300, 100350, 100400, 100430, 
    100440, 100460, 100440, 100410, 100420, 100390, 100380, 100320, 100270, 
    100210, 100160, 100130, 100080, 100010, 99990, 100010, 100030, 100050, 
    100090, 100140, 100190, 100210, 100250, 100260, 100300, 100330, 100390, 
    100430, 100480, 100520, 100570, 100620, 100650, 100680, 100720, 100760, 
    _, 100820, 100850, 100870, 100890, 100890, 100900, 100960, 100990, 
    100960, 100990, _, 101000, 101030, 101030, 101050, 101080, 101140, 
    101210, 101280, 101330, 101360, 101370, 101420, 101450, 101480, 101520, 
    101530, 101540, 101550, 101570, 101590, 101590, 101580, 101570, 101560, 
    101540, 101540, 101540, 101530, 101530, 101510, 101460, 101490, 101510, 
    101520, 101490, 101480, 101470, 101470, 101430, 101420, 101420, 101450, 
    101440, 101460, 101440, 101440, 101420, 101420, 101420, 101420, 101440, 
    101450, 101470, 101450, 101460, 101440, 101450, 101450, 101420, 101420, 
    101410, 101410, 101390, 101410, 101420, 101430, 101420, 101430, 101450, 
    101450, 101430, 101410, 101400, 101380, 101380, 101350, 101340, 101330, 
    101310, 101300, 101280, 101250, 101220, 101180, 101140, 101130, 101100, 
    101070, 101050, 101020, 101010, 100990, 100970, 100940, 100930, 100890, 
    100870, 100840, 100810, 100770, 100770, 100760, 100740, 100730, 100700, 
    100710, 100690, 100660, 100640, 100650, 100650, 100630, 100620, 100620, 
    100630, 100640, 100660, 100660, 100650, 100660, 100660, 100660, 100650, 
    100640, 100630, 100630, 100600, 100620, 100630, 100610, 100610, 100600, 
    100570, 100570, 100570, 100600, 100610, 100610, 100640, 100650, 100650, 
    100670, 100650, 100650, 100640, 100640, 100650, 100620, 100610, 100630, 
    100580, 100570, 100580, 100560, 100550, 100530, 100520, 100510, 100510, 
    100530, 100540, 100550, 100530, 100550, 100530, 100500, 100480, 100440, 
    100380, 100300, 100320, 100330, 100280, 100320, 100360, 100370, 100320, 
    100340, 100400, 100400, 100380, 100360, 100310, 100250, 100120, 100080, 
    100130, 100180, 100180, 100200, 100210, 100210, 100220, 100280, 100330, 
    100390, 100430, 100500, 100570, 100600, 100630, 100660, 100670, 100660, 
    100630, 100670, 100660, 100640, 100620, 100630, 100620, 100630, 100640, 
    100690, 100690, 100670, 100680, 100670, 100660, 100640, 100600, 100600, 
    100590, 100600, 100650, 100680, 100720, 100720, 100720, 100720, 100720, 
    100710, 100700, 100690, 100690, 100660, 100700, 100690, 100670, 100640, 
    100610, 100550, 100530, 100500, 100450, 100400, 100340, 100310, 100260, 
    100180, 100100, 100040, 99960, 99910, 99880, 99870, 99870, 99860, 99920, 
    99990, 100040, 100060, 100070, 100020, 100020, 99980, 99980, 99970, 
    99970, 99980, 100030, 100080, 100130, 100190, 100240, 100280, 100340, 
    100360, 100400, 100440, 100480, 100470, 100510, 100540, 100580, 100590, 
    100590, 100590, 100580, 100590, 100600, 100610, 100630, 100640, 100660, 
    100700, 100740, 100770, 100840, 100880, 100900, 100960, 100990, 101030, 
    101050, 101060, 101100, 101100, 101120, 101120, 101130, 101130, 101120, 
    101130, 101130, 101140, 101140, 101170, 101170, 101180, 101150, 101170, 
    101190, 101160, 101150, 101150, 101190, 101220, 101250, 101260, 101290, 
    101340, 101360, 101400, 101400, 101420, 101440, 101480, 101500, 101530, 
    101580, 101590, 101560, 101550, 101570, 101650, 101690, 101700, 101700, 
    101710, 101720, 101730, 101740, 101760, 101760, 101770, 101750, 101730, 
    101730, 101680, 101610, 101540, 101500, 101460, 101440, 101410, 101370, 
    101330, 101270, 101230, 101200, 101180, 101120, 101070, 101070, 101060, 
    101020, 100990, 101000, 101000, 100990, 101000, 101020, 101050, 101040, 
    101050, 101040, 101060, 101090, 101100, 101120, 101140, 101150, 101140, 
    101170, 101180, 101180, 101220, 101210, 101230, 101240, 101230, 101220, 
    101180, 101170, 101130, 101110, 101080, 101050, 100980, 100940, 100890, 
    100820, 100800, 100740, 100700, 100670, 100610, 100600, 100560, 100540, 
    100470, 100400, 100340, 100290, 100340, 100320, 100330, 100340, 100360, 
    100400, 100380, 100390, 100430, 100420, 100450, 100430, 100430, 100440, 
    100460, 100420, 100390, 100370, 100320, 100260, 100230, 100170, 100120, 
    100040, 99970, 99850, 99780, 99600, 99410, 99270, 99110, 98960, 98880, 
    98820, 98830, 98810, 98840, 98860, 98890, 98880, 98940, 98940, 99030, 
    99070, 99230, 99450, 99520, 99660, 99800, 99940, 100080, 100110, 100140, 
    100230, 100190, 100130, 100080, 99990, 99890, 99780, 99570, 99360, 99110, 
    98880, 98710, 98470, 98350, 98260, 98250, 98250, 98370, 98420, 98520, 
    98680, 98790, 98890, 99030, 99140, 99300, 99440, 99480, 99570, 99630, 
    99690, 99770, 99850, 99890, 99940, 99900, 99960, 100000, 100040, 100040, 
    100010, 100010, 100010, 100010, 100010, 99990, 100010, 99990, 99970, 
    99960, 99950, 99950, 99990, 100010, 100010, 100040, 100110, 100150, 
    100200, 100250, 100300, 100360, 100430, 100490, 100530, 100560, 100620, 
    100680, 100720, 100740, 100780, 100820, 100860, 100900, 100940, 100950, 
    100920, 100900, 100940, 100850, 100800, 100820, 100760, 100690, 100670, 
    100670, 100640, 100720, 100730, 100730, 100720, 100740, 100740, 100780, 
    100780, 100820, 100820, 100780, 100800, 100830, 100800, 100740, 100740, 
    100730, 100780, 100790, 100780, 100730, 100700, 100670, 100640, 100600, 
    100570, 100550, 100500, 100480, 100480, 100510, 100540, 100550, 100540, 
    100540, 100570, 100540, 100560, 100580, 100610, 100630, 100630, 100670, 
    100700, 100720, 100700, 100670, 100680, 100680, 100710, 100730, 100710, 
    100670, 100690, 100680, 100710, 100710, 100710, 100700, 100700, 100680, 
    100690, 100650, 100640, 100620, 100610, 100600, 100510, 100430, 100390, 
    100400, 100410, 100360, 100310, 100290, 100280, 100220, 100200, 100220, 
    100220, 100210, 100210, 100190, 100180, 100200, 100160, 100150, 100150, 
    100140, 100130, 100150, 100140, 100130, 100130, 100130, 100120, 100140, 
    100130, 100140, 100140, 100150, 100170, 100220, 100250, 100270, 100260, 
    100300, 100320, 100360, 100400, 100420, 100450, 100470, 100480, 100520, 
    100540, 100550, 100560, 100560, 100590, 100580, 100610, 100620, 100620, 
    100620, 100620, 100620, 100630, 100650, 100650, 100660, 100670, 100690, 
    100700, 100710, 100720, 100720, 100740, 100740, 100750, 100750, 100760, 
    100750, 100760, 100760, 100760, 100770, 100760, 100760, 100770, 100790, 
    100810, 100810, 100800, 100810, 100800, 100810, 100820, 100810, 100800, 
    100770, 100780, 100770, 100750, 100740, 100720, 100680, 100610, 100550, 
    100440, 100410, 100390, 100390, 100390, 100390, 100380, 100380, 100370, 
    100340, 100320, 100290, 100240, 100220, 100210, 100250, 100240, 100280, 
    100300, 100310, 100310, 100340, 100360, 100380, 100390, 100410, 100410, 
    100400, 100430, 100440, 100470, 100470, 100450, 100420, 100410, 100400, 
    100380, 100360, 100340, 100310, 100300, 100300, 100270, 100280, 100260, 
    100240, 100230, 100230, 100190, 100140, 100100, 100050, 100020, 100010, 
    99950, 99870, 99810, 99760, 99670, 99610, 99540, 99450, 99360, 99270, 
    99180, 99120, 99080, 98950, 98810, 98670, 98460, 98330, 98280, 98290, 
    98250, 98250, 98200, 98150, 98090, 98020, 97990, 97940, 97900, 97890, 
    97920, 97950, 97960, 97850, 97870, 98000, 98180, 98170, 98320, 98330, 
    98290, 98320, 98350, 98400, 98440, 98500, 98510, 98600, 98690, 98710, 
    98730, 98810, 98990, 99070, 99120, 99170, 99220, 99260, 99280, 99280, 
    99330, 99330, 99330, 99330, 99310, 99290, 99290, 99290, 99300, 99330, 
    99330, 99350, 99340, 99360, 99360, 99340, 99350, 99360, 99360, 99360, 
    99380, 99390, 99370, 99370, 99380, 99410, 99430, 99430, 99430, 99460, 
    99480, 99510, 99520, 99560, 99600, 99620, 99650, 99710, 99730, 99770, 
    99820, 99830, 99830, 99880, 99930, 99980, 100000, 100010, 100070, 100110, 
    100180, 100230, 100270, 100300, 100320, 100360, 100420, 100470, 100540, 
    100610, 100670, 100730, 100810, 100850, 100910, 100930, 100980, 101010, 
    101040, 101090, 101130, 101180, 101240, 101270, 101300, 101320, 101340, 
    101350, 101380, 101420, 101450, 101460, 101470, 101490, 101490, 101520, 
    101520, 101510, 101520, 101520, 101520, 101520, 101500, 101520, 101520, 
    101520, 101510, 101530, 101490, 101500, 101480, 101490, 101470, 101440, 
    101430, 101430, 101450, 101480, 101490, 101500, 101500, 101500, 101470, 
    101470, 101460, 101490, 101510, 101520, 101540, 101570, 101590, 101590, 
    101610, 101610, 101620, 101610, 101630, 101650, 101660, 101650, 101710, 
    101750, 101770, 101780, 101770, 101780, 101780, 101780, 101790, 101810, 
    101820, 101850, 101870, 101900, 101900, 101890, 101860, 101840, 101840, 
    101820, 101820, 101810, 101770, 101760, 101760, 101770, 101760, 101720, 
    101710, 101690, 101650, 101620, 101600, 101590, 101550, 101530, 101500, 
    101480, 101470, 101460, 101430, 101390, 101380, 101350, 101350, 101350, 
    101350, 101340, 101350, 101360, 101380, 101380, 101390, 101410, 101450, 
    101440, 101470, 101480, 101520, 101520, 101510, 101510, 101510, 101500, 
    101490, 101520, 101530, 101540, 101560, 101560, 101580, 101610, 101630, 
    101650, 101640, 101650, 101670, 101670, 101660, 101670, 101710, 101720, 
    101750, 101760, 101770, 101800, 101820, 101830, 101830, 101820, 101830, 
    101840, 101830, 101830, 101820, 101810, 101810, 101810, 101790, 101770, 
    101700, 101690, 101660, 101670, 101670, 101650, 101630, 101610, 101590, 
    101570, 101570, 101530, 101470, 101460, 101440, 101400, 101370, 101340, 
    101340, 101310, 101280, 101250, 101250, 101220, 101170, 101140, 101110, 
    101110, 101100, 101070, 101030, 101010, 101030, 101070, 101090, 101130, 
    101140, 101190, 101230, 101290, 101310, 101320, 101340, 101360, 101360, 
    101350, 101310, 101270, 101240, 101220, 101230, 101250, 101260, 101260, 
    101260, 101250, 101270, 101290, 101250, 101240, 101230, 101190, 101180, 
    101100, 101040, 100950, 100920, 100910, 100850, 100880, 100830, 100830, 
    100860, 100900, 100940, 100970, 100980, 100970, 100970, 101000, 101010, 
    101050, 101110, 101090, 101110, 101110, 101120, 101120, 101140, 101120, 
    101160, 101210, 101220, 101250, 101260, 101270, 101280, 101320, 101300, 
    101260, 101210, 101150, 101220, 101210, 101200, 101170, 101130, 101140, 
    101060, 101030, 101000, 100940, 100870, 100830, 100780, 100790, 100770, 
    100770, 100800, 100770, 100780, 100780, 100760, 100740, 100690, 100660, 
    100670, 100630, 100570, 100530, 100590, 100620, 100580, 100550, 100570, 
    100550, 100610, 100610, 100710, 100740, 100760, 100760, 100790, 100800, 
    100810, 100870, 100840, 100860, 100870, 100870, 100950, 100990, 100940, 
    100930, 100980, 100970, 100950, 100990, 100970, 100970, 100960, 100960, 
    100970, 100990, 100990, 101040, 101060, 101020, 101000, 101010, 100980, 
    100970, 100990, 100990, 101110, 101090, 101110, 101100, 101100, 101060, 
    101120, 101180, 101180, 101160, 101180, 101210, 101200, 101230, 101240, 
    101260, 101270, 101290, 101300, 101320, 101330, 101350, 101350, 101360, 
    101370, 101400, 101420, 101420, 101420, 101410, 101390, 101390, 101390, 
    101370, 101350, 101360, 101350, 101350, 101340, 101330, 101320, 101320, 
    101300, 101290, 101280, 101270, 101240, 101230, 101220, 101190, 101170, 
    101150, 101130, 101120, 101120, 101090, 101050, 101030, 101000, 100970, 
    100950, 100910, 100880, 100810, 100730, 100670, 100560, 100500, 100430, 
    100340, 100280, 100220, 100160, 100040, 99990, 99930, 99890, 99810, 
    99760, 99720, 99640, 99540, 99500, 99510, 99490, 99490, 99490, 99500, 
    99510, 99520, 99530, 99550, 99550, 99550, 99580, 99600, 99610, 99630, 
    99650, 99670, 99680, 99700, 99730, 99750, 99780, 99790, 99820, 99860, 
    99910, 99930, 99960, 99990, 100070, 100130, 100160, 100270, 100380, 
    100420, 100500, 100550, 100590, 100630, 100670, 100700, 100750, 100800, 
    100870, 100960, 101000, 101040, 101100, 101130, 101210, 101280, 101350, 
    101420, 101490, 101560, 101640, 101680, 101750, 101770, 101800, 101840, 
    101880, 101910, 101950, 101990, 102020, 102030, 102000, 102010, 102010, 
    102010, 101980, 101970, 101980, 101940, 101940, 101900, 101830, 101790, 
    101760, 101710, 101700, 101700, 101700, 101650, 101640, 101630, 101610, 
    _, 101610, 101620, 101610, 101590, 101580, 101530, 101500, 101460, 
    101450, 101430, _, 101350, 101310, _, 101230, 101180, 101130, 101130, 
    101090, 101060, 101000, 100990, 101000, 100980, 100960, 101000, 101040, 
    101050, 101070, 101090, 101110, 101140, 101200, 101270, 101340, 101390, 
    101460, 101520, 101560, 101600, 101650, 101670, 101710, 101730, 101760, 
    101790, 101830, 101850, 101870, 101870, 101820, 101850, 101910, 101930, 
    101880, 101890, 101900, 101950, 102010, 102060, 102130, 102180, 102280, 
    102320, 102370, 102460, 102540, 102630, 102750, 102880, 103000, _, 
    103170, 103240, 103320, 103380, 103470, 103540, 103610, 103690, 103730, 
    103800, _, 103860, 103890, 103940, 103970, 103970, 103960, 103980, 
    104000, 104020, 104020, 104060, 104040, 104010, 103990, 103960, 103910, 
    103900, 103870, 103810, 103780, 103700, 103740, 103630, 103690, 103660, 
    103640, 103640, 103630, 103610, 103600, 103580, 103560, 103560, 103530, 
    103510, _, 103480, 103470, 103440, 103410, 103350, 103280, 103240, 
    103190, 103150, 103120, 103090, 103060, 103010, 102970, 102950, 102910, 
    102860, 102880, 102870, 102860, 102870, 102890, 102900, 102930, _, 
    103030, 103050, 103080, 103120, 103130, 103170, 103170, 103220, 103250, 
    103270, 103310, 103340, 103370, 103380, 103370, 103380, 103390, 103350, 
    103330, 103280, 103260, 103230, 103190, _, 103140, 103130, 103160, 
    103150, 103130, 103130, 103110, 103120, 103100, 103080, 103080, 103070, 
    103040, 103000, 102990, 102960, 102920, 102860, 102810, 102730, 102660, 
    102590, 102540, 102440, 102340, 102230, 102160, 102080, 102030, 101930, 
    101820, 101780, 101740, 101730, 101650, 101620, 101590, 101540, 101510, 
    101500, 101510, 101530, 101510, 101530, 101540, 101540, 101570, 101570, 
    101610, 101600, 101620, 101690, 101730, 101740, 101780, 101780, 101840, 
    101850, 101910, 101970, 101990, 102020, 102070, 102100, 102140, 102160, 
    102200, 102210, 102240, 102270, 102310, 102360, 102400, 102430, 102450, 
    102470, 102490, 102500, 102500, 102520, 102540, 102580, 102620, 102640, 
    102650, 102680, 102700, 102720, 102720, 102730, 102720, 102730, 102730, 
    102740, 102760, 102780, 102780, 102790, 102800, 102780, 102780, 102770, 
    102780, 102760, 102750, 102760, 102770, 102780, 102790, 102780, 102790, 
    102780, 102790, 102780, 102750, 102750, 102780, 102740, 102740, 102740, 
    102750, 102760, 102750, 102750, 102740, 102730, 102730, 102740, 102750, 
    102770, 102790, 102800, 102810, 102810, 102820, 102820, 102800, 102790, 
    102800, 102790, 102770, 102750, 102750, _, 102730, 102740, 102740, 
    102690, 102670, 102640, 102620, 102600, 102580, 102570, 102580, 102580, 
    102580, 102550, 102510, 102500, 102490, 102450, 102450, 102440, 102410, 
    102420, 102370, 102360, 102380, 102350, 102320, 102290, 102270, 102270, 
    102260, 102230, 102190, 102180, 102170, 102190, 102230, 102220, 102210, 
    102200, 102110, 102080, 102070, 102060, 102040, 102060, 102020, 102010, 
    101990, 101950, 101930, 101900, 101880, 101860, 101850, 101870, 101870, 
    101930, 101960, _, 102030, 101940, 101960, 101980, 101990, 101990, 
    101990, 102070, 102050, 101990, 102010, 102070, 102100, 102080, 102080, 
    102070, 102070, 102070, 102070, 102090, 102100, 102100, 102120, 102090, 
    102120, 102120, 102130, 102130, 102130, 102120, 102110, 102100, 102060, 
    102050, 102030, 102010, 102000, 102010, 102010, 102000, 101990, 101980, 
    101990, 101990, 101980, 101990, 102000, 102020, 102020, 102050, 102040, 
    102040, 102060, 102040, 102050, 102040, 102030, 102040, 102040, 102040, 
    102050, 102060, 102060, 102070, 102070, 102070, 102070, 102070, 102090, 
    102090, 102080, 102070, 102090, 102100, 102110, 102080, 102030, 102030, 
    102020, 101980, 101920, 101920, 101910, 101860, 101820, 101790, 101720, 
    101700, 101670, 101640, 101590, 101530, 101540, 101540, 101560, 101580, 
    101600, 101610, 101680, 101700, 101730, 101780, 101840, 101860, 101890, 
    101890, 101890, 101920, 101950, 101980, 102000, 102000, 102020, 102050, 
    102070, 102050, 102040, 102060, 102080, 102080, 102060, 102070, 102050, 
    102060, 102040, 102020, 102000, 102000, 101970, 101970, 101930, 101930, 
    101880, 101850, 101820, 101820, 101770, 101750, 101710, 101660, 101630, 
    101580, 101550, 101520, 101510, 101480, 101430, 101420, 101350, 101290, 
    101240, 101190, 101120, 101040, 100950, 100870, 100840, 100750, 100640, 
    100510, 100480, 100440, 100430, 100440, 100430, 100430, 100390, 100400, 
    100430, 100470, 100470, 100460, 100460, 100430, 100450, 100420, 100430, 
    100440, 100430, 100470, 100480, 100460, 100410, 100390, 100400, 100350, 
    100300, 100270, 100250, 100210, 100110, 100080, 100150, 100070, 100030, 
    99980, 100030, 100020, 100050, 100100, 100100, 100080, 100070, 100090, 
    100100, 100110, 100110, 100110, 100120, 100120, 100130, 100150, 100170, 
    100190, 100220, 100230, 100250, 100270, 100250, 100250, 100250, 100260, 
    100250, 100260, 100240, 100230, 100230, 100200, 100190, 100170, 100160, 
    100140, 100100, 100070, 100050, 100010, 99990, 99980, 99960, 99950, 
    99940, 99910, 99880, 99860, 99830, 99810, 99790, 99770, 99740, 99730, 
    99700, 99690, 99670, 99660, 99650, 99640, 99630, 99620, 99640, 99620, 
    99630, 99640, 99660, 99690, 99720, 99740, 99750, 99780, 99800, 99820, 
    99860, 99860, 99900, 99930, 99960, 100000, 100050, 100080, 100100, 
    100120, 100150, 100160, 100180, 100220, 100230, 100270, 100300, 100320, 
    100340, 100360, 100350, 100360, 100380, 100410, 100440, 100470, 100460, 
    100460, 100460, 100450, 100520, 100590, 100620, 100680, 100770, 100820, 
    100910, 101010, 101030, 101110, 101190, 101250, 101310, 101380, 101420, 
    101450, 101480, 101500, 101540, 101530, 101540, 101560, 101570, 101590, 
    101620, 101650, 101690, 101730, 101750, 101780, 101790, 101820, 101850, 
    101880, 101920, 101930, 101970, 102000, 102010, 102010, 102020, 102020, 
    102010, 102000, 102000, 101980, 101990, 101980, 101970, 101980, 101950, 
    101930, 101900, 101860, 101830, 101810, 101800, 101790, 101790, 101790, 
    101790, 101780, 101780, 101810, 101780, 101770, 101750, 101750, 101730, 
    101770, 101790, 101760, 101730, 101680, 101630, 101620, 101640, 101640, 
    101590, 101690, 101700, 101700, 101680, 101650, 101610, 101510, 101450, 
    101360, 101430, 101380, 101370, 101420, 101480, 101440, 101450, 101490, 
    101540, 101510, 101510, 101480, 101510, 101560, 101530, 101530, 101530, 
    101480, 101490, 101470, 101460, 101470, 101450, 101460, 101470, 101470, 
    101500, 101490, 101520, 101530, 101540, 101510, 101510, 101520, 101510, 
    101540, 101550, 101580, 101570, 101580, 101600, 101630, 101640, 101650, 
    101660, 101670, 101690, 101710, 101700, 101720, 101710, 101690, 101700, 
    101680, 101680, 101700, 101690, 101680, 101650, 101650, 101650, 101660, 
    101590, 101620, 101590, 101550, 101500, 101460, 101410, 101320, 101280, 
    101180, 101120, 101010, 100900, 100830, 100730, 100650, 100620, 100580, 
    100610, 100530, 100490, 100440, 100410, 100350, 100340, 100280, 100260, 
    100250, 100300, 100340, 100370, 100420, 100470, 100530, 100590, 100670, 
    100760, 100880, 101000, 101080, 101200, 101330, 101490, 101660, 101840, 
    101970, 102100, 102230, 102330, 102430, 102540, 102650, 102750, 102820, 
    102880, 102980, 103020, 103070, 103140, 103190, 103200, 103220, 103250, 
    103260, 103260, 103270, 103280, 103290, 103260, 103260, 103240, 103210, 
    103190, 103150, 103120, 103100, 103080, 103070, 103070, 103030, 103020, 
    103000, 102950, 102900, 102850, 102800, 102760, 102710, 102670, 102620, 
    102570, 102520, 102500, 102440, 102370, 102310, 102250, 102210, 102140, 
    102080, 102010, 101960, 101910, 101870, 101830, 101780, 101730, 101670, 
    101610, 101590, 101540, 101480, 101470, 101440, 101430, 101380, 101360, 
    101340, 101330, 101310, 101320, 101400, 101450, 101540, 101590, 101650, 
    101770, 101840, 101900, 101960, 101960, 101990, 102020, 102020, 102010, 
    101990, 101990, 101980, 101970, 101940, 101920, 101890, 101820, 101750, 
    101670, 101620, 101560, 101500, 101430, 101380, 101310, 101260, 101210, 
    101160, 101120, 101090, 101010, 100970, 100930, 100880, 100820, 100760, 
    100690, 100690, 100720, 100690, 100720, 100720, 100700, 100700, 100750, 
    100770, 100810, 100830, 100840, 100860, 100860, 100880, 100880, 100890, 
    100860, 100840, 100880, 100850, 100860, 100880, 100910, 100920, 100930, 
    100910, 100940, 100920, 100930, 100920, 100870, 100830, 100880, 100980, 
    101020, 101060, 101150, 101210, 101250, 101280, 101330, 101320, 101370, 
    101420, 101520, 101590, 101600, 101610, 101670, 101700, 101710, 101730, 
    101750, 101780, 101800, 101790, 101810, 101870, 101890, 101910, 101940, 
    101950, 101940, 101940, 101920, 101940, 101930, 101900, 101920, 101880, 
    101870, 101850, 101850, 101820, 101800, 101790, 101760, 101710, 101690, 
    101680, 101630, 101610, 101580, 101540, 101490, 101430, 101380, 101360, 
    101300, 101230, 101190, 101150, 101110, 101090, 101030, 100990, 100950, 
    100910, 100880, 100850, 100920, 100810, 100820, 100820, 100830, 100820, 
    100830, 100830, 100860, 100860, 100830, 100820, 100810, 100850, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 101050, 101050, 101030, 101040, 
    101050, 101070, 101120, 101120, 101140, 101130, 101110, 101090, 101050, 
    100990, 100960, 100920, 100890, 100840, 100800, 100750, 100710, 100700, 
    100680, 100650, 100670, 100680, 100690, 100690, 100680, 100680, 100670, 
    100670, 100680, 100710, 100700, 100690, 100690, 100710, 100700, 100690, 
    100690, _, _, _, _, 100630, _, 100550, _, 100430, 100380, 100310, 100280, 
    _, 100190, _, 100040, 99960, _, 99960, _, _, 100050, _, _, 100080, _, 
    100110, 100140, 100200, 100270, 100300, _, 100370, 100440, 100480, 
    100520, 100520, _, _, 100590, _, 100640, 100660, 100670, 100710, 100720, 
    100730, _, _, 100770, 100780, _, 100800, 100850, _, 100880, 100880, 
    100900, 100900, _, _, _, _, 100970, _, 101020, _, 101060, 101060, _, _, 
    101130, _, 101170, _, 101200, _, 101290, 101320, _, 101380, 101410, 
    101450, 101460, _, 101540, 101560, 101600, 101650, _, 101730, 101780, _, 
    101830, _, 101880, 101890, 101940, 101960, 101980, 102010, 102050, 
    102080, 102110, 102120, 102120, 102150, 102150, _, 102170, 102170, 
    102160, 102130, 102110, _, 102060, _, _, 101980, 101890, 101840, 101750, 
    101660, 101590, _, 101370, _, 101330, 101260, _, 101020, _, 100890, 
    100800, 100770, 100760, _, 100900, 100710, _, 100840, _, 100870, 100890, 
    100910, _, _, 100930, _, 100970, 101010, _, 101000, 101000, 101000, 
    101000, _, 100990, 100990, 101040, 101120, _, 101160, 101160, 101200, 
    101240, 101220, 101210, 101180, 101170, 101100, 101070, 101060, 101050, 
    101040, 101040, 101040, 101050, 101060, 101060, 101080, 101100, 101110, 
    101140, 101160, 101160, 101150, 101200, _, 101190, 101200, 101180, 
    101200, _, 101190, 101170, 101170, 101160, _, 101150, 101120, 101070, 
    101020, _, 100910, 100850, _, 100650, _, 100510, 100460, 100380, 100280, 
    _, 100170, 100120, 100070, 100010, _, 99970, 99970, 99970, 99980, _, 
    100010, 100000, 100000, 100000, _, 100020, 100040, 100040, 100030, _, _, 
    100020, 100010, 99980, 99950, 99920, _, 99900, 99900, 99900, 99900, 
    99900, 99920, 99960, 99990, 100000, 100040, _, _, 100150, 100130, _, 
    100160, 100190, 100180, 100200, _, 100200, 100250, 100220, 100240, _, 
    100270, 100310, 100320, 100390, _, 100490, 100550, 100580, 100630, _, 
    100690, 100680, 100730, 100710, _, 100690, 100710, 100760, 100780, _, 
    100790, 100790, 100790, 100790, 100790, 100760, 100770, _, 100800, _, 
    100820, 100820, 100830, 100790, _, 100800, 100780, 100760, 100750, 
    100730, 100710, _, 100680, 100640, 100610, 100590, 100530, 100520, 
    100490, 100470, 100470, 100450, 100450, 100460, 100440, 100430, _, 
    100390, 100350, 100320, 100320, 100350, 100370, 100410, 100440, 100510, 
    100520, 100550, 100540, 100570, 100600, 100620, 100610, 100600, 100610, 
    100590, 100620, 100660, 100680, 100680, 100680, 100700, 100740, 100750, 
    100750, 100780, 100800, 100840, 100860, 100890, 100930, 100970, 101010, 
    101050, 101090, 101130, 101170, 101210, 101240, 101300, 101350, 101380, 
    101420, 101470, 101490, 101510, 101530, 101540, 101560, 101580, 101610, 
    101630, 101660, 101650, 101660, 101660, 101660, 101680, 101660, 101670, 
    101670, 101660, 101670, 101670, 101680, 101650, 101610, 101620, 101580, 
    101540, 101480, 101460, 101440, 101370, 101320, 101250, 101220, 101180, 
    101140, 101070, 101030, 100990, 100940, 100900, 100840, 100810, 100780, 
    100750, 100730, 100730, 100730, 100730, 100750, 100720, 100760, 100750, 
    100760, 100780, 100830, 100870, 100870, 100880, 100910, 100930, 100920, 
    100940, 100930, 100950, 100940, 100960, 101020, 101030, 101060, 101110, 
    101130, 101160, 101200, 101230, 101250, 101260, 101300, 101290, 101330, 
    101350, 101370, 101370, 101400, 101400, 101420, 101420, 101430, 101440, 
    101460, 101470, 101480, 101500, 101520, 101510, 101550, 101560, 101570, 
    101580, 101600, 101620, 101630, 101630, 101660, 101670, 101690, 101690, 
    101700, 101690, 101690, 101720, 101690, 101680, 101670, 101660, 101650, 
    101660, 101650, 101620, 101620, 101610, 101610, 101590, 101570, 101540, 
    101530, 101510, 101490, 101480, 101470, 101460, 101440, 101420, 101400, 
    101380, 101340, 101320, 101310, 101300, 101300, 101340, 101310, 101300, 
    101310, 101330, 101350, 101340, 101350, 101370, 101370, 101380, 101390, 
    101400, 101440, 101430, 101420, 101410, 101420, 101420, 101410, 101400, 
    101390, 101400, 101410, 101420, 101430, 101430, 101440, 101430, 101430, 
    101410, 101400, 101380, 101360, 101350, 101330, 101320, 101270, 101240, 
    101230, 101200, 101160, 101110, 101030, 100990, 100880, 100950, 100890, 
    100860, 100800, 100790, 100760, _, 100750, _, _, _, _, _, _, _, _, _, _, 
    99760, _, _, _, _, _, _, _, _, _, 99050, 99090, 99210, 99310, 99370, 
    99500, 99560, 99670, 99750, 99850, 99940, 100020, 100150, 100250, 100370, 
    100440, 100510, 100580, 100640, 100680, 100730, 100780, 100850, 100920, 
    100970, 101030, 101070, 101130, 101180, 101220, 101240, 101300, 101350, 
    101420, 101470, 101530, 101620, 101640, 101710, 101750, 101770, 101790, 
    101860, 101890, 101890, 101910, 101960, 102000, 102050, 102050, 102100, 
    102120, 102120, 102110, 102110, 102140, 102160, 102170, 102180, 102180, 
    102190, 102220, 102220, 102230, 102220, 102220, 102200, 102190, 102180, 
    102200, 102210, 102210, 102230, 102250, 102250, 102240, 102230, 102210, 
    102200, 102170, 102200, 102200, 102210, 102210, 102230, 102230, 102220, 
    102220, 102250, 102250, 102260, 102250, 102290, 102310, 102330, 102360, 
    102390, 102430, 102430, 102450, 102450, 102450, 102460, 102480, 102500, 
    102490, 102510, 102520, 102510, 102500, 102500, 102490, 102490, 102460, 
    102450, 102440, 102390, 102390, 102400, 102360, 102310, 102280, 102270, 
    102280, 102260, 102250, 102190, 102150, 102130, 102110, 102140, 102120, 
    102050, 102040, 102060, 102070, 102060, 102000, 101990, 101970, 101970, 
    101970, 101980, 102000, 102000, 101940, 101990, 101990, 101980, 101970, 
    101950, 101950, 101930, 101900, 101900, 101890, 101900, 101850, 101880, 
    101900, 101880, 101860, 101860, 101820, 101830, 101810, 101690, 101730, 
    101810, 101700, 101660, 101630, 101670, 101690, 101690, 101670, 101620, 
    101600, 101570, 101630, 101610, 101610, 101580, 101570, 101650, 101680, 
    101640, 101590, 101650, 101610, 101660, 101680, 101600, 101530, 101590, 
    101610, 101610, 101630, 101630, 101590, 101480, 101570, 101460, 101440, 
    101430, 101390, 101340, 101290, 101250, 101360, 101320, 101300, 101300, 
    101340, 101360, 101330, 101370, 101350, 101370, 101350, 101330, 101320, 
    101310, 101290, 101290, 101260, 101270, 101230, 101210, 101220, 101180, 
    101140, 101120, 101110, 101100, 101070, 101070, 101050, 101040, 101040, 
    101020, 101000, 100980, 100980, 100970, 100980, 100940, 100930, 100940, 
    100910, 100910, 100920, 100940, 100930, 100900, 100900, 100890, 100910, 
    100920, 100880, 100880, 100900, 100920, 100870, 100870, 100870, 100880, 
    100890, 100860, 100860, 100890, 100860, 100840, 100800, 100780, 100750, 
    100740, 100740, 100720, 100750, 100740, 100720, 100670, 100670, 100610, 
    100590, 100590, 100570, 100550, 100530, 100540, 100530, 100520, 100510, 
    100500, 100520, 100530, 100530, 100560, 100570, 100600, 100620, 100670, 
    100700, 100730, 100740, 100760, 100850, 100900, 100920, 100920, 100990, 
    101050, 101080, 101140, 101170, 101170, 101190, 101180, 101190, 101230, 
    101240, 101250, 101250, 101270, 101270, 101250, 101270, 101270, 101260, 
    101230, 101190, 101160, 101150, 101150, 101130, 101160, 101160, 101140, 
    101130, 101110, 101010, 100970, 100930, 100930, 100840, 100810, 100850, 
    100850, 100730, 100640, 100550, 100480, 100410, 100290, 100230, 100190, 
    100120, 100090, 100130, 100160, 100210, 100340, 100290, 100310, 100280, 
    100290, 100240, 100210, 100220, 100200, 100170, 100130, 100100, 100100, 
    100080, 100060, 100040, 100040, 100010, 99960, 99960, 99950, 99960, 
    99960, 100000, 100020, 99980, 99990, 99970, 99950, 99900, 99880, 99840, 
    99830, 99840, 99910, 99910, 99930, 99950, 99980, 100030, 100050, 100070, 
    100100, 100160, 100190, 100220, 100260, 100300, 100370, 100410, 100460, 
    100500, 100520, 100540, 100600, 100670, 100740, 100780, 100800, 100850, 
    100920, 100980, 101030, 101040, 101070, 101100, 101160, 101240, 101300, 
    101370, 101430, 101440, 101470, 101480, 101500, 101530, 101540, 101520, 
    101560, 101560, 101570, 101570, 101570, 101580, 101590, 101590, 101590, 
    101600, 101590, 101570, 101590, 101600, 101620, 101640, 101660, 101650, 
    101660, 101690, 101710, 101710, 101720, 101710, 101710, 101720, 101710, 
    101710, 101690, 101690, 101670, 101640, 101610, 101610, 101580, 101560, 
    101540, 101530, 101510, 101490, 101480, 101450, 101400, 101430, 101350, 
    101330, 101280, 101250, 101240, 101220, 101200, 101200, 101200, 101180, 
    101150, 101140, 101140, 101160, 101170, 101170, 101200, 101200, 101220, 
    101260, 101290, 101310, 101350, 101380, 101420, 101480, 101510, 101530, 
    101540, 101570, 101590, 101610, 101650, 101640, 101590, 101610, 101660, 
    101690, 101720, 101750, 101770, 101810, 101830, 101880, 101930, 101990, 
    102030, 102060, 102090, 102130, 102140, 102170, 102190, 102180, 102200, 
    102220, 102260, 102270, 102270, 102260, 102250, 102270, 102250, 102250, 
    102250, 102250, 102240, 102260, 102250, 102250, 102250, 102240, 102220, 
    102200, 102210, 102200, 102180, 102160, 102130, 102130, 102150, 102110, 
    102070, 102080, 102060, 102050, 102050, 102010, 101990, 101960, 101950, 
    101950, 101950, 101940, 101920, 101880, 101870, 101840, 101840, 101810, 
    101770, 101730, 101720, 101700, 101670, 101630, 101600, 101570, 101550, 
    101530, 101490, 101460, 101410, 101380, 101380, 101350, 101330, 101310, 
    101270, 101250, 101220, 101190, 101170, 101140, 101120, 101100, 101080, 
    101060, 101060, 101040, 101020, 101000, 100980, 100950, 100930, 100910, 
    100890, 100870, 100870, 100890, 100920, 100920, 100900, 100880, 100880, 
    100860, 100840, 100770, 100720, 100700, 100680, 100660, 100640, 100620, 
    100600, 100610, 100600, 100600, 100610, 100610, 100600, 100610, 100620, 
    100670, 100710, 100740, 100750, 100780, 100780, 100800, 100820, 100830, 
    100850, 100860, 100870, 100880, 100880, 100900, 100910, 100900, 100880, 
    100870, 100860, 100850, 100830, 100820, 100810, 100810, 100800, 100810, 
    100830, 100830, 100850, 100880, 100910, 100940, 100990, 101020, 101020, 
    101050, 101090, 101100, 101110, 101140, 101150, 101150, 101150, 101140, 
    101150, 101150, 101140, 101170, 101190, 101220, 101210, 101190, 101190, 
    101200, 101190, 101160, 101140, 101100, 101080, 101040, 101010, 100980, 
    100960, 100940, 100920, 100910, 100900, 100890, 100850, 100820, 100820, 
    100820, 100830, 100830, 100850, 100840, 100830, 100800, 100790, 100770, 
    100750, 100750, 100730, 100730, 100740, 100720, 100720, 100690, 100670, 
    100670, 100670, 100640, 100610, 100600, 100600, 100610, 100620, 100640, 
    100650, 100650, 100660, 100640, 100630, 100600, 100580, 100560, 100560, 
    100540, 100540, 100510, 100500, 100510, 100510, 100520, 100480, 100440, 
    100410, 100400, 100420, 100420, 100420, 100440, 100430, 100430, 100420, 
    100410, 100390, 100370, 100330, 100320, 100310, 100310, 100310, 100300, 
    100300, 100280, 100270, 100240, 100230, 100220, 100220, 100230, 100240, 
    100270, 100280, 100280, 100290, 100290, 100290, 100300, 100310, 100320, 
    100330, 100330, 100340, 100350, 100350, 100370, 100370, 100390, 100370, 
    100360, 100340, 100330, 100280, 100280, 100270, 100260, 100230, 100210, 
    100150, 100060, 100070, 100050, 100030, 100010, 99990, 99970, 99960, 
    99990, 99990, 99970, 99960, 99940, 99940, 99930, 99910, 99910, 99900, 
    99920, 99930, 99940, 99960, 99960, 99980, 99990, 100010, 100020, 100040, 
    100060, 100100, 100140, 100170, 100200, 100230, 100260, 100260, 100260, 
    100270, 100280, 100280, 100280, 100280, 100300, 100280, 100300, 100340, 
    100350, 100350, 100350, 100360, 100340, 100350, 100350, 100340, 100340, 
    100280, 100270, 100280, 100260, 100200, 100180, 100200, 100160, 100120, 
    100110, 100090, 100060, 100060, 100060, 100060, 100040, 100030, 100010, 
    100010, 100000, 100000, 100010, 100000, 100010, 100040, 100050, 100040, 
    100040, 100070, 100080, 100110, 100110, 100140, 100150, 100190, 100210, 
    100230, 100260, 100290, 100320, 100370, 100390, 100410, 100430, 100450, 
    100460, 100490, 100530, 100550, 100570, 100570, 100590, 100610, 100630, 
    100640, 100660, 100660, 100670, 100690, 100690, 100690, 100690, 100680, 
    100680, 100660, 100660, 100650, 100640, 100630, 100620, 100610, 100600, 
    100590, 100590, 100580, 100570, 100590, 100590, 100590, 100590, 100570, 
    100570, 100560, 100590, 100600, 100620, 100610, 100620, 100640, 100660, 
    100670, 100680, 100690, 100690, 100690, 100680, 100680, 100700, 100700, 
    100720, 100710, 100690, 100650, 100620, 100570, 100550, 100530, 100520, 
    100500, 100470, 100430, 100390, 100360, 100320, 100260, 100230, 100200, 
    100170, 100190, 100210, 100270, 100360, 100480, 100590, 100640, 100690, 
    100700, 100760, 100800, 100860, 100900, 100940, 100990, 101020, 101070, 
    101110, 101170, 101200, 101230, 101240, 101270, 101300, 101300, 101300, 
    101300, 101290, 101260, 101240, 101240, 101230, 101210, 101200, 101230, 
    101220, 101230, 101250, 101280, 101320, 101330, 101350, 101400, 101420, 
    101430, 101440, 101460, 101480, 101480, 101480, 101450, 101440, 101470, 
    101480, 101460, 101450, 101410, 101360, 101340, 101300, 101280, 101230, 
    101180, 101120, 101060, 100980, 100910, 100790, 100710, 100630, 100510, 
    100380, 100280, 100210, 100170, 100160, 100150, 100210, 100260, 100320, 
    100390, 100450, 100530, 100620, 100720, 100790, 100880, 100930, 101030, 
    101100, 101180, 101180, 101190, 101100, 101110, 101030, 101010, 100990, 
    100860, 100810, 100750, 100710, 100640, 100600, 100620, 100570, 100570, 
    100590, 100620, 100730, 100820, 100860, 100900, 100960, 101040, 101110, 
    101100, 101070, 101030, 100990, 100970, 100960, 100950, 100930, 100910, 
    100900, 100850, 100810, 100800, 100750, 100730, 100720, 100710, 100720, 
    100690, 100680, 100640, 100650, 100630, 100580, 100500, 100420, 100360, 
    100370, 100290, 100210, 100150, 100100, 100020, 99950, 99890, 99830, 
    99760, 99710, 99630, 99600, 99610, 99630, 99630, 99690, 99700, 99730, 
    99750, 99760, 99760, 99760, 99780, 99810, 99820, 99850, 99880, 99850, 
    99920, 99980, 100040, 100080, 100160, 100200, 100240, 100290, 100370, 
    100420, 100450, 100480, 100510, 100530, 100490, 100460, 100400, 100360, 
    100270, 100220, 100140, 100100, 100020, 100040, 99980, 100110, 100290, 
    100410, 100470, 100540, 100610, 100660, 100690, 100690, 100760, 100780, 
    100840, 100940, 100970, 100970, 100990, 101070, 101110, 101130, 101160, 
    101180, 101220, 101240, 101240, 101250, 101300, 101330, 101310, 101290, 
    101320, 101320, 101300, 101290, 101260, 101210, 101110, 101040, 101000, 
    100960, 100910, 100790, 100700, 100620, 100580, 100540, 100500, 100470, 
    100420, 100400, 100360, 100310, 100280, 100210, 100180, 100130, 100070, 
    100020, 100030, 100000, 99990, 99970, 99960, 99970, 99950, 99930, 99910, 
    99890, 99860, 99870, 99880, 99860, 99850, 99810, 99780, 99780, 99750, 
    99750, 99740, 99730, 99810, 99900, 100020, 100090, 100160, 100250, 
    100300, 100340, 100400, 100420, 100420, 100430, 100430, 100440, 100410, 
    100410, 100370, 100330, 100300, 100240, 100150, 100080, 99990, 99960, 
    99890, 99830, 99790, 99730, 99660, 99600, 99520, 99520, 99480, 99460, 
    99370, 99280, 99180, 99080, 99040, 98950, 98840, 98750, 98710, 98710, 
    98680, 98640, 98640, 98580, 98530, 98510, 98450, 98400, 98350, 98310, 
    98290, 98260, 98170, 98140, 98050, 98010, 97950, 97890, 97840, 97770, 
    97720, 97670, 97620, 97580, 97530, 97490, 97460, 97440, 97450, 97430, 
    97430, 97470, 97520, 97590, 97650, 97700, 97750, 97800, 97850, 97940, 
    98000, 98090, 98170, 98290, 98390, 98490, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 99340, 99340, 99360, 99370, 99370, 99380, _, 99390, 
    99360, 99360, 99350, 99320, 99300, 99300, 99300, 99280, 99270, 99270, 
    99250, 99220, 99180, 99140, 99110, 99080, 99090, 99070, 99050, 99060, 
    99060, 99070, 99100, 99110, 99120, 99100, 99090, 99080, 99080, 99100, 
    99090, 99080, 99050, 99000, 98950, 98900, 98790, 98790, 98750, 98740, 
    98760, 98770, 98780, 98800, 98810, 98800, 98780, 98720, 98640, 98590, 
    98540, 98470, 98450, 98460, 98500, 98540, 98610, 98720, 98840, 98980, 
    99080, 99170, 99280, 99420, 99560, 99680, 99770, 99860, 99950, 100020, 
    100080, 100120, 100170, 100210, 100280, 100320, 100380, 100450, 100510, 
    100570, 100630, 100690, 100750, 100800, 100860, 100890, 100950, 100980, 
    101000, 101030, 101060, 101080, 101090, 101080, 101070, 101060, 101080, 
    101070, 101070, 101050, 101050, 101070, 101030, 101010, 100990, 100980, 
    100970, 100960, 100960, 100960, 100910, 100880, 100880, 100860, 100850, 
    100870, 100870, 100870, 100890, 100930, 100960, 100990, 101030, 101060, 
    101090, 101120, 101140, 101180, 101210, 101240, 101260, 101270, 101310, 
    101340, 101360, 101390, 101390, 101400, 101380, 101380, 101370, 101360, 
    101350, 101340, 101320, 101310, 101300, 101260, 101240, 101210, 101180, 
    101170, 101120, 101100, 101080, 101040, 101020, 101000, 100970, 100930, 
    100890, 100870, 100840, 100830, 100780, 100760, 100710, 100680, 100650, 
    100620, 100590, 100560, 100530, 100510, 100490, 100460, 100440, 100440, 
    100460, 100490, 100530, 100560, 100590, 100650, 100690, 100740, 100770, 
    100810, 100870, 100920, 101000, 101060, 101120, 101140, 101190, 101230, 
    101300, 101330, 101340, 101390, 101440, 101490, 101530, 101550, 101610, 
    101620, 101650, 101660, 101660, 101680, 101680, 101700, 101690, 101740, 
    101750, 101750, 101760, 101790, 101790, 101810, 101820, 101820, 101810, 
    101840, 101840, 101810, 101880, 101890, 101920, 101940, 101940, 101930, 
    101920, 101910, 101930, 101960, 101930, 101940, 101990, 101980, 102000, 
    102050, 102000, 102000, 102010, 101980, 101960, 101960, 101960, 101940, 
    101940, 101940, 101910, 101900, 101910, 101860, 101840, 101850, 101850, 
    101780, 101750, 101770, 101780, 101770, 101720, 101710, 101690, 101670, 
    101650, 101620, 101620, 101610, 101620, 101590, 101600, 101630, 101620, 
    101620, 101590, 101600, 101600, 101580, 101560, 101560, 101570, 101580, 
    101560, 101550, 101560, 101540, 101500, 101480, 101400, 101380, 101330, 
    101370, 101400, 101400, 101400, 101390, 101390, 101380, 101360, 101350, 
    101400, 101410, 101420, 101370, 101420, 101430, 101420, 101420, 101420, 
    101470, 101410, 101410, 101510, 101520, 101440, 101480, 101460, 101450, 
    101470, 101430, 101420, 101370, 101350, 101250, 101190, 101120, 101080, 
    101030, 100880, 100820, 100770, 100650, 100490, 100420, 100340, 100230, 
    100110, 99990, 99930, 99830, 99700, 99580, 99520, 99500, 99430, 99300, 
    99350, 99290, 99220, 99150, 99180, 99130, 99090, 99140, 99160, 99170, 
    99230, 99270, 99360, 99460, 99570, 99660, 99760, 99860, 99970, 100070, 
    100200, 100330, 100440, 100480, 100600, 100710, 100780, 100880, 100960, 
    101040, 101130, 101200, 101310, 101370, 101420, 101500, 101570, 101640, 
    101700, 101720, 101760, 101830, 101890, 101890, 101940, 101940, 101940, 
    101950, 101950, 101980, 101950, 101930, 101900, 101860, 101850, 101830, 
    101780, 101730, 101690, 101650, 101600, 101560, 101540, 101470, 101410, 
    101380, 101320, 101250, 101210, 101170, 101160, 101130, 101130, 101100, 
    101080, 101050, 101020, 100990, 100870, 100870, 100870, 100800, 100750, 
    100770, 100690, 100640, 100620, 100620, 100570, 100590, 100570, 100570, 
    100580, 100520, 100500, 100440, 100340, 100210, 100130, 100010, 99750, 
    99620, 99490, 99500, 99250, 99130, 99070, 98940, 98960, 99040, 99100, 
    99230, 99350, 99530, 99690, 99850, 100080, 100210, 100250, 100360, 
    100350, 100390, 100460, 100490, 100550, 100550, 100610, 100670, 100760, 
    100840, 100920, 100980, 101030, 101120, 101160, 101240, 101260, 101390, 
    101390, 101470, 101490, 101540, 101550, 101560, 101550, 101550, 101570, 
    101580, 101580, 101620, 101640, 101660, 101670, 101670, 101690, 101640, 
    101630, 101590, 101540, 101500, 101410, 101350, 101240, 101060, 100820, 
    100620, 100560, 100520, 100490, 100460, 100480, 100520, 100580, 100620, 
    100700, 100760, 100800, 100910, 100990, 101070, 101070, 101010, 100990, 
    101060, 101000, 100960, 100910, 100910, 100910, 100870, 100900, 100980, 
    101040, 101130, 101210, 101280, 101330, 101420, 101500, 101590, 101670, 
    101740, 101760, 101780, 101780, 101770, 101820, 101820, 101840, 101840, 
    101810, 101800, 101790, 101750, 101730, 101720, 101690, 101670, 101670, 
    101690, 101700, 101720, 101750, 101770, 101810, 101800, 101860, 101870, 
    101930, 101950, 101980, 102000, 101990, 102000, 101980, 101970, 101940, 
    101920, 101890, 101830, 101740, 101690, 101670, 101640, 101600, 101590, 
    101600, 101570, 101580, 101580, 101590, 101570, 101600, 101600, 101600, 
    101620, 101630, 101650, 101670, 101680, 101680, 101710, 101710, 101690, 
    101690, 101700, 101710, 101730, 101740, 101720, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 100820, 100720, 100700, 100640, 100650, 100620, 100620, 
    100610, 100600, 100570, 100520, 100500, 100450, 100410, 100400, 100360, 
    100330, 100290, 100260, 100210, 100200, 100170, 100170, 100170, 100210, 
    100200, 100180, 100170, 100170, 100170, 100160, 100170, 100180, 100190, 
    100220, 100240, 100260, 100250, 100300, 100300, 100320, 100350, 100350, 
    100350, 100390, 100490, 100470, 100460, 100440, _, 100390, 100330, 
    100330, 100230, 100180, 100150, 100050, 99940, 99940, 99860, 99800, 
    99750, 99630, 99440, 99310, 99120, 99040, 98980, 98870, 98800, 98780, 
    98800, 98830, 98860, 98880, 98890, 98930, 98940, 98940, 98970, 99010, 
    99050, 99100, 99130, 99150, 99190, 99190, 99190, 99180, 99150, 99190, 
    99150, 99180, 99200, 99230, 99250, 99260, 99290, 99320, 99310, 99300, 
    99300, 99310, 99320, 99320, 99350, 99420, 99450, 99410, 99370, 99390, 
    99410, 99430, 99450, 99460, 99470, 99500, 99520, 99540, 99620, 99630, 
    99670, 99690, 99700, 99700, 99770, 99830, 99890, 99930, 99930, 99960, 
    99990, 99990, 100020, 100030, 100050, 100080, 100170, 100260, 100340, 
    100410, 100500, 100570, 100650, 100720, 100780, 100850, 100900, 100920, 
    100970, 101020, 101110, 101170, 101260, 101340, 101420, 101520, 101570, 
    101670, 101760, 101850, 101950, 102030, 102110, 102170, 102190, 102240, 
    102270, 102280, 102290, 102240, 102170, 102110, 102050, 102010, 101980, 
    101910, 101790, 101720, 101640, 101560, 101470, 101400, 101330, 101250, 
    101220, 101140, 101080, 101030, 100940, 100860, 100750, 100660, 100520, 
    100440, 100380, 100330, 100300, 100290, 100330, 100370, 100420, 100480, 
    100560, 100650, 100750, 100850, 101040, 101260, 101450, 101570, 101690, 
    101820, 101970, 102050, 102170, 102260, 102350, 102440, 102540, 102510, 
    102540, 102520, 102520, 102480, 102390, 102390, 102310, 102200, 102090, 
    101980, 101880, 101730, 101600, 101420, 101260, 101070, 100970, 100800, 
    100680, 100540, 100420, 100390, 100280, 100280, 100310, 100320, 100300, 
    100340, 100390, 100430, 100520, 100610, 100700, 100750, 100860, 100960, 
    100980, 101180, 101210, 101350, 101460, 101540, 101680, 101810, 101950, 
    102050, 102180, 102220, 102290, 102340, 102390, 102380, 102430, 102450, 
    102430, 102420, 102410, 102440, 102450, 102490, 102540, 102550, 102550, 
    102570, 102580, 102600, 102590, 102600, 102560, 102520, 102470, 102390, 
    102320, 102230, 102190, 102140, 102100, 102090, 102020, 101970, 101920, 
    101860, 101810, 101730, 101680, 101620, 101550, 101520, 101440, 101430, 
    101400, 101390, 101340, 101340, 101320, 101280, 101250, 101240, 101220, 
    101240, 101260, 101310, 101340, 101420, 101450, 101470, 101410, 101450, 
    101440, 101410, 101380, 101340, 101310, 101300, 101270, 101190, 101120, 
    101060, 100990, 100930, 100880, 100840, 100810, 100810, 100840, 100850, 
    100880, 100910, 100930, 100970, 101020, 101080, 101120, 101140, 101170, 
    101200, 101220, 101250, 101290, 101330, 101380, 101410, 101440, 101480, 
    101490, 101510, 101550, 101570, 101600, 101630, 101680, 101710, 101730, 
    101740, 101780, 101800, 101840, 101870, 101900, 101930, 101940, 101980, 
    102030, 102070, 102080, 102070, 102090, 102080, 102100, 102110, 102080, 
    102060, 102060, 102060, 102050, 102020, 101990, 101970, 101930, 101930, 
    101840, 101810, 101800, 101710, 101700, 101630, 101570, 101490, 101390, 
    101270, 101120, 101000, 100880, 100730, 100580, 100450, 100360, 100270, 
    100180, 100130, 100060, 100030, 99980, 99980, 99950, 99900, 99860, 99770, 
    99700, 99590, 99530, 99440, 99410, 99380, 99410, 99480, 99550, 99490, 
    99440, 99360, 99320, 99310, 99200, 99230, 99220, 99280, 99360, 99490, 
    99620, 99750, 99850, 100040, 100090, 100250, 100310, 100400, 100530, 
    100670, 100770, 100880, 100900, 100940, 100980, 100980, 101050, 101190, 
    101260, 101270, 101320, 101350, 101380, 101410, 101430, 101420, 101440, 
    101450, 101480, 101510, 101540, 101550, 101590, 101600, 101610, 101630, 
    101630, 101610, 101610, 101590, 101570, 101550, 101500, 101490, 101450, 
    101420, 101400, 101370, 101370, 101350, 101340, 101340, 101350, 101350, 
    101390, 101390, 101400, 101420, 101440, 101440, 101460, 101460, 101440, 
    101440, 101470, 101430, 101430, 101450, 101440, 101400, 101360, 101320, 
    101310, 101320, 101320, 101310, 101290, 101340, 101350, 101350, 101340, 
    101340, 101320, 101310, 101310, 101280, 101250, 101230, 101180, 101170, 
    101140, 101120, 101110, 101090, 101080, 101070, 101040, 101040, 101040, 
    101040, 101080, 101090, 101080, 101150, 101180, 101180, 101180, 101180, 
    101200, 101200, 101190, 101170, 101120, 101100, 101040, 101020, 100910, 
    100860, 100830, 100760, 100660, 100630, 100530, 100490, 100430, 100420, 
    100410, 100420, 100470, 100600, 100640, 100660, 100700, 100770, 100910, 
    100930, 100990, 101100, 101200, 101300, 101370, 101460, 101500, 101540, 
    101550, 101610, 101650, 101700, 101780, 101870, 101960, 102030, 102110, 
    102220, 102340, 102420, 102510, 102600, 102690, 102800, 102880, 102960, 
    103030, 103050, 103090, 103110, 103100, 103130, 103130, 103130, 103090, 
    103100, 103040, 103010, 103060, 103010, 102950, 102940, 102870, 102820, 
    102810, 102750, 102720, 102670, 102640, 102560, 102580, 102590, 102580, 
    102580, 102550, 102560, 102580, 102560, 102540, 102570, 102530, 102520, 
    102540, 102510, 102500, 102460, 102400, 102340, 102330, 102340, 102250, 
    102300, 102210, 102170, 102150, 102090, 102050, 102010, 101950, 101900, 
    101850, 101800, 101780, 101750, 101700, 101680, 101650, 101610, 101570, 
    101530, 101490, 101420, 101390, 101350, 101300, 101260, 101230, 101190, 
    101150, 101120, 101070, 101040, 101030, 100980, 100940, 100930, 100900, 
    100800, 100840, 100900, 100880, 100890, 100970, 101020, 101040, 101100, 
    101110, 101120, 101130, 101170, 101190, 101180, 101180, 101210, 101250, 
    101240, 101270, 101270, 101270, 101310, 101320, 101340, 101360, 101390, 
    101420, 101450, 101440, 101430, 101410, 101410, 101410, 101420, 101440, 
    101460, 101480, 101510, 101550, 101580, 101610, 101600, 101600, 101610, 
    101620, 101650, 101640, 101670, 101660, 101660, 101710, 101740, 101750, 
    101750, 101760, 101800, 101810, 101820, 101830, 101860, 101930, 101960, 
    101960, 101960, 102040, 102070, 102070, 102050, 102140, 102270, 102330, 
    102380, 102430, 102470, 102510, 102640, 102680, 102710, 102780, 102860, 
    102910, 102950, 102980, 103030, 103070, 103100, 103140, 103150, 103200, 
    103230, 103250, 103270, 103290, 103290, 103300, 103310, 103320, 103320, 
    103350, 103380, 103390, 103420, 103420, 103430, 103410, 103430, 103430, 
    103430, 103440, 103440, 103440, 103430, 103440, 103440, 103430, 103400, 
    103390, 103380, 103370, 103340, 103320, 103320, 103320, 103330, 103320, 
    103330, 103330, 103320, 103320, 103340, 103320, 103310, 103320, 103330, 
    103330, 103320, 103300, 103300, 103280, 103280, 103250, 103230, 103190, 
    103170, 103160, 103150, 103140, 103130, 103090, 103070, 103030, 103000, 
    102970, 102930, 102910, 102890, 102860, 102830, 102800, 102770, 102760, 
    102730, 102710, 102690, 102680, 102670, 102670, 102680, 102690, 102680, 
    102690, 102700, 102730, 102750, 102720, 102710, 102730, 102750, 102770, 
    102790, 102790, 102800, 102810, 102830, 102840, 102840, 102830, 102820, 
    102850, 102850, 102860, 102860, 102860, 102870, 102860, 102900, 102900, 
    102900, 102890, 102880, 102860, 102860, 102860, 102850, 102840, 102850, 
    102830, 102800, 102790, 102770, 102740, 102720, 102680, 102650, 102630, 
    102620, 102580, 102540, 102540, 102520, 102480, 102460, 102410, 102370, 
    102300, 102270, 102240, 102200, 102150, 102110, 102070, 102010, 101970, 
    101950, 101920, 101900, 101890, 101900, 101920, 101970, 102010, 102030, 
    102060, 102070, 102080, 102100, 102100, 102100, 102100, 102100, 102110, 
    102110, 102080, 102060, 102050, 102020, 101990, 101950, 101910, 101840, 
    101790, 101740, 101650, 101580, 101490, 101420, 101350, 101270, 101190, 
    101130, 101070, 101010, 100940, 100880, 100830, 100750, 100680, 100620, 
    100570, 100510, 100450, 100390, 100350, 100290, 100220, 100160, 100090, 
    100020, 99920, 99870, 99800, 99700, 99630, 99540, 99450, 99370, 99250, 
    99220, 99080, 98970, 98920, 98810, 98690, 98570, 98510, 98410, 98270, 
    98120, 98030, 97980, 97910, 97900, 97920, 98080, 98230, 98330, 98460, 
    98640, 98600, 98840, 98670, 98810, 98930, 99050, 99160, 99430, 99470, 
    99440, 99580, 99710, 99740, 99670, 99760, 99870, 99910, 99960, 99980, 
    100140, 100240, 100300, 100410, 100440, 100600, 100670, 100760, 100760, 
    100830, 100980, 101040, 101140, 101190, 101250, 101320, 101350, 101390, 
    101470, 101500, 101540, 101550, 101590, 101620, 101690, 101740, 101760, 
    101780, 101810, 101860, 101870, 101900, 101950, 101990, 102020, 102040, 
    102070, 102090, 102120, 102130, 102130, 102130, 102140, 102160, 102140, 
    102140, 102110, 102080, 102070, 102050, 102020, 101990, 101970, 101930, 
    101900, 101860, 101820, 101760, 101720, 101710, 101690, 101680, 101690, 
    101700, 101690, 101610, 101560, 101510, 101460, 101420, 101410, 101370, 
    101360, 101360, 101350, 101310, 101280, 101200, 101180, 101150, 101100, 
    101050, 101000, 100970, 100920, 100880, 100850, 100820, 100770, 100730, 
    100700, 100660, 100620, 100570, 100500, 100440, 100390, 100350, 100320, 
    100300, 100290, 100250, 100160, 100120, 100080, 100050, 100020, 99990, 
    99960, 99940, 99930, 99950, 99930, 99910, 99870, 99830, 99770, 99730, 
    99660, 99560, 99500, 99380, 99330, 99270, 99230, 99080, 98900, 98800, 
    98710, 98560, 98450, 98280, 98120, 97960, 97850, 97730, 97630, 97600, 
    97510, 97430, 97450, 97540, 97630, 97760, 97810, 97900, 97950, 98030, 
    98090, 98140, 98190, 98220, 98310, 98410, 98470, 98560, 98660, 98740, 
    98830, 98900, 98970, 99000, 99010, 99040, 99040, 99020, 98980, 98890, 
    98820, 98740, 98690, 98630, 98590, 98580, 98570, 98610, 98640, 98680, 
    98700, 98730, 98730, 98760, 98760, 98810, 98850, 98870, 98900, 99050, 
    99200, 99320, 99450, 99650, 99780, 99980, 100190, 100350, 100500, 100630, 
    100700, 100860, 101000, 101050, 101110, 101210, 101280, 101310, 101390, 
    101430, 101500, 101550, 101570, 101630, 101670, 101710, 101710, 101760, 
    101800, 101830, 101850, 101850, 101880, 101880, 101870, 101850, 101840, 
    101820, 101830, 101810, 101810, 101810, 101760, 101700, 101670, 101690, 
    101640, 101600, 101570, 101520, 101480, 101430, 101360, 101350, 101280, 
    101240, 101240, 101200, 101180, 101130, 101080, 101040, 101000, 100920, 
    100870, 100860, 100800, 100780, 100720, 100700, 100660, 100610, 100640, 
    100560, 100530, 100530, 100570, 100610, 100610, 100650, 100640, 100630, 
    100610, 100600, 100700, 100730, 100740, 100740, 100750, 100760, 100790, 
    100790, 100790, 100780, 100850, 100870, 100910, 100920, 100950, 100950, 
    101000, 101020, 101050, 101090, 101090, 101120, 101130, 101120, 101130, 
    101160, 101160, 101180, 101170, 101190, 101200, 101220, 101230, 101240, 
    101260, 101290, 101290, 101310, 101310, 101330, 101340, 101380, 101410, 
    101460, 101490, 101530, 101550, 101570, 101580, 101590, 101610, 101640, 
    101680, 101690, 101720, 101720, 101740, 101750, 101760, 101760, 101750, 
    101780, 101770, 101780, 101810, 101850, 101870, 101870, 101880, 101880, 
    101860, 101890, 101900, 101870, 101870, 101870, 101870, 101860, 101870, 
    101840, 101830, 101790, 101750, 101700, 101650, 101620, 101630, 101640, 
    101710, 101760, 101790, 101790, 101790, 101790, 101800, 101790, 101790, 
    101770, 101760, 101740, 101740, 101720, 101710, 101710, 101710, 101690, 
    101680, 101640, 101630, 101570, 101510, 101510, 101470, 101460, 101460, 
    101450, 101440, 101390, 101370, 101330, 101280, 101220, 101240, 101220, 
    101190, 101180, 101190, 101180, 101160, 101120, 101110, 101100, 101080, 
    101060, 101040, 101020, 101010, 100980, 100960, 100980, 100960, 100970, 
    100980, 101000, 101030, 101060, 101110, 101140, 101190, 101230, 101250, 
    101300, 101290, 101270, 101380, 101410, 101510, 101590, 101620, 101680, 
    101710, 101730, 101730, 101760, 101800, 101790, 101760, 101770, 101750, 
    101750, 101730, 101700, 101680, 101670, 101670, 101650, 101620, 101590, 
    101560, 101530, 101510, 101470, 101460, 101450, 101430, 101440, 101430, 
    101410, 101380, 101390, 101370, 101360, 101340, 101310, 101310, 101250, 
    101250, 101260, 101290, 101270, 101260, _, 101250, 101220, 101230, 
    101190, 101220, 101190, 101160, 101160, 101180, 101190, 101190, 101190, 
    101140, 101150, 101170, 101170, 101150, 101160, 101130, 101120, 101070, 
    101050, 101060, 101050, 101090, 101060, 101120, 101130, 101150, 101160, 
    101180, 101200, 101210, 101250, 101220, 101230, 101220, 101220, 101250, 
    101260, 101270, 101300, 101290, 101320, 101350, 101390, 101410, 101390, 
    101420, 101420, 101450, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 101510, 101510, 101470, 101430, 101380, 
    101360, 101280, 101230, 101220, 101200, 101240, 101180, 101130, 101090, 
    101050, 101020, 100970, 100930, 100890, 100860, 100840, 100800, 100770, 
    100740, 100700, 100680, 100680, 100650, 100620, 100590, 100550, 100510, 
    100490, 100470, 100450, 100440, 100450, 100450, 100470, 100490, 100520, 
    100530, 100550, 100560, 100570, 100560, 100550, 100630, 100560, 100550, 
    100570, 100570, 100560, 100480, 100420, 100380, 100310, 100190, 100120, 
    100010, 99830, 99740, 99590, 99420, 99270, 99260, 99300, 99450, 99560, 
    99660, 99760, 99870, 99930, 100020, 100090, 100120, 100120, 100170, 
    100180, 100260, 100290, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 100620, 100590, 100550, 100520, 100470, 100420, 100380, 
    100320, 100300, 100240, 100180, 100120, 100070, 100020, 99970, 99920, 
    99840, 99800, 99800, 99820, 99840, 99870, 99890, 99930, 99980, 100000, 
    100040, 100050, 100080, 100090, 100130, 100120, 100120, 100120, 100090, 
    100040, 100020, 99990, 99960, 99870, 99830, 99760, 99740, 99760, 99770, 
    99780, 99780, _, 99820, 99860, 99920, 99950, 99980, 100060, 100050, 
    100110, 100160, 100160, 100170, 100130, 100120, 100090, 100100, 100050, 
    99970, 100010, 100050, 100060, 100080, 100070, 100050, 100040, 100030, 
    100010, 100000, 100020, 100010, 100010, 99970, 99930, 99900, 99870, 
    99850, 99830, 99800, 99760, 99720, 99720, 99630, 99550, 99610, 99580, 
    99560, 99550, 99510, 99480, 99450, 99430, 99400, 99350, 99350, 99350, 
    99370, 99370, 99410, 99470, 99520, 99560, 99600, 99630, 99650, 99650, 
    99660, 99610, 99520, 99430, 99460, 99410, 99320, 99210, 99110, 99000, 
    98820, 98660, 98400, 98120, 97820, 97460, 97080, 96630, 96350, 96130, 
    95920, 95880, 95900, 96020, 96110, 96280, 96520, 96680, 96910, 97070, 
    97250, 97360, 97520, 97630, 97770, 97850, 97950, 98040, 98080, 98180, 
    98250, 98310, 98350, 98320, 98280, 98230, 98160, 98100, 98050, 97940, 
    97760, 97560, 97270, 96950, 96740, 96700, 96690, 96660, 96720, 96750, 
    96760, 96820, 96840, 96800, 96730, 96740, 96790, 96760, 96740, 96800, 
    96880, 96950, 97000, 97060, 97190, 97290, 97360, 97380, 97340, 97320, 
    97330, 97370, 97350, 97370, 97390, 97400, 97380, 97370, 97350, 97290, 
    97200, 97160, 97100, 97060, 97050, 97010, 97010, 96990, 96980, 97020, 
    97020, 97020, 97050, 97040, 97050, 97060, 97050, 97040, 97040, 97080, 
    97080, 97180, 97230, 97280, 97330, 97370, 97420, 97460, 97480, 97540, 
    97560, 97580, 97560, 97630, 97680, 97690, 97720, 97700, 97730, 97750, 
    97750, 97770, 97770, 97800, 97810, 97820, 97810, 97820, 97850, 97880, 
    97870, 97910, 97960, 97980, 98020, 98050, 98070, 98040, 98030, 98030, 
    98020, 98030, 98030, 98040, 98030, 98020, 98020, 97980, 97960, 97930, 
    97910, 97950, 97920, 97870, 97820, 97870, 97860, 97870, 97910, 97990, 
    97970, 97920, 97950, 98070, 98160, 98240, 98300, 98370, 98460, 98530, 
    98600, 98680, 98810, 98850, 98960, 99070, 99120, 99180, 99360, 99560, 
    99720, 99830, 99940, 100050, 100170, 100270, 100370, 100460, 100550, 
    100620, 100690, 100760, 100800, 100850, 100870, 100910, 100950, 101020, 
    101040, 101070, 101130, 101220, 101270, 101350, 101400, 101410, 101380, 
    101440, 101470, 101470, 101400, 101340, 101320, 101250, 101130, 101040, 
    100970, 100870, 100710, 100510, 100420, 100320, 100180, 100090, 100010, 
    99910, 99920, 99840, 99810, 99750, 99700, 99590, 99620, 99740, 99860, 
    99970, 100010, 100100, 100100, 100170, 100310, 100380, 100460, 100530, 
    100570, 100640, 100690, 100740, 100810, 100870, 100890, 100930, 100940, 
    100960, 100940, 100940, 100990, 101050, 101100, 101080, 101050, 101030, 
    101020, 101050, 101020, 101000, 100990, 100950, 100970, 101000, 101010, 
    101030, 101030, 101040, 101070, 101060, 101110, 101170, 101190, 101240, 
    101310, 101360, 101420, 101510, 101610, 101660, 101700, 101790, 101880, 
    101940, 101990, 102010, 102070, 102130, 102170, 102230, 102230, 102240, 
    102260, 102290, 102300, 102310, 102310, 102330, 102370, 102400, 102430, 
    102450, 102470, 102440, 102470, 102460, 102480, 102490, 102520, 102520, 
    102550, 102500, 102510, 102520, 102530, 102500, 102490, 102420, 102390, 
    102380, 102370, 102380, 102340, 102320, 102260, 102260, 102230, 102180, 
    102140, 102140, 102120, 102120, 102090, 102060, 102050, 102030, 102050, 
    102050, 102040, 102010, 102010, 102000, 102000, 102000, 101960, 101970, 
    101960, 101990, 101970, 101950, 101930, 101920, 101910, 101890, 101870, 
    101850, 101790, 101760, 101740, 101680, 101640, 101550, 101530, 101500, 
    101440, 101410, 101370, 101300, 101270, 101240, 101230, 101230, 101190, 
    101130, 101130, 101080, 101070, 101020, 100950, 100880, 100800, 100720, 
    100670, 100630, 100600, 100560, 100560, 100540, 100520, 100490, 100460, 
    100430, 100370, 100320, 100280, 100200, 100070, 99880, 99810, 99680, 
    99520, 99380, 99160, 99000, 98840, 98810, 98700, 98590, 98470, 98380, 
    98300, 98250, 98220, 98200, 98200, 98240, 98290, 98360, 98390, 98470, 
    98550, 98620, 98690, 98780, 98820, 98860, 98850, 98850, 98810, 98790, 
    98760, 98790, 98740, 98660, 98610, 98650, 98660, 98630, 98580, 98570, 
    98570, 98540, 98560, 98590, 98570, 98580, 98610, 98620, 98620, 98640, 
    98670, 98670, 98660, 98670, 98720, 98790, 98810, 98830, 98860, 98880, 
    98930, 98950, 98980, 99000, 99030, 99040, 99080, 99140, 99160, 99180, 
    99210, 99220, 99230, 99230, 99240, 99210, 99230, 99230, 99230, 99250, 
    99280, 99280, 99270, 99250, 99240, 99220, 99240, 99220, 99220, 99190, 
    99180, 99140, 99160, 99120, 99040, 99020, 98970, 98970, 98910, 98880, 
    98830, 98730, 98660, 98630, 98590, 98520, 98410, 98340, 98280, 98190, 
    98090, 98000, 97990, 97990, 98000, 97980, 98080, 98050, 98070, 98040, 
    98060, 98060, 98050, 98070, 98060, 98100, 98120, 98160, 98190, 98230, 
    98250, 98280, 98290, 98340, 98350, 98340, 98370, 98370, 98390, 98380, 
    98400, 98430, 98450, 98450, 98440, 98450, 98430, 98460, 98460, 98500, 
    98500, 98530, 98550, 98560, 98580, 98600, 98620, 98630, 98640, 98660, 
    98690, 98720, 98760, 98810, 98890, 98910, 98960, 98960, 99000, 99020, 
    99050, 99060, 99080, 99100, 99100, 99120, 99110, 99120, 99110, 99110, 
    99060, 99070, 99040, 99040, 99050, 99080, 99130, 99200, 99250, 99310, 
    99350, 99390, 99410, 99450, 99470, 99480, 99540, 99570, 99600, 99630, 
    99680, 99690, 99730, 99760, 99770, 99770, 99740, 99740, 99740, 99750, 
    99730, 99710, 99720, 99690, 99670, 99680, 99660, 99580, 99620, 99570, 
    99570, 99610, 99520, 99530, 99540, 99570, 99580, 99570, 99590, 99630, 
    99660, 99660, 99680, 99720, 99740, 99780, 99790, 99840, 99870, 99910, 
    99930, 99940, 99960, 99980, 100010, 100050, 100070, 100120, 100150, 
    100220, 100270, 100340, 100350, 100350, 100310, 100290, 100260, 100180, 
    100080, 99960, 99840, 99740, 99590, 99440, 99270, 99110, 98930, 98740, 
    98510, 98280, 98070, 97950, 97810, 97630, 97490, 97390, 97360, 97370, 
    97370, 97370, 97290, 97180, 97120, 97050, 97020, 96930, 96880, 96880, 
    96850, 96740, 96660, 96650, 96660, 96690, 96670, 96720, 96910, 97050, 
    97170, 97270, 97350, 97370, 97460, 97520, 97580, 97650, 97670, 97680, 
    97750, 97780, 97780, 97800, 97800, 97750, 97710, 97710, 97650, 97650, 
    97640, 97650, 97700, 97730, 97770, 97800, 97830, 97820, 97790, 97770, 
    97780, 97750, 97700, 97650, 97600, 97550, 97530, 97500, 97430, 97470, 
    97510, 97500, 97520, 97540, 97570, 97600, 97610, 97640, 97630, 97590, 
    97540, 97530, 97520, 97510, 97520, 97550, 97550, 97630, 97730, 97840, 
    97940, 97980, 98040, 98100, 98140, 98170, 98220, 98270, 98350, 98420, 
    98520, 98570, 98630, 98680, 98730, 98750, 98820, 98880, 98910, 98960, 
    99090, 99270, 99420, 99560, 99700, 99830, 99930, 100050, 100160, 100240, 
    100330, 100390, 100510, 100590, 100630, 100680, 100750, 100790, 100830, 
    100860, 100900, 100940, 100910, 100920, 100950, 100940, 100940, 100960, 
    100980, 100990, 100980, 100980, 100970, 100990, 101000, 101000, 101000, 
    101000, 101010, 101010, 100970, 100940, 100910, 100870, 100860, 100840, 
    100800, 100790, 100770, 100770, 100770, 100740, 100710, 100670, 100680, 
    100630, 100590, 100580, 100520, 100480, 100420, 100410, 100370, 100330, 
    100300, 100250, 100190, 100090, 99960, 99830, 99690, 99540, 99450, 99350, 
    99290, 99170, 99000, 98870, 98740, 98570, 98440, 98260, 98120, 98080, 
    98040, 97990, 97980, 97940, 98000, 98020, 98010, 98050, 98070, 98130, 
    98180, 98240, 98130, 98210, 98270, 98320, 98370, 98380, 98350, 98340, 
    98340, 98350, 98350, 98390, 98440, 98530, 98610, 98700, 98800, 98880, 
    98970, 99090, 99210, 99340, 99420, 99570, 99660, 99790, 99900, 99960, 
    100000, 100090, 100120, 100140, 100170, 100190, 100150, 100210, 100310, 
    100300, 100320, 100360, 100350, 100310, 100290, 100220, 100180, 100140, 
    100100, 100020, 100010, 100010, 100000, 99950, 99920, 99860, 99750, 
    99720, 99640, 99600, 99510, 99480, 99510, 99510, 99520, 99580, 99620, 
    99640, 99680, 99740, 99810, 99850, 99950, 100020, 100100, 100110, 100120, 
    100130, 100130, 100110, 100100, 100060, 100040, 100020, 100000, 99980, 
    100000, 100010, 100060, 100060, 100070, 100110, 100100, 100070, 100040, 
    100090, 100040, 100030, 100000, 99980, 99970, 99920, 99870, 99830, 99770, 
    99700, 99650, 99600, 99570, 99540, 99520, 99510, 99480, 99450, 99440, 
    99410, 99410, 99420, 99400, 99440, 99420, 99420, 99430, 99450, 99460, 
    99480, 99490, 99490, 99480, 99520, 99640, 99680, 99720, 99760, 99840, 
    99900, 99920, 99930, 99970, 99950, 99900, 99910, 100000, 100050, 100150, 
    100190, 100210, 100310, 100380, 100450, 100510, 100550, 100610, 100670, 
    100770, 100860, 100920, 100920, 100930, 100960, 100950, 100930, 100930, 
    100900, 100960, 101000, 101090, 101120, 101150, 101190, 101260, 101300, 
    101340, 101380, 101380, 101430, 101550, 101500, 101510, 101480, 101520, 
    101510, 101500, 101480, 101460, 101440, 101400, 101350, 101270, 101220, 
    101190, 101140, 101120, 101090, 101050, 101030, 101020, 101000, 100980, 
    100950, 100940, 100920, 100900, 100870, 100830, 100830, 100810, 100780, 
    100790, 100820, 100830, 100830, 100820, 100820, 100790, 100750, 100740, 
    100760, 100760, 100740, 100760, 100750, 100770, 100780, 100750, 100710, 
    100660, 100630, 100600, 100530, 100480, 100420, 100400, 100360, 100320, 
    100300, 100260, 100250, 100250, 100260, 100290, 100310, 100330, 100390, 
    100400, 100400, 100440, 100430, 100470, 100530, 100600, 100620, 100690, 
    100730, 100710, 100750, 100740, 100730, 100670, 100640, 100570, 100520, 
    100420, 100430, 100390, 100370, 100340, 100330, 100310, 100350, 100330, 
    100320, 100310, 100280, 100290, 100290, 100240, 100190, 100250, 100340, 
    100380, 100450, 100500, 100560, 100650, 100670, 100740, 100790, 100800, 
    100850, 100870, 100920, 100970, 101040, 101020, 101050, 101020, 101060, 
    101120, 101130, 101180, 101200, 101240, 101260, 101290, 101280, 101260, 
    101230, 101190, 101140, 101100, 101100, 101080, 101040, 101030, 101070, 
    101090, 101090, 101090, 101110, 101160, 101220, 101290, 101330, 101400, 
    101480, 101540, 101600, 101730, 101840, 101920, 102000, 102070, 102160, 
    102200, 102270, 102340, 102420, 102480, 102520, 102590, 102680, 102740, 
    102740, 102780, 102760, 102720, 102730, 102710, 102680, 102660, 102630, 
    102620, 102630, 102620, 102620, 102610, 102650, 102650, 102640, 102650, 
    102620, 102640, 102640, 102650, 102690, 102650, 102660, 102640, 102640, 
    102610, 102600, 102620, 102600, 102600, 102720, 102720, 102700, 102720, 
    102710, 102670, 102670, 102650, 102610, 102610, 102570, 102570, 102540, 
    102500, 102440, 102390, 102350, 102260, 102120, 102020, 101910, 101810, 
    101640, 101520, 101400, 101320, 101190, 101100, 101080, 100940, 100870, 
    100820, 100840, 100870, 100910, 100910, 100870, 100880, 100870, 100800, 
    100750, 100670, 100600, 100480, 100360, 100240, 100110, 99980, 99880, 
    99740, 99580, 99440, 99330, 99200, 99060, 98900, 98770, 98650, 98510, 
    98400, 98320, 98250, 98210, 98170, 98110, 98120, 98140, 98240, 98330, 
    98360, 98490, 98570, 98720, 98880, 99030, 99130, 99180, 99310, 99370, 
    99400, 99380, 99340, 99410, 99340, 99450, 99590, 99630, 99690, 99760, 
    99840, 99940, 100030, 100120, 100250, 100360, 100430, 100520, 100600, 
    100700, 100760, 100870, 101060, 101160, 101280, 101410, 101500, 101570, 
    101630, 101680, 101760, 101820, 101860, 101890, 101930, 101910, 101880, 
    101860, 101820, 101800, 101740, 101690, 101670, 101620, 101570, 101510, 
    101460, 101350, 101280, 101190, 101120, 101080, 101030, 100990, 100940, 
    100900, 100860, 100740, 100680, 100640, 100610, 100590, 100610, 100600, 
    100550, 100570, 100570, 100550, 100510, 100540, 100510, 100500, 100520, 
    100540, 100480, 100420, 100470, 100540, 100560, 100550, 100560, 100530, 
    100490, 100500, 100520, 100560, 100560, 100540, 100590, 100630, 100630, 
    100630, 100660, 100640, 100640, 100620, 100630, 100610, 100610, 100590, 
    100610, 100620, 100660, 100690, 100690, 100670, 100630, 100640, 100630, 
    100620, 100630, 100620, 100630, 100680, 100680, 100710, 100700, 100690, 
    100650, 100610, 100580, 100580, 100580, 100550, 100550, 100530, 100540, 
    100520, 100510, 100500, 100490, 100470, 100450, 100440, 100390, 100340, 
    100310, 100270, 100240, 100200, 100180, 100120, 100080, 100000, 99980, 
    99910, 99860, 99810, 99750, 99710, 99670, 99650, 99560, 99440, 99350, 
    99270, 99170, 99070, 98960, 98820, 98670, 98590, 98520, 98420, 98330, 
    98380, 98440, 98500, 98530, 98580, 98650, 98730, 98720, 98750, 98870, 
    98930, 98910, 98880, 98900, 98960, 98970, 99040, 99130, 99150, 99180, 
    99250, 99290, 99270, 99330, 99510, 99540, 99540, 99640, 99740, 99700, 
    99680, 99740, 99840, 99960, 100120, 100220, 100170, 100190, 100220, 
    100170, 100200, 100190, 100170, 100160, 100140, 100110, 100060, 100030, 
    99990, 99960, 99930, 99890, 99850, 99790, 99760, 99740, 99720, 99680, 
    99620, 99600, 99640, 99650, 99650, 99630, 99610, 99600, 99560, 99560, 
    99530, 99530, 99540, 99530, 99510, 99480, 99450, 99410, 99350, 99350, 
    99300, 99290, 99270, 99300, 99370, 99420, 99430, 99360, 99370, 99370, 
    99440, 99580, 99470, 99430, 99500, 99490, 99450, 99430, 99360, 99320, 
    99300, 99270, 99310, 99340, 99370, 99390, 99400, 99450, 99460, 99510, 
    99560, 99600, 99570, 99640, 99710, 99760, 99770, 99830, 99870, 99870, 
    99870, 99980, 100000, 100050, 100090, 100110, 100110, 100160, 100190, 
    100270, 100340, 100390, 100430, 100520, 100590, 100650, 100690, 100780, 
    100840, 100870, 100910, 100960, 101020, 101080, 101130, 101190, 101220, 
    101260, 101300, 101340, 101360, 101370, 101390, 101410, 101450, 101480, 
    101510, 101540, 101550, 101570, 101590, 101600, 101580, 101590, 101680, 
    101750, 101780, 101780, 101750, 101760, 101720, 101660, 101640, 101670, 
    101710, 101710, 101690, 101710, 101740, 101740, 101720, 101700, 101660, 
    101630, 101630, 101580, 101520, 101450, 101430, 101390, 101350, 101280, 
    101180, 101160, 101150, 101090, 101010, 100960, 100900, 100870, 100820, 
    100770, 100730, 100720, 100690, 100620, 100570, 100520, 100500, 100570, 
    100540, 100520, 100470, 100450, 100400, 100380, 100350, 100320, 100330, 
    100320, 100340, 100350, 100350, 100350, 100350, 100380, 100390, 100430, 
    100460, 100450, 100500, 100520, 100520, 100540, 100560, 100580, 100590, 
    100620, 100650, 100660, 100680, 100690, 100660, 100670, 100690, 100750, 
    100750, 100740, 100730, 100740, 100760, 100750, 100820, 100850, 100870, 
    100920, 100950, 100990, 100990, 101020, 101090, 101130, 101200, 101230, 
    101240, 101280, 101290, 101310, 101380, 101410, 101420, 101390, 101420, 
    101440, 101480, 101480, 101500, 101470, 101470, 101460, 101460, 101450, 
    101460, 101460, 101420, 101410, 101400, 101380, 101370, 101340, 101320, 
    101290, 101230, 101230, 101270, 101210, 101180, 101170, 101180, 101170, 
    101130, 101130, 101120, 101100, 101100, 101100, 101090, 101080, 101050, 
    100990, 100950, 100910, 100900, 100800, 100720, 100650, 100600, 100510, 
    100520, 100480, 100350, 100350, 100290, 100260, 100250, 100260, 100350, 
    100370, 100480, 100550, 100620, 100670, 100690, 100750, 100830, 100900, 
    100960, 100860, 100820, 100930, 100980, 101060, 101040, 101030, 101040, 
    101080, 101130, 101150, 101190, 101200, 101220, 101250, 101280, 101300, 
    101280, 101290, 101300, 101330, 101360, 101360, 101380, 101420, 101430, 
    101450, 101460, 101450, 101470, 101500, 101490, 101500, 101520, 101550, 
    101570, 101560, 101550, 101510, 101480, 101450, 101390, 101260, 101170, 
    101110, 101060, 100930, 100780, 100740, 100720, 100730, 100670, 100700, 
    100630, 100620, 100630, 100620, 100660, 100680, 100710, 100750, 100800, 
    100870, 100920, 100950, 100980, 101020, 101070, 101120, 101180, 101260, 
    101310, 101370, 101410, 101450, 101450, 101450, 101460, 101470, 101460, 
    101480, 101480, 101490, 101470, 101460, 101460, 101450, 101440, 101410, 
    101360, 101290, 101240, 101180, 101140, 101090, 101040, 101020, 100950, 
    100860, 100720, 100600, 100480, 100350, 100180, 99990, 99890, 99770, 
    99560, 99350, 99180, 99040, 98890, 98700, 98520, 98220, 97810, 97440, 
    97200, 97270, 97190, 97290, 97380, 97450, 97450, 97350, 97370, 97350, 
    97280, 97230, 97200, 97190, 97260, 97290, 97350, 97410, 97500, 97620, 
    97730, 97900, 98070, 98280, 98470, 98640, 98810, 98950, 99070, 99190, 
    99310, 99410, 99460, 99580, 99710, 99850, 99980, 100070, 100170, 100220, 
    100330, 100420, 100550, 100560, 100610, 100630, 100690, 100720, 100700, 
    100700, 100700, 100630, 100530, 100440, 100330, 100280, 100180, 100080, 
    99890, 99830, 99760, 99700, 99590, 99570, 99540, 99570, 99610, 99580, 
    99580, 99530, 99570, 99540, 99540, 99530, 99530, 99540, 99530, 99490, 
    99460, 99440, 99380, 99320, 99200, 99120, 99020, 98920, 98750, 98600, 
    98460, 98430, 98290, 98250, 98170, 98140, 98070, 97950, 97890, 97880, 
    97860, 97840, 97780, 97730, 97670, 97660, 97660, 97680, 97650, 97660, 
    97690, 97720, 97750, 97790, 97870, 97890, 97910, 97940, 97990, 98000, 
    98000, 98030, 98060, 98050, 98050, 98040, 98050, 98040, 98030, 98020, 
    98010, 98000, 97980, 97970, 97920, 97910, 97910, 97860, 97840, 97790, 
    97760, 97730, 97680, 97630, 97620, 97580, 97540, 97510, 97510, 97500, 
    97470, 97460, 97430, 97410, 97380, 97420, 97410, 97420, 97440, 97470, 
    97490, 97530, 97570, 97600, 97620, 97650, 97680, 97720, 97770, 97810, 
    97870, 97920, 97970, 98010, 98020, 98020, 98030, 98040, 98060, 98070, 
    98060, 98070, 98090, 98080, 98080, 98080, 98080, 98100, 98080, 98070, 
    98060, 98100, 98120, 98120, 98150, 98170, 98180, 98210, 98230, 98260, 
    98270, 98270, 98280, 98300, 98350, 98400, 98420, 98400, 98410, 98440, 
    98470, 98450, 98450, 98460, 98460, 98450, 98450, 98450, 98450, 98450, 
    98460, 98480, 98500, 98500, 98520, 98530, 98550, 98570, 98590, 98640, 
    98670, 98720, 98780, 98830, 98880, 98950, 98990, 99060, 99110, 99170, 
    99250, 99290, 99360, 99420, 99470, 99510, 99600, 99680, 99730, 99800, 
    99850, 99900, 99930, 100020, 100060, 100080, 100140, 100220, 100250, 
    100260, 100300, 100330, 100350, 100380, 100400, 100420, 100430, 100430, 
    100440, 100440, 100400, 100420, 100420, 100410, 100390, 100390, 100400, 
    100410, 100390, 100380, 100390, 100400, 100360, 100300, 100280, 100270, 
    100200, 100110, 100040, 100040, 99940, 99960, 99870, 99660, 99640, 99520, 
    99290, 99270, 99240, 99150, 99050, 98980, 98960, 99000, 98940, 98890, 
    98860, 98850, 98880, 98910, 98950, 99000, 99050, 99120, 99190, 99230, 
    99330, 99370, 99440, 99460, 99510, 99520, 99560, 99600, 99620, 99660, 
    99660, 99660, 99710, 99750, 99730, 99740, 99710, 99720, 99660, 99670, 
    99600, 99610, 99620, 99620, 99600, 99590, 99580, 99550, 99600, 99640, 
    99650, 99610, 99700, 99770, 99750, 99780, 99780, 99690, 99650, 99650, 
    99630, 99600, 99510, 99400, 99370, 99300, 99160, 99130, 99010, 98970, 
    98970, 98930, 98870, 98840, 98790, 98840, 98860, 98930, 98890, 98900, 
    98940, 99010, 99080, 99140, 99210, 99280, 99300, 99280, 99350, 99420, 
    99460, 99500, 99520, 99530, 99540, 99550, 99630, 99570, 99520, 99570, 
    99530, 99610, 99630, 99710, 99760, 99740, 99750, 99810, 99870, 99920, 
    100000, 100080, 100040, 100000, 100020, 100100, 100200, 100300, 100360, 
    100430, 100510, 100550, 100610, 100650, 100690, 100710, 100710, 100690, 
    100700, 100740, 100740, 100740, 100710, 100680, 100710, 100720, 100700, 
    100680, 100660, 100690, 100710, 100740, 100730, 100650, 100670, 100630, 
    100650, 100630, 100600, 100570, 100590, 100590, 100610, 100590, 100510, 
    100470, 100440, 100410, 100410, 100410, 100410, 100370, 100360, 100370, 
    100360, 100360, 100290, 100240, 100230, 100190, 100200, 100190, 100180, 
    100220, 100210, 100220, 100230, 100230, 100240, 100260, 100260, 100260, 
    100270, 100300, 100290, 100280, 100290, 100300, 100310, 100320, 100320, 
    100330, 100350, 100360, 100350, 100380, 100390, 100410, 100420, 100460, 
    100500, 100520, 100540, 100550, 100540, 100550, 100560, 100560, 100550, 
    100550, 100580, 100570, 100580, 100600, 100610, 100620, 100650, 100650, 
    100640, 100650, 100650, 100670, 100700, 100730, 100760, 100770, 100770, 
    100810, 100810, 100840, 100830, 100860, 100880, 100870, 100870, 100930, 
    100970, 101000, 100990, 100990, 101010, 101040, 101040, 101010, 101010, 
    101010, 101030, 101050, 101070, 101100, 101140, 101190, 101210, 101190, 
    101130, 101120, 101090, 101090, 101060, 101040, 101000, 100990, 100970, 
    100950, 100880, 100820, 100800, 100760, 100720, 100710, 100700, 100670, 
    100640, 100580, 100550, 100520, 100460, 100430, 100380, 100350, 100340, 
    100320, 100310, 100330, 100280, 100330, 100350, 100360, 100390, 100430, 
    100430, 100450, 100500, 100540, 100560, 100600, 100660, 100660, 100690, 
    100710, 100760, 100770, 100820, 100860, 100870, 100850, 100860, 100890, 
    100970, 101020, 100980, 101110, 101160, 101180, 101200, 101200, 101210, 
    101260, 101260, 101260, 101280, 101280, 101250, 101220, 101230, 101270, 
    101300, 101300, 101310, 101310, 101270, 101210, 101290, 101290, 101270, 
    101230, 101230, 101270, 101290, 101310, 101340, 101360, 101360, 101450, 
    101490, 101490, 101510, 101480, 101430, 101440, 101460, 101510, 101660, 
    101690, 101710, 101700, 101700, 101720, 101700, 101740, 101750, 101780, 
    101810, 101870, 101880, 101880, 101920, 101920, 101960, 101950, 101950, 
    101960, 101970, 101980, 101970, 101960, 101930, 101950, 101950, 101950, 
    101930, 101910, 101840, 101840, 101840, 101830, 101760, 101710, 101680, 
    101640, 101650, 101680, 101700, 101720, 101720, 101690, 101700, 101730, 
    101740, 101730, 101730, 101720, 101720, 101730, 101740, 101700, 101680, 
    101640, 101640, 101620, 101610, 101600, 101580, 101580, 101580, 101570, 
    101570, 101560, 101560, 101550, 101540, 101510, 101520, 101500, 101490, 
    101470, 101470, 101440, 101430, 101400, 101370, 101360, 101360, 101350, 
    101340, 101330, 101330, 101320, 101340, 101330, 101340, 101360, 101380, 
    101370, 101390, 101410, 101400, 101420, 101430, 101430, 101440, 101490, 
    101500, 101510, 101550, 101560, 101580, 101580, 101590, 101600, 101640, 
    101650, 101690, 101750, 101760, 101790, 101820, 101850, 101880, 101910, 
    101910, 101930, 101930, 101950, 101980, 102000, 102030, 102060, 102080, 
    102100, 102130, 102150, 102180, 102180, 102200, 102220, 102240, 102270, 
    102270, 102270, 102270, 102280, 102290, 102290, 102270, 102260, 102250, 
    102240, 102230, 102220, 102190, 102170, 102170, 102150, 102130, 102110, 
    102090, 102060, 102070, 102050, 102030, 102030, 102020, 102010, 101980, 
    101960, 101920, 101860, 101770, 101720, 101660, 101610, 101560, 101540, 
    101530, 101550, 101630, 101620, 101650, 101680, 101690, 101730, 101750, 
    101670, 101850, 101770, 101970, 101970, 101960, 101960, 101910, 101860, 
    101890, 101920, 101910, 101950, 101990, 101920, 101960, 101950, 101970, 
    101930, 101900, 101910, 101860, 101840, 101860, 101850, 101820, 101740, 
    101750, 101630, 101580, 101580, 101500, 101470, 101530, 101500, 101480, 
    101530, 101540, 101600, 101640, 101660, 101670, 101690, 101720, 101750, 
    101770, 101780, 101780, 101760, 101780, 101800, 101840, 101880, 101920, 
    101930, 101930, 101950, 101950, 101960, 101950, 101970, 101970, 101980, 
    101990, 102010, 102030, 102020, 102030, 102050, 102050, 102060, 102070, 
    102080, 102090, 102110, 102120, 102150, 102150, 102160, 102150, 102150, 
    102140, 102120, 102100, 102060, 102040, 102100, 102080, 102050, 102030, 
    102030, 102020, 102000, 101980, 101960, 101940, 101920, 101930, 101920, 
    101900, 101890, 101880, 101840, 101840, 101810, 101800, 101780, 101750, 
    101740, 101730, 101720, 101740, 101730, 101750, 101770, 101790, 101790, 
    101800, 101810, 101830, 101840, 101840, 101770, 101830, 101820, 101810, 
    101780, 101780, 101710, 101590, 101470, 101470, 101480, 101490, 101500, 
    101510, 101510, 101500, 101520, 101540, 101530, 101620, 101650, 101610, 
    101600, 101640, 101630, 101640, 101600, 101530, 101510, 101550, 101530, 
    101560, 101580, 101630, 101590, 101530, 101500, 101500, 101500, 101480, 
    101490, 101440, 101390, 101360, 101360, 101450, 101460, 101480, 101510, 
    101530, 101560, 101570, 101580, 101600, 101590, 101610, 101630, 101660, 
    101660, 101680, 101720, 101760, 101770, 101760, 101760, 101760, 101780, 
    101750, 101750, 101770, 101810, 101790, 101810, 101790, 101770, 101750, 
    101730, 101680, 101560, 101560, 101600, 101620, 101610, 101600, 101600, 
    101590, 101600, 101560, 101540, 101520, 101490, 101480, 101470, 101450, 
    101440, 101420, 101410, 101430, 101390, 101330, 101330, 101300, 101310, 
    101310, 101280, 101270, 101280, 101280, 101240, 101220, 101180, 101170, 
    101160, 101160, 101150, 101140, 101140, 101090, 101110, 101130, 101150, 
    101190, 101190, 101190, 101200, 101190, 101230, 101250, 101250, 101260, 
    101260, 101240, 101230, 101200, 101230, 101220, 101240, 101220, 101180, 
    101150, 101160, 101130, 101110, 101110, 101120, 101120, 101130, 101150, 
    101190, 101210, 101200, 101230, 101230, 101230, 101280, 101320, 101320, 
    101350, 101380, 101400, 101380, 101400, 101420, 101430, 101430, 101450, 
    101460, 101490, 101510, 101500, 101530, 101520, 101500, 101490, 101480, 
    101450, 101440, 101410, 101390, 101310, 101240, 101170, 101080, 101010, 
    100930, 100880, 100820, 100750, 100710, 100720, 100810, 100790, 100820, 
    100840, 100860, 100920, 100990, 101030, 101030, 101070, 101080, 101080, 
    101090, 101070, 101090, 101040, 101020, 100990, 100930, 100920, 100860, 
    100810, 100780, 100730, 100690, 100660, 100620, 100600, 100540, 100580, 
    100590, 100590, 100610, 100650, 100660, 100690, 100680, 100720, 100740, 
    100720, 100750, 100750, 100780, 100780, 100820, 100840, 100910, 101050, 
    101140, 101280, 101400, 101480, 101560, 101650, 101710, 101830, 101900, 
    102000, 102090, 102140, 102260, 102340, 102450, 102520, 102560, 102630, 
    102670, 102740, 102780, 102810, 102850, 102920, 102940, 102950, 103020, 
    103050, 103060, 103090, 103080, 103070, 103090, 103070, 103060, 103040, 
    103020, 102990, 102970, 102930, 102900, 102850, 102800, 102770, 102720, 
    102680, 102630, 102550, 102510, 102470, 102440, 102420, 102370, 102310, 
    102260, 102200, 102170, 102060, 102030, 101990, 102000, 102000, 102000, 
    102010, 101990, 101970, 101980, 101980, 101990, 102040, 102100, 102150, 
    102170, 102210, 102230, 102250, 102270, 102320, 102340, 102340, 102340, 
    102340, 102350, 102380, 102410, 102430, 102450, 102470, 102490, 102520, 
    102520, 102480, 102460, 102500, 102490, 102480, 102450, 102420, 102370, 
    102340, 102240, 102150, 102080, 101980, 101880, 101780, 101670, 101550, 
    101490, 101400, 101280, 101200, 101210, 101120, 101100, 101090, 101020, 
    100990, 100970, 100960, 100980, 100940, 100970, 100990, 101020, 101060, 
    101070, 101140, 101180, 101210, 101280, 101350, 101410, 101440, 101470, 
    101510, 101520, 101560, 101590, 101650, 101690, 101720, 101740, 101780, 
    101800, 101790, 101840, 101920, 102020, 102080, 102100, 102120, 102130, 
    102140, 102170, 102210, 102200, 102220, 102230, 102250, 102270, 102230, 
    102230, 102220, 102170, 102160, 102130, 102150, 102160, 102160, 102170, 
    102200, 102210, 102180, 102200, 102280, 102190, 102190, 102200, 102250, 
    102240, 102230, 102270, 102210, 102300, 102330, 102290, 102320, 102390, 
    102560, 102490, 102470, 102490, 102530, 102540, 102630, 102640, 102640, 
    102650, 102680, 102720, 102750, 102770, 102790, 102810, 102810, 102840, 
    102840, 102820, 102810, 102790, 102830, 102830, 102850, 102860, 102870, 
    102870, 102890, 102890, 102910, 102930, 102960, 102960, 102960, 102960, 
    102940, 102920, 102910, 102910, 102900, 102870, 102870, 102840, 102830, 
    102800, 102800, 102790, 102780, 102770, 102770, 102760, 102790, 102850, 
    102880, 102930, 102940, 102990, 103020, 103060, 103080, 103110, 103140, 
    103160, 103180, 103180, 103220, 103230, 103230, 103230, 103230, 103230, 
    103220, 103230, 103220, 103230, 103240, 103220, 103210, 103200, 103190, 
    103170, 103160, 103150, 103110, 103100, 103070, 103060, 103080, 103070, 
    103040, 103030, 103030, 103010, 103000, 102980, 102960, 102950, 102940, 
    102970, 102960, 102990, 102980, 102990, 102980, 102970, 102950, 102940, 
    102950, 102950, 102930, 102940, 102960, 102960, 102970, 102950, 102960, 
    102940, 102930, 102920, 102900, 102910, 102920, 102940, 102950, 102960, 
    102980, 102980, 102970, 102960, 102960, 102930, 102930, 102910, 102900, 
    102900, 102900, 102880, 102870, 102860, 102830, 102800, 102800, 102780, 
    102770, 102750, 102770, 102770, 102780, 102770, 102800, 102810, 102790, 
    102810, 102820, 102820, 102820, 102800, 102780, 102760, 102790, 102760, 
    102760, 102740, 102710, 102690, 102680, 102660, 102630, 102620, 102620, 
    102640, 102640, 102620, 102620, 102630, 102600, 102580, 102570, 102550, 
    102500, 102430, 102360, 102290, 102230, 102180, 102110, 102050, 101950, 
    101860, 101790, 101710, 101630, 101530, 101460, 101400, 101310, 101250, 
    101170, 101130, 101100, 101130, 101180, 101230, 101270, 101310, 101310, 
    101320, 101370, 101410, 101450, 101480, 101440, 101430, 101460, 101470, 
    101460, 101450, 101440, 101430, 101420, 101420, 101450, 101430, 101400, 
    101380, 101390, 101410, 101430, 101420, 101400, 101440, 101410, 101480, 
    101530, 101560, 101650, 101670, 101660, 101660, 101710, 101720, 101760, 
    101730, 101790, 101950, 101970, 101970, 101920, 101940, 102030, 102050, 
    102070, 102070, 102070, 102090, 102070, 102080, 102120, 102070, 102090, 
    102090, 102090, 102080, 102080, 102080, 102080, 102100, 102110, 102110, 
    102090, 102100, 102110, 102120, 102120, 102110, 102090, 102080, 102040, 
    102030, 102040, 102040, 102030, 102010, 102000, 101990, 102000, 102000, 
    101980, 101980, 101980, 101990, 101990, 102020, 102030, 102020, 102000, 
    102000, 101990, 101980, 101970, 101970, 101960, 101950, 101940, 101940, 
    101930, 101930, 101900, 101910, 101910, 101910, 101890, 101850, 101850, 
    101860, 101850, 101860, 101870, 101880, 101850, 101830, 101810, 101770, 
    101760, 101730, 101700, 101690, 101660, 101630, 101590, 101570, 101530, 
    101510, 101470, 101420, 101350, 101290, 101240, 101200, 101180, 101150, 
    101110, 101060, 101020, 100990, 100940, 100890, 100840, 100780, 100730, 
    100710, 100670, 100630, 100600, 100580, 100590, 100580, 100560, 100530, 
    100510, 100490, 100460, 100430, 100410, 100400, 100390, 100380, 100390, 
    100350, 100310, 100260, 100220, 100210, 100180, 100170, 100170, 100190, 
    100210, 100240, 100260, 100280, 100280, 100300, 100330, 100350, 100370, 
    100400, 100430, 100470, 100520, 100540, 100570, 100590, 100610, 100640, 
    100650, 100680, 100690, 100710, 100720, 100740, 100760, 100780, 100790, 
    100810, 100820, 100840, 100860, 100870, 100870, 100870, 100900, 100900, 
    100920, 100940, 100950, 100980, 101000, 101010, 101050, 101090, 101110, 
    101110, 101110, 101100, 101100, 101080, 101080, 101050, 101020, 100990, 
    100980, 100930, 100990, 101030, 101050, 101070, 101080, 101080, 101110, 
    101130, 101130, 101120, 101120, 101140, 101140, 101130, 101130, 101130, 
    101120, 101140, 101150, 101150, 101150, 101170, 101180, 101200, 101190, 
    101210, 101240, 101260, 101300, 101320, 101350, 101370, 101410, 101420, 
    101430, 101430, 101440, 101440, 101460, 101490, 101530, 101570, 101610, 
    101640, 101670, 101690, 101720, 101740, 101790, 101840, 101870, 101910, 
    101950, 101990, 102020, 102050, 102080, 102080, 102110, 102120, 102140, 
    102130, 102150, 102160, 102180, 102200, 102200, 102210, 102210, 102180, 
    102150, 102120, 102140, 102130, 102120, 102120, 102090, 102120, 102110, 
    102070, 102060, 102010, 101980, 101960, 101900, 101880, 101840, 101810, 
    101800, 101710, 101610, 101590, 101520, 101480, 101400, 101280, 101220, 
    101220, 101150, 101090, 101120, 101090, 101110, 101090, 101060, 101030, 
    101050, 101060, 101080, 101110, 101150, 101190, 101230, 101270, 101290, 
    101300, 101330, 101330, 101340, 101370, 101360, 101380, 101410, 101450, 
    101420, 101450, 101480, 101530, 101560, 101640, 101690, 101700, 101710, 
    101740, 101820, 101850, 101910, 101880, 101880, 101910, 101900, 101970, 
    101950, 101980, 102020, 102030, 102070, 102080, 102100, 102100, 102140, 
    102210, 102210, 102260, 102280, 102320, 102360, 102390, 102430, 102440, 
    102480, 102500, 102530, 102580, 102590, 102620, 102640, 102650, 102670, 
    102690, 102760, 102790, 102790, 102830, 102860, 102880, 102900, 102930, 
    102930, 102940, 102990, 103000, 102990, 103000, 102980, 102970, 102960, 
    102940, 102960, 102940, 102920, 102910, 102890, 102870, 102880, 102870, 
    102840, 102830, 102820, 102800, 102780, 102750, 102720, 102700, 102680, 
    102650, 102600, 102550, 102510, 102470, 102450, 102400, 102370, 102320, 
    102290, 102260, 102230, 102250, 102210, 102200, 102210, 102180, 102180, 
    102190, 102200, 102190, 102190, 102210, 102200, 102210, 102220, 102230, 
    102250, 102250, 102260, 102270, 102280, 102310, 102330, 102340, 102350, 
    102340, 102350, 102380, 102380, 102380, 102400, 102410, 102400, 102430, 
    102420, 102430, 102430, 102440, 102420, 102410, 102370, 102350, 102330, 
    102320, 102310, 102300, 102300, 102260, 102260, 102240, 102260, 102240, 
    102250, 102240, 102220, 102230, 102250, 102230, 102210, 102210, 102190, 
    102180, 102190, 102180, 102160, 102130, 102140, 102140, 102100, 102110, 
    102110, 102120, 102110, 102110, 102120, 102110, 102110, 102100, 102110, 
    102110, 102110, 102120, 102140, 102110, 102090, 102090, 102090, 102050, 
    102030, 102040, 102040, 102010, 102010, 102020, 102030, 101990, 101940, 
    101950, 101970, 101990, 101990, 101980, 102000, 101990, 101980, 101960, 
    101970, 101970, 101980, 101980, 101990, 101990, 102030, 102060, 102090, 
    102110, 102130, 102190, 102240, 102270, 102310, 102360, 102420, 102490, 
    102540, 102600, 102630, 102650, 102690, 102720, 102740, 102770, 102790, 
    102810, 102800, 102820, 102830, 102820, 102840, 102820, 102790, 102800, 
    102770, 102770, 102760, 102720, 102730, 102710, 102690, 102680, 102640, 
    102620, 102620, 102600, 102540, 102510, 102460, 102430, 102470, 102440, 
    102410, 102410, 102350, 102340, 102310, 102280, 102240, 102250, 102250, 
    102250, 102300, 102350, 102360, 102380, 102390, 102390, 102350, 102330, 
    102300, 102230, 102180, 102120, 102040, 101960, 101840, 101720, 101650, 
    101560, 101510, 101480, 101440, 101420, 101460, 101480, 101470, 101460, 
    101480, 101480, 101510, 101480, 101470, 101480, 101470, 101440, 101410, 
    101370, 101320, 101280, 101270, 101230, 101210, 101200, 101170, 101120, 
    101040, 101010, 100970, 100940, 100900, 100920, 100920, 100900, 100900, 
    100910, 100900, 100880, 100880, 100850, 100850, 100810, 100810, 100790, 
    100740, 100730, 100690, 100720, 100700, 100680, 100650, 100590, 100540, 
    100530, 100560, 100520, 100480, 100420, 100430, 100430, 100360, 100320, 
    100280, 100120, 100110, 100100, 100080, 100050, 100020, 100010, 99920, 
    99850, 99800, 99770, 99720, 99710, 99720, 99780, 99820, 99890, 99910, 
    99930, 100010, 100060, 100110, 100180, 100200, 100180, 100230, 100280, 
    100300, 100330, 100340, 100350, 100360, 100370, 100380, 100380, 100380, 
    100380, 100370, 100390, 100380, 100400, 100400, 100400, 100370, 100370, 
    100370, 100370, 100330, 100330, 100320, 100320, 100310, 100320, 100320, 
    100330, 100340, 100320, 100330, 100330, 100350, 100370, 100370, 100400, 
    100410, 100440, 100470, 100510, 100530, 100540, 100550, 100550, 100580, 
    100590, 100580, 100580, 100590, 100610, 100630, 100630, 100620, 100590, 
    100570, 100580, 100580, 100580, 100580, 100570, 100580, 100600, 100610, 
    100610, 100620, 100610, 100610, 100600, 100620, 100610, 100600, 100570, 
    100570, 100590, 100590, 100610, 100620, 100610, 100600, 100590, 100580, 
    100580, 100560, 100560, 100570, 100590, 100600, 100610, 100600, 100610, 
    100600, 100630, 100620, 100600, 100600, 100590, 100580, 100580, 100570, 
    100560, 100570, 100560, 100540, 100490, 100470, 100450, 100420, 100410, 
    100410, 100430, 100430, 100390, 100380, 100360, 100350, 100330, 100330, 
    100330, 100350, 100360, 100370, 100390, 100400, 100420, 100430, 100450, 
    100460, 100470, 100500, 100520, 100520, 100560, 100570, 100620, 100650, 
    100670, 100670, 100690, 100690, 100700, 100720, 100730, 100730, 100730, 
    100750, 100750, 100750, 100770, 100760, 100770, 100770, 100770, 100760, 
    100760, 100780, 100800, 100810, 100820, 100820, 100830, 100830, 100840, 
    100850, 100860, 100850, 100870, 100880, 100850, 100850, 100850, 100860, 
    100880, 100880, 100860, 100860, 100850, 100850, 100850, 100830, 100860, 
    100860, 100870, 100870, 100880, 100910, 100910, 100900, 100890, 100890, 
    100900, 100900, 100910, 100920, 100910, 100910, 100910, 100890, 100900, 
    100910, 100910, 100920, 100910, 100880, 100890, 100900, 100930, 100930, 
    100930, 100930, 100920, 100900, 100910, 100890, 100900, 100900, 100910, 
    100900, 100890, 100900, 100910, 100920, 100920, 100920, 100920, 100910, 
    100900, 100900, 100920, 100930, 100930, 100940, 100940, 100940, 100940, 
    100960, 100950, 100950, 100940, 100950, 100940, 100950, 100960, 100980, 
    100980, 100980, 100960, 100960, 100950, 100950, 100940, 100920, 100930, 
    100940, 100950, 100970, 100960, 100930, 100910, 100880, 100860, 100860, 
    100850, 100830, 100810, 100780, 100780, 100750, 100740, 100710, 100680, 
    100660, 100640, 100620, 100590, 100580, 100570, 100560, 100580, 100570, 
    100560, 100540, 100530, 100510, 100500, 100460, 100450, 100460, 100440, 
    100440, 100400, 100350, 100330, 100290, 100260, 100230, 100240, 100220, 
    100250, 100210, 100210, 100230, 100250, 100240, 100260, 100260, 100250, 
    100220, 100220, 100230, 100240, 100220, 100230, 100240, 100270, 100270, 
    100280, 100290, 100310, 100330, 100330, 100350, 100340, 100350, 100370, 
    100380, 100360, 100330, 100330, 100360, 100350, 100330, 100300, 100270, 
    100220, 100170, 100130, 100100, 100070, 100060, 100040, 100000, 99990, 
    99970, 99980, 99980, 99980, 100000, 100030, 100070, 100110, 100140, 
    100210, 100250, 100300, 100350, 100400, 100450, 100500, 100530, 100540, 
    100620, 100680, 100740, 100820, 100880, 100930, 100960, 100980, 101030, 
    101040, 101070, 101100, 101150, 101180, 101230, 101260, 101280, 101300, 
    101300, 101300, 101300, 101280, 101250, 101290, 101300, 101360, 101390, 
    101420, 101430, 101430, 101390, 101390, 101370, 101380, 101410, 101390, 
    101390, 101390, 101410, 101470, 101510, 101540, 101540, 101480, 101490, 
    101450, 101470, 101490, 101530, 101550, 101550, 101530, 101500, 101500, 
    101490, 101480, 101480, 101470, 101460, 101440, 101470, 101500, 101480, 
    101480, 101480, 101490, 101480, 101490, 101470, 101470, 101480, 101480, 
    101470, 101490, 101490, 101480, 101480, 101470, 101460, 101470, 101450, 
    101450, 101420, 101400, 101420, 101400, 101430, 101410, 101410, 101380, 
    101350, 101320, 101300, 101250, 101230, 101200, 101160, 101140, 101100, 
    101060, 101010, 100980, 100910, 100840, 100810, 100770, 100700, 100680, 
    100640, 100590, 100550, 100540, 100490, 100450, 100380, 100330, 100260, 
    100210, 100180, 100140, 100100, 100060, 100060, 100050, 100020, 100010, 
    99990, 99990, 100000, 100000, 99990, 100000, 100030, 100050, 100070, 
    100110, 100130, 100150, 100170, 100200, 100180, 100180, 100230, 100270, 
    100310, 100340, 100380, 100400, 100410, 100410, 100410, 100440, 100440, 
    100460, 100490, 100470, 100480, 100550, 100610, 100660, 100670, 100670, 
    100730, 100730, 100730, 100750, 100780, 100780, 100780, 100820, 100800, 
    100800, 100810, 100800, 100780, 100750, 100760, 100750, 100770, 100800, 
    100780, 100790, 100780, 100780, 100740, 100700, 100660, 100630, 100590, 
    100540, 100480, 100430, 100340, 100250, 100190, 100080, 99990, 99950, 
    99860, 99810, 99710, 99640, 99630, 99550, 99520, 99520, 99500, 99530, 
    99540, 99570, 99630, 99650, 99720, 99760, 99780, 99790, 99840, 99880, 
    99910, 99940, 99990, 100020, 100040, 100090, 100130, 100160, 100210, 
    100260, 100320, 100340, 100400, 100450, 100470, 100480, 100510, 100530, 
    100560, 100580, 100610, 100620, 100640, 100650, 100690, 100690, 100700, 
    100690, 100690, 100680, 100690, 100700, 100720, 100730, 100750, 100780, 
    100780, 100810, 100820, 100830, 100850, 100860, 100880, 100900, 100910, 
    100930, 100940, 100950, 100950, 100970, 100980, 100990, 100980, 100960, 
    100970, 100990, 100980, 101000, 101000, 100990, 101010, 101030, 101020, 
    101010, 101010, 101000, 101000, 100970, 100940, 100930, 100910, 100910, 
    100910, 100900, 100880, 100880, 100870, 100870, 100860, 100870, 100880, 
    100880, 100890, 100880, 100900, 100910, 100920, 100940, 100940, 100910, 
    100920, 100950, 100970, 101000, 100980, 100970, 101010, 100990, 100970, 
    101000, 100980, 100910, 100960, 100950, 100920, 100880, 100840, 100800, 
    100770, 100700, 100570, 100430, 100330, 100210, 100170, 100020, 99840, 
    99760, 99550, 99530, 99410, 99380, 99440, 99450, 99480, 99490, 99540, 
    99590, 99650, 99710, 99740, 99760, 99780, 99810, 99890, 99940, 99970, 
    100010, 100060, 100150, 100200, 100230, 100300, 100370, 100470, 100530, 
    100600, 100670, 100760, 100850, 100940, 101000, 101060, 101140, 101190, 
    101260, 101330, 101370, 101380, 101390, 101410, 101460, 101480, 101500, 
    101490, 101500, 101490, 101470, 101430, 101460, 101440, 101390, 101360, 
    101300, 101300, 101230, 101150, 101060, 100960, 100900, 100770, 100700, 
    100590, 100460, 100380, 100190, 100290, 100240, 100280, 100240, 100270, 
    100300, 100320, 100350, 100400, 100450, 100490, 100540, 100570, 100600, 
    100600, 100630, 100680, 100740, 100730, 100730, 100730, 100730, 100740, 
    100760, 100730, 100760, 100780, 100800, 100820, 100850, 100940, 100940, 
    100980, 101070, 101070, 101100, 101160, 101190, 101220, 101220, 101270, 
    101280, 101280, 101330, 101310, 101280, 101310, 101300, 101270, 101240, 
    101220, 101210, 101210, 101220, 101200, 101190, 101110, 101030, 100910, 
    100910, 100840, 100800, 100790, 100700, 100660, 100640, 100570, 100560, 
    100510, 100510, 100540, 100540, 100550, 100550, 100550, 100580, 100580, 
    100600, 100630, 100670, 100740, 100790, 100800, 100780, 100790, 100860, 
    100900, 100920, 100920, 100930, 100920, 100880, 100860, 100800, 100720, 
    100630, 100580, 100560, 100550, 100530, 100520, 100500, 100520, 100550, 
    100570, 100590, 100620, 100640, 100670, 100700, 100770, 100800, 100880, 
    100910, 100960, 101030, 101090, 101150, 101200, 101250, 101300, 101370, 
    101400, 101460, 101530, 101580, 101630, 101680, 101730, 101760, 101790, 
    101800, 101810, 101730, 101780, 101780, 101760, 101760, 101740, 101710, 
    101670, 101620, 101540, 101490, 101450, 101360, 101310, 101260, 101180, 
    101090, 101040, 100980, 100920, 100930, 100920, 100950, 100970, 101030, 
    101090, 101150, 101250, 101310, 101390, 101440, 101490, 101490, 101540, 
    101540, 101630, 101660, 101700, 101710, 101750, 101740, 101750, 101720, 
    101720, 101680, 101660, 101650, 101640, 101600, 101570, 101560, 101560, 
    101550, 101530, 101560, 101530, 101500, 101470, 101430, 101400, 101390, 
    101390, 101350, 101330, 101310, 101300, 101240, 101280, 101270, 101270, 
    101260, 101240, 101230, 101190, 101210, 101220, 101270, 101300, 101330, 
    101350, 101360, 101370, 101400, 101420, 101440, 101460, 101480, 101500, 
    101500, 101510, 101550, 101560, 101560, 101560, 101540, 101530, 101530, 
    101540, 101500, 101480, 101470, 101450, 101450, 101400, 101370, 101340, 
    101310, 101260, 101240, 101210, 101170, 101170, 101140, 101090, 101080, 
    101040, 101000, 100940, 100910, 100880, 100870, 100820, 100760, 100760, 
    100710, 100710, 100690, 100670, 100640, 100590, 100570, 100520, 100490, 
    100460, 100440, 100430, 100420, 100420, 100400, 100400, 100390, 100380, 
    100370, 100390, 100400, 100410, 100420, 100440, 100480, 100520, 100510, 
    100520, 100540, 100560, 100590, 100610, 100600, 100620, 100660, 100640, 
    100670, 100640, 100640, 100760, 100810, 100820, 100830, 100800, 100800, 
    100810, 100930, 100950, 100940, 100970, 101010, 101060, 101060, 101040, 
    101110, 101110, 101160, 101200, 101230, 101260, 101280, 101220, 101220, 
    101210, 101230, 101210, 101210, 101200, 101180, 101180, 101170, 101160, 
    101150, 101140, 101130, 101120, 101090, 101090, 101080, 101070, 101070, 
    101060, 101080, 101040, 101020, 101020, 101030, 101020, 101000, 100940, 
    100900, 100850, 100790, 100770, 100770, 100750, 100740, 100720, 100700, 
    100640, 100630, 100600, 100580, 100550, 100560, 100580, 100580, 100620, 
    100630, 100630, 100630, 100590, 100620, 100640, 100700, 100680, 100630, 
    100660, 100670, 100710, 100740, 100750, 100750, 100750, 100720, 100710, 
    100710, 100670, 100690, 100680, 100680, 100690, 100670, 100690, 100690, 
    100680, 100640, 100640, 100630, 100640, 100640, 100640, 100650, 100660, 
    100690, 100710, 100730, 100730, 100730, 100720, 100740, 100750, 100780, 
    100800, 100820, 100870, 100890, 100910, 100930, 100900, 100890, 100890, 
    100890, 100890, 100860, 100860, 100870, 100870, 100850, 100880, 100880, 
    100870, 100880, 100880, 100870, 100870, 100880, 100910, 100920, 100950, 
    100940, 100960, 100940, 100950, 100930, 100930, 100930, 100930, 100950, 
    100960, 100990, 101010, 101050, 101060, 101090, 101100, 101110, 101110, 
    101110, 101110, 101100, 101110, 101110, 101120, 101120, 101120, 101110, 
    101120, 101090, 101090, 101090, 101080, 101080, 101050, 101100, 101110, 
    101120, 101140, 101170, 101180, 101200, 101220, 101230, 101260, 101300, 
    101320, 101360, 101380, 101410, 101440, 101480, 101490, 101510, 101520, 
    101520, 101530, 101550, 101570, 101600, 101620, 101620, 101650, 101660, 
    101670, 101680, 101670, 101670, 101650, 101640, 101620, 101620, 101600, 
    101600, 101610, 101590, 101590, 101570, 101560, 101560, 101530, 101520, 
    101510, 101500, 101490, 101500, 101500, 101530, 101530, 101550, 101550, 
    101540, 101530, 101530, 101500, 101480, 101480, 101490, 101490, 101510, 
    101500, 101510, 101510, 101490, 101490, 101480, 101480, 101510, 101550, 
    101600, 101650, 101690, 101700, 101750, 101770, 101800, 101810, 101830, 
    101840, 101850, 101880, 101890, 101920, 101950, 101980, 102000, 102010, 
    102030, 102040, 102060, 102050, 102090, 102100, 102120, 102150, 102160, 
    102150, 102130, 102110, 102120, 102100, 102090, 102080, 102050, 102080, 
    102080, 102050, 102050, 102010, 101970, 101950, 101910, 101880, 101860, 
    101840, 101850, 101850, 101850, 101850, 101830, 101860, 101850, 101840, 
    101830, 101830, 101840, 101850, 101830, 101830, 101830, 101830, 101830, 
    101820, 101800, 101760, 101740, 101730, 101720, 101720, 101730, 101700, 
    101720, 101730, 101700, 101680, 101640, 101620, 101590, 101570, 101520, 
    101510, 101480, 101430, 101390, 101360, 101330, 101280, 101250, 101220, 
    101190, 101180, 101160, 101120, 101130, 101100, 101100, 101090, 101060, 
    101020, 100980, 100960, 100960, 100910, 100880, 100860, 100860, 100840, 
    100810, 100770, 100740, 100770, 100680, 100640, 100680, 100660, 100630, 
    100660, 100650, 100560, 100570, 100510, 100500, 100490, 100460, 100460, 
    100410, 100400, 100310, 100290, 100260, 100210, 100110, 100050, 100030, 
    100010, 99980, 99890, 99850, 99810, 99740, 99740, 99710, 99610, 99600, 
    99580, 99580, 99520, 99460, 99430, 99360, 99300, 99200, 99280, 99310, 
    99330, 99290, 99260, 99220, 99200, 99170, 99130, 99090, 99080, 99070, 
    99060, 99030, 99030, 99040, 99040, 99060, 99090, 99130, 99100, 99160, 
    99160, 99130, 99180, 99210, 99250, 99250, 99280, 99300, 99320, 99350, 
    99350, 99330, 99350, 99370, 99400, 99420, 99460, 99440, 99500, 99550, 
    99560, 99590, 99590, 99620, 99660, 99740, 99810, 99850, 99890, 99970, 
    100050, 100140, 100190, 100250, 100280, 100280, 100280, 100270, 100280, 
    100290, 100290, 100280, 100250, 100230, 100210, 100220, 100240, 100250, 
    100260, 100280, 100360, 100400, 100440, 100470, 100490, 100470, 100480, 
    100530, 100550, 100570, 100520, 100600, 100660, 100690, 100690, 100690, 
    100730, 100810, 100790, 100810, 100820, 100830, 100850, 100880, 100920, 
    100930, 100980, 100990, 100970, 100950, 100920, 100940, 100910, 100870, 
    100860, 100850, 100850, 100860, 100860, 100850, 100860, 100850, 100840, 
    100840, 100840, 100790, 100760, 100730, 100710, 100670, 100650, 100640, 
    100650, 100640, 100660, 100680, 100680, 100690, 100690, 100710, 100720, 
    100700, 100730, 100740, 100740, 100740, 100730, 100730, 100700, 100640, 
    100620, 100610, 100550, 100530, 100490, 100460, 100420, 100390, 100340, 
    100350, 100340, 100320, 100290, 100250, 100220, 100210, 100220, 100230, 
    100230, 100250, 100240, 100220, 100200, 100190, 100180, 100190, 100180, 
    100130, 100180, 100200, 100230, 100240, 100290, 100380, 100490, 100580, 
    100650, 100720, 100780, 100830, 100920, 100990, 101050, 101110, 101160, 
    101200, 101220, 101260, 101270, 101290, 101330, 101360, 101390, 101420, 
    101450, 101480, 101510, 101520, 101520, 101500, 101510, 101510, 101520, 
    101520, 101510, 101520, 101560, 101580, 101610, 101630, 101650, 101650, 
    101660, 101660, 101670, 101670, 101680, 101670, 101680, 101680, 101670, 
    101670, 101670, 101650, 101620, 101630, 101640, 101670, 101660, 101670, 
    101660, 101640, 101650, 101620, 101600, 101560, 101530, 101510, 101500, 
    101450, 101420, 101380, 101360, 101350, 101350, 101310, 101300, 101260, 
    101240, 101220, 101220, 101210, 101200, 101190, 101170, 101130, 101130, 
    101130, 101090, 101030, 101010, 100990, 100940, 100910, 100860, 100830, 
    100840, 100840, 100790, 100750, 100710, 100680, 100630, 100580, 100560, 
    100520, 100500, 100440, 100380, 100330, 100280, 100210, 100150, 100140, 
    100150, 100140, 100150, 100170, 100190, 100230, 100290, 100320, 100360, 
    100370, 100400, 100430, 100450, 100470, 100480, 100520, 100560, 100590, 
    100630, 100640, 100630, 100590, 100610, 100600, 100580, 100550, 100550, 
    100520, 100490, 100470, 100430, 100400, 100350, 100310, 100230, 100140, 
    100000, 99930, 99880, 99880, 99850, 99880, 99890, 99920, 99930, 99920, 
    99900, 99890, 99870, 99850, 99810, 99780, 99730, 99700, 99650, 99640, 
    99630, 99630, 99610, 99590, 99570, 99540, 99540, 99550, 99540, 99550, 
    99550, 99560, 99590, 99600, 99590, 99580, 99540, 99520, 99510, 99510, 
    99500, 99480, 99450, 99410, 99380, 99320, 99230, 99150, 99100, 99060, 
    99000, 98920, 98860, 98840, 98790, 98800, 98780, 98760, 98760, 98770, 
    98800, 98800, 98800, 98850, 98860, 98880, 98910, 98950, 98950, 99000, 
    99010, 99050, 99080, 99110, 99170, 99220, 99300, 99290, 99360, 99410, 
    99480, 99560, 99610, 99710, 99760, 99770, 99820, 99890, 99960, 100000, 
    100120, 100220, 100260, 100330, 100360, 100360, 100390, 100460, 100490, 
    100510, 100520, 100580, 100600, 100620, 100650, 100660, 100680, 100680, 
    100700, 100710, 100720, 100730, 100730, 100770, 100770, 100800, 100810, 
    100830, 100840, 100860, 100870, 100900, 100920, 100930, 100980, 101000, 
    101030, 101040, 101040, 101040, 101030, 101030, 101030, 101030, 101040, 
    101030, 101010, 101010, 101010, 101000, 100980, 100940, 100900, 100880, 
    100870, 100800, 100770, 100720, 100680, 100640, 100550, 100440, 100320, 
    100290, 100180, 100110, 99980, 99890, 99810, 99710, 99730, 99680, 99690, 
    99760, 99820, 99890, 99960, 100100, 100160, 100230, 100310, 100370, 
    100460, 100550, 100620, 100690, 100730, 100770, 100830, 100880, 100920, 
    100980, 101050, 101140, 101180, 101210, 101310, 101290, 101370, 101410, 
    101410, 101460, 101560, 101640, 101750, 101850, 101940, 102020, 102070, 
    102100, 102180, 102230, 102280, 102310, 102380, 102370, 102420, 102450, 
    102460, 102500, 102520, 102540, 102540, 102540, 102540, 102560, 102550, 
    102550, 102540, 102560, 102570, 102560, 102560, 102560, 102540, 102540, 
    102530, 102520, 102490, 102480, 102440, 102470, 102470, 102470, 102470, 
    102440, 102400, 102370, 102390, 102380, 102350, 102330, 102330, 102330, 
    102310, 102280, 102260, 102220, 102190, 102200, 102190, 102180, 102140, 
    102110, 102080, 102090, 102090, 102080, 102070, 102060, 102050, 102070, 
    102050, 101990, 102000, 102000, 101980, 101970, 101990, 101970, 101980, 
    101990, 101990, 101990, 102000, 102000, 102020, 102030, 102030, 102030, 
    102070, 102070, 102070, 102060, 102060, 102050, 102040, 102040, 102030, 
    102030, 102020, 102050, 102070, 102070, 102080, 102130, 102150, 102120, 
    102110, 102100, 102100, 102100, 102080, 102080, 102040, 102050, 102070, 
    102070, 102050, 102040, 102050, 102040, 102000, 101990, 102000, 102010, 
    102000, 102000, 102020, 102010, 101990, 101970, 102000, 101980, 101970, 
    101950, 101950, 101940, 101940, 101960, 101980, 101990, 101970, 101950, 
    101940, 101920, 101900, 101910, 101910, 101900, 101920, 101910, 101940, 
    101940, 101940, 101940, 101950, 101880, 101870, 101830, 101820, 101840, 
    101810, 101810, 101820, 101870, 101860, 101870, 101880, 101880, 101830, 
    101830, 101850, 101870, 101900, 101920, 101940, 101960, 101960, 101960, 
    101910, 101920, 101920, 101950, 102000, 102020, 102040, 102030, 102040, 
    102070, 102070, 102070, 102080, 102120, 102120, 102150, 102160, 102180, 
    102210, 102250, 102270, 102250, 102260, 102300, 102270, 102310, 102350, 
    102390, 102440, 102440, 102430, 102460, 102470, 102460, 102470, 102430, 
    102480, 102500, 102510, 102510, 102520, 102510, 102500, 102480, 102460, 
    102460, 102440, 102430, 102390, 102360, 102380, 102340, 102340, 102320, 
    102310, 102290, 102270, 102260, 102220, 102200, 102180, 102160, 102130, 
    102140, 102120, 102080, 102070, 102080, 102080, 102020, 101990, 101960, 
    101950, 101950, 101880, 101870, 101840, 101810, 101770, 101740, 101710, 
    101670, 101660, 101600, 101570, 101560, 101540, 101480, 101470, 101430, 
    101390, 101360, 101370, 101300, 101280, 101230, 101170, 101100, 101030, 
    100990, 100930, 100870, 100820, 100790, 100760, 100750, 100720, 100680, 
    100640, 100630, 100650, 100670, 100690, 100720, 100770, 100820, 100880, 
    100910, 100940, 101020, 101060, 101120, 101200, 101260, 101290, 101330, 
    101390, 101430, 101450, 101480, 101490, 101530, 101560, 101530, 101510, 
    101490, 101410, 101330, 101270, 101280, 101180, 101110, 101080, 101040, 
    101040, 100950, 100880, 100780, 100800, 100760, 100750, 100780, 100780, 
    100810, 100890, 100880, 100900, 100890, 100910, 100910, 100920, 100980, 
    101060, 101150, 101250, 101400, 101480, 101620, 101720, 101800, 101900, 
    102030, 102130, 102200, 102270, 102330, 102460, 102540, 102610, 102640, 
    102710, 102750, 102770, 102830, 102870, 102860, 102920, 102970, 102990, 
    103030, 103060, 103060, 103040, 103050, 103060, 103050, 103020, 103010, 
    102970, 102950, 102940, 102910, 102860, 102820, 102790, 102780, 102740, 
    102740, 102720, 102730, 102710, 102710, 102720, 102730, 102740, 102750, 
    102740, 102730, 102690, 102710, 102680, 102660, 102630, 102600, 102540, 
    102490, 102430, 102360, 102280, 102200, 102120, 102040, 101990, 101930, 
    101880, 101810, 101760, 101700, 101670, 101620, 101560, 101530, 101450, 
    101440, 101410, 101410, 101380, 101400, 101410, 101400, 101400, 101420, 
    101390, 101370, 101320, 101310, 101240, 101210, 101150, 101060, 101000, 
    100950, 100830, 100810, 100680, 100660, 100610, 100590, 100590, 100590, 
    100560, 100570, 100630, 100720, 100850, 100980, 101100, 101240, 101400, 
    101560, 101670, 101790, 101940, 102030, 102140, 102260, 102330, 102420, 
    102490, 102570, 102620, 102670, 102750, 102780, 102830, 102850, 102880, 
    102850, 102820, 102810, 102770, 102770, 102690, 102600, 102510, 102470, 
    102410, 102350, 102270, 102170, 102130, 102020, 101960, 101880, 101810, 
    101710, 101660, 101590, 101550, 101520, 101480, 101460, 101430, 101370, 
    101360, 101370, 101420, 101430, 101440, 101480, 101540, 101610, 101610, 
    101640, 101640, 101730, 101770, 101840, 101880, 101920, 101930, 101940, 
    101950, 101920, 101940, 101910, 101900, 101880, 101840, 101870, 101880, 
    101910, 101930, 101970, 102030, 102080, 102100, 102130, 102190, 102220, 
    102250, 102260, 102260, 102310, 102320, 102340, 102340, 102380, 102350, 
    102340, 102320, 102260, 102290, 102200, 102220, 102240, 102230, 102280, 
    102270, 102280, 102310, 102330, 102340, 102360, 102380, 102390, 102410, 
    102440, 102400, 102430, 102400, 102380, 102390, 102410, 102430, 102410, 
    102410, 102400, 102420, 102390, 102400, 102400, 102430, 102420, 102410, 
    102390, 102380, 102330, 102330, 102320, 102290, 102270, 102240, 102190, 
    102220, 102190, 102190, 102200, 102210, 102190, 102210, 102210, 102180, 
    102150, 102240, 102250, 102250, 102320, 102310, 102350, 102360, 102390, 
    102370, 102400, 102460, 102480, 102480, 102520, 102520, 102530, 102550, 
    102560, 102550, 102580, 102580, 102600, 102610, 102600, 102550, 102550, 
    102520, 102490, 102480, 102440, 102390, 102440, 102460, 102370, 102300, 
    102300, 102260, 102180, 102200, 102160, 102110, 102050, 102030, 102030, 
    101980, 101920, 101910, 101920, 101890, 101880, 101890, 101880, 101810, 
    101750, 101680, 101650, 101580, 101540, 101480, 101400, 101320, 101270, 
    101210, 101150, 101080, 101020, 100930, 100840, 100800, 100750, 100680, 
    100630, 100600, 100580, 100530, 100490, 100460, 100400, 100360, 100330, 
    100290, 100250, 100200, 100130, 100090, 100070, 100070, 100030, 99990, 
    99950, 99920, 99920, 99910, 99910, 99890, 99870, 99880, 99880, 99890, 
    99910, 99930, 99940, 99940, 99960, 99970, 99970, 99970, 99960, 100000, 
    100000, 100020, 100060, 100080, 100090, 100120, 100140, 100160, 100150, 
    100180, 100170, 100210, 100250, 100300, 100360, 100420, 100450, 100450, 
    100470, 100500, 100530, 100570, 100590, 100600, 100650, 100690, 100720, 
    100750, 100790, 100810, 100850, 100850, 100870, 100910, 100930, 100950, 
    100950, 100980, 101000, 101040, 101060, 101100, 101130, 101120, 101090, 
    101110, 101140, 101140, 101160, 101190, 101190, 101230, 101240, 101230, 
    101230, 101250, 101290, 101290, 101290, 101290, 101300, 101310, 101310, 
    101310, 101310, 101310, 101340, 101340, 101350, 101360, 101350, 101340, 
    101340, 101360, 101380, 101410, 101410, 101410, 101410, 101420, 101420, 
    101420, 101430, 101430, 101440, 101470, 101490, 101510, 101540, 101570, 
    101580, 101590, 101610, 101610, 101620, 101620, 101610, 101620, 101650, 
    101650, 101640, 101630, 101620, 101630, 101620, 101630, 101630, 101620, 
    101610, 101600, 101600, 101600, 101580, 101560, 101520, 101490, 101470, 
    101420, 101430, 101420, 101420, 101410, 101400, 101430, 101440, 101440, 
    101460, 101480, 101490, 101490, 101480, 101500, 101490, 101480, 101480, 
    101490, 101480, 101460, 101440, 101440, 101450, 101460, 101470, 101450, 
    101480, 101510, 101530, 101550, 101580, 101570, 101600, 101610, 101600, 
    101610, 101640, 101630, 101620, 101620, 101650, 101640, 101630, 101630, 
    101630, 101620, 101580, 101620, 101630, 101610, 101620, 101630, 101650, 
    101630, 101650, 101650, 101640, 101640, 101660, 101680, 101680, 101690, 
    101720, 101740, 101770, 101810, 101810, 101820, 101840, 101840, 101850, 
    101890, 101920, 101920, 101920, 101940, 101930, 101930, 101940, 101950, 
    101950, 101940, 101980, 101980, 102000, 102020, 102030, 102040, 102050, 
    102060, 102050, 102030, 102030, 102030, 102030, 102010, 102000, 102000, 
    101990, 101970, 101980, 101970, 101970, 101960, 101960, 101960, 101940, 
    101940, 101940, 101940, 101940, 101920, 101940, 101940, 101920, 101900, 
    101920, 101890, 101860, 101750, 101780, 101840, 101890, 101920, 101950, 
    101970, 101970, 101970, 101910, 101940, 101910, 101890, 101850, 101850, 
    101870, 101900, 101920, 101940, 101960, 101950, 101920, 101900, 101900, 
    101890, 101870, 101880, 101890, 101850, 101800, 101800, 101740, 101690, 
    101660, 101630, 101590, 101540, 101510, 101480, 101470, 101440, 101450, 
    101440, 101430, 101430, 101450, 101440, 101440, 101430, 101410, 101440, 
    101460, 101480, 101490, 101500, 101520, 101550, 101550, 101550, 101550, 
    101540, 101520, 101520, 101560, 101600, 101630, 101650, 101680, 101700, 
    101700, 101720, 101750, 101760, 101780, 101810, 101840, 101870, 101880, 
    101900, 101910, 101920, 101920, 101940, 101950, 101960, 101990, 102000, 
    102020, 102040, 102050, 102060, 102040, 102070, 102070, 102070, 102050, 
    102040, 102030, 102030, 102040, 102050, 102060, 102050, 102030, 102000, 
    102000, 102000, 101990, 102000, 101950, 101950, 101940, 101930, 101910, 
    101890, 101860, 101840, 101840, 101820, 101810, 101800, 101780, 101750, 
    101730, 101720, 101730, 101730, 101680, 101650, 101610, 101630, 101640, 
    101630, 101600, 101620, 101600, 101640, 101630, 101670, 101680, 101690, 
    101710, 101740, 101720, 101750, 101770, 101780, 101820, 101830, 101830, 
    101850, 101860, 101870, 101880, 101880, 101880, 101900, 101880, 101900, 
    101910, 101940, 101950, 101940, 101940, 101960, 101970, 101950, 101990, 
    101980, 101990, 101980, 101990, 101980, 101960, 101950, 101930, 101890, 
    101870, 101830, 101820, 101770, 101770, 101680, 101640, 101630, 101570, 
    101460, 101340, 101270, 101150, 101100, 101030, 100980, 100910, 100840, 
    100820, 100740, 100670, 100600, 100560, 100510, 100450, 100430, 100440, 
    100430, 100430, 100440, 100440, 100470, 100460, 100420, 100400, 100380, 
    100330, 100350, 100370, 100390, 100430, 100420, 100450, 100460, 100460, 
    100480, 100540, 100550, 100580, 100630, 100670, 100690, 100690, 100730, 
    100760, 100780, 100820, 100840, 100860, 100870, 100860, 100790, 100760, 
    100750, 100740, 100710, 100700, 100720, 100680, 100630, 100630, 100620, 
    100590, 100590, 100600, 100600, 100560, 100570, 100550, 100560, 100560, 
    100590, 100590, 100600, 100580, 100570, 100570, 100550, 100540, 100570, 
    100570, 100560, 100540, 100550, 100520, 100510, 100500, 100450, 100440, 
    100400, 100370, 100320, 100300, 100240, 100240, 100210, 100180, 100140, 
    100060, 100000, 99960, 99910, 99860, 99790, 99720, 99670, 99600, 99550, 
    99490, 99440, 99370, 99310, 99240, 99170, 99140, 99090, 98980, 99000, 
    98970, 98900, 98890, 98840, 98800, 98790, 98750, 98610, 98550, 98570, 
    98570, 98530, 98480, 98410, 98380, 98350, 98300, 98250, 98230, 98180, 
    98120, 98180, 98120, 98170, 98160, 98060, 98040, 98010, 98020, 97980, 
    98050, 98130, 98200, 98260, 98340, 98400, 98430, 98460, 98490, 98510, 
    98580, 98560, 98540, 98590, 98610, 98660, 98650, 98660, 98700, 98700, 
    98670, 98670, 98720, 98740, 98760, 98830, 98860, 98860, 98900, 98910, 
    98920, 98970, 98980, 98970, 98970, 98970, 99010, 99020, 99040, 99090, 
    99100, 99090, 99080, 99050, 98970, 98920, 98850, 98810, 98810, 98790, 
    98720, 98780, 98770, 98840, 98860, 98890, 98860, 98890, 98890, 98910, 
    98910, 98930, 98910, 98910, 98940, 98930, 98940, 98980, 98990, 98990, 
    99010, 99030, 99030, 99050, 99070, 99070, 99100, 99110, 99130, 99140, 
    99160, 99170, 99200, 99210, 99230, 99250, 99280, 99300, 99330, 99360, 
    99380, 99400, 99400, 99420, 99400, 99390, 99400, 99410, 99400, 99400, 
    99400, 99380, 99380, 99380, 99340, 99320, 99310, 99290, 99270, 99240, 
    99220, 99200, 99160, 99140, 99120, 99110, 99070, 99030, 98980, 98920, 
    98840, 98790, 98710, 98700, 98660, 98630, 98580, 98570, 98560, 98550, 
    98560, 98560, 98510, 98510, 98540, 98490, 98520, 98490, 98480, 98400, 
    98360, 98330, 98320, 98340, 98380, 98390, 98420, 98440, 98460, 98510, 
    98560, 98590, 98640, 98710, 98860, 98860, 98960, 99060, 99150, 99240, 
    99290, 99340, 99360, 99380, 99430, 99490, 99490, 99500, 99510, 99520, 
    99520, 99530, 99540, 99620, 99750, 99780, 99800, 99850, 99880, 99940, 
    99990, 100050, 100070, 100120, 100190, 100230, 100300, 100330, 100380, 
    100430, 100450, 100540, 100590, 100650, 100680, 100720, 100760, 100810, 
    100850, 100910, 100930, 100970, 101010, 101050, 101090, 101100, 101140, 
    101180, 101220, 101270, 101290, 101330, 101370, 101390, 101420, 101450, 
    101470, 101480, 101520, 101540, 101560, 101620, 101650, 101670, 101700, 
    101710, 101730, 101770, 101800, 101800, 101840, 101870, 101920, 101970, 
    101970, 102020, 102080, 102110, 102140, 102190, 102210, 102250, 102260, 
    102300, 102330, 102370, 102380, 102400, 102400, 102410, 102400, 102410, 
    102410, 102400, 102420, 102370, 102370, 102370, 102340, 102310, 102290, 
    102240, 102200, 102160, 102120, 102110, 102060, 102010, 101980, 101950, 
    101900, 101810, 101760, 101680, 101620, 101580, 101580, 101560, 101520, 
    101510, 101490, 101470, 101460, 101450, 101430, 101400, 101370, 101310, 
    101280, 101220, 101130, 101060, 100990, 101020, 101030, 101050, 101120, 
    101180, 101080, 101070, 101180, 101220, 101250, 101260, 101230, 101150, 
    101170, 101130, 101160, 101300, 101360, 101320, 101300, 101250, 101210, 
    101140, 101080, 101110, 101140, 101070, 101030, 101010, 100950, 100850, 
    100790, 100730, 100770, 100740, 100750, 100760, 100760, 100760, 100740, 
    100690, 100620, 100580, 100550, 100620, 100550, 100440, 100400, 100280, 
    100400, 100470, 100460, 100440, 100440, 100400, 100330, 100200, 100200, 
    100230, 100250, 100300, 100320, 100330, 100370, 100360, 100360, 100360, 
    100330, 100310, 100300, 100230, 100160, 100140, 100150, 100190, 100210, 
    100250, 100290, 100340, 100370, 100410, 100440, 100460, 100530, 100520, 
    100550, 100560, 100560, 100590, 100600, 100590, 100580, 100540, 100540, 
    100580, 100590, 100610, 100630, 100640, 100620, 100590, 100620, 100640, 
    100660, 100670, 100710, 100750, 100780, 100810, 100820, 100860, 100890, 
    100920, 100930, 100990, 101010, 101050, 101100, 101180, 101200, 101190, 
    101170, 101200, 101200, 101190, 101220, 101270, 101210, 101230, 101300, 
    101360, 101370, 101410, 101470, 101530, 101540, 101590, 101640, 101630, 
    101620, 101590, 101550, 101690, 101710, 101700, 101710, 101730, 101740, 
    101730, 101730, 101720, 101740, 101760, 101780, 101790, 101770, 101830, 
    101840, 101840, 101830, 101870, 101840, 101910, 101860, 101850, 101890, 
    101910, 101910, 101920, 101910, 101890, 101870, 101850, 101840, 101840, 
    101820, 101790, 101770, 101720, 101700, 101760, 101770, 101760, 101760, 
    101640, 101770, 101830, 101910, 101920, 101910, 101930, 101970, 101990, 
    102030, 102050, 102050, 102070, 102070, 102110, 102110, 102100, 102120, 
    102140, 102150, 102220, 102250, 102260, 102270, 102230, 102310, 102320, 
    102320, 102330, 102330, 102250, 102320, 102340, 102380, 102380, 102400, 
    102410, 102430, 102440, 102440, 102460, 102470, 102490, 102510, 102550, 
    102610, 102650, 102670, 102690, 102710, 102740, 102760, 102770, 102780, 
    102790, 102830, 102870, 102870, 102900, 102900, 102900, 103000, 103030, 
    103010, 103030, 103080, 103100, 103140, 103250, 103290, 103220, 103420, 
    103400, 103390, 103460, 103480, 103510, 103530, 103550, 103600, 103650, 
    103680, 103750, 103750, 103780, 103770, 103780, 103790, 103830, 103830, 
    103850, 103840, 103830, 103860, 103890, 103990, 103980, 103930, 103960, 
    103980, 104010, 103980, 104020, 103990, 104020, 104030, 103980, 103970, 
    104050, 104060, 104110, 104130, 104110, 104100, 104090, 104090, 104110, 
    104140, 104160, 104150, 104160, 104120, 104140, 104160, 104160, 104160, 
    104160, 104170, 104190, 104170, 104180, 104200, 104200, 104200, 104190, 
    104220, 104210, 104180, 104160, 104150, 104140, 104140, 104110, 104060, 
    104040, 103980, 103960, 103940, 103900, 103880, 103850, 103800, 103770, 
    103730, 103690, 103670, 103620, 103560, 103490, 103470, 103440, 103410, 
    103370, 103350, 103330, 103320, 103280, 103240, 103200, 103160, 103120, 
    103090, 103070, 103060, 103020, 102930, 102880, 102840, 102810, 102740, 
    102690, 102640, 102600, 102540, 102470, 102420, 102360, 102310, 102260, 
    102240, 102170, 102120, 102060, 101980, 101890, 101830, 101770, 101710, 
    101650, 101580, 101520, 101440, 101370, 101300, 101220, 101160, 101070, 
    100970, 100900, 100830, 100750, 100680, 100620, 100550, 100500, 100440, 
    100350, 100280, 100250, 100250, 100230, 100230, 100230, 100240, 100240, 
    100240, 100230, 100250, 100230, 100210, 100170, 100160, 100160, 100180, 
    100220, 100220, 100220, 100230, 100240, 100180, 100190, 100220, 100250, 
    100270, 100350, 100420, 100440, 100450, 100460, 100460, 100520, 100520, 
    100500, 100540, 100550, 100520, 100570, 100570, 100590, 100680, 100910, 
    100960, 100990, 101030, 101050, 101070, 101120, 101150, 101140, 101160, 
    101200, 101200, 101180, 101160, 101230, 101220, 101210, 101180, 101170, 
    101150, 101110, 101130, 101130, 101110, 101130, 101180, 101160, 101160, 
    101150, 101160, 101180, 101210, 101230, 101230, 101280, 101280, 101300, 
    101310, 101320, 101310, 101300, 101230, 101240, 101250, 101230, 101220, 
    101200, 101190, 101190, 101190, 101200, 101220, 101190, 101160, 101130, 
    101140, 101120, 101100, 101100, 101090, 101080, 101060, 101040, 100970, 
    100910, 100820, 100710, 100650, 100520, 100340, 100160, 100000, 99790, 
    99590, 99380, 99240, 99230, 99260, 99250, 99240, 99220, 99190, 99220, 
    99240, 99290, 99320, 99380, 99410, 99440, 99450, 99460, 99480, 99460, 
    99450, 99420, 99390, 99340, 99300, 99290, 99280, 99220, 99180, 99150, 
    99140, 99140, 99160, 99170, 99200, 99200, 99200, 99190, 99220, 99240, 
    99290, 99310, 99340, 99340, 99310, 99330, 99340, 99360, 99380, 99300, 
    99320, 99310, 99360, 99430, 99500, 99570, 99630, 99680, 99750, 99770, 
    99810, 99860, 99870, 99900, 99880, 99870, 99850, 99930, 99930, 99960, 
    99980, 100040, 100110, 100110, 100210, 100250, 100310, 100340, 100350, 
    100390, 100410, 100440, 100450, 100440, 100460, 100450, 100460, 100430, 
    100430, 100440, 100420, 100420, 100460, 100480, 100540, 100580, 100530, 
    100590, 100590, 100630, 100650, 100610, 100700, 100670, 100680, 100690, 
    100710, 100690, 100580, 100640, 100600, 100730, 100740, 100800, 100920, 
    100930, 100890, 100990, 101040, 101070, 101110, 101130, 101150, 101200, 
    101260, 101280, 101270, 101330, 101350, 101360, 101440, 101440, 101440, 
    101420, 101480, 101440, 101500, 101520, 101500, 101520, 101490, 101490, 
    101530, 101520, 101460, 101430, 101470, 101430, 101580, 101660, 101700, 
    101710, 101700, 101740, 101790, 101810, 101830, 101850, 101870, 101890, 
    101910, 101920, 101940, 101910, 101910, 101900, 101990, 102050, 102060, 
    102120, 102140, 102150, 102140, 102180, 102230, 102230, 102280, 102250, 
    102270, 102280, 102320, 102330, 102350, 102360, 102360, 102350, 102340, 
    102330, 102310, 102310, 102290, 102290, 102320, 102290, 102260, 102220, 
    102160, 102140, 102130, 102120, 102110, 102070, 102000, 102020, 101990, 
    101970, 101940, 101890, 101870, 101870, 101840, 101810, 101790, 101760, 
    101750, 101730, 101730, 101720, 101690, 101620, 101620, 101620, 101610, 
    101620, 101650, 101660, 101660, 101670, 101660, 101650, 101650, 101600, 
    101630, 101570, 101560, 101590, 101600, 101570, 101570, 101600, 101610, 
    101580, 101560, 101580, 101560, 101550, 101520, 101520, 101470, 101440, 
    101380, 101350, 101280, 101280, 101230, 101200, 101120, 101070, 101040, 
    101010, 100970, 100910, 100830, 100800, 100780, 100670, 100570, 100510, 
    100420, 100330, 100240, 100060, 100190, 99880, 99820, 99770, 99560, 
    99550, 99520, 99470, 99400, 99460, 99350, 99310, 99300, 99290, 99340, 
    99360, 99440, 99480, 99520, 99550, 99580, 99600, 99640, 99680, 99740, 
    99760, 99780, 99780, 99650, 99590, 99600, 99600, 99590, 99610, 99640, 
    99600, 99770, 99940, 99950, 99940, 99970, 99970, 99970, 99960, 99940, 
    99920, 99890, 99860, 99830, 99840, 99880, 99880, 99860, 99820, 99840, 
    99860, 99900, 100090, 100120, 100150, 100140, 100160, 100210, 100190, 
    100040, 100020, 100150, 100170, 100200, 100230, 100230, 100000, 99950, 
    99930, 99980, 100040, 100120, 100200, 100170, 100200, 100250, 100280, 
    100270, 100300, 100300, 100310, 100300, 100320, 100350, 100370, 100340, 
    100330, 100330, 100350, 100340, 100330, 100270, 100280, 100240, 100230, 
    100240, 100250, 100230, 100210, 100220, 100220, 100160, 100190, 100160, 
    100150, 100160, 100120, 100100, 100040, 100030, 99980, 99940, 99880, 
    99890, 99920, 99940, 99970, 100010, 99990, 100020, 100040, 100050, 
    100070, 100080, 100080, 100070, 100080, 100080, 100110, 100140, 100150, 
    100160, 100190, 100220, 100240, 100270, 100340, 100370, 100380, 100410, 
    100420, 100450, 100470, 100480, 100490, 100530, 100500, 100490, 100470, 
    100420, 100390, 100340, 100310, 100300, 100240, 100200, 100180, 100170, 
    100060, 99910, 99770, 99620, 99400, 99250, 99050, 98860, 98650, 98450, 
    98250, 98000, 97720, 97460, 97180, 96900, 96630, 96500, 96460, 96440, 
    96410, 96390, 96360, 96270, 96200, 96130, 96110, 96110, 96140, 96170, 
    96160, 96160, 96140, 96150, 96130, 96210, 96300, 96380, 96480, 96580, 
    96650, 96720, 96790, 96850, 96960, 97090, 97220, 97300, 97370, 97420, 
    97470, 97480, 97570, 97600, 97730, 97860, 97940, 98060, 98150, 98230, 
    98310, 98420, 98510, 98600, 98690, 98700, 98780, 98820, 98810, 98820, 
    98680, 98710, 98740, 98770, 98820, 98870, 98840, 98850, 98900, 98980, 
    99010, 99030, 99020, 99100, 99110, 99150, 99130, 99170, 99250, 99320, 
    99410, 99480, 99540, 99580, 99660, 99710, 99760, 99840, 99890, 99910, 
    99930, 99960, 99980, 100000, 100040, 100070, 100120, 100160, 100180, 
    100210, 100210, 100240, 100240, 100240, 100210, 100270, 100280, 100320, 
    100320, 100300, 100240, 100300, 100290, 100300, 100260, 100260, 100300, 
    100310, 100330, 100400, 100550, 100620, 100660, 100670, 100730, 100830, 
    100930, 100980, 101050, 101130, 101180, 101180, 101220, 101250, 101330, 
    101400, 101410, 101370, 101390, 101450, 101450, 101480, 101490, 101560, 
    101510, 101490, 101560, 101530, 101500, 101480, 101430, 101350, 101210, 
    101040, 100810, 100680, 100660, 100480, 100360, 100290, 100190, 100130, 
    100040, 100020, 99960, 100030, 100070, 100050, 100090, 100150, 100220, 
    100250, 100250, 100290, 100260, 100230, 100220, 100190, 100220, 100210, 
    100200, 100100, 99990, 99960, 99920, 99850, 99740, 99590, 99390, 99250, 
    99050, 98840, 98580, 98360, 98130, 97960, 97900, 97830, 97790, 97780, 
    97770, 97810, 97850, 97920, 97970, 98000, 98020, 98070, 98140, 98190, 
    98290, 98320, 98380, 98430, 98510, 98560, 98590, 98600, 98660, 98700, 
    98760, 98790, 98810, 98780, 98760, 98860, 98830, 98790, 98770, 98760, 
    98740, 98840, 98920, 98940, 98990, 99030, 99050, 99130, 99260, 99400, 
    99500, 99520, 99740, 99800, 99930, 100000, 100010, 100090, 100260, 
    100380, 100450, 100520, 100480, 100540, 100570, 100630, 100650, 100710, 
    100730, 100690, 100730, 100770, 100750, 100780, 100750, 100730, 100730, 
    100770, 100780, 100790, 100760, 100760, 100760, 100770, 100780, 100770, 
    100780, 100820, 100810, 100790, 100810, 100850, 100820, 100810, 100830, 
    100820, 100840, 100810, 100840, 100850, 100830, 100830, 100840, 100810, 
    100790, 100780, 100770, 100750, 100750, 100730, 100720, 100700, 100630, 
    100620, 100620, 100600, 100590, 100570, 100520, 100500, 100490, 100490, 
    100480, 100470, 100460, 100420, 100400, 100380, 100340, 100320, 100290, 
    100270, 100240, 100240, 100240, 100240, 100230, 100220, 100200, 100210, 
    100230, 100220, 100220, 100250, 100280, 100290, 100290, 100260, 100250, 
    100210, 100200, 100180, 100200, 100180, 100180, 100220, 100220, 100250, 
    100270, 100290, 100300, 100310, 100310, 100330, 100350, 100390, 100430, 
    100430, 100440, 100460, 100550, 100510, 100530, 100590, 100610, 100610, 
    100610, 100640, 100670, 100680, 100710, 100730, 100750, 100800, 100810, 
    100800, 100780, 100860, 100830, 100880, 100900, 100900, 100920, 100930, 
    100970, 100970, 101000, 101010, 101020, 101010, 101010, 100990, 101020, 
    101090, 101080, 101100, 101090, 101120, 101150, 101110, 101100, 101090, 
    101120, 101090, 101090, 101100, 101110, 101100, 101090, 101050, 101020, 
    100980, 100960, 100860, 100740, 100550, 100500, 100450, 100360, 100390, 
    100360, 100390, 100420, 100450, 100460, 100500, 100510, 100490, 100500, 
    100500, 100490, 100480, 100480, 100500, 100500, 100500, 100480, 100450, 
    100370, 100350, 100330, 100310, 100310, 100220, 100220, 100200, 100170, 
    100180, 100140, 100120, 100080, 100020, 99980, 99940, 99920, 99970, 
    100060, 100070, 100110, 100150, 100210, 100250, 100310, 100380, 100430, 
    100500, 100560, 100610, 100670, 100730, 100780, 100810, 100860, 100890, 
    100930, 100930, 100980, 101040, 101060, 101060, 101070, 101090, 101120, 
    101120, 101150, 101150, 101160, 101170, 101200, 101220, 101260, 101310, 
    101290, 101310, 101300, 101360, 101380, 101370, 101390, 101400, 101420, 
    101420, 101430, 101440, 101440, 101430, 101440, 101470, 101480, 101460, 
    101460, 101460, 101440, 101440, 101440, 101460, 101450, 101440, 101400, 
    101400, 101380, 101330, 101320, 101320, 101290, 101270, 101260, 101270, 
    101260, 101250, 101230, 101180, 101170, 101130, 101110, 101090, 101070, 
    101050, 101060, 101030, 101020, 101050, 101020, 100990, 100980, 100950, 
    100920, 100930, 100910, 100870, 100830, 100790, 100800, 100770, 100750, 
    100730, 100710, 100710, 100650, 100630, 100600, 100580, 100590, 100570, 
    100540, 100460, 100380, 100320, 100330, 100330, 100400, 100380, 100430, 
    100480, 100500, 100530, 100550, 100620, 100580, 100570, 100500, 100420, 
    100350, 100210, 100080, 99970, 99860, 99720, 99610, 99460, 99260, 99140, 
    98980, 98820, 98700, 98610, 98550, 98510, 98390, 98330, 98290, 98240, 
    98200, 98220, 98280, 98290, 98340, 98400, 98530, 98640, 98720, 98840, 
    98950, 99030, 99110, 99150, 99230, 99250, 99250, 99270, 99310, 99350, 
    99390, 99390, 99440, 99480, 99500, 99500, 99500, 99530, 99510, 99510, 
    99470, 99480, 99490, 99490, 99490, 99540, 99580, 99620, 99590, 99610, 
    99610, 99670, 99680, 99700, 99750, 99770, 99810, 99840, 99850, 99860, 
    99870, 99870, 99880, 99920, 99940, 99970, 100010, 100040, 100090, 100150, 
    100190, 100150, 100180, 100220, 100230, 100270, 100280, 100280, 100340, 
    100450, 100530, 100610, 100660, 100760, 100780, 100850, 100890, 100970, 
    101050, 101110, 101170, 101230, 101290, 101350, 101370, 101370, 101420, 
    101460, 101470, 101550, 101570, 101630, 101680, 101710, 101670, 101720, 
    101720, 101710, 101710, 101720, 101770, 101810, 101840, 101880, 101910, 
    101920, 101890, 101860, 101860, 101790, 101770, 101720, 101650, 101640, 
    101620, 101650, 101640, 101710, 101770, 101840, 101890, 101910, 101940, 
    101950, 101980, 102000, 102040, 102080, 102120, 102170, 102210, 102250, 
    102250, 102260, 102280, 102310, 102280, 102240, 102220, 102200, 102200, 
    102220, 102200, 102170, 102080, 102010, 101930, 101870, 101790, 101730, 
    101640, 101560, 101450, 101410, 101470, 101400, 101360, 101320, 101290, 
    101250, 101250, 101200, 101120, 100960, 100850, 100840, 100820, 100790, 
    100870, 100990, 101190, 101360, 101440, 101530, 101610, 101670, 101760, 
    101800, 101830, 101850, 101840, 101820, 101850, 101860, 101890, 101940, 
    101990, 101980, 101980, 101990, 101980, 101980, 101980, 101980, 101990, 
    101980, 101950, 101960, 101970, 101960, 101980, 102010, 102030, 102040, 
    102050, 102050, 102050, 102040, 102050, 102050, 102050, 102050, 102070, 
    102070, 102100, 102090, 102110, 102090, 102120, 102140, 102140, 102160, 
    102160, 102170, 102170, 102170, 102170, 102190, 102160, 102180, 102160, 
    102160, 102140, 102140, 102110, 102090, 102070, 102060, 102030, 101990, 
    101940, 101910, 101850, 101810, 101810, 101780, 101730, 101690, 101650, 
    101630, 101590, 101530, 101490, 101500, 101480, 101460, 101430, 101370, 
    101360, 101360, 101350, 101330, 101300, 101270, 101240, 101210, 101240, 
    101200, 101170, 101160, 101120, 101140, 101130, 101110, 101120, 101080, 
    101070, 101060, 101030, 101020, 101020, 101010, 101020, 101010, 101030, 
    100980, 100980, 100900, 100830, 100840, 100850, 100740, 100720, 100670, 
    100620, 100580, 100540, 100510, 100460, 100440, 100380, 100340, 100370, 
    100390, 100400, 100410, 100350, 100390, 100430, 100510, 100540, 100610, 
    100650, 100680, 100700, 100680, 100700, 100730, 100730, 100740, 100750, 
    100770, 100800, 100830, 100830, 100850, 100940, 101000, 100980, 101000, 
    101020, 101000, 101000, 101000, 101010, 101000, 100970, 100940, 100930, 
    100910, 100880, 100850, 100810, 100830, 100860, 100890, 100870, 100910, 
    100950, 100970, 101010, 101040, 101060, 101070, 101080, 101100, 101120, 
    101170, 101210, 101240, 101270, 101310, 101300, 101330, 101350, 101380, 
    101380, 101410, 101490, 101520, 101540, 101580, 101610, 101610, 101640, 
    101680, 101680, 101680, 101690, 101720, 101740, 101790, 101800, 101810, 
    101820, 101830, 101840, 101850, 101860, 101860, 101850, 101860, 101880, 
    101930, 101940, 101950, 101960, 101980, 101960, 101980, 101990, 101970, 
    101970, 101980, 101990, 102030, 102010, 102060, 102020, 102010, 102070, 
    102070, 102070, 102070, 102070, 102120, 102160, 102200, 102230, 102250, 
    102290, 102320, 102330, 102370, 102380, 102400, 102450, 102490, 102520, 
    102560, 102600, 102630, 102630, 102650, 102690, 102710, 102700, 102700, 
    102720, 102750, 102780, 102790, 102780, 102770, 102750, 102740, 102720, 
    102680, 102640, 102620, 102570, 102530, 102500, 102480, 102450, 102390, 
    102360, 102280, 102220, 102180, 102100, 102030, 102000, 101970, 101960, 
    101920, 101880, 101830, 101780, 101690, 101610, 101580, 101550, 101510, 
    101470, 101460, 101430, 101430, 101450, 101420, 101420, 101430, 101430, 
    101420, 101420, 101440, 101430, 101430, 101440, 101470, 101460, 101460, 
    101480, 101410, 101430, 101430, 101400, 101360, 101330, 101300, 101290, 
    101210, 101180, 101110, 101060, 101020, 100940, 100870, 100770, 100680, 
    100540, 100420, 100380, 100310, 100240, 100110, 100000, 99940, 99820, 
    99690, 99560, 99470, 99400, 99420, 99360, 99200, 99010, 98860, 98670, 
    98320, 98080, 97830, 97380, 97170, 97040, 97030, 97050, 97110, 97160, 
    97210, 97320, 97420, 97460, 97610, 97750, 97910, 98060, 98240, 98430, 
    98540, 98710, 98840, 98950, 99100, 99210, 99310, 99420, 99550, 99750, 
    99900, 100120, 100270, 100430, 100580, 100640, 100730, 100760, 100800, 
    100850, 100850, 100770, 100680, 100700, 100730, 100830, 100910, 100920, 
    100900, 100900, 100910, 100870, 100820, 100770, 100600, 100400, 100230, 
    100070, 99950, 99620, 99400, 99300, 99150, 99020, 98890, 98780, 98720, 
    98710, 98700, 98680, 98650, 98620, 98640, 98640, 98600, 98620, 98600, 
    98590, 98590, 98610, 98630, 98680, 98720, 98730, 98760, 98810, 98830, 
    98840, 98840, 98900, 98970, 98990, 99040, 99110, 99160, 99200, 99270, 
    99330, 99400, 99450, 99480, 99520, 99560, 99620, 99670, 99700, 99740, 
    99730, 99780, 99810, 99830, 99840, 99900, 99960, 99980, 100040, 100100, 
    100130, 100150, 100130, 100150, 100120, 100130, 100130, 100080, 100090, 
    100080, 100120, 100100, 100040, 99970, 99920, 99840, 99760, 99660, 99550, 
    99450, 99370, 99300, 99200, 99130, 98990, 98930, 98800, 98820, 98960, 
    99120, 99240, 99380, 99420, 99520, 99590, 99650, 99670, 99720, 99740, 
    99760, 99770, 99780, 99810, 99870, 99940, 100020, 100090, 100180, 100250, 
    100340, 100410, 100470, 100510, 100570, 100620, 100640, 100680, 100720, 
    100750, 100820, 100860, 100900, 100900, 100920, 100950, 100970, 101000, 
    101020, 101050, 101070, 101120, 101160, 101170, 101190, 101210, 101220, 
    101250, 101260, 101280, 101260, 101270, 101280, 101310, 101330, 101320, 
    101320, 101290, 101290, 101260, 101270, 101280, 101290, 101300, 101320, 
    101340, 101370, 101380, 101400, 101410, 101420, 101440, 101440, 101450, 
    101450, 101470, 101500, 101520, 101550, 101570, 101570, 101580, 101570, 
    101580, 101580, 101580, 101590, 101600, 101590, 101580, 101580, 101590, 
    101600, 101600, 101590, 101590, 101590, 101560, 101590, 101610, 101610, 
    101630, 101670, 101700, 101730, 101740, 101760, 101790, 101790, 101830, 
    101860, 101860, 101890, 101930, 101970, 101990, 102000, 102020, 102050, 
    102050, 102060, 102060, 102050, 102060, 102070, 102100, 102130, 102130, 
    102150, 102160, 102170, 102190, 102210, 102200, 102230, 102250, 102280, 
    102340, 102410, 102440, 102450, 102480, 102540, 102630, 102680, 102730, 
    102730, 102760, 102790, 102850, 102890, 102930, 102990, 103010, 103030, 
    103070, 103120, 103160, 103160, 103180, 103190, 103220, 103250, 103260, 
    103270, 103270, 103280, 103290, 103280, 103270, 103230, 103210, 103200, 
    103190, 103210, 103210, 103200, 103210, 103190, 103200, 103200, 103180, 
    103150, 103140, 103120, 103110, 103110, 103110, 103090, 103060, 103050, 
    103030, 103010, 103000, 102990, 102990, 102970, 102970, 103000, 103030, 
    103040, 103050, 103040, 103050, 103060, 103050, 103020, 103050, 103060, 
    103070, 103070, 103100, 103100, 103110, 103130, 103170, 103200, 103180, 
    103170, 103180, 103250, 103300, 103350, 103390, 103420, 103460, 103470, 
    103470, 103490, 103510, 103520, 103520, 103530, 103510, 103500, 103560, 
    103560, 103510, 103500, 103490, 103490, 103490, 103460, 103440, 103410, 
    103410, 103430, 103460, 103450, 103440, 103460, 103490, 103480, 103510, 
    103520, 103480, 103460, 103490, 103520, 103550, 103580, 103580, 103670, 
    103640, 103660, 103670, 103670, 103670, 103700, 103720, 103750, 103800, 
    103840, 103860, 103900, 103930, 103940, 103950, 104000, 104010, 104040, 
    104060, 104080, 104110, 104130, 104130, 104130, 104130, 104160, 104140, 
    104110, 104070, 104070, 104040, 104030, 104040, 104020, 103970, 103940, 
    103920, 103910, 103910, 103870, 103810, 103760, 103770, 103770, 103760, 
    103790, 103740, 103720, 103730, 103770, 103750, 103800, 103860, 103870, 
    103910, 103970, 104020, 104110, 104170, 104240, 104270, 104300, 104320, 
    104340, 104350, 104350, 104350, 104330, 104300, 104300, 104260, 104220, 
    104190, 104160, 104120, 104090, 104060, 104000, 103990, 103940, 103940, 
    103900, 103850, 103740, 103700, 103730, 103690, 103670, 103560, 103600, 
    103540, 103480, 103400, 103410, 103350, 103320, 103270, 103250, 103170, 
    103160, 103130, 103120, 103160, 103160, 103180, 103200, 103160, 103070, 
    102970, 103030, 102910, 102840, 102680, 102590, 102440, 102320, 102190, 
    102110, 102060, 101970, 101920, 101810, 101720, 101650, 101570, 101530, 
    101490, 101460, 101460, 101380, 101290, 101270, 101200, 101190, 101190, 
    101200, 101180, 101180, 101240, 101250, 101290, 101350, 101380, 101430, 
    101480, 101540, 101600, 101600, 101630, 101660, 101720, 101810, 101940, 
    102000, 102090, 102160, 102260, 102330, 102430, 102500, 102550, 102570, 
    102600, 102650, 102680, 102690, 102720, 102730, 102740, 102760, 102780, 
    102740, 102700, 102670, 102660, 102620, 102600, 102610, 102580, 102550, 
    102470, 102380, 102350, 102320, 102300, 102320, 102240, 102190, 102130, 
    102130, 102110, 102070, 102090, 102090, 102060, 102000, 102010, 102000, 
    101900, 101970, 101950, 102000, 102020, 102080, 102090, 102140, 102110, 
    102130, 102160, 102170, 102220, 102260, 102310, 102350, 102400, 102440, 
    102470, 102510, 102510, 102530, 102550, 102580, 102640, 102700, 102720, 
    102770, 102800, 102790, 102830, 102870, 102930, 102960, 102990, 103030, 
    103070, 103080, 103100, 103130, 103110, 103130, 103140, 103150, 103160, 
    103170, 103170, 103200, 103200, 103200, 103270, 103210, 103210, 103130, 
    103110, 103100, 103180, 103330, 103270, 103220, 103200, 103260, 103290, 
    103300, 103250, 103230, 103200, 103170, 103170, 103150, 103130, 103130, 
    103110, 103110, 103100, 103100, 103050, 103050, 103040, 103030, 103020, 
    103020, 103040, 103040, 103020, 103040, 103050, 103090, 103080, 103080, 
    103070, 103070, 103060, 103060, 103060, 103040, 103050, 103070, 103090, 
    103100, 103100, 103070, 103070, 103070, 103070, 103070, 103060, 103060, 
    103070, 103080, 103080, 103060, 103040, 103050, 103030, 103030, 103020, 
    103030, 103010, 103000, 103000, 103010, 103020, 103040, 103020, 103030, 
    103040, 103050, 103040, 103050, 103030, 103030, 103030, 103070, 103070, 
    103070, 103070, 103070, 103050, 103060, 103060, 103060, 103060, 103060, 
    103070, 103100, 103120, 103110, 103120, 103120, 103130, 103150, 103150, 
    103130, 103140, 103140, 103170, 103180, 103190, 103190, 103200, 103200, 
    103200, 103200, 103210, 103210, 103210, 103250, 103250, 103290, 103290, 
    103290, 103280, 103300, 103320, 103320, 103330, 103310, 103310, 103310, 
    103310, 103300, 103290, 103260, 103260, 103230, 103220, 103200, 103200, 
    103180, 103180, 103170, 103160, 103140, 103130, 103100, 103110, 103090, 
    103090, 103050, 103060, 103060, 103070, 103040, 103050, 103060, 103060, 
    103040, 102990, 102950, 102920, 102900, 102850, 102810, 102760, 102750, 
    102710, 102670, 102640, 102590, 102550, 102510, 102470, 102490, 102480, 
    102480, 102480, 102510, 102520, 102520, 102500, 102440, 102430, 102410, 
    102380, 102340, 102330, 102310, 102290, 102270, 102260, 102250, 102220, 
    102240, 102270, 102270, 102260, 102230, 102240, 102260, 102250, 102270, 
    102270, 102290, 102320, 102320, 102310, 102330, 102330, 102310, 102290, 
    102310, 102290, 102310, 102330, 102340, 102350, 102350, 102360, 102370, 
    102320, 102360, 102360, 102370, 102360, 102360, 102360, 102390, 102390, 
    102400, 102410, 102440, 102440, 102410, 102450, 102460, 102430, 102460, 
    102500, 102530, 102540, 102520, 102520, 102540, 102560, 102580, 102610, 
    102610, 102610, 102610, 102600, 102600, 102590, 102560, 102540, 102510, 
    102530, 102520, 102520, 102540, 102540, 102550, 102560, 102560, 102610, 
    102580, 102590, 102600, 102610, 102610, 102610, 102540, 102530, 102540, 
    102460, 102530, 102530, 102440, 102410, 102410, 102340, 102290, 102300, 
    102270, 102240, 102170, 102150, 102120, 102090, 102040, 101980, 101900, 
    101890, 101810, 101760, 101700, 101640, 101570, 101510, 101420, 101290, 
    101200, 101070, 100960, 100890, 100830, 100740, 100650, 100560, 100460, 
    100400, 100350, 100260, 100210, 100170, 100120, 100140, 100150, 100200, 
    100240, 100140, 100200, 100270, 100270, 100420, 100570, 100620, 100670, 
    100580, 100700, 100820, 101080, 101210, 101240, 101280, 101300, 101290, 
    101370, 101370, 101520, 101570, 101630, 101690, 101730, 101830, 101980, 
    102020, 102070, 102080, 102150, 102120, 102030, 102020, 102040, 102100, 
    102150, 102200, 102200, 102190, 102180, 102170, 102170, 102140, 102140, 
    102150, 102120, 102130, 102100, 102080, 102040, 102020, 101990, 101980, 
    101950, 101900, 101860, 101860, 101830, 101810, 101800, 101780, 101740, 
    101720, 101710, 101700, 101660, 101640, 101620, 101570, 101540, 101510, 
    101470, 101440, 101390, 101330, 101290, 101260, 101210, 101200, 101120, 
    101070, 101030, 100960, 100940, 100890, 100830, 100760, 100710, 100680, 
    100620, 100570, 100530, 100450, 100380, 100340, 100280, 100220, 100160, 
    100130, 100110, 100080, 100010, 99970, 99890, 99850, 99820, 99790, 99810, 
    99900, 99930, 99890, 99840, 99840, 99780, 99700, 99700, 99730, 99790, 
    99850, 99890, 99920, 99980, 100050, 100140, 100210, 100230, 100220, 
    100180, 100120, 100160, 100200, 100270, 100330, 100380, 100410, 100480, 
    100520, 100520, 100540, 100590, 100560, 100530, 100660, 100720, 100700, 
    100770, 100760, 100780, 100860, 100880, 100940, 101030, 101060, 101080, 
    101120, 101120, 101100, 101110, 101170, 101190, 101220, 101250, 101300, 
    101350, 101380, 101420, 101500, 101480, 101590, 101600, 101570, 101590, 
    101570, 101540, 101570, 101580, 101630, 101680, 101670, 101680, 101660, 
    101650, 101640, 101650, 101640, 101610, 101580, 101480, 101380, 101350, 
    101190, 101000, 100820, 100710, 100650, 100620, 100630, 100650, 100640, 
    100690, 100700, 100740, 100770, _, 100750, 100730, 100720, 100720, 
    100690, 100640, 100610, 100550, 100530, 100560, 100610, 100630, 100630, 
    100650, 100670, 100730, 100740, 100760, 100780, 100770, 100770, 100770, 
    100770, 100750, 100750, 100710, 100700, 100700, 100690, 100670, 100650, 
    100650, 100620, 100610, 100600, 100580, 100530, 100500, 100480, 100460, 
    100440, 100420, 100400, 100400, 100370, 100350, 100380, 100380, 100380, 
    100380, 100400, 100440, 100470, 100510, 100500, 100530, 100550, 100570, 
    100580, 100590, 100600, 100610, _, 100680, 100720, 100750, _, 100780, 
    100780, 100770, 100810, _, 100840, 100850, 100880, 100930, 100960, 
    100990, 101010, 101010, 101010, 101000, 101010, 101000, 101010, 101010, 
    101000, 101030, 101030, 101030, 101020, 100990, 101000, 100990, 100980, 
    100980, 100960, 100950, 100970, _, 101000, _, 101010, 100990, 100990, 
    100960, 100970, 100970, _, 101000, 101030, 101040, 101050, 101070, 
    101090, 101110, 101100, 101130, 101140, 101140, 101120, 101160, 101200, 
    101250, _, 101290, 101310, 101350, 101380, 101430, 101450, 101480, 
    101520, 101540, 101570, 101620, 101640, 101670, 101770, 101820, 101860, 
    101900, 101920, _, 101980, 102030, 102070, 102110, 102170, 102200, 
    102220, 102230, 102240, 102240, 102250, _, 102300, 102320, 102350, 
    102400, 102430, 102480, 102500, 102550, 102580, 102610, 102620, 102670, 
    102710, _, _, 102820, 102840, _, 102930, 102950, 102960, 102960, 102990, 
    103010, 103030, 103040, 103040, 103080, 103090, 103080, 103080, 103090, 
    103080, 103080, 103080, 103060, 103060, 103040, 103050, 103040, 103040, 
    103050, 103050, 103020, 103000, _, 102990, 102980, 102990, 102960, 
    102970, 102950, 102970, 102960, 102920, _, 102840, 102830, 102840, _, 
    102810, 102800, 102780, 102740, 102740, 102720, 102690, 102670, 102610, 
    102600, 102590, _, 102520, 102490, 102460, 102440, 102410, 102390, 
    102370, 102340, 102310, 102270, 102240, 102200, 102190, 102160, 102150, 
    102120, 102100, _, 102070, 102030, 102000, 101970, 101940, 101920, 
    101920, 101920, 101910, 101890, 101870, 101850, 101850, 101840, 101830, 
    101830, 101810, 101820, 101840, 101860, 101880, 101850, 101880, 101900, 
    101890, 101890, 101880, 101860, 101840, 101850, 101880, 101870, 101900, 
    101880, 101890, 101850, 101830, 101880, 101820, 101820, 101820, 101800, 
    101780, 101750, 101730, 101710, 101670, 101630, 101590, 101630, 101550, 
    101500, _, 101470, 101460, 101450, 101440, 101410, 101390, 101370, 
    101350, 101340, 101290, 101260, 101210, 101140, 101100, 100990, 100930, 
    100820, 100760, _, 100830, 100830, 100840, 100850, 100840, 100850, _, 
    100850, 100830, 100810, 100820, 100820, 100820, 100810, 100790, 100770, 
    100730, 100680, 100640, 100630, 100590, 100570, 100540, 100530, 100520, 
    100510, 100480, 100460, 100410, 100350, 100280, 100190, 100130, 100060, 
    99980, 99930, 99860, 99800, 99710, 99630, 99580, _, 99530, 99550, 99570, 
    99650, 99780, 99860, 100050, 100190, 100260, 100330, _, 100440, 100520, 
    100530, 100630, 100710, 100740, 100740, 100750, 100740, 100730, 100700, 
    100680, 100630, 100610, 100650, 100680, 100700, 100710, _, 100690, 
    100710, 100700, 100700, 100690, 100650, 100670, 100690, 100700, 100770, 
    100780, 100840, 100840, 100890, 100930, 100980, 101000, 101000, 101000, 
    100980, 100980, 100980, 100950, 100930, 100880, 100820, 100730, 100630, 
    100510, 100360, 100290, 100130, 100030, 99920, 99880, 99870, 99870, 
    99890, 99930, 99980, 100020, 100030, 100020, 100040, 100060, 100090, 
    100110, 100120, 100110, 100160, 100170, 100270, 100410, 100520, 100630, 
    100730, 100840, 100880, 100920, 101000, 100970, 100990, 101070, 101100, 
    101140, 101090, 101170, 101230, _, 101290, 101280, 101310, 101320, 
    101320, 101340, _, 101370, 101380, 101350, 101350, 101350, 101360, 
    101360, 101380, 101410, 101460, 101510, 101570, 101620, 101650, 101740, 
    101780, 101820, 101880, 101920, 101940, 101920, 101940, 101960, 101940, 
    101900, _, 101790, 101750, 101720, 101690, 101650, 101580, 101540, 
    101480, 101450, _, 101390, 101340, 101300, 101290, 101290, 101300, 
    101310, 101280, 101240, 101210, 101180, 101140, 101120, 101060, 100970, 
    100900, _, 100760, 100730, 100650, 100620, 100610, 100580, 100550, 
    100510, 100480, 100470, 100490, 100500, 100540, 100570, 100550, 100460, 
    100350, 100270, _, 100440, 100700, 100830, 100890, 101050, 101130, 
    101250, 101280, 101190, 101320, 101320, 101430, 101390, 101460, 101480, 
    101480, 101550, 101550, 101620, 101670, 101760, 101710, 101760, 101850, 
    101920, 101990, 102040, 102080, 102130, 102170, 102200, 102250, 102280, 
    102290, 102300, 102310, 102310, 102290, 102290, 102310, 102320, 102330, 
    102350, 102370, 102370, _, 102360, 102350, 102330, 102290, 102260, 
    102250, 102240, 102190, 102170, 102170, 102130, 102120, 102090, 102050, 
    102020, 101970, 101910, 101860, 101790, 101740, 101700, 101710, 101670, 
    101600, 101620, 101570, 101520, 101470, 101430, 101390, 101340, 101290, 
    101250, 101210, 101150, 101080, 101060, _, 100930, 100890, 100850, 
    100800, 100770, 100740, 100690, 100670, 100590, 100530, 100420, 100410, 
    100360, 100330, 100270, 100220, 100210, 100150, 100170, 100150, 100180, 
    100200, 100210, 100280, 100350, 100410, 100470, 100560, 100610, 100650, 
    100710, 100730, _, 100780, 100770, 100770, 100780, _, 100730, 100710, 
    100710, 100710, 100700, _, 100780, 100790, 100820, 100820, 100820, 
    100840, 100850, _, 100880, 100890, 100920, 100940, 100940, _, 100930, 
    100910, 100900, 100890, 100880, 100870, 100890, 100890, 100880, 100870, 
    100850, 100840, 100830, _, 100800, 100790, 100790, 100790, 100780, 
    100780, 100770, 100760, 100760, 100750, 100740, 100720, 100700, 100700, 
    100700, 100700, 100690, 100690, 100670, 100660, 100660, 100660, _, 
    100640, 100640, 100640, 100640, 100680, 100670, 100670, 100700, 100710, 
    _, 100730, 100740, 100760, 100760, 100770, 100790, 100810, 100830, 
    100850, 100870, 100870, 100880, 100920, 100930, 100920, 100930, 100940, 
    100960, 100990, 101030, 101050, 101070, 101100, 101130, _, 101170, 
    101150, 101190, 101230, 101250, 101280, 101300, 101300, 101300, 101310, 
    101330, 101340, 101340, 101350, 101350, 101360, 101390, 101400, 101420, 
    101440, 101450, 101460, 101480, 101480, 101470, 101470, 101480, 101480, 
    101470, 101490, 101490, 101480, 101470, 101460, 101450, 101440, 101410, 
    101400, _, 101370, 101350, 101340, 101330, 101310, 101290, 101240, 
    101220, 101180, 101160, 101120, 101080, 101030, 100990, 100960, 100920, 
    100900, 100860, 100830, 100800, 100790, 100790, 100780, 100770, 100760, 
    100770, 100780, 100810, 100820, 100830, 100850, 100860, _, 100890, 
    100910, 100910, 100930, 100920, 100920, 100940, 100960, 100970, 100960, 
    100980, 101010, 101020, 101040, 101040, 101060, 101070, 101090, 101120, 
    101150, 101180, 101220, 101230, 101260, 101270, 101310, 101320, 101310, 
    101330, 101340, 101370, 101360, 101370, 101400, 101400, 101450, 101500, 
    101530, 101530, 101510, 101560, 101610, _, 101680, 101720, 101770, 
    101820, 101840, 101870, 101910, 101930, 101970, 101960, 101980, 102030, 
    102060, 102080, 102080, 102100, 102070, 102090, 102100, 102070, 102070, 
    102070, 102080, 102060, 102050, 102090, 102090, 102080, _, 102120, 
    102090, 102080, 102070, 102070, 102070, 102110, 102100, 102120, 102110, 
    102080, 102090, 102070, _, 102070, 102050, 102060, 102040, 102030, 
    102010, 102040, 102030, 101990, 101980, 101970, 101970, 101980, 101970, 
    101950, 101960, 101960, 101950, 101980, 102010, 101990, 101980, 101940, 
    101890, 101840, 101780, 101680, 101660, 101630, 101580, 101580, 101510, 
    101510, 101490, 101490, 101420, 101340, 101290, 101300, 101260, 101230, 
    101260, 101250, 101250, 101260, 101190, 101190, 101170, 101140, 101110, 
    101050, 101000, 100960, 100970, 100920, 100880, 100880, _, 100770, 
    100720, 100670, 100620, 100570, 100480, 100420, 100370, 100320, 100270, 
    100240, 100210, 100160, 100160, 100120, 100150, 100180, 100170, 100190, 
    100170, 100150, 100120, 100080, 100010, 99950, 99880, 99810, 99770, 
    99700, 99650, 99600, 99570, 99540, 99490, 99460, 99440, 99440, 99420, 
    99410, 99420, 99470, 99500, 99540, 99610, 99680, 99780, 99870, _, 100090, 
    100190, 100270, 100380, 100460, 100520, 100590, 100650, 100680, 100700, 
    100710, 100730, 100730, 100740, 100720, 100740, 100720, 100730, 100730, 
    100700, 100680, 100660, 100630, _, 100530, 100420, 100350, 100270, 
    100240, 100270, 100250, 100300, 100300, 100300, 100330, 100410, 100460, 
    100540, 100590, 100650, 100670, 100770, 100800, 100840, 100880, 100880, 
    100880, 100850, 100810, 100680, 100640, 100590, 100440, 100380, 100260, 
    100140, 100050, 99950, 99820, 99720, 99670, 99610, 99510, 99500, 99570, 
    99680, 99700, 99850, 99970, 100070, 100180, 100300, 100460, 100540, 
    100620, 100700, 100790, 100880, 100940, 101010, 101070, 101110, 101180, 
    101280, 101340, 101370, 101410, 101440, 101510, 101560, 101600, 101610, 
    101630, 101640, 101640, 101650, 101620, 101550, 101470, 101400, 101310, 
    101160, 100960, 100800, 100660, 100400, 100260, 100040, 99870, 99820, 
    99760, 99760, 99780, 99850, 99960, 100070, 100200, 100340, 100470, 
    100560, _, 100730, 100820, 100890, 100970, 101090, 101180, 101280, 
    101350, 101450, 101530, 101600, 101640, 101750, 101770, 101790, 101780, 
    101800, 101790, 101760, 101740, 101660, 101590, 101530, 101440, 101310, 
    101230, 101120, 101090, 101060, 101140, 101250, 101310, 101450, 101560, 
    101750, 102060, 102160, 102270, 102400, 102450, 102530, 102610, 102690, 
    102690, 102710, 102750, 102780, 102790, 102770, 102710, 102680, 102660, 
    102620, 102610, 102560, 102530, 102500, 102410, 102380, 102340, 102260, 
    102160, 102110, 102020, 101990, 101970, 101950, 101910, 101880, 101840, 
    101830, 101800, 101760, 101710, 101660, 101640, 101620, 101630, 101610, 
    101600, 101580, 101620, 101560, 101560, 101550, 101510, 101490, 101470, 
    101490, 101490, 101480, 101500, 101540, 101550, 101520, 101540, 101580, 
    101590, 101600, 101630, 101610, 101630, 101660, 101660, 101620, 101600, 
    101600, 101590, 101530, 101460, 101480, 101440, 101420, 101320, 101300, 
    101360, 101360, 101320, 101260, 101190, 101120, 101070, 100980, 100900, 
    100940, 100970, 100980, 100950, 100950, 100950, 100950, 100890, 100890, 
    100870, 100870, 100840, 100870, 100870, 100860, 100840, 100820, 100760, 
    100720, 100690, 100700, 100630, 100530, 100510, 100500, 100530, 100550, 
    100540, 100510, 100470, 100450, 100420, 100380, 100340, _, 100200, 
    100220, 100240, 100220, 100200, 100200, 100200, 100180, 100160, 100100, 
    100120, 100080, 100010, 100040, 100090, 100140, 100060, 100000, 100040, 
    100070, 100060, _, 99970, 100060, 100040, 100090, 100170, 100230, 100270, 
    100320, 100340, 100340, 100330, 100330, 100330, 100290, 100230, 100130, 
    100100, 100090, 100030, 100020, 100040, 99980, 99970, 99940, 99950, 
    99930, 99920, 99930, 99970, 100040, 100080, _, 100170, 100220, 100270, 
    100330, 100370, 100410, 100450, _, 100540, 100580, 100610, 100650, 
    100670, 100680, 100710, 100730, 100750, 100750, 100750, 100750, 100770, 
    100780, 100790, 100800, 100830, 100830, 100830, 100830, 100820, 100810, 
    100800, 100780, 100800, 100810, 100810, 100810, 100840, 100870, 100890, 
    100910, 100930, 100950, _, 101050, 101110, 101160, 101200, 101230, 
    101260, 101280, 101320, 101330, 101320, 101310, 101290, 101290, 101300, 
    101310, 101310, 101310, 101260, 101280, 101230, 101190, 101140, 101100, 
    101040, 100990, 100960, 100950, 100910, 100860, 100840, 100790, 100730, 
    100700, 100680, 100640, 100610, 100630, 100630, 100630, 100630, 100630, 
    100630, 100630, 100640, 100630, 100650, 100680, 100720, 100770, 100820, 
    100830, 100870, 100890, 100900, 100900, 100880, 100840, 100790, 100760, 
    100690, 100650, 100590, 100550, 100510, 100440, 100380, 100300, 100240, 
    100200, 100170, 100140, _, 100130, 100160, 100200, 100260, 100310, 
    100370, 100410, 100450, 100480, 100530, 100570, 100600, 100630, 100650, 
    100670, 100690, 100730, 100770, 100830, 100900, 100940, 100970, 100990, 
    101020, 101070, 101130, 101180, 101230, 101230, 101250, 101260, 101250, 
    101210, 101190, 101170, 101140, 101130, 101100, 101090, 101050, 101050, 
    101040, 101040, 101060, 101070, 101080, 101110, 101150, 101200, 101250, 
    101300, 101350, 101440, 101480, 101510, 101550, 101600, 101620, 101660, 
    101680, _, 101740, 101790, 101820, 101850, 101870, 101850, 101840, 
    101850, 101850, 101880, _, 101910, 101950, 101980, 101990, 101960, 
    102000, 102010, 102020, 102020, 102010, 102010, 102010, 102000, 102010, 
    102010, 102000, 101990, 102000, 102000, 101990, 102010, 102010, 102030, 
    102060, 102110, 102140, 102140, 102160, 102180, 102190, 102190, 102190, 
    102180, 102170, 102160, 102160, _, 102110, 102100, 102100, 102070, _, 
    102010, 101990, 101960, 101920, 101900, 101880, 101840, 101770, 101720, 
    101670, 101600, 101570, 101520, 101430, 101360, 101300, 101260, 101200, 
    101150, 101080, 101040, 100980, 100930, 100900, 100880, 100870, 100860, 
    100860, 100810, _, 100830, 100830, 100830, 100840, 100840, 100810, 
    100800, 100750, 100720, 100690, 100700, 100700, 100700, 100700, 100660, 
    100630, 100600, 100560, 100540, 100520, 100470, 100440, 100410, 100400, 
    100380, 100370, 100350, 100360, 100350, 100360, 100350, 100340, 100340, 
    100300, 100270, 100230, 100170, 100160, 100130, 100120, 100100, _, 
    100080, 100070, 100050, 100020, 100030, 100050, 100090, 100110, 100140, 
    100130, _, 100130, 100100, 100120, 100050, 100110, 100190, 100250, 
    100320, _, 100400, 100460, 100540, 100530, 100640, 100740, 100810, 
    100860, 100970, 101020, 101070, 101100, 101180, 101220, 101280, 101320, 
    101370, 101400, 101390, 101410, 101420, 101440, 101440, 101450, 101440, 
    101420, 101400, 101380, 101370, 101360, 101350, 101270, 101260, 101220, 
    101230, 101240, 101220, 101150, 101170, 101100, 101130, 101150, 101010, 
    101070, 101030, 100930, 100960, 100840, 100790, 100800, 100680, 100590, 
    100580, 100510, 100490, 100490, 100460, 100410, 100480, 100460, 100430, 
    100410, _, _, 100370, 100360, 100330, 100290, 100280, 100260, 100220, 
    100140, 100050, 99880, 99800, 99750, 99710, 99590, 99480, 99450, 99230, 
    99120, 99020, 98830, 98670, _, 98440, 98270, 98160, 98030, 97970, 97950, 
    97960, 98010, 98010, 97980, 98070, 98190, 98280, 98350, 98400, 98470, 
    98530, 98570, 98470, 98640, 98770, 98840, 98910, 99000, 99140, 99320, 
    99320, 99500, 99600, 99730, 99850, 99990, 100100, 100230, 100300, 100390, 
    100490, 100590, 100670, 100700, 100790, 100850, 100910, 100950, 101010, 
    101070, _, 101170, 101210, 101260, 101300, 101330, 101340, 101350, 
    101350, 101360, 101370, 101390, 101390, 101410, 101410, 101420, 101430, 
    101450, 101450, 101450, 101450, 101470, 101470, 101480, 101490, 101510, 
    101510, 101520, 101530, 101530, 101530, 101520, 101490, 101500, 101470, 
    101480, 101460, 101430, 101410, 101390, 101350, 101300, 101220, 101140, 
    101140, 101100, 101080, 101090, 101020, 100930, 100850, 100820, 100830, 
    100780, 100720, 100630, 100610, 100570, 100550, 100490, 100450, _, 
    100380, 100360, 100370, 100360, 100350, 100360, 100330, 100360, 100350, 
    100350, _, 100300, 100260, 100230, _, 100130, 100070, 99990, 99900, 
    99850, 99810, 99750, 99730, 99660, 99660, 99620, 99600, 99510, 99500, 
    99560, 99560, 99550, 99550, 99530, 99520, 99510, 99510, 99480, 99500, 
    99480, 99490, 99520, _, 99540, 99570, 99610, 99660, 99700, 99750, 99820, 
    99840, 99890, 99950, 100020, 100070, 100110, 100170, 100230, 100260, 
    100320, 100380, 100430, 100500, 100560, 100600, 100640, 100670, 100680, 
    100710, 100710, 100730, 100770, 100840, 100890, 100920, 100960, 101020, 
    101070, 101090, 101140, 101220, 101240, _, 101330, 101320, 101340, 
    101370, 101350, 101330, 101330, 101310, _, 101230, 101220, 101230, 
    101230, 101230, 101180, 101160, 101140, 101080, 100990, 100870, 100800, 
    100680, _, 100620, 100560, 100480, 100500, 100450, 100340, 100310, 
    100300, 100260, 100220, 100220, 100250, 100240, 100250, 100230, 100180, 
    100160, 100170, 100090, 100060, 100020, 99970, 99920, 99900, 99870, 
    99860, 99830, 99800, 99760, 99720, 99710, 99710, 99740, 99740, 99760, 
    99820, 99850, 99910, 99920, 100000, 100060, 100110, 100180, 100240, 
    100270, 100360, 100450, 100560, 100640, 100720, 100790, 100890, 100960, 
    101000, 101040, 101100, 101130, 101150, 101180, 101210, 101190, 101200, 
    101190, 101180, 101170, 101150, 101140, 101110, 101080, 101070, 101060, 
    _, 100970, 100940, 100900, 100850, 100770, 100740, 100710, 100670, 
    100570, 100400, 100240, 100140, 100080, _, 99800, 99630, 99600, 99590, 
    99610, 99540, 99590, 99590, 99620, 99670, 99700, 99720, 99730, 99760, 
    99810, 99870, 99950, 100060, _, 100250, 100330, 100400, 100460, 100530, 
    100560, 100600, 100660, 100670, 100710, 100730, 100740, 100760, 100820, 
    100850, 100880, 100900, 100930, 100950, 100960, 100970, 100990, 101010, 
    101010, 101020, 101040, 101040, 101050, 101050, 101050, 101040, 101030, 
    101040, 101060, 101050, 101070, 101090, 101090, _, 101140, 101170, 
    101220, 101210, 101230, 101250, 101270, 101290, 101290, 101300, 101320, 
    101330, 101350, 101340, 101320, 101350, 101350, 101330, 101330, 101310, 
    101310, 101310, 101300, 101320, 101330, 101340, 101330, 101310, 101270, 
    101260, 101230, 101160, 101210, 101280, 101230, 101160, 101070, 101120, 
    101060, 100820, 100940, 100910, 100860, 100840, 100730, 100620, 100580, 
    100420, _, 100350, 100220, 100180, 100070, 100010, 99930, 99930, 99910, 
    99850, 99840, 99790, 99780, 99950, 99920, 99890, 99840, 99850, 99780, 
    99790, 99740, 99730, 99720, _, 99680, 99660, 99630, 99630, 99620, 99580, 
    99540, 99510, 99480, 99440, 99460, 99420, 99390, _, 99350, 99320, 99300, 
    99290, 99270, 99280, 99250, 99230, 99250, 99240, 99250, 99220, 99240, 
    99220, 99190, 99180, 99150, 99110, 99070, 99040, 99030, 99020, 99000, 
    98970, 98950, 98930, 98900, 98880, 98860, 98850, 98870, 98890, 98910, 
    98940, 99010, 99060, 99100, 99140, 99160, 99200, 99230, 99240, 99280, 
    99310, 99360, 99390, 99430, 99440, 99490, 99510, 99520, 99560, 99570, 
    99570, 99590, 99570, 99600, _, 99640, _, 99690, 99710, 99700, 99690, 
    99710, 99720, 99730, 99720, 99710, 99740, 99730, 99730, _, 99710, 99710, 
    99670, 99650, 99650, 99690, 99720, 99760, 99780, 99810, 99830, 99850, 
    99880, 99880, 99900, 99920, 99930, 99930, 99960, 99960, 100000, 100010, 
    100050, 100090, 99990, 99960, 100000, 100080, 100160, 100200, 100200, 
    100280, 100300, 100320, 100390, 100440, 100410, 100450, 100480, 100500, 
    100510, 100500, 100480, 100460, 100420, 100370, 100350, 100350, 100320, 
    100300, 100250, 100210, 100200, 100190, 100220, 100210, 100180, 100180, 
    100180, 100150, 100160, 100170, 100140, 100160, 100170, 100160, 100150, 
    _, _, 100110, 100120, 100180, 100230, 100290, 100340, 100430, 100490, 
    100560, 100610, 100660, 100710, 100770, 100830, 100870, 100900, 100930, 
    100970, 100970, 100980, 100990, 100990, 101010, 101070, 101100, _, 
    101070, _, 101100, 101110, 101090, 101100, 101070, 101080, 101100, 
    101160, 101210, 101240, 101270, 101260, 101310, 101340, 101350, 101340, 
    101360, 101360, 101330, 101310, 101340, 101340, 101330, 101330, 101300, 
    101330, 101320, 101320, 101280, _, 101200, 101210, 101230, 101260, 
    101240, 101210, 101210, 101210, 101210, 101200, 101150, 101140, 101170, 
    101130, 101130, 101110, 101120, 101110, 101130, 101130, 101110, 101110, 
    101100, 101100, 101110, 101120, 101130, 101150, 101180, 101170, 101180, 
    101200, 101180, 101190, 101160, 101170, 101200, 101200, 101190, 101190, 
    101200, 101210, 101210, 101200, 101210, 101230, 101250, 101250, 101270, 
    101310, 101340, 101390, 101430, 101440, 101460, 101490, 101530, 101530, 
    101530, 101540, 101570, 101590, 101580, 101580, 101600, 101610, 101620, 
    101610, 101590, 101580, 101580, 101590, _, 101570, 101550, 101540, 
    101500, 101440, 101420, 101370, 101330, 101290, 101260, 101200, 101180, 
    101130, 101110, 101080, 101080, 101110, 101090, 101050, 101000, 100970, 
    100950, 100930, 100900, 100880, 100860, 100820, 100810, 100740, 100710, 
    100640, 100570, 100590, 100520, 100540, 100520, 100500, 100440, 100390, 
    100370, 100340, 100330, 100310, 100300, 100290, 100290, 100280, 100250, 
    100260, 100250, 100300, 100350, 100420, 100450, 100460, 100490, 100520, 
    100500, 100450, 100430, 100420, 100360, 100320, 100280, 100250, 100200, 
    100180, 100160, 100140, 100130, 100100, 100070, 100070, 100030, _, 99900, 
    99910, 99860, 99830, 99770, 99730, 99720, 99680, 99680, 99680, 99620, 
    99610, 99590, 99630, 99640, 99660, 99730, 99800, 99880, 99950, _, 100100, 
    100170, 100230, 100300, 100340, 100340, 100340, 100350, 100380, 100360, 
    100390, 100380, 100410, 100440, 100470, 100500, 100550, 100600, 100580, 
    100590, 100650, 100630, 100610, 100580, 100560, 100530, 100460, 100470, 
    100400, 100310, 100240, 100160, 100030, 99940, 99870, 99780, 99770, 
    99750, 99760, 99790, 99860, 99930, 99980, 100020, 100070, 100110, 100160, 
    100200, 100250, 100320, 100380, 100450, 100490, 100540, 100600, 100660, 
    100700, 100740, 100790, 100810, 100820, 100800, 100820, 100810, 100790, 
    100760, 100700, 100620, 100600, 100560, 100510, 100460, 100420, 100380, 
    100310, 100230, 100190, 100130, 100100, 100050, 100050, 100040, 100080, 
    100140, 100200, 100280, 100350, 100460, 100540, 100620, 100670, 100700, 
    100770, 100820, 100850, 100910, 100950, 100990, 101020, 101000, 101010, 
    101010, 101010, 100960, 100980, 100940, 100890, 100820, 100810, 100760, 
    100730, 100640, 100570, 100490, 100440, 100380, 100350, 100360, 100320, 
    100310, 100320, 100330, 100350, 100350, 100380, 100410, 100410, 100440, 
    100490, 100550, 100600, 100640, 100730, 100770, 100830, 100890, 100980, 
    101030, 101060, 101130, 101170, 101200, 101250, 101280, 101360, 101370, 
    101380, 101410, 101440, 101450, 101440, 101450, 101450, 101470, 101460, 
    101460, 101480, 101500, 101520, 101540, 101590, 101630, 101660, 101690, 
    101740, 101770, 101820, 101850, 101880, 101900, 101930, 101970, 101990, 
    101960, 101930, 101960, 101930, 101930, 101880, 101860, 101810, 101780, 
    101770, 101730, 101680, 101640, 101640, 101630, 101590, 101600, 101600, 
    101610, 101600, 101580, 101600, 101580, 101540, 101490, 101490, 101440, 
    101380, 101330, 101250, 101180, 100910, 100980, 100850, 100730, 100590, 
    100470, 100420, 100330, 100230, 100180, 100150, 100120, 100130, 100110, 
    100140, 100160, 100160, 100190, 100190, 100140, 100130, _, 100100, 
    100120, 100150, 100160, 100180, 100200, 100220, 100210, 100230, 100250, 
    100310, 100270, 100320, 100360, 100400, 100450, 100470, 100490, 100530, 
    100570, 100580, 100610, 100670, 100700, _, 100790, 100860, 100900, 
    100940, 101010, 101050, 101070, 101100, 101110, 101090, 101120, 101130, 
    101110, 101080, 101050, 101020, 101020, 100990, 100940, 100900, 100900, 
    100870, 100800, 100760, 100700, 100670, 100680, 100650, 100650, 100640, 
    100610, 100600, 100550, 100490, 100500, 100470, 100480, 100470, 100440, 
    100420, 100440, 100410, 100400, _, 100430, 100450, 100410, 100410, 
    100400, 100400, 100400, 100350, 100340, 100310, 100300, 100270, 100250, 
    100240, 100220, 100200, 100190, 100180, 100170, 100160, 100170, 100160, 
    100150, 100140, 100140, 100130, 100130, _, 100170, 100180, 100210, 
    100240, 100280, 100310, 100360, 100390, 100410, 100480, 100580, 100630, 
    100690, 100800, 100870, 100900, 100940, 100980, 101020, 101030, 101000, 
    100990, 100960, 100930, 100880, 100830, 100820, 100800, 100750, 100690, 
    100660, 100590, 100530, 100520, 100480, 100470, 100510, 100480, 100440, 
    100480, 100520, 100550, 100580, 100600, 100600, 100640, _, 100740, _, 
    100810, 100780, 100800, 100850, 100880, 100880, 100880, 100900, _, 
    100950, 100960, 101020, 101060, 101110, 101170, 101220, 101280, 101320, 
    101360, 101400, 101430, 101470, 101480, 101500, 101450, 101410, 101390, 
    101330, 101310, 101240, 101170, 101130, 101070, 101060, 101030, 101030, 
    101040, 101070, 101060, 101060, 101090, 101100, 101090, 101080, 101120, 
    101180, 101180, 101240, 101270, 101320, 101320, 101330, 101320, 101370, 
    101370, 101350, 101350, 101330, 101320, 101280, 101320, 101350, 101400, 
    101430, 101410, _, 101460, 101490, 101540, 101570, 101610, 101670, 
    101750, 101760, 101810, 101840, 101850, 101860, 101890, 101920, 101970, 
    102000, 102050, 102080, 102160, 102190, 102220, 102190, 102250, 102230, 
    102280, 102270, 102240, 102230, _, 102240, 102250, 102230, 102200, 
    102180, 102200, 102140, 102110, 102070, 102050, 102000, 101990, 101970, 
    101980, 101970, 101960, 101960, 101930, 101900, 101910, 101890, 101860, 
    _, 101850, 101850, 101850, 101840, 101820, 101830, 101820, 101790, 
    101750, 101710, 101730, 101730, 101760, 101750, 101780, 101800, 101810, 
    101830, 101850, 101890, 101870, 101850, 101850, 101920, 101920, 102010, 
    102030, 102060, 102120, 102090, 102130, 102170, 102240, 102330, _, 
    102360, 102390, 102410, 102420, 102450, 102490, 102530, 102530, 102510, 
    102530, 102530, 102530, 102510, 102500, 102510, 102500, 102500, 102490, 
    102460, 102440, 102430, 102400, 102380, 102350, 102320, 102320, 102280, 
    102260, 102260, 102250, 102220, 102180, 102130, 102130, 102110, 102060, 
    _, 102000, 101960, 101930, 101910, _, 101860, 101830, 101800, 101760, 
    101730, 101680, 101660, 101650, 101620, 101610, 101600, 101600, 101600, 
    101550, 101520, 101540, 101510, 101490, 101480, 101450, 101460, 101440, 
    101420, 101430, 101390, 101370, 101400, 101420, 101460, _, 101500, 
    101540, 101550, 101560, 101560, 101570, 101550, 101500, 101470, 101370, 
    101290, 101210, 101230, 101190, 101200, 101120, 100970, 100910, 100890, 
    100900, 100850, 100850, 100790, 100730, 100700, 100630, 100610, 100550, 
    100460, 100390, 100310, _, 100380, 100290, 100230, 100220, 100180, 
    100180, 100180, 100070, 99980, 99910, 99850, 99750, 99650, 99620, 99560, 
    99550, 99500, 99470, 99480, 99420, 99470, 99460, _, 99470, 99430, 99430, 
    99420, 99400, 99370, 99410, 99410, 99420, 99530, 99560, 99620, 99660, 
    99710, 99730, 99770, _, 99790, 99790, 99770, 99760, 99800, 99820, 99860, 
    99890, 99920, 99960, 100030, 100050, 100040, 100050, 100080, 100120, 
    100150, 100180, 100170, 100180, 100190, 100210, 100230, 100220, 100230, 
    100250, 100290, 100320, 100360, 100370, 100390, 100400, 100420, 100440, 
    100460, 100470, 100470, 100480, 100500, 100520, 100540, 100570, 100590, 
    100620, 100610, 100630, 100640, 100640, 100650, 100670, 100690, 100750, 
    100790, 100810, 100830, 100840, 100870, 100900, 100910, 100940, 100940, 
    100950, 100960, 101030, 101040, 101020, 101030, 101020, 101010, 101000, 
    101010, 101020, 100990, 100970, 100950, 100980, 100970, 100960, 100980, 
    100920, 100910, 100900, 100900, 100900, 100940, 100900, 100860, 100800, 
    100780, 100730, 100710, 100710, 100650, 100610, _, 100580, 100580, 
    100530, 100520, 100520, 100530, 100570, 100570, 100580, 100580, 100570, 
    100580, 100590, 100600, 100570, 100510, 100570, 100600, 100560, 100570, 
    100530, 100560, 100590, 100560, 100530, 100510, 100470, 100480, 100480, 
    _, 100490, 100490, 100530, 100500, 100480, 100460, 100450, 100420, 
    100370, 100350, 100370, 100370, 100380, 100370, 100380, 100360, 100350, 
    100370, 100340, 100320, 100330, 100320, 100300, 100290, 100280, 100310, 
    100380, 100400, 100390, 100450, 100470, 100500, 100490, 100470, 100480, 
    100520, 100570, 100540, 100530, 100560, 100580, _, 100630, 100620, 
    100660, 100660, 100690, 100700, 100730, 100760, 100800, 100820, 100800, 
    100810, 100810, _, 100830, 100830, 100850, 100860, 100880, 100890, 
    100900, 100920, 100950, 100950, 100960, 100980, 101010, 101020, 101040, 
    101050, 101070, 101080, 101080, 101080, 101100, 101090, 101060, 101070, 
    101070, 101090, 101100, 101100, 101070, 101070, 101080, 101080, 101070, 
    101050, 101020, 101000, 100990, 100990, 100950, 100950, 100910, 100880, 
    100840, 100820, 100770, 100740, 100710, 100650, 100610, 100510, 100480, 
    100410, 100290, 100090, 99930, 99790, 99700, _, 99330, 99210, 99120, 
    98940, 98770, 98660, 98650, 98750, 98770, 98850, 98910, 98940, 98950, 
    98970, 98970, 98950, 98980, 98980, 98970, 98990, 98970, 98940, 98910, 
    98870, 98860, 98810, 98810, 98790, 98780, 98770, 98750, 98740, 98750, 
    98770, 98780, 98790, 98800, 98800, 98790, 98770, 98730, 98620, 98620, 
    98630, 98630, 98650, 98670, 98710, 98650, 98700, 98730, 98750, 98670, 
    98690, 98660, 98720, 98780, 98720, 98760, 98840, 98860, 98840, 98900, 
    98860, 98830, 98880, 98900, 98930, _, _, 98880, _, 98910, 98900, 98940, 
    99020, _, 99040, _, 99080, 99060, 99110, 99150, 99150, 99180, 99180, 
    99180, 99200, 99220, 99300, 99340, 99340, 99350, 99390, 99430, 99480, 
    99530, 99580, 99630, 99670, 99700, 99730, 99800, 99900, 99940, 99990, 
    100040, 100080, _, 100180, 100220, 100280, 100330, 100370, 100390, 
    100440, 100480, 100530, 100560, 100590, 100600, 100650, 100690, 100700, 
    100720, 100750, 100770, 100790, 100820, 100860, 100890, 100860, _, 
    100850, 100850, 100870, 100820, 100820, 100810, 100860, 100850, 100830, 
    100790, _, 100800, 100800, 100780, 100760, _, 100770, 100780, 100780, 
    100770, _, 100740, 100740, 100720, 100680, 100700, 100730, 100750, 
    100760, 100790, 100790, 100840, 100860, 100850, 100850, 100830, 100790, 
    100790, 100770, 100800, _, 100840, 100820, 100810, 100760, 100700, 
    100700, 100660, 100640, 100560, 100510, 100440, 100350, 100300, 100230, 
    100130, 100020, 99960, 99870, 99790, 99730, 99680, 99630, 99600, 99550, 
    99550, 99530, 99550, 99570, 99600, 99620, 99660, 99720, 99780, 99840, 
    99920, 99980, 100040, 100110, 100200, 100250, _, 100350, 100390, 100460, 
    100500, 100560, 100590, 100610, _, 100670, 100700, 100720, 100740, 
    100760, 100750, 100780, 100780, 100770, 100770, 100770, 100760, 100750, 
    100760, 100770, 100750, 100740, 100750, 100800, 100810, 100820, 100850, 
    100870, 100910, 100930, 100970, 101000, 101030, 101040, 101080, 101090, 
    101140, 101170, 101200, 101220, 101250, 101290, 101320, 101350, 101360, 
    101360, 101340, 101320, 101300, 101270, 101250, 101210, 101190, 101200, 
    101190, 101170, 101170, 101150, 101140, 101140, 101150, 101150, _, 
    101120, 101100, 101070, 101050, 100990, 100920, 100850, 100730, 100660, 
    100600, 100500, _, 100300, 100200, 100110, 100020, 99910, 99760, _, 
    99450, 99270, 99150, 99040, 99010, 98980, 98940, 99030, 99020, 98990, 
    99010, 98990, 98880, 98740, 98700, 98710, 98650, 98650, 98680, 98700, 
    98750, 98750, 98870, 98970, 99110, 99260, 99400, 99590, 99720, 99730, 
    99870, 100080, 100280, 100410, 100480, 100560, 100630, 100720, 100800, 
    100870, 100940, 101010, 101080, 101150, 101190, 101210, 101210, 101210, 
    101200, 101210, 101190, 101160, 101120, 101060, 101010, 100980, 100920, 
    100910, 100880, 100850, 100830, 100770, 100760, 100710, 100690, 100640, 
    100560, 100520, 100440, 100370, 100260, 100180, 100140, 100090, 100050, 
    99990, 99950, 99910, 99880, 99840, 99810, 99800, _, 99740, 99740, 99730, 
    99720, 99700, 99700, 99730, 99650, 99530, 99480, 99350, 99250, 99130, 
    99050, 99010, 98940, 98950, 98950, 99030, 99120, 99230, 99370, 99500, 
    99650, 99770, 99880, 99970, 100080, 100220, 100340, 100450, 100570, 
    100670, 100740, 100830, 100940, 101020, 101100, 101180, 101260, 101300, 
    101350, 101390, 101390, 101390, 101400, 101410, 101440, 101450, 101470, 
    101530, 101570, 101600, 101630, 101620, 101640, 101620, 101600, 101530, 
    101480, 101440, 101370, 101290, 101220, 101170, 101130, 101060, 100980, 
    100870, _, 100750, _, 100610, 100560, 100530, 100530, 100560, 100600, 
    100640, 100690, 100750, 100800, 100880, 100980, 101080, 101140, 101180, 
    101230, 101270, 101310, 101380, 101400, 101420, 101470, 101480, 101510, 
    101520, 101530, 101570, 101640, 101650, 101630, 101650, 101620, 101570, 
    101560, 101530, 101500, 101440, 101400, 101370, 101320, 101310, 101310, 
    101310, 101310, 101340, 101360, 101340, 101350, 101360, 101380, 101400, 
    101400, 101390, 101420, 101450, 101420, 101410, 101400, 101370, 101350, 
    101280, 101230, 101240, 101170, 101140, 101080, 101070, 101060, 101020, 
    101010, 101000, 101020, 101030, 101040, 101030, 101050, 101080, 101100, 
    101130, 101130, 101160, 101200, 101230, 101260, 101260, 101320, 101340, 
    101370, 101380, 101400, 101420, 101420, 101430, 101480, 101490, 101520, 
    101550, 101530, 101540, 101530, 101570, 101610, 101620, 101640, 101660, 
    101670, 101700, 101700, 101710, 101720, 101750, 101760, 101790, 101790, 
    101810, 101800, 101820, 101820, 101830, 101810, 101810, 101830, 101830, 
    101830, 101800, 101810, 101830, 101780, 101740, 101770, 101790, 101730, 
    101670, 101660, 101610, 101580, 101560, 101540, 101500, 101450, 101420, 
    101390, 101380, 101370, 101320, 101280, 101260, 101270, 101230, 101220, 
    101190, 101200, 101230, 101240, 101210, 101180, 101140, 101110, 101090, 
    101060, 101000, 100970, 100920, 100860, 100790, 100760, 100700, 100630, 
    100560, 100470, 100390, 100320, 100280, 100240, 100210, 100170, 100130, 
    100100, 100060, 100020, 99990, 99940, 99910, 99880, 99870, 99880, 99910, 
    99930, 99930, 99900, 99880, 99880, 99850, 99830, 99850, 99870, 99920, 
    99980, 100060, 100130, 100190, 100250, 100310, 100400, 100440, 100490, 
    100540, 100600, 100670, 100730, 100790, 100830, 100860, 100870, 100900, 
    100940, 100970, 100990, 101010, 101000, 101030, 101030, 101080, 101100, 
    101080, 101100, 101090, 101060, 101080, 101100, 101100, 101080, 101110, 
    101120, 101150, 101190, 101210, 101250, 101300, 101340, 101400, 101450, 
    101470, 101490, 101510, 101570, 101590, 101620, 101690, 101720, 101720, 
    101730, 101750, 101770, 101790, 101810, 101820, 101830, 101810, 101820, 
    101810, 101800, 101780, 101780, 101780, 101780, 101780, 101780, 101770, 
    101760, 101730, 101710, 101700, 101660, 101640, 101620, 101580, 101560, 
    101540, 101500, 101480, 101460, 101430, 101400, 101370, 101350, 101340, 
    101330, 101320, 101300, 101290, 101290, 101290, 101290, 101290, 101300, 
    101310, 101320, 101340, 101330, 101340, 101350, 101360, 101350, 101340, 
    101370, 101390, 101400, 101400, 101400, 101400, 101400, 101440, 101430, 
    101440, 101430, 101430, 101430, 101450, 101460, 101470, 101450, 101450, 
    101470, 101470, 101460, 101440, 101440, 101440, 101430, 101420, 101380, 
    101360, 101350, 101330, 101320, 101310, 101300, 101290, 101250, 101230, 
    101210, 101200, 101170, 101180, 101150, 101150, 101100, 101110, 101080, 
    101040, 101010, 100920, 100910, 100870, 100820, 100800, 100740, 100730, 
    100710, 100700, 100660, 100650, 100630, 100600, 100590, 100580, 100570, 
    100560, 100550, 100540, 100560, 100560, 100530, 100510, 100500, 100440, 
    100390, 100380, 100390, 100390, 100400, 100370, 100310, 100270, 100270, 
    100240, 100310, 100330, 100330, 100390, 100440, 100450, 100420, 100420, 
    100460, 100390, 100340, 100290, 100290, 100270, 100290, 100270, 100220, 
    100180, 100220, 100170, 100140, 100040, 99970, 99860, 99810, 99710, 
    99500, 99340, 99270, 99190, 99220, 99180, 98900, 98930, 98930, 98820, 
    98670, 98510, 98450, 98230, 98110, 98130, 98110, 98180, 98190, 98150, 
    98150, 98120, 98050, 98060, 98060, 98090, 98060, 98050, 97990, 97940, 
    97880, 97890, 97830, 97830, 97860, 97820, 97850, 97870, 97850, 97820, 
    97820, 97800, 97780, 97760, 97730, 97730, 97750, 97760, 97780, 97790, 
    97800, 97790, 97780, 97800, 97790, 97770, 97770, 97760, 97760, 97770, 
    97790, 97820, 97850, 97850, 97870, 97930, 97980, 98020, 98050, 98070, 
    98120, 98130, 98190, 98230, 98290, 98310, 98340, 98360, 98380, 98400, 
    98420, 98440, 98450, 98460, 98490, 98520, 98520, 98550, 98550, 98570, 
    98580, 98580, 98590, 98600, 98600, 98630, 98670, 98720, 98780, 98810, 
    98830, 98840, 98870, 98900, 98930, 98950, 98970, 99000, 99010, 99040, 
    99070, 99060, 99070, 99080, 99100, 99110, 99130, 99150, 99170, 99180, 
    99200, 99240, 99290, 99330, 99360, 99370, 99370, 99370, 99380, 99360, 
    99360, 99380, 99390, 99420, 99460, 99500, 99510, 99540, 99550, 99580, 
    99600, 99620, 99640, 99700, 99730, 99770, 99810, 99840, 99860, 99890, 
    99890, 99890, 99900, 99880, 99890, 99890, 99900, 99900, 99910, 99900, 
    99880, 99850, 99850, 99840, 99840, 99870, 99900, 99950, 99990, 100020, 
    100060, 100110, 100180, 100200, 100220, 100230, 100260, 100240, 100210, 
    100210, 100190, 100100, 100080, 100080, 99990, 99950, 99920, 99840, 
    99760, 99700, 99690, 99590, 99630, 99610, 99560, 99650, 99590, 99530, 
    99470, 99520, 99560, 99570, 99550, 99580, 99580, 99540, 99530, 99440, 
    99450, 99450, 99440, 99460, 99580, 99590, 99640, 99650, 99670, 99690, 
    99790, 99810, 99830, 99850, 99850, 99850, 99850, 99880, 99910, 99930, 
    99950, 99990, 100000, 99990, 99950, 99970, 99950, 99950, 99900, 99940, 
    99970, 100000, 99970, 99970, 100040, 100110, 100110, 100160, 100150, 
    100180, 100160, 100140, 100090, 100030, 100020, 99980, 99970, 99960, 
    99970, 100000, 100020, 100000, 100020, 99980, 100010, 100000, 100000, 
    100010, 100010, 100020, 100010, 100000, 99970, 99960, 99920, 99870, 
    99820, 99770, 99730, 99690, 99650, 99590, 99520, 99430, 99330, 99240, 
    99140, 99060, 99010, 98950, 98910, 98860, 98820, 98770, 98720, 98670, 
    98610, 98580, 98540, 98500, 98440, 98430, 98420, 98410, 98410, 98390, 
    98410, 98410, 98400, 98400, 98380, 98390, 98420, 98460, 98500, 98540, 
    98550, 98600, 98600, 98640, 98670, 98650, 98580, 98580, 98570, 98590, 
    98600, 98640, 98620, 98600, 98600, 98570, 98550, 98540, 98510, 98500, 
    98480, 98480, 98490, 98490, 98490, 98520, 98520, 98530, 98540, 98550, 
    98570, 98590, 98580, 98600, 98580, 98590, 98580, 98550, 98510, 98500, 
    98440, 98400, 98380, 98350, 98330, 98340, 98360, 98370, 98370, 98380, 
    98400, 98420, 98410, 98420, 98440, 98440, 98460, 98490, 98510, 98550, 
    98560, 98550, 98550, 98550, 98550, 98540, 98530, 98540, 98560, 98570, 
    98580, 98600, 98620, 98620, 98620, 98610, 98600, 98590, 98580, 98580, 
    98590, 98580, 98580, 98590, 98580, 98600, 98620, 98640, 98650, 98660, 
    98680, 98720, 98750, 98770, 98810, 98860, 98930, 99000, 99040, 99130, 
    99160, 99200, 99240, 99260, 99310, 99360, 99410, 99470, 99580, 99660, 
    99730, 99790, 99910, 99970, 100060, 100150, 100210, 100310, 100410, 
    100490, 100580, 100660, 100750, 100840, 100880, 100950, 101020, 101100, 
    101160, 101230, 101290, 101370, 101420, 101440, 101490, 101500, 101500, 
    101500, 101500, 101490, 101510, 101510, 101510, 101490, 101520, 101520, 
    101520, 101520, 101550, 101590, 101600, 101620, 101640, 101680, 101720, 
    101750, 101750, 101750, 101740, 101730, 101710, 101650, 101640, 101580, 
    101510, 101500, 101450, 101390, 101370, 101320, 101290, 101280, 101190, 
    101110, 101060, 100990, 100910, 100800, 100740, 100660, 100540, 100510, 
    100440, 100340, 100240, 100200, 100200, 100140, 100030, 99980, 99930, 
    99850, 99790, 99720, 99680, 99580, 99630, 99630, 99570, 99490, 99460, 
    99490, 99470, 99500, 99520, 99540, 99530, 99460, 99310, 99370, 99430, 
    99370, 99310, 99280, 99260, 99280, 99290, 99240, 99270, 99280, 99310, 
    99320, 99360, 99390, 99410, 99450, 99510, 99520, 99520, 99550, 99610, 
    99610, 99620, 99650, 99670, 99680, 99730, 99750, 99790, 99820, 99850, 
    99890, 99910, 99930, 99950, 99990, 100010, 100070, 100090, 100100, 
    100140, 100170, 100170, 100210, 100250, 100260, 100280, 100300, 100310, 
    100350, 100360, 100360, 100380, 100420, 100420, 100410, 100400, 100390, 
    100380, 100340, 100320, 100290, 100230, 100200, 100170, 100160, 100130, 
    100100, 100070, 100050, 100000, 99960, 99930, 99900, 99890, 99870, 99850, 
    99850, 99870, 99870, 99850, 99840, 99840, 99820, 99820, 99820, 99830, 
    99830, 99850, 99880, 99910, 99930, 99940, 99970, 99990, 100030, 100060, 
    100090, 100120, 100150, 100220, 100280, 100340, 100420, 100460, 100520, 
    100570, 100620, 100690, 100740, 100770, 100810, 100840, 100900, 100950, 
    101000, 101020, 101030, 101060, 101050, 101040, 101030, 101050, 101080, 
    101080, 101060, 101040, 101030, 100990, 100950, 100910, 100880, 100830, 
    100790, 100740, 100650, 100600, 100560, 100510, 100430, 100390, 100310, 
    100250, 100190, 100180, 100140, 100110, 100070, 100030, 100000, 99930, 
    99840, 99780, 99710, 99660, 99630, 99600, 99570, 99520, 99450, 99400, 
    99330, 99300, 99260, 99250, 99230, 99200, 99200, 99230, 99250, 99280, 
    99310, 99350, 99380, 99410, 99400, 99430, 99440, 99450, 99500, 99560, 
    99590, 99630, 99650, 99700, 99770, 99820, 99860, 99900, 99940, 99980, 
    100050, 100130, 100200, 100270, 100340, 100390, 100450, 100500, 100550, 
    100590, 100660, 100690, 100720, 100780, 100830, 100880, 100920, 100970, 
    101010, 101030, 101040, 101070, 101110, 101150, 101150, 101200, 101240, 
    101300, 101360, 101400, 101440, 101450, 101470, 101480, 101510, 101490, 
    101500, 101540, 101570, 101590, 101630, 101640, 101660, 101670, 101670, 
    101700, 101730, 101750, 101760, 101760, 101770, 101830, 101850, 101890, 
    101930, 101970, 101990, 102030, 102050, 102070, 102140, 102140, 102190, 
    102230, 102250, 102320, 102370, 102390, 102410, 102440, 102460, 102510, 
    102550, 102590, 102620, 102660, 102670, 102690, 102730, 102730, 102750, 
    102760, 102750, 102750, 102730, 102700, 102640, 102580, 102530, 102440, 
    102400, 102380, 102360, 102330, 102280, 102280, 102270, 102240, 102240, 
    102230, 102230, 102190, 102160, 102100, 101990, 101910, 101870, 101830, 
    101800, 101750, 101700, 101670, 101640, 101570, 101520, 101480, 101400, 
    101380, 101330, 101360, 101360, 101370, 101340, 101300, 101290, 101300, 
    101290, 101270, 101240, 101250, 101220, 101190, 101170, 101130, 101080, 
    101050, 100990, 101000, 100950, 100890, 100840, 100800, 100750, 100720, 
    100650, 100560, 100490, 100430, 100330, 100280, 100210, 100210, 100220, 
    100230, 100220, 100230, 100210, 100220, 100210, 100210, 100200, 100210, 
    100230, 100250, 100230, 100280, 100310, 100410, 100520, 100600, 100660, 
    100720, 100850, 101020, 101180, 101370, 101430, 101580, 101690, 101730, 
    101870, 101950, 101980, 102010, 102040, 102070, 102070, 102060, 102030, 
    101980, 101890, 101850, 101760, 101680, 101600, 101520, 101460, 101390, 
    101330, 101270, 101210, 101130, 101070, 101010, 100960, 100910, 100860, 
    100840, 100830, 100810, 100770, 100740, 100740, 100730, 100750, 100770, 
    100830, 100910, 100980, 101010, 101050, 101200, 101280, 101310, 101370, 
    101400, 101440, 101470, 101530, 101570, 101600, 101610, 101650, 101690, 
    101710, 101740, 101770, 101760, 101750, 101720, 101680, 101620, 101710, 
    101760, 101810, 101880, 101930, 101910, 101940, 101960, 102010, 102060, 
    102060, 102050, 102070, 102080, 102090, 102090, 102090, 102080, 102080, 
    102070, 102040, 102020, 102000, 101990, 101990, 101980, 101990, 101970, 
    101960, 101920, 101920, 101910, 101860, 101840, 101810, 101780, 101770, 
    101760, 101760, 101740, 101710, 101710, 101660, 101620, 101600, 101570, 
    101530, 101520, 101500, 101450, 101420, 101390, 101360, 101350, 101320, 
    101280, 101220, 101150, 101120, 101070, 100960, 100910, 100860, 100810, 
    100750, 100740, 100680, 100670, 100620, 100590, 100580, 100520, 100510, 
    100480, 100480, 100510, 100640, 100630, 100650, 100680, 100720, 100720, 
    100750, 100780, 100790, 100820, 100880, 100940, 100990, 101040, 101110, 
    101150, 101180, 101220, 101270, 101320, 101380, 101420, 101480, 101540, 
    101620, 101670, 101750, 101780, 101820, 101850, 101880, 101910, 101940, 
    102020, 102090, 102140, 102190, 102250, 102310, 102360, 102410, 102440, 
    102520, 102570, 102620, 102650, 102690, 102750, 102830, 102880, 102910, 
    102940, 102960, 102980, 103000, 103010, 103030, 103060, 103080, 103110, 
    103130, 103140, 103150, 103180, 103170, 103160, 103160, 103160, 103150, 
    103130, 103130, 103160, 103160, 103130, 103120, 103100, 103090, 103060, 
    103000, 102980, 102930, 102870, 102860, 102820, 102800, 102770, 102730, 
    102680, 102670, 102630, 102580, 102510, 102460, 102440, 102400, 102400, 
    102340, 102310, 102250, 102160, 102090, 102040, 101990, 101910, 101860, 
    101810, 101770, 101720, 101680, 101630, 101560, 101490, 101420, 101360, 
    101330, 101230, 101180, 101110, 101050, 101060, 100970, 100940, 100900, 
    100820, 100770, 100700, 100620, 100600, 100500, 100450, 100380, 100350, 
    100320, 100280, 100240, 100160, 100150, 100170, 100160, 100120, 100110, 
    100130, 100160, 100210, 100240, 100260, 100180, 100170, 100220, 100230, 
    100160, 100100, 100080, 100020, 100060, 100040, 100050, 100080, 100060, 
    100030, 99960, 99940, 99910, 99850, 99800, 99780, 99740, 99680, 99570, 
    99560, 99470, 99420, 99320, 99260, 99060, 99080, 99150, 99250, 99270, 
    99340, 99510, 99700, 99840, 99930, 100050, 100200, 100280, 100400, 
    100500, 100590, 100670, 100710, 100780, 100830, 100880, 100900, 100950, 
    101000, 101050, 101090, 101140, 101190, 101260, 101290, 101340, 101390, 
    101410, 101420, 101420, 101450, 101470, 101460, 101470, 101400, 101400, 
    101390, 101370, 101280, 101220, 101160, 101050, 100960, 100900, 100850, 
    100800, 100750, 100660, 100620, 100580, 100490, 100430, 100370, 100310, 
    100290, 100330, 100270, 100300, 100320, 100370, 100390, 100450, 100480, 
    100490, 100510, 100540, 100550, 100570, 100620, 100640, 100680, 100700, 
    100780, 100810, 100850, 100900, 100940, 100970, 101040, 101100, 101180, 
    101240, 101310, 101400, 101470, 101520, 101500, 101560, 101580, 101640, 
    101650, 101700, 101740, 101760, 101760, 101800, 101830, 101850, 101880, 
    101910, 101910, 101930, 101990, 102040, 102080, 102090, 102100, 102140, 
    102220, 102240, 102360, 102440, 102440, 102430, 102530, 102520, 102510, 
    102400, 102400, 102430, 102330, 102320, 102190, 102080, 101930, 101820, 
    101710, 101570, 101430, 101260, 101110, 100960, 100900, 100730, 100650, 
    100560, 100460, 100430, 100370, 100370, 100320, 100300, 100190, 100110, 
    99980, 99920, 99750, 99590, 99390, 99260, 99120, 98960, 98870, 98810, 
    98840, 98830, 98860, 98970, 98940, 98930, 98960, 98940, 98910, 98870, 
    99130, 99550, 99880, 100140, 100340, 100580, 100780, 100970, 101080, 
    101140, 101210, 101280, 101390, 101420, 101430, 101470, 101540, 101580, 
    101670, 101770, 101890, 101900, 101860, 101830, 101810, 101760, 101760, 
    101880, 101830, 101770, 101750, 101690, 101650, 101580, 101520, 101460, 
    101420, 101370, 101340, 101330, 101290, 101240, 101250, 101240, 101250, 
    101200, 101250, 101310, 101380, 101470, 101510, 101590, 101640, 101630, 
    101650, 101660, 101690, 101700, 101690, 101680, 101640, 101630, 101620, 
    101580, 101540, 101500, 101470, 101440, 101340, 101290, 101220, 101150, 
    101080, 100990, 100890, 100840, 100790, 100690, 100620, 100540, 100440, 
    100400, 100350, 100320, 100280, 100290, 100290, 100280, 100320, 100360, 
    100380, 100420, 100460, 100480, 100480, 100530, 100540, 100560, 100560, 
    100580, 100600, 100630, 100640, 100620, 100630, 100660, 100670, 100670, 
    100660, 100690, 100710, 100710, 100730, 100760, 100780, 100810, 100820, 
    100850, 100870, 100870, 100900, 100890, 100910, 100930, 100950, 100990, 
    101020, 101050, 101050, 101060, 101070, 101080, 101080, 101090, 101150, 
    101180, 101210, 101240, 101260, 101250, 101250, 101250, 101250, 101260, 
    101270, 101280, 101280, 101300, 101310, 101320, 101330, 101330, 101330, 
    101370, 101400, 101420, 101420, 101440, 101480, 101520, 101540, 101550, 
    101570, 101550, 101570, 101560, 101550, 101550, 101520, 101520, 101520, 
    101500, 101500, 101520, 101510, 101490, 101450, 101410, 101390, 101360, 
    101320, 101270, 101250, 101220, 101190, 101160, 101120, 101070, 101000, 
    100940, 100860, 100830, 100720, 100690, 100620, 100540, 100510, 100420, 
    100340, 100320, 100220, 100200, 100180, 100170, 100160, 100120, 100130, 
    100230, 100300, 100330, 100220, 100260, 100270, 100430, 100410, 100430, 
    100440, 100430, 100470, 100520, 100570, 100620, 100600, 100600, 100640, 
    100610, 100590, 100610, 100640, 100630, 100620, 100590, 100620, 100650, 
    100680, 100650, 100620, 100590, 100610, 100560, 100550, 100530, 100410, 
    100420, 100600, 100670, 100660, 100690, 100610, 100610, 100520, 100580, 
    100570, 100630, 100670, 100690, 100820, 100920, 101000, 101070, 101160, 
    101090, 101100, 101140, 101090, 101090, 101070, 101150, 101160, 101160, 
    101140, 101160, 101120, 101100, 101080, 101060, 101020, 101030, 101050, 
    101020, 101040, 101030, 101040, 101030, 100990, 100980, 100950, 100920, 
    100870, 100840, 100760, 100700, 100660, 100610, 100540, 100400, 100220, 
    100180, 100110, 100110, 100020, 99960, 99820, 99880, 99850, 99820, 99810, 
    99790, 99770, 99730, 99670, 99600, 99520, 99530, 99560, 99580, 99570, 
    99610, 99670, 99680, 99690, 99700, 99730, 99750, 99740, 99750, 99760, 
    99790, 99790, 99820, 99830, 99830, 99850, 99780, 99750, 99730, 99650, 
    99670, 99620, 99600, 99590, 99550, 99590, 99620, 99630, 99560, 99510, 
    99570, 99560, 99570, 99560, 99560, 99550, 99530, 99550, 99520, 99530, 
    99480, 99530, 99580, 99590, 99620, 99620, 99670, 99680, 99720, 99720, 
    99710, 99680, 99620, 99570, 99550, 99520, 99480, 99470, 99470, 99460, 
    99460, 99440, 99410, 99370, 99360, 99350, 99320, 99290, 99270, 99270, 
    99230, 99220, 99240, 99290, 99320, 99380, 99410, 99440, 99450, 99460, 
    99470, 99490, 99530, 99570, 99600, 99620, 99620, 99620, 99620, 99610, 
    99600, 99580, 99580, 99550, 99500, 99490, 99500, 99460, 99520, 99500, 
    99450, 99440, 99360, 99270, 99250, 99270, 99220, 99180, 99200, 99180, 
    99190, 99180, 99110, 99080, 99050, 99060, 99150, 99050, 99020, 99020, 
    99050, 99020, 99020, 99050, 99010, 98990, 98980, 98960, 98940, 98930, 
    98910, 98910, 98900, 98920, 98920, 98910, 98910, 98920, 98940, 98950, 
    98950, 98960, 98980, 99000, 99030, 99040, 99040, 99040, 99040, 99060, 
    99080, 99110, 99160, 99190, 99220, 99280, 99320, 99350, 99390, 99410, 
    99440, 99490, 99520, 99560, 99600, 99610, 99650, 99680, 99720, 99780, 
    99810, 99830, 99880, 99930, 99980, 100040, 100090, 100150, 100220, 
    100340, 100400, 100460, 100520, 100540, 100530, 100500, 100490, 100460, 
    100430, 100400, 100340, 100280, 100280, 100250, 100310, 100310, 100270, 
    100270, 100290, 100260, 100200, 100130, 100030, 99940, 99820, 99730, 
    99610, 99440, 99330, 99220, 99130, 99140, 99240, 99290, 99390, 99550, 
    99640, 99700, 99830, 99950, 100020, 100030, 100040, 100040, 100090, 
    100150, 100220, 100280, 100340, 100410, 100420, 100420, 100430, 100400, 
    100360, 100290, 100200, 100070, 99990, 99920, 99830, 99740, 99650, 99500, 
    99350, 99200, 99090, 98950, 98870, 98780, 98740, 98740, 98810, 98870, 
    98940, 98990, 99070, 99120, 99150, 99170, 99180, 99180, 99200, 99240, 
    99220, 99220, 99230, 99260, 99310, 99390, 99480, 99580, 99640, 99740, 
    99810, 99890, 99950, 100000, 100060, 100060, 100050, 100030, 100010, 
    99990, 99960, 99960, 99960, 99930, 99920, 99910, 99830, 99740, 99630, 
    99520, 99490, 99390, 99330, 99260, 99230, 99180, 99120, 99100, 99110, 
    99120, 99110, 99120, 99120, 99140, 99090, 99060, 99010, 98990, 98900, 
    98870, 98990, 99090, 99200, 99270, 99350, 99440, 99520, 99570, 99640, 
    99580, 99700, 99740, 99690, 99700, 99660, 99560, 99480, 99450, 99410, 
    99370, 99380, 99380, 99400, 99440, 99460, 99560, 99570, 99710, 99820, 
    99900, 100060, 100120, 100240, 100400, 100550, 100650, 100730, 100880, 
    101000, 101100, 101220, 101360, 101480, 101580, 101690, 101800, 101950, 
    101980, 102040, 102110, 102140, 102190, 102200, 102220, 102230, 102240, 
    102240, 102260, 102260, 102260, 102260, 102290, 102260, 102240, 102140, 
    102060, 101970, 101920, 101810, 101680, 101560, 101480, 101380, 101280, 
    101190, 101130, 101060, 101010, 100960, 100930, 100860, 100840, 100840, 
    100810, 100780, 100770, 100790, 100780, 100770, 100780, 100810, 100740, 
    100740, 100780, 100770, 100800, 100820, 100860, 100850, 100910, 100960, 
    100990, 101020, 101020, 101040, 101070, 101100, 101150, 101200, 101170, 
    101210, 101210, 101230, 101190, 101190, 101160, 101150, 101130, 101110, 
    101050, 100990, 100950, 100910, 100870, 100840, 100810, 100770, 100720, 
    100690, 100640, 100600, 100560, 100520, 100470, 100410, 100370, 100320, 
    100270, 100210, 100170, 100120, 100100, 100060, 100000, 99920, 99860, 
    99790, 99720, 99710, 99670, 99650, 99620, 99560, 99500, 99440, 99330, 
    99210, 99010, 98830, 98570, 98490, 98290, 98060, 98050, 98030, 97950, 
    97890, 97820, 97770, 97760, 97820, 97860, 97900, 98000, 98100, 98290, 
    98450, 98580, 98760, 98920, 99060, 99110, 99210, 99300, 99380, 99470, 
    99560, 99660, 99750, 99770, 99820, 99890, 99910, 99970, 100030, 100030, 
    100040, 100030, 99990, 99960, 99900, 99900, 99870, 99890, 99920, 99930, 
    99900, 99960, 99910, 99900, 99920, 99910, 99900, 99920, 99960, 99950, 
    100020, 100030, 100030, 100040, 100050, 100060, 100090, 100100, 100130, 
    100150, 100180, 100190, 100190, 100210, 100220, 100220, 100210, 100210, 
    100170, 100170, 100110, 100120, 100110, 100100, 100050, 100040, 100030, 
    99990, 99960, 99930, 99900, 99890, 99870, 99860, 99830, 99820, 99760, 
    99750, 99760, 99750, 99710, 99670, 99680, 99680, 99650, 99620, 99640, 
    99640, 99640, 99670, 99680, 99730, 99780, 99810, 99780, 99710, 99740, 
    99750, 99800, 99820, 99840, 99860, 99870, 99890, 99950, 99970, 99990, 
    100010, 100080, 100070, 100080, 100100, 100050, 100020, 99980, 99990, 
    99960, 99930, 99900, 99840, 99820, 99770, 99740, 99690, 99640, 99570, 
    99500, 99430, 99370, 99320, 99250, 99190, 99140, 99100, 99060, 99010, 
    98980, 98940, 98910, 98910, 98920, 98950, 98930, 98950, 98960, 99000, 
    99010, 99060, 99090, 99100, 99080, 99010, 98970, 98940, 98960, 98970, 
    99000, 99010, 99040, 99060, 99120, 99160, 99220, 99380, 99490, 99530, 
    99540, 99590, 99620, 99630, 99740, 99830, 99850, 99900, 99920, 99980, 
    99980, 99980, 99960, 99930, 99930, 99960, 100010, 100070, 100080, 100130, 
    100180, 100190, 100200, 100180, 100140, 100120, 100100, 100090, 100070, 
    100030, 100020, 100000, 99970, 99950, 99900, 99880, 99850, 99840, 99820, 
    99800, 99800, 99810, 99800, 99780, 99750, 99750, 99790, 99810, 99840, 
    99840, 99880, 99940, 100000, 100020, 100040, 100090, 100120, 100190, 
    100240, 100250, 100220, 100240, 100290, 100330, 100400, 100500, 100580, 
    100620, 100660, 100690, 100740, 100790, 100840, 100870, 100930, 100990, 
    101060, 101140, 101190, 101220, 101240, 101210, 101210, 101240, 101330, 
    101340, 101330, 101290, 101280, 101240, 101180, 101100, 101040, 100980, 
    100910, 100810, 100770, 100700, 100660, 100630, 100590, 100540, 100530, 
    100510, 100490, 100500, 100510, 100470, 100470, 100470, 100450, 100440, 
    100410, 100390, 100360, 100330, 100340, 100310, 100310, 100300, 100330, 
    100370, 100410, 100440, 100510, 100530, 100580, 100610, 100690, 100730, 
    100720, 100750, 100730, 100720, 100730, 100780, 100800, 100820, 100800, 
    100790, 100830, 100840, 100850, 100860, 100880, 100880, 100880, 100870, 
    100850, 100880, 100880, 100830, 100850, 100810, 100790, 100810, 100760, 
    100740, 100680, 100660, 100620, 100650, 100660, 100630, 100620, 100670, 
    100640, 100690, 100700, 100740, 100680, 100710, 100730, 100740, 100740, 
    100720, 100730, 100720, 100680, 100680, 100680, 100590, 100630, 100660, 
    100650, 100630, 100650, 100630, 100600, 100600, 100550, 100580, 100580, 
    100520, 100600, 100620, 100600, 100630, 100650, 100690, 100720, 100780, 
    100790, 100830, 100990, 101070, 101210, 101230, 101120, 101100, 101140, 
    101360, 101440, 101500, 101550, 101560, 101550, 101550, 101560, 101600, 
    101620, 101630, 101640, 101630, 101630, 101620, 101610, 101600, 101590, 
    101550, 101510, 101460, 101390, 101320, 101290, 101240, 101170, 101080, 
    100990, 100910, 100810, 100740, 100700, 100660, 100620, 100580, 100540, 
    100480, 100410, 100380, 100320, 100320, 100260, 100220, 100170, 100140, 
    100070, 100000, 99970, 99950, 99980, 99900, 99810, 99760, 99920, 99900, 
    99820, 99860, 99860, 99850, 99750, 99600, 99590, 99540, 99440, 99230, 
    99310, 99490, 99630, 99970, 100110, 100190, 100240, 100180, 100170, 
    100140, 100130, 100070, 100140, 100110, 100100, 100060, 100150, 100190, 
    100090, 100070, 100300, 100400, 100410, 100370, 100400, 100320, 100290, 
    100260, 100250, 100270, 100370, 100350, 100290, 100300, 100300, 100290, 
    100240, 100210, 100180, 100140, 100100, 100070, 100050, 99980, 99900, 
    99840, 99790, 99740, 99680, 99580, 99590, 99560, 99560, 99570, 99540, 
    99470, 99470, 99430, 99270, 99220, 99290, 99350, 99330, 99360, 99420, 
    99460, 99450, 99440, 99430, 99430, 99450, 99410, 99430, 99430, 99440, 
    99460, 99470, 99500, 99500, 99510, 99520, 99570, 99600, 99630, 99670, 
    99670, 99710, 99750, 99790, 99810, 99820, 99870, 99890, 99930, 99960, 
    99990, 100010, 100030, 100000, 100050, 100100, 100070, 100090, 100110, 
    100140, 100150, 100150, 100140, 100120, 100090, 100090, 100100, 100130, 
    100160, 100150, 100160, 100140, 100150, 100160, 100180, 100180, 100160, 
    100160, 100160, 100160, 100170, 100170, 100170, 100200, 100140, 100160, 
    100190, 100190, 100190, 100120, 100070, 100050, 100120, 100140, 100250, 
    100250, 100240, 100210, 100120, 100300, 100310, 100270, 100310, 100340, 
    100350, 100370, 100360, 100350, 100320, 100330, 100330, 100340, 100340, 
    100330, 100340, 100370, 100390, 100380, 100360, 100360, 100350, 100350, 
    100400, 100370, 100370, 100370, 100350, 100330, 100320, 100310, 100320, 
    100280, 100270, 100260, 100250, 100230, 100190, 100160, 100150, 100140, 
    100140, 100130, 100170, 100120, 100100, _, 100030, 100020, 100000, 
    100000, 99940, 99950, 99980, 99960, 99910, 99970, 99930, 99950, 99960, 
    99960, 99970, 99960, 100000, 100030, 100080, 100070, 100100, 100110, 
    100140, 100160, 100190, 100240, _, 100280, _, 100340, 100400, 100430, 
    100520, 100560, 100610, 100630, 100620, 100680, 100710, 100710, 100770, 
    100820, 100870, 100890, _, 100960, 100980, 101030, 101060, 101090, 
    101090, 101130, 101180, 101210, 101250, 101270, 101320, 101360, 101390, 
    101390, 101420, 101440, 101510, 101550, 101610, 101640, 101650, 101660, 
    101650, 101660, 101690, 101720, 101760, 101790, 101800, 101810, 101830, 
    101820, 101900, 101940, 101970, 101990, 101990, 102020, 102040, 102050, 
    102090, 102120, 102140, 102210, 102250, 102250, 102300, 102350, 102360, 
    102370, 102410, 102420, 102460, 102470, 102500, 102530, 102560, 102590, 
    102580, 102590, 102580, 102600, 102600, 102610, 102620, 102630, 102640, 
    102660, 102650, 102630, 102610, 102600, 102590, 102580, 102550, 102540, 
    102520, 102520, 102490, 102460, 102450, 102430, 102420, 102410, 102400, 
    102380, 102370, 102360, 102340, 102350, 102360, 102360, 102330, 102330, 
    102320, 102320, 102310, 102300, 102300, 102280, 102280, 102290, 102290, 
    102300, 102300, 102280, 102230, 102190, 102210, 102190, 102140, 102170, 
    102130, 102120, 102120, 102120, 102110, 102090, 102070, 102040, 102010, 
    102020, 102010, 102020, 102030, 102010, 102020, 102020, 102050, 102030, 
    102060, 102070, 102100, 102080, 102060, 102030, 102040, 102030, 101960, 
    101930, 101950, 101940, 101900, 101870, 101830, 101800, 101780, 101800, 
    101770, 101740, 101700, 101670, 101660, 101620, 101590, 101560, 101540, 
    101490, 101470, 101430, 101380, 101350, 101340, 101380, 101370, 101370, 
    101370, 101370, 101400, 101390, 101390, 101390, 101410, 101430, 101450, 
    101500, 101530, 101550, 101570, 101570, 101590, 101600, 101620, 101620, 
    101610, 101620, 101640, 101660, 101690, 101680, 101700, 101700, 101720, 
    101760, 101800, 101820, 101850, 101870, 101920, 101940, 101960, 101990, 
    102000, 101980, 101980, 102000, 102000, 102020, _, 102040, 102070, 
    102110, 102130, 102120, _, 102110, 102090, 102080, 102050, 102020, 
    101980, 101960, 101920, 101930, 101890, 101860, 101840, 101820, 101830, 
    101800, 101800, 101770, 101770, 101770, 101780, 101790, 101790, 101800, 
    101820, 101780, 101740, 101720, 101720, 101700, 101690, 101660, 101660, 
    101650, 101650, 101670, 101620, 101610, 101600, 101600, 101620, 101630, 
    101650, 101700, 101770, 101850, 101930, 101990, 102060, 102120, 102160, 
    102220, 102270, 102310, 102380, 102440, 102480, 102540, 102580, 102630, 
    102650, 102670, 102690, 102720, 102740, 102770, 102790, 102840, 102860, 
    102900, 102930, 102970, 102990, 103000, 103010, 103020, 103040, 103040, 
    103090, 103110, 103120, 103140, 103170, 103180, 103170, 103170, 103170, 
    103180, 103190, 103190, 103180, 103200, 103230, 103240, 103260, 103280, 
    103270, 103250, 103240, 103230, 103210, 103190, 103170, 103160, 103140, 
    103100, 103070, 103040, 103010, 102950, 102880, 102850, 102820, 102790, 
    102720, 102720, 102730, 102740, 102730, 102730, 102710, 102690, 102680, 
    102670, 102640, 102650, 102640, 102640, 102630, 102670, 102640, 102630, 
    102620, 102600, 102580, 102530, 102490, 102470, 102420, 102410, 102350, 
    102400, 102380, 102390, 102410, 102370, 102360, 102310, 102290, 102270, 
    102250, 102210, 102200, 102210, 102200, 102190, 102160, 102160, 102140, 
    102160, 102150, 102150, 102160, 102160, 102190, 102210, 102240, 102260, 
    102270, 102280, 102280, 102300, 102310, 102300, 102300, 102330, 102330, 
    102320, 102300, 102310, 102290, 102280, 102270, 102240, 102220, 102200, 
    102180, 102170, 102170, 102160, 102120, 102090, 102030, 101990, 101940, 
    101910, 101880, 101840, 101790, 101750, 101760, 101710, 101670, 101620, 
    101580, 101530, 101490, 101460, 101440, 101410, 101380, 101350, 101330, 
    101320, 101290, 101260, 101280, 101240, 101200, 101180, 101140, 101130, 
    101100, 101080, 101070, 101030, 101010, 100970, 100890, 100880, 100860, 
    100840, 100830, 100810, 100790, 100800, 100800, 100800, 100800, 100740, 
    100710, 100710, 100640, 100620, 100590, 100580, 100650, 100670, 100620, 
    100610, 100560, 100490, 100510, 100480, 100430, 100390, 100310, 100230, 
    100210, 100170, 100140, 100170, 100160, 100120, 100120, 100090, 100110, 
    100100, 100150, 100140, 100110, 100080, 100050, 100040, 100070, 100090, 
    100130, 100100, 100020, 100010, 99970, 99940, 99920, 99870, 99810, 99810, 
    99850, 99850, 99900, 99940, 99960, 99930, 99950, 99990, 100020, 100030, 
    100020, 100030, 99970, 99930, 99910, 99960, 100010, 100060, 100100, 
    100120, 100170, 100210, 100260, 100310, 100350, 100370, 100390, 100410, 
    100410, 100450, 100480, 100500, 100510, 100510, 100550, 100580, 100570, 
    100590, 100600, 100610, 100620, 100640, 100630, 100630, 100600, 100580, 
    100570, 100540, 100520, 100480, 100460, 100470, 100470, 100460, 100460, 
    100450, 100420, 100420, 100390, 100360, 100320, 100300, 100260, 100230, 
    100230, 100180, 100140, 100110, 100080, 100080, 100100, 100100, 100050, 
    100030, 100010, 100000, 99970, 99970, 99940, 99890, 99860, 99830, 99810, 
    99790, 99770, 99780, 99760, 99720, 99710, 99680, 99670, 99640, 99620, 
    99600, 99610, 99590, 99580, 99550, 99510, 99460, 99430, 99440, 99420, 
    99430, 99400, 99400, 99420, 99430, 99450, 99490, 99520, 99550, 99630, 
    99630, 99670, 99690, 99750, 99770, 99810, 99890, 99900, 99940, 99960, 
    99980, 100030, 99990, 99980, 99930, 99910, 99910, 99920, 100060, 100150, 
    100230, 100230, 100230, 100270, 100300, 100260, 100260, 100250, 100220, 
    100240, 100280, 100280, 100290, 100290, 100290, 100280, 100260, 100240, 
    100230, 100210, 100220, 100270, 100320, 100350, 100340, 100380, 100410, 
    100420, 100430, 100420, 100440, 100460, 100490, 100520, 100580, 100630, 
    100670, 100710, 100770, 100770, 100740, 100780, 100810, 100840, 100850, 
    100860, 100870, 100890, 100930, 100840, 100810, 100800, 100850, 100810, 
    100760, 100820, 100860, 100830, 100870, 100850, 100820, 100770, 100750, 
    100720, 100700, 100660, 100670, 100620, 100550, 100510, 100430, 100320, 
    100330, 100310, 100290, 100190, 100130, 100090, 100050, 99970, 99920, 
    99880, 99860, 99830, 99800, 99780, 99760, 99720, 99660, 99610, 99540, 
    99540, 99500, 99460, 99440, 99440, 99450, 99470, 99490, 99510, 99520, 
    99570, 99610, 99620, 99670, 99710, 99780, 99850, 99870, 99890, 99910, 
    99920, 99990, 100000, 100010, 100030, 100040, 100050, 100070, 100100, 
    100140, 100170, 100190, 100200, 100250, 100270, 100300, 100390, 100400, 
    100420, 100480, 100530, 100570, 100520, 100570, 100540, 100500, 100420, 
    100300, 100150, 100020, 99860, 99760, 99650, 99530, 99410, 99290, 99200, 
    99060, 99010, 98940, 98900, 98910, 98870, 98820, 98780, 98700, 98570, 
    98450, 98390, 98290, 98200, 98080, 98070, 98060, 98030, 98060, 98080, 
    98110, 98110, 98170, 98220, 98270, 98370, 98420, 98540, 98600, 98730, 
    98840, 98930, 99010, 99140, 99210, 99300, 99350, 99510, 99520, 99590, 
    99620, 99690, 99680, 99740, 99730, 99740, 99750, 99670, 99680, 99680, 
    99630, 99560, 99520, 99510, 99520, 99540, 99550, 99540, 99540, 99610, 
    99680, 99700, 99850, 99980, 100120, 100210, 100260, 100330, 100410, 
    100520, 100600, 100730, 100820, 100870, 100850, 100900, 100900, 100930, 
    100930, 100980, 100980, 100970, 101000, 101000, 100970, 100960, 100920, 
    100860, 100860, 100850, 100820, 100860, 100860, 100820, 100820, 100830, 
    100750, 100780, 100790, 100780, 100780, 100830, 100820, 100880, 100880, 
    100820, 100870, 100870, 100870, 100880, 100780, 100730, 100660, 100700, 
    100680, 100650, 100680, 100660, 100650, 100630, 100570, 100570, 100610, 
    100590, 100590, 100520, 100450, 100580, 100570, 100530, 100510, 100510, 
    100530, 100520, 100460, 100260, 100200, 100320, 100360, 100380, 100300, 
    100280, 100230, 100260, 100260, 100200, 100210, 100260, 100290, 100430, 
    100520, 100540, 100570, 100620, 100680, 100720, 100730, 100830, 100800, 
    100830, 100830, 100860, 100880, 100950, 100920, 100920, 100900, 100910, 
    100930, 100920, 100840, 100810, 100750, 100620, _, 100520, 100470, 
    100400, 100370, 100350, 100270, 100210, 100150, 100040, 99940, 99920, 
    99840, 99870, 99760, 99650, 99630, 99580, 99570, 99530, 99480, 99420, 
    99430 ;

 air_temperature_2m = 250.65, 250.65, 250.35, 249.65, 249.45, 249.15, 248.65, 
    248.55, 248.45, 248.25, 248.25, 248.25, 248.35, 248.55, 248.95, 249.35, 
    249.85, 251.15, 251.45, 251.65, 252.05, 254.05, 255.05, 256.85, 257.65, 
    258.25, 258.85, 259.25, 260.15, 261.75, 261.95, 261.45, 261.15, 261.15, 
    261.25, 262.75, 263.25, 263.15, 262.05, 261.05, 260.55, 260.65, 262.25, 
    262.75, 263.95, 264.35, 264.95, 265.15, 265.25, 265.05, 264.85, 265.15, 
    265.55, 266.85, 266.35, 264.85, 264.45, 261.95, 260.85, 260.95, 258.95, 
    257.95, 256.85, 256.45, 256.45, 256.85, 258.25, 259.45, 260.05, 260.45, 
    260.85, 260.95, 260.95, 260.45, 259.75, 259.65, 259.65, 259.45, 258.95, 
    258.35, 258.25, 257.15, 254.45, 253.55, 252.75, 251.55, 250.85, 250.35, 
    249.35, 249.25, 249.35, 249.45, 249.55, 249.45, 249.35, 249.35, 249.35, 
    249.45, 249.45, 249.55, 249.55, 249.85, 250.15, 251.65, 252.35, 252.85, 
    253.85, 254.35, 254.65, 254.95, 254.85, 254.75, 254.75, 255.45, 256.05, 
    256.35, 256.75, 256.95, 257.25, 257.45, 257.35, 257.05, 256.75, 255.85, 
    255.45, 255.15, 254.75, 254.55, 253.85, 253.55, 253.15, 253.15, 252.85, 
    252.85, 252.85, 252.95, 252.95, 252.55, 252.45, 252.25, 252.05, 252.05, 
    252.15, 266.15, 256.45, 243.55, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 281.15, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 275.15, 275.15, 275.05, 275.45, 
    275.25, 275.15, 275.25, 275.35, 275.45, 275.25, 275.15, 275.15, 275.05, 
    275.05, 275.05, 274.85, 274.95, 274.85, 274.85, 274.85, 274.85, 274.85, 
    274.95, 275.05, 275.15, 275.25, 275.35, 274.65, 274.35, 274.55, 274.75, 
    274.65, 274.45, 274.25, 273.75, 273.45, 273.45, 273.35, 273.15, 273.15, 
    273.35, 273.55, 273.65, 273.65, 273.55, 273.55, 273.85, 273.95, 273.85, 
    273.85, 274.15, 274.15, 274.05, 274.35, 273.85, 274.05, 274.15, 273.85, 
    273.65, 273.45, 273.35, 273.35, 273.15, 273.25, 273.25, 273.65, 273.75, 
    273.85, 273.75, 273.85, 273.75, 273.85, 274.45, 274.65, 274.75, 274.85, 
    275.05, 274.65, 274.35, 274.45, 274.25, 273.95, 274.25, 273.95, 273.65, 
    274.25, 274.85, 274.95, 274.75, 274.45, 274.75, 274.85, 274.75, 274.55, 
    274.55, 274.45, 274.65, 274.65, 274.65, 274.55, 275.05, 274.85, 275.65, 
    275.35, 275.75, 275.75, 275.75, 275.75, 275.95, 275.55, 275.25, 274.65, 
    274.35, 274.05, 273.65, 273.85, 274.05, 274.15, 274.15, 274.65, 274.65, 
    274.25, 274.35, 273.95, 273.95, 273.75, 273.35, 272.85, 272.55, 272.55, 
    272.65, 273.15, 274.05, 274.25, 274.35, 274.65, 274.85, 275.35, 274.75, 
    274.85, 275.35, 275.65, 276.05, 276.15, 276.05, 274.85, 275.95, 275.75, 
    275.65, 275.65, 275.75, 275.15, 275.25, 275.35, 274.85, 274.65, 275.05, 
    275.35, 274.85, 276.05, 275.95, 275.95, 276.05, 276.95, 276.95, 276.95, 
    276.85, 277.05, 276.45, 276.65, 276.85, 276.65, 276.05, 276.25, 276.25, 
    276.25, 276.25, 276.15, 276.25, 275.85, 275.95, 275.65, 275.75, 275.75, 
    275.15, 275.35, 274.85, 275.55, 274.15, 274.15, 274.55, 274.55, 274.55, 
    274.05, 274.05, 274.15, 273.25, 272.45, 272.35, 271.95, 271.55, 271.25, 
    270.85, 270.65, 270.55, 270.65, 271.05, 271.45, 271.85, 272.25, 272.65, 
    273.45, 273.55, 273.45, 274.85, 274.85, 275.55, 273.15, 273.15, 272.35, 
    272.85, 272.05, 272.15, 272.45, 273.45, 272.15, 271.35, 271.75, 271.85, 
    271.95, 273.25, 272.55, 272.65, 274.15, 273.25, 273.45, 273.45, 273.45, 
    274.05, 274.65, 275.05, 275.45, 274.85, 274.65, 274.45, 274.35, 275.35, 
    274.65, 274.95, 275.25, 274.35, 273.65, 272.95, 272.35, 272.25, 272.55, 
    272.75, 272.75, 272.95, 273.65, 273.75, 273.75, 273.75, 273.75, 273.75, 
    273.75, 274.15, 274.15, 274.25, 273.75, 273.55, 273.15, 272.95, 272.45, 
    271.95, 272.15, 271.75, 271.15, 272.25, 271.45, 271.65, 271.95, 272.05, 
    271.85, 272.25, 272.35, 272.25, 272.45, 272.35, 272.75, 272.45, 272.75, 
    272.35, 272.25, 272.55, 271.85, 272.15, 272.45, 272.05, 271.85, 271.65, 
    271.75, 272.05, 272.05, 272.25, 272.35, 271.95, 272.25, 272.95, 272.45, 
    273.25, 273.05, 273.45, 273.35, 273.35, 273.55, 273.05, 273.15, 272.95, 
    272.85, 272.95, 272.85, 272.75, 272.55, 272.35, 272.45, 272.35, 272.05, 
    271.85, 272.15, 272.35, 272.45, 272.55, 272.05, 272.15, 272.25, 272.85, 
    272.65, 272.85, 273.15, 272.95, 272.95, 273.25, 273.25, 273.45, 273.95, 
    274.05, 274.05, 274.35, 274.35, 274.25, 274.25, 274.15, 273.95, 273.85, 
    274.05, 274.45, 274.75, 274.65, 274.65, 274.95, 275.25, 275.05, 274.95, 
    274.75, 275.15, 275.45, 275.45, 275.05, 275.05, 274.95, 274.95, 275.05, 
    275.15, 274.95, 274.95, 274.85, 274.95, 275.05, 274.85, 275.25, 275.55, 
    275.85, 275.95, 276.35, 276.25, 276.15, 276.65, 276.95, 276.55, 275.75, 
    275.35, 274.85, 274.65, 274.75, 274.55, 274.65, 274.55, 274.45, 274.55, 
    274.55, 274.65, 274.55, 274.45, 274.55, 274.95, 275.35, 275.65, 275.15, 
    274.85, 274.95, 275.25, 275.15, 275.55, 275.05, 274.25, 274.15, 273.85, 
    272.95, 272.45, 271.95, 271.55, 270.95, 270.85, 271.25, 271.15, 271.45, 
    271.65, 272.75, 272.15, 272.95, 272.55, 273.35, 273.55, 273.75, 274.35, 
    274.55, 274.85, 275.65, 275.75, 276.35, 275.45, 275.95, 276.35, 276.35, 
    275.55, 275.25, 276.25, 276.55, 276.75, 277.45, 277.05, 276.25, 275.25, 
    275.05, 274.85, 276.15, 276.25, 276.45, 276.15, 275.85, 275.95, 275.75, 
    275.35, 275.15, 275.35, 275.15, 275.35, 275.55, 276.55, 276.65, 275.75, 
    275.65, 275.65, 275.35, 275.15, 274.75, 274.45, 274.35, 273.35, 273.65, 
    273.55, 274.65, 276.35, 276.15, 275.95, 276.25, 276.05, 275.35, 275.45, 
    275.65, 275.35, 276.35, 275.25, 274.55, 275.25, 274.75, 274.65, 274.55, 
    274.15, 274.15, 275.05, 274.85, 274.95, 275.15, 275.15, 274.85, 275.15, 
    274.75, 274.45, 274.45, 274.35, 274.85, 275.25, 275.25, 275.75, 276.35, 
    276.35, 276.75, 276.65, 276.55, 276.25, 276.75, 276.65, 276.75, 277.35, 
    277.15, 276.75, 276.55, 276.75, 276.65, 277.05, 276.85, 276.85, 276.95, 
    276.45, 275.45, 275.35, 275.25, 275.05, 274.15, 274.35, 274.45, 275.05, 
    274.85, 274.55, 274.25, 274.05, 274.05, 274.05, 274.25, 274.05, 274.35, 
    274.55, 274.85, 274.65, 274.85, 274.55, 274.65, 274.65, 274.75, 274.55, 
    274.45, 274.35, 274.45, 274.45, 274.05, 274.05, 274.05, 274.45, 275.05, 
    275.75, 275.55, 276.35, 277.05, 276.95, 275.55, 276.05, 275.95, 276.35, 
    276.15, 275.65, 276.15, 278.45, 279.65, 277.65, 277.95, 277.75, 276.95, 
    276.35, 276.85, 276.75, 276.35, 275.85, 275.35, 275.15, 274.85, 275.35, 
    275.35, 275.25, 275.25, 275.05, 275.25, 275.15, 275.15, 274.95, 275.15, 
    275.35, 275.25, 275.35, 275.35, 275.55, 275.35, 275.55, 275.85, 276.05, 
    275.65, 275.55, 275.65, 275.65, 276.05, 276.05, 275.95, 276.15, 276.05, 
    276.05, 275.65, 275.35, 275.55, 274.35, 274.15, 273.85, 273.45, 273.25, 
    272.95, 272.75, 272.45, 271.85, 271.75, 271.45, 271.15, 270.95, 270.85, 
    270.35, 270.45, 270.35, 270.55, 270.35, 270.85, 270.35, 270.25, 270.35, 
    270.15, 270.15, 270.15, 270.15, 270.35, 270.35, 270.85, 270.85, 270.95, 
    271.75, 272.15, 272.75, 272.95, 273.05, 273.65, 274.45, 274.85, 274.85, 
    274.85, 275.35, 275.25, 275.95, 276.05, 276.75, 277.25, 276.35, 276.45, 
    276.35, 276.25, 276.35, 276.65, 276.55, 276.55, 276.45, 276.45, 276.75, 
    276.55, 277.05, 276.65, 276.35, 276.95, 276.55, 276.65, 275.95, 276.05, 
    276.55, 278.15, 276.55, 275.95, 275.85, 275.95, 277.35, 276.65, 277.05, 
    276.25, 276.45, 276.75, 277.45, 277.95, 278.15, 278.45, 278.15, 277.55, 
    278.05, 277.15, 279.05, 277.75, 279.35, 275.15, 275.95, 275.65, 275.45, 
    275.65, 275.25, 274.75, 275.15, 275.15, 274.35, 274.55, 274.45, 274.55, 
    274.65, 274.55, 274.75, 274.85, 274.75, 274.65, 274.65, 273.95, 273.85, 
    273.85, 273.65, 273.75, 273.95, 273.85, 273.75, 273.45, 273.35, 273.35, 
    273.15, 273.15, 273.05, 272.85, 272.75, 272.35, 272.15, 272.15, 272.05, 
    271.95, 271.85, 271.45, 271.35, 271.25, 270.95, 271.45, 271.95, 272.35, 
    272.65, 272.85, 272.75, 272.85, 273.05, 273.35, 273.35, 273.25, 273.05, 
    272.75, 272.95, 273.15, 273.35, 273.45, 273.55, 273.75, 273.75, 274.35, 
    274.45, 274.45, 275.05, 275.05, 274.95, 274.85, 275.05, 276.05, 275.25, 
    277.55, 277.05, 275.85, 275.15, 275.25, 274.95, 274.35, 274.15, 273.75, 
    273.65, 273.35, 273.75, 275.05, 274.75, 273.35, 272.95, 272.45, 273.35, 
    273.95, 274.25, 274.65, 274.75, 274.95, 274.65, 274.75, 274.75, 274.85, 
    274.35, 274.15, 274.05, 273.75, 273.95, 273.95, 273.55, 272.55, 273.35, 
    273.25, 273.35, 273.55, 273.65, 273.35, 272.95, 272.95, 272.95, 273.35, 
    273.55, 273.75, 273.65, 273.65, 273.75, 273.75, 273.65, 273.95, 274.55, 
    275.05, 275.25, 275.15, 275.05, 275.45, 275.15, 275.25, 275.05, 274.45, 
    274.45, 274.35, 274.35, 274.25, 274.45, 274.25, 274.25, 274.25, 274.05, 
    274.05, 273.85, 273.55, 273.25, 273.15, 272.85, 272.85, 272.75, 273.15, 
    273.65, 273.75, 274.05, 274.65, 274.75, 274.65, 274.65, 274.15, 273.15, 
    273.35, 273.25, 273.45, 273.55, 273.95, 274.55, 274.85, 275.15, 274.95, 
    275.45, 275.25, 275.25, 274.75, 275.05, 274.55, 274.55, 274.35, 274.25, 
    274.15, 273.75, 272.95, 272.65, 272.65, 272.75, 272.95, 273.05, 272.95, 
    273.25, 273.35, 272.65, 272.95, 275.15, 273.85, 274.05, 274.25, 274.25, 
    274.45, 274.35, 274.45, 273.85, 273.65, 273.35, 273.35, 273.55, 273.55, 
    273.75, 273.95, 274.35, 274.55, 274.35, 274.35, 274.55, 274.65, 275.15, 
    275.45, 275.45, 275.25, 275.35, 275.85, 275.95, 275.55, 275.25, 274.95, 
    275.05, 274.75, 274.95, 274.95, 275.25, 275.25, 274.95, 274.95, 274.85, 
    274.85, 274.95, 274.95, 274.85, 274.85, 274.85, 275.05, 274.75, 274.75, 
    274.95, 275.35, 275.15, 275.35, 275.05, 274.85, 274.55, 274.95, 274.65, 
    274.55, 275.45, 275.55, 275.75, 275.55, 275.35, 274.95, 274.85, 275.05, 
    275.45, 274.95, 274.75, 275.35, 275.35, 275.25, 275.55, 275.75, 275.65, 
    275.55, 275.55, 276.05, 276.45, 276.05, 276.05, 276.15, 276.45, 276.05, 
    275.55, 275.85, 275.35, 275.15, 275.15, 275.45, 275.15, 275.15, 275.55, 
    275.65, 275.75, 275.85, 276.15, 275.95, 275.35, 274.85, 274.95, 274.75, 
    275.05, 275.25, 275.25, 275.45, 275.25, 276.05, 275.55, 275.35, 275.15, 
    275.15, 274.55, 274.55, 274.35, 274.35, 274.15, 274.05, 274.05, 273.85, 
    273.75, 273.35, 272.95, 272.65, 272.45, 272.05, 271.85, 271.25, 270.65, 
    269.75, 268.85, 268.75, 268.95, 268.75, 268.95, 268.55, 268.55, 268.75, 
    269.35, 269.05, 268.15, 268.25, 268.15, 267.95, 268.05, 267.95, 267.95, 
    267.95, 268.15, 268.55, 268.75, 269.45, 269.65, 269.95, 270.15, 270.55, 
    271.05, 270.85, 271.15, 271.25, 271.15, 271.15, 271.05, 271.15, 271.05, 
    271.05, 270.95, 270.85, 270.95, 270.55, 271.05, 271.45, 271.55, 271.75, 
    271.85, 271.65, 271.65, 272.15, 272.45, 272.35, 272.45, 272.45, 272.45, 
    272.75, 272.55, 272.25, 271.85, 271.65, 271.25, 270.95, 271.25, 271.05, 
    270.45, 270.35, 270.45, 270.45, 269.45, 268.85, 268.65, 268.55, 268.15, 
    268.25, 267.85, 267.85, 268.05, 268.25, 268.55, 268.65, 268.95, 269.45, 
    269.45, 269.35, 269.25, 268.95, 268.55, 268.05, 267.85, 267.65, 267.65, 
    267.75, 267.75, 267.95, 267.85, 267.65, 266.65, 266.95, 267.95, 269.05, 
    269.65, 270.35, 270.85, 270.95, 270.85, 270.55, 270.95, 270.35, 269.95, 
    270.05, 269.95, 269.95, 268.45, 269.55, 269.85, 270.05, 269.75, 269.15, 
    268.95, 270.15, 270.05, 270.15, 270.25, 270.45, 270.45, 270.35, 270.05, 
    270.15, 270.35, 270.45, 270.65, 270.15, 270.15, 270.35, 270.45, 270.35, 
    270.45, 269.65, 269.85, 269.85, 268.65, 269.55, 269.05, 269.15, 269.25, 
    268.75, 268.25, 268.55, 268.75, 269.25, 269.85, 270.45, 270.65, 270.75, 
    270.55, 270.25, 269.45, 268.95, 269.25, 269.05, 268.35, 269.35, 268.65, 
    268.85, 269.65, 269.75, 269.65, 269.55, 269.45, 269.35, 269.15, 268.95, 
    268.95, 268.45, 268.35, 269.45, 269.25, 269.35, 269.35, 269.35, 269.35, 
    269.35, 268.85, 268.05, 267.55, 266.95, 266.05, 265.65, 265.25, 264.85, 
    264.55, 264.25, 263.65, 263.55, 263.55, 263.45, 263.35, 262.15, 261.35, 
    261.05, 261.25, 261.85, 262.65, 263.45, 265.25, 266.05, 265.95, 265.25, 
    264.75, 264.55, 264.35, 263.45, 263.35, 262.85, 262.95, 262.95, 262.65, 
    261.85, 262.05, 261.75, 261.75, 261.35, 261.25, 261.15, 261.45, 261.65, 
    261.35, 261.75, 262.05, 262.45, 262.95, 263.75, 264.35, 264.65, 265.15, 
    265.65, 266.05, 266.55, 266.85, 267.25, 267.65, 267.85, 268.05, 268.05, 
    268.15, 268.25, 268.55, 268.55, 268.25, 267.95, 268.45, 268.95, 269.25, 
    269.15, 268.95, 268.85, 268.55, 268.65, 268.55, 269.05, 268.25, 268.35, 
    268.35, 268.25, 267.95, 268.05, 267.95, 267.95, 267.85, 267.75, 267.95, 
    267.95, 267.65, 267.95, 268.25, 268.15, 268.25, 268.35, 268.25, 268.25, 
    268.35, 268.35, 268.55, 268.55, 268.65, 268.75, 268.75, 268.75, 268.75, 
    269.05, 269.35, 269.35, 269.35, 269.85, 269.85, 269.85, 269.85, 270.35, 
    270.75, 270.65, 269.85, 270.35, 269.95, 269.75, 269.75, 268.95, 268.95, 
    268.95, 268.95, 269.15, 268.85, 268.45, 268.35, 268.15, 268.25, 268.05, 
    267.95, 267.85, 267.45, 267.65, 267.45, 267.25, 267.35, 267.25, 267.45, 
    267.35, 267.65, 267.55, 267.75, 268.15, 268.35, 268.45, 268.75, 268.25, 
    268.75, 267.95, 267.85, 268.25, 268.05, 267.55, 267.05, 267.05, 266.95, 
    267.15, 267.05, 267.45, 267.45, 267.25, 267.15, 266.95, 266.55, 266.15, 
    266.95, 267.55, 268.15, 268.45, 268.55, 269.15, 269.05, 269.65, 270.25, 
    270.85, 271.05, 271.55, 271.75, 271.85, 272.05, 272.45, 273.15, 272.15, 
    272.45, 272.65, 272.65, 272.85, 272.85, 272.45, 272.45, 272.15, 271.75, 
    271.65, 271.95, 272.15, 271.85, 271.65, 271.85, 271.85, 272.05, 271.95, 
    271.75, 271.95, 272.05, 271.85, 271.55, 271.35, 270.95, 270.65, 270.75, 
    270.85, 270.85, 270.75, 270.65, 270.75, 270.85, 270.75, 270.55, 270.55, 
    270.45, 270.35, 270.15, 270.05, 269.85, 269.55, 269.45, 269.25, 269.15, 
    269.15, 269.75, 269.75, 270.35, 270.65, 271.05, 270.95, 270.75, 270.55, 
    270.35, 270.05, 269.75, 269.35, 269.15, 269.15, 268.85, 268.85, 268.65, 
    268.65, 268.65, 268.55, 268.15, 268.15, 267.95, 267.85, 267.95, 267.95, 
    268.15, 268.15, 268.45, 268.45, 268.35, 268.25, 268.55, 268.75, 269.25, 
    269.65, 269.75, 269.75, 269.65, 269.55, 269.35, 269.15, 269.05, 269.55, 
    269.85, 270.05, 269.85, 270.25, 270.15, 270.05, 270.55, 270.55, 270.85, 
    270.85, 270.55, 270.05, 270.25, 270.65, 270.65, 270.65, 270.65, 270.75, 
    270.55, 270.15, 270.35, 270.75, 271.05, 271.35, 271.55, 271.55, 271.25, 
    271.15, 271.35, 271.25, 271.25, 271.15, 270.85, 271.05, 271.15, 271.25, 
    271.35, 271.15, 271.25, 271.25, 271.55, 271.45, 271.45, 271.25, 270.95, 
    270.75, 270.35, 270.05, 269.85, 269.65, 269.65, 269.55, 269.45, 269.25, 
    269.25, 268.75, 268.55, 268.55, 268.25, 268.65, 268.55, 268.65, 268.55, 
    268.65, 268.55, 268.25, 267.05, 265.95, 265.95, 266.25, 266.35, 267.15, 
    267.05, 267.35, 266.55, 266.35, 265.35, 266.25, 268.45, 267.75, 268.15, 
    268.25, 268.55, 267.95, 267.45, 268.05, 267.45, 268.55, 268.95, 268.55, 
    268.85, 268.55, 268.95, 268.95, 268.85, 269.15, 269.25, 269.45, 270.05, 
    270.05, 270.05, 270.45, 270.45, 270.55, 270.65, 270.75, 270.75, 270.75, 
    270.75, 270.75, 270.65, 270.45, 270.45, 270.25, 270.55, 270.85, 270.75, 
    270.55, 270.95, 271.45, 271.75, 271.95, 272.05, 271.85, 271.55, 271.75, 
    272.05, 272.35, 272.75, 272.95, 273.15, 273.25, 273.25, 273.25, 273.15, 
    273.05, 273.05, 272.65, 272.85, 273.05, 273.25, 273.15, 272.95, 272.95, 
    272.85, 272.75, 272.15, 272.15, 271.65, 271.65, 271.55, 271.65, 271.45, 
    270.95, 270.65, 270.55, 270.75, 270.75, 270.65, 270.45, 270.55, 270.35, 
    270.25, 270.15, 270.05, 269.95, 270.05, 269.95, 269.95, 269.85, 269.55, 
    269.25, 269.15, 268.95, 268.55, 268.25, 267.85, 267.15, 267.55, 267.25, 
    267.25, 267.15, 267.45, 267.75, 268.05, 268.15, 268.55, 268.35, 268.35, 
    268.95, 269.45, 270.25, 270.15, 270.45, 270.75, 270.55, 270.55, 270.45, 
    270.75, 270.85, 271.05, 271.25, 271.15, 271.35, 271.25, 270.95, 270.85, 
    270.95, 271.15, 270.85, 270.85, 271.05, 270.95, 270.85, 270.75, 270.85, 
    270.75, 270.85, 271.15, 271.55, 271.85, 272.25, 272.35, 272.45, 272.45, 
    272.45, 272.45, 272.45, 272.35, 272.25, 272.35, 272.65, 272.95, 272.95, 
    272.95, 272.95, 272.95, 273.05, 273.05, 273.25, 273.15, 273.15, 273.15, 
    273.05, 272.85, 272.25, 271.75, 272.05, 272.65, 272.25, 271.85, 271.65, 
    272.25, 272.45, 271.75, 271.05, 270.55, 270.95, 271.65, 270.95, 269.75, 
    269.65, 269.15, 268.75, 268.45, 267.95, 267.65, 267.45, 267.25, 266.95, 
    266.75, 266.45, 266.35, 265.85, 265.25, 265.05, 264.25, 264.25, 264.15, 
    263.45, 263.45, 263.15, 262.85, 262.35, 262.05, 261.95, 261.55, 261.35, 
    260.95, 260.75, 260.65, 260.15, 260.25, 260.75, 260.65, 260.55, 260.15, 
    259.75, 259.45, 259.65, 259.05, 259.25, 259.65, 259.65, 259.85, 259.65, 
    259.65, 259.75, 259.95, 259.85, 260.25, 260.35, 260.75, 261.05, 260.95, 
    260.85, 261.55, 261.95, 261.85, 262.05, 262.25, 262.15, 262.45, 262.45, 
    262.75, 263.15, 262.85, 262.95, 263.05, 263.05, 263.15, 263.25, 263.25, 
    263.35, 263.15, 263.45, 263.65, 263.65, 264.05, 263.65, 264.25, 264.25, 
    264.55, 264.25, 266.25, 265.25, 266.75, 265.65, 266.55, 267.05, 265.85, 
    265.65, 264.75, 264.35, 264.25, 264.55, 264.55, 265.55, 264.05, 264.05, 
    264.05, 264.55, 263.65, 264.95, 265.05, 265.85, 265.25, 266.15, 266.75, 
    266.35, 265.85, 266.75, 266.35, 266.45, 266.35, 266.45, 266.75, 266.35, 
    266.75, 267.15, 267.15, 266.95, 266.25, 265.85, 266.05, 265.95, 269.25, 
    269.05, 269.55, 270.15, 270.25, 270.15, 270.45, 270.35, 270.35, 270.65, 
    270.95, 271.05, 271.35, 271.85, 271.95, 271.75, 271.85, 272.05, 272.65, 
    272.85, 272.65, 272.75, 272.95, 273.05, 273.05, 273.05, 272.65, 272.95, 
    273.35, 273.25, 273.15, 273.05, 273.15, 272.95, 272.95, 272.95, 272.95, 
    272.95, 272.85, 272.75, 272.85, 272.95, 272.95, 272.95, 273.15, 273.05, 
    273.05, 272.75, 273.15, 273.35, 273.05, 273.05, 272.65, 272.95, 273.45, 
    273.25, 273.25, 273.75, 273.75, 273.75, 273.65, 273.65, 273.55, 273.45, 
    273.05, 272.85, 272.75, 273.55, 273.95, 272.05, 272.95, 272.75, 272.95, 
    273.25, 273.05, 273.05, 273.05, 273.05, 273.25, 273.55, 273.65, 273.55, 
    273.55, 273.35, 273.25, 273.45, 273.55, 273.45, 273.35, 273.35, 273.85, 
    273.15, 272.75, 272.35, 272.35, 272.05, 271.95, 272.25, 271.15, 270.35, 
    269.85, 269.25, 268.45, 267.85, 267.15, 267.05, 266.75, 266.25, 265.95, 
    265.85, 265.85, 265.75, 265.45, 265.35, 265.25, 265.25, 265.35, 265.35, 
    265.35, 265.15, 265.15, 265.05, 264.95, 264.95, 264.95, 264.95, 264.85, 
    264.85, 264.95, 264.85, 264.75, 264.85, 264.85, 264.95, 264.95, 265.25, 
    264.85, 264.65, 264.15, 264.05, 263.85, 263.85, 263.75, 264.05, 264.25, 
    264.45, 264.25, 264.25, 264.15, 264.25, 263.25, 262.35, 260.65, 260.15, 
    261.35, 261.35, 261.25, 260.95, 260.45, 259.95, 259.25, 258.95, 258.55, 
    258.15, 257.85, 258.55, 258.65, 259.05, 259.85, 260.65, 261.55, 263.65, 
    264.05, 264.25, 264.35, 264.35, 263.95, 263.05, 262.85, 262.65, 262.45, 
    261.95, 261.45, 258.25, 257.75, 257.45, 257.35, 257.15, 257.15, 256.65, 
    256.75, 256.95, 256.95, 256.75, 256.55, 256.35, 256.25, 256.05, 255.85, 
    255.65, 255.35, 254.45, 254.25, 254.05, 253.95, 253.95, 253.85, 253.95, 
    253.85, 253.85, 253.75, 253.85, 253.95, 253.95, 254.05, 254.15, 254.25, 
    254.35, 254.45, 254.95, 254.95, 255.15, 255.15, 255.25, 255.25, 255.25, 
    255.35, 255.35, 255.25, 255.25, 255.05, 254.75, 254.75, 254.75, 254.75, 
    254.65, 254.75, 255.15, 255.15, 255.15, 255.15, 255.15, 255.15, 255.25, 
    255.35, 255.35, 255.35, 255.25, 255.05, 253.25, 253.15, 253.05, 252.95, 
    252.85, 252.65, 252.95, 252.95, 253.05, 252.95, 252.75, 252.55, 252.55, 
    252.65, 252.65, 252.45, 252.25, 252.25, 252.25, 252.15, 252.05, 251.95, 
    251.95, 251.85, 249.45, 249.35, 249.35, 249.25, 249.35, 249.65, 249.85, 
    250.55, 251.55, 252.45, 253.75, 254.95, 256.95, 258.05, 259.15, 260.45, 
    261.45, 262.45, 263.35, 264.25, 265.05, 265.75, 266.35, 266.95, 267.45, 
    267.95, 268.45, 268.85, 269.25, 269.35, 268.85, 269.05, 268.95, 268.75, 
    268.85, 268.95, 269.05, 269.25, 269.55, 269.85, 270.05, 270.35, 270.55, 
    270.85, 271.15, 271.25, 271.35, 271.05, 270.55, 269.75, 269.25, 268.75, 
    268.25, 267.95, 268.45, 268.85, 269.35, 269.65, 270.05, 270.45, 269.05, 
    269.75, 269.95, 269.75, 269.25, 268.75, 268.05, 267.15, 266.55, 266.65, 
    267.45, 268.25, 268.85, 269.75, 271.05, 271.75, 272.05, 271.85, 271.95, 
    271.95, 272.05, 272.15, 272.05, 272.15, 272.05, 271.85, 271.55, 270.85, 
    269.95, 269.05, 268.35, 267.95, 267.35, 266.55, 265.75, 265.45, 265.15, 
    264.95, 264.75, 264.55, 264.15, 264.55, 264.15, 263.95, 263.85, 263.75, 
    263.75, 263.15, 262.95, 262.65, 262.55, 262.35, 262.15, 263.25, 263.15, 
    262.75, 262.25, 261.65, 261.35, 261.05, 261.05, 261.15, 261.15, 260.95, 
    260.85, 263.65, 263.65, 263.25, 262.65, 262.15, 261.85, 260.35, 260.05, 
    259.75, 259.35, 259.15, 259.15, 259.85, 260.05, 260.15, 260.05, 260.25, 
    260.45, 260.65, 260.55, 260.65, 260.55, 260.35, 260.35, 260.45, 260.45, 
    260.55, 260.55, 260.55, 260.65, 259.85, 259.85, 259.85, 259.85, 259.95, 
    259.95, 260.55, 260.75, 261.05, 261.25, 261.45, 261.65, 263.25, 263.55, 
    263.85, 264.15, 264.35, 264.55, 265.45, 265.45, 265.45, 265.55, 265.55, 
    265.55, 264.85, 264.75, 264.65, 264.55, 264.45, 264.35, 263.75, 263.75, 
    263.75, 263.75, 263.65, 263.55, 263.45, 263.35, 263.15, 263.05, 262.75, 
    262.25, 261.65, 261.25, 260.85, 260.55, 260.05, 259.65, 258.55, 257.95, 
    257.55, 257.25, 256.75, 256.45, 256.85, 256.75, 256.55, 256.15, 256.15, 
    256.55, 256.25, 256.75, 256.85, 257.75, 259.05, 259.85, 259.35, 260.15, 
    260.45, 260.35, 260.35, 260.25, 260.25, 260.75, 261.15, 261.45, 261.55, 
    261.75, 260.95, 261.25, 261.75, 262.45, 263.55, 264.55, 265.95, 267.05, 
    267.95, 268.75, 269.25, 269.65, 270.15, 270.35, 270.65, 270.75, 270.85, 
    270.85, 270.35, 269.75, 269.65, 269.95, 270.05, 270.05, 270.55, 270.45, 
    270.35, 269.95, 269.55, 269.35, 268.75, 269.45, 269.95, 270.45, 270.65, 
    270.85, 270.95, 270.85, 270.55, 270.25, 269.75, 269.25, 269.75, 269.35, 
    269.15, 268.95, 268.85, 268.75, 268.35, 268.35, 268.45, 268.65, 268.85, 
    269.25, 268.95, 269.15, 269.35, 269.35, 269.25, 269.15, 268.75, 268.15, 
    267.35, 266.55, 265.65, 264.85, 264.95, 264.45, 264.05, 263.75, 263.35, 
    263.15, 263.75, 263.65, 263.55, 263.25, 262.95, 262.75, 262.75, 262.35, 
    261.85, 261.45, 260.95, 260.45, 258.75, 258.25, 257.85, 257.45, 257.35, 
    257.25, 256.35, 256.35, 256.35, 256.45, 256.45, 256.45, 256.65, 256.65, 
    256.65, 256.75, 256.75, 256.85, 257.15, 257.15, 257.15, 257.25, 257.15, 
    256.95, 256.35, 255.85, 255.45, 254.95, 254.55, 254.25, 253.85, 253.45, 
    253.05, 252.75, 252.45, 252.35, 253.15, 252.95, 252.75, 252.65, 252.65, 
    252.75, 253.35, 253.25, 253.35, 253.45, 253.55, 253.75, 253.65, 253.95, 
    254.15, 254.45, 254.75, 255.05, 255.35, 255.65, 255.95, 256.25, 256.55, 
    256.95, 257.25, 257.75, 258.25, 258.75, 259.35, 259.95, 269.25, 269.15, 
    269.05, 268.95, 268.75, 268.85, 268.95, 268.95, 268.85, 268.85, 268.85, 
    268.15, 268.25, 268.25, 268.05, 267.85, 267.55, 266.75, 266.55, 266.35, 
    266.15, 266.05, 265.35, 265.75, 265.95, 265.55, 264.75, 263.85, 263.05, 
    265.15, 264.65, 263.85, 263.25, 262.75, 262.45, 262.75, 262.35, 262.05, 
    261.95, 261.85, 261.75, 260.85, 260.55, 260.45, 260.55, 260.45, 260.45, 
    260.45, 260.55, 260.75, 260.75, 260.85, 260.85, 260.55, 260.75, 260.75, 
    260.65, 260.45, 260.35, 260.15, 260.15, 260.15, 259.95, 259.95, 259.85, 
    259.35, 259.05, 258.85, 258.75, 258.55, 256.25, 255.75, 255.85, 256.05, 
    256.05, 256.05, 255.05, 255.15, 255.25, 255.35, 255.45, 255.25, 253.55, 
    253.85, 254.05, 254.25, 254.25, 254.45, 253.95, 254.05, 254.35, 254.55, 
    254.95, 255.15, 253.95, 254.35, 254.85, 255.35, 255.75, 256.35, 256.15, 
    256.35, 256.95, 257.65, 258.35, 258.85, 258.15, 258.05, 258.15, 258.25, 
    258.35, 258.25, 261.05, 260.95, 261.25, 261.25, 261.45, 261.45, 260.55, 
    260.35, 260.15, 260.35, 260.35, 260.35, 260.55, 260.35, 260.05, 259.55, 
    259.05, 258.55, 257.15, 256.65, 255.95, 255.45, 255.15, 255.05, 251.95, 
    251.25, 250.65, 250.25, 249.85, 249.45, 249.35, 249.15, 248.85, 248.75, 
    248.95, 249.45, 265.85, 266.05, 266.45, 267.05, 254.15, 253.95, 253.75, 
    254.05, 254.15, 254.35, 254.75, 254.65, 254.65, 254.85, 254.75, 254.95, 
    255.65, 255.95, 256.15, 256.45, 256.65, 256.95, 255.35, 255.25, 255.25, 
    255.15, 255.15, 255.15, 255.65, 255.85, 256.05, 256.15, 256.35, 256.65, 
    256.25, 256.45, 256.45, 256.75, 256.95, 257.25, 258.85, 258.95, 259.05, 
    259.05, 258.95, 258.85, 258.85, 258.85, 258.85, 258.95, 258.85, 259.05, 
    259.45, 259.15, 259.35, 259.85, 260.25, 260.45, 260.75, 261.15, 261.15, 
    261.45, 262.15, 262.75, 263.95, 264.15, 264.35, 264.25, 264.55, 264.45, 
    263.65, 263.35, 263.35, 263.85, 264.35, 265.15, 266.15, 266.75, 267.25, 
    267.95, 268.55, 269.05, 269.85, 269.95, 270.05, 269.95, 269.95, 269.85, 
    269.65, 269.75, 269.85, 270.15, 270.55, 270.95, 270.95, 271.25, 271.35, 
    271.45, 271.55, 271.65, 271.85, 271.95, 271.95, 271.95, 271.95, 271.95, 
    272.05, 272.05, 271.95, 271.95, 271.85, 271.85, 271.75, 271.65, 271.55, 
    271.45, 271.25, 270.95, 270.35, 269.25, 268.25, 267.25, 266.35, 265.75, 
    264.15, 263.45, 262.65, 262.15, 262.45, 263.05, 263.05, 263.25, 264.05, 
    264.65, 265.35, 265.75, 265.35, 265.65, 265.55, 266.05, 266.35, 266.55, 
    266.55, 266.75, 266.95, 267.15, 267.25, 267.45, 267.85, 268.15, 267.95, 
    267.95, 268.15, 268.35, 269.15, 269.35, 269.35, 269.25, 268.75, 267.85, 
    269.95, 268.95, 267.85, 266.85, 265.95, 265.05, 266.35, 265.75, 265.15, 
    264.35, 263.55, 262.75, 263.25, 262.45, 261.65, 260.95, 260.25, 259.65, 
    257.95, 257.35, 256.85, 256.35, 255.85, 255.55, 255.05, 255.05, 255.15, 
    255.45, 255.75, 255.85, 253.95, 253.85, 253.65, 253.55, 253.45, 253.25, 
    252.65, 252.55, 252.55, 252.55, 252.65, 252.75, 252.75, 252.85, 252.95, 
    252.95, 253.05, 253.15, 253.15, 253.15, 253.15, 253.25, 253.45, 253.65, 
    252.85, 253.15, 253.25, 253.25, 253.15, 253.05, 252.65, 252.65, 252.85, 
    252.95, 253.05, 253.25, 252.45, 252.65, 252.95, 253.35, 253.75, 254.05, 
    253.25, 253.45, 253.75, 254.05, 254.15, 254.35, 253.35, 253.75, 254.05, 
    254.05, 254.05, 253.95, 253.35, 253.65, 253.55, 253.55, 252.95, 252.75, 
    252.15, 252.15, 254.65, 255.65, 255.45, 255.35, 255.95, 255.85, 255.85, 
    255.75, 255.85, 256.05, 256.35, 257.75, 258.55, 258.65, 258.85, 259.15, 
    260.35, 260.65, 260.95, 261.35, 261.75, 262.05, 262.45, 262.65, 262.85, 
    262.85, 263.15, 263.05, 262.15, 262.55, 262.95, 263.35, 263.45, 262.95, 
    261.35, 260.95, 260.35, 260.65, 261.25, 262.25, 264.05, 264.55, 265.05, 
    265.75, 266.45, 267.45, 268.85, 269.25, 269.85, 270.15, 270.45, 270.65, 
    270.45, 270.55, 270.85, 270.95, 270.65, 270.65, 270.65, 270.55, 270.45, 
    270.55, 270.55, 270.65, 270.85, 271.15, 271.05, 271.15, 271.25, 270.95, 
    270.55, 270.35, 270.25, 270.45, 270.65, 270.35, 270.15, 270.05, 269.95, 
    269.95, 270.15, 270.85, 270.95, 271.05, 271.25, 271.55, 271.65, 271.25, 
    271.25, 271.15, 270.85, 270.75, 270.35, 270.05, 269.85, 269.35, 268.85, 
    268.45, 268.35, 268.25, 268.15, 267.95, 267.45, 267.05, 266.75, 266.25, 
    266.15, 266.05, 265.75, 265.45, 265.15, 265.75, 265.25, 264.85, 264.25, 
    263.95, 263.55, 263.05, 262.75, 262.55, 262.45, 262.25, 261.95, 261.35, 
    261.35, 262.15, 262.55, 262.25, 262.55, 261.25, 261.25, 261.25, 260.85, 
    260.55, 261.55, 261.95, 261.65, 262.45, 262.85, 262.95, 262.75, 262.35, 
    262.35, 262.75, 263.25, 263.45, 263.55, 263.65, 263.75, 263.85, 263.95, 
    264.05, 264.15, 263.25, 263.35, 263.45, 263.55, 263.65, 263.75, 260.15, 
    260.35, 260.85, 261.25, 261.65, 262.05, 260.25, 260.65, 260.95, 261.45, 
    261.85, 262.25, 261.05, 260.75, 260.75, 260.75, 260.55, 260.45, 259.75, 
    259.75, 260.15, 260.45, 260.65, 260.95, 259.55, 259.55, 259.55, 259.55, 
    259.55, 259.75, 258.45, 258.55, 258.75, 258.75, 258.75, 258.45, 255.25, 
    255.55, 255.65, 255.55, 255.45, 255.55, 251.15, 251.15, 251.15, 251.35, 
    251.45, 251.55, 248.85, 249.65, 250.25, 250.85, 251.35, 251.55, 247.25, 
    247.85, 248.45, 248.85, 249.35, 249.35, 250.15, 250.75, 251.35, 251.85, 
    252.15, 252.35, 248.95, 248.85, 248.95, 249.15, 249.05, 249.05, 249.25, 
    249.65, 250.35, 250.95, 251.65, 252.35, 258.95, 259.35, 259.75, 260.35, 
    260.75, 261.15, 261.75, 262.25, 255.65, 255.35, 255.75, 256.45, 256.95, 
    256.75, 255.15, 254.95, 254.85, 255.15, 255.85, 256.75, 256.35, 256.85, 
    257.45, 257.95, 258.55, 259.05, 260.85, 261.85, 262.65, 263.25, 263.65, 
    263.65, 262.25, 261.75, 261.65, 261.75, 262.55, 263.25, 263.55, 264.95, 
    266.65, 268.25, 269.15, 269.75, 270.15, 270.45, 270.75, 271.15, 271.55, 
    271.75, 271.95, 271.95, 271.95, 272.05, 272.05, 272.05, 271.75, 271.75, 
    271.85, 271.85, 271.95, 271.95, 271.85, 271.85, 271.85, 271.85, 271.85, 
    271.55, 270.75, 270.15, 269.95, 270.15, 270.45, 269.85, 269.85, 268.85, 
    267.85, 266.85, 266.05, 266.05, 264.45, 264.55, 264.75, 265.05, 265.35, 
    265.55, 265.25, 264.65, 264.65, 264.85, 264.95, 263.85, 258.55, 258.85, 
    259.85, 260.45, 261.15, 262.75, 263.25, 264.65, 266.05, 267.45, 268.15, 
    269.15, 268.95, 269.55, 269.95, 270.35, 270.55, 270.55, 269.45, 269.65, 
    269.75, 269.65, 268.85, 268.65, 268.35, 268.25, 267.55, 266.55, 265.25, 
    264.35, 266.45, 266.85, 267.15, 267.25, 267.65, 267.75, 267.55, 267.85, 
    268.05, 268.25, 268.25, 268.35, 268.75, 268.95, 268.85, 268.75, 268.45, 
    267.85, 269.45, 269.35, 268.65, 268.35, 268.55, 268.75, 266.95, 266.85, 
    266.85, 266.25, 265.75, 265.75, 268.45, 268.45, 268.55, 268.65, 268.75, 
    268.75, 269.45, 269.45, 268.95, 268.85, 268.75, 268.45, 269.75, 269.65, 
    269.35, 269.05, 268.85, 268.65, 268.25, 268.45, 268.65, 268.75, 268.65, 
    268.35, 264.95, 264.45, 263.95, 263.35, 262.85, 262.45, 267.15, 266.85, 
    266.55, 266.05, 265.75, 265.55, 265.65, 265.45, 265.25, 264.45, 263.45, 
    262.65, 260.45, 259.65, 258.85, 258.15, 257.55, 257.15, 260.55, 260.25, 
    260.05, 259.85, 259.55, 259.25, 261.75, 262.45, 262.85, 262.45, 261.85, 
    262.05, 260.25, 259.95, 260.55, 261.25, 261.75, 262.35, 262.95, 263.45, 
    264.25, 264.95, 264.95, 264.65, 263.45, 263.05, 262.65, 262.25, 261.75, 
    261.15, 260.45, 260.15, 259.65, 259.15, 258.85, 258.25, 258.75, 258.55, 
    258.35, 257.95, 257.55, 257.15, 257.75, 257.55, 257.25, 256.95, 256.85, 
    256.55, 253.95, 253.95, 254.55, 255.25, 255.85, 256.15, 256.55, 256.65, 
    256.55, 256.55, 256.75, 256.95, 255.15, 255.75, 256.05, 256.55, 257.05, 
    257.45, 258.15, 258.55, 259.05, 259.45, 259.85, 260.15, 261.15, 261.25, 
    261.25, 261.05, 260.85, 260.75, 260.55, 260.35, 260.25, 260.25, 260.35, 
    260.35, 260.95, 260.95, 260.95, 260.85, 260.85, 260.85, 261.55, 261.45, 
    261.25, 261.05, 260.95, 261.15, 259.35, 259.25, 259.15, 258.65, 257.95, 
    257.35, 254.75, 254.05, 253.75, 254.35, 255.05, 255.75, 254.95, 255.35, 
    255.75, 256.25, 256.25, 256.05, 257.85, 257.45, 257.75, 258.85, 259.55, 
    260.15, 259.25, 259.35, 259.65, 260.65, 262.05, 263.75, 262.25, 263.65, 
    265.45, 267.55, 269.65, 270.95, 271.45, 271.55, 271.65, 271.75, 271.85, 
    271.85, 271.95, 271.95, 271.75, 271.45, 271.65, 271.65, 271.25, 271.35, 
    271.55, 271.45, 271.55, 271.45, 271.65, 271.65, 271.75, 271.65, 271.35, 
    270.75, 270.35, 270.35, 270.85, 271.35, 271.85, 272.25, 272.25, 271.65, 
    269.45, 268.15, 267.15, 266.25, 265.35, 264.85, 264.45, 263.95, 263.95, 
    263.85, 265.25, 264.85, 264.25, 263.85, 263.65, 263.75, 263.85, 264.55, 
    265.15, 265.75, 266.15, 266.75, 265.85, 266.65, 267.55, 268.35, 268.55, 
    268.65, 269.35, 269.85, 270.45, 271.05, 271.45, 271.85, 272.25, 272.25, 
    272.35, 272.55, 272.65, 272.75, 272.95, 272.95, 273.05, 273.05, 273.05, 
    273.25, 273.45, 273.45, 273.45, 273.45, 273.45, 273.55, 273.55, 273.45, 
    273.25, 273.15, 272.85, 272.55, 272.35, 272.25, 272.15, 271.95, 271.85, 
    271.95, 271.75, 271.65, 271.55, 271.55, 271.85, 271.85, 271.65, 271.35, 
    271.25, 271.35, 271.75, 271.95, 272.05, 272.15, 272.15, 272.15, 272.25, 
    272.35, 272.65, 272.65, 272.55, 272.15, 271.75, 271.25, 270.35, 269.85, 
    269.25, 269.05, 269.45, 270.05, 270.15, 271.45, 272.35, 272.75, 273.05, 
    273.15, 273.15, 273.15, 273.25, 272.95, 270.35, 268.35, 268.15, 266.95, 
    266.25, 265.55, 264.75, 264.05, 262.25, 261.95, 261.85, 261.75, 261.65, 
    261.75, 260.95, 260.95, 260.85, 260.85, 260.85, 260.85, 260.75, 260.65, 
    260.85, 260.85, 260.95, 261.45, 262.35, 263.65, 265.25, 267.25, 269.75, 
    271.65, 272.45, 272.55, 272.55, 272.45, 272.35, 271.75, 271.25, 271.15, 
    270.95, 270.75, 270.75, 271.25, 270.65, 270.45, 270.25, 270.25, 267.95, 
    267.55, 266.65, 265.95, 265.45, 265.15, 264.85, 265.15, 264.95, 264.85, 
    264.95, 264.85, 264.85, 265.45, 265.75, 265.65, 265.75, 265.95, 266.25, 
    265.75, 266.75, 267.75, 268.85, 270.25, 271.35, 272.15, 272.35, 272.25, 
    271.95, 271.55, 271.15, 271.05, 270.65, 270.35, 269.95, 269.55, 269.05, 
    269.35, 268.95, 268.55, 268.35, 268.35, 268.15, 266.85, 267.35, 267.75, 
    268.05, 268.15, 268.55, 267.45, 267.95, 268.85, 269.75, 270.45, 271.15, 
    271.35, 271.05, 270.85, 270.65, 270.45, 270.15, 269.25, 269.05, 268.85, 
    268.45, 268.05, 267.85, 267.85, 268.05, 267.95, 267.95, 267.95, 267.95, 
    267.15, 266.95, 266.95, 266.75, 266.95, 267.15, 267.45, 267.45, 267.55, 
    267.65, 267.85, 267.75, 267.85, 268.15, 268.15, 268.45, 268.75, 269.05, 
    268.95, 268.85, 268.85, 269.15, 269.45, 269.75, 269.75, 269.85, 269.95, 
    270.15, 270.35, 270.65, 270.85, 271.35, 271.65, 271.45, 271.35, 271.65, 
    271.05, 271.25, 271.45, 271.75, 271.95, 272.05, 272.25, 272.45, 272.75, 
    272.95, 273.05, 273.05, 273.15, 273.15, 273.25, 273.25, 273.15, 273.05, 
    272.95, 272.85, 272.25, 271.05, 270.05, 269.05, 269.15, 268.55, 268.25, 
    268.15, 267.95, 266.55, 266.25, 266.05, 265.85, 265.55, 265.15, 265.25, 
    264.95, 264.75, 264.55, 264.25, 264.05, 263.75, 263.55, 263.45, 263.35, 
    263.15, 263.15, 263.15, 263.15, 263.05, 262.95, 262.95, 263.05, 263.05, 
    263.15, 263.35, 263.45, 263.55, 263.75, 263.75, 263.75, 263.85, 263.85, 
    263.85, 263.95, 263.35, 263.35, 263.35, 263.25, 263.25, 263.25, 263.45, 
    263.45, 263.45, 263.35, 263.35, 263.35, 263.65, 263.65, 263.55, 263.55, 
    263.35, 263.35, 263.75, 263.75, 263.75, 263.75, 263.75, 263.75, 263.95, 
    263.95, 263.95, 263.95, 263.95, 263.75, 264.05, 263.95, 263.75, 263.75, 
    263.65, 263.45, 263.55, 263.45, 263.45, 263.45, 263.35, 263.35, 262.95, 
    262.35, 261.85, 261.45, 261.15, 260.95, 261.65, 261.85, 261.95, 262.05, 
    262.15, 262.05, 262.35, 262.25, 262.15, 261.95, 261.75, 261.65, 261.65, 
    261.65, 261.65, 261.45, 261.35, 261.15, 261.55, 261.25, 261.05, 260.85, 
    260.85, 260.85, 260.95, 260.85, 260.75, 260.65, 260.75, 261.05, 260.55, 
    260.75, 260.95, 261.05, 261.35, 261.75, 260.25, 260.25, 260.05, 260.15, 
    260.45, 260.65, 260.95, 260.95, 261.15, 261.45, 261.85, 262.25, 263.45, 
    263.85, 264.35, 265.05, 265.85, 266.15, 265.95, 266.25, 266.65, 266.65, 
    266.75, 266.45, 266.25, 265.75, 265.45, 265.45, 265.35, 265.15, 264.95, 
    265.55, 266.05, 264.85, 263.65, 263.05, 262.55, 262.25, 262.05, 262.05, 
    262.05, 262.05, 262.45, 262.45, 262.35, 262.05, 261.75, 261.55, 260.95, 
    261.15, 261.25, 261.35, 260.95, 260.55, 259.35, 259.65, 259.75, 259.65, 
    259.25, 258.75, 258.35, 258.35, 258.45, 258.35, 258.45, 258.55, 258.65, 
    258.95, 259.25, 260.05, 261.15, 262.25, 259.95, 260.65, 261.55, 262.45, 
    263.25, 263.85, 265.05, 265.05, 265.05, 265.25, 265.45, 265.65, 264.65, 
    264.45, 264.65, 264.75, 264.75, 264.85, 264.45, 264.65, 265.05, 265.65, 
    266.15, 266.35, 265.55, 265.85, 266.25, 266.55, 267.05, 267.35, 266.85, 
    267.35, 267.75, 268.15, 268.45, 268.85, 268.55, 268.75, 268.95, 269.05, 
    269.05, 269.05, 268.05, 267.95, 267.85, 267.95, 267.95, 267.75, 267.45, 
    267.55, 267.75, 267.95, 268.05, 268.35, 268.25, 268.65, 269.05, 269.15, 
    268.95, 269.15, 267.85, 267.95, 268.05, 268.25, 268.45, 268.55, 267.75, 
    268.15, 267.95, 268.05, 268.25, 268.45, 268.45, 268.65, 268.85, 268.95, 
    269.05, 269.15, 269.25, 269.35, 269.45, 269.55, 269.65, 269.65, 269.95, 
    269.85, 269.55, 268.95, 268.45, 267.85, 267.55, 267.85, 268.25, 268.65, 
    269.15, 269.55, 268.65, 268.85, 268.95, 269.15, 269.35, 269.45, 268.85, 
    268.65, 268.65, 268.15, 267.55, 267.25, 266.05, 266.15, 266.15, 265.45, 
    265.25, 265.75, 265.55, 265.95, 266.45, 266.65, 266.85, 267.25, 267.05, 
    267.35, 267.55, 267.65, 267.65, 268.15, 268.25, 268.55, 268.75, 268.55, 
    268.35, 267.75, 267.35, 267.25, 267.25, 267.25, 267.25, 267.35, 265.15, 
    265.25, 265.25, 264.95, 264.55, 264.35, 264.45, 265.15, 265.65, 266.15, 
    266.65, 266.85, 267.25, 267.35, 267.45, 267.85, 268.35, 268.65, 267.35, 
    267.25, 266.55, 265.95, 265.55, 265.75, 266.45, 266.35, 266.45, 266.55, 
    266.75, 266.95, 267.95, 267.95, 268.05, 268.15, 268.25, 268.05, 265.55, 
    265.95, 266.35, 266.75, 267.15, 267.35, 267.65, 267.75, 267.55, 267.65, 
    267.95, 268.15, 268.15, 268.35, 268.55, 268.75, 268.95, 269.05, 268.45, 
    268.65, 268.85, 269.05, 269.25, 269.45, 268.95, 268.65, 268.35, 267.95, 
    267.55, 267.15, 267.05, 266.95, 266.75, 266.45, 266.25, 266.25, 265.85, 
    265.85, 265.75, 265.65, 265.55, 265.45, 264.65, 264.65, 264.55, 264.45, 
    264.45, 264.35, 265.25, 265.35, 265.45, 265.65, 265.85, 266.05, 264.95, 
    264.85, 264.55, 264.05, 263.35, 262.75, 265.75, 265.35, 265.45, 265.65, 
    265.65, 265.55, 265.05, 265.15, 265.25, 265.45, 265.45, 265.25, 264.45, 
    264.75, 264.65, 264.55, 264.05, 263.55, 264.15, 263.75, 263.65, 263.75, 
    263.95, 263.95, 263.15, 264.15, 264.85, 265.05, 264.95, 265.25, 266.35, 
    266.25, 265.95, 265.65, 265.05, 264.55, 264.15, 263.75, 263.45, 263.15, 
    262.65, 262.25, 262.35, 262.05, 261.65, 261.25, 260.95, 260.85, 260.15, 
    259.95, 259.95, 260.15, 260.45, 260.75, 261.35, 261.75, 262.25, 262.75, 
    263.15, 263.85, 265.15, 265.85, 266.75, 267.25, 267.35, 267.25, 267.55, 
    267.15, 266.75, 266.85, 266.95, 267.05, 266.95, 266.15, 265.55, 264.85, 
    264.35, 264.05, 264.35, 264.05, 263.75, 263.45, 263.25, 263.15, 263.25, 
    263.15, 263.05, 263.05, 262.95, 262.95, 261.55, 261.45, 261.35, 261.25, 
    261.25, 261.25, 261.45, 261.45, 261.55, 261.65, 261.75, 261.85, 262.05, 
    262.15, 262.15, 262.25, 262.35, 262.55, 262.85, 263.25, 263.35, 263.55, 
    265.45, 265.75, 264.85, 264.95, 264.85, 264.75, 264.65, 264.25, 264.55, 
    264.25, 263.65, 263.15, 262.95, 262.65, 261.85, 261.65, 262.65, 263.45, 
    264.35, 265.35, 265.35, 266.45, 267.45, 268.45, 269.25, 269.65, 269.95, 
    272.15, 269.55, 269.55, 269.95, 270.35, 271.65, 271.65, 271.65, 271.35, 
    271.25, 271.05, 270.85, 270.65, 270.75, 270.85, 271.25, 271.35, 271.15, 
    270.85, 270.75, 270.95, 270.75, 270.75, 270.75, 271.65, 271.75, 271.85, 
    272.05, 272.35, 272.25, 272.25, 271.85, 271.75, 271.85, 271.35, 271.35, 
    271.45, 271.25, 271.55, 271.95, 271.85, 271.65, 271.35, 271.65, 271.65, 
    271.65, 271.65, 271.25, 270.55, 270.65, 270.45, 270.55, 269.75, 269.45, 
    270.65, 270.85, 271.15, 269.95, 269.25, 269.45, 269.55, 268.25, 268.85, 
    268.75, 267.55, 268.35, 266.45, 270.85, 271.25, 269.15, 269.35, 268.75, 
    269.85, 270.15, 271.35, 271.15, 271.45, 272.25, 271.85, 272.65, 272.05, 
    272.45, 272.45, 271.65, 271.45, 270.85, 271.45, 271.55, 271.55, 271.25, 
    271.45, 271.35, 271.45, 271.45, 271.65, 271.75, 271.65, 271.75, 271.55, 
    271.05, 270.95, 271.15, 271.25, 271.35, 271.25, 271.15, 270.95, 270.75, 
    270.65, 270.65, 270.45, 270.35, 270.05, 269.95, 269.75, 269.75, 269.55, 
    269.45, 269.45, 269.15, 269.35, 269.25, 268.85, 269.05, 269.15, 269.15, 
    268.95, 268.75, 268.35, 268.15, 268.15, 268.25, 267.85, 267.65, 267.45, 
    267.55, 266.75, 266.75, 266.85, 267.15, 267.05, 267.15, 267.15, 266.95, 
    267.15, 267.15, 267.05, 267.05, 267.15, 267.25, 267.25, 267.55, 268.15, 
    268.85, 269.55, 270.15, 270.35, 270.95, 271.15, 271.95, 272.05, 271.95, 
    272.45, 271.95, 271.85, 271.85, 272.05, 271.65, 271.15, 271.05, 270.75, 
    270.95, 270.95, 270.95, 271.15, 271.15, 270.95, 270.95, 270.75, 270.55, 
    270.35, 270.15, 269.95, 269.85, 269.75, 269.65, 269.45, 269.45, 269.55, 
    269.55, 269.25, 268.95, 268.55, 267.75, 267.65, 267.85, 268.25, 268.25, 
    268.15, 268.35, 268.65, 268.75, 268.95, 268.95, 268.85, 269.25, 268.15, 
    268.35, 268.75, 269.45, 268.55, 267.65, 266.85, 266.35, 265.85, 265.55, 
    265.25, 265.05, 264.95, 264.65, 264.55, 264.65, 264.55, 264.45, 264.35, 
    264.55, 264.45, 264.35, 264.35, 264.35, 264.15, 264.05, 263.85, 263.75, 
    263.45, 263.45, 263.05, 263.05, 263.05, 262.85, 262.75, 262.65, 262.55, 
    262.55, 262.25, 261.95, 261.95, 262.05, 261.95, 262.05, 261.65, 261.45, 
    261.05, 260.75, 260.55, 260.05, 260.45, 261.15, 261.15, 261.45, 260.35, 
    261.35, 261.55, 261.85, 261.65, 260.45, 260.05, 261.45, 262.15, 262.75, 
    263.35, 263.35, 263.35, 263.85, 264.35, 264.85, 265.15, 265.55, 265.45, 
    265.95, 265.95, 266.55, 267.55, 268.35, 268.75, 268.75, 269.05, 269.35, 
    269.55, 269.85, 269.95, 269.65, 269.65, 269.45, 269.55, 269.55, 269.45, 
    269.35, 269.15, 269.05, 268.85, 268.95, 268.85, 268.35, 268.35, 268.25, 
    268.05, 267.85, 267.75, 267.85, 267.85, 267.75, 267.95, 267.65, 267.15, 
    266.95, 267.35, 267.25, 267.15, 267.05, 267.05, 267.15, 266.45, 266.55, 
    266.35, 265.65, 265.85, 265.05, 265.05, 265.15, 265.05, 265.05, 264.65, 
    264.65, 264.45, 264.35, 264.35, 264.05, 263.85, 264.05, 263.65, 263.75, 
    263.75, 263.85, 263.35, 263.25, 263.25, 262.95, 262.45, 261.85, 261.75, 
    260.95, 260.05, 258.95, 258.25, 258.05, 257.95, 257.85, 257.75, 257.85, 
    258.05, 257.85, 257.75, 257.65, 257.65, 257.25, 257.45, 257.55, 257.05, 
    257.05, 257.15, 257.05, 257.45, 257.65, 257.65, 257.75, 257.65, 257.75, 
    258.15, 258.05, 258.55, 258.65, 258.65, 258.75, 259.05, 258.95, 258.95, 
    259.05, 258.95, 258.95, 259.05, 258.95, 258.95, 258.75, 259.65, 259.25, 
    259.25, 259.45, 259.45, 259.85, 259.95, 259.85, 260.05, 261.35, 261.05, 
    260.95, 260.95, 260.55, 261.05, 260.75, 261.15, 260.95, 260.85, 259.95, 
    259.95, 259.55, 259.65, 259.85, 259.55, 259.15, 259.15, 259.15, 258.75, 
    258.55, 258.25, 258.05, 257.45, 257.55, 258.05, 257.95, 258.35, 257.95, 
    257.75, 257.45, 257.65, 257.55, 257.65, 256.95, 257.65, 257.05, 256.75, 
    257.95, 256.85, 257.85, 257.75, 258.15, 257.95, 257.65, 257.85, 257.95, 
    257.25, 257.15, 257.15, 257.75, 257.95, 257.05, 256.65, 257.35, 256.85, 
    256.05, 256.95, 256.15, 256.15, 256.45, 256.55, 256.55, 258.85, 256.95, 
    256.05, 256.75, 256.55, 256.05, 256.35, 256.65, 256.75, 256.35, 257.55, 
    256.25, 254.95, 254.95, 254.95, 254.35, 254.25, 254.25, 255.15, 254.95, 
    255.15, 255.55, 256.15, 255.95, 256.35, 256.35, 256.25, 256.15, 256.05, 
    256.25, 256.15, 255.65, 255.95, 256.25, 257.65, 258.75, 257.95, 257.85, 
    258.05, 257.55, 257.45, 257.25, 256.65, 256.55, 256.55, 256.25, 256.25, 
    255.75, 256.25, 256.85, 256.35, 256.75, 256.65, 257.25, 257.65, 256.25, 
    257.65, 257.35, 258.75, 258.45, 258.05, 258.05, 258.35, 259.25, 259.35, 
    259.45, 259.35, 259.75, 259.55, 259.55, 259.25, 259.25, 259.55, 259.75, 
    259.65, 259.45, 259.45, 259.75, 260.15, 260.45, 260.45, 260.95, 261.05, 
    261.45, 261.15, 261.05, 260.95, 260.05, 260.35, 260.35, 260.15, 259.65, 
    259.65, 259.45, 259.25, 258.55, 259.05, 258.25, 258.35, 258.65, 257.95, 
    257.65, 257.05, 256.95, 257.65, 258.35, 258.05, 258.85, 258.45, 258.15, 
    258.25, 258.45, 258.35, 258.35, 258.25, 258.05, 258.15, 258.35, 258.75, 
    258.85, 259.05, 260.05, 259.85, 261.05, 260.05, 261.05, 262.25, 260.95, 
    261.55, 261.55, 261.45, 260.55, 260.65, 261.05, 260.75, 261.05, 260.85, 
    260.65, 260.75, 261.15, 261.25, 260.15, 260.25, 260.85, 260.65, 260.75, 
    259.45, 259.35, 259.45, 259.25, 259.15, 259.05, 259.05, 259.25, 259.65, 
    259.95, 262.15, 262.45, 262.45, 262.25, 261.85, 262.05, 261.95, 262.15, 
    261.95, 261.15, 260.75, 260.25, 260.25, 259.75, 259.55, 259.05, 258.75, 
    258.95, 258.65, 258.65, 258.55, 258.55, 258.65, 258.55, 258.35, 258.25, 
    258.35, 258.15, 258.15, 258.55, 258.65, 258.55, 258.85, 258.85, 258.95, 
    259.05, 259.75, 259.95, 260.45, 260.85, 261.95, 262.75, 263.45, 262.95, 
    261.65, 262.55, 263.65, 263.75, 263.85, 263.55, 264.05, 265.15, 266.45, 
    265.85, 265.15, 264.85, 264.35, 264.45, 264.65, 264.75, 264.25, 264.45, 
    264.05, 263.55, 263.25, 263.75, 264.35, 264.65, 264.65, 264.15, 263.65, 
    263.25, 263.25, 263.05, 262.75, 262.85, 262.75, 262.35, 262.25, 262.45, 
    261.75, 261.55, 261.65, 261.55, 261.75, 261.45, 260.25, 260.35, 261.25, 
    261.95, 260.35, 261.05, 262.15, 262.15, 260.25, 259.75, 259.25, 257.95, 
    258.45, 258.45, 258.55, 258.65, 258.95, 259.45, 259.95, 260.05, 259.85, 
    260.75, 260.25, 259.95, 260.05, 260.25, 260.55, 261.05, 260.75, 260.85, 
    261.05, 261.25, 261.35, 261.45, 261.25, 260.25, 259.25, 258.95, 258.75, 
    258.75, 258.45, 258.45, 258.55, 258.75, 259.05, 259.45, 259.75, 260.05, 
    260.75, 261.15, 261.45, 262.05, 262.55, 262.85, 263.25, 263.55, 263.85, 
    264.35, 264.45, 264.55, 264.55, 264.85, 264.95, 265.25, 265.35, 265.75, 
    266.05, 266.05, 265.95, 265.15, 265.25, 265.45, 266.55, 266.55, 267.35, 
    267.45, 267.55, 267.55, 267.95, 268.25, 268.05, 266.95, 267.15, 265.65, 
    266.45, 266.35, 265.55, 265.55, 265.65, 266.35, 266.45, 266.45, 266.25, 
    265.25, 265.75, 266.35, 266.35, 265.95, 265.75, 266.15, 266.15, 267.25, 
    266.65, 265.65, 264.75, 264.95, 267.15, 266.55, 266.25, 266.45, 265.05, 
    263.55, 262.95, 260.95, 260.85, 260.55, 260.25, 261.35, 263.35, 262.05, 
    261.75, 262.45, 262.55, 262.35, 262.95, 261.45, 261.85, 263.05, 262.55, 
    262.95, 262.75, 263.15, 264.05, 263.45, 262.85, 262.85, 261.95, 260.65, 
    260.15, 260.55, 259.65, 261.85, 263.35, 264.25, 264.15, 264.35, 264.75, 
    265.25, 265.05, 265.05, 264.55, 264.35, 263.75, 263.25, 263.25, 263.35, 
    263.25, 263.25, 263.45, 263.45, 262.65, 263.05, 262.25, 261.25, 261.05, 
    263.55, 263.65, 263.85, 263.65, 263.85, 264.45, 264.35, 264.25, 264.05, 
    264.35, 264.15, 264.15, 264.15, 263.95, 263.85, 263.85, 263.45, 262.95, 
    262.45, 261.85, 262.05, 261.35, 261.35, 261.45, 260.45, 260.05, 259.65, 
    258.95, 258.55, 258.35, 258.55, 259.05, 259.05, 259.95, 260.95, 261.35, 
    261.95, 261.05, 260.65, 260.45, 260.15, 260.55, 259.95, 259.75, 260.95, 
    260.65, 260.65, 260.05, 258.35, 259.35, 260.05, 259.85, 260.35, 260.35, 
    261.05, 261.25, 262.35, 261.85, 261.15, 260.65, 259.85, 260.05, 259.05, 
    258.65, 259.05, 258.65, 258.45, 257.55, 257.75, 258.35, 258.45, 259.35, 
    259.05, 259.45, 259.35, 259.95, 260.75, 260.85, 260.75, 260.75, 260.95, 
    261.25, 261.45, 262.05, 262.55, 262.35, 262.25, 262.15, 262.15, 261.75, 
    261.95, 261.45, 261.15, 261.35, 260.85, 260.65, 260.45, 259.75, 259.35, 
    259.55, 260.05, 259.75, 259.35, 258.95, 259.05, 258.75, 258.75, 259.05, 
    259.15, 258.95, 259.15, 259.25, 258.65, 258.65, 258.45, 258.45, 258.95, 
    258.45, 258.65, 258.15, 258.15, 258.05, 258.05, 257.85, 258.15, 258.05, 
    258.25, 258.25, 257.85, 257.55, 257.15, 257.35, 257.35, 258.05, 258.05, 
    257.95, 258.15, 258.35, 258.95, 259.55, 259.85, 259.65, 259.35, 259.75, 
    259.95, 259.75, 259.55, 259.25, 259.25, 259.25, 259.05, 258.85, 258.85, 
    259.05, 259.35, 259.75, 260.35, 259.75, 259.35, 259.15, 258.95, 258.55, 
    258.75, 258.85, 258.55, 258.25, 258.35, 257.55, 257.35, 257.45, 257.55, 
    257.25, 257.35, 257.15, 256.85, 256.65, 256.15, 256.45, 256.15, 256.25, 
    256.15, 255.95, 255.85, 255.75, 256.55, 255.85, 256.45, 256.65, 257.15, 
    255.55, 256.35, 258.05, 257.35, 257.25, 257.45, 257.75, 257.95, 257.75, 
    258.25, 258.85, 259.65, 259.85, 260.35, 260.35, 259.75, 259.25, 258.35, 
    258.85, 259.35, 257.35, 258.05, 258.15, 257.25, 257.65, 257.55, 257.45, 
    256.85, 257.45, 257.45, 257.15, 257.05, 256.55, 256.85, 256.35, 256.35, 
    256.25, 256.25, 255.75, 255.85, 255.95, 256.35, 256.45, 256.65, 256.85, 
    257.15, 256.85, 256.35, 256.25, 256.05, 255.85, 255.85, 256.15, 256.15, 
    256.05, 255.85, 255.75, 255.75, 255.85, 255.95, 256.15, 256.75, 256.95, 
    257.15, 257.45, 257.25, 257.75, 257.55, 257.05, 256.95, 256.85, 257.15, 
    257.25, 257.25, 257.45, 257.35, 257.55, 257.45, 257.25, 257.05, 257.25, 
    257.55, 257.75, 258.25, 258.45, 258.85, 258.95, 259.05, 259.25, 259.95, 
    259.85, 259.75, 259.75, 259.75, 259.75, 259.55, 259.65, 259.55, 259.65, 
    259.75, 260.05, 260.15, 259.95, 260.05, 259.85, 259.75, 259.65, 259.35, 
    259.15, 259.15, 259.35, 260.05, 260.75, 261.05, 260.85, 260.85, 260.45, 
    260.85, 260.95, 260.85, 260.45, 260.55, 260.55, 259.95, 260.15, 260.45, 
    261.25, 261.45, 260.95, 260.65, 260.95, 261.35, 261.05, 261.85, 262.25, 
    262.35, 262.45, 262.45, 263.15, 262.45, 263.55, 264.65, 265.05, 265.45, 
    265.85, 265.95, 266.15, 266.75, 266.55, 266.45, 266.35, 265.95, 264.15, 
    264.25, 265.05, 264.45, 264.55, 265.45, 266.35, 266.55, 266.45, 266.95, 
    267.45, 267.45, 267.45, 268.25, 269.05, 268.55, 268.55, 268.25, 267.65, 
    267.55, 267.35, 267.75, 266.65, 266.85, 267.35, 268.35, 268.75, 266.95, 
    268.05, 268.65, 269.35, 269.55, 269.55, 269.45, 269.05, 268.55, 268.35, 
    267.75, 267.45, 267.85, 267.95, 267.95, 267.55, 267.05, 266.45, 266.25, 
    266.85, 267.35, 267.45, 267.55, 267.65, 267.15, 267.15, 267.45, 267.55, 
    267.85, 267.95, 268.25, 268.15, 268.15, 268.25, 268.25, 268.35, 268.35, 
    268.55, 268.95, 269.15, 269.45, 269.85, 270.25, 270.65, 270.75, 271.25, 
    271.75, 271.85, 270.85, 270.05, 270.25, 271.05, 270.35, 269.75, 269.55, 
    269.35, 269.45, 269.55, 269.25, 268.95, 268.15, 268.35, 269.15, 268.45, 
    268.15, 267.75, 267.85, 267.85, 268.55, 268.75, 268.55, 268.55, 269.35, 
    268.85, 269.15, 269.35, 269.45, 269.15, 269.25, 269.05, 269.05, 269.35, 
    269.45, 269.35, 268.95, 269.05, 268.65, 268.05, 268.05, 267.85, 267.65, 
    267.35, 267.15, 266.85, 266.65, 266.55, 266.25, 266.25, 264.55, 262.75, 
    262.15, 261.75, 261.15, 260.75, 261.15, 260.55, 260.55, 259.95, 260.15, 
    260.05, 259.25, 259.25, 259.85, 260.35, 260.55, 260.75, 260.75, 262.15, 
    262.65, 262.95, 262.35, 262.65, 262.85, 263.15, 263.45, 264.65, 264.55, 
    264.95, 265.35, 265.25, 265.65, 266.15, 265.55, 265.55, 266.15, 266.55, 
    267.55, 267.85, 269.95, 270.15, 269.95, 269.75, 269.45, 269.75, 269.85, 
    270.05, 270.05, 270.05, 270.25, 270.35, 270.25, 270.55, 270.35, 270.25, 
    269.95, 269.85, 269.65, 269.35, 269.15, 268.95, 269.05, 269.05, 268.95, 
    269.35, 269.45, 269.65, 269.75, 270.05, 270.35, 270.85, 271.65, 271.85, 
    271.85, 272.05, 271.85, 272.15, 271.95, 271.95, 271.85, 271.75, 271.55, 
    271.25, 270.85, 270.35, 269.75, 269.55, 270.05, 270.05, 270.05, 269.65, 
    269.65, 269.75, 269.75, 270.05, 270.35, 270.05, 270.35, 270.05, 269.95, 
    269.95, 269.75, 269.75, 269.15, 268.65, 268.05, 267.55, 267.55, 266.85, 
    267.65, 267.45, 267.65, 267.95, 268.25, 268.75, 268.65, 268.85, 269.45, 
    268.95, 269.45, 269.25, 268.95, 268.85, 268.65, 268.75, 268.25, 268.15, 
    268.15, 268.15, 267.65, 267.45, 267.15, 267.15, 267.65, 267.65, 267.55, 
    267.55, 267.25, 267.45, 267.65, 268.05, 268.55, 268.45, 269.35, 268.85, 
    268.65, 267.75, 266.95, 266.65, 265.95, 266.25, 266.05, 265.05, 264.55, 
    264.15, 263.65, 263.45, 263.75, 263.75, 264.25, 264.05, 263.85, 264.15, 
    264.15, 264.15, 264.15, 264.25, 264.55, 265.05, 265.45, 265.65, 265.65, 
    265.75, 265.65, 265.65, 265.55, 265.55, 265.45, 265.45, 265.45, 265.35, 
    265.25, 265.25, 265.05, 264.55, 264.45, 264.55, 264.55, 264.75, 265.05, 
    265.55, 264.85, 265.45, 265.65, 265.45, 264.85, 264.85, 265.15, 265.25, 
    265.05, 265.25, 265.05, 264.65, 264.25, 263.95, 263.95, 263.85, 264.05, 
    264.05, 264.05, 264.45, 264.75, 264.95, 264.95, 264.85, 264.75, 264.75, 
    264.65, 265.25, 265.55, 265.95, 266.15, 266.05, 266.05, 265.95, 265.95, 
    265.85, 266.05, 266.25, 266.45, 266.75, 266.85, 266.95, 267.25, 267.65, 
    268.35, 268.75, 268.25, 268.95, 268.85, 268.85, 268.75, 268.75, 268.45, 
    268.35, 268.15, 267.85, 267.55, 267.45, 267.35, 267.25, 267.55, 267.45, 
    267.75, 267.65, 267.65, 267.85, 267.35, 268.55, 268.85, 269.05, 269.35, 
    269.45, 269.85, 270.25, 270.25, 270.25, 270.25, 270.25, 270.05, 269.95, 
    269.85, 269.35, 268.95, 268.35, 268.75, 268.05, 267.45, 267.05, 266.15, 
    266.15, 265.85, 265.75, 265.65, 266.95, 267.35, 267.25, 268.45, 269.55, 
    269.55, 270.05, 269.95, 269.85, 269.45, 269.45, 269.55, 269.65, 269.85, 
    269.45, 269.35, 269.25, 268.95, 268.95, 268.95, 269.35, 269.35, 269.45, 
    270.05, 270.95, 270.95, 271.45, 271.15, 270.85, 270.95, 270.75, 271.35, 
    270.25, 269.65, 269.35, 268.55, 267.95, 267.15, 267.25, 267.25, 267.05, 
    266.75, 266.45, 267.35, 268.15, 268.15, 268.05, 268.15, 268.45, 268.85, 
    269.35, 269.45, 269.05, 269.05, 269.05, 269.15, 268.85, 268.65, 268.75, 
    269.65, 269.55, 268.15, 268.35, 267.75, 265.85, 266.05, 265.65, 265.25, 
    265.95, 266.25, 267.05, 265.65, 265.45, 265.25, 265.45, 266.05, 266.25, 
    266.65, 266.35, 265.65, 264.15, 262.95, 263.05, 263.25, 263.55, 263.55, 
    263.55, 262.95, 262.55, 262.35, 262.45, 262.55, 262.75, 263.15, 262.65, 
    262.65, 262.95, 263.55, 263.65, 264.25, 264.25, 263.65, 263.85, 263.35, 
    263.35, 263.25, 262.85, 262.05, 262.25, 262.05, 262.35, 262.15, 262.25, 
    262.35, 261.45, 261.15, 261.65, 262.05, 262.05, 262.65, 262.45, 263.25, 
    263.85, 265.05, 264.25, 264.85, 265.95, 264.65, 264.25, 264.35, 264.85, 
    264.25, 263.85, 263.95, 264.15, 263.85, 263.65, 263.55, 263.45, 263.55, 
    263.55, 263.85, 263.55, 263.45, 264.05, 264.45, 264.25, 264.45, 264.45, 
    264.45, 264.25, 264.25, 264.15, 264.05, 264.05, 264.25, 264.15, 264.25, 
    264.35, 264.15, 263.75, 263.95, 264.05, 264.15, 264.35, 264.35, 264.85, 
    265.05, 265.15, 265.05, 265.65, 265.95, 266.15, 266.45, 267.75, 267.65, 
    267.55, 267.85, 267.55, 267.55, 266.95, 266.95, 266.25, 265.35, 265.15, 
    264.95, 264.45, 264.45, 264.55, 265.85, 265.05, 265.05, 265.85, 266.65, 
    267.15, 265.75, 265.95, 267.05, 267.45, 267.85, 268.05, 267.95, 267.95, 
    268.15, 268.25, 268.55, 268.55, 268.45, 268.35, 268.25, 268.35, 267.75, 
    267.25, 267.75, 268.15, 268.65, 268.85, 268.25, 269.15, 270.35, 270.35, 
    269.45, 268.75, 268.45, 268.95, 268.95, 268.65, 268.75, 268.35, 268.15, 
    267.45, 266.85, 266.55, 266.75, 267.25, 266.15, 267.55, 268.25, 268.75, 
    268.95, 269.05, 268.95, 268.85, 269.25, 269.35, 269.25, 269.45, 269.15, 
    269.15, 268.85, 269.25, 268.65, 268.45, 268.15, 267.65, 267.35, 266.95, 
    266.95, 266.95, 266.45, 266.35, 266.45, 266.45, 266.55, 266.65, 266.85, 
    267.05, 267.35, 267.55, 267.85, 268.15, 268.45, 268.55, 268.75, 269.05, 
    268.85, 269.25, 269.75, 270.15, 270.75, 270.45, 270.35, 270.35, 270.35, 
    270.55, 270.35, 270.25, 269.95, 270.85, 271.75, 271.55, 272.15, 272.05, 
    272.35, 271.95, 271.75, 271.65, 271.85, 271.65, 271.55, 271.85, 272.35, 
    272.75, 273.15, 273.15, 272.65, 273.15, 272.65, 272.15, 271.75, 271.65, 
    270.95, 270.95, 270.95, 270.95, 270.95, 271.05, 271.75, 271.95, 271.55, 
    271.95, 270.85, 270.85, 269.85, 269.55, 269.25, 268.95, 268.05, 267.75, 
    266.85, 266.15, 265.65, 264.95, 264.95, 265.35, 265.75, 265.55, 265.55, 
    265.95, 266.35, 266.45, 266.85, 266.55, 267.75, 266.75, 266.45, 266.75, 
    267.05, 266.85, 266.95, 267.35, 268.25, 267.95, 268.25, 268.55, 268.95, 
    269.45, 269.85, 269.75, 269.95, 269.95, 270.25, 270.35, 270.35, 270.25, 
    270.55, 270.45, 270.25, 270.15, 270.25, 270.15, 269.95, 269.75, 269.35, 
    269.25, 269.05, 268.75, 268.65, 268.85, 268.45, 268.45, 268.95, 268.85, 
    268.95, 268.75, 268.95, 268.65, 268.65, 269.05, 269.45, 269.65, 270.05, 
    270.05, 269.65, 270.05, 270.05, 270.05, 269.85, 269.85, 270.15, 270.65, 
    270.85, 271.55, 271.75, 271.75, 271.65, 271.65, 271.65, 271.65, 271.05, 
    270.45, 270.15, 270.15, 270.05, 270.25, 270.35, 270.55, 270.75, 270.55, 
    270.25, 270.15, 270.05, 270.45, 270.55, 270.65, 270.95, 270.75, 270.75, 
    270.25, 269.85, 270.45, 270.85, 270.85, 270.75, 270.55, 270.25, 269.85, 
    269.85, 269.65, 269.55, 269.15, 268.85, 268.45, 268.25, 268.45, 268.75, 
    269.15, 269.35, 269.55, 269.35, 269.25, 268.95, 268.85, 268.75, 268.85, 
    269.25, 269.55, 269.55, 269.35, 269.25, 269.25, 269.45, 269.45, 269.65, 
    269.65, 269.65, 269.65, 269.55, 269.85, 269.95, 270.05, 270.15, 270.25, 
    270.35, 270.35, 270.05, 270.25, 270.35, 270.55, 270.45, 270.55, 270.95, 
    271.45, 271.75, 271.75, 271.95, 272.05, 272.15, 271.95, 271.95, 271.95, 
    271.85, 272.15, 272.05, 271.95, 271.85, 271.45, 271.05, 270.95, 270.85, 
    271.05, 270.65, 270.65, 270.35, 270.45, 270.75, 270.75, 270.85, 270.95, 
    271.05, 271.25, 271.15, 271.15, 271.45, 271.15, 271.25, 271.15, 271.05, 
    270.95, 271.05, 271.05, 271.05, 271.15, 271.15, 271.15, 271.05, 271.05, 
    271.15, 271.25, 271.45, 271.65, 271.85, 271.95, 271.65, 272.05, 271.85, 
    271.95, 271.75, 271.75, 271.55, 271.35, 271.25, 271.25, 271.25, 271.35, 
    271.45, 271.85, 271.75, 271.65, 271.75, 271.85, 271.95, 272.05, 271.95, 
    272.35, 271.95, 272.05, 271.95, 271.65, 271.25, 270.75, 270.45, 270.25, 
    270.45, 270.65, 270.85, 271.05, 271.15, 271.15, 271.85, 271.75, 271.75, 
    271.75, 271.85, 271.75, 271.75, 271.85, 271.75, 271.65, 271.65, 272.05, 
    272.15, 272.15, 272.15, 271.95, 271.85, 271.85, 272.05, 271.65, 271.75, 
    271.95, 271.65, 271.45, 271.35, 271.35, 271.35, 271.25, 271.25, 271.35, 
    271.55, 271.65, 271.65, 271.85, 272.25, 272.35, 272.45, 272.65, 272.65, 
    272.65, 272.65, 272.85, 272.75, 272.75, 272.95, 272.95, 272.45, 272.45, 
    272.15, 271.75, 271.25, 271.15, 271.65, 271.95, 271.95, 271.85, 271.55, 
    271.65, 271.75, 271.65, 271.55, 272.25, 271.95, 272.05, 272.15, 271.75, 
    272.05, 272.15, 272.45, 273.15, 273.35, 273.35, 273.15, 273.05, 273.35, 
    273.35, 273.35, 273.15, 272.85, 272.95, 272.55, 271.85, 271.45, 271.35, 
    271.05, 271.65, 271.65, 271.65, 271.65, 271.45, 271.25, 271.25, 270.95, 
    271.05, 271.55, 271.75, 271.75, 272.05, 272.25, 271.85, 271.65, 271.55, 
    271.25, 271.25, 270.95, 270.75, 271.55, 271.95, 272.55, 272.45, 272.75, 
    271.85, 271.95, 271.65, 271.45, 271.25, 271.15, 271.45, 271.05, 271.15, 
    271.05, 271.15, 271.15, 271.35, 271.55, 271.65, 271.55, 271.75, 272.15, 
    272.15, 271.95, 272.15, 272.05, 272.05, 271.85, 271.65, 271.45, 271.15, 
    271.35, 271.35, 270.95, 270.65, 269.85, 269.55, 270.55, 270.05, 270.35, 
    270.35, 270.45, 270.25, 270.05, 270.25, 270.15, 270.35, 270.55, 270.75, 
    270.55, 270.45, 270.55, 270.75, 270.85, 271.05, 270.75, 270.75, 270.85, 
    270.85, 270.45, 269.75, 270.35, 270.45, 270.45, 270.25, 270.35, 270.55, 
    270.55, 270.85, 271.05, 271.15, 271.35, 271.45, 271.55, 271.55, 271.45, 
    271.45, 271.45, 271.35, 271.95, 272.05, 272.05, 271.95, 271.75, 271.65, 
    272.05, 272.05, 271.15, 271.55, 271.25, 271.35, 271.25, 271.75, 271.65, 
    271.65, 271.45, 271.95, 272.25, 272.35, 272.35, 272.15, 272.05, 271.55, 
    271.75, 272.35, 272.55, 271.15, 270.65, 271.75, 270.65, 270.55, 270.85, 
    271.75, 272.15, 272.35, 272.75, 273.35, 273.85, 273.55, 274.35, 274.15, 
    274.35, 274.55, 275.15, 274.05, 273.55, 273.15, 273.25, 273.05, 273.05, 
    272.75, 272.05, 272.35, 272.25, 272.65, 272.55, 272.35, 272.35, 272.95, 
    272.55, 273.75, 273.95, 273.95, 274.65, 273.45, 273.65, 274.15, 274.35, 
    274.65, 274.65, 275.05, 274.25, 274.35, 274.45, 274.35, 274.85, 274.55, 
    274.05, 274.45, 273.75, 273.25, 273.85, 273.85, 272.85, 272.65, 272.55, 
    272.65, 272.95, 273.45, 273.55, 273.35, 274.15, 273.85, 273.75, 274.05, 
    273.35, 273.75, 273.05, 272.85, 272.75, 271.85, 271.05, 271.15, 270.95, 
    270.85, 270.85, 270.65, 272.75, 272.75, 272.95, 273.15, 273.55, 274.05, 
    274.35, 275.55, 274.25, 275.25, 274.25, 276.35, 275.45, 275.45, 275.15, 
    274.75, 275.05, 274.25, 273.35, 273.15, 274.05, 274.35, 274.55, 274.65, 
    275.45, 274.65, 274.35, 274.55, 275.15, 275.35, 274.85, 274.65, 274.45, 
    275.85, 275.75, 274.55, 272.35, 271.75, 271.45, 271.15, 271.75, 271.55, 
    271.25, 271.55, 271.05, 272.55, 273.85, 273.75, 273.85, 274.05, 274.15, 
    274.55, 274.25, 274.15, 273.95, 274.15, 274.55, 274.45, 274.15, 273.85, 
    273.75, 273.55, 273.35, 273.05, 272.75, 272.45, 272.15, 271.95, 272.15, 
    272.15, 272.05, 271.75, 271.25, 271.55, 271.65, 271.45, 271.65, 271.85, 
    271.95, 271.85, 271.95, 272.15, 272.55, 272.65, 272.85, 272.95, 272.75, 
    273.05, 273.35, 273.35, 273.35, 273.45, 273.55, 273.65, 273.65, 273.45, 
    273.45, 273.45, 273.45, 273.45, 273.45, 273.55, 273.65, 273.55, 273.55, 
    273.55, 273.55, 273.35, 273.35, 273.35, 273.35, 273.35, 273.35, 273.45, 
    273.45, 273.35, 273.45, 273.45, 273.55, 273.65, 273.85, 273.45, 273.65, 
    273.35, 273.55, 274.85, 273.65, 274.15, 274.55, 274.15, 275.45, 275.65, 
    275.35, 274.75, 274.15, 274.25, 274.35, 274.15, 273.85, 273.95, 273.85, 
    273.85, 273.85, 273.85, 273.85, 273.85, 273.75, 273.65, 273.45, 273.85, 
    273.85, 273.95, 274.25, 273.75, 273.25, 273.15, 272.95, 272.95, 273.05, 
    273.05, 273.05, 273.65, 273.25, 273.65, 273.45, 273.65, 273.75, 273.95, 
    274.25, 274.15, 274.25, 274.45, 274.65, 274.45, 274.65, 274.55, 275.05, 
    276.05, 275.25, 274.95, 275.05, 275.15, 274.95, 275.05, 275.05, 274.65, 
    274.95, 275.35, 275.05, 274.45, 274.35, 274.15, 274.05, 274.35, 273.55, 
    274.25, 275.05, 274.75, 274.75, 273.55, 273.45, 273.55, 273.15, 273.25, 
    274.25, 273.05, 273.05, 273.05, 272.95, 272.55, 272.55, 272.55, 272.55, 
    272.45, 272.45, 272.25, 272.25, 272.35, 272.25, 272.45, 272.55, 272.55, 
    272.85, 272.75, 272.25, 272.25, 272.05, 272.15, 272.35, 272.35, 272.25, 
    272.75, 273.25, 272.95, 273.25, 273.05, 273.45, 273.35, 273.35, 273.65, 
    274.15, 273.75, 274.55, 274.65, 274.35, 275.35, 274.05, 274.25, 274.25, 
    273.75, 274.05, 273.55, 273.35, 273.65, 273.25, 273.85, 273.55, 273.35, 
    272.95, 272.85, 272.75, 272.45, 272.75, 272.55, 272.05, 272.55, 271.95, 
    272.45, 272.45, 272.35, 272.35, 272.35, 272.75, 272.65, 272.75, 272.85, 
    272.65, 273.05, 273.05, 272.75, 272.55, 272.55, 272.35, 272.85, 272.85, 
    273.25, 273.45, 273.65, 274.05, 273.95, 273.45, 272.95, 273.45, 274.15, 
    274.55, 274.85, 274.95, 274.85, 273.75, 272.85, 272.55, 273.45, 273.55, 
    273.05, 273.05, 271.75, 272.15, 272.05, 272.45, 272.45, 272.65, 273.05, 
    273.15, 273.25, 273.35, 273.75, 274.15, 274.25, 274.25, 274.65, 274.65, 
    273.95, 274.25, 273.95, 273.95, 273.75, 273.35, 273.15, 272.95, 273.25, 
    273.05, 273.15, 273.15, 273.25, 273.15, 273.45, 273.35, 273.55, 273.65, 
    273.35, 273.25, 273.35, 273.45, 273.45, 273.15, 273.15, 273.05, 272.95, 
    272.95, 272.95, 273.05, 272.95, 272.75, 272.95, 272.75, 272.85, 272.85, 
    272.95, 273.15, 273.25, 273.25, 273.35, 273.55, 273.75, 273.75, 273.35, 
    273.45, 273.25, 273.15, 272.95, 272.85, 272.75, 272.35, 272.35, 271.95, 
    272.25, 271.55, 271.75, 271.55, 271.55, 271.65, 271.75, 271.75, 272.15, 
    272.55, 272.85, 273.05, 273.15, 273.55, 273.65, 273.55, 273.75, 273.85, 
    274.05, 274.45, 274.45, 274.55, 274.55, 274.35, 274.45, 274.95, 274.85, 
    274.75, 274.95, 275.15, 274.85, 274.65, 274.65, 274.75, 274.85, 274.75, 
    275.25, 275.25, 275.15, 275.25, 276.25, 276.35, 275.15, 275.65, 276.05, 
    274.75, 274.75, 275.55, 275.15, 274.55, 274.75, 275.35, 274.75, 275.65, 
    276.25, 275.75, 276.75, 275.55, 275.45, 275.15, 274.75, 273.85, 274.25, 
    274.55, 275.35, 275.25, 275.05, 274.85, 274.45, 274.25, 274.35, 274.25, 
    274.05, 274.15, 274.05, 273.85, 273.85, 273.85, 273.85, 273.85, 274.05, 
    273.95, 273.85, 273.75, 273.85, 273.95, 273.95, 273.95, 274.05, 273.85, 
    273.85, 273.85, 273.45, 273.35, 272.55, 272.45, 272.45, 272.35, 272.05, 
    272.35, 272.05, 272.05, 271.75, 272.05, 272.05, 272.45, 272.45, 272.45, 
    272.35, 272.25, 272.75, 272.95, 272.85, 272.55, 272.55, 273.15, 273.35, 
    273.35, 273.15, 273.25, 273.35, 273.45, 273.55, 273.85, 273.85, 273.85, 
    274.15, 274.05, 274.05, 274.05, 274.15, 274.35, 274.65, 275.65, 275.65, 
    275.25, 274.95, 274.25, 274.95, 275.25, 274.95, 275.05, 275.15, 275.45, 
    275.65, 275.95, 275.95, 275.25, 275.45, 275.55, 275.55, 275.45, 275.35, 
    275.25, 275.65, 274.25, 275.35, 274.15, 273.95, 273.65, 273.85, 274.15, 
    274.45, 273.55, 273.45, 273.45, 273.35, 273.25, 273.25, 273.25, 273.15, 
    273.25, 273.15, 273.15, 273.25, 273.35, 273.35, 273.45, 273.25, 273.05, 
    273.15, 273.35, 273.45, 273.45, 273.45, 273.45, 273.55, 273.45, 273.35, 
    273.35, 273.35, 273.35, 273.35, 273.25, 273.15, 273.15, 273.15, 273.35, 
    273.35, 273.35, 273.35, 273.35, 273.45, 273.55, 273.75, 273.45, 273.75, 
    273.65, 273.75, 273.55, 273.65, 273.75, 273.45, 273.65, 273.45, 273.55, 
    273.55, 273.55, 273.55, 273.45, 273.55, 273.55, 273.65, 273.55, 273.55, 
    273.65, 273.55, 273.45, 273.45, 273.45, 273.45, 273.75, 273.75, 273.95, 
    273.85, 274.05, 273.75, 273.65, 273.55, 272.65, 272.75, 272.65, 272.75, 
    272.75, 272.65, 272.85, 272.85, 273.15, 273.55, 273.35, 273.75, 273.75, 
    274.35, 274.55, 274.85, 275.15, 275.35, 275.65, 276.95, 280.15, 279.55, 
    276.45, 276.25, 279.45, 279.15, 276.25, 275.75, 275.45, 275.15, 275.35, 
    275.55, 275.75, 275.85, 275.55, 275.75, 276.35, 276.05, 275.85, 276.25, 
    276.35, 276.05, 275.55, 275.35, 274.65, 274.75, 274.95, 274.95, 275.15, 
    275.05, 275.05, 275.15, 275.25, 275.25, 275.65, 275.85, 275.85, 276.45, 
    275.35, 275.25, 275.05, 275.15, 275.45, 275.55, 275.45, 275.25, 275.35, 
    275.55, 275.65, 275.75, 275.75, 275.55, 275.45, 275.55, 275.25, 275.35, 
    274.35, 274.25, 273.75, 273.55, 273.45, 273.65, 273.95, 274.25, 274.75, 
    274.75, 274.65, 274.55, 275.15, 274.85, 274.95, 275.35, 275.05, 275.45, 
    274.85, 274.45, 274.25, 273.45, 273.65, 273.75, 273.35, 273.15, 272.75, 
    272.75, 272.75, 272.95, 273.25, 273.15, 273.05, 273.15, 273.25, 273.35, 
    273.45, 273.85, 274.25, 274.05, 274.15, 274.15, 273.95, 273.95, 273.65, 
    273.55, 273.55, 273.65, 273.85, 273.35, 273.15, 272.75, 272.35, 272.35, 
    272.85, 272.95, 273.25, 273.55, 273.75, 273.45, 273.75, 273.65, 274.05, 
    274.15, 273.65, 273.85, 274.15, 273.65, 273.25, 273.05, 272.85, 272.65, 
    271.85, 271.95, 272.55, 272.55, 272.65, 272.75, 272.55, 272.35, 272.15, 
    274.35, 272.25, 272.25, 272.75, 273.05, 273.55, 273.45, 274.05, 274.05, 
    273.75, 273.55, 273.55, 274.05, 274.05, 274.15, 274.15, 274.05, 274.15, 
    274.25, 274.25, 274.15, 274.25, 274.35, 274.35, 274.35, 274.45, 274.45, 
    274.55, 274.55, 274.95, 274.85, 274.65, 274.85, 274.95, 274.15, 274.05, 
    273.85, 273.65, 273.05, 272.85, 272.95, 273.25, 273.45, 273.35, 273.35, 
    274.45, 274.95, 273.65, 274.45, 274.45, 274.65, 275.45, 275.05, 274.95, 
    274.95, 275.15, 274.25, 274.05, 273.65, 273.35, 272.75, 275.35, 276.05, 
    277.95, 277.25, 278.05, 278.05, 277.55, 277.15, 276.75, 276.45, 276.25, 
    276.35, 275.75, 275.75, 275.75, 276.05, 275.95, 275.95, 276.75, 276.45, 
    276.15, 276.85, 276.15, 277.05, 276.25, 275.75, 275.55, 275.25, 275.05, 
    275.05, 275.25, 275.95, 278.15, 278.05, 277.75, 278.45, 278.25, 276.85, 
    276.65, 276.75, 276.75, 276.55, 276.45, 276.55, 276.85, 276.35, 275.95, 
    277.05, 277.95, 277.85, 277.65, 276.95, 276.65, 276.55, 276.15, 276.15, 
    276.25, 276.15, 276.35, 276.35, 276.35, 276.05, 276.25, 276.35, 276.25, 
    276.15, 275.95, 275.75, 275.75, 275.65, 275.85, 275.75, 275.65, 275.65, 
    275.65, 275.65, 275.65, 275.55, 275.55, 275.75, 275.65, 275.65, 275.65, 
    275.65, 275.75, 275.85, 275.95, 276.05, 276.25, 276.25, 276.15, 276.15, 
    275.75, 275.75, 275.95, 275.75, 275.65, 275.25, 276.25, 275.65, 276.05, 
    275.55, 275.75, 277.75, 277.15, 277.05, 277.05, 276.95, 276.45, 278.15, 
    278.25, 277.85, 277.55, 277.05, 277.45, 278.05, 278.45, 278.15, 278.45, 
    277.85, 278.45, 278.45, 278.25, 278.65, 277.55, 277.15, 277.75, 277.65, 
    278.05, 277.25, 277.55, 278.25, 278.05, 278.55, 277.55, 278.05, 278.05, 
    277.75, 277.25, 276.95, 277.55, 277.75, 277.15, 277.05, 277.85, 278.15, 
    276.85, 279.15, 277.85, 277.55, 277.35, 277.35, 276.85, 276.75, 277.55, 
    278.25, 278.15, 278.05, 277.15, 278.05, 277.05, 277.55, 277.05, 276.85, 
    276.65, 277.25, 276.85, 277.15, 277.45, 277.15, 277.55, 276.85, 277.25, 
    277.05, 276.65, 275.45, 276.35, 274.85, 274.95, 275.85, 274.85, 274.75, 
    274.85, 274.75, 274.85, 275.15, 275.35, 275.05, 274.95, 274.85, 274.55, 
    274.45, 274.45, 274.45, 274.25, 274.35, 274.25, 274.35, 274.25, 274.25, 
    275.05, 274.65, 275.25, 275.85, 276.15, 276.35, 275.75, 275.45, 275.15, 
    275.95, 276.35, 276.45, 276.05, 276.15, 275.85, 275.65, 275.85, 275.65, 
    275.65, 275.55, 275.35, 275.05, 275.35, 275.75, 276.65, 276.55, 276.45, 
    276.55, 276.65, 276.05, 275.55, 275.45, 275.25, 275.05, 274.65, 274.95, 
    274.85, 274.85, 274.85, 274.55, 273.95, 273.95, 273.95, 274.05, 274.15, 
    274.45, 274.25, 274.15, 273.95, 274.05, 273.85, 273.85, 273.85, 274.05, 
    274.15, 274.05, 274.05, 273.95, 274.05, 273.95, 273.55, 273.35, 272.85, 
    272.85, 272.95, 272.55, 272.95, 273.15, 273.25, 273.15, 273.15, 273.05, 
    272.95, 273.05, 273.65, 273.75, 273.75, 274.55, 274.55, 276.35, 276.05, 
    276.35, 276.25, 276.35, 276.35, 276.25, 276.05, 275.95, 275.85, 275.85, 
    273.95, 273.95, 275.05, 275.45, 277.25, 276.85, 276.65, 276.65, 278.05, 
    278.65, 277.75, 278.65, 278.65, 278.55, 278.75, 279.05, 278.75, 278.45, 
    277.55, 277.95, 277.15, 277.15, 277.15, 277.05, 277.05, 276.65, 276.45, 
    276.15, 275.35, 274.85, 277.15, 277.05, 275.25, 275.25, 275.25, 275.55, 
    275.45, 275.35, 275.45, 275.25, 275.25, 275.45, 275.35, 275.15, 275.25, 
    275.15, 275.15, 275.05, 275.25, 275.25, 275.35, 275.35, 275.65, 275.55, 
    275.65, 275.85, 275.95, 275.85, 275.95, 275.95, 275.95, 275.75, 275.75, 
    275.55, 275.55, 275.65, 275.45, 275.35, 275.35, 275.55, 275.55, 275.45, 
    275.35, 275.35, 275.45, 275.45, 275.85, 276.05, 275.05, 274.85, 275.05, 
    274.85, 274.95, 275.15, 275.15, 275.25, 275.55, 275.15, 274.65, 274.75, 
    274.65, 274.65, 274.45, 274.45, 274.15, 274.25, 274.15, 273.95, 274.15, 
    274.15, 274.25, 274.25, 274.25, 274.35, 274.45, 274.65, 274.65, 274.45, 
    274.45, 274.25, 274.25, 274.05, 273.95, 274.05, 273.85, 273.95, 273.95, 
    274.05, 274.05, 274.05, 273.95, 274.05, 274.05, 273.95, 273.75, 273.55, 
    273.45, 273.75, 274.05, 274.05, 274.15, 274.25, 274.25, 274.25, 274.05, 
    274.25, 274.55, 274.65, 274.65, 274.75, 275.05, 275.25, 275.45, 275.35, 
    275.35, 275.75, 275.75, 275.95, 276.05, 276.55, 276.35, 276.25, 275.25, 
    274.75, 274.65, 274.65, 274.55, 275.25, 275.05, 274.95, 275.35, 275.55, 
    275.75, 275.45, 275.35, 275.25, 275.15, 275.15, 274.95, 274.95, 274.85, 
    275.05, 275.35, 276.15, 276.65, 276.85, 277.35, 277.05, 277.45, 278.35, 
    278.15, 278.75, 278.15, 278.05, 279.35, 278.25, 276.45, 276.85, 275.05, 
    274.75, 275.35, 274.75, 274.45, 275.05, 275.45, 277.25, 277.65, 277.15, 
    277.55, 277.25, 277.65, 278.15, 278.55, 277.95, 277.05, 276.35, 276.15, 
    276.15, 276.25, 276.55, 276.65, 276.35, 276.25, 276.45, 276.05, 276.05, 
    276.05, 276.25, 276.35, 276.05, 275.85, 275.95, 276.05, 275.95, 276.75, 
    276.35, 276.45, 276.95, 277.35, 277.05, 277.05, 276.35, 275.85, 275.55, 
    275.25, 275.05, 275.15, 275.05, 274.75, 275.55, 275.25, 275.05, 275.15, 
    274.95, 275.15, 274.95, 274.85, 274.85, 274.75, 274.75, 274.85, 275.15, 
    275.05, 274.55, 274.15, 273.35, 273.45, 273.35, 273.05, 273.15, 273.25, 
    272.45, 272.25, 272.15, 272.15, 272.25, 272.35, 272.45, 272.55, 272.85, 
    272.85, 273.35, 273.25, 273.35, 273.65, 273.75, 273.75, 273.75, 274.15, 
    273.55, 273.75, 273.75, 273.75, 274.05, 274.15, 273.85, 273.05, 273.15, 
    273.65, 273.75, 273.95, 273.75, 273.65, 273.45, 273.35, 273.35, 273.25, 
    273.35, 273.45, 273.45, 273.35, 273.45, 273.65, 274.35, 275.15, 275.25, 
    275.55, 276.05, 276.45, 276.15, 276.05, 275.65, 275.85, 275.65, 276.15, 
    276.05, 275.75, 276.35, 276.55, 276.55, 276.75, 277.15, 277.65, 277.55, 
    277.65, 277.75, 278.15, 277.85, 277.25, 276.25, 275.45, 274.95, 274.95, 
    275.05, 275.35, 275.45, 275.75, 276.15, 275.95, 276.15, 275.45, 275.35, 
    275.45, 275.35, 275.25, 274.65, 274.45, 273.75, 273.35, 273.25, 272.95, 
    272.95, 272.85, 272.85, 272.25, 272.45, 272.55, 272.85, 272.65, 272.85, 
    273.05, 273.15, 273.15, 273.25, 273.35, 273.35, 273.35, 273.45, 273.35, 
    273.25, 273.35, 273.45, 273.35, 273.45, 273.35, 273.25, 273.45, 273.45, 
    273.45, 273.45, 273.55, 273.55, 273.55, 273.55, 273.85, 274.05, 274.05, 
    274.15, 274.15, 274.45, 274.15, 274.05, 273.85, 273.85, 274.25, 274.45, 
    274.65, 274.85, 274.85, 274.75, 274.75, 274.45, 274.55, 274.45, 274.45, 
    274.45, 274.55, 274.55, 274.55, 274.45, 274.55, 274.45, 274.55, 274.55, 
    274.45, 274.65, 274.75, 274.95, 275.15, 275.05, 275.35, 275.35, 275.65, 
    275.55, 275.55, 275.45, 275.25, 275.55, 275.35, 275.55, 275.35, 275.15, 
    275.05, 275.35, 275.35, 274.65, 273.65, 272.95, 273.45, 272.85, 272.45, 
    273.05, 273.45, 273.85, 274.05, 273.85, 273.85, 273.35, 273.65, 273.55, 
    273.25, 272.95, 272.65, 272.45, 272.55, 272.55, 272.75, 272.75, 272.45, 
    272.65, 273.45, 273.75, 273.45, 273.55, 273.55, 273.55, 273.45, 273.25, 
    273.25, 273.35, 273.35, 273.15, 272.95, 273.05, 273.15, 273.25, 273.25, 
    273.15, 273.15, 273.15, 273.35, 273.45, 273.45, 273.45, 273.65, 273.85, 
    273.95, 273.95, 274.15, 274.95, 274.65, 274.95, 274.85, 274.45, 274.65, 
    274.25, 274.25, 273.85, 273.65, 273.75, 273.45, 273.25, 273.15, 273.25, 
    273.35, 273.75, 274.25, 274.05, 274.05, 274.55, 274.45, 274.65, 274.75, 
    275.35, 275.55, 275.45, 275.45, 275.55, 275.55, 275.55, 275.55, 275.55, 
    275.45, 274.95, 274.95, 274.55, 274.55, 274.15, 274.25, 274.35, 274.25, 
    274.35, 274.25, 275.25, 274.95, 274.65, 274.95, 275.25, 275.25, 275.15, 
    274.45, 274.85, 275.25, 274.85, 274.65, 274.25, 274.15, 274.05, 273.95, 
    273.95, 273.95, 273.75, 273.65, 273.35, 273.35, 273.35, 273.35, 273.05, 
    272.95, 273.25, 273.45, 273.35, 273.45, 273.55, 273.85, 273.85, 273.55, 
    273.75, 273.85, 273.45, 273.25, 273.45, 273.55, 273.25, 273.25, 273.25, 
    273.65, 273.25, 273.15, 273.15, 273.35, 273.35, 273.25, 273.45, 274.05, 
    274.35, 274.95, 275.25, 274.85, 274.55, 275.05, 275.65, 275.95, 275.65, 
    275.65, 275.65, 275.25, 275.25, 275.15, 275.35, 274.95, 275.15, 274.95, 
    275.05, 274.85, 274.85, 274.95, 275.35, 275.35, 275.35, 275.65, 275.65, 
    275.65, 275.55, 275.15, 275.55, 275.05, 274.85, 274.55, 274.55, 274.25, 
    274.05, 274.15, 273.95, 274.25, 273.95, 273.95, 274.35, 274.55, 274.55, 
    274.55, 274.75, 274.85, 275.15, 275.25, 275.35, 275.45, 275.95, 276.05, 
    275.65, 275.35, 275.05, 274.75, 274.25, 274.05, 274.25, 274.45, 274.25, 
    274.25, 274.05, 274.45, 274.85, 275.15, 275.25, 275.45, 275.35, 275.45, 
    275.55, 276.45, 275.95, 276.15, 276.35, 276.15, 275.85, 275.75, 275.95, 
    275.95, 276.15, 276.35, 276.55, 276.55, 276.45, 276.45, 276.15, 276.15, 
    276.05, 276.35, 276.15, 276.05, 275.75, 276.75, 276.55, 276.75, 276.55, 
    276.75, 276.95, 277.35, 277.55, 276.85, 277.45, 276.75, 276.45, 276.15, 
    276.45, 276.15, 275.15, 274.75, 275.65, 275.95, 275.55, 276.15, 276.15, 
    275.65, 275.85, 277.15, 276.75, 277.75, 278.25, 276.95, 276.55, 276.05, 
    276.25, 277.05, 277.05, 277.25, 276.15, 276.65, 276.25, 276.15, 276.65, 
    276.65, 276.85, 276.65, 276.45, 276.25, 275.95, 275.95, 275.75, 275.75, 
    275.25, 275.35, 276.15, 276.35, 276.45, 276.45, 275.95, 275.45, 275.15, 
    275.05, 274.95, 274.95, 274.95, 274.15, 274.15, 274.25, 274.05, 273.45, 
    273.65, 274.75, 275.25, 275.25, 275.45, 275.65, 275.55, 275.85, 276.05, 
    276.55, 276.95, 276.25, 276.15, 276.45, 276.65, 276.55, 276.35, 276.05, 
    275.95, 275.95, 275.95, 275.95, 275.65, 275.65, 275.75, 275.55, 275.75, 
    275.85, 275.55, 275.35, 275.65, 275.85, 276.15, 276.25, 276.55, 276.05, 
    275.55, 275.95, 275.35, 277.15, 276.85, 276.25, 276.65, 276.55, 276.75, 
    277.25, 277.35, 277.05, 276.75, 276.55, 276.45, 276.55, 276.75, 276.45, 
    276.95, 277.05, 275.95, 276.15, 276.15, 276.05, 276.15, 275.95, 276.15, 
    276.05, 276.05, 275.85, 275.55, 276.05, 275.85, 276.05, 276.05, 275.75, 
    275.55, 275.75, 275.75, 275.45, 275.75, 275.75, 275.55, 275.55, 275.35, 
    275.35, 275.35, 275.15, 275.35, 275.95, 276.35, 275.65, 275.25, 275.25, 
    275.85, 274.85, 274.75, 274.65, 274.65, 274.45, 274.65, 275.15, 275.05, 
    274.65, 274.75, 274.75, 274.75, 275.05, 275.05, 274.85, 275.05, 275.85, 
    276.45, 275.95, 276.55, 276.35, 276.65, 276.45, 276.25, 276.35, 276.35, 
    276.35, 276.45, 276.35, 276.55, 276.45, 276.45, 276.45, 276.35, 276.65, 
    276.55, 276.45, 276.45, 276.15, 276.25, 276.45, 276.55, 276.85, 276.65, 
    276.45, 278.35, 275.55, 274.95, 273.85, 274.45, 275.35, 274.75, 274.05, 
    274.25, 273.45, 273.85, 273.95, 273.95, 274.35, 274.15, 274.45, 274.85, 
    276.05, 275.65, 274.85, 275.05, 275.85, 275.45, 275.65, 275.95, 275.95, 
    275.65, 275.75, 276.55, 275.25, 276.85, 276.35, 275.75, 275.75, 275.75, 
    275.75, 275.75, 276.55, 276.35, 276.35, 275.35, 275.45, 275.95, 275.65, 
    275.65, 274.85, 274.75, 274.55, 274.65, 274.95, 275.15, 274.15, 274.75, 
    274.45, 274.25, 274.35, 274.25, 274.35, 274.25, 274.25, 274.35, 274.25, 
    274.25, 274.35, 274.25, 274.25, 274.25, 274.25, 274.45, 274.35, 274.35, 
    274.25, 274.25, 274.25, 274.15, 274.15, 274.15, 274.15, 274.05, 273.95, 
    273.85, 273.85, 273.75, 273.65, 273.55, 273.85, 274.25, 274.25, 274.45, 
    274.65, 274.85, 275.05, 274.95, 274.85, 274.45, 274.25, 274.35, 273.95, 
    273.95, 274.25, 275.45, 275.65, 275.65, 275.15, 275.15, 275.15, 275.45, 
    275.55, 275.55, 275.95, 276.15, 276.15, 276.35, 276.15, 275.65, 275.75, 
    275.65, 275.85, 275.95, 275.95, 275.95, 275.85, 276.15, 276.05, 276.35, 
    276.25, 275.75, 275.65, 274.95, 274.15, 274.25, 274.35, 274.35, 274.25, 
    274.25, 274.55, 274.45, 274.65, 274.85, 275.25, 275.45, 275.35, 275.55, 
    276.25, 275.55, 275.55, 275.85, 275.65, 275.45, 274.95, 274.65, 274.95, 
    275.45, 275.05, 274.85, 274.75, 274.85, 275.05, 275.45, 275.55, 275.55, 
    275.45, 275.75, 275.85, 276.05, 275.85, 275.75, 275.75, 275.75, 275.75, 
    275.75, 275.85, 275.95, 276.15, 276.15, 275.95, 276.05, 276.25, 276.35, 
    276.35, 276.65, 276.25, 275.95, 275.95, 276.05, 276.45, 276.55, 276.55, 
    276.45, 276.25, 276.05, 275.95, 276.25, 276.15, 276.35, 276.55, 276.15, 
    276.05, 275.95, 276.15, 276.35, 276.25, 276.45, 276.45, 276.35, 276.15, 
    276.25, 276.25, 276.55, 276.65, 276.55, 276.55, 276.15, 276.25, 276.55, 
    276.75, 276.95, 276.85, 276.35, 275.95, 276.75, 276.95, 276.55, 276.65, 
    276.75, 276.75, 276.95, 277.55, 276.75, 276.55, 276.35, 276.15, 275.75, 
    275.45, 275.15, 275.05, 274.85, 274.75, 274.65, 274.85, 274.85, 274.85, 
    274.75, 274.85, 274.65, 274.45, 274.45, 274.65, 274.65, 274.75, 274.65, 
    274.65, 274.55, 274.65, 275.05, 275.35, 275.25, 275.15, 275.05, 274.75, 
    274.65, 274.45, 274.45, 274.25, 273.95, 273.85, 273.85, 273.75, 273.75, 
    274.15, 273.75, 273.55, 273.45, 273.45, 273.55, 273.35, 273.25, 273.15, 
    273.15, 273.75, 274.05, 273.95, 274.25, 274.05, 273.75, 273.75, 273.65, 
    273.55, 273.55, 273.85, 273.95, 274.05, 274.15, 274.15, 274.25, 274.45, 
    274.15, 274.15, 273.75, 273.55, 273.35, 273.45, 273.65, 273.65, 274.15, 
    274.25, 274.25, 274.05, 274.25, 274.55, 274.85, 274.75, 274.75, 274.65, 
    274.55, 274.45, 273.85, 274.25, 274.25, 273.85, 273.85, 273.85, 273.95, 
    273.75, 273.85, 273.95, 273.95, 273.85, 273.95, 273.85, 273.95, 273.75, 
    273.55, 273.55, 273.65, 273.45, 273.55, 273.35, 273.35, 273.05, 273.05, 
    272.85, 272.25, 272.05, 272.15, 272.25, 272.65, 272.45, 272.55, 272.65, 
    272.45, 271.95, 271.65, 271.25, 271.65, 271.75, 271.55, 271.95, 272.05, 
    271.85, 271.35, 271.25, 271.45, 271.15, 271.15, 271.45, 271.35, 271.25, 
    271.05, 271.25, 271.15, 271.15, 271.45, 271.25, 271.85, 271.65, 272.05, 
    272.25, 271.95, 272.05, 272.15, 272.25, 272.05, 272.05, 272.05, 272.05, 
    272.05, 272.05, 271.55, 271.65, 271.45, 271.75, 271.55, 271.65, 272.15, 
    271.55, 272.55, 272.55, 272.75, 272.55, 272.25, 272.55, 272.45, 272.65, 
    272.65, 272.85, 272.85, 272.95, 273.15, 273.45, 273.65, 273.35, 273.45, 
    272.45, 272.25, 271.85, 271.45, 271.15, 270.85, 270.85, 271.05, 271.15, 
    271.25, 271.25, 271.25, 271.05, 270.55, 271.25, 270.95, 270.95, 271.15, 
    271.15, 271.35, 271.15, 271.15, 271.35, 271.45, 271.65, 271.55, 271.15, 
    271.55, 272.05, 272.25, 272.65, 272.75, 272.65, 272.25, 272.65, 272.15, 
    272.15, 272.25, 271.85, 270.25, 271.95, 271.65, 271.95, 272.15, 271.45, 
    270.75, 270.85, 270.85, 271.05, 271.05, 271.05, 271.15, 271.35, 270.85, 
    270.15, 271.05, 270.95, 272.25, 272.15, 271.65, 271.45, 271.15, 271.05, 
    271.45, 271.65, 272.05, 271.85, 272.25, 272.05, 272.25, 271.35, 270.65, 
    270.75, 271.55, 271.95, 271.65, 271.95, 272.25, 271.85, 271.95, 272.35, 
    272.45, 272.75, 272.75, 272.95, 272.85, 272.45, 272.25, 272.35, 273.35, 
    272.45, 273.15, 273.35, 273.05, 273.45, 273.05, 273.25, 272.75, 272.65, 
    272.75, 273.15, 273.35, 273.65, 273.85, 273.65, 273.75, 273.65, 273.85, 
    273.95, 273.95, 273.35, 273.35, 273.45, 273.55, 273.75, 273.85, 273.85, 
    273.85, 274.05, 274.25, 274.25, 274.25, 274.35, 274.45, 274.35, 274.35, 
    274.65, 274.35, 274.25, 274.05, 273.95, 272.95, 273.25, 273.45, 272.45, 
    272.85, 272.15, 272.55, 272.45, 272.25, 272.35, 272.55, 272.95, 272.85, 
    272.75, 272.85, 272.75, 272.35, 272.15, 272.65, 272.35, 272.15, 272.15, 
    272.85, 272.55, 273.05, 273.55, 272.95, 272.95, 272.55, 272.25, 271.45, 
    271.65, 272.85, 271.95, 271.05, 271.65, 271.65, 273.05, 273.15, 273.15, 
    273.25, 274.45, 274.55, 274.95, 275.05, 274.95, 274.75, 274.85, 274.85, 
    274.75, 274.65, 274.75, 274.75, 274.75, 274.95, 274.85, 274.75, 274.65, 
    274.05, 273.85, 273.95, 273.65, 273.65, 273.35, 273.05, 273.25, 273.25, 
    272.95, 272.75, 272.95, 273.15, 273.05, 273.15, 273.05, 272.95, 272.85, 
    272.05, 272.35, 271.95, 271.75, 271.05, 270.55, 268.75, 267.85, 268.15, 
    268.45, 268.85, 269.15, 269.05, 269.55, 268.35, 268.25, 267.45, 267.65, 
    267.45, 268.45, 267.25, 267.85, 268.35, 267.75, 267.15, 268.35, 268.55, 
    268.75, 269.45, 269.45, 269.45, 269.65, 269.75, 269.75, 269.75, 269.75, 
    270.05, 270.35, 270.75, 270.85, 270.95, 270.95, 271.15, 271.35, 271.65, 
    271.85, 272.25, 272.55, 272.95, 273.05, 273.05, 273.65, 273.45, 273.35, 
    273.55, 272.15, 271.35, 270.65, 270.05, 269.55, 269.05, 268.55, 268.15, 
    268.05, 267.75, 267.45, 267.25, 267.25, 267.45, 267.65, 267.65, 267.65, 
    267.95, 267.95, 268.35, 268.25, 268.25, 268.15, 268.15, 268.25, 268.15, 
    268.25, 268.25, 268.45, 268.35, 268.45, 268.35, 268.15, 268.15, 268.45, 
    268.35, 268.95, 269.45, 270.55, 270.75, 271.45, 271.35, 271.15, 270.75, 
    270.75, 271.15, 271.15, 271.15, 271.15, 271.35, 271.35, 271.25, 270.65, 
    271.15, 271.15, 271.05, 270.05, 271.45, 271.45, 271.35, 271.65, 271.85, 
    271.75, 272.15, 272.25, 272.15, 272.65, 272.15, 272.65, 272.15, 272.05, 
    272.15, 272.35, 272.75, 273.05, 273.15, 273.35, 273.05, 273.35, 273.55, 
    273.35, 273.75, 274.05, 274.15, 274.15, 274.05, 274.15, 274.25, 274.15, 
    274.35, 274.35, 274.55, 274.45, 274.25, 274.35, 274.35, 274.35, 274.45, 
    274.45, 274.45, 274.35, 274.35, 274.45, 274.45, 274.45, 274.55, 274.55, 
    274.55, 274.55, 274.55, 274.25, 274.25, 274.35, 274.25, 274.15, 274.45, 
    274.05, 274.15, 274.15, 274.15, 273.85, 273.85, 273.55, 273.45, 272.75, 
    273.25, 272.45, 272.55, 272.75, 272.75, 272.65, 272.65, 272.85, 272.85, 
    272.75, 272.85, 273.25, 272.05, 270.55, 269.95, 269.05, 268.45, 268.25, 
    267.95, 267.75, 268.05, 268.15, 268.35, 268.15, 268.45, 267.85, 267.65, 
    267.55, 267.35, 267.35, 265.95, 265.85, 266.45, 266.85, 266.75, 266.85, 
    267.25, 268.25, 270.25, 270.75, 270.65, 270.85, 271.15, 271.25, 271.35, 
    271.35, 271.35, 271.65, 271.75, 271.85, 271.85, 271.75, 271.95, 272.15, 
    272.25, 272.45, 272.65, 272.75, 272.95, 273.05, 273.25, 273.15, 273.15, 
    273.45, 273.75, 274.65, 273.55, 273.15, 272.75, 272.15, 271.55, 271.25, 
    271.35, 271.45, 271.65, 271.55, 271.45, 271.45, 271.95, 272.25, 273.05, 
    273.15, 272.95, 273.45, 272.75, 272.95, 272.35, 273.75, 273.25, 273.65, 
    273.25, 273.25, 273.45, 272.95, 273.15, 272.15, 272.05, 271.45, 271.65, 
    272.05, 271.35, 272.05, 271.15, 271.15, 271.95, 271.85, 272.15, 271.95, 
    271.85, 272.15, 272.85, 273.15, 272.75, 272.65, 272.45, 272.25, 272.55, 
    272.25, 271.85, 272.15, 272.75, 272.45, 272.25, 272.45, 272.35, 272.65, 
    272.95, 273.05, 272.75, 272.95, 273.05, 273.05, 272.85, 272.45, 272.45, 
    272.55, 272.35, 272.45, 272.35, 272.45, 272.55, 272.65, 272.55, 272.75, 
    272.95, 273.15, 273.35, 273.55, 273.45, 273.45, 273.45, 273.65, 274.05, 
    273.85, 273.95, 273.95, 273.95, 273.95, 274.05, 274.15, 274.15, 273.95, 
    273.95, 274.05, 273.85, 273.45, 273.25, 273.55, 273.35, 273.55, 273.65, 
    273.55, 273.35, 273.15, 273.15, 273.05, 272.85, 272.85, 272.75, 272.45, 
    272.45, 272.45, 272.35, 272.35, 272.85, 273.35, 273.35, 273.55, 273.45, 
    273.45, 272.85, 272.65, 272.25, 273.45, 273.35, 273.35, 274.25, 273.95, 
    274.15, 274.35, 274.25, 273.95, 273.95, 273.85, 274.25, 274.25, 274.35, 
    274.35, 274.25, 274.15, 273.75, 273.65, 273.35, 273.25, 273.85, 273.65, 
    273.65, 272.85, 272.65, 273.05, 273.05, 272.95, 272.95, 273.05, 273.35, 
    273.75, 273.55, 273.65, 273.45, 273.55, 273.45, 273.25, 273.25, 273.55, 
    273.35, 273.25, 273.75, 273.55, 273.05, 272.85, 272.85, 272.45, 272.35, 
    272.05, 271.85, 271.65, 271.15, 271.55, 271.25, 271.45, 270.95, 271.45, 
    271.45, 271.55, 271.65, 271.95, 271.95, 271.85, 272.05, 271.65, 271.75, 
    271.35, 271.85, 271.55, 271.45, 271.25, 271.35, 271.25, 270.75, 270.65, 
    270.75, 270.85, 270.75, 270.75, 270.65, 269.85, 269.45, 269.45, 269.15, 
    269.05, 269.25, 269.55, 269.45, 269.05, 269.45, 269.45, 269.15, 269.35, 
    269.45, 269.85, 270.55, 270.05, 269.75, 269.35, 269.35, 268.95, 268.45, 
    268.35, 267.95, 267.55, 267.45, 267.05, 266.65, 266.45, 265.95, 265.65, 
    264.95, 264.35, 264.05, 263.95, 263.95, 263.55, 263.65, 263.75, 263.75, 
    263.95, 263.75, 263.65, 263.45, 263.45, 263.75, 263.95, 264.45, 264.35, 
    264.55, 265.05, 265.15, 265.45, 264.95, 264.65, 264.75, 264.35, 264.25, 
    264.65, 264.65, 264.85, 265.05, 265.25, 265.55, 265.95, 266.45, 266.25, 
    266.55, 266.65, 267.25, 267.85, 268.45, 269.65, 270.35, 269.95, 269.65, 
    270.35, 271.95, 271.85, 270.35, 270.95, 270.05, 270.05, 269.65, 269.05, 
    268.95, 270.25, 269.75, 269.95, 269.75, 270.35, 270.65, 271.05, 270.55, 
    270.35, 270.85, 270.75, 270.45, 270.25, 270.55, 270.45, 270.25, 268.75, 
    269.15, 269.75, 270.15, 269.65, 269.85, 270.25, 270.55, 270.05, 270.35, 
    269.45, 269.75, 270.05, 269.25, 270.05, 269.35, 269.45, 269.85, 270.25, 
    268.25, 269.95, 270.45, 270.75, 270.75, 270.25, 270.25, 270.15, 269.65, 
    269.55, 270.05, 270.65, 271.15, 271.65, 271.05, 271.25, 269.75, 268.95, 
    270.15, 270.75, 270.55, 270.35, 270.35, 270.25, 269.85, 269.65, 269.75, 
    269.75, 269.75, 269.65, 269.55, 269.55, 269.55, 269.45, 269.05, 269.15, 
    269.05, 268.85, 268.95, 268.95, 269.15, 269.45, 269.85, 269.55, 270.05, 
    270.15, 269.65, 270.05, 269.95, 270.85, 270.55, 270.05, 269.75, 269.65, 
    268.85, 268.35, 269.85, 268.65, 268.95, 270.15, 269.25, 269.25, 269.45, 
    269.75, 269.35, 269.45, 268.05, 268.55, 268.85, 268.05, 267.35, 267.45, 
    267.25, 266.85, 267.25, 268.75, 268.75, 269.05, 267.75, 268.85, 268.75, 
    268.65, 268.75, 268.65, 267.25, 267.45, 266.85, 266.95, 267.45, 268.75, 
    269.05, 269.45, 270.45, 270.35, 269.95, 270.35, 270.75, 271.05, 271.75, 
    272.45, 272.95, 273.05, 273.35, 273.35, 273.35, 272.75, 273.05, 273.05, 
    273.15, 273.25, 273.45, 273.45, 273.35, 272.95, 273.05, 272.75, 272.45, 
    272.55, 272.45, 272.15, 271.65, 271.55, 271.65, 271.65, 271.45, 271.15, 
    270.95, 271.15, 271.05, 271.25, 271.25, 271.35, 271.45, 271.65, 271.75, 
    271.75, 271.85, 271.65, 271.65, 271.85, 271.55, 271.55, 271.85, 271.75, 
    271.85, 272.05, 272.35, 272.15, 272.25, 272.15, 272.35, 272.35, 272.35, 
    272.45, 272.05, 272.45, 271.85, 272.55, 272.75, 272.75, 272.75, 272.75, 
    272.85, 272.85, 273.05, 273.15, 273.15, 273.15, 273.15, 273.15, 273.15, 
    273.15, 273.15, 273.15, 273.25, 273.25, 273.25, 273.15, 273.15, 273.15, 
    273.15, 273.35, 273.55, 273.45, 273.55, 273.45, 273.35, 273.35, 273.25, 
    273.15, 273.15, 273.05, 272.95, 272.75, 272.75, 272.85, 272.95, 273.05, 
    273.15, 272.95, 272.95, 273.05, 273.35, 273.55, 273.35, 273.15, 271.45, 
    270.35, 269.15, 268.55, 268.05, 267.45, 266.65, 266.75, 266.35, 266.45, 
    266.55, 266.05, 265.75, 265.45, 265.65, 265.85, 265.95, 266.15, 266.35, 
    266.75, 267.15, 267.35, 267.85, 268.15, 268.55, 268.95, 269.15, 269.35, 
    269.45, 269.45, 269.45, 268.85, 268.15, 267.55, 267.35, 267.35, 267.05, 
    266.75, 266.75, 266.35, 265.85, 265.95, 265.75, 265.45, 265.25, 265.45, 
    265.15, 264.95, 265.05, 265.05, 265.05, 264.85, 264.95, 264.75, 264.65, 
    264.55, 264.55, 264.65, 264.35, 264.55, 264.45, 264.45, 264.45, 264.55, 
    264.65, 264.65, 264.55, 264.45, 264.35, 264.25, 263.95, 264.15, 263.85, 
    263.65, 263.65, 263.55, 263.45, 263.75, 263.95, 263.75, 263.25, 263.05, 
    262.95, 262.25, 262.05, 261.95, 262.05, 261.75, 261.75, 261.85, 261.95, 
    261.65, 261.45, 261.75, 261.45, 261.45, 261.65, 261.45, 261.35, 261.55, 
    261.35, 261.45, 261.95, 261.85, 261.95, 261.95, 261.75, 261.55, 261.65, 
    261.75, 262.05, 262.65, 262.35, 262.85, 262.85, 263.25, 262.55, 263.15, 
    262.85, 262.65, 262.55, 262.65, 262.55, 262.75, 262.95, 263.35, 263.65, 
    263.65, 263.85, 264.15, 264.45, 264.45, 264.25, 264.55, 264.45, 264.45, 
    264.65, 264.55, 264.75, 264.55, 264.85, 264.85, 265.35, 265.65, 265.75, 
    265.75, 266.05, 265.95, 266.15, 266.15, 265.55, 265.55, 264.85, 264.35, 
    263.15, 262.95, 263.25, 263.55, 263.65, 264.45, 264.95, 265.45, 265.65, 
    266.45, 266.35, 267.55, 268.25, 268.55, 269.15, 269.35, 269.65, 269.75, 
    269.95, 269.85, 270.35, 270.35, 270.55, 270.75, 271.15, 271.35, 271.55, 
    271.35, 271.25, 270.75, 270.65, 271.15, 270.55, 270.05, 269.85, 269.35, 
    268.95, 268.55, 268.15, 267.65, 267.25, 266.85, 266.95, 267.05, 267.15, 
    267.05, 266.75, 266.05, 266.05, 265.95, 265.95, 265.65, 265.75, 265.95, 
    266.15, 264.25, 262.85, 263.05, 263.35, 263.55, 262.55, 262.85, 262.75, 
    263.15, 263.15, 263.45, 263.25, 263.35, 263.65, 263.95, 264.45, 265.35, 
    266.05, 266.45, 266.65, 266.55, 266.95, 267.05, 267.15, 267.25, 267.35, 
    267.35, 267.45, 267.45, 267.85, 267.75, 267.75, 267.25, 268.15, 267.65, 
    267.55, 267.15, 266.85, 267.85, 268.15, 267.85, 268.35, 267.15, 269.05, 
    269.85, 269.85, 270.35, 269.75, 271.15, 271.25, 270.95, 270.95, 270.85, 
    270.75, 270.35, 270.25, 269.85, 269.55, 270.35, 270.15, 269.75, 269.65, 
    269.15, 268.95, 269.05, 269.05, 269.05, 269.05, 269.25, 269.15, 269.15, 
    268.85, 268.35, 268.25, 268.25, 268.15, 267.45, 267.65, 266.75, 266.45, 
    266.15, 266.85, 266.45, 266.15, 266.15, 266.55, 266.45, 264.65, 264.85, 
    264.45, 264.65, 265.25, 265.55, 265.55, 265.35, 265.25, 265.15, 264.35, 
    264.75, 264.75, 264.65, 265.85, 265.65, 265.15, 266.15, 265.55, 265.55, 
    266.65, 265.95, 265.05, 265.15, 265.35, 266.55, 265.95, 266.25, 266.05, 
    266.45, 266.25, 266.35, 266.65, 266.95, 267.35, 265.35, 265.65, 264.65, 
    263.95, 262.85, 262.55, 263.55, 263.55, 263.15, 262.75, 263.05, 262.75, 
    262.75, 262.95, 263.15, 262.95, 262.65, 262.55, 262.55, 262.35, 262.25, 
    262.35, 262.55, 262.95, 263.25, 263.75, 264.15, 263.85, 263.65, 264.25, 
    264.05, 263.75, 263.65, 263.25, 262.65, 262.45, 262.25, 262.25, 261.15, 
    260.65, 260.05, 259.75, 259.65, 259.85, 259.95, 260.15, 260.35, 260.25, 
    260.25, 260.45, 260.45, 260.75, 260.65, 260.35, 260.05, 259.45, 259.95, 
    260.45, 259.85, 260.35, 260.25, 260.35, 260.65, 260.95, 261.05, 261.05, 
    260.75, 260.65, 259.95, 260.15, 260.05, 260.35, 260.25, 260.85, 261.85, 
    262.25, 261.65, 261.55, 261.15, 261.15, 261.75, 261.45, 260.75, 259.45, 
    259.15, 258.75, 258.45, 258.35, 258.15, 257.85, 257.65, 257.85, 258.15, 
    258.15, 258.15, 257.85, 257.45, 257.15, 257.35, 257.45, 257.05, 257.45, 
    257.25, 257.05, 257.35, 257.35, 257.75, 257.95, 258.25, 258.35, 259.05, 
    259.05, 259.05, 258.75, 258.95, 259.15, 258.85, 258.45, 258.05, 257.15, 
    256.65, 257.95, 257.75, 257.95, 258.95, 259.55, 259.05, 260.15, 260.25, 
    260.05, 259.05, 260.25, 260.65, 261.15, 260.85, 262.45, 262.95, 263.35, 
    263.25, 263.85, 263.85, 263.65, 263.95, 263.75, 264.55, 264.75, 264.75, 
    265.65, 265.25, 266.15, 266.25, 266.15, 264.95, 265.35, 265.75, 265.95, 
    266.75, 266.75, 266.85, 266.65, 266.55, 266.55, 266.15, 265.65, 266.15, 
    265.95, 265.65, 263.65, 261.95, 262.15, 263.25, 263.05, 261.35, 263.35, 
    262.35, 261.75, 262.15, 263.25, 264.05, 264.25, 263.75, 263.85, 263.65, 
    263.75, 263.75, 263.35, 263.55, 262.55, 262.95, 262.95, 261.45, 261.15, 
    261.55, 263.15, 264.25, 264.75, 265.15, 265.45, 265.45, 266.05, 266.55, 
    266.75, 267.35, 267.05, 267.15, 267.65, 267.75, 267.35, 268.05, 268.55, 
    268.95, 268.65, 268.75, 268.45, 268.25, 267.55, 266.45, 265.55, 265.15, 
    264.75, 264.45, 263.85, 264.25, 264.25, 262.55, 263.05, 264.05, 265.15, 
    264.55, 264.45, 264.65, 264.75, 264.45, 264.75, 264.95, 264.35, 264.05, 
    262.95, 262.35, 262.45, 262.45, 262.95, 262.25, 262.15, 262.75, 262.45, 
    262.85, 262.95, 262.85, 260.65, 262.15, 262.75, 263.05, 263.35, 263.75, 
    264.55, 265.05, 265.75, 266.15, 266.25, 266.75, 266.95, 267.05, 266.55, 
    267.25, 266.85, 266.55, 266.55, 267.15, 267.35, 268.15, 268.35, 268.75, 
    268.85, 268.75, 269.25, 269.25, 269.15, 269.15, 269.15, 268.75, 268.35, 
    268.45, 268.35, 268.55, 267.45, 268.65, 268.95, 269.75, 269.85, 270.35, 
    270.85, 271.05, 271.05, 271.25, 271.05, 270.85, 270.65, 270.65, 270.35, 
    270.35, 270.05, 270.75, 271.05, 271.05, 270.85, 271.15, 271.15, 271.25, 
    271.45, 271.55, 271.55, 271.85, 271.65, 270.75, 270.55, 270.95, 271.15, 
    271.55, 271.05, 270.55, 270.15, 270.05, 269.85, 269.45, 269.75, 270.15, 
    270.25, 270.85, 267.85, 269.45, 267.45, 267.85, 268.45, 268.95, 269.05, 
    269.25, 269.25, 269.45, 269.35, 269.25, 268.85, 268.05, 268.85, 269.45, 
    269.25, 268.55, 268.45, 268.45, 268.25, 268.25, 266.35, 265.75, 264.35, 
    265.45, 267.35, 266.65, 265.45, 265.35, 265.35, 265.05, 265.05, 265.35, 
    265.75, 266.25, 267.15, 267.55, 267.15, 267.05, 267.05, 266.45, 266.95, 
    266.95, 266.35, 266.05, 265.55, 265.25, 265.05, 264.35, 263.65, 263.65, 
    262.25, 261.65, 261.45, 260.95, 260.25, 259.95, 259.95, 260.15, 259.95, 
    258.35, 258.15, 258.35, 258.75, 259.35, 259.55, 260.15, 260.05, 259.95, 
    259.65, 259.35, 259.05, 259.05, 259.05, 259.25, 259.45, 259.65, 259.35, 
    259.05, 258.55, 258.55, 257.45, 257.95, 257.15, 257.55, 257.55, 257.55, 
    257.35, 257.75, 258.65, 258.55, 259.35, 259.05, 259.65, 259.35, 259.35, 
    259.65, 260.05, 260.05, 260.85, 261.45, 261.85, 262.55, 262.55, 262.65, 
    262.85, 262.95, 263.35, 263.55, 263.85, 264.15, 264.45, 264.55, 264.75, 
    264.95, 265.05, 265.25, 265.45, 265.25, 265.95, 267.05, 268.55, 267.85, 
    266.85, 267.95, 268.45, 268.65, 268.65, 268.05, 268.15, 267.75, 267.55, 
    268.05, 268.85, 268.15, 267.75, 267.25, 267.55, 268.55, 268.85, 269.25, 
    270.25, 269.95, 271.15, 271.55, 271.55, 271.45, 271.45, 271.45, 271.35, 
    271.45, 271.75, 272.45, 272.55, 272.55, 272.55, 272.55, 272.55, 272.55, 
    272.45, 272.55, 272.55, 272.45, 272.45, 272.45, 272.45, 272.15, 272.25, 
    272.35, 272.45, 272.35, 272.35, 272.35, 272.35, 272.35, 272.25, 272.35, 
    272.25, 272.05, 272.25, 272.05, 272.15, 272.05, 271.95, 272.05, 272.15, 
    272.15, 272.15, 272.05, 272.15, 272.15, 272.15, 272.15, 272.15, 272.15, 
    272.15, 272.05, 271.95, 271.65, 271.75, 271.55, 271.35, 271.25, 271.25, 
    271.25, 271.15, 271.35, 271.65, 271.55, 271.25, 271.15, 271.05, 271.15, 
    271.05, 270.95, 270.95, 270.85, 271.25, 270.95, 270.95, 271.25, 271.15, 
    271.15, 271.05, 271.15, 269.45, 270.95, 271.05, 271.15, 271.25, 271.25, 
    271.25, 271.35, 271.35, 271.25, 271.25, 270.95, 270.75, 270.95, 270.65, 
    270.85, 270.75, 270.75, 270.75, 271.25, 270.95, 270.55, 270.75, 270.85, 
    271.25, 270.95, 270.75, 270.85, 270.55, 270.45, 269.85, 269.85, 270.35, 
    270.85, 271.45, 271.45, 271.35, 271.45, 271.25, 271.55, 271.55, 271.45, 
    271.55, 271.45, 271.35, 271.35, 271.35, 271.15, 270.95, 271.45, 271.25, 
    271.45, 271.15, 270.95, 270.15, 270.05, 271.05, 271.55, 272.15, 272.05, 
    272.05, 271.95, 271.85, 271.55, 271.65, 271.65, 272.15, 272.45, 272.45, 
    272.45, 272.35, 272.35, 272.35, 272.25, 272.35, 272.25, 272.15, 271.95, 
    271.75, 271.65, 271.35, 271.25, 271.05, 270.55, 270.15, 270.05, 269.35, 
    268.15, 266.35, 264.65, 263.35, 263.05, 262.75, 262.65, 262.65, 262.25, 
    261.75, 261.55, 261.25, 260.75, 260.05, 259.85, 259.75, 259.45, 259.15, 
    259.05, 258.95, 258.55, 258.75, 258.75, 258.65, 258.35, 258.15, 258.15, 
    258.15, 257.75, 257.75, 257.55, 257.55, 257.95, 257.75, 257.45, 258.15, 
    257.45, 257.75, 257.25, 257.25, 257.95, 257.65, 257.65, 257.65, 257.85, 
    258.25, 258.15, 259.15, 260.75, 261.45, 262.15, 263.15, 263.75, 264.45, 
    265.35, 266.05, 267.05, 267.95, 268.65, 269.75, 270.35, 270.35, 270.75, 
    269.85, 270.05, 268.05, 267.55, 266.25, 265.75, 266.55, 267.85, 268.85, 
    268.25, 268.25, 267.25, 266.75, 266.15, 265.75, 265.05, 264.35, 263.65, 
    263.15, 262.35, 262.05, 261.95, 261.95, 262.15, 262.25, 262.35, 262.95, 
    263.25, 262.75, 262.45, 261.75, 261.75, 261.45, 261.05, 260.45, 258.75, 
    259.15, 257.35, 258.05, 258.05, 259.25, 259.75, 259.05, 259.25, 259.15, 
    258.75, 258.85, 259.05, 259.95, 260.35, 260.65, 261.45, 262.55, 263.35, 
    264.05, 265.05, 265.95, 267.35, 268.55, 269.65, 271.35, 270.35, 269.25, 
    268.45, 268.05, 267.45, 267.05, 266.85, 266.45, 266.15, 265.55, 265.55, 
    265.55, 265.95, 266.35, 266.55, 265.85, 266.45, 267.25, 267.45, 265.85, 
    264.65, 263.65, 262.95, 263.65, 264.35, 264.05, 263.65, 263.75, 263.05, 
    262.95, 263.25, 263.55, 262.95, 262.75, 262.35, 262.45, 262.15, 262.15, 
    261.75, 261.15, 261.05, 260.65, 260.75, 260.95, 260.15, 259.85, 260.15, 
    259.75, 260.85, 260.95, 261.15, 261.45, 261.75, 261.85, 262.25, 262.15, 
    262.35, 262.05, 261.35, 260.35, 258.65, 257.85, 257.55, 257.35, 257.15, 
    257.05, 257.45, 257.55, 258.15, 258.55, 258.25, 257.75, 257.75, 257.25, 
    256.95, 256.95, 256.95, 256.35, 256.15, 255.95, 256.05, 255.75, 255.85, 
    255.65, 255.45, 255.75, 255.65, 255.95, 255.35, 254.85, 255.85, 255.75, 
    257.45, 258.65, 258.55, 258.45, 259.05, 258.85, 258.95, 258.55, 257.05, 
    256.15, 256.25, 256.55, 256.45, 255.75, 255.65, 255.05, 256.25, 256.65, 
    257.45, 256.55, 257.15, 257.65, 258.45, 259.35, 260.05, 260.05, 261.25, 
    266.55, 267.45, 267.05, 266.45, 266.75, 267.85, 266.25, 266.65, 265.15, 
    264.35, 264.05, 263.45, 263.55, 263.45, 263.95, 263.85, 263.85, 263.15, 
    262.65, 262.95, 262.85, 263.65, 263.05, 263.35, 264.35, 264.35, 264.35, 
    264.15, 263.95, 264.25, 264.75, 266.15, 266.15, 264.55, 264.85, 265.15, 
    265.15, 264.95, 264.65, 264.95, 265.15, 264.75, 264.65, 264.95, 265.35, 
    265.55, 265.55, 266.15, 265.05, 264.45, 265.75, 265.85, 266.85, 267.95, 
    268.75, 269.45, 270.35, 270.35, 270.45, 270.25, 270.35, 270.45, 270.25, 
    270.05, 270.15, 269.95, 270.25, 269.95, 270.25, 270.15, 269.95, 270.05, 
    270.25, 269.75, 269.95, 269.65, 269.55, 269.75, 269.45, 269.45, 269.65, 
    268.35, 268.25, 268.55, 268.35, 268.15, 268.15, 268.25, 268.15, 267.75, 
    266.15, 266.75, 266.55, 266.65, 267.05, 267.95, 268.05, 268.45, 268.65, 
    269.05, 269.65, 269.85, 270.25, 271.25, 271.15, 270.65, 270.55, 270.45, 
    270.05, 270.35, 270.85, 270.75, 270.35, 270.65, 270.75, 270.55, 270.05, 
    269.45, 269.45, 269.65, 269.75, 269.45, 269.05, 268.75, 268.55, 268.75, 
    268.95, 268.75, 268.95, 269.25, 269.35, 269.15, 269.35, 269.15, 269.15, 
    269.15, 269.25, 269.35, 269.45, 269.45, 269.05, 269.15, 269.25, 269.45, 
    269.45, 269.55, 269.75, 270.25, 270.65, 270.85, 270.75, 270.65, 270.55, 
    270.65, 270.55, 270.55, 270.55, 270.55, 270.55, 270.55, 270.35, 270.55, 
    270.45, 270.45, 270.45, 270.25, 270.55, 270.55, 270.45, 270.35, 270.55, 
    270.55, 270.75, 270.75, 270.55, 270.35, 270.35, 270.25, 270.15, 270.15, 
    270.25, 270.65, 270.85, 270.65, 270.65, 270.65, 270.65, 270.65, 270.55, 
    270.45, 270.55, 270.55, 270.35, 270.25, 269.95, 269.85, 269.85, 269.55, 
    269.55, 269.55, 269.45, 269.45, 269.15, 268.75, 268.35, 268.15, 267.85, 
    268.55, 268.95, 269.05, 268.75, 268.55, 268.55, 268.35, 268.05, 267.45, 
    267.45, 267.45, 266.95, 267.25, 267.35, 267.95, 268.05, 266.85, 267.15, 
    266.35, 266.25, 266.25, 266.35, 266.75, 266.55, 266.45, 267.15, 266.75, 
    266.55, 266.55, 266.65, 267.95, 267.35, 267.05, 267.25, 267.65, 268.45, 
    267.55, 267.15, 267.55, 267.45, 267.55, 267.95, 268.55, 267.95, 268.75, 
    269.45, 268.55, 269.15, 268.75, 268.45, 268.35, 268.65, 268.75, 268.65, 
    269.05, 269.25, 269.35, 269.65, 269.45, 269.65, 270.15, 270.85, 271.15, 
    271.25, 271.35, 271.45, 271.65, 271.65, 272.05, 272.15, 272.25, 272.35, 
    272.25, 272.25, 272.15, 272.15, 272.25, 272.35, 272.25, 272.25, 272.25, 
    272.25, 272.15, 271.95, 271.65, 271.15, 271.95, 271.75, 271.65, 271.55, 
    271.45, 270.85, 270.75, 270.35, 270.25, 270.45, 270.35, 270.35, 271.05, 
    270.35, 269.25, 268.35, 268.15, 268.05, 268.95, 268.75, 268.45, 268.55, 
    268.05, 270.35, 270.15, 269.75, 269.45, 269.45, 269.25, 269.35, 269.15, 
    269.05, 269.15, 269.35, 268.95, 268.05, 267.95, 268.05, 268.15, 267.75, 
    267.55, 267.25, 267.35, 267.25, 267.05, 267.05, 267.05, 266.75, 266.75, 
    266.75, 266.55, 266.65, 266.75, 266.75, 266.15, 267.05, 267.45, 267.35, 
    267.65, 268.05, 268.45, 269.05, 270.35, 270.95, 271.05, 270.95, 270.95, 
    270.95, 271.15, 271.15, 270.95, 271.05, 270.95, 271.25, 270.75, 270.75, 
    270.45, 270.35, 270.05, 269.95, 269.95, 269.65, 269.35, 268.75, 268.35, 
    268.15, 268.25, 268.45, 268.55, 268.75, 269.15, 268.95, 269.05, 268.25, 
    267.65, 266.95, 266.65, 266.65, 266.25, 265.05, 263.85, 262.45, 261.95, 
    260.35, 259.75, 261.45, 261.25, 261.95, 262.55, 263.65, 263.55, 263.65, 
    263.35, 263.25, 263.65, 263.95, 263.95, 264.25, 264.45, 264.35, 263.85, 
    264.05, 263.95, 262.95, 262.95, 262.55, 262.35, 261.95, 262.55, 262.15, 
    262.75, 263.25, 263.45, 263.45, 263.55, 263.85, 264.05, 264.35, 264.55, 
    263.95, 264.45, 264.35, 265.05, 265.25, 264.65, 264.35, 264.15, 264.35, 
    263.95, 263.45, 263.85, 262.45, 261.85, 262.65, 262.55, 261.95, 262.05, 
    262.35, 262.55, 262.65, 262.75, 262.35, 261.15, 261.85, 262.15, 261.75, 
    262.35, 262.65, 262.15, 262.35, 262.55, 263.45, 262.25, 262.35, 262.45, 
    262.95, 262.55, 262.55, 262.25, 262.05, 261.65, 262.95, 260.45, 260.35, 
    260.95, 261.15, 260.25, 261.15, 261.35, 261.85, 261.55, 261.75, 261.55, 
    261.55, 261.65, 262.15, 262.85, 262.55, 262.75, 262.15, 261.85, 261.45, 
    261.75, 261.35, 260.35, 259.95, 260.75, 261.55, 260.95, 260.65, 260.45, 
    261.15, 260.95, 260.25, 259.85, 260.05, 260.05, 260.25, 260.55, 260.35, 
    260.15, 259.95, 259.45, 258.65, 258.55, 259.05, 259.45, 259.35, 260.15, 
    260.75, 260.85, 260.65, 260.45, 259.95, 259.25, 259.25, 259.25, 259.35, 
    259.35, 259.15, 259.25, 259.45, 259.75, 259.95, 260.25, 260.55, 260.65, 
    260.45, 259.95, 259.85, 260.25, 259.65, 259.65, 259.55, 259.25, 259.05, 
    259.35, 259.35, 259.15, 259.05, 260.15, 260.95, 261.15, 260.65, 260.75, 
    260.55, 260.25, 259.95, 259.55, 258.85, 258.45, 256.85, 257.15, 256.05, 
    256.05, 256.15, 255.35, 254.15, 253.55, 253.75, 255.75, 255.05, 256.05, 
    258.15, 258.35, 258.25, 257.85, 257.65, 257.65, 257.05, 256.25, 254.85, 
    255.05, 254.65, 253.95, 254.55, 255.85, 255.35, 255.55, 255.45, 255.85, 
    256.75, 257.05, 257.65, 258.65, 259.05, 259.65, 259.95, 259.75, 259.75, 
    259.25, 258.55, 258.25, 257.45, 256.75, 255.85, 255.15, 254.55, 253.95, 
    253.45, 253.15, 252.85, 252.65, 252.75, 252.95, 252.85, 252.65, 252.15, 
    251.95, 252.05, 252.75, 253.05, 253.75, 253.55, 253.95, 254.35, 254.45, 
    255.15, 255.55, 255.95, 256.35, 256.85, 256.55, 257.35, 257.45, 257.25, 
    257.35, 257.25, 256.75, 256.35, 256.05, 255.95, 255.85, 255.75, 255.65, 
    255.35, 255.85, 255.65, 256.35, 256.75, 257.15, 257.65, 258.05, 258.25, 
    257.85, 258.15, 259.15, 261.35, 262.45, 263.15, 263.35, 262.75, 261.95, 
    261.65, 261.55, 261.85, 262.05, 262.35, 262.65, 262.45, 262.85, 262.45, 
    261.45, 260.25, 259.45, 259.35, 259.15, 259.45, 259.55, 259.85, 258.85, 
    259.35, 259.45, 259.45, 258.85, 258.35, 258.55, 258.45, 259.05, 258.65, 
    258.85, 258.45, 258.25, 258.15, 259.35, 259.85, 260.05, 259.75, 259.25, 
    259.85, 260.25, 258.75, 257.75, 258.25, 256.35, 256.75, 257.25, 257.15, 
    257.15, 257.65, 257.55, 257.85, 258.85, 258.65, 258.35, 257.55, 258.55, 
    258.55, 258.85, 258.85, 259.35, 259.95, 259.15, 258.95, 258.95, 258.45, 
    257.55, 257.45, 257.35, 256.65, 257.65, 257.15, 257.95, 258.25, 258.45, 
    258.35, 258.35, 257.85, 256.75, 255.95, 257.15, 257.45, 257.75, 257.55, 
    257.65, 256.25, 258.15, 258.75, 259.15, 258.95, 258.75, 258.65, 257.65, 
    257.65, 257.35, 258.05, 257.65, 257.35, 257.55, 257.45, 257.25, 257.35, 
    258.35, 258.55, 258.25, 258.25, 258.05, 257.85, 257.65, 258.05, 258.15, 
    257.85, 257.45, 258.25, 258.65, 258.65, 258.15, 258.55, 258.05, 256.25, 
    258.25, 258.25, 257.25, 258.15, 259.05, 258.75, 259.25, 258.95, 259.35, 
    259.75, 259.05, 259.45, 259.35, 258.85, 258.35, 258.05, 257.55, 256.85, 
    256.95, 257.15, 257.25, 256.75, 256.25, 256.05, 255.75, 255.75, 255.05, 
    253.95, 254.75, 254.15, 254.75, 255.05, 253.85, 255.55, 254.55, 254.35, 
    254.65, 253.15, 254.05, 254.35, 255.05, 254.15, 254.75, 254.45, 254.15, 
    253.95, 253.85, 253.65, 253.55, 253.55, 254.05, 255.25, 255.25, 255.85, 
    257.35, 258.95, 258.45, 258.55, 257.95, 257.65, 257.95, 257.85, 257.95, 
    257.95, 257.55, 258.25, 258.65, 259.45, 259.85, 260.25, 259.45, 260.05, 
    260.15, 260.75, 259.95, 260.25, 260.15, 261.95, 263.45, 265.15, 263.95, 
    262.75, 262.55, 262.15, 261.85, 261.75, 261.65, 260.55, 260.35, 260.55, 
    260.75, 261.55, 261.25, 260.95, 260.55, 260.95, 260.95, 260.75, 260.95, 
    261.15, 261.65, 261.35, 261.05, 260.75, 260.45, 260.55, 260.65, 260.65, 
    260.25, 260.05, 258.75, 258.75, 256.55, 257.35, 258.55, 258.25, 258.85, 
    258.85, 258.85, 259.75, 259.85, 259.15, 258.85, 259.05, 258.45, 259.25, 
    259.25, 259.25, 258.45, 258.05, 257.75, 257.65, 257.85, 258.95, 258.55, 
    258.65, 258.85, 259.15, 259.25, 259.15, 259.35, 259.35, 259.45, 259.45, 
    259.55, 259.95, 259.75, 259.65, 260.25, 260.55, 260.75, 261.85, 262.55, 
    264.85, 263.75, 264.75, 265.65, 266.25, 265.95, 266.75, 267.45, 267.55, 
    267.75, 268.25, 268.45, 269.35, 269.85, 269.75, 269.25, 269.85, 269.85, 
    270.05, 269.65, 269.55, 269.55, 269.45, 269.05, 269.15, 268.15, 267.85, 
    267.95, 268.15, 267.65, 267.65, 267.95, 267.85, 267.55, 267.85, 267.95, 
    267.75, 267.85, 267.65, 267.65, 267.25, 267.25, 267.15, 267.25, 267.55, 
    267.65, 267.95, 266.55, 266.35, 267.35, 268.15, 269.05, 269.55, 269.15, 
    269.15, 269.35, 269.55, 269.05, 269.05, 269.05, 269.05, 268.75, 268.35, 
    268.65, 268.85, 268.75, 268.55, 268.75, 268.75, 268.55, 268.25, 267.75, 
    268.35, 267.55, 267.65, 267.65, 268.25, 267.45, 267.65, 267.05, 266.85, 
    267.05, 266.75, 266.75, 266.55, 266.25, 265.55, 266.95, 266.55, 266.15, 
    265.85, 265.85, 265.85, 266.05, 265.25, 265.15, 263.25, 265.45, 261.75, 
    261.25, 262.45, 262.55, 262.85, 263.85, 263.45, 264.25, 264.85, 265.25, 
    264.65, 264.05, 264.75, 264.65, 264.05, 264.05, 263.75, 263.85, 263.55, 
    262.85, 263.75, 263.55, 262.25, 262.45, 262.65, 262.35, 263.05, 263.35, 
    264.05, 264.25, 264.65, 264.95, 265.15, 265.55, 265.95, 266.65, 266.65, 
    267.75, 267.85, 268.55, 268.75, 268.95, 269.45, 269.45, 269.35, 270.05, 
    270.25, 270.35, 270.15, 270.25, 270.55, 270.65, 270.85, 270.65, 270.65, 
    270.95, 271.05, 271.25, 271.45, 271.55, 271.25, 270.45, 270.75, 270.45, 
    270.25, 268.75, 268.85, 268.25, 267.05, 266.25, 265.45, 265.25, 264.75, 
    266.25, 267.45, 267.75, 267.05, 266.05, 266.65, 267.15, 267.35, 266.55, 
    267.65, 267.55, 268.05, 266.45, 266.25, 265.25, 264.95, 264.65, 264.35, 
    264.45, 264.25, 264.55, 264.55, 264.75, 264.95, 265.45, 265.95, 266.15, 
    266.35, 266.75, 267.45, 267.75, 267.35, 267.95, 266.95, 267.65, 268.85, 
    267.85, 265.75, 265.75, 264.25, 263.85, 262.75, 262.95, 263.85, 264.15, 
    264.45, 264.65, 265.35, 266.45, 267.75, 268.15, 267.85, 268.05, 267.95, 
    267.95, 267.75, 267.55, 267.75, 267.35, 267.75, 269.05, 269.25, 268.85, 
    268.15, 267.95, 267.75, 268.25, 267.75, 266.75, 266.15, 264.75, 265.25, 
    266.25, 266.35, 266.65, 269.75, 270.75, 269.15, 269.95, 270.55, 269.45, 
    268.55, 270.05, 270.45, 271.15, 271.65, 267.15, 267.15, 267.05, 266.25, 
    269.05, 269.05, 269.55, 268.95, 268.75, 267.65, 267.45, 266.95, 266.75, 
    266.65, 266.85, 267.45, 267.65, 267.65, 267.95, 268.35, 268.65, 268.65, 
    268.95, 268.85, 268.75, 268.45, 268.65, 267.95, 266.45, 265.15, 264.55, 
    263.85, 263.45, 262.95, 262.35, 261.45, 261.25, 261.15, 261.15, 261.35, 
    261.45, 261.85, 261.45, 261.15, 260.75, 260.75, 260.45, 260.35, 260.05, 
    259.65, 259.25, 257.75, 257.55, 257.65, 257.35, 257.25, 257.35, 258.45, 
    258.75, 258.85, 259.05, 259.55, 260.05, 260.75, 260.95, 259.55, 259.65, 
    259.75, 259.75, 259.75, 260.55, 260.75, 260.45, 260.35, 260.45, 260.15, 
    259.85, 260.05, 259.35, 260.35, 260.55, 260.05, 259.75, 260.65, 261.45, 
    261.95, 262.75, 262.75, 263.55, 264.45, 262.25, 260.65, 259.15, 258.15, 
    255.95, 255.15, 254.45, 252.65, 251.85, 251.45, 250.95, 250.05, 250.15, 
    249.95, 250.15, 249.65, 249.95, 249.45, 248.15, 247.95, 248.65, 249.55, 
    248.85, 248.05, 248.65, 248.05, 247.95, 247.65, 248.35, 248.85, 248.75, 
    249.55, 250.65, 251.35, 251.85, 252.75, 253.95, 254.85, 255.85, 256.85, 
    255.25, 254.35, 252.85, 251.15, 249.95, 248.55, 247.65, 247.75, 248.05, 
    248.55, 249.65, 249.65, 250.45, 250.35, 250.55, 249.75, 249.25, 249.95, 
    247.95, 247.35, 247.35, 247.45, 246.75, 246.45, 246.35, 246.05, 245.75, 
    245.15, 244.95, 244.75, 243.85, 242.65, 241.85, 241.05, 240.05, 239.85, 
    239.85, 240.25, 240.35, 240.35, 241.05, 241.25, 241.65, 241.85, 241.65, 
    241.85, 242.25, 242.25, 242.25, 242.25, 242.25, 242.55, 243.05, 243.25, 
    243.35, 243.65, 243.95, 244.35, 244.25, 243.15, 243.15, 243.35, 242.95, 
    243.25, 243.65, 245.05, 243.75, 243.35, 242.95, 243.45, 244.35, 243.25, 
    243.35, 244.75, 244.55, 243.85, 242.85, 243.55, 242.75, 242.85, 243.05, 
    243.45, 244.35, 244.45, 245.45, 246.55, 249.65, 250.25, 249.65, 252.35, 
    251.55, 250.85, 248.35, 247.95, 247.65, 249.05, 248.15, 247.25, 246.85, 
    246.55, 245.35, 245.45, 246.55, 245.35, 245.15, 244.95, 243.95, 244.05, 
    243.65, 243.45, 243.75, 244.05, 245.65, 246.45, 247.65, 248.75, 245.85, 
    245.75, 245.95, 245.65, 245.05, 245.85, 246.15, 245.45, 245.95, 245.75, 
    245.65, 245.25, 245.05, 244.95, 245.75, 246.55, 246.55, 247.05, 246.85, 
    247.75, 249.15, 249.45, 249.75, 249.95, 250.85, 250.85, 250.55, 250.45, 
    250.85, 251.05, 250.65, 249.85, 249.75, 249.65, 249.25, 248.45, 248.25, 
    248.45, 248.25, 247.95, 247.85, 248.65, 248.25, 248.85, 248.95, 249.15, 
    249.15, 249.35, 249.45, 249.05, 248.95, 249.45, 249.75, 249.95, 250.05, 
    249.95, 250.25, 249.85, 249.25, 249.35, 249.05, 249.35, 249.75, 250.15, 
    250.25, 249.65, 249.35, 249.75, 249.05, 249.25, 249.45, 249.85, 249.45, 
    249.15, 248.75, 248.85, 247.85, 247.95, 248.35, 248.15, 248.65, 248.95, 
    249.05, 248.55, 247.35, 248.95, 248.85, 247.95, 248.25, 248.65, 248.25, 
    246.85, 248.25, 248.45, 247.85, 246.75, 248.15, 249.25, 248.75, 249.45, 
    249.55, 250.15, 249.75, 249.25, 249.55, 249.15, 249.25, 249.95, 248.25, 
    248.45, 249.65, 249.85, 249.15, 248.25, 248.95, 248.65, 249.05, 249.65, 
    249.55, 250.35, 250.35, 249.85, 250.65, 250.75, 250.85, 251.05, 251.25, 
    251.35, 251.85, 251.85, 252.05, 252.05, 252.25, 252.25, 252.35, 252.45, 
    252.05, 252.15, 251.95, 252.45, 251.95, 251.85, 252.35, 252.05, 252.35, 
    252.55, 252.75, 252.75, 252.95, 252.85, 253.05, 252.65, 252.95, 252.75, 
    252.85, 253.05, 253.25, 253.55, 253.85, 254.15, 254.35, 253.65, 253.95, 
    254.35, 255.25, 254.85, 251.85, 251.95, 251.15, 249.75, 248.05, 245.65, 
    245.05, 243.95, 243.35, 244.05, 243.75, 243.65, 243.15, 242.95, 243.35, 
    242.95, 242.65, 242.75, 243.15, 243.15, 243.45, 243.75, 244.45, 246.25, 
    246.35, 246.35, 246.45, 246.65, 247.55, 248.15, 248.75, 248.05, 247.85, 
    247.55, 248.55, 248.35, 248.45, 246.25, 245.45, 244.65, 245.05, 244.85, 
    244.75, 244.85, 245.05, 244.35, 244.35, 244.05, 243.45, 242.95, 243.45, 
    244.15, 244.15, 244.65, 245.65, 245.85, 246.35, 246.85, 246.65, 246.95, 
    248.05, 248.05, 247.45, 246.95, 246.25, 246.05, 246.25, 246.85, 247.35, 
    246.95, 246.85, 246.85, 246.75, 246.55, 246.45, 246.25, 245.55, 245.75, 
    245.65, 245.95, 246.45, 246.45, 247.15, 247.45, 246.95, 246.65, 246.95, 
    246.95, 246.55, 246.55, 247.05, 246.55, 246.85, 246.65, 246.05, 246.95, 
    246.15, 246.95, 246.95, 247.65, 247.05, 247.15, 248.95, 247.35, 247.15, 
    246.85, 246.45, 246.45, 246.75, 246.05, 245.55, 245.65, 245.35, 244.95, 
    244.25, 244.45, 245.55, 247.05, 247.65, 249.75, 249.65, 250.05, 251.95, 
    252.55, 255.25, 255.05, 254.15, 251.75, 252.15, 252.75, 253.25, 253.85, 
    254.15, 254.85, 255.25, 255.55, 255.75, 254.95, 254.65, 253.85, 253.35, 
    253.25, 253.15, 253.05, 252.75, 252.75, 252.45, 251.65, 251.85, 251.65, 
    251.35, 251.15, 250.75, 250.95, 251.15, 251.05, 250.75, 250.65, 249.75, 
    249.95, 250.25, 250.75, 250.85, 250.85, 250.95, 250.65, 250.35, 249.15, 
    249.75, 249.45, 250.45, 249.65, 249.45, 249.15, 249.05, 248.85, 249.75, 
    248.95, 248.75, 249.25, 251.25, 250.25, 248.55, 249.05, 250.85, 249.35, 
    250.95, 248.45, 248.55, 247.05, 246.85, 247.05, 245.85, 245.15, 246.25, 
    246.35, 246.45, 246.45, 246.45, 247.55, 247.75, 248.35, 248.65, 248.65, 
    248.55, 246.25, 245.45, 246.15, 245.85, 246.25, 246.15, 246.45, 246.45, 
    246.85, 247.35, 248.35, 246.95, 249.15, 247.45, 248.65, 247.85, 247.75, 
    249.35, 248.85, 248.65, 248.95, 249.65, 250.25, 250.65, 251.75, 252.65, 
    254.35, 254.65, 254.25, 252.05, 251.15, 251.05, 251.25, 251.15, 250.85, 
    250.45, 250.45, 250.05, 250.05, 250.05, 250.15, 250.55, 250.75, 250.65, 
    250.05, 249.25, 247.75, 247.25, 247.55, 247.65, 247.05, 246.55, 246.55, 
    246.15, 244.75, 244.95, 244.75, 245.55, 245.95, 246.55, 247.55, 248.85, 
    248.15, 248.65, 249.45, 250.45, 251.05, 250.65, 249.85, 249.85, 250.65, 
    251.65, 251.95, 252.45, 252.55, 252.45, 252.55, 252.65, 252.75, 252.95, 
    253.85, 254.15, 253.75, 253.95, 254.15, 253.65, 253.65, 253.35, 253.85, 
    252.85, 252.85, 252.05, 251.45, 250.65, 250.45, 252.55, 251.35, 251.85, 
    251.95, 251.95, 253.25, 253.25, 253.35, 254.25, 254.05, 254.55, 255.05, 
    255.55, 255.15, 255.25, 255.55, 255.75, 256.15, 256.85, 257.15, 257.45, 
    258.15, 259.85, 260.65, 261.25, 262.75, 264.25, 263.65, 264.15, 264.45, 
    265.15, 265.05, 264.85, 264.65, 265.25, 263.95, 263.85, 264.45, 264.35, 
    263.55, 262.85, 262.75, 262.75, 263.35, 264.55, 265.15, 264.35, 265.15, 
    264.95, 265.25, 265.35, 265.65, 265.05, 264.45, 264.75, 264.95, 264.75, 
    264.05, 263.95, 263.55, 262.45, 263.85, 261.35, 260.25, 261.25, 260.75, 
    260.05, 259.15, 259.05, 257.85, 257.65, 257.15, 257.45, 257.65, 257.35, 
    258.45, 258.15, 256.95, 256.35, 256.35, 257.15, 256.55, 255.85, 255.15, 
    255.05, 254.25, 254.65, 254.85, 255.65, 255.65, 256.85, 257.65, 257.45, 
    257.65, 256.95, 257.35, 256.65, 257.45, 257.45, 257.55, 257.35, 256.85, 
    257.85, 259.75, 259.65, 260.05, 260.55, 260.15, 260.25, 259.75, 259.95, 
    258.65, 260.45, 258.45, 261.65, 260.85, 261.15, 261.15, 260.75, 260.15, 
    259.45, 258.25, 258.75, 259.05, 258.85, 258.75, 258.25, 259.05, 258.65, 
    258.75, 258.75, 260.15, 259.75, 258.65, 258.75, 258.75, 258.55, 258.95, 
    258.05, 258.75, 258.95, 260.05, 257.45, 260.65, 259.25, 260.35, 260.35, 
    259.55, 261.05, 261.75, 261.55, 261.35, 261.85, 263.15, 264.75, 264.65, 
    264.55, 264.45, 264.55, 265.25, 264.55, 262.75, 261.75, 261.75, 261.65, 
    261.45, 260.65, 260.45, 259.45, 259.25, 259.25, 259.05, 258.85, 258.25, 
    257.45, 256.85, 256.85, 256.95, 256.95, 256.55, 256.25, 255.15, 254.65, 
    254.65, 254.65, 254.75, 254.45, 254.35, 254.05, 253.45, 253.15, 252.95, 
    252.45, 252.25, 252.15, 251.45, 250.65, 250.55, 250.55, 249.95, 249.25, 
    249.75, 249.85, 250.05, 250.35, 249.85, 249.95, 250.25, 250.15, 249.65, 
    253.05, 253.25, 252.85, 249.45, 248.95, 248.45, 248.55, 248.25, 248.25, 
    250.25, 250.55, 254.15, 249.15, 248.55, 250.45, 248.85, 250.25, 250.95, 
    251.85, 254.95, 256.15, 254.75, 254.85, 254.95, 254.95, 256.45, 257.35, 
    257.85, 258.05, 257.65, 257.75, 257.25, 256.35, 256.05, 255.65, 256.05, 
    254.35, 254.15, 254.55, 255.45, 255.35, 255.25, 255.25, 255.15, 255.15, 
    255.35, 254.75, 254.65, 254.45, 256.15, 255.95, 256.45, 256.95, 257.35, 
    259.65, 260.05, 262.55, 263.55, 263.35, 263.05, 262.55, 262.25, 262.65, 
    263.65, 262.75, 263.45, 263.25, 264.05, 263.95, 263.55, 263.65, 263.65, 
    263.65, 263.75, 263.55, 263.25, 262.95, 262.65, 262.55, 262.65, 262.55, 
    262.45, 262.35, 262.05, 262.05, 262.45, 261.95, 261.45, 261.35, 260.45, 
    260.25, 260.75, 260.75, 260.45, 259.95, 260.55, 260.25, 259.75, 259.35, 
    259.15, 258.95, 258.25, 257.85, 257.45, 257.25, 256.65, 256.65, 257.05, 
    256.95, 257.65, 258.85, 257.85, 258.05, 258.35, 257.65, 259.05, 259.25, 
    259.15, 260.45, 260.75, 260.55, 260.45, 260.25, 260.15, 259.85, 260.35, 
    260.55, 260.95, 260.95, 261.05, 261.95, 262.25, 262.35, 262.45, 262.35, 
    261.85, 261.65, 261.45, 261.75, 262.75, 263.15, 263.05, 262.45, 262.05, 
    261.75, 261.85, 261.65, 260.35, 260.45, 260.55, 260.95, 260.95, 261.25, 
    262.55, 261.55, 260.95, 261.05, 261.35, 260.95, 259.85, 260.65, 261.15, 
    261.25, 261.55, 261.65, 261.45, 261.95, 262.55, 263.15, 263.85, 264.45, 
    264.65, 264.35, 264.65, 265.05, 264.75, 264.55, 263.85, 263.45, 263.25, 
    263.45, 263.95, 263.85, 263.75, 264.15, 265.55, 266.55, 266.75, 266.05, 
    266.65, 266.85, 267.25, 267.35, 267.75, 266.15, 265.35, 264.85, 264.25, 
    265.45, 265.95, 265.35, 264.65, 263.85, 263.25, 262.65, 261.95, 260.75, 
    260.25, 259.45, 261.95, 263.55, 264.15, 264.75, 266.75, 267.65, 267.65, 
    267.55, 267.55, 266.75, 264.05, 263.05, 263.05, 263.15, 263.15, 262.65, 
    263.15, 263.45, 262.65, 262.55, 262.35, 261.25, 261.85, 262.55, 261.95, 
    261.95, 262.35, 262.95, 262.65, 262.85, 263.75, 263.95, 263.65, 263.95, 
    263.75, 263.45, 263.45, 263.25, 263.15, 262.85, 263.15, 261.55, 260.45, 
    259.85, 262.15, 262.05, 262.65, 262.55, 262.95, 262.85, 263.95, 264.25, 
    263.65, 263.35, 263.95, 264.25, 264.45, 264.05, 263.65, 263.05, 262.15, 
    262.25, 261.45, 258.85, 258.65, 256.15, 254.15, 254.25, 253.55, 253.05, 
    253.05, 253.05, 253.25, 253.35, 253.15, 254.15, 255.05, 255.85, 255.65, 
    255.85, 255.45, 255.05, 254.55, 254.05, 253.65, 253.45, 253.25, 253.05, 
    252.65, 252.05, 251.35, 250.95, 250.35, 250.05, 249.45, 249.35, 249.35, 
    250.05, 250.25, 250.55, 250.85, 251.55, 251.85, 251.95, 251.75, 251.65, 
    251.35, 251.15, 251.05, 250.55, 249.95, 250.25, 251.05, 250.95, 250.25, 
    250.15, 250.55, 250.75, 250.15, 250.55, 250.45, 250.65, 250.65, 250.35, 
    249.45, 248.35, 248.35, 248.25, 248.65, 248.75, 248.45, 248.35, 248.35, 
    248.25, 248.25, 248.15, 248.15, 248.15, 248.05, 247.85, 247.65, 247.45, 
    247.35, 247.45, 247.45, 247.25, 247.15, 247.05, 247.25, 247.65, 248.35, 
    248.85, 249.05, 248.95, 248.85, 248.75, 248.45, 248.45, 248.15, 248.15, 
    248.05, 248.35, 248.05, 247.85, 247.85, 247.95, 248.65, 249.05, 249.15, 
    249.25, 249.45, 249.65, 249.95, 250.45, 250.55, 251.15, 251.55, 251.75, 
    251.95, 252.15, 252.05, 251.75, 251.45, 251.15, 250.85, 250.85, 251.05, 
    251.15, 251.25, 251.45, 251.45, 251.75, 251.95, 252.35, 252.65, 252.95, 
    253.05, 253.55, 254.15, 254.85, 255.65, 255.95, 256.25, 256.15, 255.65, 
    254.85, 253.85, 254.05, 253.05, 252.65, 252.25, 252.25, 251.45, 251.35, 
    251.05, 250.95, 251.05, 251.05, 250.55, 250.65, 250.75, 251.15, 251.85, 
    251.95, 252.05, 251.85, 251.65, 251.55, 251.45, 251.25, 250.15, 250.05, 
    249.75, 249.65, 250.85, 250.55, 250.05, 250.35, 251.15, 250.65, 251.85, 
    253.25, 255.15, 255.25, 255.85, 256.25, 257.15, 257.35, 257.35, 257.45, 
    257.65, 257.25, 257.35, 257.75, 257.45, 257.55, 257.45, 257.35, 256.85, 
    256.85, 256.85, 256.35, 256.45, 257.15, 257.05, 257.45, 258.35, 257.65, 
    257.85, 259.05, 258.75, 259.95, 259.65, 259.55, 259.45, 260.05, 260.05, 
    260.05, 259.95, 259.05, 258.75, 258.35, 258.65, 258.95, 258.55, 258.25, 
    257.75, 258.85, 258.75, 258.35, 260.15, 259.85, 259.95, 260.45, 259.55, 
    259.85, 259.45, 259.35, 259.05, 257.95, 256.95, 255.35, 255.75, 254.35, 
    253.65, 253.45, 252.85, 254.15, 254.35, 254.95, 254.25, 254.95, 253.95, 
    254.55, 254.95, 255.85, 257.35, 258.15, 258.55, 259.65, 258.95, 259.05, 
    259.75, 261.25, 259.95, 257.95, 256.35, 255.65, 254.65, 253.65, 252.05, 
    251.75, 251.55, 250.95, 251.55, 251.65, 251.35, 252.05, 252.05, 253.35, 
    253.85, 254.15, 254.55, 254.65, 254.75, 254.45, 254.15, 253.75, 253.25, 
    252.75, 251.85, 251.25, 250.85, 251.75, 251.45, 250.65, 250.55, 250.05, 
    250.45, 250.85, 250.95, 251.45, 251.45, 251.75, 251.85, 252.05, 252.05, 
    251.75, 251.95, 251.95, 251.75, 252.05, 251.75, 251.45, 251.15, 250.85, 
    250.35, 249.75, 249.15, 248.85, 249.75, 249.45, 249.65, 250.35, 250.25, 
    250.15, 250.15, 251.25, 251.95, 252.25, 252.65, 252.55, 252.85, 253.55, 
    253.85, 253.55, 253.45, 252.95, 252.75, 252.65, 251.55, 250.95, 250.85, 
    250.75, 250.25, 249.65, 249.15, 249.65, 249.75, 250.15, 250.55, 250.95, 
    251.65, 252.35, 252.75, 253.35, 253.55, 253.65, 253.75, 253.65, 253.75, 
    253.55, 253.75, 253.05, 252.85, 252.65, 252.45, 254.25, 254.45, 255.85, 
    256.45, 256.05, 255.75, 255.25, 255.45, 254.85, 255.35, 256.35, 257.15, 
    258.25, 260.55, 259.55, 259.35, 258.45, 258.75, 257.95, 257.55, 257.15, 
    256.75, 255.55, 255.95, 255.65, 257.55, 257.15, 256.45, 257.95, 257.45, 
    257.55, 258.35, 258.85, 259.85, 260.15, 261.15, 261.25, 261.65, 261.65, 
    261.65, 261.65, 261.65, 262.05, 261.65, 261.55, 261.35, 261.25, 261.75, 
    263.25, 264.15, 263.55, 264.35, 265.25, 265.85, 266.65, 267.05, 267.65, 
    267.95, 268.45, 268.85, 269.05, 269.35, 269.55, 269.65, 269.65, 269.75, 
    269.55, 269.65, 269.65, 269.75, 269.85, 270.15, 270.35, 270.65, 271.05, 
    271.45, 271.65, 271.65, 271.75, 271.95, 272.05, 272.25, 272.35, 272.35, 
    272.55, 272.95, 273.25, 273.35, 273.25, 273.25, 273.05, 272.95, 272.95, 
    273.05, 273.05, 272.95, 272.75, 272.85, 272.55, 272.15, 272.05, 272.25, 
    272.45, 272.65, 272.65, 272.85, 272.75, 272.95, 272.95, 272.95, 272.95, 
    272.95, 272.95, 273.05, 272.95, 272.95, 272.85, 272.85, 272.85, 272.85, 
    272.85, 272.75, 272.65, 272.55, 272.55, 272.65, 272.75, 272.75, 272.65, 
    272.65, 272.85, 272.85, 272.95, 273.05, 273.15, 273.05, 273.05, 272.95, 
    272.95, 272.95, 272.85, 273.05, 272.95, 272.85, 272.75, 272.45, 272.55, 
    272.75, 272.65, 272.65, 272.55, 272.75, 272.55, 272.55, 272.75, 272.75, 
    272.75, 272.55, 272.55, 272.35, 272.35, 272.35, 272.35, 272.25, 272.25, 
    271.95, 271.75, 272.05, 272.15, 272.15, 271.85, 271.15, 270.75, 270.85, 
    270.65, 270.85, 270.95, 271.25, 271.15, 271.55, 271.75, 272.05, 271.65, 
    271.45, 271.45, 271.15, 270.85, 270.75, 270.55, 270.55, 270.35, 270.35, 
    270.05, 270.05, 269.85, 269.75, 269.85, 269.65, 269.95, 269.35, 269.35, 
    268.45, 269.15, 270.15, 269.65, 269.75, 270.35, 270.05, 269.05, 268.85, 
    268.25, 268.55, 268.75, 268.85, 268.85, 269.15, 269.55, 269.85, 270.35, 
    270.75, 270.95, 271.35, 271.45, 271.55, 271.55, 271.25, 271.35, 271.35, 
    271.45, 270.65, 270.65, 270.85, 270.45, 270.15, 269.75, 269.85, 269.85, 
    270.15, 270.25, 269.25, 268.75, 269.15, 268.75, 268.45, 268.55, 268.25, 
    269.05, 269.05, 269.05, 269.35, 269.65, 269.45, 270.25, 271.65, 271.35, 
    270.95, 269.95, 269.85, 270.25, 269.55, 269.05, 268.65, 268.05, 269.05, 
    267.95, 267.95, 267.15, 267.15, 267.05, 268.25, 269.05, 269.35, 269.55, 
    269.75, 269.55, 270.35, 269.45, 269.65, 269.35, 268.95, 268.85, 268.65, 
    268.35, 268.35, 268.35, 267.95, 267.85, 267.65, 268.15, 267.55, 266.85, 
    267.05, 267.15, 267.45, 267.55, 267.15, 267.05, 267.15, 267.75, 267.55, 
    267.45, 266.95, 266.45, 266.35, 266.35, 266.35, 266.05, 265.55, 265.25, 
    265.45, 265.65, 265.75, 265.65, 265.75, 265.75, 265.85, 265.85, 265.95, 
    266.05, 266.35, 266.35, 266.45, 266.45, 266.45, 266.45, 266.75, 266.85, 
    266.85, 266.95, 267.05, 267.15, 267.15, 267.15, 267.25, 267.35, 267.55, 
    267.95, 268.35, 268.45, 268.55, 268.55, 268.75, 269.05, 268.85, 268.55, 
    267.85, 267.65, 267.25, 266.65, 265.95, 265.65, 265.65, 265.85, 265.65, 
    265.25, 264.85, 265.45, 266.05, 266.05, 265.65, 265.55, 265.65, 265.45, 
    265.65, 265.75, 265.75, 265.95, 265.95, 265.75, 265.95, 265.05, 264.45, 
    264.65, 264.75, 264.75, 264.75, 264.15, 263.65, 263.15, 263.15, 262.75, 
    262.35, 261.95, 261.55, 261.25, 261.25, 261.55, 261.15, 260.75, 261.35, 
    261.75, 261.25, 261.45, 261.75, 262.25, 262.85, 263.75, 264.05, 264.15, 
    264.15, 264.95, 264.65, 264.15, 264.15, 264.15, 263.15, 263.95, 263.55, 
    263.55, 261.85, 263.35, 263.55, 264.25, 264.85, 265.75, 265.15, 265.15, 
    267.15, 267.15, 268.05, 268.45, 268.15, 268.25, 268.55, 268.55, 268.45, 
    268.45, 268.45, 268.95, 269.25, 269.35, 269.35, 269.35, 269.35, 269.05, 
    269.05, 268.95, 268.45, 268.55, 268.75, 268.85, 268.85, 269.05, 269.25, 
    269.45, 269.85, 269.25, 268.85, 269.45, 268.65, 267.85, 267.85, 267.45, 
    267.15, 267.25, 267.15, 266.85, 266.05, 266.05, 266.35, 266.75, 266.35, 
    266.45, 266.35, 266.75, 266.95, 266.95, 267.55, 267.75, 268.05, 267.75, 
    267.35, 267.35, 266.95, 266.45, 265.85, 266.35, 265.05, 265.35, 265.05, 
    266.95, 267.35, 267.55, 267.35, 267.75, 267.95, 268.15, 268.25, 267.85, 
    267.95, 268.85, 269.25, 269.35, 269.85, 269.55, 269.85, 270.35, 270.85, 
    271.05, 271.35, 271.05, 270.85, 270.45, 271.65, 271.45, 270.55, 269.25, 
    269.65, 269.35, 269.95, 269.85, 270.35, 270.35, 270.55, 270.35, 270.95, 
    271.15, 271.15, 271.25, 271.35, 271.65, 271.15, 270.95, 270.35, 270.25, 
    270.35, 270.05, 269.55, 269.65, 269.95, 269.85, 269.55, 269.35, 269.55, 
    269.35, 269.25, 269.15, 269.05, 268.55, 268.55, 268.25, 268.55, 268.15, 
    268.05, 267.65, 267.45, 267.45, 267.65, 267.45, 267.55, 267.75, 267.75, 
    267.75, 268.05, 267.85, 267.95, 267.95, 267.95, 268.15, 267.85, 267.95, 
    267.65, 267.55, 267.25, 266.65, 266.35, 266.15, 266.25, 266.35, 266.35, 
    266.65, 266.55, 265.95, 265.85, 265.65, 265.35, 265.25, 265.05, 264.55, 
    264.55, 264.75, 265.05, 265.35, 265.55, 265.95, 266.95, 266.55, 267.15, 
    266.65, 266.85, 267.25, 266.85, 267.75, 266.55, 266.25, 265.85, 265.75, 
    265.55, 265.25, 264.85, 264.75, 265.05, 265.55, 265.95, 265.95, 266.25, 
    266.75, 266.15, 266.25, 266.25, 266.15, 266.05, 266.35, 266.65, 266.45, 
    266.15, 266.25, 265.75, 265.45, 265.25, 265.05, 265.55, 265.15, 265.05, 
    265.15, 265.45, 265.25, 264.95, 264.65, 265.05, 265.45, 265.85, 265.65, 
    265.95, 265.95, 265.95, 266.25, 266.35, 266.85, 266.85, 266.65, 266.05, 
    266.05, 265.95, 265.95, 266.05, 266.05, 266.15, 266.25, 266.45, 266.35, 
    266.35, 266.55, 266.75, 266.95, 268.05, 268.55, 269.35, 270.35, 270.75, 
    270.85, 270.95, 270.95, 270.85, 270.75, 270.65, 270.35, 270.25, 270.15, 
    270.15, 270.15, 269.95, 270.15, 269.95, 270.05, 270.35, 270.55, 270.75, 
    270.85, 271.15, 271.75, 271.85, 272.25, 272.05, 272.45, 272.15, 272.25, 
    272.55, 272.75, 273.25, 272.25, 272.15, 271.95, 271.65, 271.75, 271.65, 
    271.55, 271.15, 271.25, 271.25, 271.15, 270.75, 270.35, 270.25, 270.25, 
    270.15, 270.35, 270.35, 270.45, 270.35, 270.45, 270.55, 270.25, 270.25, 
    270.25, 270.25, 269.85, 269.55, 269.65, 269.55, 270.05, 270.25, 270.45, 
    270.75, 270.75, 271.35, 271.55, 271.85, 271.45, 272.15, 272.25, 272.25, 
    272.45, 272.45, 272.65, 272.55, 272.45, 272.25, 272.25, 272.05, 271.85, 
    271.75, 271.75, 271.85, 271.85, 271.75, 271.85, 272.15, 272.75, 271.25, 
    270.05, 269.35, 268.15, 267.65, 267.15, 267.15, 266.85, 266.85, 266.95, 
    266.95, 266.95, 266.85, 266.45, 267.15, 265.85, 265.85, 267.05, 267.45, 
    266.85, 266.55, 266.25, 265.95, 265.65, 265.65, 265.45, 265.85, 266.55, 
    266.35, 266.45, 266.25, 266.45, 265.65, 265.15, 265.25, 265.65, 266.05, 
    266.15, 266.35, 266.45, 266.35, 266.25, 266.35, 266.05, 266.35, 266.35, 
    266.95, 266.85, 266.75, 266.95, 266.85, 266.75, 266.75, 266.75, 266.75, 
    266.85, 266.85, 266.85, 267.05, 267.45, 267.85, 268.25, 268.75, 269.05, 
    269.45, 269.85, 270.15, 270.35, 270.55, 270.75, 270.95, 271.15, 271.15, 
    271.35, 271.75, 271.95, 271.95, 271.95, 272.05, 272.45, 272.25, 272.35, 
    272.25, 272.25, 272.15, 272.25, 272.25, 271.65, 271.65, 271.45, 271.25, 
    271.15, 270.35, 268.85, 267.55, 267.25, 266.75, 266.75, 266.45, 265.75, 
    265.65, 265.75, 265.75, 265.55, 265.25, 265.05, 265.05, 265.15, 265.15, 
    265.25, 265.85, 266.25, 266.75, 267.25, 267.25, 267.35, 267.25, 267.65, 
    267.95, 268.05, 268.15, 268.25, 268.25, 268.35, 268.25, 268.15, 268.35, 
    268.75, 268.55, 268.35, 268.35, 268.25, 267.95, 268.15, 268.25, 267.95, 
    267.85, 268.55, 268.55, 268.65, 268.85, 269.05, 269.55, 269.55, 269.65, 
    269.25, 269.65, 269.85, 269.85, 270.15, 270.35, 270.45, 270.75, 270.75, 
    270.55, 270.45, 270.45, 270.45, 270.05, 269.85, 269.65, 269.95, 269.15, 
    269.25, 269.05, 268.35, 269.05, 268.55, 268.55, 269.15, 269.15, 269.05, 
    269.15, 269.35, 269.85, 270.05, 270.35, 270.55, 270.65, 270.85, 271.05, 
    271.05, 271.15, 271.05, 271.05, 271.05, 270.95, 270.95, 270.75, 270.05, 
    269.75, 269.65, 269.95, 270.05, 270.35, 271.25, 271.45, 272.25, 272.95, 
    272.95, 272.85, 272.65, 272.85, 272.35, 271.95, 272.25, 272.55, 272.45, 
    272.65, 272.85, 273.35, 271.65, 272.05, 272.45, 271.85, 272.75, 273.45, 
    272.75, 272.45, 272.15, 272.35, 273.55, 273.05, 272.55, 272.65, 272.55, 
    272.55, 272.75, 272.75, 272.95, 272.85, 272.85, 272.85, 272.95, 272.25, 
    272.15, 272.05, 271.95, 271.95, 271.85, 272.05, 272.15, 272.55, 274.45, 
    273.75, 273.35, 273.65, 273.55, 272.85, 272.85, 272.55, 272.85, 272.25, 
    272.15, 271.95, 271.85, 271.95, 272.05, 272.25, 272.75, 272.85, 272.85, 
    272.95, 272.45, 272.25, 272.25, 272.25, 271.95, 271.95, 272.05, 272.15, 
    271.75, 271.95, 271.85, 271.75, 271.65, 272.15, 272.45, 272.25, 271.65, 
    271.65, 271.65, 271.75, 271.45, 271.55, 271.55, 271.75, 271.55, 271.45, 
    271.55, 271.65, 271.75, 271.75, 271.95, 272.05, 272.15, 272.25, 272.35, 
    272.55, 272.45, 272.45, 272.55, 272.45, 272.45, 272.35, 272.25, 272.25, 
    272.25, 272.05, 271.95, 271.65, 271.45, 271.65, 271.35, 271.75, 272.45, 
    272.05, 272.45, 272.65, 273.05, 273.45, 273.75, 273.55, 273.75, 273.75, 
    273.75, 273.65, 273.65, 273.65, 273.75, 273.75, 273.85, 273.85, 273.95, 
    274.25, 274.25, 274.15, 273.95, 273.65, 273.55, 273.55, 273.75, 274.15, 
    274.45, 274.35, 274.65, 274.85, 274.55, 274.25, 274.05, 273.95, 273.95, 
    273.85, 273.75, 273.05, 273.65, 272.35, 272.15, 273.05, 274.85, 273.05, 
    274.05, 274.35, 274.15, 274.45, 274.75, 274.85, 274.85, 275.45, 275.55, 
    275.65, 275.85, 276.05, 276.35, 276.45, 275.55, 274.65, 274.95, 274.85, 
    274.75, 274.15, 274.05, 273.95, 273.55, 273.55, 273.85, 274.15, 274.65, 
    273.35, 273.45, 275.25, 275.95, 275.15, 274.85, 273.15, 274.45, 273.25, 
    271.45, 273.15, 273.95, 273.45, 272.85, 272.45, 272.85, 272.55, 276.35, 
    276.15, 275.75, 274.75, 274.15, 273.75, 273.45, 273.95, 273.25, 272.25, 
    271.05, 271.15, 270.25, 270.05, 269.95, 270.05, 270.25, 270.65, 270.45, 
    270.55, 270.55, 270.55, 271.05, 271.25, 271.55, 271.65, 271.85, 272.05, 
    272.05, 272.05, 272.05, 271.75, 271.75, 271.35, 271.55, 271.65, 271.95, 
    272.55, 273.25, 272.75, 272.75, 272.65, 272.55, 272.25, 272.15, 272.25, 
    272.45, 272.25, 272.45, 272.35, 272.45, 272.75, 272.55, 272.75, 272.75, 
    272.85, 272.65, 272.75, 273.05, 272.25, 272.25, 272.05, 270.55, 269.85, 
    269.35, 269.25, 268.75, 268.35, 268.15, 268.25, 268.75, 269.15, 269.25, 
    269.85, 270.55, 270.95, 271.15, 271.55, 271.55, 271.55, 271.75, 271.65, 
    271.35, 271.35, 271.85, 272.25, 272.25, 271.85, 272.05, 272.25, 272.05, 
    272.05, 271.95, 271.95, 271.75, 271.65, 271.65, 271.55, 271.45, 271.35, 
    271.45, 270.55, 269.65, 269.95, 269.85, 269.75, 270.05, 270.35, 270.45, 
    271.15, 271.55, 272.25, 272.45, 272.55, 272.55, 272.45, 272.25, 271.65, 
    270.95, 270.85, 270.65, 270.35, 269.95, 269.35, 269.35, 269.25, 269.85, 
    270.05, 269.95, 270.25, 270.55, 270.55, 270.75, 270.75, 270.75, 270.75, 
    271.05, 270.85, 270.45, 270.55, 270.95, 270.75, 271.05, 271.15, 271.15, 
    271.25, 271.25, 270.95, 270.85, 270.65, 270.55, 270.55, 270.85, 271.15, 
    271.15, 271.55, 271.05, 271.05, 270.85, 271.05, 271.55, 271.45, 271.45, 
    270.75, 270.75, 270.35, 270.65, 271.15, 271.25, 270.55, 270.15, 270.35, 
    270.25, 270.35, 270.95, 271.15, 271.15, 271.35, 271.85, 271.15, 271.45, 
    271.55, 271.15, 271.25, 271.45, 271.05, 271.15, 270.85, 270.85, 270.85, 
    270.85, 270.45, 270.65, 270.45, 270.65, 270.55, 270.35, 270.65, 270.75, 
    270.95, 270.85, 270.85, 271.15, 270.85, 270.95, 270.05, 270.85, 270.85, 
    270.55, 270.35, 270.35, 270.65, 270.45, 270.35, 270.15, 270.05, 269.75, 
    269.75, 269.85, 269.65, 269.65, 269.85, 270.15, 270.25, 270.35, 270.45, 
    270.45, 270.45, 270.95, 270.35, 270.35, 270.25, 270.65, 270.95, 270.55, 
    270.25, 270.45, 270.35, 270.55, 270.65, 271.05, 271.25, 271.65, 272.25, 
    272.45, 272.75, 273.15, 273.45, 273.25, 273.25, 273.65, 273.65, 273.25, 
    273.35, 273.35, 273.55, 273.15, 272.95, 273.25, 272.65, 273.15, 273.25, 
    272.65, 272.75, 272.75, 272.65, 272.55, 272.45, 272.65, 272.35, 272.55, 
    272.65, 272.75, 273.35, 272.95, 273.75, 273.15, 273.95, 273.85, 273.75, 
    274.25, 274.55, 274.75, 274.45, 274.25, 275.15, 275.65, 275.45, 275.75, 
    274.55, 274.45, 274.35, 273.45, 274.65, 274.95, 273.75, 273.85, 274.35, 
    274.65, 274.15, 274.05, 274.05, 274.85, 274.45, 274.15, 273.95, 272.65, 
    274.75, 274.45, 275.15, 275.45, 275.85, 274.75, 274.85, 275.55, 274.75, 
    274.45, 274.65, 274.65, 274.75, 274.85, 274.75, 274.85, 274.65, 274.75, 
    274.95, 274.35, 274.05, 274.05, 274.25, 273.95, 273.95, 274.05, 274.35, 
    274.55, 274.75, 274.55, 274.45, 274.85, 275.35, 275.25, 274.85, 273.85, 
    277.15, 277.05, 277.25, 277.45, 277.25, 277.15, 277.55, 277.15, 277.05, 
    276.55, 275.25, 275.95, 274.65, 274.15, 274.15, 274.85, 274.75, 274.95, 
    274.65, 274.15, 274.45, 274.45, 274.85, 275.75, 276.45, 276.65, 275.65, 
    274.95, 274.75, 276.05, 276.55, 276.35, 275.95, 276.35, 276.25, 276.05, 
    276.25, 275.65, 276.15, 276.45, 275.55, 275.25, 274.75, 274.65, 274.85, 
    275.85, 275.95, 276.05, 277.25, 278.55, 278.25, 277.25, 275.95, 273.95, 
    273.75, 273.55, 273.65, 274.05, 274.15, 275.55, 276.25, 276.05, 274.25, 
    274.15, 273.95, 273.95, 273.55, 273.25, 273.55, 272.85, 272.65, 272.85, 
    272.95, 273.05, 272.85, 272.95, 272.65, 272.45, 272.45, 272.55, 272.55, 
    272.55, 272.55, 272.45, 272.45, 272.45, 272.45, 272.45, 272.45, 272.45, 
    272.55, 272.85, 274.15, 274.85, 273.35, 273.55, 275.25, 274.65, 275.55, 
    276.05, 275.65, 275.25, 276.45, 275.85, 275.85, 275.35, 275.15, 272.25, 
    272.35, 272.65, 272.65, 272.35, 272.05, 272.65, 272.95, 272.65, 273.25, 
    273.15, 273.25, 273.45, 273.45, 273.55, 273.85, 273.75, 273.75, 273.75, 
    273.75, 273.35, 273.35, 273.35, 273.45, 273.35, 273.15, 272.95, 272.75, 
    272.65, 272.45, 272.65, 273.05, 275.75, 274.25, 275.05, 274.45, 275.65, 
    277.05, 277.35, 278.35, 277.05, 277.45, 276.75, 276.45, 276.25, 276.35, 
    276.25, 275.95, 275.95, 276.75, 276.95, 279.45, 280.05, 279.05, 277.35, 
    277.65, 276.55, 276.55, 276.35, 275.85, 275.65, 276.35, 276.45, 276.35, 
    276.25, 276.25, 276.35, 277.15, 276.55, 275.35, 275.05, 275.25, 275.35, 
    275.45, 276.15, 277.85, 277.85, 277.45, 277.35, 275.05, 275.25, 275.75, 
    275.85, 275.35, 275.65, 275.45, 275.35, 276.85, 276.45, 275.15, 274.65, 
    274.05, 274.15, 274.35, 275.25, 274.55, 274.05, 274.85, 273.95, 274.05, 
    274.25, 275.25, 275.75, 275.65, 276.95, 274.85, 275.05, 274.95, 275.75, 
    275.25, 275.55, 275.85, 275.75, 276.05, 276.05, 275.95, 276.45, 276.15, 
    277.05, 275.75, 275.25, 275.05, 275.65, 276.15, 276.05, 275.95, 275.85, 
    275.65, 275.45, 274.95, 275.95, 275.75, 276.35, 276.45, 275.75, 277.05, 
    277.25, 277.55, 278.05, 278.05, 277.75, 278.05, 277.15, 277.05, 276.55, 
    276.25, 275.85, 275.35, 275.05, 275.35, 275.35, 275.75, 275.85, 277.05, 
    277.65, 278.55, 278.25, 274.65, 275.05, 275.05, 275.55, 276.45, 277.45, 
    276.05, 275.05, 274.85, 273.65, 273.15, 275.55, 274.75, 275.15, 275.85, 
    275.65, 275.35, 275.05, 276.95, 276.75, 277.45, 277.35, 276.85, 276.75, 
    277.25, 277.25, 277.05, 277.05, 277.75, 277.15, 277.85, 277.35, 277.35, 
    277.45, 278.25, 278.45, 277.95, 278.55, 277.75, 277.05, 276.75, 276.35, 
    275.95, 275.95, 277.05, 275.35, 275.25, 275.65, 275.45, 275.25, 274.95, 
    274.85, 275.05, 275.25, 275.35, 275.45, 275.95, 275.95, 275.75, 275.55, 
    275.65, 275.65, 275.45, 275.35, 275.45, 275.45, 275.95, 275.75, 275.95, 
    276.25, 276.15, 276.25, 276.35, 276.25, 276.35, 276.15, 276.25, 276.25, 
    276.05, 275.45, 275.65, 275.45, 275.35, 275.65, 275.85, 275.95, 276.75, 
    276.55, 276.75, 276.55, 275.95, 275.85, 275.75, 275.55, 275.85, 276.05, 
    276.75, 277.15, 278.55, 278.35, 277.45, 278.75, 276.85, 277.55, 277.35, 
    278.25, 278.25, 278.15, 280.15, 279.25, 279.55, 279.65, 276.25, 275.85, 
    276.15, 276.85, 275.95, 275.95, 275.65, 276.25, 277.05, 277.15, 277.25, 
    278.05, 278.05, 277.35, 276.95, 276.75, 276.45, 276.25, 276.55, 276.65, 
    276.95, 276.25, 276.35, 275.85, 275.55, 274.85, 274.85, 275.75, 276.85, 
    276.65, 275.75, 277.05, 277.45, 277.55, 278.15, 277.35, 277.15, 277.45, 
    277.85, 276.95, 275.55, 276.15, 276.95, 275.45, 274.45, 274.35, 274.95, 
    274.95, 274.25, 274.35, 274.95, 274.95, 275.05, 274.65, 274.25, 273.95, 
    273.85, 273.75, 273.55, 273.65, 273.55, 273.85, 273.45, 273.25, 273.15, 
    273.15, 273.25, 273.25, 273.45, 273.85, 274.25, 274.35, 274.55, 274.85, 
    274.85, 274.25, 274.85, 275.45, 275.35, 275.35, 275.65, 275.45, 275.35, 
    275.75, 276.25, 275.75, 275.85, 275.95, 276.45, 276.25, 276.45, 277.75, 
    276.65, 276.35, 275.55, 275.95, 274.55, 274.15, 274.65, 275.65, 276.95, 
    275.95, 275.75, 274.85, 275.05, 274.35, 275.75, 274.95, 274.65, 274.45, 
    274.15, 273.65, 273.65, 273.65, 273.55, 273.45, 273.35, 273.55, 273.35, 
    273.05, 273.25, 273.65, 273.65, 273.65, 273.85, 273.95, 273.65, 273.95, 
    273.35, 273.65, 273.25, 273.25, 273.15, 273.05, 272.95, 272.85, 272.65, 
    272.65, 272.95, 272.75, 272.85, 272.75, 272.65, 272.75, 272.55, 272.55, 
    273.05, 272.95, 272.55, 272.95, 273.45, 273.25, 273.85, 273.75, 273.65, 
    274.25, 273.85, 273.75, 274.15, 273.95, 273.45, 273.45, 273.05, 272.65, 
    272.45, 272.35, 272.65, 272.85, 272.45, 272.25, 272.45, 272.65, 272.85, 
    272.85, 273.45, 274.05, 273.85, 274.35, 274.15, 273.65, 273.55, 273.45, 
    273.25, 273.05, 272.95, 273.05, 272.95, 273.05, 272.95, 272.95, 272.95, 
    272.95, 272.85, 272.85, 272.85, 272.95, 272.95, 272.95, 273.15, 273.15, 
    273.35, 273.45, 273.15, 273.25, 273.25, 273.15, 273.05, 272.95, 272.95, 
    272.95, 273.05, 273.05, 273.05, 273.05, 272.95, 272.95, 272.85, 272.85, 
    272.85, 272.95, 272.95, 272.95, 272.95, 272.95, 272.95, 273.05, 273.15, 
    273.25, 273.45, 273.15, 273.25, 273.25, 273.25, 273.25, 273.25, 273.35, 
    273.25, 273.25, 273.25, 273.35, 273.35, 273.55, 273.45, 273.45, 273.55, 
    273.75, 273.85, 274.15, 274.05, 274.25, 274.45, 274.55, 275.05, 275.35, 
    275.65, 275.45, 274.85, 274.45, 274.35, 274.65, 274.75, 275.05, 275.85, 
    276.15, 275.15, 276.65, 277.75, 277.15, 278.25, 278.55, 278.85, 278.95, 
    277.75, 278.05, 278.65, 276.75, 279.35, 278.65, 278.35, 280.45, 277.35, 
    276.55, 277.05, 276.45, 276.85, 275.55, 276.05, 276.35, 275.85, 276.05, 
    276.55, 276.45, 276.15, 278.05, 278.05, 277.85, 277.85, 278.05, 278.75, 
    277.15, 277.25, 278.35, 280.25, 279.35, 278.55, 278.15, 278.35, 277.65, 
    276.65, 276.45, 276.45, 276.45, 276.25, 275.95, 275.75, 275.95, 275.75, 
    275.65, 276.35, 275.55, 275.65, 275.95, 275.55, 275.95, 275.15, 275.15, 
    275.25, 275.45, 275.55, 275.75, 275.95, 275.95, 275.75, 275.35, 275.75, 
    275.65, 275.25, 275.25, 275.65, 275.65, 275.95, 276.35, 276.25, 276.15, 
    276.15, 275.95, 275.75, 275.75, 275.95, 275.85, 276.15, 275.95, 275.95, 
    275.65, 275.25, 274.95, 274.75, 274.65, 274.55, 274.55, 274.65, 274.75, 
    274.75, 275.35, 275.65, 275.95, 275.95, 276.05, 276.25, 276.65, 276.45, 
    276.55, 276.45, 276.45, 276.45, 276.35, 276.95, 276.55, 276.55, 276.35, 
    276.25, 275.95, 275.85, 276.05, 276.05, 276.05, 276.55, 276.55, 276.25, 
    276.25, 276.35, 276.35, 276.45, 276.75, 276.55, 277.75, 277.65, 277.65, 
    277.25, 277.25, 275.85, 275.85, 276.55, 276.35, 276.15, 276.25, 275.75, 
    275.95, 275.75, 275.85, 276.25, 275.95, 275.65, 276.05, 276.65, 276.95, 
    275.65, 275.95, 276.05, 276.15, 275.95, 275.75, 275.75, 275.85, 275.55, 
    276.75, 275.85, 276.25, 275.75, 275.15, 275.35, 275.55, 275.65, 275.35, 
    275.25, 275.25, 275.65, 275.75, 275.55, 276.05, 276.45, 276.05, 275.85, 
    275.25, 275.25, 275.15, 274.95, 274.75, 274.85, 274.55, 274.35, 274.75, 
    274.85, 274.55, 274.25, 274.35, 274.25, 274.25, 274.65, 274.65, 274.55, 
    274.55, 274.75, 274.85, 275.05, 275.15, 275.05, 274.65, 274.85, 275.45, 
    276.15, 275.85, 276.25, 275.95, 276.45, 276.45, 276.45, 276.15, 276.05, 
    276.65, 276.65, 276.65, 276.45, 275.95, 276.15, 275.85, 276.35, 276.05, 
    276.05, 276.15, 275.95, 276.45, 276.25, 276.85, 276.35, 276.45, 276.65, 
    275.95, 276.15, 276.25, 276.45, 276.55, 276.55, 276.55, 276.25, 276.05, 
    276.15, 276.25, 276.15, 276.05, 275.35, 275.05, 274.95, 275.45, 276.35, 
    278.15, 277.85, 278.45, 278.45, 277.45, 277.25, 277.75, 277.95, 278.15, 
    277.85, 277.55, 277.75, 277.15, 276.65, 276.85, 276.35, 276.65, 276.65, 
    277.05, 277.25, 276.75, 276.65, 276.95, 276.35, 276.85, 276.65, 276.85, 
    275.85, 275.95, 276.05, 275.55, 275.35, 276.95, 279.25, 279.05, 278.75, 
    279.05, 279.15, 278.95, 279.05, 278.85, 278.65, 278.35, 277.95, 278.05, 
    277.25, 277.15, 277.45, 276.65, 277.15, 277.45, 277.65, 276.85, 276.75, 
    276.75, 277.65, 277.95, 278.15, 278.35, 278.15, 277.45, 277.65, 277.25, 
    276.55, 275.45, 275.55, 275.75, 276.45, 278.05, 277.75, 276.65, 276.35, 
    276.25, 276.35, 276.55, 276.85, 277.55, 278.15, 276.45, 277.95, 277.25, 
    277.15, 277.75, 277.65, 277.65, 277.95, 277.25, 277.25, 277.85, 278.05, 
    278.05, 277.15, 277.25, 277.75, 278.05, 278.05, 278.45, 279.25, 278.65, 
    277.75, 278.35, 280.25, 279.15, 277.45, 277.55, 276.85, 280.15, 277.75, 
    277.75, 278.05, 277.65, 276.85, 276.85, 277.15, 277.45, 277.25, 277.35, 
    277.25, 277.15, 277.25, 277.05, 277.35, 277.15, 276.55, 276.85, 276.45, 
    275.95, 275.95, 275.45, 275.05, 275.05, 274.95, 274.85, 274.75, 274.85, 
    274.85, 274.85, 274.85, 274.85, 274.75, 274.55, 274.45, 274.45, 274.65, 
    274.35, 274.25, 274.25, 273.95, 273.55, 273.65, 273.65, 273.15, 273.05, 
    272.95, 273.05, 272.95, 272.75, 272.95, 272.95, 273.45, 273.45, 273.45, 
    273.45, 273.35, 273.35, 273.55, 274.95, 274.45, 274.95, 274.95, 274.85, 
    274.05, 274.15, 273.45, 273.65, 273.15, 272.95, 273.15, 272.95, 272.45, 
    272.15, 271.65, 271.45, 271.65, 271.35, 271.45, 272.05, 273.25, 273.15, 
    272.95, 273.05, 273.15, 273.15, 273.65, 274.05, 273.95, 274.15, 274.15, 
    274.35, 274.25, 274.25, 273.45, 273.55, 273.25, 272.25, 271.95, 271.75, 
    272.15, 272.05, 272.05, 272.55, 273.05, 272.95, 273.15, 272.95, 272.75, 
    274.45, 274.85, 274.45, 274.75, 274.85, 275.25, 275.55, 276.05, 276.15, 
    275.75, 275.85, 276.15, 276.05, 276.15, 276.35, 276.25, 276.35, 275.85, 
    276.15, 276.75, 276.65, 277.15, 277.15, 277.25, 277.35, 277.35, 276.65, 
    276.65, 276.65, 276.95, 276.85, 276.95, 278.05, 277.65, 276.85, 276.35, 
    277.05, 276.95, 275.85, 275.15, 274.85, 274.55, 274.55, 274.55, 274.45, 
    273.75, 273.75, 273.95, 274.15, 273.65, 273.55, 273.45, 272.85, 272.55, 
    271.95, 271.75, 271.75, 271.85, 271.15, 271.05, 270.95, 271.15, 271.15, 
    271.35, 271.55, 271.75, 271.95, 272.05, 272.45, 272.05, 272.45, 272.45, 
    272.85, 272.65, 272.95, 272.65, 272.75, 273.05, 273.85, 274.05, 273.95, 
    274.05, 274.25, 274.25, 274.15, 274.35, 274.55, 274.55, 274.55, 274.65, 
    274.15, 274.25, 274.45, 274.65, 274.55, 274.65, 274.35, 274.05, 273.25, 
    273.15, 273.05, 272.55, 271.55, 271.25, 271.05, 271.35, 271.45, 271.75, 
    272.35, 272.25, 272.95, 272.35, 272.85, 273.15, 273.55, 273.75, 274.35, 
    273.85, 274.15, 273.95, 274.15, 274.65, 274.65, 274.75, 274.75, 274.65, 
    274.95, 274.95, 274.85, 274.75, 274.55, 274.65, 274.45, 274.45, 274.15, 
    273.95, 274.55, 275.25, 275.25, 275.25, 275.15, 274.45, 274.25, 274.15, 
    274.15, 274.35, 274.75, 273.65, 273.55, 274.45, 274.35, 274.35, 275.05, 
    275.45, 274.05, 273.95, 273.35, 273.05, 273.05, 273.05, 273.15, 273.45, 
    273.65, 273.75, 273.75, 274.55, 274.55, 274.65, 274.15, 274.35, 274.05, 
    274.05, 273.95, 273.95, 273.45, 272.95, 272.45, 272.15, 271.65, 271.35, 
    271.35, 271.25, 271.25, 271.55, 271.35, 271.25, 271.05, 270.85, 270.85, 
    270.95, 271.15, 271.35, 271.55, 271.45, 271.65, 271.65, 271.95, 272.15, 
    273.45, 274.95, 275.25, 274.95, 275.35, 275.65, 275.75, 275.55, 275.65, 
    275.85, 275.65, 275.65, 275.95, 275.95, 276.15, 276.75, 276.25, 275.95, 
    276.45, 276.65, 276.55, 276.55, 276.55, 276.35, 276.35, 276.05, 275.95, 
    275.85, 276.05, 275.85, 276.15, 277.25, 277.05, 276.85, 276.45, 276.25, 
    276.65, 276.55, 276.85, 277.15, 276.95, 277.15, 277.05, 276.95, 276.85, 
    277.25, 277.15, 277.15, 276.75, 276.85, 276.45, 276.25, 276.25, 276.25, 
    276.25, 276.25, 276.35, 276.25, 276.55, 276.75, 276.75, 276.95, 277.05, 
    277.35, 277.55, 277.15, 277.15, 277.35, 277.15, 278.35, 279.05, 278.55, 
    278.75, 277.25, 277.15, 276.75, 276.35, 276.15, 277.15, 277.85, 277.95, 
    278.05, 278.45, 278.65, 278.75, 278.65, 278.05, 277.65, 278.55, 277.75, 
    278.25, 278.95, 278.75, 278.35, 278.25, 278.25, 277.25, 276.45, 276.65, 
    277.05, 276.65, 277.35, 277.25, 277.85, 277.65, 277.95, 278.35, 278.45, 
    278.35, 278.45, 278.55, 278.15, 277.75, 277.85, 278.35, 278.75, 278.05, 
    278.15, 277.85, 277.35, 278.05, 277.85, 277.95, 277.75, 277.35, 277.25, 
    277.35, 277.35, 277.35, 277.45, 277.75, 277.35, 277.75, 277.35, 277.45, 
    278.25, 278.35, 277.55, 277.75, 278.05, 278.35, 277.65, 277.95, 278.05, 
    277.45, 277.05, 276.75, 277.05, 276.65, 276.25, 276.05, 277.05, 277.05, 
    277.25, 276.15, 276.05, 275.75, 276.15, 276.75, 277.05, 276.45, 276.35, 
    275.85, 275.85, 275.95, 276.75, 277.65, 278.15, 277.55, 278.25, 278.85, 
    278.15, 278.45, 277.65, 277.75, 277.05, 276.85, 276.65, 276.55, 277.85, 
    277.05, 277.45, 277.25, 277.15, 276.55, 276.75, 277.65, 276.65, 277.75, 
    278.25, 278.15, 276.65, 276.85, 278.65, 277.95, 278.05, 278.35, 278.45, 
    277.65, 278.15, 277.85, 277.85, 277.55, 276.65, 277.65, 276.75, 277.45, 
    278.25, 277.65, 277.15, 276.45, 276.55, 276.95, 277.05, 276.65, 277.05, 
    277.55, 277.75, 277.25, 276.45, 276.95, 276.85, 277.15, 277.25, 277.25, 
    277.55, 277.65, 277.15, 276.85, 276.35, 276.85, 276.65, 277.05, 277.45, 
    277.25, 277.75, 277.85, 276.85, 276.15, 275.65, 274.45, 274.75, 274.95, 
    275.05, 275.45, 275.45, 274.95, 275.15, 275.55, 275.55, 275.65, 275.75, 
    275.85, 275.65, 275.75, 275.65, 275.55, 275.55, 275.85, 276.05, 275.75, 
    276.05, 276.05, 275.85, 275.75, 276.05, 275.75, 276.05, 276.05, 276.15, 
    276.15, 276.55, 276.15, 276.35, 276.15, 276.15, 276.15, 276.75, 276.15, 
    276.05, 276.05, 276.05, 276.15, 276.65, 276.35, 276.15, 276.65, 276.35, 
    276.75, 277.05, 276.85, 277.35, 277.05, 276.95, 277.05, 276.85, 276.65, 
    276.65, 275.75, 275.65, 275.75, 275.65, 275.75, 275.75, 275.55, 275.55, 
    275.45, 275.45, 275.45, 275.35, 275.25, 275.15, 275.05, 275.05, 275.05, 
    275.05, 275.05, 275.05, 275.05, 274.75, 275.15, 275.15, 275.25, 275.55, 
    275.55, 275.75, 275.95, 275.95, 275.85, 275.75, 275.95, 275.75, 276.15, 
    275.85, 276.15, 276.35, 275.85, 275.95, 276.05, 276.35, 275.25, 276.15, 
    276.45, 276.15, 276.55, 276.45, 276.55, 276.05, 276.05, 276.35, 276.55, 
    275.65, 275.65, 275.55, 275.15, 275.15, 274.85, 274.75, 274.85, 275.05, 
    275.15, 275.25, 275.35, 275.35, 275.45, 275.55, 275.55, 275.25, 275.35, 
    275.55, 275.05, 275.05, 275.15, 274.85, 274.35, 274.15, 273.85, 273.85, 
    273.65, 273.75, 273.55, 273.15, 273.05, 273.45, 273.45, 273.55, 273.35, 
    273.35, 273.35, 273.45, 273.35, 272.95, 272.75, 272.65, 272.65, 272.75, 
    272.75, 272.75, 273.15, 273.75, 274.15, 274.25, 274.35, 274.25, 274.25, 
    274.35, 274.25, 274.25, 274.05, 273.95, 274.05, 273.85, 273.85, 273.85, 
    273.85, 273.85, 273.85, 273.85, 273.85, 273.95, 273.75, 273.55, 273.45, 
    273.85, 274.05, 274.25, 274.25, 274.25, 274.15, 273.95, 273.45, 273.65, 
    273.85, 273.65, 273.55, 273.75, 273.85, 274.25, 274.05, 274.35, 274.35, 
    274.65, 274.95, 274.95, 274.35, 274.05, 274.35, 274.25, 274.25, 274.45, 
    274.45, 274.25, 274.25, 273.85, 273.85, 273.05, 272.95, 272.65, 272.55, 
    272.45, 271.75, 271.75, 272.05, 272.85, 273.25, 273.65, 273.75, 273.35, 
    273.35, 273.85, 274.05, 274.35, 274.65, 274.85, 274.55, 274.45, 274.15, 
    274.35, 274.35, 274.95, 274.65, 274.85, 275.05, 275.25, 275.45, 275.25, 
    275.55, 275.65, 275.75, 275.75, 275.85, 275.95, 276.05, 276.55, 276.65, 
    277.35, 277.25, 277.25, 277.05, 276.55, 276.25, 275.55, 274.85, 274.75, 
    275.05, 275.45, 275.35, 274.95, 275.05, 275.25, 275.45, 275.15, 274.55, 
    274.35, 275.25, 274.65, 274.55, 274.75, 274.75, 274.55, 275.05, 275.65, 
    276.05, 275.95, 276.15, 276.15, 276.05, 275.85, 275.45, 275.05, 275.55, 
    275.65, 275.75, 275.45, 275.75, 275.35, 275.25, 275.45, 275.35, 275.15, 
    275.25, 275.35, 275.95, 276.45, 276.05, 275.95, 275.65, 275.65, 275.55, 
    275.85, 275.65, 275.85, 275.85, 275.95, 275.95, 275.85, 275.55, 275.85, 
    275.65, 275.85, 276.05, 275.55, 275.15, 275.25, 275.35, 275.85, 275.85, 
    275.75, 275.75, 276.35, 275.45, 275.25, 274.45, 273.75, 273.95, 273.65, 
    273.55, 273.45, 273.45, 272.65, 272.95, 273.75, 273.85, 273.85, 273.75, 
    273.85, 274.05, 274.05, 274.25, 274.25, 274.45, 274.65, 274.75, 274.75, 
    274.65, 275.15, 274.55, 274.35, 274.15, 274.05, 273.85, 273.55, 273.35, 
    273.45, 273.35, 273.35, 273.15, 272.95, 272.45, 272.95, 273.05, 273.05, 
    273.15, 273.45, 273.75, 273.95, 274.25, 273.85, 274.05, 273.35, 273.35, 
    273.75, 273.75, 273.15, 272.25, 271.95, 272.05, 272.55, 272.55, 273.35, 
    273.15, 272.85, 272.65, 272.65, 272.45, 272.25, 272.05, 272.15, 272.05, 
    272.35, 272.35, 272.15, 271.95, 271.85, 271.55, 271.75, 272.15, 270.95, 
    270.65, 269.85, 270.45, 270.55, 270.25, 270.75, 271.35, 271.65, 271.75, 
    272.25, 272.55, 272.55, 272.85, 273.05, 273.25, 273.35, 273.45, 273.35, 
    273.45, 273.35, 272.95, 272.95, 272.95, 273.15, 273.45, 273.65, 274.05, 
    274.15, 274.05, 273.85, 273.35, 273.35, 273.35, 273.15, 273.25, 273.35, 
    273.25, 273.05, 273.05, 272.85, 272.85, 273.25, 273.55, 273.55, 273.65, 
    273.65, 273.35, 273.35, 272.35, 272.35, 273.05, 272.85, 272.95, 272.85, 
    272.85, 273.05, 273.15, 273.25, 273.35, 273.25, 273.45, 273.75, 273.85, 
    273.95, 274.05, 274.15, 274.15, 273.75, 273.85, 273.55, 273.75, 273.55, 
    273.35, 273.45, 273.65, 273.85, 274.05, 274.05, 274.05, 274.15, 274.25, 
    274.75, 275.25, 275.45, 275.65, 275.85, 275.85, 276.55, 276.35, 276.05, 
    275.45, 274.75, 274.85, 275.65, 275.85, 276.35, 275.95, 275.75, 275.65, 
    276.35, 277.05, 277.75, 277.55, 276.85, 276.65, 276.15, 275.95, 275.95, 
    275.65, 275.55, 275.35, 274.85, 274.55, 274.25, 273.85, 273.55, 273.85, 
    273.75, 273.35, 273.25, 273.35, 273.35, 273.35, 273.45, 273.45, 274.45, 
    274.45, 274.45, 273.85, 273.35, 273.55, 274.25, 275.05, 275.15, 275.25, 
    275.25, 275.55, 275.75, 275.75, 275.65, 275.15, 274.95, 275.15, 275.15, 
    274.25, 273.95, 274.05, 274.25, 273.85, 273.75, 273.65, 272.85, 274.65, 
    274.55, 274.75, 275.15, 275.95, 275.45, 276.15, 275.55, 275.55, 275.25, 
    275.85, 275.85, 275.75, 275.75, 276.55, 277.95, 278.95, 278.85, 276.95, 
    276.05, 275.85, 275.65, 275.15, 275.05, 275.35, 275.75, 276.15, 275.95, 
    276.35, 277.55, 275.75, 275.45, 276.15, 275.65, 276.35, 277.45, 278.85, 
    276.95, 276.75, 276.85, 277.05, 277.15, 276.15, 275.55, 275.15, 274.85, 
    275.45, 274.75, 274.85, 274.65, 274.35, 274.25, 274.15, 274.65, 274.75, 
    274.65, 275.15, 275.15, 274.95, 274.35, 273.65, 273.75, 273.35, 273.35, 
    273.45, 273.75, 275.65, 276.35, 274.95, 274.85, 274.55, 274.35, 274.45, 
    274.65, 276.85, 276.75, 276.55, 276.75, 276.35, 276.35, 276.65, 276.85, 
    276.85, 276.05, 275.55, 275.35, 275.35, 275.35, 275.35, 274.95, 274.45, 
    274.55, 274.65, 274.95, 274.85, 274.95, 274.85, 274.55, 274.35, 274.25, 
    273.95, 273.75, 273.55, 273.85, 274.15, 274.35, 274.35, 274.25, 274.25, 
    273.85, 273.85, 273.95, 273.85, 273.95, 273.65, 273.85, 273.65, 273.65, 
    273.55, 273.65, 274.15, 273.95, 273.85, 273.75, 273.65, 273.55, 273.85, 
    273.75, 273.75, 274.05, 274.35, 274.35, 274.05, 274.15, 273.95, 273.95, 
    274.15, 274.55, 274.15, 273.95, 274.45, 274.35, 274.15, 274.05, 274.25, 
    274.25, 274.25, 273.65, 273.45, 273.45, 273.45, 273.95, 274.25, 274.25, 
    274.45, 274.55, 274.75, 274.65, 274.25, 273.85, 273.75, 274.05, 273.95, 
    274.15, 273.65, 273.85, 273.75, 274.05, 273.75, 273.75, 274.05, 273.95, 
    274.45, 274.05, 273.95, 273.85, 273.75, 273.75, 274.15, 273.95, 273.75, 
    274.25, 274.35, 274.25, 274.05, 273.75, 273.55, 273.65, 273.65, 273.55, 
    273.45, 273.45, 273.35, 273.85, 274.25, 273.45, 273.35, 273.65, 273.65, 
    273.55, 273.45, 273.65, 273.75, 273.45, 273.75, 273.05, 272.85, 272.95, 
    272.95, 272.95, 272.45, 272.35, 272.65, 272.85, 272.55, 272.95, 272.95, 
    273.05, 273.25, 273.25, 273.15, 273.15, 273.15, 273.15, 273.45, 273.25, 
    273.35, 273.35, 273.05, 273.25, 273.15, 272.85, 272.95, 272.95, 272.65, 
    272.55, 272.25, 272.15, 272.25, 272.35, 272.45, 272.65, 272.45, 272.45, 
    272.65, 273.15, 273.05, 273.05, 273.05, 273.05, 273.35, 273.45, 273.45, 
    272.35, 273.55, 273.35, 273.75, 273.65, 273.65, 273.95, 274.05, 273.85, 
    273.85, 273.85, 273.55, 273.45, 273.65, 273.15, 273.75, 273.75, 273.75, 
    273.85, 274.15, 274.25, 273.65, 273.55, 273.75, 273.85, 273.85, 273.95, 
    274.25, 273.55, 273.75, 273.85, 273.65, 273.45, 273.35, 273.05, 272.85, 
    272.85, 272.85, 272.75, 272.65, 273.55, 273.55, 273.75, 273.85, 273.95, 
    274.25, 274.35, 274.55, 274.65, 274.85, 275.05, 275.05, 275.15, 274.65, 
    274.95, 275.05, 274.75, 275.15, 274.95, 275.25, 275.35, 275.45, 275.35, 
    275.55, 275.55, 275.55, 275.75, 275.55, 275.35, 275.25, 274.85, 274.85, 
    275.05, 275.05, 274.85, 274.85, 274.95, 274.95, 275.05, 275.25, 275.25, 
    275.35, 275.35, 275.35, 275.55, 275.55, 275.65, 275.65, 275.85, 275.75, 
    275.65, 275.65, 275.35, 275.15, 274.95, 275.15, 275.35, 275.15, 274.95, 
    274.65, 274.65, 274.55, 274.65, 274.05, 273.35, 273.25, 273.45, 273.55, 
    273.65, 274.45, 274.45, 274.55, 274.45, 273.75, 274.25, 274.25, 273.85, 
    273.65, 274.05, 274.25, 274.05, 273.85, 273.65, 273.85, 274.15, 273.55, 
    273.85, 273.55, 273.65, 273.35, 273.25, 273.35, 273.75, 273.65, 273.75, 
    273.85, 273.45, 273.05, 272.65, 272.85, 272.65, 272.85, 272.85, 272.55, 
    272.65, 272.25, 272.15, 271.75, 271.75, 271.65, 271.65, 271.85, 272.35, 
    272.95, 273.15, 273.05, 273.05, 272.95, 272.35, 272.55, 271.95, 271.65, 
    271.65, 271.55, 271.65, 271.35, 271.45, 271.15, 271.05, 271.05, 271.05, 
    271.15, 271.35, 271.35, 271.45, 271.75, 271.95, 272.25, 272.55, 272.85, 
    272.85, 273.05, 272.95, 272.75, 272.95, 272.75, 272.55, 272.35, 272.25, 
    271.45, 271.55, 271.55, 271.85, 271.85, 271.35, 271.55, 271.85, 271.85, 
    271.45, 271.45, 270.85, 269.75, 269.65, 270.25, 270.25, 269.85, 268.75, 
    268.85, 269.75, 269.95, 269.95, 270.05, 269.95, 269.75, 269.55, 269.35, 
    269.25, 269.25, 269.15, 269.15, 269.15, 269.65, 269.35, 269.45, 269.45, 
    269.45, 269.15, 269.35, 269.75, 269.65, 269.45, 269.35, 269.45, 269.45, 
    269.45, 269.65, 269.15, 269.05, 269.25, 269.35, 269.25, 269.45, 269.55, 
    269.25, 269.25, 268.95, 269.15, 268.95, 269.65, 269.55, 269.55, 269.25, 
    268.95, 268.75, 268.55, 268.45, 268.05, 268.05, 268.05, 268.65, 268.95, 
    270.15, 270.95, 270.25, 269.55, 268.75, 268.45, 271.15, 270.85, 271.05, 
    271.35, 271.65, 271.75, 271.55, 271.65, 271.75, 271.75, 272.15, 272.05, 
    272.25, 271.85, 271.45, 271.95, 271.15, 270.25, 271.15, 272.25, 271.75, 
    271.35, 271.35, 271.15, 271.15, 271.35, 270.85, 269.65, 269.75, 270.25, 
    271.05, 271.45, 271.75, 272.35, 272.55, 273.15, 273.25, 273.45, 273.45, 
    273.85, 273.75, 274.15, 274.05, 274.55, 274.35, 274.35, 274.35, 274.15, 
    274.05, 273.75, 273.75, 273.75, 273.55, 273.35, 273.45, 273.55, 273.45, 
    272.95, 272.75, 272.65, 272.55, 272.25, 272.35, 272.45, 272.05, 272.05, 
    272.25, 271.55, 271.95, 271.65, 270.95, 270.65, 270.75, 270.95, 271.85, 
    270.55, 270.45, 270.45, 270.15, 269.85, 270.35, 270.55, 271.25, 271.25, 
    270.75, 271.45, 271.25, 271.65, 271.75, 271.85, 271.65, 271.35, 271.25, 
    270.55, 270.55, 270.15, 270.15, 270.45, 270.45, 270.35, 270.05, 270.25, 
    269.95, 270.25, 269.85, 269.45, 269.35, 269.55, 268.85, 268.25, 267.95, 
    267.45, 267.15, 266.55, 267.65, 267.45, 267.15, 267.45, 266.65, 267.05, 
    267.05, 267.75, 267.65, 268.85, 266.25, 266.75, 267.15, 267.45, 267.65, 
    267.65, 267.05, 266.75, 266.35, 265.85, 265.35, 266.25, 265.85, 267.05, 
    267.15, 267.25, 267.55, 267.45, 267.95, 267.35, 267.35, 267.95, 267.55, 
    268.05, 266.35, 266.95, 267.25, 266.35, 266.55, 265.35, 265.35, 266.45, 
    266.35, 266.35, 267.05, 266.65, 266.05, 266.45, 266.45, 266.65, 266.45, 
    266.85, 265.55, 266.35, 267.45, 265.45, 266.95, 267.05, 267.45, 267.95, 
    266.85, 266.55, 265.05, 265.65, 264.15, 266.35, 265.55, 265.15, 265.35, 
    266.25, 267.45, 268.55, 269.75, 268.35, 269.15, 268.85, 268.65, 268.05, 
    268.25, 267.95, 266.25, 267.05, 268.15, 268.75, 267.85, 267.25, 266.65, 
    266.15, 265.35, 265.45, 265.05, 264.95, 264.85, 264.05, 264.85, 264.55, 
    263.15, 262.95, 262.85, 263.05, 263.65, 264.25, 264.85, 264.65, 264.25, 
    264.95, 265.25, 266.75, 267.75, 268.05, 268.35, 266.85, 266.95, 267.15, 
    266.85, 266.65, 266.25, 266.95, 266.45, 265.55, 265.25, 265.95, 265.35, 
    267.05, 266.65, 267.25, 267.25, 267.15, 267.35, 267.05, 266.55, 266.15, 
    265.65, 266.05, 265.95, 265.35, 265.15, 265.35, 265.65, 265.55, 265.25, 
    264.95, 264.65, 264.85, 265.15, 265.55, 265.15, 265.85, 265.25, 266.15, 
    265.35, 265.25, 265.15, 265.85, 265.55, 265.85, 265.35, 265.45, 265.45, 
    265.35, 265.05, 266.25, 266.15, 266.15, 266.15, 265.45, 266.35, 265.65, 
    265.85, 265.55, 265.05, 265.45, 265.65, 265.65, 265.35, 265.45, 265.05, 
    265.25, 264.85, 264.15, 264.65, 265.35, 266.15, 266.35, 265.55, 267.25, 
    266.45, 266.65, 267.85, 268.55, 268.85, 269.35, 269.95, 269.35, 269.65, 
    268.65, 268.05, 267.25, 265.95, 265.35, 265.95, 267.75, 266.75, 266.45, 
    266.55, 266.45, 266.25, 266.05, 266.05, 266.15, 266.35, 266.75, 267.15, 
    267.95, 268.65, 269.45, 269.55, 268.95, 268.15, 267.95, 267.75, 267.25, 
    266.35, 265.95, 265.85, 265.25, 264.65, 263.85, 265.25, 265.25, 265.25, 
    264.95, 264.75, 264.35, 264.05, 263.95, 263.95, 263.65, 263.45, 263.05, 
    263.25, 264.05, 264.15, 264.05, 264.35, 264.25, 264.25, 264.35, 264.45, 
    264.35, 264.25, 264.05, 264.45, 264.65, 264.45, 264.65, 263.55, 263.55, 
    263.75, 264.15, 263.75, 263.65, 263.25, 263.05, 262.85, 262.75, 262.65, 
    263.15, 263.15, 262.95, 263.05, 263.05, 262.85, 263.05, 262.85, 262.85, 
    263.05, 262.95, 263.15, 263.05, 263.35, 263.45, 263.35, 263.05, 262.35, 
    261.85, 262.05, 261.95, 262.45, 262.55, 262.75, 262.95, 263.15, 263.35, 
    263.55, 263.65, 263.45, 263.75, 263.25, 263.15, 262.75, 262.15, 261.85, 
    261.95, 262.15, 262.15, 262.55, 262.55, 262.45, 262.85, 262.95, 262.95, 
    263.15, 263.35, 263.35, 263.75, 264.15, 264.25, 264.45, 264.75, 264.35, 
    264.15, 264.15, 264.35, 264.25, 264.25, 264.15, 264.25, 264.05, 263.85, 
    263.65, 263.65, 263.45, 263.45, 263.15, 263.05, 263.25, 263.05, 263.15, 
    263.25, 263.25, 263.05, 261.65, 261.35, 261.35, 261.25, 261.25, 260.75, 
    261.25, 260.75, 259.45, 259.95, 260.85, 261.05, 261.55, 261.45, 261.15, 
    260.85, 262.35, 261.25, 261.75, 261.85, 261.45, 261.85, 262.55, 262.45, 
    263.85, 262.95, 261.85, 262.45, 262.75, 261.55, 261.35, 261.65, 261.35, 
    260.45, 259.55, 260.05, 261.05, 260.55, 260.35, 259.95, 260.95, 261.65, 
    262.95, 262.95, 261.45, 261.85, 262.95, 262.05, 262.25, 262.85, 262.15, 
    262.55, 261.75, 262.05, 262.25, 262.15, 262.95, 262.15, 262.15, 262.25, 
    262.55, 262.35, 262.55, 262.85, 263.15, 263.25, 263.65, 263.95, 263.75, 
    263.65, 263.75, 263.35, 262.95, 263.65, 263.05, 263.15, 263.75, 261.65, 
    262.15, 263.35, 262.65, 262.95, 262.65, 262.45, 262.35, 262.25, 262.45, 
    262.25, 261.95, 262.05, 262.05, 262.15, 262.05, 261.75, 261.35, 261.35, 
    261.35, 261.45, 261.35, 261.55, 261.35, 261.25, 261.25, 261.35, 261.25, 
    261.65, 261.25, 261.35, 261.85, 260.45, 260.15, 259.85, 260.15, 260.25, 
    260.75, 260.85, 261.65, 260.75, 261.35, 260.45, 262.15, 261.75, 262.35, 
    262.55, 262.75, 263.15, 263.15, 263.25, 263.95, 263.25, 263.65, 263.85, 
    264.55, 265.15, 264.95, 265.15, 264.55, 265.65, 265.75, 265.85, 265.95, 
    266.05, 266.25, 266.55, 266.85, 266.95, 267.45, 267.85, 268.15, 268.15, 
    268.25, 268.45, 268.85, 269.25, 269.55, 269.75, 269.75, 269.85, 270.05, 
    270.85, 271.45, 270.75, 270.75, 270.85, 270.65, 270.85, 270.55, 270.15, 
    270.05, 270.55, 269.05, 267.45, 268.55, 270.45, 270.45, 270.25, 269.25, 
    268.75, 269.15, 268.25, 267.95, 267.65, 267.15, 266.75, 266.75, 266.75, 
    266.75, 266.75, 266.55, 266.25, 265.55, 265.65, 265.35, 265.05, 265.15, 
    264.95, 265.45, 265.55, 265.95, 265.95, 266.35, 266.55, 266.85, 267.05, 
    267.55, 267.85, 268.15, 268.45, 268.45, 269.05, 269.75, 270.05, 270.35, 
    270.85, 271.15, 271.45, 271.85, 272.15, 272.45, 272.85, 273.05, 272.85, 
    272.35, 271.75, 270.95, 270.75, 270.65, 270.65, 270.45, 270.45, 270.65, 
    271.15, 269.95, 269.55, 269.35, 269.05, 269.15, 269.05, 269.25, 269.15, 
    269.25, 269.05, 269.05, 269.15, 269.05, 268.85, 268.75, 269.35, 268.85, 
    268.35, 268.75, 269.05, 268.75, 268.55, 268.45, 268.25, 268.45, 268.45, 
    268.25, 267.65, 267.35, 267.35, 267.35, 267.65, 267.75, 268.15, 268.45, 
    267.75, 267.65, 266.45, 266.85, 266.55, 267.85, 267.15, 266.95, 266.65, 
    266.35, 265.55, 264.25, 263.75, 263.65, 263.75, 263.85, 264.55, 264.65, 
    264.55, 264.05, 263.75, 263.65, 263.55, 263.35, 263.35, 263.15, 263.15, 
    263.25, 263.45, 263.55, 263.65, 263.85, 263.95, 263.85, 262.75, 262.45, 
    262.45, 262.75, 264.25, 265.55, 265.85, 265.95, 265.85, 266.35, 266.35, 
    267.75, 266.55, 267.15, 268.15, 268.35, 267.55, 269.55, 269.85, 269.85, 
    270.15, 270.45, 270.55, 270.55, 270.85, 270.95, 270.75, 270.65, 270.65, 
    270.35, 270.35, 270.05, 270.25, 270.85, 270.55, 270.55, 270.75, 270.75, 
    270.35, 270.25, 270.55, 270.75, 270.85, 270.75, 270.35, 270.75, 270.85, 
    271.15, 271.35, 271.65, 272.05, 272.15, 271.15, 269.95, 268.65, 267.75, 
    266.75, 266.15, 266.05, 265.95, 265.65, 265.55, 265.15, 264.95, 264.55, 
    264.45, 264.65, 264.55, 264.75, 264.75, 264.95, 264.95, 264.95, 264.75, 
    265.05, 264.55, 264.75, 264.55, 264.75, 265.15, 265.25, 264.95, 265.15, 
    265.05, 264.75, 264.35, 264.65, 264.95, 264.05, 263.85, 263.65, 264.95, 
    265.25, 265.55, 265.75, 265.85, 265.15, 264.85, 264.35, 264.05, 263.65, 
    263.45, 263.95, 263.55, 263.25, 263.15, 262.95, 263.15, 262.85, 262.85, 
    262.75, 262.65, 262.65, 262.75, 262.75, 262.75, 262.75, 262.45, 262.65, 
    262.75, 262.45, 262.55, 262.45, 262.35, 262.25, 262.45, 262.35, 262.65, 
    262.55, 262.55, 262.95, 263.25, 263.85, 263.75, 265.05, 265.75, 265.15, 
    266.75, 267.45, 267.85, 268.45, 268.45, 268.25, 268.15, 268.05, 268.45, 
    268.75, 268.85, 269.25, 269.75, 270.15, 270.25, 270.85, 271.45, 271.75, 
    271.85, 272.05, 272.15, 272.25, 272.45, 272.45, 272.45, 272.45, 272.45, 
    272.45, 272.45, 272.45, 272.45, 272.45, 272.35, 272.15, 271.05, 270.75, 
    269.45, 268.95, 268.65, 268.35, 267.85, 267.65, 267.45, 267.55, 267.85, 
    267.85, 268.35, 268.45, 269.35, 271.25, 272.45, 272.45, 272.45, 272.45, 
    272.55, 272.45, 272.45, 272.65, 271.95, 270.35, 267.45, 267.25, 266.85, 
    266.95, 266.85, 266.45, 266.85, 266.85, 266.85, 267.25, 267.25, 267.65, 
    268.05, 268.05, 268.15, 268.35, 268.35, 268.25, 268.15, 268.15, 267.95, 
    267.75, 267.85, 267.65, 267.45, 267.25, 267.45, 267.55, 267.55, 267.85, 
    267.85, 267.95, 267.65, 267.65, 267.25, 266.85, 267.15, 266.95, 266.75, 
    266.95, 267.15, 267.35, 267.75, 267.95, 267.65, 267.95, 267.35, 268.05, 
    268.25, 268.25, 268.25, 268.55, 268.85, 268.75, 268.15, 267.45, 266.75, 
    266.45, 266.05, 266.45, 266.25, 265.85, 265.45, 265.25, 265.05, 264.55, 
    264.75, 264.65, 264.45, 264.45, 264.45, 264.25, 263.65, 263.35, 263.75, 
    264.15, 263.45, 263.35, 263.75, 264.05, 264.05, 263.75, 263.55, 263.75, 
    263.35, 263.65, 262.85, 263.25, 262.45, 263.45, 263.55, 263.25, 263.25, 
    262.55, 263.35, 263.15, 261.75, 262.05, 262.45, 261.45, 262.05, 262.65, 
    263.85, 264.25, 265.65, 266.05, 266.85, 267.75, 268.35, 269.75, 269.75, 
    269.75, 269.35, 269.55, 270.35, 270.95, 271.35, 271.15, 271.15, 271.15, 
    270.95, 270.55, 269.95, 270.15, 270.05, 270.15, 270.05, 270.05, 270.55, 
    270.95, 271.25, 271.45, 271.25, 271.05, 270.85, 271.15, 271.35, 271.65, 
    271.75, 271.55, 271.45, 271.45, 271.65, 271.75, 271.75, 271.85, 272.05, 
    272.05, 271.95, 271.95, 271.85, 271.65, 271.45, 271.35, 271.05, 270.75, 
    270.75, 270.65, 270.55, 270.15, 270.25, 270.25, 269.85, 269.75, 269.75, 
    269.55, 269.55, 268.95, 269.05, 268.85, 268.65, 268.45, 268.35, 268.15, 
    267.75, 266.95, 266.75, 266.75, 266.75, 266.35, 265.85, 265.15, 264.65, 
    264.55, 263.85, 263.85, 263.45, 263.25, 263.25, 262.55, 262.55, 262.65, 
    262.25, 262.35, 262.15, 261.75, 261.85, 261.85, 261.85, 261.55, 261.35, 
    261.25, 261.25, 260.55, 260.55, 260.15, 260.15, 260.05, 259.75, 259.65, 
    259.15, 258.75, 258.45, 258.25, 258.25, 258.55, 258.95, 258.95, 258.85, 
    259.15, 258.85, 259.35, 259.45, 259.65, 259.55, 259.75, 259.85, 259.95, 
    259.85, 259.85, 259.75, 259.85, 260.25, 260.15, 260.55, 260.45, 261.05, 
    259.75, 257.85, 257.45, 258.45, 258.15, 258.45, 258.15, 258.05, 258.95, 
    258.95, 261.15, 260.35, 260.15, 260.45, 260.65, 260.75, 260.65, 261.15, 
    260.65, 260.55, 260.45, 260.65, 260.35, 260.15, 259.85, 259.85, 259.95, 
    259.65, 259.85, 259.75, 260.05, 260.25, 260.15, 259.65, 259.15, 259.05, 
    258.55, 257.95, 257.65, 257.65, 257.75, 257.85, 257.85, 257.85, 257.95, 
    258.35, 258.55, 258.85, 258.75, 258.65, 259.05, 259.25, 259.35, 259.15, 
    259.25, 259.35, 259.15, 258.95, 258.95, 259.05, 259.35, 258.95, 258.65, 
    258.25, 258.35, 258.45, 257.55, 257.25, 256.85, 257.05, 257.35, 256.65, 
    256.85, 256.65, 256.65, 256.65, 256.45, 255.15, 254.55, 253.75, 254.65, 
    255.35, 255.05, 256.15, 256.25, 256.55, 256.75, 257.05, 256.35, 256.45, 
    257.35, 255.85, 255.75, 255.25, 255.85, 256.95, 256.55, 257.05, 256.95, 
    257.55, 257.65, 257.45, 257.75, 257.45, 257.15, 256.95, 256.75, 256.55, 
    256.35, 256.25, 256.05, 256.55, 256.25, 257.45, 258.05, 258.25, 258.05, 
    258.25, 259.05, 259.45, 259.55, 259.35, 259.45, 260.15, 260.85, 260.45, 
    260.55, 260.45, 260.25, 260.15, 262.45, 262.35, 262.15, 262.35, 262.65, 
    263.25, 263.55, 263.45, 263.45, 262.85, 262.85, 262.85, 262.85, 262.75, 
    262.65, 262.95, 262.75, 262.65, 262.35, 262.15, 261.95, 261.45, 260.95, 
    260.75, 260.15, 259.65, 259.25, 258.65, 258.65, 258.15, 258.15, 257.75, 
    256.95, 257.45, 256.95, 256.85, 254.85, 254.35, 253.55, 253.55, 253.55, 
    253.55, 253.35, 253.45, 253.45, 253.35, 253.15, 253.95, 253.55, 252.85, 
    253.15, 253.55, 253.95, 254.45, 255.05, 255.85, 256.75, 256.05, 256.75, 
    258.15, 259.05, 256.45, 256.55, 256.35, 256.25, 257.75, 257.85, 257.25, 
    256.35, 256.45, 256.65, 256.65, 257.65, 257.45, 257.45, 256.75, 256.75, 
    255.95, 256.05, 255.55, 255.35, 254.95, 254.45, 254.45, 254.55, 254.25, 
    254.05, 254.45, 254.25, 254.45, 254.45, 254.85, 254.95, 255.15, 255.95, 
    256.25, 256.55, 255.25, 257.25, 257.55, 257.05, 257.35, 257.45, 257.25, 
    257.85, 257.95, 257.85, 257.65, 256.85, 256.85, 257.15, 257.15, 257.15, 
    256.45, 256.45, 258.25, 259.15, 259.85, 260.35, 260.25, 260.45, 260.15, 
    259.85, 259.75, 259.95, 259.85, 259.85, 259.45, 259.15, 258.15, 257.85, 
    257.45, 257.35, 257.05, 257.95, 258.65, 259.55, 259.45, 259.35, 258.85, 
    258.55, 258.55, 258.35, 258.15, 258.05, 257.95, 258.05, 258.05, 258.05, 
    258.25, 257.95, 257.95, 257.85, 257.95, 257.55, 257.45, 257.55, 257.85, 
    257.25, 256.55, 255.95, 256.15, 256.25, 256.45, 257.05, 258.15, 257.75, 
    257.65, 258.55, 260.75, 261.55, 262.25, 263.35, 265.05, 265.05, 264.45, 
    263.15, 262.45, 261.85, 262.15, 262.05, 260.35, 259.15, 258.05, 257.35, 
    257.55, 261.35, 259.35, 262.05, 257.55, 258.95, 259.35, 260.05, 259.45, 
    258.85, 257.15, 257.35, 256.65, 258.05, 256.95, 257.55, 256.85, 256.55, 
    255.65, 257.95, 260.05, 259.25, 260.75, 262.35, 261.85, 261.35, 261.15, 
    261.05, 260.75, 260.65, 260.85, 261.25, 262.25, 262.45, 264.05, 265.05, 
    265.45, 266.05, 266.55, 266.75, 266.35, 265.35, 264.45, 263.25, 263.05, 
    263.15, 263.15, 263.55, 263.65, 263.25, 262.75, 262.35, 261.95, 261.65, 
    262.15, 262.75, 260.45, 260.55, 260.75, 260.85, 260.85, 259.95, 259.55, 
    258.55, 258.25, 258.65, 260.15, 260.65, 260.25, 260.45, 260.65, 260.45, 
    259.95, 259.45, 260.15, 258.75, 258.85, 259.25, 259.25, 259.15, 259.75, 
    259.55, 259.85, 260.35, 260.75, 261.25, 261.25, 261.85, 263.05, 262.65, 
    263.25, 263.05, 263.25, 263.45, 264.25, 265.05, 266.15, 267.05, 267.45, 
    267.95, 268.25, 269.15, 269.45, 269.45, 269.75, 270.15, 270.05, 270.55, 
    270.55, 270.45, 270.55, 270.05, 270.05, 267.65, 269.15, 268.15, 267.35, 
    267.95, 268.05, 267.65, 267.45, 267.55, 268.15, 268.85, 268.45, 268.35, 
    268.75, 268.75, 269.35, 269.75, 270.15, 270.55, 270.75, 271.05, 271.15, 
    271.55, 271.65, 271.65, 271.65, 271.75, 271.85, 272.05, 272.15, 272.25, 
    272.25, 272.25, 272.85, 273.15, 272.95, 272.85, 272.55, 272.35, 272.25, 
    272.15, 272.25, 272.25, 272.25, 272.45, 272.55, 272.65, 272.75, 272.75, 
    272.55, 272.35, 272.45, 272.55, 272.45, 272.25, 272.35, 272.05, 272.15, 
    272.35, 272.25, 272.25, 272.25, 272.25, 272.15, 272.15, 272.15, 272.15, 
    272.15, 272.05, 271.55, 271.25, 271.35, 271.35, 270.05, 269.55, 269.05, 
    268.85, 268.55, 269.15, 269.35, 269.45, 268.85, 268.45, 268.35, 267.45, 
    268.05, 267.95, 267.85, 267.65, 267.05, 267.45, 267.35, 267.35, 268.35, 
    268.05, 267.95, 268.15, 267.85, 268.35, 267.55, 267.35, 266.85, 266.95, 
    266.75, 266.85, 268.25, 268.75, 268.95, 269.15, 269.15, 269.25, 269.35, 
    269.25, 269.05, 269.25, 269.45, 269.65, 269.55, 269.35, 268.85, 268.35, 
    268.45, 268.85, 269.05, 269.45, 269.65, 268.85, 268.95, 268.75, 269.05, 
    269.25, 269.35, 268.85, 268.75, 268.75, 268.65, 268.55, 268.05, 267.85, 
    267.15, 266.65, 267.05, 267.15, 266.65, 267.25, 267.55, 267.45, 267.15, 
    266.35, 266.95, 267.35, 267.35, 267.75, 267.85, 267.75, 267.65, 268.05, 
    267.65, 267.85, 268.05, 268.15, 268.05, 267.85, 267.95, 267.55, 267.75, 
    267.55, 266.95, 265.95, 264.85, 264.35, 263.35, 262.35, 261.85, 261.55, 
    261.05, 261.15, 260.95, 261.15, 261.15, 261.05, 261.65, 261.85, 261.65, 
    261.95, 261.85, 261.85, 261.65, 261.65, 261.95, 261.85, 261.65, 261.55, 
    261.35, 261.15, 261.15, 261.05, 260.55, 260.05, 259.65, 259.75, 259.45, 
    259.25, 258.85, 258.55, 258.45, 258.25, 258.05, 257.65, 257.65, 257.75, 
    257.85, 257.75, 257.75, 258.35, 258.85, 258.95, 258.65, 258.85, 258.05, 
    257.45, 258.15, 257.55, 257.65, 256.25, 256.35, 256.55, 257.25, 256.85, 
    257.05, 258.85, 258.35, 256.05, 255.35, 255.65, 256.85, 257.05, 257.45, 
    257.75, 257.95, 258.45, 258.75, 258.65, 259.35, 259.15, 259.05, 259.25, 
    258.95, 259.35, 259.55, 259.55, 259.65, 259.55, 259.45, 259.45, 259.35, 
    259.35, 258.95, 259.15, 258.55, 258.75, 258.65, 259.05, 259.55, 259.45, 
    259.15, 259.05, 258.65, 259.15, 258.85, 259.05, 258.65, 258.85, 259.25, 
    258.75, 258.85, 258.85, 258.65, 259.05, 258.85, 260.15, 259.05, 259.35, 
    259.35, 259.05, 258.25, 257.95, 257.75, 255.85, 254.45, 255.55, 256.45, 
    255.65, 254.55, 255.45, 256.05, 256.35, 256.65, 257.25, 257.35, 257.85, 
    258.15, 258.35, 258.05, 258.15, 258.45, 258.35, 258.75, 258.55, 259.15, 
    259.25, 258.95, 258.45, 258.35, 257.45, 257.05, 257.15, 256.95, 256.85, 
    256.85, 257.35, 256.75, 257.05, 257.55, 257.15, 257.35, 256.85, 257.25, 
    257.65, 257.65, 256.35, 256.95, 256.55, 255.15, 254.95, 256.25, 256.35, 
    256.35, 257.05, 256.55, 255.85, 257.05, 256.75, 256.45, 254.35, 258.25, 
    254.35, 257.25, 256.65, 257.15, 255.55, 255.85, 256.45, 255.75, 256.05, 
    255.75, 255.15, 254.85, 254.65, 255.15, 254.85, 254.85, 254.35, 254.55, 
    254.95, 255.55, 254.75, 255.65, 254.85, 254.35, 254.25, 254.55, 253.95, 
    253.75, 253.75, 252.85, 252.95, 253.25, 252.95, 253.35, 253.75, 253.65, 
    254.45, 255.35, 254.65, 255.05, 255.35, 255.55, 256.95, 257.75, 257.55, 
    257.45, 257.35, 257.55, 258.15, 258.45, 258.85, 258.95, 259.55, 260.05, 
    260.35, 259.85, 259.45, 259.45, 260.15, 260.05, 259.75, 260.15, 259.95, 
    259.75, 258.45, 260.55, 260.75, 260.55, 260.85, 260.65, 260.85, 261.25, 
    261.75, 261.95, 262.15, 262.55, 263.65, 264.65, 265.95, 266.75, 266.95, 
    267.25, 267.65, 268.05, 268.25, 268.05, 268.05, 266.25, 266.75, 266.95, 
    267.25, 266.85, 264.85, 266.35, 266.35, 266.05, 265.55, 265.45, 265.15, 
    264.75, 264.95, 264.55, 264.15, 264.55, 264.15, 265.05, 265.25, 266.05, 
    266.35, 266.75, 267.15, 267.65, 265.35, 264.25, 263.95, 263.75, 263.55, 
    263.65, 263.75, 262.75, 263.05, 262.35, 262.45, 262.15, 262.15, 261.95, 
    261.65, 261.25, 261.15, 261.25, 261.05, 260.85, 260.95, 260.55, 260.15, 
    259.95, 259.75, 259.25, 258.15, 257.45, 257.95, 258.15, 258.65, 257.55, 
    257.95, 259.25, 258.45, 258.25, 258.45, 258.85, 258.35, 258.25, 258.05, 
    258.45, 258.35, 258.95, 259.65, 259.75, 259.35, 259.25, 259.05, 258.85, 
    258.55, 258.55, 258.75, 258.65, 258.45, 258.15, 257.85, 257.75, 257.55, 
    257.25, 257.05, 256.45, 256.25, 256.15, 256.65, 257.15, 256.85, 256.65, 
    253.55, 253.45, 252.55, 252.55, 253.75, 252.45, 253.95, 254.45, 254.05, 
    253.85, 252.95, 253.15, 252.55, 253.35, 253.75, 253.75, 253.95, 253.75, 
    253.55, 253.35, 253.05, 252.45, 252.35, 251.95, 252.85, 252.15, 252.95, 
    253.15, 253.35, 252.75, 252.15, 253.35, 253.25, 251.15, 252.05, 252.65, 
    253.65, 254.35, 253.25, 254.15, 256.65, 256.95, 257.75, 256.65, 256.75, 
    255.85, 254.95, 254.75, 254.15, 254.25, 254.45, 254.35, 255.35, 254.15, 
    253.75, 253.95, 253.45, 253.05, 252.65, 252.95, 253.25, 253.05, 253.35, 
    253.65, 253.05, 252.75, 253.25, 252.55, 252.15, 252.05, 252.55, 253.75, 
    253.95, 254.25, 254.45, 256.15, 257.05, 256.75, 256.45, 256.35, 255.55, 
    255.25, 255.35, 256.55, 256.95, 258.05, 257.85, 258.45, 259.15, 259.95, 
    260.65, 261.45, 262.55, 263.55, 264.25, 264.95, 265.65, 266.15, 266.35, 
    266.45, 266.55, 266.75, 267.05, 267.15, 267.25, 267.65, 267.75, 267.85, 
    267.75, 267.65, 267.65, 267.75, 267.65, 267.65, 267.45, 267.15, 267.55, 
    267.95, 267.75, 268.15, 267.55, 266.95, 267.55, 267.25, 266.95, 266.65, 
    266.95, 267.35, 267.65, 268.05, 268.45, 268.55, 268.55, 268.55, 268.45, 
    268.55, 268.15, 267.15, 267.75, 266.55, 267.45, 267.65, 266.85, 266.55, 
    267.55, 267.75, 268.65, 268.95, 268.95, 269.15, 269.55, 269.95, 269.95, 
    270.55, 270.85, 271.05, 270.85, 270.95, 270.65, 269.75, 269.85, 270.15, 
    269.05, 267.85, 267.65, 267.75, 268.05, 267.65, 268.45, 268.35, 268.95, 
    268.95, 268.55, 268.45, 267.75, 266.45, 266.65, 267.45, 266.65, 267.15, 
    266.95, 264.05, 263.85, 264.75, 265.65, 265.35, 267.25, 269.35, 266.95, 
    266.65, 265.55, 264.95, 264.35, 263.75, 262.45, 262.85, 264.05, 264.35, 
    264.15, 263.45, 264.15, 264.75, 264.95, 263.95, 263.05, 264.15, 264.25, 
    261.65, 262.05, 261.55, 262.15, 261.75, 261.15, 260.65, 260.75, 261.35, 
    262.15, 263.05, 263.55, 262.85, 263.15, 263.55, 264.05, 264.05, 265.45, 
    265.75, 266.25, 265.85, 265.05, 266.05, 265.95, 266.45, 266.45, 266.65, 
    266.85, 266.35, 266.35, 265.15, 265.25, 265.85, 266.25, 265.05, 265.75, 
    266.35, 266.35, 267.15, 266.15, 266.55, 267.05, 267.55, 267.55, 267.55, 
    268.05, 268.25, 268.65, 268.85, 269.15, 269.15, 268.75, 268.65, 268.85, 
    269.15, 269.45, 269.45, 269.45, 269.75, 269.25, 269.35, 268.75, 268.55, 
    268.35, 268.35, 268.85, 268.45, 268.25, 268.85, 268.55, 267.95, 268.75, 
    269.25, 268.15, 268.35, 268.45, 268.85, 269.25, 269.55, 269.85, 270.35, 
    269.65, 268.75, 268.65, 268.85, 268.75, 269.05, 269.45, 269.65, 269.55, 
    269.85, 269.95, 270.05, 269.95, 267.75, 265.95, 264.75, 264.15, 263.75, 
    263.55, 263.55, 263.95, 263.85, 263.75, 263.75, 263.45, 263.45, 263.45, 
    263.35, 263.35, 263.35, 263.65, 263.95, 264.05, 264.55, 264.95, 264.95, 
    265.25, 265.45, 265.25, 265.25, 265.45, 265.15, 265.15, 265.35, 265.65, 
    265.75, 265.75, 265.75, 265.75, 265.85, 266.45, 265.55, 265.45, 264.95, 
    264.15, 262.65, 262.65, 262.45, 263.35, 264.15, 263.65, 263.55, 262.95, 
    263.05, 263.55, 264.05, 264.05, 264.25, 264.35, 264.85, 265.45, 266.15, 
    266.65, 266.95, 267.25, 268.55, 268.15, 268.15, 269.15, 269.45, 269.25, 
    269.25, 267.35, 263.75, 262.55, 262.15, 261.55, 260.65, 260.35, 260.45, 
    260.15, 260.95, 261.95, 262.55, 261.65, 261.05, 261.65, 261.95, 262.85, 
    264.05, 264.55, 264.95, 265.45, 265.45, 265.55, 265.95, 265.95, 265.75, 
    266.75, 267.35, 267.65, 268.55, 269.25, 269.55, 269.65, 269.95, 270.35, 
    271.05, 270.75, 270.55, 270.15, 269.95, 270.25, 270.45, 270.35, 271.45, 
    271.35, 271.45, 271.85, 272.15, 271.75, 271.45, 271.05, 271.75, 270.25, 
    269.85, 269.65, 269.15, 268.65, 268.35, 268.25, 267.95, 267.85, 267.85, 
    267.65, 267.55, 267.55, 267.45, 267.25, 267.55, 267.55, 267.65, 267.65, 
    268.25, 268.45, 268.45, 268.85, 268.55, 266.85, 266.65, 267.55, 266.55, 
    266.65, 266.05, 266.15, 266.05, 266.65, 266.55, 266.75, 267.25, 266.25, 
    266.55, 266.65, 267.05, 267.95, 268.05, 268.15, 268.15, 267.65, 267.15, 
    266.35, 265.95, 265.45, 264.85, 264.15, 264.15, 263.75, 263.75, 264.35, 
    264.15, 263.95, 263.95, 263.95, 264.15, 264.15, 264.25, 264.25, 264.85, 
    265.55, 266.05, 266.55, 266.55, 267.75, 269.65, 270.35, 270.55, 270.55, 
    270.35, 270.15, 270.15, 269.95, 269.75, 269.75, 269.75, 269.65, 268.35, 
    267.75, 267.55, 267.45, 267.15, 267.15, 267.15, 266.85, 266.95, 266.95, 
    266.35, 266.25, 266.65, 267.05, 267.55, 267.85, 267.85, 267.75, 267.55, 
    267.55, 267.65, 267.55, 267.65, 267.65, 267.65, 267.35, 267.65, 267.25, 
    267.05, 267.05, 266.55, 266.05, 265.85, 266.95, 265.05, 265.85, 266.15, 
    267.25, 267.65, 268.15, 268.15, 268.15, 267.35, 267.65, 267.85, 267.85, 
    267.95, 267.85, 267.85, 267.75, 267.75, 268.15, 268.15, 267.85, 267.45, 
    267.25, 267.35, 267.35, 267.25, 267.25, 267.45, 267.45, 267.45, 267.55, 
    267.95, 268.35, 268.55, 268.45, 268.35, 268.45, 268.35, 268.35, 267.55, 
    267.25, 267.85, 268.55, 268.55, 268.45, 268.35, 268.15, 268.25, 268.15, 
    267.95, 267.65, 267.35, 267.25, 267.55, 267.35, 268.15, 267.85, 266.85, 
    266.45, 267.05, 267.65, 267.65, 267.75, 267.65, 267.35, 267.65, 266.65, 
    267.45, 266.25, 265.75, 266.45, 266.85, 266.75, 267.05, 267.35, 267.25, 
    267.45, 267.45, 267.95, 267.95, 269.05, 268.85, 268.55, 268.35, 269.15, 
    269.55, 268.65, 269.05, 269.45, 269.45, 268.95, 268.25, 267.75, 267.95, 
    268.65, 267.65, 268.45, 266.85, 268.15, 268.45, 266.65, 266.85, 266.65, 
    266.75, 267.15, 267.05, 267.65, 267.75, 267.75, 269.05, 269.65, 269.85, 
    269.45, 269.45, 269.55, 269.95, 269.95, 269.25, 268.75, 268.45, 267.65, 
    268.05, 268.25, 269.15, 269.35, 270.05, 270.25, 270.15, 270.15, 270.15, 
    270.25, 270.35, 270.55, 270.45, 270.35, 270.35, 270.35, 270.15, 270.05, 
    269.95, 269.95, 269.95, 269.95, 269.95, 269.85, 269.75, 269.85, 269.85, 
    269.95, 269.65, 269.85, 269.95, 270.15, 270.25, 270.45, 270.55, 270.75, 
    270.85, 271.05, 271.15, 271.25, 271.35, 271.35, 271.35, 271.25, 271.25, 
    271.25, 271.15, 271.05, 270.45, 270.25, 270.15, 269.75, 269.55, 269.45, 
    269.85, 270.15, 270.55, 270.25, 270.15, 270.35, 270.15, 269.45, 268.25, 
    268.05, 267.55, 268.35, 269.15, 269.65, 269.75, 269.85, 269.55, 269.55, 
    269.55, 269.65, 268.95, 268.85, 268.75, 269.15, 269.55, 269.75, 269.85, 
    269.25, 269.45, 269.45, 269.25, 269.45, 269.25, 268.85, 268.65, 268.85, 
    268.95, 269.05, 269.05, 269.05, 268.95, 269.05, 269.15, 269.35, 269.25, 
    269.15, 268.85, 268.55, 268.05, 268.15, 268.25, 268.05, 268.25, 268.95, 
    269.35, 268.95, 268.85, 268.65, 268.25, 268.75, 268.35, 268.35, 269.05, 
    269.85, 269.95, 270.15, 270.35, 270.45, 270.15, 270.05, 269.75, 269.65, 
    269.45, 269.45, 269.45, 269.45, 269.75, 270.35, 270.55, 270.45, 270.65, 
    270.55, 270.25, 270.35, 270.35, 270.25, 269.55, 268.95, 269.05, 268.75, 
    268.55, 268.55, 268.65, 268.55, 268.75, 268.65, 268.75, 268.85, 268.95, 
    269.05, 269.05, 269.05, 268.95, 269.05, 269.15, 269.55, 269.45, 269.45, 
    269.45, 269.45, 269.35, 269.35, 269.25, 269.25, 269.25, 269.05, 269.15, 
    269.85, 270.15, 270.25, 270.55, 270.45, 270.65, 270.75, 270.85, 270.85, 
    270.95, 270.85, 270.85, 270.85, 270.95, 270.85, 271.05, 271.35, 271.75, 
    272.05, 272.15, 272.25, 272.45, 272.45, 272.55, 272.55, 272.65, 272.75, 
    272.75, 273.25, 273.45, 273.45, 273.25, 273.35, 273.15, 273.25, 273.45, 
    273.55, 273.65, 273.55, 273.65, 273.65, 273.55, 273.45, 273.25, 273.25, 
    273.05, 272.95, 272.85, 272.85, 272.65, 272.95, 273.15, 273.15, 272.95, 
    273.15, 272.95, 272.85, 272.85, 272.85, 272.95, 273.05, 272.85, 272.85, 
    273.15, 272.85, 272.75, 272.75, 272.85, 272.85, 272.75, 272.45, 272.25, 
    272.05, 271.65, 271.35, 271.85, 272.15, 272.05, 271.85, 271.65, 271.45, 
    270.75, 270.95, 271.45, 270.95, 270.45, 271.05, 270.65, 270.35, 269.95, 
    269.95, 269.65, 269.65, 269.05, 269.25, 268.85, 268.75, 268.95, 269.05, 
    269.05, 269.05, 268.95, 269.05, 268.75, 268.85, 268.85, 268.85, 268.95, 
    268.95, 269.05, 268.95, 269.05, 269.05, 269.05, 268.95, 268.85, 269.05, 
    268.85, 269.05, 268.95, 269.05, 268.95, 269.35, 269.25, 269.15, 269.35, 
    269.45, 269.55, 269.45, 269.45, 269.75, 269.85, 270.15, 270.25, 270.15, 
    270.05, 270.05, 270.35, 270.85, 271.55, 271.55, 271.35, 271.35, 271.15, 
    271.15, 271.05, 270.95, 270.95, 270.85, 270.75, 270.85, 271.05, 271.15, 
    271.35, 271.25, 271.25, 271.55, 271.55, 271.55, 271.45, 271.65, 271.35, 
    271.45, 271.55, 271.45, 271.45, 271.55, 271.45, 271.65, 271.35, 271.55, 
    271.45, 271.35, 271.35, 271.25, 271.25, 272.05, 272.05, 272.05, 272.05, 
    271.95, 272.05, 271.85, 271.65, 271.65, 271.05, 270.65, 270.65, 270.55, 
    270.15, 270.55, 269.75, 270.35, 270.45, 270.35, 270.35, 269.95, 270.15, 
    270.15, 269.85, 269.95, 269.45, 269.35, 269.25, 268.75, 268.85, 269.05, 
    268.75, 268.45, 268.45, 268.55, 267.65, 267.95, 268.15, 266.75, 267.45, 
    267.65, 268.25, 266.25, 266.75, 266.25, 266.55, 266.75, 265.95, 264.95, 
    266.55, 266.45, 266.75, 266.55, 265.45, 265.65, 264.75, 264.35, 264.35, 
    264.75, 264.85, 265.55, 265.35, 266.25, 266.55, 268.15, 268.15, 268.15, 
    268.55, 268.75, 268.55, 268.55, 268.75, 268.85, 269.05, 269.05, 269.35, 
    269.45, 269.65, 269.75, 269.85, 269.45, 270.45, 270.55, 270.55, 270.35, 
    270.05, 269.45, 269.75, 269.95, 269.75, 270.25, 269.75, 269.55, 269.15, 
    268.65, 268.45, 268.45, 268.55, 268.75, 268.55, 269.15, 268.85, 268.35, 
    270.85, 271.15, 271.35, 271.25, 270.05, 270.55, 270.65, 270.85, 269.75, 
    269.75, 270.05, 269.95, 270.25, 269.75, 269.65, 269.75, 269.25, 268.65, 
    268.65, 268.15, 268.25, 267.85, 268.05, 268.25, 268.15, 268.15, 268.45, 
    268.95, 269.45, 269.95, 269.65, 268.85, 267.95, 269.15, 270.25, 270.65, 
    270.55, 270.15, 270.05, 269.95, 270.05, 270.05, 269.65, 269.65, 268.95, 
    269.65, 269.95, 269.15, 268.75, 268.45, 267.55, 268.25, 268.25, 269.25, 
    269.05, 268.65, 269.35, 268.65, 268.85, 268.55, 268.35, 268.85, 269.45, 
    270.05, 270.35, 270.25, 270.35, 270.35, 270.15, 270.25, 270.15, 270.25, 
    270.15, 269.75, 270.05, 270.05, 270.35, 270.35, 270.35, 270.75, 270.85, 
    270.85, 270.75, 271.15, 270.85, 270.65, 270.25, 270.25, 270.55, 270.65, 
    271.05, 271.35, 271.45, 271.35, 271.05, 270.85, 270.65, 270.35, 269.95, 
    269.85, 269.85, 269.55, 269.65, 269.75, 269.75, 269.75, 269.65, 269.65, 
    269.65, 269.45, 269.15, 268.95, 268.85, 268.75, 269.25, 268.95, 268.85, 
    268.55, 268.55, 268.15, 267.65, 267.45, 267.35, 267.35, 266.95, 266.55, 
    266.25, 265.95, 265.65, 265.45, 265.45, 265.25, 265.25, 265.35, 265.45, 
    265.25, 265.25, 265.45, 265.45, 265.65, 266.25, 266.55, 266.95, 266.85, 
    266.95, 267.15, 267.55, 267.35, 268.25, 268.15, 267.15, 267.25, 266.35, 
    265.55, 265.25, 264.65, 264.15, 263.65, 261.65, 260.85, 259.55, 257.55, 
    256.05, 254.95, 254.25, 253.15, 252.65, 252.35, 252.65, 252.55, 252.55, 
    252.35, 252.05, 252.15, 252.25, 252.65, 252.55, 252.85, 253.05, 253.65, 
    254.25, 254.05, 253.75, 253.95, 253.85, 254.05, 253.85, 253.85, 254.25, 
    254.25, 254.45, 254.75, 254.85, 254.45, 254.55, 255.15, 255.75, 256.35, 
    256.65, 255.85, 255.25, 255.85, 256.85, 256.75, 256.55, 256.45, 256.25, 
    256.25, 256.45, 256.65, 256.65, 256.55, 256.35, 255.25, 254.85, 254.95, 
    255.25, 255.35, 255.95, 256.75, 256.95, 257.35, 259.15, 258.35, 257.95, 
    258.45, 258.25, 258.15, 258.55, 259.15, 260.15, 260.85, 260.95, 262.15, 
    264.05, 265.95, 267.05, 267.45, 268.05, 269.15, 269.25, 269.55, 269.95, 
    269.85, 270.25, 270.45, 270.95, 271.05, 271.35, 271.45, 270.05, 269.35, 
    268.75, 268.05, 268.05, 266.75, 264.55, 263.25, 262.55, 261.85, 261.45, 
    261.15, 260.75, 260.35, 259.25, 258.85, 258.45, 258.25, 258.05, 258.35, 
    257.85, 258.35, 258.75, 258.05, 257.95, 258.75, 258.25, 259.65, 260.85, 
    261.25, 262.45, 264.55, 264.85, 265.05, 265.35, 265.45, 265.65, 265.85, 
    266.15, 266.55, 266.55, 267.65, 268.95, 269.45, 270.15, 269.35, 268.95, 
    268.45, 267.25, 267.95, 267.75, 267.85, 268.75, 269.35, 268.95, 268.85, 
    268.65, 268.35, 268.45, 268.55, 268.75, 269.05, 268.75, 268.15, 269.05, 
    269.95, 270.15, 269.65, 270.35, 270.35, 270.45, 270.35, 269.95, 269.85, 
    270.05, 270.35, 270.65, 270.85, 271.05, 271.15, 271.45, 271.45, 271.55, 
    271.75, 272.25, 272.35, 271.85, 271.85, 271.85, 271.65, 271.65, 271.75, 
    271.85, 271.85, 271.85, 271.75, 271.85, 271.85, 271.85, 271.75, 271.65, 
    271.55, 271.55, 271.55, 271.65, 271.55, 271.45, 271.45, 271.55, 271.45, 
    271.55, 271.45, 271.45, 271.55, 271.45, 271.35, 271.25, 271.05, 271.05, 
    270.85, 270.65, 270.55, 270.65, 270.65, 270.45, 270.35, 269.85, 269.55, 
    269.25, 269.05, 269.05, 269.05, 268.85, 269.45, 269.95, 269.65, 269.35, 
    269.15, 269.05, 268.35, 268.05, 267.65, 267.35, 267.05, 266.45, 264.05, 
    264.75, 263.55, 265.15, 265.35, 264.95, 265.25, 264.85, 264.15, 263.45, 
    264.25, 265.55, 264.95, 263.75, 265.35, 264.75, 263.75, 264.85, 263.45, 
    263.35, 262.75, 262.15, 262.15, 262.15, 262.15, 262.55, 262.65, 262.55, 
    262.55, 262.35, 261.95, 262.65, 262.35, 261.55, 261.45, 261.35, 261.15, 
    261.35, 261.45, 261.15, 260.45, 259.75, 259.55, 259.65, 259.35, 259.45, 
    259.25, 258.75, 258.65, 258.45, 258.05, 258.65, 258.85, 259.55, 259.05, 
    258.35, 257.75, 258.95, 258.75, 258.85, 257.95, 258.05, 257.75, 257.55, 
    257.65, 257.85, 257.85, 257.75, 257.65, 257.45, 256.75, 256.55, 256.15, 
    256.45, 256.45, 256.35, 256.25, 256.05, 256.05, 256.05, 255.45, 255.15, 
    256.25, 256.05, 254.85, 254.55, 254.65, 254.25, 254.55, 255.75, 256.35, 
    256.75, 256.75, 257.05, 257.35, 258.35, 257.55, 258.25, 257.75, 257.65, 
    259.85, 259.95, 259.75, 260.25, 259.95, 260.05, 260.65, 260.25, 259.85, 
    258.85, 258.95, 256.55, 255.05, 255.35, 256.15, 255.35, 254.95, 254.15, 
    253.45, 252.75, 252.25, 251.95, 251.75, 251.65, 251.55, 251.65, 251.65, 
    251.75, 251.65, 251.65, 251.75, 251.45, 251.25, 251.35, 251.35, 251.15, 
    251.05, 250.95, 251.15, 251.15, 251.15, 250.95, 251.05, 251.05, 251.25, 
    251.45, 251.75, 251.95, 251.95, 252.15, 252.35, 252.45, 252.45, 252.05, 
    251.85, 251.65, 252.05, 252.35, 252.75, 253.15, 253.55, 253.75, 253.55, 
    252.35, 252.05, 251.75, 251.75, 251.75, 251.95, 252.45, 252.85, 253.35, 
    253.15, 253.95, 254.55, 254.85, 254.85, 255.05, 255.55, 256.45, 257.05, 
    257.15, 256.35, 256.35, 256.35, 256.25, 256.35, 256.45, 256.55, 256.85, 
    257.15, 257.35, 257.65, 257.45, 257.45, 257.45, 257.15, 257.35, 257.25, 
    257.05, 256.85, 257.05, 257.15, 257.05, 257.45, 257.95, 258.35, 259.15, 
    259.25, 258.85, 259.05, 259.15, 259.05, 258.95, 258.95, 259.55, 259.85, 
    259.75, 259.45, 259.05, 258.55, 258.75, 258.45, 258.35, 258.25, 258.15, 
    258.05, 258.55, 258.85, 258.65, 258.75, 258.65, 258.55, 258.45, 258.15, 
    257.95, 257.75, 257.65, 257.15, 257.15, 257.05, 256.55, 256.15, 256.05, 
    255.85, 256.55, 256.25, 256.55, 256.65, 256.75, 256.65, 256.65, 256.55, 
    256.05, 256.25, 255.85, 256.15, 257.05, 256.65, 256.25, 256.05, 255.95, 
    255.15, 256.85, 256.95, 256.75, 256.65, 256.25, 255.75, 255.05, 255.15, 
    255.45, 255.95, 256.45, 256.05, 256.25, 256.95, 257.25, 257.15, 256.85, 
    256.95, 256.95, 257.15, 257.05, 256.45, 257.15, 257.55, 256.15, 255.95, 
    255.35, 255.25, 255.15, 254.85, 254.75, 253.95, 253.95, 253.35, 253.35, 
    254.25, 253.65, 254.05, 253.55, 255.15, 255.35, 256.45, 256.55, 256.95, 
    257.15, 257.65, 257.55, 257.65, 257.35, 255.85, 256.45, 256.85, 256.35, 
    255.75, 255.35, 255.35, 256.05, 255.55, 255.15, 255.35, 254.45, 254.15, 
    253.55, 253.05, 252.55, 252.65, 252.85, 254.45, 254.45, 254.65, 254.75, 
    255.05, 255.65, 255.65, 255.65, 255.85, 255.95, 256.25, 256.35, 256.75, 
    256.85, 257.15, 257.45, 257.65, 257.75, 257.95, 258.25, 258.85, 259.25, 
    259.55, 259.85, 259.85, 259.85, 260.15, 260.35, 260.75, 260.85, 260.75, 
    260.55, 260.35, 260.25, 260.25, 260.25, 260.65, 260.45, 260.55, 259.25, 
    258.35, 258.15, 256.85, 255.45, 255.05, 254.45, 256.15, 255.85, 255.85, 
    256.35, 256.55, 257.05, 258.05, 258.05, 257.25, 257.05, 257.15, 256.85, 
    255.55, 256.95, 258.75, 258.45, 258.05, 257.35, 256.95, 256.45, 256.85, 
    256.75, 256.75, 256.65, 256.55, 256.75, 256.85, 256.95, 257.15, 257.05, 
    257.55, 257.05, 256.95, 255.55, 255.05, 256.05, 256.55, 256.25, 255.75, 
    255.75, 256.65, 257.05, 257.95, 258.25, 259.05, 259.85, 258.85, 260.45, 
    260.65, 261.35, 262.05, 262.15, 261.75, 261.25, 261.25, 261.15, 261.85, 
    262.45, 263.05, 262.85, 262.85, 263.25, 264.35, 265.35, 266.05, 267.05, 
    267.95, 268.95, 269.25, 267.55, 267.55, 268.35, 269.45, 268.85, 267.85, 
    267.55, 267.45, 267.55, 267.15, 266.75, 266.95, 267.45, 266.35, 264.75, 
    263.05, 263.15, 263.95, 263.95, 262.95, 261.35, 259.65, 258.25, 257.75, 
    257.35, 256.65, 256.65, 256.95, 256.75, 257.25, 258.95, 259.65, 260.55, 
    260.55, 260.25, 260.45, 260.15, 259.25, 258.35, 258.25, 258.15, 258.05, 
    258.25, 258.15, 258.25, 258.65, 259.25, 259.45, 259.15, 259.45, 259.55, 
    259.45, 260.15, 260.35, 260.75, 260.05, 259.95, 257.95, 256.05, 254.25, 
    253.65, 253.75, 253.95, 253.95, 253.65, 253.65, 253.65, 253.75, 254.05, 
    253.55, 253.85, 253.85, 254.05, 254.35, 254.45, 254.35, 253.85, 254.05, 
    253.85, 253.55, 253.25, 252.95, 252.95, 253.35, 253.55, 253.75, 253.75, 
    253.85, 253.55, 253.55, 253.35, 253.05, 253.35, 253.85, 253.35, 253.15, 
    253.55, 253.85, 254.15, 254.85, 255.35, 255.55, 255.85, 255.85, 255.85, 
    255.65, 255.45, 255.35, 255.35, 253.85, 253.25, 253.05, 252.85, 252.55, 
    252.25, 251.95, 251.65, 251.55, 251.55, 251.55, 251.55, 251.55, 251.85, 
    252.35, 252.25, 252.55, 252.85, 252.95, 252.95, 253.05, 253.15, 252.75, 
    252.55, 252.55, 252.35, 252.25, 252.45, 252.65, 252.85, 253.75, 254.75, 
    255.35, 255.75, 255.95, 255.85, 256.45, 256.35, 256.25, 257.05, 257.25, 
    257.95, 258.55, 258.15, 258.25, 258.45, 258.95, 257.85, 257.95, 257.95, 
    258.05, 256.75, 256.55, 256.65, 256.85, 256.85, 256.85, 257.15, 257.25, 
    257.25, 257.35, 257.45, 257.55, 257.85, 258.05, 258.25, 258.15, 257.95, 
    258.25, 257.55, 257.15, 256.75, 257.55, 257.95, 258.05, 257.75, 258.25, 
    257.95, 256.95, 255.85, 256.45, 256.95, 256.35, 256.65, 255.45, 254.85, 
    255.05, 255.35, 255.45, 255.25, 255.15, 255.05, 255.75, 255.35, 255.55, 
    254.85, 255.75, 255.75, 255.75, 254.95, 255.05, 255.45, 255.65, 256.75, 
    257.25, 256.75, 256.65, 256.55, 256.65, 256.15, 256.15, 256.25, 255.95, 
    255.85, 256.05, 255.95, 255.85, 255.95, 255.85, 255.55, 254.45, 253.35, 
    252.25, 251.85, 251.65, 250.95, 251.05, 250.75, 250.55, 250.05, 250.25, 
    250.75, 251.45, 252.35, 253.05, 253.45, 253.35, 252.85, 252.65, 252.45, 
    252.35, 252.05, 251.85, 251.85, 250.85, 250.45, 250.05, 250.35, 250.55, 
    250.25, 250.35, 250.25, 249.95, 249.75, 249.25, 249.25, 249.35, 251.15, 
    251.25, 252.05, 253.45, 254.15, 255.05, 255.95, 256.65, 257.55, 258.45, 
    258.75, 258.85, 258.75, 260.65, 261.15, 261.35, 261.75, 262.05, 262.25, 
    262.55, 262.85, 263.25, 263.65, 264.35, 266.15, 263.35, 261.95, 261.25, 
    260.85, 260.85, 260.45, 260.75, 260.55, 260.55, 260.85, 261.45, 261.55, 
    259.35, 259.65, 260.05, 260.55, 259.95, 260.55, 261.65, 261.05, 261.55, 
    261.75, 262.95, 264.15, 265.95, 266.25, 267.15, 267.75, 267.55, 264.45, 
    264.25, 261.25, 262.05, 261.15, 260.45, 259.55, 257.35, 256.15, 255.25, 
    253.35, 252.15, 250.85, 250.35, 249.85, 250.55, 250.75, 252.55, 253.75, 
    253.25, 253.65, 253.05, 253.35, 254.55, 254.95, 255.15, 255.45, 256.15, 
    256.25, 256.15, 256.15, 255.95, 256.05, 256.45, 256.45, 256.15, 255.15, 
    254.65, 253.75, 253.55, 254.45, 254.05, 253.75, 253.25, 253.35, 253.15, 
    253.45, 252.75, 252.25, 251.85, 251.55, 251.35, 250.85, 250.25, 250.05, 
    250.15, 249.65, 249.35, 248.65, 248.65, 248.35, 249.85, 249.75, 249.55, 
    249.35, 248.15, 248.05, 247.95, 248.05, 248.65, 248.95, 248.95, 249.35, 
    249.55, 249.55, 250.05, 249.55, 249.95, 250.15, 249.95, 250.35, 250.05, 
    250.35, 250.25, 249.85, 249.85, 249.45, 248.65, 250.35, 250.35, 251.55, 
    252.35, 254.05, 254.85, 255.35, 255.95, 256.35, 256.85, 257.15, 258.55, 
    257.85, 257.45, 257.15, 256.95, 257.25, 255.95, 255.65, 254.95, 254.75, 
    254.45, 255.85, 254.65, 257.05, 257.75, 258.45, 259.35, 259.95, 260.75, 
    261.65, 261.65, 262.35, 262.55, 262.95, 263.15, 263.35, 262.55, 262.85, 
    262.25, 262.95, 263.15, 262.35, 262.85, 261.15, 262.25, 261.35, 263.35, 
    262.35, 262.45, 263.65, 264.15, 264.75, 265.45, 266.25, 266.85, 266.95, 
    267.05, 267.15, 267.35, 267.75, 269.15, 269.95, 270.15, 270.85, 270.95, 
    270.85, 270.85, 270.65, 270.55, 270.65, 270.75, 270.75, 270.85, 271.25, 
    271.45, 272.55, 272.45, 272.45, 271.85, 271.55, 271.45, 270.75, 267.55, 
    262.65, 261.45, 259.75, 259.35, 258.35, 258.25, 257.45, 256.35, 255.55, 
    254.75, 254.95, 254.75, 254.65, 254.85, 254.95, 255.35, 255.35, 255.15, 
    255.45, 255.65, 255.45, 255.95, 256.05, 255.75, 255.95, 255.85, 256.15, 
    255.95, 255.35, 255.25, 254.95, 255.15, 254.95, 255.25, 255.35, 255.25, 
    255.05, 254.95, 254.95, 255.15, 255.65, 256.05, 256.35, 256.35, 256.05, 
    256.45, 256.75, 257.15, 257.95, 258.15, 257.65, 258.15, 258.35, 258.15, 
    257.85, 257.65, 256.45, 256.95, 256.85, 256.85, 256.85, 256.65, 256.75, 
    257.55, 258.75, 259.45, 259.85, 260.15, 260.05, 260.35, 259.95, 259.75, 
    259.45, 259.55, 259.85, 259.75, 258.85, 258.35, 256.35, 257.15, 256.95, 
    257.75, 258.25, 259.05, 259.15, 260.35, 261.05, 261.25, 261.25, 260.65, 
    260.45, 260.25, 259.65, 259.05, 257.55, 256.95, 257.25, 256.85, 256.65, 
    256.95, 256.95, 256.95, 257.15, 257.15, 257.35, 257.15, 257.05, 257.05, 
    257.45, 257.15, 257.15, 257.05, 257.05, 257.25, 257.05, 257.05, 258.05, 
    258.25, 258.35, 257.65, 257.55, 257.45, 257.75, 257.95, 257.75, 257.75, 
    257.55, 257.35, 257.35, 257.25, 257.45, 257.45, 256.75, 257.05, 257.45, 
    257.85, 258.05, 257.95, 257.35, 257.55, 257.85, 257.75, 257.55, 257.45, 
    257.35, 257.05, 256.95, 257.35, 256.85, 255.95, 255.25, 255.15, 254.95, 
    255.05, 255.65, 256.25, 256.15, 256.55, 257.15, 257.55, 258.05, 258.45, 
    258.25, 258.95, 258.65, 258.75, 258.85, 258.95, 259.15, 259.15, 258.85, 
    258.15, 257.95, 257.85, 257.45, 257.75, 257.75, 257.45, 257.45, 257.45, 
    257.75, 258.05, 257.95, 258.15, 258.05, 258.25, 258.35, 258.05, 258.65, 
    258.85, 258.55, 258.65, 258.85, 259.05, 259.05, 259.15, 259.15, 259.05, 
    258.85, 258.55, 257.95, 257.65, 257.55, 257.65, 257.85, 258.15, 258.65, 
    258.65, 258.85, 258.95, 258.95, 258.85, 258.75, 258.75, 258.85, 258.95, 
    258.95, 259.05, 259.15, 259.45, 259.45, 259.55, 259.45, 259.55, 259.85, 
    260.15, 260.15, 260.65, 261.05, 261.25, 261.65, 262.05, 262.45, 262.45, 
    262.55, 262.35, 260.45, 261.15, 260.95, 261.65, 262.25, 261.55, 260.25, 
    260.85, 261.65, 263.25, 262.75, 262.35, 262.15, 262.65, 263.25, 263.45, 
    263.55, 263.35, 263.85, 264.05, 263.95, 263.75, 263.35, 263.05, 262.95, 
    263.15, 262.85, 262.45, 262.75, 261.85, 261.75, 261.15, 259.95, 259.55, 
    260.05, 260.35, 260.55, 260.95, 261.25, 261.55, 261.95, 262.45, 262.85, 
    263.25, 263.35, 263.65, 264.25, 264.65, 265.05, 265.15, 265.05, 264.95, 
    264.75, 264.45, 264.15, 264.05, 263.85, 264.55, 265.05, 265.15, 265.05, 
    265.05, 265.05, 265.15, 265.15, 265.25, 265.35, 265.35, 265.55, 265.75, 
    265.15, 265.55, 265.95, 265.85, 265.65, 265.45, 265.05, 264.85, 264.95, 
    264.55, 264.55, 264.65, 264.65, 264.75, 264.55, 264.55, 264.45, 264.85, 
    264.55, 264.45, 264.65, 264.65, 264.85, 264.95, 265.35, 265.35, 265.55, 
    265.45, 265.05, 265.05, 264.65, 264.45, 264.75, 264.95, 264.85, 264.75, 
    264.95, 264.95, 264.65, 265.15, 264.85, 264.75, 264.75, 264.75, 264.45, 
    263.95, 263.65, 263.25, 263.65, 264.05, 263.75, 263.45, 263.35, 262.85, 
    262.35, 262.15, 262.25, 261.95, 261.85, 261.55, 261.55, 261.45, 261.85, 
    261.85, 261.65, 261.15, 260.35, 259.35, 258.95, 258.65, 258.65, 258.75, 
    259.15, 259.55, 260.15, 260.45, 260.45, 260.35, 260.55, 260.95, 261.05, 
    260.15, 259.75, 259.55, 259.75, 259.55, 259.35, 259.65, 259.45, 259.25, 
    259.15, 259.55, 260.05, 259.65, 259.55, 259.25, 260.05, 260.25, 259.65, 
    259.75, 260.05, 259.75, 259.85, 259.95, 260.35, 260.95, 261.15, 261.35, 
    261.35, 261.65, 262.25, 262.85, 263.45, 263.95, 264.35, 264.85, 264.45, 
    265.65, 266.85, 267.15, 267.55, 268.25, 268.25, 267.95, 267.75, 267.35, 
    267.35, 266.85, 266.15, 265.85, 265.35, 265.15, 264.35, 264.05, 265.05, 
    265.15, 265.25, 265.25, 266.05, 266.75, 267.35, 267.45, 268.55, 268.75, 
    268.35, 268.85, 269.05, 269.05, 269.15, 269.45, 268.95, 269.75, 269.05, 
    269.75, 270.65, 270.65, 271.25, 271.85, 272.25, 270.35, 272.05, 271.75, 
    270.35, 271.85, 272.65, 272.95, 272.75, 271.45, 271.05, 271.35, 271.45, 
    271.45, 271.65, 271.05, 270.95, 270.95, 270.95, 270.65, 269.95, 269.75, 
    270.05, 270.45, 270.75, 270.95, 271.75, 269.25, 266.65, 265.15, 264.85, 
    264.85, 264.95, 265.25, 265.65, 265.65, 266.05, 266.25, 266.25, 266.15, 
    265.95, 265.85, 265.65, 265.55, 265.45, 265.45, 264.95, 264.75, 264.95, 
    264.95, 264.85, 265.45, 265.75, 266.25, 265.95, 266.05, 266.65, 266.75, 
    267.35, 267.65, 267.15, 267.15, 267.45, 266.55, 266.25, 265.75, 265.55, 
    265.05, 264.95, 264.65, 264.65, 264.65, 264.15, 264.15, 264.35, 263.75, 
    263.35, 263.25, 263.95, 264.55, 264.55, 264.75, 265.15, 263.65, 263.35, 
    263.25, 262.95, 262.65, 262.55, 262.85, 262.85, 262.55, 262.05, 262.05, 
    262.85, 262.95, 262.85, 262.95, 262.95, 262.65, 262.65, 262.85, 263.25, 
    263.55, 264.05, 264.55, 264.45, 264.25, 263.75, 263.65, 263.25, 263.15, 
    263.15, 263.05, 262.95, 261.85, 262.85, 263.25, 263.45, 263.05, 262.85, 
    262.75, 262.45, 262.85, 263.25, 264.55, 265.25, 265.25, 265.55, 265.25, 
    264.95, 264.25, 263.65, 263.35, 263.15, 262.95, 262.95, 262.95, 262.85, 
    262.95, 263.45, 263.35, 263.45, 263.75, 263.95, 263.05, 262.55, 262.75, 
    263.35, 263.15, 262.95, 263.75, 263.45, 263.45, 264.05, 264.15, 264.35, 
    263.85, 263.85, 263.85, 263.45, 262.95, 262.45, 262.45, 261.65, 261.05, 
    260.85, 260.85, 260.85, 261.05, 262.15, 262.75, 263.15, 263.45, 262.95, 
    264.25, 264.05, 264.25, 264.35, 264.85, 264.15, 263.35, 263.35, 262.85, 
    262.75, 263.25, 262.35, 262.05, 261.45, 261.05, 260.75, 260.35, 260.35, 
    260.95, 260.95, 260.75, 260.35, 260.55, 260.75, 260.85, 261.25, 261.45, 
    261.65, 261.75, 261.95, 262.15, 261.65, 261.55, 262.25, 262.65, 262.95, 
    263.15, 263.35, 263.35, 262.95, 263.25, 263.05, 263.75, 264.05, 264.25, 
    264.65, 265.15, 265.95, 266.95, 268.15, 268.65, 268.95, 269.25, 269.15, 
    269.35, 269.65, 269.95, 269.25, 269.35, 269.55, 270.45, 270.95, 271.25, 
    271.25, 271.75, 271.95, 272.25, 272.75, 272.85, 272.85, 272.55, 272.85, 
    272.75, 272.65, 272.65, 272.95, 273.25, 272.05, 270.65, 269.75, 268.85, 
    267.85, 267.35, 266.25, 265.55, 264.95, 264.25, 264.15, 263.75, 263.25, 
    262.75, 262.75, 262.65, 262.55, 262.65, 262.75, 263.05, 263.45, 263.75, 
    263.75, 264.05, 264.25, 264.05, 264.45, 264.55, 264.55, 264.45, 264.35, 
    264.35, 264.25, 264.15, 264.55, 264.95, 264.65, 265.15, 266.25, 266.25, 
    266.35, 266.55, 266.05, 265.25, 264.55, 264.25, 264.55, 266.35, 264.95, 
    267.75, 267.55, 267.35, 267.65, 269.05, 268.85, 268.65, 268.55, 268.65, 
    268.65, 267.25, 268.05, 267.05, 266.35, 266.35, 265.95, 265.05, 264.85, 
    264.65, 264.65, 265.05, 265.15, 265.45, 265.95, 266.15, 266.35, 266.55, 
    266.35, 266.25, 266.55, 266.85, 267.15, 265.95, 265.55, 265.85, 265.75, 
    265.85, 265.95, 265.95, 266.25, 266.55, 267.05, 266.55, 266.05, 266.25, 
    265.75, 265.55, 265.65, 265.75, 265.95, 266.15, 265.85, 265.45, 265.05, 
    265.15, 265.45, 265.65, 265.85, 265.55, 266.05, 266.55, 266.25, 266.45, 
    266.55, 266.35, 266.55, 267.05, 266.45, 266.95, 267.05, 267.25, 267.25, 
    267.75, 267.55, 267.35, 267.25, 266.95, 266.65, 267.45, 267.15, 267.05, 
    266.75, 266.55, 266.65, 266.35, 267.05, 267.45, 268.15, 268.15, 268.15, 
    268.45, 268.75, 268.55, 268.75, 268.45, 268.15, 267.55, 267.35, 267.05, 
    266.85, 266.85, 266.85, 266.95, 266.75, 265.65, 265.25, 264.85, 265.35, 
    264.85, 264.25, 264.25, 263.85, 263.95, 263.85, 264.45, 265.25, 265.75, 
    266.15, 266.65, 266.25, 266.25, 266.25, 266.25, 266.15, 266.15, 266.05, 
    266.05, 266.05, 266.05, 265.85, 265.75, 265.85, 265.95, 266.05, 266.25, 
    266.35, 266.25, 266.35, 266.45, 266.95, 266.95, 267.05, 267.25, 267.25, 
    267.25, 267.15, 266.95, 266.65, 266.65, 266.65, 266.55, 266.45, 266.15, 
    265.85, 265.55, 264.65, 264.15, 263.45, 263.25, 263.95, 264.65, 265.15, 
    265.55, 266.15, 266.45, 266.45, 266.35, 266.15, 266.25, 266.55, 266.55, 
    266.65, 267.05, 267.55, 267.95, 268.15, 268.75, 269.55, 269.25, 269.45, 
    269.75, 269.65, 269.45, 269.65, 270.15, 270.15, 269.85, 269.55, 269.25, 
    269.55, 269.55, 270.05, 271.05, 271.85, 272.65, 273.55, 272.85, 272.75, 
    272.65, 272.65, 272.45, 273.05, 272.95, 271.75, 272.95, 272.85, 273.45, 
    273.45, 273.25, 273.15, 272.85, 273.25, 272.85, 272.15, 271.55, 271.15, 
    271.25, 271.15, 271.15, 271.65, 271.25, 270.95, 271.15, 270.75, 270.85, 
    271.05, 271.15, 271.15, 271.85, 272.75, 271.45, 271.75, 272.15, 272.45, 
    272.95, 273.35, 274.55, 273.95, 274.25, 274.75, 275.85, 273.75, 274.05, 
    273.45, 273.35, 273.45, 273.45, 273.45, 273.85, 272.85, 272.65, 273.65, 
    274.45, 273.35, 273.55, 273.85, 273.45, 274.15, 273.35, 275.25, 273.95, 
    273.45, 273.65, 273.25, 272.95, 272.75, 272.65, 272.75, 272.55, 272.15, 
    272.65, 272.05, 272.05, 271.95, 271.45, 271.25, 271.15, 271.25, 271.15, 
    271.35, 271.15, 269.95, 270.15, 269.95, 269.65, 269.55, 268.95, 269.65, 
    269.65, 269.55, 270.25, 270.45, 270.75, 270.55, 270.45, 269.85, 269.75, 
    269.65, 269.55, 269.75, 269.65, 269.65, 269.75, 270.05, 270.15, 270.05, 
    269.95, 269.75, 269.85, 270.25, 269.95, 270.25, 270.35, 270.45, 270.65, 
    270.55, 269.95, 268.65, 269.05, 268.45, 268.35, 268.25, 268.15, 267.75, 
    267.65, 267.65, 267.25, 267.25, 267.25, 267.15, 267.15, 268.15, 269.55, 
    270.85, 269.75, 269.75, 270.45, 271.15, 271.45, 271.35, 271.25, 271.45, 
    271.75, 271.85, 271.85, 271.95, 272.05, 272.05, 272.15, 272.35, 272.75, 
    272.55, 272.85, 271.75, 270.55, 271.45, 271.25, 270.95, 270.65, 270.55, 
    270.65, 270.55, 270.75, 270.55, 270.65, 270.65, 270.55, 270.05, 269.55, 
    268.95, 268.75, 268.45, 269.25, 269.45, 269.35, 268.95, 268.45, 268.15, 
    268.65, 268.95, 269.55, 269.25, 269.55, 270.25, 272.55, 271.85, 270.65, 
    269.75, 269.35, 269.75, 269.45, 269.25, 269.15, 269.15, 269.25, 270.35, 
    271.05, 271.65, 271.85, 272.05, 272.05, 271.95, 271.85, 271.65, 271.65, 
    271.75, 271.75, 271.75, 271.85, 271.95, 272.05, 272.05, 272.15, 272.35, 
    272.45, 272.45, 272.45, 272.45, 272.45, 272.55, 272.65, 272.75, 272.95, 
    273.05, 273.35, 273.95, 274.45, 274.25, 273.25, 273.15, 273.05, 273.05, 
    273.15, 273.15, 273.15, 272.55, 272.25, 271.65, 271.25, 270.95, 270.85, 
    269.55, 269.45, 269.55, 270.35, 271.25, 271.45, 272.25, 273.75, 272.55, 
    272.65, 273.55, 272.55, 272.35, 272.05, 271.95, 271.45, 271.15, 270.95, 
    270.75, 270.75, 271.35, 271.45, 271.55, 272.05, 272.45, 272.65, 272.65, 
    272.85, 272.85, 273.05, 273.05, 273.05, 273.05, 273.15, 273.25, 273.25, 
    273.35, 273.35, 273.15, 272.75, 272.65, 272.75, 272.25, 272.65, 272.65, 
    272.45, 272.75, 273.25, 273.15, 272.85, 272.75, 272.95, 273.05, 273.15, 
    272.85, 272.55, 272.15, 271.65, 271.25, 270.85, 270.75, 270.35, 270.45, 
    270.05, 270.55, 270.65, 270.55, 270.55, 270.75, 270.85, 270.95, 271.05, 
    270.85, 270.85, 271.25, 271.25, 271.25, 271.35, 271.25, 271.35, 271.45, 
    271.55, 271.55, 271.45, 271.95, 271.65, 271.95, 272.05, 271.95, 272.15, 
    272.35, 272.25, 272.15, 271.75, 272.25, 271.35, 271.35, 271.15, 270.75, 
    270.75, 270.75, 270.35, 270.45, 270.35, 270.85, 270.05, 269.55, 269.45, 
    269.55, 269.45, 269.65, 269.85, 270.15, 270.25, 270.15, 271.35, 271.45, 
    270.95, 270.55, 270.55, 270.65, 270.35, 270.95, 270.75, 270.85, 271.45, 
    271.65, 270.75, 270.05, 269.75, 270.15, 270.25, 269.95, 269.75, 269.25, 
    269.05, 269.55, 269.35, 269.25, 269.05, 268.65, 268.45, 268.15, 268.55, 
    268.65, 268.95, 269.65, 269.95, 270.05, 270.15, 270.45, 270.75, 271.25, 
    271.45, 271.85, 272.75, 273.05, 274.25, 274.05, 273.25, 272.95, 273.05, 
    272.85, 272.65, 272.45, 272.25, 272.05, 271.85, 271.75, 270.35, 269.95, 
    269.05, 268.85, 268.85, 268.85, 268.95, 269.25, 269.25, 269.25, 268.35, 
    268.15, 268.45, 268.45, 268.55, 268.95, 269.25, 269.35, 269.15, 268.95, 
    269.05, 270.15, 268.75, 268.85, 267.35, 268.05, 269.65, 268.45, 268.15, 
    268.65, 268.85, 268.55, 268.55, 269.35, 272.45, 272.25, 272.65, 273.15, 
    272.95, 272.75, 272.65, 272.85, 272.45, 272.05, 272.15, 272.55, 272.55, 
    272.55, 272.55, 271.45, 272.15, 270.65, 271.85, 272.95, 272.15, 272.05, 
    272.45, 272.25, 272.05, 272.05, 272.45, 272.55, 272.45, 272.25, 272.35, 
    272.05, 272.25, 271.75, 271.65, 271.65, 271.15, 271.35, 271.45, 271.45, 
    271.65, 271.65, 271.85, 272.05, 272.25, 272.45, 272.55, 272.15, 272.35, 
    272.45, 272.25, 272.35, 272.25, 271.85, 271.35, 271.35, 271.45, 271.25, 
    270.75, 270.15, 269.95, 269.65, 269.05, 269.15, 269.65, 269.75, 269.75, 
    269.85, 269.65, 269.55, 269.55, 269.75, 269.85, 270.05, 270.15, 270.05, 
    270.05, 269.95, 269.95, 270.05, 269.95, 269.35, 269.05, 269.15, 268.95, 
    269.05, 268.95, 269.05, 269.15, 269.15, 269.15, 269.25, 269.55, 269.75, 
    269.75, 269.95, 270.15, 270.15, 270.25, 270.45, 270.45, 270.45, 270.55, 
    270.65, 270.35, 270.25, 270.35, 270.65, 270.45, 270.75, 270.75, 270.45, 
    270.55, 270.35, 270.75, 271.55, 271.75, 271.55, 272.25, 272.15, 271.85, 
    271.65, 271.55, 271.45, 271.85, 271.65, 271.65, 271.65, 271.95, 271.85, 
    271.75, 271.35, 271.25, 271.15, 271.45, 271.25, 270.85, 270.45, 270.65, 
    271.05, 271.35, 271.15, 271.05, 270.75, 271.25, 271.45, 271.65, 271.35, 
    271.25, 271.35, 271.25, 271.25, 270.95, 270.55, 270.25, 270.15, 270.05, 
    269.85, 269.55, 269.65, 269.35, 269.15, 269.15, 269.05, 268.95, 268.95, 
    269.35, 269.55, 269.55, 269.65, 269.85, 270.05, 269.85, 270.25, 270.75, 
    270.75, 271.25, 271.45, 271.55, 271.85, 271.75, 271.75, 271.85, 271.95, 
    272.15, 272.05, 272.15, 272.25, 271.95, 272.25, 272.25, 272.05, 272.35, 
    272.55, 272.55, 272.45, 272.45, 272.35, 271.65, 271.85, 271.35, 271.25, 
    271.25, 270.75, 269.95, 269.55, 268.75, 268.45, 268.55, 268.75, 268.25, 
    268.75, 268.55, 269.75, 270.35, 270.65, 270.65, 270.75, 271.25, 271.35, 
    272.15, 272.15, 272.75, 274.15, 273.35, 273.45, 273.35, 273.35, 273.45, 
    273.55, 273.55, 273.45, 273.55, 273.45, 273.55, 273.55, 273.65, 273.45, 
    273.55, 273.65, 273.85, 273.65, 273.85, 273.95, 274.45, 274.75, 274.05, 
    274.35, 274.45, 275.45, 275.15, 275.35, 275.55, 274.95, 275.15, 275.65, 
    274.35, 275.45, 274.55, 274.25, 275.45, 275.35, 274.75, 274.35, 275.15, 
    275.35, 274.85, 274.65, 274.45, 274.05, 273.65, 273.45, 273.25, 273.15, 
    273.05, 273.15, 273.45, 273.15, 273.35, 273.25, 272.85, 272.55, 272.85, 
    272.85, 272.35, 272.85, 272.55, 272.95, 272.45, 272.35, 272.25, 272.55, 
    272.45, 272.35, 272.25, 272.25, 271.95, 272.05, 271.85, 271.95, 272.05, 
    272.05, 271.75, 271.85, 271.85, 272.05, 272.35, 272.35, 272.25, 272.15, 
    272.55, 272.65, 272.75, 272.95, 273.05, 273.25, 273.25, 273.25, 272.95, 
    272.85, 272.85, 272.85, 272.65, 272.65, 272.55, 272.25, 272.15, 271.85, 
    271.95, 272.25, 272.65, 273.05, 272.85, 272.95, 273.05, 272.95, 272.95, 
    273.05, 273.15, 273.05, 273.15, 272.85, 272.85, 272.85, 272.65, 272.55, 
    272.05, 272.05, 272.35, 272.35, 272.35, 272.75, 272.75, 272.55, 272.65, 
    272.85, 272.75, 273.05, 273.05, 273.35, 273.85, 273.55, 273.85, 273.95, 
    274.55, 274.25, 274.35, 274.15, 273.95, 273.95, 274.05, 274.25, 274.15, 
    274.25, 274.15, 273.95, 273.75, 273.65, 273.55, 273.55, 273.45, 273.55, 
    273.55, 273.45, 273.45, 273.35, 273.45, 273.45, 273.35, 273.35, 273.25, 
    273.15, 273.15, 273.15, 273.15, 273.25, 273.25, 273.35, 273.35, 273.55, 
    274.15, 274.55, 273.45, 273.95, 273.75, 273.85, 274.25, 274.25, 274.45, 
    274.45, 275.15, 274.35, 273.85, 274.45, 273.95, 273.15, 272.35, 272.55, 
    272.55, 272.05, 272.35, 272.05, 271.45, 271.15, 271.15, 271.35, 272.15, 
    273.05, 272.05, 272.85, 274.15, 274.15, 273.85, 273.25, 273.25, 273.55, 
    273.35, 273.15, 273.15, 273.65, 274.35, 275.15, 273.35, 273.35, 273.75, 
    273.45, 273.45, 273.45, 273.35, 273.45, 273.35, 273.45, 273.25, 273.35, 
    273.35, 273.45, 273.75, 273.55, 273.55, 273.25, 273.25, 273.25, 273.35, 
    273.15, 273.05, 273.05, 272.85, 272.35, 271.45, 271.65, 271.65, 271.85, 
    272.15, 272.25, 272.55, 272.75, 272.85, 272.85, 273.05, 272.95, 272.75, 
    272.95, 273.15, 272.65, 272.85, 272.85, 272.95, 272.65, 272.75, 273.05, 
    272.25, 272.75, 271.25, 271.65, 271.65, 272.05, 272.95, 273.35, 273.95, 
    274.55, 274.65, 275.15, 274.55, 274.55, 275.05, 274.55, 274.25, 273.95, 
    274.05, 273.35, 273.15, 273.65, 274.05, 274.15, 273.65, 273.65, 274.15, 
    275.15, 274.55, 274.05, 273.35, 273.25, 272.85, 272.75, 272.85, 272.55, 
    273.15, 273.15, 273.55, 273.75, 273.85, 273.35, 272.75, 273.75, 273.35, 
    272.85, 272.85, 272.75, 272.55, 272.45, 272.45, 272.25, 272.15, 272.25, 
    272.45, 272.45, 272.55, 272.55, 272.45, 272.35, 272.35, 272.35, 272.35, 
    272.75, 273.75, 274.15, 273.85, 273.85, 273.25, 272.45, 271.85, 272.15, 
    271.65, 271.75, 272.35, 273.95, 273.95, 275.15, 275.45, 275.05, 274.95, 
    274.65, 274.65, 274.65, 274.65, 274.95, 274.95, 274.95, 275.55, 276.15, 
    275.95, 276.15, 276.85, 275.35, 275.05, 275.55, 275.25, 274.75, 273.75, 
    274.45, 275.55, 276.15, 279.05, 277.95, 279.45, 279.25, 279.45, 278.45, 
    277.45, 278.65, 275.75, 276.25, 275.75, 278.55, 278.85, 277.15, 276.55, 
    276.15, 275.95, 275.25, 275.15, 275.05, 274.65, 273.75, 273.55, 273.65, 
    273.35, 273.65, 273.55, 273.75, 273.65, 273.55, 273.85, 273.75, 273.75, 
    273.85, 274.15, 274.15, 273.95, 274.55, 274.55, 274.75, 275.45, 275.35, 
    276.65, 275.35, 274.95, 274.65, 274.85, 276.55, 274.05, 274.05, 274.45, 
    274.35, 273.95, 273.45, 273.35, 273.35, 273.35, 273.35, 273.25, 273.05, 
    273.15, 272.95, 272.95, 273.05, 273.05, 273.05, 273.05, 273.05, 273.05, 
    273.05, 273.15, 272.95, 272.95, 273.05, 273.05, 273.05, 273.15, 273.25, 
    273.25, 273.35, 273.35, 273.25, 273.35, 273.25, 273.25, 273.05, 273.15, 
    273.15, 273.15, 273.15, 273.15, 273.25, 273.25, 273.15, 273.05, 273.05, 
    272.95, 272.95, 273.05, 272.95, 273.05, 273.15, 273.15, 273.25, 273.35, 
    273.35, 273.35, 273.25, 273.35, 273.25, 273.25, 273.15, 273.15, 273.05, 
    273.05, 272.85, 272.85, 272.85, 272.95, 273.15, 273.15, 273.15, 273.25, 
    273.35, 273.45, 273.45, 273.25, 273.05, 273.25, 273.55, 273.55, 273.55, 
    273.55, 273.65, 273.65, 273.55, 273.55, 273.35, 272.55, 273.75, 273.95, 
    274.15, 274.25, 274.65, 274.55, 274.75, 275.75, 275.45, 275.45, 275.55, 
    275.65, 274.75, 274.05, 273.65, 273.45, 273.95, 273.85, 274.15, 274.35, 
    274.15, 274.15, 274.55, 274.55, 274.55, 274.45, 274.45, 274.25, 274.15, 
    274.25, 274.25, 273.95, 274.35, 274.65, 274.75, 274.45, 274.55, 274.55, 
    274.55, 274.55, 274.65, 274.65, 275.35, 274.75, 274.45, 275.25, 273.75, 
    274.45, 274.05, 273.75, 273.45, 274.05, 274.55, 273.65, 273.75, 273.75, 
    273.75, 273.75, 275.95, 273.75, 274.05, 275.05, 274.85, 274.75, 274.45, 
    274.45, 275.35, 275.75, 276.15, 276.05, 276.05, 276.95, 276.05, 276.35, 
    276.15, 275.75, 276.15, 276.45, 275.65, 275.45, 274.95, 274.85, 274.15, 
    273.75, 274.85, 274.65, 274.25, 276.15, 275.25, 275.65, 274.05, 273.65, 
    273.55, 275.45, 276.45, 276.95, 276.55, 276.65, 276.25, 276.05, 275.95, 
    276.45, 276.25, 276.65, 275.85, 276.35, 277.05, 277.05, 275.05, 275.95, 
    276.65, 276.15, 276.65, 276.55, 276.55, 276.55, 275.25, 275.35, 275.95, 
    276.05, 275.75, 275.95, 275.75, 275.55, 275.35, 275.95, 276.15, 274.25, 
    273.05, 274.25, 273.85, 273.85, 276.35, 276.95, 276.85, 276.25, 275.95, 
    274.75, 274.15, 273.55, 273.35, 273.35, 273.25, 273.25, 273.05, 272.85, 
    272.95, 272.85, 273.05, 273.15, 273.05, 273.25, 273.45, 273.55, 273.65, 
    273.65, 273.45, 273.35, 273.35, 273.45, 273.75, 274.25, 273.85, 274.45, 
    274.45, 274.45, 274.95, 275.15, 275.55, 275.45, 274.65, 274.25, 274.35, 
    274.25, 274.25, 274.25, 274.35, 274.45, 274.45, 274.55, 274.65, 274.85, 
    274.85, 274.95, 275.15, 275.35, 275.65, 275.95, 275.45, 275.75, 275.35, 
    275.35, 275.15, 276.35, 274.95, 278.55, 278.95, 277.75, 275.55, 274.15, 
    276.45, 278.85, 275.65, 276.05, 275.95, 275.25, 275.65, 274.95, 275.25, 
    277.95, 277.85, 275.45, 275.15, 276.55, 274.35, 274.65, 273.55, 274.15, 
    274.15, 275.85, 275.95, 274.85, 274.85, 274.35, 274.05, 273.55, 273.75, 
    273.75, 273.65, 273.65, 273.75, 273.65, 273.55, 273.05, 272.95, 273.05, 
    272.95, 273.05, 272.95, 272.85, 272.85, 272.85, 272.95, 273.05, 273.15, 
    273.15, 273.35, 273.25, 273.75, 273.15, 273.95, 274.15, 274.25, 273.25, 
    273.05, 273.45, 273.35, 273.65, 273.75, 273.65, 273.85, 273.95, 274.05, 
    273.95, 273.75, 273.75, 273.55, 273.35, 273.05, 273.05, 273.05, 273.05, 
    273.35, 273.25, 273.35, 273.35, 273.25, 273.35, 273.25, 273.35, 273.15, 
    273.55, 273.25, 273.15, 273.15, 273.15, 272.65, 272.25, 272.05, 271.85, 
    271.65, 271.55, 271.65, 271.95, 271.85, 271.85, 272.05, 271.95, 272.15, 
    272.35, 272.45, 272.75, 272.95, 273.05, 273.15, 272.95, 272.85, 272.75, 
    272.75, 272.75, 272.65, 272.75, 272.45, 272.35, 272.35, 272.15, 272.15, 
    272.05, 271.95, 271.85, 271.85, 272.05, 272.25, 272.35, 272.55, 272.65, 
    272.45, 272.75, 272.65, 272.85, 272.75, 272.75, 272.75, 272.65, 272.95, 
    272.95, 272.75, 272.55, 272.45, 272.45, 272.45, 272.45, 272.55, 272.65, 
    272.75, 272.75, 272.75, 273.05, 273.05, 273.15, 273.15, 272.85, 272.85, 
    272.75, 272.65, 272.85, 272.45, 272.45, 272.15, 272.35, 272.05, 271.95, 
    272.15, 272.15, 272.35, 272.35, 272.45, 272.45, 272.65, 272.75, 272.95, 
    273.45, 273.85, 273.85, 273.65, 274.05, 274.35, 274.25, 274.05, 274.05, 
    274.25, 274.15, 274.05, 273.95, 274.55, 275.05, 274.75, 274.65, 273.85, 
    274.05, 273.65, 273.65, 273.65, 273.35, 272.35, 272.95, 272.85, 272.35, 
    272.55, 272.95, 273.05, 273.45, 272.85, 272.55, 272.45, 272.15, 272.05, 
    272.45, 272.75, 272.55, 272.75, 272.85, 272.95, 273.15, 273.15, 273.15, 
    273.35, 273.35, 273.35, 273.35, 273.35, 273.45, 273.45, 273.35, 273.55, 
    273.45, 273.45, 273.45, 273.45, 273.65, 273.55, 273.45, 273.45, 273.35, 
    273.35, 273.45, 273.45, 273.45, 273.55, 273.55, 273.55, 272.65, 272.85, 
    272.95, 273.05, 273.15, 273.15, 273.15, 273.25, 273.25, 273.25, 273.05, 
    272.85, 272.65, 272.65, 272.55, 272.45, 272.35, 272.35, 272.25, 272.25, 
    272.35, 272.45, 272.55, 272.55, 272.95, 273.05, 271.85, 271.75, 273.45, 
    271.45, 271.95, 273.05, 272.85, 272.65, 272.45, 272.35, 272.95, 272.75, 
    272.55, 272.45, 272.35, 272.35, 272.25, 272.25, 272.25, 272.45, 272.55, 
    272.75, 273.05, 273.05, 272.45, 273.15, 273.45, 274.05, 274.65, 275.15, 
    275.05, 275.45, 275.45, 275.35, 275.25, 275.35, 274.75, 273.85, 273.35, 
    273.05, 272.95, 273.05, 272.95, 273.05, 273.45, 273.35, 273.35, 273.15, 
    272.85, 272.45, 272.25, 272.25, 272.45, 272.65, 272.65, 272.65, 272.75, 
    272.75, 272.75, 272.15, 272.25, 271.65, 270.65, 269.75, 269.45, 268.45, 
    269.95, 270.55, 271.05, 271.15, 271.15, 271.25, 271.25, 271.25, 270.75, 
    270.25, 270.35, 270.55, 270.75, 270.35, 270.55, 270.05, 270.05, 270.35, 
    270.55, 270.95, 271.25, 271.15, 271.05, 271.05, 270.95, 270.85, 271.55, 
    272.05, 272.35, 272.35, 272.55, 272.95, 273.45, 273.45, 273.65, 273.55, 
    273.55, 273.55, 273.35, 273.35, 273.35, 273.25, 273.25, 273.15, 273.15, 
    273.05, 273.05, 273.05, 273.05, 273.15, 273.15, 273.15, 273.05, 273.05, 
    272.35, 272.35, 272.35, 272.45, 272.35, 272.45, 272.55, 272.45, 272.45, 
    272.55, 272.95, 272.95, 272.95, 272.85, 272.85, 272.85, 272.65, 272.45, 
    272.85, 274.35, 274.55, 274.25, 274.25, 274.15, 274.05, 274.05, 274.35, 
    275.95, 275.85, 275.15, 275.15, 275.85, 273.85, 274.85, 273.95, 273.85, 
    273.85, 273.85, 273.85, 273.75, 273.75, 273.75, 273.85, 273.65, 273.35, 
    273.25, 273.25, 273.85, 273.95, 274.05, 274.85, 275.25, 274.95, 274.75, 
    274.55, 274.45, 274.75, 275.25, 275.75, 276.15, 276.25, 276.15, 276.05, 
    275.85, 275.75, 275.75, 275.25, 275.05, 275.15, 275.15, 275.35, 275.05, 
    274.15, 273.75, 273.95, 273.95, 273.35, 272.75, 272.25, 272.05, 271.75, 
    271.55, 271.35, 271.15, 270.75, 270.55, 270.85, 270.95, 271.15, 271.45, 
    271.75, 272.05, 272.35, 272.75, 273.05, 273.35, 273.65, 273.95, 273.65, 
    274.05, 273.55, 273.65, 273.65, 273.45, 273.35, 273.35, 273.35, 273.25, 
    273.15, 273.05, 273.15, 273.15, 273.15, 273.15, 272.75, 272.95, 273.15, 
    272.95, 272.95, 273.25, 273.35, 273.45, 273.35, 273.55, 273.25, 273.45, 
    273.45, 273.45, 273.35, 273.35, 272.55, 271.85, 271.65, 271.45, 271.35, 
    271.25, 272.05, 272.25, 272.55, 272.75, 272.95, 273.25, 273.25, 273.05, 
    272.75, 272.35, 272.25, 272.45, 272.45, 272.55, 272.45, 272.45, 272.35, 
    272.15, 272.05, 271.85, 271.65, 271.65, 271.35, 271.55, 271.35, 271.25, 
    271.35, 271.65, 272.15, 272.45, 272.95, 273.25, 273.35, 273.25, 273.15, 
    272.45, 271.95, 271.75, 271.75, 272.15, 271.95, 271.35, 271.25, 270.95, 
    270.65, 270.05, 270.05, 270.45, 270.55, 270.85, 271.25, 271.05, 270.75, 
    270.25, 270.15, 270.45, 270.85, 271.05, 271.65, 272.25, 272.45, 272.65, 
    272.75, 272.75, 272.75, 272.65, 272.55, 272.35, 272.15, 272.05, 272.25, 
    272.05, 271.85, 271.65, 271.75, 271.95, 272.25, 272.45, 272.55, 272.45, 
    272.25, 272.35, 272.15, 272.45, 272.35, 272.35, 272.35, 272.35, 272.35, 
    272.35, 272.15, 272.05, 271.95, 271.85, 271.85, 271.75, 271.65, 271.65, 
    271.45, 271.15, 270.75, 270.75, 271.05, 271.55, 271.75, 272.05, 272.15, 
    272.55, 272.45, 272.55, 272.65, 272.55, 272.45, 272.25, 272.05, 271.75, 
    271.05, 270.65, 270.15, 269.65, 269.15, 268.45, 268.25, 268.65, 268.85, 
    269.05, 268.95, 268.75, 268.55, 268.05, 268.25, 268.45, 268.45, 268.45, 
    268.85, 268.85, 268.75, 269.55, 269.25, 268.45, 268.15, 268.15, 268.35, 
    268.75, 268.75, 268.85, 268.85, 268.35, 268.05, 267.75, 270.15, 268.75, 
    269.05, 269.25, 269.45, 270.65, 269.95, 270.05, 269.85, 269.95, 270.75, 
    270.65, 270.45, 270.35, 270.15, 270.15, 270.25, 270.25, 270.35, 270.35, 
    270.25, 271.75, 271.85, 271.95, 272.45, 272.55, 272.85, 273.05, 273.15, 
    273.05, 273.05, 272.95, 272.95, 272.95, 272.75, 272.65, 272.65, 272.55, 
    272.45, 272.25, 272.05, 271.95, 271.95, 271.65, 271.65, 271.55, 271.45, 
    271.35, 271.25, 271.45, 271.45, 271.75, 271.75, 271.65, 271.45, 271.25, 
    271.15, 271.35, 271.45, 271.55, 271.55, 271.65, 271.75, 272.25, 271.85, 
    271.25, 270.65, 270.35, 270.35, 270.75, 270.75, 270.75, 270.75, 270.75, 
    270.75, 270.65, 270.65, 271.05, 271.05, 271.15, 271.25, 271.15, 271.15, 
    271.05, 271.15, 271.35, 271.55, 271.65, 271.75, 271.75, 271.85, 271.85, 
    271.65, 271.65, 270.95, 271.35, 271.85, 271.95, 272.15, 272.25, 272.45, 
    272.55, 272.55, 272.45, 272.05, 271.65, 271.25, 271.05, 270.85, 270.75, 
    270.65, 270.75, 270.85, 270.85, 270.75, 270.95, 271.05, 271.05, 271.15, 
    271.45, 271.05, 271.05, 270.85, 270.75, 271.25, 271.25, 271.25, 271.35, 
    271.55, 271.65, 271.85, 271.95, 271.55, 271.45, 271.05, 270.85, 270.95, 
    270.85, 270.85, 270.55, 270.75, 271.05, 271.45, 271.45, 272.35, 273.45, 
    274.95, 274.05, 274.75, 275.25, 275.25, 275.05, 274.95, 274.75, 274.55, 
    274.35, 274.15, 274.35, 274.35, 274.65, 275.05, 274.85, 274.95, 275.05, 
    275.05, 275.05, 274.95, 274.65, 274.75, 274.75, 274.55, 274.65, 274.75, 
    274.85, 274.45, 274.25, 274.25, 274.15, 274.55, 274.45, 274.45, 274.45, 
    274.35, 274.45, 274.55, 274.45, 274.15, 273.75, 273.45, 273.15, 273.15, 
    273.55, 273.95, 274.15, 274.95, 274.85, 274.45, 274.85, 274.65, 274.45, 
    274.05, 273.75, 273.25, 273.35, 272.65, 272.45, 271.85, 271.85, 271.25, 
    271.65, 271.75, 271.65, 270.35, 270.45, 270.15, 269.95, 269.65, 270.15, 
    270.15, 270.35, 270.15, 270.75, 271.25, 271.45, 271.75, 272.05, 272.25, 
    272.25, 272.85, 272.95, 272.15, 272.05, 272.05, 272.25, 272.25, 272.25, 
    272.25, 272.25, 271.15, 270.85, 271.05, 271.05, 270.95, 271.45, 271.75, 
    271.85, 271.85, 271.95, 271.95, 272.05, 272.15, 272.25, 272.05, 271.85, 
    271.45, 271.25, 270.85, 270.75, 270.95, 271.05, 271.05, 270.45, 270.25, 
    270.05, 269.85, 269.95, 270.45, 270.65, 270.75, 270.35, 270.65, 270.75, 
    271.25, 271.55, 270.85, 269.55, 268.65, 269.15, 269.05, 268.65, 268.85, 
    269.05, 268.95, 268.35, 268.65, 268.65, 268.15, 268.45, 268.25, 268.05, 
    267.95, 268.15, 268.65, 269.05, 270.15, 269.55, 269.25, 269.15, 268.25, 
    267.85, 268.15, 268.45, 268.75, 269.05, 269.35, 269.65, 269.55, 269.55, 
    268.95, 267.85, 266.95, 267.55, 268.15, 268.85, 269.45, 268.85, 268.15, 
    267.65, 268.05, 268.95, 268.85, 268.95, 268.25, 268.35, 269.15, 268.95, 
    268.75, 268.65, 268.45, 268.25, 268.05, 267.95, 267.75, 267.55, 267.85, 
    268.45, 269.05, 269.25, 269.15, 270.05, 270.05, 270.35, 270.05, 269.65, 
    269.25, 268.85, 268.55, 268.15, 267.75, 267.35, 267.05, 266.75, 266.75, 
    266.95, 267.15, 266.75, 266.65, 266.45, 266.75, 267.05, 267.35, 267.95, 
    268.85, 268.95, 268.65, 268.65, 268.85, 267.95, 268.15, 268.75, 269.15, 
    269.45, 269.85, 270.35, 270.65, 270.75, 271.35, 271.45, 271.35, 271.35, 
    271.55, 271.75, 271.95, 272.25, 272.55, 272.85, 273.05, 273.35, 273.45, 
    273.95, 274.05, 274.05, 273.85, 273.85, 273.85, 273.85, 273.75, 273.75, 
    273.75, 273.85, 273.75, 273.45, 273.15, 272.45, 271.75, 270.95, 270.35, 
    269.95, 269.75, 269.45, 269.15, 268.85, 268.95, 268.25, 267.15, 266.15, 
    266.05, 265.55, 265.25, 265.35, 265.75, 265.85, 265.75, 265.65, 265.45, 
    265.65, 266.25, 266.65, 266.95, 267.55, 267.85, 268.15, 268.15, 268.05, 
    268.05, 268.45, 268.65, 268.35, 268.15, 268.45, 268.65, 269.05, 269.35, 
    269.55, 269.75, 269.85, 269.85, 269.05, 270.05, 270.45, 270.75, 270.75, 
    270.75, 270.75, 270.75, 271.25, 271.45, 271.15, 271.55, 271.55, 271.55, 
    271.65, 271.35, 271.15, 271.35, 271.45, 272.45, 272.15, 272.55, 272.85, 
    271.35, 271.15, 271.05, 270.95, 270.85, 270.75, 270.45, 270.45, 270.45, 
    270.55, 270.75, 269.75, 269.85, 270.05, 270.35, 270.75, 270.75, 271.05, 
    271.55, 271.95, 272.55, 272.15, 272.35, 271.95, 271.65, 271.35, 271.15, 
    270.85, 270.55, 270.25, 270.05, 269.65, 269.45, 269.55, 270.35, 271.55, 
    271.05, 270.35, 269.85, 269.15, 268.65, 268.15, 267.95, 268.45, 268.45, 
    268.45, 267.85, 267.75, 267.65, 267.65, 267.85, 267.95, 268.15, 268.15, 
    267.75, 267.85, 267.45, 267.35, 267.75, 268.05, 268.55, 269.05, 269.55, 
    269.85, 269.95, 269.55, 269.15, 268.95, 269.05, 269.75, 269.85, 269.75, 
    269.55, 269.75, 270.25, 270.65, 270.65, 271.45, 272.05, 273.05, 273.75, 
    273.85, 273.85, 273.85, 273.95, 274.05, 274.05, 274.35, 274.45, 274.55, 
    274.45, 274.45, 274.85, 275.05, 275.05, 275.25, 275.15, 274.85, 274.25, 
    274.15, 273.85, 273.75, 273.75, 273.75, 273.35, 272.95, 273.15, 273.25, 
    272.95, 273.45, 273.35, 272.75, 272.55, 271.95, 271.85, 271.75, 271.55, 
    271.25, 271.15, 271.05, 270.95, 271.05, 271.05, 271.05, 271.15, 271.45, 
    271.75, 271.55, 271.15, 271.35, 271.35, 271.45, 271.65, 271.75, 271.65, 
    271.35, 271.25, 271.15, 270.95, 270.65, 270.35, 270.15, 270.15, 270.35, 
    270.35, 270.45, 270.55, 270.65, 270.85, 271.65, 271.85, 272.25, 272.55, 
    272.65, 272.95, 273.25, 273.55, 273.75, 273.75, 273.85, 274.25, 274.25, 
    273.85, 274.25, 274.45, 274.45, 274.55, 274.55, 274.55, 274.65, 275.15, 
    274.65, 274.65, 273.65, 273.75, 273.85, 273.45, 273.45, 273.55, 273.65, 
    273.65, 273.55, 273.75, 273.75, 272.65, 271.85, 271.35, 271.05, 270.85, 
    270.75, 270.55, 270.35, 270.35, 269.35, 269.55, 269.35, 269.15, 269.25, 
    269.05, 268.95, 268.85, 268.75, 268.65, 268.15, 268.55, 269.15, 270.05, 
    270.05, 270.05, 269.85, 269.75, 269.65, 269.55, 269.45, 269.45, 269.35, 
    269.25, 269.05, 269.05, 269.15, 268.95, 268.95, 269.15, 269.35, 269.45, 
    269.35, 269.15, 268.95, 268.85, 269.85, 270.05, 269.55, 270.15, 270.15, 
    269.95, 269.45, 269.15, 269.55, 269.55, 269.65, 269.65, 269.75, 269.75, 
    269.85, 269.85, 269.65, 269.95, 270.65, 270.35, 270.35, 270.25, 270.45, 
    270.15, 269.55, 269.05, 268.75, 268.65, 268.65, 268.85, 269.05, 269.65, 
    270.25, 270.25, 269.85, 269.45, 269.45, 270.35, 270.65, 270.45, 270.95, 
    271.65, 272.05, 272.15, 272.25, 272.35, 272.35, 272.45, 272.55, 272.55, 
    272.45, 272.25, 272.15, 272.05, 271.85, 271.75, 271.65, 271.55, 271.35, 
    271.25, 271.15, 271.05, 270.95, 270.75, 270.65, 270.55, 270.45, 270.35, 
    270.45, 270.35, 270.75, 270.65, 270.85, 270.85, 270.85, 270.75, 270.75, 
    270.85, 270.75, 270.65, 270.55, 270.55, 270.55, 270.55, 270.65, 270.75, 
    270.75, 270.75, 270.75, 270.75, 270.55, 270.65, 270.75, 270.55, 270.85, 
    270.95, 271.05, 271.15, 271.25, 271.15, 270.95, 271.25, 271.35, 271.25, 
    271.05, 270.85, 270.75, 270.85, 270.75, 271.25, 271.25, 271.15, 271.45, 
    271.55, 271.25, 271.15, 271.45, 271.75, 272.05, 272.05, 272.55, 273.05, 
    273.15, 273.35, 272.95, 273.05, 272.75, 272.75, 273.05, 272.75, 272.65, 
    272.45, 272.35, 272.15, 271.95, 271.85, 271.75, 271.65, 271.65, 272.45, 
    272.45, 272.45, 272.35, 272.35, 272.15, 272.15, 272.25, 272.45, 272.25, 
    272.25, 271.95, 272.05, 272.05, 272.05, 272.05, 272.15, 272.25, 272.35, 
    272.35, 272.25, 272.25, 272.25, 272.25, 272.25, 272.25, 272.45, 272.65, 
    272.15, 271.95, 271.85, 272.15, 271.25, 271.35, 273.25, 273.25, 273.15, 
    273.05, 273.05, 273.05, 273.15, 273.15, 273.05, 272.35, 272.45, 272.45, 
    271.85, 271.65, 271.45, 271.45, 271.45, 271.45, 271.35, 271.15, 271.15, 
    271.15, 271.15, 271.25, 271.25, 271.25, 271.35, 271.35, 271.35, 271.25, 
    271.15, 270.95, 270.75, 270.65, 270.45, 270.15, 270.15, 270.05, 269.85, 
    269.75, 269.85, 269.85, 269.65, 269.55, 269.45, 269.35, 269.25, 269.15, 
    269.45, 269.65, 269.15, 268.65, 268.45, 268.25, 268.15, 267.95, 267.85, 
    267.75, 267.35, 267.25, 266.95, 266.55, 266.35, 265.85, 265.45, 265.55, 
    265.95, 266.35, 266.55, 266.65, 266.65, 266.55, 267.15, 266.85, 266.95, 
    267.15, 267.25, 267.15, 266.85, 266.85, 266.95, 266.95, 266.55, 266.35, 
    266.15, 266.05, 266.05, 266.05, 265.95, 265.45, 265.25, 265.95, 264.95, 
    266.55, 266.65, 267.15, 267.35, 267.45, 267.65, 268.05, 268.65, 268.95, 
    267.85, 267.35, 266.95, 266.55, 266.25, 266.65, 266.65, 266.75, 266.75, 
    266.85, 266.85, 266.65, 266.95, 267.55, 267.75, 267.55, 267.35, 267.85, 
    268.25, 268.45, 268.55, 268.25, 266.85, 266.35, 265.65, 265.35, 265.25, 
    265.55, 266.35, 266.95, 267.65, 268.05, 268.25, 268.45, 268.65, 270.05, 
    270.55, 271.05, 272.05, 272.25, 272.55, 272.95, 273.35, 273.45, 273.45, 
    273.85, 273.85, 273.15, 272.95, 272.85, 272.85, 272.85, 272.65, 272.25, 
    271.75, 271.35, 270.85, 270.35, 270.25, 269.95, 269.65, 269.05, 268.55, 
    268.45, 268.55, 268.65, 268.25, 267.75, 267.55, 267.55, 267.25, 266.75, 
    266.15, 265.65, 265.15, 264.75, 265.65, 267.45, 267.65, 267.35, 267.15, 
    267.05, 266.55, 266.95, 267.45, 267.75, 268.05, 268.95, 270.05, 269.45, 
    271.05, 270.25, 270.85, 271.45, 272.15, 272.75, 273.25, 273.45, 274.25, 
    275.05, 274.75, 274.65, 275.75, 275.65, 275.15, 274.85, 274.55, 274.25, 
    273.85, 273.55, 273.25, 272.95, 272.45, 272.35, 272.35, 272.75, 273.35, 
    274.05, 274.35, 274.55, 275.05, 274.85, 274.35, 273.95, 273.85, 273.75, 
    272.85, 272.85, 272.85, 272.65, 272.55, 272.45, 272.35, 272.25, 272.15, 
    272.05, 271.95, 271.65, 271.75, 271.65, 271.55, 271.45, 271.35, 270.95, 
    270.15, 269.45, 269.15, 269.05, 269.35, 269.45, 269.55, 269.55, 269.55, 
    269.65, 269.85, 270.05, 270.25, 270.35, 270.45, 270.65, 270.75, 270.75, 
    270.45, 270.15, 269.95, 269.45, 268.85, 268.95, 269.05, 269.05, 268.55, 
    268.35, 268.25, 267.85, 267.05, 266.95, 267.25, 267.25, 267.25, 267.55, 
    267.55, 267.45, 267.35, 267.15, 267.15, 266.85, 266.85, 266.65, 266.85, 
    267.15, 267.45, 267.65, 267.45, 267.35, 267.35, 266.95, 266.95, 266.95, 
    266.75, 266.65, 266.65, 266.55, 266.55, 266.45, 266.35, 266.45, 266.55, 
    266.45, 267.35, 268.15, 267.95, 267.95, 267.95, 268.05, 268.25, 268.45, 
    268.55, 268.75, 268.95, 269.05, 269.25, 269.45, 269.65, 269.65, 269.85, 
    270.05, 270.25, 270.55, 270.85, 270.75, 269.95, 269.15, 268.25, 266.95, 
    266.45, 266.05, 265.35, 264.55, 263.85, 263.55, 263.65, 264.25, 264.75, 
    265.55, 265.55, 265.25, 265.25, 265.35, 265.55, 266.15, 265.15, 264.95, 
    264.85, 265.05, 264.55, 264.35, 264.45, 264.55, 264.65, 264.45, 263.75, 
    262.95, 262.45, 261.85, 261.05, 261.05, 261.25, 261.55, 261.75, 261.65, 
    261.85, 261.85, 261.45, 260.95, 260.45, 260.45, 260.35, 260.25, 260.05, 
    259.95, 259.85, 259.55, 260.15, 260.65, 261.35, 261.35, 261.35, 261.45, 
    261.55, 261.95, 261.85, 262.45, 262.05, 261.35, 260.95, 260.65, 260.65, 
    260.95, 261.45, 262.25, 262.25, 261.55, 263.25, 264.05, 263.55, 263.05, 
    262.95, 262.75, 262.35, 261.95, 260.65, 260.95, 261.25, 261.75, 262.15, 
    262.15, 261.65, 261.15, 260.75, 260.25, 259.85, 259.35, 258.05, 258.15, 
    257.85, 257.65, 258.25, 258.35, 258.75, 258.75, 258.15, 258.15, 257.65, 
    256.85, 256.65, 256.75, 255.25, 255.25, 255.75, 255.95, 257.35, 258.55, 
    259.55, 260.15, 259.95, 260.25, 260.45, 261.25, 262.15, 262.75, 263.25, 
    263.55, 263.75, 263.95, 263.95, 264.15, 264.35, 264.05, 263.45, 263.25, 
    263.25, 263.25, 263.15, 263.15, 263.15, 263.15, 263.05, 263.25, 261.95, 
    262.75, 262.45, 262.65, 262.95, 262.95, 262.65, 262.55, 262.55, 262.65, 
    262.75, 262.35, 262.25, 261.65, 261.65, 261.75, 261.85, 262.05, 262.15, 
    262.15, 261.75, 260.65, 260.05, 262.05, 262.95, 263.55, 264.45, 265.55, 
    266.35, 266.25, 266.55, 268.35, 269.95, 267.85, 266.95, 267.45, 265.65, 
    264.55, 263.75, 263.45, 263.85, 264.55, 264.55, 264.35, 263.75, 263.75, 
    263.65, 263.65, 263.75, 263.85, 263.85, 263.95, 264.15, 263.75, 263.55, 
    263.45, 263.35, 263.35, 263.35, 263.25, 262.85, 262.55, 262.35, 262.05, 
    261.75, 261.55, 261.25, 260.85, 260.75, 261.65, 262.05, 260.95, 261.15, 
    260.85, 261.35, 261.95, 262.75, 262.55, 261.85, 261.95, 262.25, 262.65, 
    262.15, 261.95, 261.85, 261.85, 261.85, 261.75, 261.75, 261.55, 261.65, 
    262.25, 262.35, 263.65, 263.15, 264.65, 262.75, 262.65, 262.25, 261.85, 
    261.55, 261.85, 262.95, 263.25, 263.15, 263.45, 265.75, 265.45, 265.25, 
    265.05, 264.85, 265.45, 265.05, 265.15, 264.85, 264.85, 264.85, 265.55, 
    265.95, 269.85, 269.25, 269.35, 269.65, 269.75, 270.15, 269.25, 268.25, 
    267.45, 267.45, 266.05, 264.35, 264.05, 264.35, 264.85, 265.25, 265.75, 
    266.15, 266.65, 266.95, 266.95, 267.45, 268.55, 268.95, 269.25, 269.75, 
    270.25, 270.65, 270.25, 270.15, 270.15, 270.35, 270.15, 269.85, 270.05, 
    270.05, 269.85, 270.05, 270.25, 270.45, 270.65, 270.75, 270.85, 270.95, 
    271.05, 271.25, 271.35, 271.45, 271.75, 271.75, 271.75, 271.75, 271.85, 
    271.95, 271.65, 271.85, 271.75, 271.85, 272.15, 272.35, 272.55, 272.85, 
    272.85, 272.85, 272.85, 272.85, 272.75, 272.75, 272.75, 272.65, 272.65, 
    272.65, 272.55, 272.45, 272.45, 272.55, 272.75, 272.85, 272.85, 272.95, 
    272.95, 272.95, 272.95, 272.85, 272.95, 272.95, 272.95, 272.95, 273.05, 
    273.05, 272.95, 272.85, 272.85, 272.65, 272.65, 272.75, 272.95, 272.95, 
    273.15, 273.35, 273.45, 273.55, 273.65, 273.65, 273.75, 273.55, 273.55, 
    273.55, 273.55, 273.45, 273.45, 273.45, 273.45, 273.35, 273.25, 273.15, 
    272.95, 272.95, 272.75, 272.85, 272.75, 272.75, 272.65, 272.55, 272.35, 
    272.25, 272.15, 272.05, 272.05, 272.05, 271.95, 272.05, 271.95, 271.95, 
    271.95, 272.05, 272.05, 272.05, 272.05, 272.15, 272.15, 272.15, 272.15, 
    272.15, 272.15, 272.05, 271.95, 272.15, 271.85, 271.45, 271.05, 270.65, 
    270.85, 270.75, 270.75, 270.75, 270.75, 270.65, 270.55, 270.45, 270.35, 
    270.35, 270.45, 270.35, 270.25, 270.15, 270.15, 270.15, 270.15, 270.15, 
    270.05, 269.85, 269.75, 269.65, 269.45, 269.25, 269.15, 269.15, 268.95, 
    269.05, 268.85, 268.65, 268.55, 268.65, 268.65, 268.65, 268.55, 268.55, 
    268.55, 268.55, 268.45, 268.45, 268.45, 268.55, 268.55, 268.15, 268.25, 
    268.25, 268.25, 268.05, 267.85, 267.85, 267.85, 267.85, 267.75, 267.75, 
    267.65, 267.65, 267.65, 267.65, 267.35, 266.95, 267.15, 266.85, 266.75, 
    266.65, 266.35, 266.35, 265.95, 265.85, 265.55, 265.35, 265.15, 265.05, 
    264.85, 264.85, 265.05, 264.85, 264.85, 265.05, 265.05, 265.05, 265.05, 
    264.95, 264.95, 264.85, 264.75, 264.65, 264.45, 264.65, 264.65, 263.45, 
    263.95, 264.45, 264.25, 264.05, 264.15, 264.85, 265.25, 265.65, 266.05, 
    266.55, 267.45, 267.75, 267.75, 268.25, 267.95, 267.15, 266.95, 265.55, 
    264.75, 264.35, 263.65, 263.25, 262.85, 262.55, 261.95, 261.05, 260.15, 
    259.35, 258.55, 257.95, 257.65, 257.25, 256.35, 255.25, 255.65, 253.85, 
    254.75, 254.55, 255.25, 255.85, 255.45, 255.35, 255.55, 255.95, 256.05, 
    256.25, 255.85, 256.25, 257.15, 257.25, 257.25, 257.45, 256.45, 256.35, 
    255.95, 255.35, 254.95, 254.35, 254.25, 253.45, 253.15, 253.55, 253.55, 
    253.85, 253.75, 254.75, 255.75, 255.95, 255.95, 255.75, 256.15, 256.15, 
    256.35, 256.65, 257.05, 257.45, 256.05, 255.45, 254.95, 254.85, 254.65, 
    254.75, 254.45, 254.45, 254.45, 254.05, 254.35, 253.95, 253.25, 253.35, 
    252.25, 251.55, 251.35, 251.45, 251.25, 251.05, 251.35, 250.95, 251.45, 
    252.25, 251.95, 253.35, 252.45, 252.45, 252.15, 254.15, 252.35, 252.75, 
    252.85, 253.55, 252.95, 252.95, 253.35, 253.75, 253.85, 255.05, 255.65, 
    256.55, 257.25, 257.65, 258.05, 258.35, 258.45, 259.35, 259.45, 259.65, 
    260.55, 260.05, 259.15, 259.95, 259.65, 259.05, 257.45, 256.55, 254.95, 
    253.65, 251.55, 251.55, 250.65, 249.55, 250.55, 251.35, 250.55, 249.25, 
    248.45, 247.75, 247.75, 248.25, 248.95, 249.35, 250.25, 250.45, 250.65, 
    250.55, 250.15, 249.55, 249.95, 250.35, 250.15, 249.95, 249.65, 250.55, 
    250.95, 250.55, 251.75, 251.75, 252.15, 251.95, 252.05, 252.55, 253.05, 
    253.95, 253.95, 253.85, 254.55, 254.85, 254.85, 254.95, 255.15, 255.35, 
    255.45, 255.85, 256.05, 256.05, 256.05, 256.05, 256.55, 257.15, 257.55, 
    257.55, 257.65, 257.95, 258.35, 258.75, 260.05, 260.45, 260.55, 260.95, 
    261.25, 261.35, 261.35, 261.25, 260.85, 261.35, 260.95, 261.05, 260.45, 
    259.95, 260.05, 260.25, 259.75, 259.25, 258.95, 258.75, 258.25, 257.85, 
    257.35, 256.65, 255.75, 254.75, 254.75, 254.45, 254.45, 254.25, 254.15, 
    253.65, 253.25, 253.05, 253.15, 253.05, 253.45, 253.45, 253.35, 253.85, 
    253.75, 253.45, 253.55, 253.75, 253.65, 253.55, 252.95, 253.25, 253.55, 
    253.85, 254.15, 254.55, 254.45, 254.55, 254.35, 254.35, 254.15, 254.45, 
    254.85, 254.25, 254.15, 254.15, 254.45, 254.65, 254.85, 254.65, 254.95, 
    255.05, 254.65, 253.75, 253.15, 252.65, 252.25, 251.45, 251.65, 251.75, 
    251.75, 251.55, 251.45, 250.85, 250.65, 250.45, 250.15, 250.35, 250.15, 
    250.55, 250.85, 251.55, 252.05, 252.45, 252.85, 253.85, 254.65, 254.45, 
    255.35, 255.75, 255.95, 256.05, 256.25, 256.35, 256.25, 256.05, 255.95, 
    256.25, 256.55, 256.25, 256.05, 255.95, 256.05, 256.85, 257.45, 258.15, 
    258.05, 258.05, 257.95, 257.75, 258.05, 258.05, 258.55, 258.95, 258.65, 
    258.25, 258.35, 258.25, 257.95, 257.95, 258.25, 257.25, 257.15, 257.05, 
    256.85, 256.35, 256.15, 255.95, 255.75, 255.25, 255.25, 255.65, 256.05, 
    255.65, 256.55, 256.55, 257.05, 257.15, 256.75, 255.75, 254.35, 254.15, 
    253.85, 254.25, 255.05, 255.85, 256.75, 257.65, 258.05, 258.75, 257.85, 
    256.85, 257.35, 257.85, 258.35, 258.95, 259.25, 260.25, 260.75, 261.75, 
    263.05, 264.05, 265.05, 266.25, 266.95, 267.65, 268.15, 268.85, 268.95, 
    266.35, 262.55, 258.95, 257.55, 257.05, 256.25, 256.35, 256.35, 256.75, 
    257.05, 256.95, 257.25, 258.35, 258.05, 257.65, 257.05, 256.15, 255.15, 
    254.65, 255.35, 256.35, 257.15, 257.35, 257.65, 260.25, 259.05, 259.55, 
    259.85, 259.75, 257.85, 256.65, 256.35, 254.55, 253.15, 253.05, 252.85, 
    253.25, 253.75, 254.25, 254.85, 254.65, 255.25, 256.05, 256.35, 256.95, 
    256.95, 256.55, 256.45, 256.35, 256.15, 256.35, 256.35, 256.15, 256.35, 
    256.65, 256.15, 256.15, 256.45, 256.35, 256.25, 256.35, 256.55, 256.65, 
    256.75, 257.05, 259.05, 258.25, 257.95, 259.25, 258.25, 259.45, 258.75, 
    258.95, 259.15, 260.75, 260.45, 258.75, 258.55, 257.75, 257.75, 257.15, 
    256.75, 255.35, 255.65, 255.75, 255.55, 255.15, 254.45, 254.25, 253.75, 
    253.45, 253.15, 252.95, 252.85, 252.35, 251.95, 251.05, 249.15, 248.15, 
    247.45, 248.35, 247.85, 246.35, 246.15, 247.45, 247.65, 248.25, 248.45, 
    248.65, 248.15, 247.55, 246.65, 246.35, 246.05, 245.75, 245.85, 246.25, 
    246.25, 246.45, 247.35, 247.85, 247.75, 247.35, 247.45, 248.25, 252.15, 
    251.55, 251.05, 250.95, 250.05, 249.95, 250.55, 251.25, 251.65, 251.25, 
    251.25, 251.65, 252.15, 252.75, 252.85, 253.95, 254.45, 255.45, 256.35, 
    256.65, 257.45, 257.55, 257.95, 258.45, 258.65, 258.95, 259.05, 259.55, 
    260.35, 260.25, 260.85, 261.45, 262.15, 262.65, 263.85, 264.35, 265.25, 
    266.35, 267.05, 268.55, 268.65, 269.05, 269.15, 269.25, 269.35, 269.45, 
    268.15, 267.45, 266.35, 266.95, 267.65, 268.45, 269.25, 269.05, 268.55, 
    268.55, 267.15, 267.25, 267.25, 268.15, 268.05, 268.45, 269.25, 269.35, 
    269.75, 269.85, 269.15, 269.05, 269.35, 269.85, 270.35, 271.25, 271.45, 
    271.85, 271.45, 271.85, 267.35, 261.55, 257.95, 256.35, 254.65, 253.75, 
    253.85, 255.05, 254.95, 254.95, 255.05, 254.85, 254.65, 254.75, 255.05, 
    255.45, 255.35, 255.15, 254.05, 253.25, 252.55, 251.65, 251.25, 250.95, 
    250.75, 250.25, 251.65, 251.85, 250.45, 249.85, 249.35, 249.05, 250.15, 
    250.75, 251.85, 252.25, 253.15, 254.35, 255.95, 257.35, 256.85, 257.35, 
    257.25, 257.55, 256.55, 257.45, 258.75, 260.65, 259.95, 260.45, 260.35, 
    260.75, 261.15, 261.65, 261.95, 262.05, 261.95, 262.65, 262.35, 262.05, 
    261.85, 262.95, 261.85, 262.85, 263.15, 262.85, 262.95, 264.75, 264.85, 
    265.75, 265.95, 266.65, 267.55, 268.25, 269.05, 269.85, 270.55, 270.85, 
    270.95, 271.05, 270.95, 270.15, 269.75, 270.45, 271.35, 272.25, 272.95, 
    272.65, 272.95, 273.15, 273.35, 273.45, 273.35, 273.55, 273.25, 271.55, 
    270.55, 269.85, 269.35, 268.75, 268.05, 267.35, 266.55, 266.35, 265.45, 
    263.95, 263.15, 262.95, 263.05, 263.05, 262.95, 262.75, 262.45, 261.55, 
    260.85, 260.35, 259.85, 260.15, 259.45, 259.15, 258.75, 258.65, 258.85, 
    258.85, 258.75, 259.35, 259.75, 259.85, 259.55, 259.25, 259.45, 259.35, 
    258.95, 258.65, 259.65, 259.35, 258.65, 260.05, 261.25, 261.15, 261.55, 
    261.45, 260.35, 259.85, 259.95, 259.95, 259.95, 259.95, 259.85, 259.95, 
    260.35, 260.75, 260.85, 260.65, 260.65, 260.75, 260.65, 261.05, 261.25, 
    261.55, 261.35, 261.75, 261.55, 261.95, 262.25, 262.65, 262.95, 263.85, 
    264.75, 265.05, 265.25, 266.05, 267.35, 267.45, 267.75, 267.35, 267.25, 
    266.85, 266.75, 266.75, 266.75, 266.15, 265.95, 265.45, 265.25, 264.55, 
    264.05, 263.25, 262.15, 260.75, 259.35, 258.15, 257.55, 256.35, 257.05, 
    256.95, 256.45, 255.05, 254.75, 255.05, 254.35, 254.55, 255.25, 255.45, 
    255.85, 256.05, 255.55, 255.35, 254.35, 254.55, 253.55, 253.55, 253.35, 
    253.55, 253.35, 253.15, 253.05, 253.65, 254.25, 254.05, 253.85, 253.25, 
    253.15, 253.55, 254.45, 255.55, 255.75, 255.75, 255.85, 256.15, 256.45, 
    256.75, 256.55, 255.95, 255.65, 255.35, 255.65, 255.05, 255.15, 255.35, 
    255.75, 255.45, 255.95, 255.55, 256.95, 255.65, 255.35, 255.65, 256.65, 
    257.85, 258.65, 259.55, 259.35, 260.05, 260.45, 260.15, 258.95, 258.95, 
    258.85, 258.85, 258.85, 259.35, 259.75, 259.75, 259.35, 258.35, 257.45, 
    257.15, 256.65, 256.65, 255.65, 256.65, 254.95, 256.45, 256.55, 256.75, 
    256.65, 256.65, 255.45, 256.35, 256.65, 256.95, 257.15, 257.25, 257.65, 
    257.75, 257.25, 256.95, 256.75, 257.45, 258.35, 258.85, 259.05, 258.55, 
    258.15, 257.85, 257.95, 257.95, 257.55, 258.75, 260.05, 261.35, 262.75, 
    263.45, 263.65, 264.25, 265.45, 266.55, 266.55, 266.25, 266.05, 266.15, 
    266.35, 266.45, 266.65, 266.65, 266.75, 266.75, 266.75, 266.65, 266.35, 
    265.55, 264.75, 264.05, 263.45, 262.75, 262.25, 262.05, 261.35, 260.95, 
    260.75, 261.05, 261.25, 261.55, 261.45, 261.35, 261.95, 262.15, 262.05, 
    262.05, 262.05, 262.25, 262.45, 262.45, 262.75, 262.45, 262.45, 262.15, 
    262.35, 262.45, 262.65, 263.25, 263.05, 262.55, 262.75, 263.05, 263.45, 
    263.15, 263.25, 263.25, 262.65, 262.75, 262.45, 263.35, 264.95, 265.05, 
    263.65, 262.85, 262.65, 261.65, 260.55, 259.55, 259.95, 258.75, 258.35, 
    257.75, 258.45, 258.05, 259.45, 260.55, 260.45, 260.25, 260.35, 260.55, 
    259.85, 260.75, 260.65, 261.15, 261.65, 261.65, 261.65, 261.35, 260.75, 
    261.35, 262.65, 262.45, 262.25, 262.25, 261.75, 260.95, 260.45, 260.15, 
    260.15, 260.15, 260.15, 260.85, 260.45, 260.75, 260.35, 260.35, 260.15, 
    260.15, 260.15, 260.95, 261.55, 261.45, 261.55, 262.45, 262.65, 262.55, 
    262.85, 263.85, 263.85, 265.05, 266.25, 265.65, 266.25, 266.05, 267.25, 
    268.85, 269.45, 269.65, 269.75, 270.05, 270.25, 270.55, 270.75, 271.05, 
    271.15, 271.25, 271.35, 271.25, 271.25, 270.95, 270.85, 271.55, 271.15, 
    270.85, 270.75, 270.45, 269.55, 269.45, 269.25, 268.15, 267.65, 267.55, 
    263.95, 263.35, 262.55, 262.25, 261.85, 261.65, 262.65, 262.95, 264.05, 
    264.75, 265.15, 265.85, 265.15, 265.15, 264.85, 265.55, 265.95, 265.85, 
    265.45, 264.95, 264.15, 263.25, 261.95, 261.55, 261.25, 260.95, 260.85, 
    260.85, 260.25, 261.05, 257.25, 255.05, 260.95, 262.15, 261.55, 262.65, 
    262.95, 262.25, 263.05, 263.45, 263.15, 263.65, 263.05, 263.25, 265.25, 
    265.85, 265.85, 267.15, 268.05, 268.65, 270.65, 271.15, 271.45, 271.35, 
    271.85, 271.65, 272.15, 271.55, 271.15, 270.85, 270.75, 270.55, 270.45, 
    269.85, 269.55, 270.05, 270.05, 270.15, 270.65, 270.05, 269.95, 269.25, 
    267.75, 266.85, 266.55, 266.25, 266.35, 266.55, 266.65, 266.95, 267.15, 
    265.15, 263.15, 264.05, 261.75, 260.45, 261.35, 261.85, 262.05, 261.95, 
    261.75, 262.25, 261.45, 263.35, 261.45, 260.65, 259.35, 258.85, 258.45, 
    257.55, 259.05, 259.95, 260.65, 261.45, 262.15, 263.05, 261.55, 262.05, 
    262.95, 263.05, 263.65, 264.35, 265.45, 265.55, 265.55, 265.15, 263.05, 
    264.15, 264.35, 264.55, 264.65, 264.15, 264.05, 263.85, 263.65, 262.75, 
    262.45, 261.95, 261.85, 261.75, 261.25, 260.65, 261.25, 260.45, 261.65, 
    261.85, 261.95, 262.75, 262.55, 261.45, 261.95, 261.65, 260.95, 259.95, 
    260.35, 257.35, 255.35, 254.25, 259.45, 252.65, 251.85, 248.65, 250.85, 
    255.05, 257.15, 257.05, 254.95, 254.85, 255.65, 256.35, 257.65, 258.35, 
    259.55, 260.35, 260.85, 261.25, 261.95, 262.05, 262.15, 261.45, 261.05, 
    260.95, 260.35, 260.35, 259.85, 259.15, 259.05, 258.65, 258.15, 257.85, 
    257.45, 256.85, 256.45, 256.55, 256.55, 256.55, 256.05, 255.85, 255.65, 
    255.45, 254.95, 254.35, 253.75, 253.95, 253.45, 253.75, 253.75, 253.35, 
    252.85, 252.65, 252.95, 252.85, 252.75, 252.35, 252.25, 251.95, 252.15, 
    252.25, 252.45, 251.75, 251.95, 251.75, 252.45, 252.25, 252.45, 252.55, 
    252.15, 253.15, 253.25, 252.65, 251.65, 250.75, 250.45, 250.65, 251.95, 
    251.05, 251.25, 251.95, 252.05, 251.15, 250.75, 250.45, 250.05, 250.95, 
    251.25, 251.55, 250.95, 251.25, 251.15, 251.35, 252.05, 252.85, 251.95, 
    251.25, 250.45, 248.95, 248.15, 248.55, 248.55, 248.65, 248.75, 249.25, 
    249.45, 248.55, 248.85, 249.35, 248.15, 247.35, 247.85, 248.05, 248.15, 
    248.55, 248.85, 248.85, 249.95, 250.65, 250.35, 249.65, 248.15, 247.05, 
    246.85, 246.95, 247.75, 247.55, 246.15, 245.55, 245.75, 246.45, 246.45, 
    247.45, 248.25, 247.95, 247.35, 247.05, 247.15, 246.55, 246.05, 245.35, 
    245.65, 245.95, 246.25, 245.45, 245.05, 245.05, 244.85, 245.25, 245.35, 
    246.35, 244.25, 244.35, 244.65, 245.45, 245.45, 245.75, 246.15, 246.55, 
    246.85, 247.25, 247.15, 247.25, 247.65, 248.65, 248.65, 248.65, 248.85, 
    249.15, 249.55, 249.75, 249.55, 249.25, 248.95, 248.25, 247.35, 247.35, 
    247.85, 248.45, 248.65, 248.15, 247.85, 248.15, 248.55, 247.75, 245.85, 
    244.95, 244.75, 245.25, 247.15, 247.45, 247.45, 247.45, 247.45, 247.05, 
    246.65, 246.45, 246.45, 246.45, 246.75, 247.05, 246.95, 246.85, 246.65, 
    246.35, 246.55, 246.65, 246.05, 245.65, 245.05, 244.55, 244.45, 243.95, 
    244.75, 244.25, 244.35, 244.45, 244.75, 244.35, 243.75, 243.45, 244.95, 
    243.95, 246.35, 248.65, 249.65, 249.65, 250.05, 249.45, 249.05, 249.05, 
    249.85, 249.85, 249.65, 249.65, 248.75, 249.15, 248.85, 249.15, 248.85, 
    250.35, 250.05, 250.25, 250.45, 250.25, 250.95, 250.15, 248.95, 249.15, 
    249.25, 249.85, 249.45, 249.75, 250.05, 249.75, 249.85, 250.05, 249.95, 
    249.95, 250.55, 251.35, 252.65, 252.45, 253.15, 253.55, 253.55, 253.55, 
    253.25, 252.95, 253.35, 253.35, 253.55, 253.85, 254.35, 254.85, 255.25, 
    256.95, 259.25, 260.65, 261.75, 262.85, 263.95, 265.15, 266.05, 266.85, 
    267.25, 266.95, 266.75, 267.25, 268.15, 268.65, 268.95, 269.45, 269.55, 
    269.75, 269.55, 269.35, 269.05, 268.65, 268.35, 267.75, 267.65, 267.65, 
    267.85, 268.15, 268.55, 268.55, 268.75, 268.75, 268.95, 269.05, 269.15, 
    269.25, 269.45, 269.55, 269.65, 269.85, 269.95, 269.95, 269.85, 269.75, 
    269.65, 269.65, 269.55, 269.45, 269.55, 269.75, 269.75, 269.75, 269.95, 
    269.95, 269.95, 269.95, 270.05, 269.95, 269.85, 269.85, 269.85, 269.85, 
    269.75, 269.75, 269.85, 270.35, 270.45, 270.35, 269.75, 269.45, 269.25, 
    269.15, 268.95, 268.85, 268.65, 268.55, 268.45, 268.45, 268.45, 268.45, 
    268.45, 268.55, 268.35, 268.15, 267.95, 268.15, 268.35, 268.05, 268.65, 
    268.55, 268.45, 268.35, 268.15, 268.15, 267.85, 267.75, 267.55, 267.55, 
    267.25, 267.35, 267.35, 267.35, 267.25, 266.55, 266.25, 266.35, 265.15, 
    264.45, 264.95, 264.35, 264.45, 263.45, 263.65, 264.45, 264.75, 265.25, 
    265.05, 264.75, 264.35, 264.65, 264.65, 264.75, 265.05, 264.85, 264.75, 
    264.75, 264.55, 265.45, 265.15, 265.35, 265.45, 265.15, 265.85, 265.65, 
    265.55, 265.85, 265.95, 266.05, 266.05, 265.95, 266.15, 266.85, 266.95, 
    266.95, 266.35, 263.45, 263.45, 262.75, 262.45, 261.65, 262.65, 262.75, 
    263.15, 263.35, 262.75, 262.95, 263.15, 262.85, 262.25, 262.55, 263.75, 
    262.35, 262.65, 263.35, 263.75, 263.45, 263.45, 263.95, 263.65, 263.55, 
    262.85, 262.05, 262.35, 263.05, 263.15, 263.95, 264.75, 265.25, 266.15, 
    267.25, 267.95, 268.25, 268.95, 269.15, 269.35, 269.55, 269.65, 269.75, 
    269.65, 269.45, 269.35, 269.35, 268.85, 268.95, 269.05, 269.25, 269.45, 
    269.65, 269.95, 270.05, 270.45, 270.15, 270.25, 270.15, 270.55, 271.15, 
    271.65, 271.45, 271.15, 270.75, 270.45, 269.55, 269.55, 269.25, 269.05, 
    268.55, 267.85, 266.45, 266.25, 266.95, 269.05, 268.85, 268.75, 267.95, 
    268.35, 269.65, 270.55, 270.45, 270.05, 269.55, 269.45, 269.45, 269.35, 
    269.05, 268.95, 269.15, 268.85, 269.55, 269.75, 269.55, 269.85, 269.95, 
    269.75, 269.95, 269.65, 269.75, 269.85, 269.65, 269.65, 269.85, 269.85, 
    269.65, 269.85, 269.85, 269.35, 269.75, 269.35, 269.65, 269.35, 269.55, 
    269.05, 267.45, 266.45, 265.35, 264.25, 263.05, 262.15, 261.35, 260.85, 
    260.45, 260.15, 258.15, 257.25, 257.05, 256.85, 256.45, 256.25, 256.05, 
    256.55, 256.65, 255.95, 256.55, 256.55, 256.45, 255.65, 258.75, 259.65, 
    259.55, 259.75, 259.85, 260.55, 260.75, 261.55, 261.15, 261.35, 261.25, 
    261.35, 260.85, 261.05, 261.05, 260.95, 260.75, 260.35, 259.65, 259.65, 
    259.95, 260.35, 260.65, 261.55, 262.65, 264.45, 264.85, 264.55, 265.45, 
    265.55, 265.75, 263.95, 260.75, 260.15, 258.95, 260.45, 260.35, 260.15, 
    261.25, 260.35, 259.45, 258.75, 257.85, 258.75, 259.75, 260.45, 260.05, 
    260.45, 260.15, 259.35, 258.85, 258.55, 258.15, 257.95, 257.35, 257.75, 
    257.15, 256.95, 257.75, 257.55, 258.35, 258.65, 257.55, 256.15, 255.95, 
    256.15, 255.85, 255.55, 255.45, 255.35, 255.45, 255.35, 255.55, 255.15, 
    255.25, 255.45, 256.05, 255.25, 255.05, 254.55, 252.45, 254.05, 253.05, 
    254.05, 253.75, 252.85, 253.45, 252.95, 253.45, 253.75, 252.15, 251.25, 
    253.55, 253.95, 253.35, 253.45, 254.05, 254.25, 255.75, 255.45, 256.65, 
    257.05, 256.55, 257.35, 255.95, 256.15, 256.55, 256.45, 256.75, 257.05, 
    255.95, 254.15, 252.35, 253.55, 253.35, 252.25, 252.05, 251.75, 251.25, 
    249.75, 249.55, 251.35, 249.05, 249.15, 248.55, 247.65, 247.55, 247.65, 
    247.55, 248.75, 248.75, 248.55, 250.35, 247.25, 246.85, 247.55, 247.65, 
    247.55, 247.25, 246.85, 246.75, 246.75, 246.55, 246.35, 246.95, 246.75, 
    246.85, 245.95, 246.45, 246.85, 247.65, 248.15, 248.65, 248.75, 248.85, 
    249.35, 250.05, 250.65, 250.35, 251.95, 256.15, 253.25, 251.85, 253.65, 
    253.65, 252.55, 255.45, 255.85, 254.55, 254.75, 254.65, 253.75, 256.05, 
    255.15, 255.05, 254.85, 253.35, 252.05, 251.15, 250.35, 249.55, 248.55, 
    248.75, 248.25, 248.35, 249.45, 249.85, 250.05, 251.55, 248.45, 248.55, 
    248.95, 250.55, 252.05, 253.45, 253.65, 254.55, 255.05, 256.25, 256.85, 
    257.55, 256.35, 256.05, 255.95, 256.65, 257.35, 257.85, 259.65, 259.75, 
    260.05, 260.15, 259.35, 259.35, 258.25, 258.45, 257.35, 257.25, 257.95, 
    255.95, 255.55, 255.15, 253.95, 254.85, 255.15, 256.15, 254.75, 255.45, 
    253.75, 254.95, 253.25, 251.65, 251.95, 252.15, 252.65, 252.45, 252.05, 
    251.95, 252.75, 253.05, 253.95, 254.85, 254.95, 255.15, 255.95, 256.75, 
    257.85, 258.65, 259.55, 260.85, 261.35, 263.05, 263.55, 263.55, 264.85, 
    265.25, 266.45, 266.95, 267.75, 268.55, 268.45, 267.85, 268.35, 270.25, 
    270.35, 269.75, 270.45, 271.05, 270.75, 270.85, 271.25, 270.85, 271.05, 
    270.65, 271.35, 271.25, 271.35, 271.85, 271.75, 272.05, 272.25, 271.85, 
    272.15, 272.25, 272.15, 271.75, 271.95, 272.15, 272.25, 272.35, 272.25, 
    272.25, 271.95, 271.55, 266.75, 269.25, 269.35, 266.55, 265.55, 266.05, 
    265.45, 265.05, 264.85, 264.05, 263.35, 263.05, 261.75, 261.65, 262.15, 
    261.45, 261.45, 261.55, 260.95, 260.15, 260.45, 261.65, 260.25, 260.65, 
    260.35, 259.75, 259.55, 259.45, 258.65, 258.55, 257.55, 256.65, 256.55, 
    256.35, 255.75, 256.15, 254.35, 255.55, 256.25, 256.35, 255.35, 255.95, 
    256.45, 255.65, 255.65, 255.35, 254.05, 255.55, 252.75, 251.35, 251.55, 
    252.95, 252.05, 251.55, 251.15, 251.05, 250.55, 252.55, 251.55, 250.45, 
    251.85, 251.05, 251.25, 251.65, 251.65, 251.45, 251.15, 250.85, 250.15, 
    250.35, 250.05, 250.65, 250.45, 250.55, 250.65, 250.65, 250.05, 250.85, 
    250.55, 250.35, 251.15, 253.25, 250.75, 250.85, 250.95, 251.65, 250.75, 
    250.25, 249.75, 249.85, 248.75, 249.15, 250.35, 249.65, 249.05, 248.45, 
    248.05, 247.95, 247.85, 247.55, 246.95, 246.25, 245.15, 245.65, 246.05, 
    246.35, 246.45, 246.45, 245.85, 248.45, 246.25, 246.05, 246.25, 246.45, 
    247.55, 247.05, 248.45, 248.25, 248.75, 248.85, 248.65, 248.05, 246.55, 
    244.85, 243.85, 243.85, 243.95, 243.95, 243.25, 244.35, 243.45, 242.95, 
    244.25, 244.45, 244.15, 244.15, 244.25, 244.45, 244.35, 244.25, 243.85, 
    245.45, 245.45, 245.55, 244.85, 243.85, 242.85, 242.75, 243.65, 244.65, 
    244.85, 244.05, 243.35, 243.55, 244.25, 244.65, 244.55, 245.05, 243.95, 
    244.25, 245.05, 244.75, 244.45, 244.65, 244.75, 245.15, 244.85, 244.55, 
    245.35, 245.35, 245.45, 245.55, 245.25, 244.85, 244.65, 244.95, 245.15, 
    245.45, 245.55, 245.35, 246.45, 246.45, 245.65, 246.85, 245.45, 246.65, 
    246.75, 246.45, 246.95, 247.35, 246.45, 246.35, 244.65, 245.05, 245.65, 
    245.25, 247.05, 245.85, 245.15, 246.95, 245.85, 246.35, 246.15, 244.45, 
    244.95, 245.85, 246.45, 245.95, 245.55, 245.45, 246.25, 245.85, 246.05, 
    246.65, 246.85, 246.45, 246.45, 246.65, 245.75, 246.85, 247.85, 248.25, 
    248.85, 249.15, 249.85, 250.35, 250.25, 250.05, 249.45, 249.55, 250.35, 
    250.15, 249.85, 250.25, 250.05, 250.65, 251.25, 252.45, 252.25, 251.65, 
    251.55, 251.55, 250.85, 250.95, 251.55, 251.55, 251.05, 250.55, 250.75, 
    249.95, 249.95, 249.95, 249.95, 249.85, 249.55, 248.95, 248.45, 249.75, 
    248.35, 249.65, 249.35, 249.95, 251.15, 253.85, 254.35, 254.65, 256.55, 
    257.75, 259.25, 260.15, 261.25, 262.85, 263.15, 263.85, 264.55, 264.75, 
    265.55, 265.75, 266.05, 266.35, 266.25, 265.65, 265.65, 265.65, 265.25, 
    265.65, 266.15, 266.65, 267.25, 268.15, 268.75, 269.25, 269.75, 269.95, 
    270.05, 270.05, 270.35, 270.35, 270.15, 270.15, 270.25, 270.35, 270.35, 
    270.35, 270.45, 270.85, 270.75, 270.55, 270.55, 270.75, 270.75, 270.85, 
    270.55, 269.95, 269.05, 268.15, 267.35, 267.15, 267.05, 266.35, 266.55, 
    263.45, 262.75, 262.35, 261.85, 261.55, 261.25, 260.95, 260.65, 260.15, 
    259.55, 259.35, 258.85, 258.45, 258.15, 257.85, 257.65, 257.45, 257.25, 
    257.05, 256.85, 256.75, 256.85, 256.75, 256.85, 257.05, 257.35, 257.75, 
    258.25, 258.85, 259.25, 260.05, 260.85, 261.65, 262.35, 261.85, 261.95, 
    261.65, 261.45, 260.25, 260.35, 260.65, 260.45, 260.75, 261.15, 260.65, 
    259.85, 259.05, 258.25, 257.95, 258.15, 257.75, 257.75, 258.05, 257.35, 
    256.55, 255.95, 255.45, 255.05, 254.85, 254.85, 254.75, 254.45, 254.15, 
    254.45, 254.35, 254.25, 254.25, 254.35, 254.05, 254.15, 254.35, 254.55, 
    254.55, 254.35, 254.35, 254.05, 254.55, 254.75, 254.85, 254.75, 254.55, 
    254.25, 254.25, 254.25, 254.05, 253.85, 253.75, 253.85, 253.65, 253.75, 
    253.35, 253.55, 253.25, 253.15, 253.05, 252.75, 252.75, 252.85, 252.75, 
    252.55, 252.35, 252.45, 251.85, 252.05, 252.05, 252.75, 252.15, 252.15, 
    252.65, 253.15, 252.75, 253.05, 253.05, 252.15, 251.75, 251.85, 252.15, 
    252.35, 252.15, 251.35, 251.05, 251.55, 251.35, 251.05, 250.95, 251.05, 
    250.75, 249.95, 250.05, 250.05, 250.25, 249.15, 248.05, 249.15, 250.25, 
    250.15, 250.45, 249.45, 247.95, 247.85, 247.95, 247.65, 247.65, 248.15, 
    248.85, 248.65, 248.25, 248.45, 248.45, 248.75, 249.15, 249.65, 249.55, 
    249.65, 250.25, 250.75, 251.15, 251.25, 251.05, 250.25, 251.35, 252.05, 
    252.65, 252.95, 252.85, 253.35, 253.55, 253.95, 254.25, 254.55, 252.95, 
    252.75, 253.55, 254.35, 253.85, 253.75, 253.85, 255.15, 254.65, 252.45, 
    252.75, 252.85, 251.55, 250.55, 249.45, 249.25, 248.65, 248.85, 248.65, 
    248.65, 248.45, 247.75, 248.25, 248.35, 248.25, 248.45, 248.55, 248.25, 
    247.95, 247.95, 248.25, 248.55, 249.35, 249.45, 249.75, 249.25, 249.95, 
    250.05, 250.05, 250.05, 249.95, 250.25, 250.85, 250.95, 249.75, 248.25, 
    248.05, 248.05, 247.95, 247.55, 247.55, 248.25, 248.45, 248.35, 248.45, 
    249.55, 249.35, 250.15, 251.65, 252.35, 252.55, 252.25, 252.25, 252.95, 
    253.45, 253.95, 254.75, 255.25, 256.05, 256.75, 257.95, 259.65, 261.35, 
    262.55, 263.45, 264.25, 265.35, 265.45, 267.35, 269.35, 270.05, 270.55, 
    271.25, 272.15, 272.05, 272.55, 272.85, 272.45, 271.85, 271.55, 272.05, 
    272.05, 272.55, 272.85, 272.35, 271.95, 271.25, 270.45, 270.05, 270.15, 
    269.95, 269.85, 269.65, 269.45, 269.65, 269.75, 270.05, 269.45, 270.15, 
    269.95, 270.65, 269.75, 269.55, 270.05, 269.85, 268.75, 268.95, 268.75, 
    268.85, 268.65, 266.35, 264.55, 263.55, 262.55, 261.75, 260.55, 259.75, 
    259.45, 258.85, 257.55, 256.75, 256.55, 256.35, 256.15, 255.95, 255.85, 
    255.85, 256.25, 255.85, 256.05, 256.15, 256.25, 256.15, 256.25, 256.15, 
    255.45, 255.55, 255.85, 256.45, 256.55, 256.55, 256.55, 256.55, 256.45, 
    256.55, 256.85, 256.15, 256.25, 256.55, 256.75, 256.75, 256.75, 256.95, 
    256.95, 256.65, 255.85, 255.15, 254.65, 254.85, 254.85, 254.85, 254.25, 
    254.05, 253.85, 253.75, 253.95, 253.65, 253.65, 252.45, 253.35, 253.25, 
    253.25, 253.25, 253.65, 253.55, 253.65, 253.75, 254.15, 253.75, 253.75, 
    252.95, 253.75, 253.75, 253.55, 253.45, 253.35, 252.95, 252.75, 252.55, 
    252.05, 251.85, 251.75, 251.55, 250.65, 250.65, 251.65, 251.35, 251.75, 
    253.25, 253.45, 252.35, 252.55, 252.85, 253.15, 252.85, 253.05, 253.15, 
    253.15, 254.05, 253.85, 252.45, 253.55, 252.85, 253.15, 253.75, 253.25, 
    252.95, 252.75, 252.95, 252.95, 253.05, 252.55, 251.35, 253.05, 253.25, 
    252.05, 251.55, 252.65, 251.65, 251.45, 252.65, 252.65, 252.35, 252.65, 
    252.55, 252.55, 252.45, 252.95, 252.55, 252.55, 252.95, 253.05, 252.85, 
    252.15, 252.45, 251.95, 252.75, 253.15, 253.05, 253.15, 253.05, 252.75, 
    251.95, 251.85, 251.75, 250.35, 252.15, 252.85, 252.65, 251.95, 253.55, 
    252.65, 253.55, 253.75, 254.15, 253.05, 253.05, 254.35, 253.75, 255.55, 
    254.45, 256.55, 254.75, 261.75, 262.35, 262.85, 263.95, 264.55, 265.05, 
    265.85, 266.35, 266.05, 265.35, 264.55, 264.25, 264.25, 264.35, 264.55, 
    265.25, 265.85, 266.15, 265.75, 265.55, 264.95, 264.65, 264.15, 263.75, 
    263.45, 263.35, 262.65, 262.65, 264.05, 263.45, 263.55, 263.85, 263.05, 
    262.95, 262.85, 262.35, 262.15, 262.55, 263.35, 263.25, 263.35, 261.95, 
    260.85, 259.85, 259.05, 258.95, 258.65, 258.25, 257.85, 257.85, 257.75, 
    257.35, 256.95, 257.35, 257.35, 257.15, 257.05, 257.55, 257.25, 257.15, 
    256.85, 255.95, 255.25, 254.75, 254.45, 253.35, 252.85, 252.95, 252.25, 
    253.35, 252.85, 254.35, 254.55, 253.45, 254.45, 255.55, 256.25, 256.25, 
    255.75, 255.55, 254.75, 255.15, 254.65, 253.55, 253.45, 254.05, 254.25, 
    254.25, 254.45, 254.55, 253.95, 254.25, 254.45, 254.55, 255.65, 254.85, 
    254.35, 254.85, 254.45, 254.55, 253.95, 255.35, 255.25, 254.05, 255.35, 
    255.65, 255.95, 255.75, 255.55, 255.35, 255.15, 255.25, 255.95, 255.45, 
    256.35, 256.65, 257.75, 257.45, 256.15, 254.95, 254.95, 255.25, 255.45, 
    254.95, 254.55, 254.75, 254.95, 254.25, 254.95, 254.75, 255.45, 255.55, 
    256.75, 256.45, 257.15, 257.35, 257.75, 257.85, 257.55, 257.95, 258.95, 
    258.65, 259.35, 260.05, 260.85, 261.05, 261.65, 262.55, 263.25, 263.65, 
    263.75, 264.35, 264.95, 265.45, 265.95, 267.05, 267.65, 267.95, 268.35, 
    269.15, 270.45, 271.35, 271.95, 272.25, 272.35, 272.45, 272.65, 272.75, 
    272.85, 272.75, 275.15, 275.25, 275.25, 275.25, 275.25, 274.25, 274.15, 
    274.15, 274.05, 274.05, 274.05, 274.05, 273.95, 274.05, 274.05, 274.05, 
    274.05, 272.15, 272.05, 271.95, 271.85, 271.85, 271.75, 271.55, 271.45, 
    271.15, 271.15, 271.15, 270.95, 270.55, 270.55, 270.75, 270.85, 270.85, 
    270.75, 270.65, 270.55, 270.45, 270.35, 270.15, 269.45, 267.75, 267.05, 
    266.25, 265.85, 265.25, 264.65, 263.65, 262.65, 261.85, 261.05, 260.55, 
    260.05, 261.95, 261.75, 261.95, 262.45, 263.15, 263.75, 264.55, 265.35, 
    266.15, 266.75, 267.55, 268.05, 268.35, 268.75, 268.95, 269.05, 269.55, 
    269.85, 270.35, 270.65, 270.85, 270.95, 271.25, 271.35, 271.35, 271.35, 
    270.85, 270.85, 270.35, 269.85, 269.15, 269.45, 269.65, 270.05, 270.45, 
    270.95, 269.35, 269.85, 270.05, 270.55, 270.35, 270.45, 270.45, 270.35, 
    270.35, 270.55, 270.75, 270.85, 270.85, 271.15, 271.25, 271.45, 271.55, 
    271.85, 271.25, 271.45, 271.55, 271.75, 271.85, 271.85, 271.75, 271.75, 
    271.75, 271.75, 271.75, 271.65, 271.55, 271.55, 271.45, 271.35, 271.35, 
    271.35, 271.35, 271.45, 271.45, 271.45, 271.55, 271.55, 271.55, 271.55, 
    271.55, 271.45, 271.35, 271.35, 271.05, 270.85, 270.55, 270.25, 269.95, 
    269.65, 269.45, 269.25, 269.15, 269.05, 269.05, 269.05, 269.35, 269.45, 
    269.65, 269.95, 270.05, 269.95, 269.75, 269.55, 269.55, 269.75, 269.85, 
    269.15, 269.25, 269.35, 269.45, 269.45, 269.35, 269.15, 268.75, 268.35, 
    267.85, 267.65, 267.55, 267.35, 267.05, 266.45, 265.75, 265.05, 264.55, 
    263.95, 263.55, 263.45, 263.35, 263.35, 263.35, 263.75, 263.65, 263.55, 
    263.55, 263.45, 263.25, 263.15, 263.05, 262.85, 262.75, 262.55, 262.45, 
    263.45, 263.45, 263.55, 263.65, 263.75, 263.85, 263.75, 263.75, 263.65, 
    263.45, 263.25, 262.85, 261.35, 260.95, 261.05, 261.25, 261.45, 261.65, 
    261.75, 261.75, 261.45, 260.95, 260.65, 260.25, 259.35, 259.45, 259.45, 
    259.45, 259.55, 259.45, 259.25, 258.95, 258.75, 258.55, 258.75, 258.95, 
    255.15, 256.15, 256.85, 257.35, 257.85, 258.15, 258.45, 258.65, 258.75, 
    258.85, 259.05, 259.25, 258.55, 259.45, 259.45, 260.85, 262.45, 263.15, 
    263.65, 263.85, 263.75, 263.65, 263.45, 263.75, 263.85, 263.75, 263.75, 
    264.25, 264.95, 265.05, 265.25, 266.15, 266.95, 268.35, 269.75, 271.55, 
    273.15, 273.45, 273.75, 273.75, 273.55, 273.35, 272.45, 271.95, 271.75, 
    271.65, 272.55, 273.25, 272.65, 272.75, 272.45, 272.25, 271.95, 270.05, 
    268.75, 267.35, 265.25, 263.05, 261.15, 260.25, 260.05, 258.25, 258.35, 
    258.45, 258.35, 258.25, 258.05, 257.95, 257.85, 257.65, 257.55, 257.45, 
    259.45, 259.25, 259.35, 259.45, 259.55, 259.55, 259.45, 259.35, 259.15, 
    259.05, 258.95, 258.85, 258.65, 258.65, 258.75, 258.85, 258.95, 258.75, 
    258.65, 258.45, 258.35, 258.05, 257.65, 257.55, 257.65, 257.85, 257.75, 
    257.65, 257.55, 257.45, 256.65, 255.45, 255.65, 255.35, 255.05, 254.85, 
    254.75, 254.05, 254.05, 254.75, 254.65, 254.65, 254.15, 253.65, 253.35, 
    252.95, 252.75, 252.15, 251.95, 251.25, 251.15, 251.25, 251.35, 251.45, 
    251.55, 251.25, 250.85, 250.65, 250.55, 250.45, 249.95, 249.75, 250.25, 
    250.25, 251.05, 251.35, 251.25, 250.35, 249.65, 248.85, 248.65, 248.35, 
    248.05, 247.85, 247.85, 247.95, 247.85, 248.25, 248.05, 248.05, 248.15, 
    248.25, 248.15, 248.25, 248.85, 249.55, 250.15, 250.75, 250.35, 250.55, 
    250.75, 251.15, 251.05, 250.95, 250.85, 250.85, 250.75, 250.75, 250.85, 
    251.05, 251.15, 251.15, 250.75, 250.65, 250.05, 250.65, 248.85, 249.05, 
    248.75, 248.95, 249.15, 249.95, 249.45, 249.55, 251.05, 250.75, 251.15, 
    249.05, 248.45, 248.25, 248.65, 248.85, 248.55, 249.15, 251.45, 251.65, 
    253.25, 253.45, 248.05, 253.05, 247.45, 247.55, 254.15, 254.65, 254.65, 
    254.95, 254.55, 255.05, 249.45, 253.65, 253.85, 249.15, 253.45, 253.25, 
    246.75, 252.95, 251.25, 246.05, 245.85, 245.85, 245.85, 253.65, 252.65, 
    252.15, 251.85, 246.25, 251.85, 252.35, 252.05, 252.15, 252.55, 252.95, 
    254.25, 255.05, 255.35, 255.05, 254.05, 253.55, 252.55, 251.85, 251.25, 
    250.95, 250.75, 250.65, 250.75, 250.25, 249.85, 249.45, 249.55, 249.55, 
    248.85, 248.25, 247.95, 247.95, 247.95, 247.75, 248.05, 248.45, 248.45, 
    248.35, 248.25, 248.15, 248.05, 247.75, 247.75, 247.55, 248.35, 248.65, 
    248.85, 249.45, 248.85, 248.75, 249.55, 250.85, 253.45, 254.45, 255.05, 
    255.35, 254.55, 255.25, 254.95, 254.55, 255.05, 255.15, 254.85, 254.65, 
    255.35, 255.65, 256.25, 257.15, 258.65, 259.75, 260.95, 262.35, 263.25, 
    264.05, 265.45, 266.55, 266.65, 266.55, 266.85, 267.65, 268.15, 268.55, 
    268.85, 268.45, 268.85, 269.55, 269.45, 270.15, 270.05, 270.35, 270.35, 
    270.55, 270.35, 270.55, 270.65, 270.75, 270.05, 269.75, 269.75, 269.75, 
    270.05, 270.35, 270.45, 269.95, 270.25, 270.55, 270.15, 269.85, 269.85, 
    269.85, 269.55, 269.35, 269.15, 269.75, 269.05, 269.05, 268.85, 269.45, 
    267.65, 268.15, 267.95, 268.15, 268.75, 269.25, 269.05, 269.05, 268.95, 
    267.15, 266.35, 265.75, 265.05, 264.25, 263.75, 262.95, 262.85, 262.75, 
    262.45, 261.95, 261.55, 261.05, 261.15, 260.65, 260.15, 260.65, 259.95, 
    259.55, 259.05, 260.45, 256.65, 256.35, 256.15, 256.05, 255.85, 255.55, 
    255.05, 254.55, 253.95, 253.75, 253.15, 252.75, 252.65, 252.75, 252.75, 
    252.85, 252.95, 253.15, 253.55, 253.95, 254.35, 254.15, 254.35, 254.75, 
    255.15, 255.55, 254.05, 254.95, 255.45, 255.75, 255.55, 255.65, 256.25, 
    257.65, 255.85, 257.95, 258.05, 258.65, 258.85, 258.35, 256.05, 256.15, 
    258.85, 259.25, 259.45, 259.65, 259.55, 260.55, 260.95, 261.25, 259.15, 
    262.15, 262.45, 262.75, 262.35, 259.65, 262.85, 262.55, 261.95, 262.25, 
    260.15, 259.95, 259.15, 257.95, 257.35, 256.65, 256.55, 256.55, 256.75, 
    257.05, 257.25, 257.05, 257.05, 257.45, 257.55, 257.45, 257.55, 257.45, 
    257.35, 257.55, 257.55, 257.55, 257.85, 258.15, 258.55, 258.85, 258.75, 
    258.65, 258.35, 258.25, 258.15, 258.35, 258.65, 258.65, 258.75, 258.35, 
    257.15, 256.45, 256.05, 255.95, 255.55, 255.45, 255.35, 255.05, 254.65, 
    254.35, 253.85, 254.05, 253.15, 252.75, 252.65, 252.55, 252.55, 252.15, 
    251.65, 251.65, 251.45, 251.45, 251.75, 251.85, 251.85, 251.85, _, 
    251.25, 250.85, 250.65, 250.75, 251.05, 251.25, 251.15, 251.25, 250.85, 
    251.25, 251.45, 251.75, 251.95, 252.05, 251.85, 251.35, 251.75, 251.45, 
    251.35, 251.65, 252.45, 252.95, 254.05, 255.85, 257.55, 257.85, 255.85, 
    255.35, 255.85, 255.65, 256.45, 255.35, 255.95, 256.25, 256.55, 258.15, 
    257.55, 257.85, 258.45, 259.35, 259.85, 259.05, 260.65, 260.05, 261.45, 
    262.95, 261.35, 261.05, 260.85, 260.55, 260.25, 260.85, 260.75, 260.25, 
    260.15, 258.35, 257.85, 257.45, 257.25, 257.25, 258.85, 259.15, 257.65, 
    257.55, 258.35, 260.35, 262.25, 261.65, 261.85, 262.45, 264.25, 264.85, 
    265.85, 266.95, 267.85, 268.85, 269.45, 269.45, 269.65, 269.75, 269.85, 
    269.95, 269.95, 270.15, 270.05, 270.35, 270.45, 270.65, 270.75, 271.05, 
    271.15, 270.95, 270.45, 270.55, 270.35, 270.25, 270.05, 269.75, 269.85, 
    270.15, 270.35, 270.35, 270.15, 270.25, 270.35, 270.55, 270.75, 270.85, 
    270.65, 271.05, 271.15, 271.35, 271.25, 270.15, 270.35, 269.75, 269.65, 
    269.75, 269.95, 270.15, 270.15, 270.05, 269.75, 269.85, 269.55, 269.45, 
    269.15, 269.15, 268.95, 268.45, 268.25, 267.95, 267.95, 267.85, 267.85, 
    267.95, 267.95, 267.85, 267.95, 267.55, 267.95, 267.65, 268.55, 269.25, 
    268.25, 267.95, 268.25, 268.15, 268.25, 268.15, 270.15, 270.55, 271.05, 
    271.45, 271.25, 271.15, 270.75, 270.45, 270.35, 270.55, 270.35, 269.75, 
    269.55, 269.75, 269.75, 269.75, 269.25, 268.65, 267.65, 268.65, 269.25, 
    269.05, 268.75, 268.35, 268.65, 268.15, 268.55, 268.15, 268.05, 268.15, 
    268.15, 268.05, 268.15, 268.05, 267.75, 267.35, 267.05, 266.95, 266.65, 
    266.95, 267.35, 267.45, 267.55, 267.55, 267.15, 266.85, 266.55, 266.35, 
    266.25, 266.35, 266.45, 266.65, 266.55, 266.45, 266.45, 266.25, 266.15, 
    266.25, 266.35, 266.25, 266.25, 266.15, 266.15, 266.05, 266.05, 266.15, 
    266.35, 266.15, 265.95, 265.75, 265.85, 265.75, 266.05, 265.95, 266.15, 
    266.15, 266.15, 266.15, 266.35, 266.35, 266.15, 266.35, 266.25, 266.05, 
    265.95, 266.05, 265.85, 265.85, 265.85, 265.75, 265.75, 265.75, 266.45, 
    266.55, 266.55, 266.65, 266.85, 267.05, 267.25, 267.35, 267.55, 267.65, 
    267.75, 267.85, 268.05, 268.25, 268.65, 269.15, 269.75, 270.25, 270.75, 
    271.25, 271.25, 271.35, 271.55, 271.65, 271.15, 271.25, 270.85, 269.95, 
    269.45, 269.25, 268.95, 268.65, 269.25, 268.65, 266.75, 267.65, 267.75, 
    268.05, 268.05, 267.65, 269.55, 270.05, 270.55, 270.95, 271.25, 272.85, 
    272.65, 272.35, 272.35, 272.35, 272.35, 272.35, 272.35, 272.25, 272.35, 
    272.35, 272.45, 272.45, 272.55, 272.65, 272.35, 272.45, 272.55, 272.85, 
    273.05, 273.15, 273.25, 272.25, 271.15, 269.25, 268.25, 266.95, 266.05, 
    266.35, 266.55, 265.65, 266.05, 265.75, 267.25, 266.45, 265.75, 266.15, 
    266.65, 266.45, 266.55, 267.35, 267.75, 268.55, 268.75, 268.95, 268.85, 
    268.85, 269.25, 269.65, 270.05, 270.15, 270.25, 270.35, 270.55, 270.55, 
    270.45, 270.25, 270.05, 269.65, 269.65, 269.25, 269.05, 268.75, 268.85, 
    267.75, 266.75, 264.85, 264.05, 262.55, 261.65, 261.05, 259.95, 259.45, 
    259.35, 259.65, 259.65, 259.65, 259.45, 260.15, 259.75, 258.55, 258.05, 
    258.75, 259.65, 260.75, 262.45, 262.15, 262.55, 262.85, 263.05, 263.05, 
    262.65, 262.85, 263.05, 262.85, 261.45, 261.55, 260.35, 259.85, 260.95, 
    261.85, 260.15, 258.55, 257.95, 256.45, 256.95, 256.95, 257.35, 258.15, 
    257.35, 260.25, 260.65, 261.25, 261.55, 262.05, 262.15, 262.65, 263.05, 
    262.65, 262.65, 262.45, 261.05, 259.45, 259.45, 259.35, 260.95, 260.55, 
    260.35, 260.25, 260.15, 260.15, 260.15, 260.45, 260.65, 261.25, 261.15, 
    261.45, 261.45, 261.75, 262.25, 261.95, 261.95, 261.85, 262.45, 262.95, 
    263.05, 262.95, 262.55, 262.55, 262.55, 262.75, 263.25, 264.05, 263.85, 
    263.55, 262.95, 261.75, 261.55, 261.25, 261.45, 262.95, 262.15, 262.65, 
    261.05, 263.55, 261.05, 261.05, 261.25, 261.15, 261.15, 261.85, 261.75, 
    261.35, 261.55, 260.75, 260.85, 260.65, 260.65, 260.45, 260.25, 259.95, 
    260.65, 260.45, 260.75, 259.55, 261.05, 261.55, 263.25, 263.05, 263.05, 
    262.65, 262.25, 261.85, 262.25, 262.95, 263.35, 262.55, 262.45, 262.65, 
    262.65, 262.65, 262.85, 262.25, 261.55, 261.35, 261.95, 261.35, 260.95, 
    261.15, 261.65, 261.55, 261.45, 261.65, 261.95, 261.85, 261.95, 261.55, 
    261.65, 261.75, 261.55, 261.25, 261.15, 260.95, 261.05, 261.05, 261.95, 
    262.55, 262.25, 262.45, 262.45, 262.35, 261.85, 261.65, 260.85, 260.55, 
    260.35, 259.95, 259.65, 259.55, 259.25, 259.25, 259.35, 259.55, 259.55, 
    259.55, 259.95, 259.95, 259.85, 259.95, 260.15, 259.95, 259.65, 259.85, 
    259.85, 259.75, 259.45, 259.05, 258.75, 258.55, 258.35, 258.15, 258.05, 
    258.45, 258.45, 258.65, 259.05, 260.75, 260.35, 260.15, 260.05, 260.55, 
    260.45, 259.85, 259.95, 261.25, 263.25, 262.25, 262.85, 263.45, 263.35, 
    263.65, 263.25, 262.35, 261.45, 260.85, 260.25, 259.45, 259.55, 258.35, 
    258.25, 258.95, 257.15, 258.35, 259.55, 260.65, 261.75, 261.55, 263.75, 
    261.25, 262.45, 261.15, 260.35, 261.25, 261.35, 260.95, 261.05, 261.05, 
    260.45, 259.85, 260.35, 260.55, 261.55, 261.65, 262.05, 262.15, 261.95, 
    262.35, 261.25, 261.15, 260.75, 261.25, 262.15, 261.15, 261.15, 260.95, 
    265.45, 265.65, 265.85, 265.75, 267.25, 265.75, 265.85, 265.15, 263.95, 
    263.35, 261.95, 263.35, 263.55, 263.55, 263.45, 263.55, 263.35, 262.45, 
    262.05, 259.75, 259.25, 258.25, 257.75, 257.35, 258.75, 259.25, 259.65, 
    260.25, 260.65, 260.75, 261.05, 260.95, 260.95, 260.65, 260.65, 259.15, 
    258.25, 258.35, 258.75, 260.65, 260.85, 261.25, 261.25, 261.05, 261.55, 
    261.75, 262.05, 262.65, 263.55, 263.25, 263.65, 264.15, 264.35, 265.25, 
    265.35, 265.55, 265.65, 265.95, 266.25, 266.75, 266.55, 267.05, 267.65, 
    268.15, 268.45, 268.75, 268.85, 269.15, 268.65, 269.25, 269.45, 269.05, 
    269.25, 269.55, 269.85, 269.75, 269.75, 269.95, 269.45, 269.05, 268.85, 
    268.75, 268.45, 267.95, 267.45, 266.95, 266.85, 266.55, 266.45, 266.45, 
    266.35, 266.15, 265.65, 265.35, 265.85, 266.25, 266.05, 265.95, 265.65, 
    265.55, 265.55, 265.45, 265.35, 265.15, 265.05, 264.65, 264.25, 263.75, 
    263.25, 262.45, 261.75, 262.25, 261.85, 261.85, 261.45, 260.25, 259.95, 
    260.65, 262.15, 260.45, 259.95, 261.05, 262.05, 261.45, 261.15, 260.15, 
    260.95, 259.75, 259.95, 259.85, 260.35, 260.25, 261.15, 261.15, 261.75, 
    263.35, 263.75, 264.35, 264.65, 264.65, 264.25, 264.65, 264.95, 265.15, 
    265.25, 265.55, 265.75, 265.65, 264.65, 264.15, 263.95, 263.55, 264.05, 
    263.45, 262.45, 262.25, 261.85, 261.25, 260.95, 260.75, 260.65, 260.35, 
    262.15, 261.85, 261.55, 261.65, 261.85, 262.75, 263.05, 263.85, 263.55, 
    263.15, 264.05, 263.85, 264.05, 264.05, 263.75, 263.35, 262.85, 262.15, 
    261.65, 261.25, 260.95, 261.25, 259.75, 259.55, 259.75, 261.05, 260.15, 
    260.35, 260.65, 260.65, 260.65, 260.85, 261.45, 261.15, 261.35, 260.75, 
    260.65, 260.95, 259.95, 259.25, 258.85, 258.25, 258.15, 257.85, 258.05, 
    258.65, 258.05, 258.15, 258.85, 258.75, 258.95, 259.85, 259.75, 260.15, 
    260.65, 260.75, 260.75, 261.05, 261.25, 261.45, 261.05, 260.55, 260.15, 
    259.65, 258.95, 257.25, 257.45, 257.55, 257.75, 257.65, 257.65, 258.55, 
    258.95, 259.05, 259.15, 259.55, 259.25, 259.55, 260.25, 259.95, 261.15, 
    261.55, 260.05, 260.55, 260.35, 260.25, 260.35, 259.95, 259.85, 259.75, 
    259.85, 259.65, 259.85, 259.85, 259.95, 259.85, 260.45, 259.95, 260.55, 
    260.95, 261.45, 261.75, 262.35, 262.15, 262.65, 262.65, 262.75, 262.55, 
    263.05, 263.25, 263.65, 264.15, 264.25, 264.35, 264.25, 264.35, 264.65, 
    264.85, 265.05, 264.55, 264.45, 264.55, 265.05, 265.35, 265.15, 265.65, 
    266.45, 266.35, 266.55, 267.05, 266.55, 266.05, 265.75, 266.45, 267.65, 
    268.95, 269.35, 269.85, 269.75, 269.85, 270.05, 270.45, 269.75, 269.85, 
    268.75, 266.75, 265.55, 264.65, 263.95, 263.45, 263.15, 262.45, 262.35, 
    262.05, 261.95, 262.35, 262.35, 262.05, 262.55, 262.25, 262.45, 262.35, 
    262.55, 262.95, 263.25, 263.45, 263.35, 263.25, 263.85, 264.45, 264.65, 
    264.75, 265.25, 265.55, 265.95, 266.65, 267.05, 266.85, 267.15, 267.15, 
    267.15, 266.85, 266.95, 266.95, 267.05, 267.35, 267.75, 269.15, 270.15, 
    270.45, 270.65, 270.95, 271.15, 271.45, 271.85, 272.15, 272.15, 272.15, 
    272.25, 272.15, 271.85, 271.75, 271.55, 271.65, 272.15, 272.45, 272.45, 
    272.55, 272.55, 272.45, 272.45, 272.55, 272.35, 272.45, 272.75, 272.95, 
    273.05, 273.05, 273.25, 273.15, 272.85, 272.95, 273.35, 273.45, 274.15, 
    273.45, 273.25, 273.15, 274.05, 272.95, 273.15, 272.55, 273.05, 273.35, 
    273.25, 273.45, 273.75, 273.35, 273.55, 273.25, 273.45, 273.65, 274.15, 
    273.95, 274.15, 273.75, 274.05, 274.05, 274.35, 274.25, 273.55, 274.05, 
    273.55, 273.75, 273.55, 273.65, 273.45, 273.55, 273.75, 273.35, 273.85, 
    273.95, 273.85, 273.85, 273.65, 274.65, 273.95, 273.65, 273.45, 274.55, 
    273.75, 273.45, 273.15, 271.55, 270.85, 269.65, 269.25, 268.85, 268.55, 
    268.05, 267.75, 267.45, 267.15, 266.85, 266.55, 266.05, 265.65, 265.55, 
    265.55, 265.55, 265.35, 265.45, 265.45, 265.25, 265.15, 264.55, 264.35, 
    264.55, 264.25, 264.15, 263.95, 263.85, 264.25, 263.95, 263.75, 263.95, 
    263.75, 263.75, 263.85, 265.05, 265.25, 265.25, 265.65, 265.65, 265.55, 
    266.05, 266.25, 266.35, 266.55, 266.75, 266.95, 267.05, 267.05, 267.25, 
    267.25, 266.75, 267.35, 267.65, 268.45, 269.15, 269.75, 269.55, 269.45, 
    269.75, 269.65, 269.55, 269.45, 269.45, 269.25, 269.25, 269.25, 269.15, 
    268.85, 269.05, 269.05, 269.35, 269.65, 270.15, 269.85, 270.15, 270.15, 
    270.45, 270.15, 270.15, 270.15, 270.75, 270.75, 270.55, 270.35, 270.15, 
    270.15, 269.45, 269.05, 268.95, 268.95, 268.85, 268.95, 269.05, 269.25, 
    269.45, 269.75, 269.65, 270.15, 270.85, 270.55, 270.75, 270.55, 270.55, 
    270.05, 269.95, 269.65, 269.55, 269.65, 269.75, 269.85, 269.95, 270.05, 
    270.15, 270.25, 270.35, 270.55, 271.05, 271.35, 271.65, 271.85, 272.95, 
    273.65, 273.45, 273.85, 273.45, 272.95, 273.05, 273.85, 274.15, 272.25, 
    271.95, 271.85, 271.15, 270.55, 269.25, 269.35, 269.05, 268.75, 268.45, 
    268.55, 268.65, 268.75, 269.05, 269.05, 268.95, 269.45, 269.95, 269.65, 
    269.15, 268.75, 268.75, 269.35, 269.25, 269.05, 268.65, 268.15, 268.65, 
    268.75, 269.35, 269.65, 269.95, 270.15, 270.85, 270.75, 270.65, 270.55, 
    270.45, 270.65, 270.95, 271.35, 271.75, 271.65, 271.65, 271.55, 271.55, 
    271.45, 271.45, 271.45, 271.85, 271.45, 271.65, 271.25, 271.15, 270.75, 
    270.55, 270.45, 269.95, 269.05, 268.95, 268.75, 269.15, 269.75, 270.25, 
    270.55, 270.45, 270.25, 270.35, 270.55, 270.85, 271.05, 271.35, 271.35, 
    271.35, 271.15, 271.15, 271.15, 271.05, 270.85, 270.55, 270.65, 270.65, 
    270.75, 270.85, 271.05, 271.35, 271.75, 272.05, 272.35, 272.85, 273.35, 
    273.25, 273.25, 273.15, 273.15, 273.05, 272.95, 272.95, 272.75, 272.85, 
    272.55, 272.25, 272.25, 272.25, 272.25, 272.35, 272.25, 272.45, 272.65, 
    272.75, 272.45, 272.75, 272.55, 272.65, 272.55, 272.45, 272.35, 272.15, 
    271.95, 271.95, 271.75, 271.55, 271.65, 271.65, 271.55, 271.45, 271.35, 
    271.15, 271.15, 271.05, 270.95, 270.95, 270.85, 271.05, 271.15, 271.45, 
    271.65, 271.85, 272.15, 272.05, 272.05, 271.95, 271.75, 271.65, 271.75, 
    271.85, 271.85, 271.85, 271.85, 271.85, 271.95, 272.05, 272.05, 272.05, 
    271.95, 272.05, 272.25, 272.55, 272.75, 272.65, 272.75, 272.95, 273.65, 
    273.35, 272.95, 272.95, 272.85, 272.85, 272.95, 272.85, 272.75, 272.75, 
    272.75, 272.75, 272.65, 272.45, 272.45, 272.45, 272.65, 272.95, 272.95, 
    273.05, 273.15, 273.05, 273.05, 273.15, 273.05, 273.05, 272.95, 272.85, 
    272.65, 272.45, 272.15, 272.15, 272.25, 272.35, 272.35, 272.35, 272.25, 
    272.45, 272.55, 272.65, 272.55, 272.75, 272.75, 272.85, 272.75, 272.75, 
    272.75, 272.75, 272.75, 272.65, 272.55, 272.65, 272.35, 272.45, 272.35, 
    271.55, 271.95, 271.55, 271.75, 272.05, 271.35, 271.25, 271.45, 271.05, 
    270.95, 270.95, 270.95, 270.85, 270.85, 270.75, 270.85, 270.55, 270.25, 
    269.95, 270.35, 270.25, 269.85, 269.75, 270.05, 270.25, 270.05, 270.75, 
    270.05, 270.35, 270.35, 271.05, 270.55, 270.45, 270.35, 270.95, 271.65, 
    271.45, 271.35, 271.85, 272.05, 271.95, 271.95, 270.95, 270.95, 270.85, 
    270.55, 271.35, 271.85, 271.85, 271.95, 271.75, 272.05, 272.55, 272.75, 
    272.85, 272.95, 272.85, 272.95, 273.05, 273.15, 273.25, 273.35, 273.45, 
    273.45, 273.55, 273.75, 273.95, 274.05, 274.15, 273.95, 273.65, 273.55, 
    273.35, 273.25, 273.35, 273.35, 273.45, 273.95, 273.95, 274.25, 274.15, 
    273.95, 274.45, 274.35, 273.85, 273.95, 274.45, 275.25, 273.85, 273.65, 
    274.35, 274.85, 272.95, 272.85, 274.25, 272.65, 272.55, 273.05, 273.55, 
    276.05, 276.15, 275.25, 273.75, 273.85, 273.95, 273.15, 272.65, 272.55, 
    272.25, 271.85, 271.45, 271.25, 271.55, 271.85, 272.25, 272.75, 272.95, 
    273.05, 273.05, 273.05, 273.05, 273.15, 273.15, 273.15, 273.05, 272.95, 
    273.15, 272.95, 273.15, 272.95, 273.25, 273.85, 273.85, 273.75, 273.75, 
    273.85, 274.15, 274.45, 274.85, 274.75, 274.45, 274.25, 274.25, 274.15, 
    274.25, 274.45, 274.35, 274.55, 274.95, 274.85, 275.35, 275.75, 276.25, 
    276.45, 276.85, 276.15, 276.35, 275.25, 274.85, 274.85, 274.55, 274.35, 
    274.35, 274.15, 274.15, 274.05, 273.95, 273.55, 273.45, 273.55, 273.35, 
    273.65, 273.65, 273.35, 273.55, 273.25, 273.75, 274.25, 274.15, 274.15, 
    273.95, 274.35, 274.55, 274.75, 274.55, 274.95, 274.75, 274.35, 274.45, 
    274.75, 274.45, 273.35, 272.75, 272.95, 273.45, 273.75, 273.45, 273.65, 
    274.05, 273.75, 273.75, 273.65, 273.35, 273.85, 273.45, 274.55, 274.55, 
    273.85, 274.35, 273.25, 273.15, 273.65, 273.35, 272.55, 272.25, 271.45, 
    271.65, 271.45, 271.65, 271.95, 272.15, 272.75, 272.25, 272.15, 272.55, 
    272.15, 272.15, 272.25, 272.25, 272.15, 272.15, 272.55, 272.75, 272.85, 
    272.85, 272.85, 272.85, 272.85, 272.85, 272.65, 272.75, 272.85, 272.85, 
    272.85, 272.85, 272.75, 272.95, 273.05, 273.05, 273.05, 273.05, 272.95, 
    272.85, 273.05, 273.05, 273.05, 273.15, 273.15, 273.05, 273.15, 273.05, 
    272.95, 272.95, 273.05, 272.95, 272.95, 272.95, 273.05, 272.95, 272.75, 
    272.85, 272.85, 272.95, 273.05, 273.45, 273.95, 273.75, 273.75, 273.55, 
    273.55, 273.25, 273.15, 273.75, 273.55, 273.25, 273.45, 273.35, 273.35, 
    273.05, 272.85, 273.05, 273.05, 273.15, 273.45, 273.55, 273.85, 273.55, 
    274.05, 273.75, 273.35, 273.15, 273.25, 273.15, 273.35, 274.65, 273.45, 
    272.45, 272.25, 271.75, 271.85, 271.45, 271.45, 271.25, 271.65, 271.95, 
    274.05, 272.95, 273.35, 273.95, 272.75, 274.95, 277.45, 274.55, 274.45, 
    274.05, 274.65, 275.25, 276.45, 274.85, 273.05, 272.25, 272.15, 272.45, 
    272.25, 271.45, 271.25, 271.15, 270.75, 270.55, 270.45, 270.45, 270.15, 
    270.15, 269.95, 269.55, 269.95, 269.75, 270.05, 270.05, 270.15, 270.55, 
    270.65, 270.15, 270.35, 270.55, 270.35, 270.55, 270.05, 269.85, 270.35, 
    270.25, 270.65, 270.85, 270.85, 270.95, 271.45, 271.15, 270.75, 271.15, 
    270.15, 270.25, 270.35, 270.45, 270.45, 270.85, 270.85, 271.15, 271.35, 
    271.65, 272.45, 273.05, 272.55, 272.65, 272.95, 272.95, 272.95, 272.95, 
    273.05, 273.05, 272.95, 272.95, 272.95, 272.95, 274.25, 274.05, 272.95, 
    272.95, 273.45, 273.45, 273.15, 273.05, 273.05, 273.15, 272.65, 271.75, 
    271.45, 271.55, 271.75, 271.85, 272.15, 272.25, 272.65, 272.85, 273.05, 
    273.15, 273.05, 273.05, 273.15, 273.15, 273.05, 273.15, 273.15, 273.15, 
    273.45, 273.55, 273.65, 273.65, 273.75, 274.25, 274.45, 274.05, 274.05, 
    274.05, 273.85, 274.15, 272.95, 273.15, 272.95, 272.85, 272.85, 272.95, 
    273.35, 273.95, 273.75, 274.25, 274.35, 274.25, 274.35, 273.95, 275.15, 
    275.55, 274.85, 274.25, 274.05, 273.85, 274.05, 274.15, 274.25, 274.25, 
    274.15, 273.65, 274.25, 273.95, 273.75, 273.85, 273.45, 273.55, 273.95, 
    273.55, 273.45, 273.25, 273.25, 273.25, 273.85, 273.95, 273.55, 272.95, 
    272.85, 273.05, 273.45, 273.15, 272.95, 272.55, 272.45, 272.25, 272.25, 
    272.25, 272.25, 272.25, 272.45, 272.35, 272.35, 272.35, 272.35, 272.35, 
    272.65, 273.15, 272.95, 273.05, 273.95, 274.25, 273.95, 273.25, 273.45, 
    273.65, 273.05, 273.75, 273.25, 273.55, 273.45, 273.35, 273.55, 273.55, 
    273.35, 273.25, 273.75, 274.15, 274.15, 273.25, 273.55, 273.45, 273.35, 
    273.15, 272.75, 272.65, 272.55, 272.55, 272.45, 272.35, 272.55, 272.55, 
    272.95, 272.65, 272.95, 272.75, 272.65, 272.65, 272.65, 272.65, 272.75, 
    272.75, 272.85, 272.85, 272.85, 272.85, 272.95, 272.95, 272.85, 272.85, 
    272.65, 272.65, 272.85, 272.95, 272.55, 272.45, 272.45, 272.55, 272.65, 
    272.75, 272.85, 272.75, 272.85, 273.25, 273.25, 274.15, 273.55, 273.65, 
    273.55, 273.45, 273.85, 273.85, 273.45, 272.95, 272.75, 272.95, 273.25, 
    273.55, 273.25, 272.55, 272.45, 272.45, 271.95, 271.85, 271.85, 271.65, 
    273.15, 273.05, 273.95, 274.75, 275.25, 275.35, 276.15, 276.55, 275.95, 
    277.15, 275.55, 274.65, 275.35, 276.15, 275.55, 274.45, 275.75, 276.35, 
    273.95, 274.25, 275.15, 275.55, 274.75, 274.95, 274.85, 274.35, 274.45, 
    274.45, 275.05, 275.95, 276.55, 275.85, 275.95, 276.15, 276.35, 275.55, 
    275.05, 274.85, 274.15, 274.35, 273.85, 273.95, 273.75, 273.45, 273.25, 
    272.85, 272.85, 272.65, 272.55, 273.25, 272.95, 273.35, 273.25, 273.55, 
    273.35, 273.35, 273.35, 273.35, 273.25, 273.15, 273.25, 273.35, 273.25, 
    273.05, 272.95, 272.75, 272.65, 272.85, 272.55, 272.65, 272.55, 272.65, 
    272.75, 272.85, 272.95, 272.95, 273.15, 273.35, 273.85, 274.25, 274.35, 
    274.15, 273.45, 273.65, 273.45, 273.45, 273.95, 273.85, 274.25, 273.05, 
    273.65, 273.15, 272.65, 272.65, 272.95, 274.05, 274.35, 273.45, 273.25, 
    273.45, 273.45, 275.15, 275.35, 275.75, 277.45, 275.65, 273.45, 274.35, 
    272.35, 272.05, 272.05, 272.35, 272.35, 272.95, 272.85, 272.75, 273.85, 
    272.75, 273.15, 273.05, 273.05, 272.95, 272.85, 272.25, 272.15, 272.55, 
    272.95, 272.85, 273.45, 273.45, 273.45, 273.35, 273.25, 272.85, 272.55, 
    272.25, 272.05, 271.85, 271.95, 271.95, 271.85, 271.75, 271.95, 272.25, 
    272.25, 272.35, 272.65, 272.55, 272.85, 272.75, 272.75, 272.75, 272.85, 
    272.85, 273.75, 274.15, 274.45, 274.85, 275.15, 274.85, 274.45, 275.85, 
    274.95, 274.25, 273.55, 274.25, 274.75, 275.05, 274.95, 274.25, 273.95, 
    273.75, 273.75, 275.75, 274.15, 274.25, 274.35, 274.65, 274.55, 273.95, 
    273.45, 273.35, 273.15, 272.95, 273.55, 274.95, 274.75, 274.45, 274.05, 
    273.65, 273.25, 272.95, 272.55, 272.75, 272.75, 273.05, 273.45, 273.55, 
    273.55, 273.45, 273.25, 273.15, 273.15, 272.95, 273.15, 273.05, 273.05, 
    272.95, 272.95, 273.05, 273.05, 273.15, 273.15, 273.05, 273.05, 273.05, 
    272.95, 272.85, 272.85, 272.75, 272.75, 272.95, 273.05, 273.25, 273.45, 
    273.45, 273.75, 273.65, 273.45, 273.75, 273.15, 273.15, 272.95, 272.75, 
    272.65, 272.45, 272.25, 272.15, 272.35, 272.75, 273.25, 273.75, 276.25, 
    274.25, 274.35, 274.65, 275.55, 275.15, 274.85, 274.95, 274.95, 274.95, 
    274.85, 274.65, 274.45, 274.25, 273.75, 273.15, 273.05, 273.55, 273.05, 
    272.65, 272.15, 271.75, 274.15, 273.05, 273.55, 273.45, 273.75, 274.95, 
    274.65, 275.25, 274.85, 275.85, 275.15, 275.05, 275.15, 274.85, 274.65, 
    274.85, 274.45, 274.45, 274.15, 273.05, 273.35, 274.95, 274.65, 274.85, 
    275.35, 275.75, 276.15, 274.95, 274.95, 274.85, 275.35, 275.45, 274.95, 
    275.25, 275.05, 274.95, 275.45, 275.15, 275.05, 275.45, 275.45, 275.15, 
    274.45, 274.45, 274.85, 275.95, 274.75, 273.35, 273.45, 273.35, 273.05, 
    272.75, 273.15, 272.65, 273.05, 273.25, 273.65, 273.85, 273.95, 274.05, 
    273.65, 273.45, 273.55, 273.55, 273.45, 273.45, 273.45, 273.35, 273.35, 
    273.35, 273.55, 273.55, 272.75, 272.75, 273.25, 273.35, 273.25, 273.15, 
    273.25, 273.25, 273.35, 273.35, 273.15, 272.95, 272.75, 272.75, 272.95, 
    273.35, 273.65, 273.75, 273.35, 273.05, 272.65, 272.95, 272.85, 272.95, 
    273.15, 273.35, 274.05, 275.95, 275.85, 275.75, 275.75, 275.85, 275.45, 
    274.85, 275.55, 275.65, 275.65, 276.35, 275.55, 274.75, 274.55, 274.95, 
    276.15, 278.35, 274.15, 273.85, 273.95, 274.05, 274.05, 274.25, 273.75, 
    274.15, 274.25, 274.05, 274.15, 275.15, 275.15, 274.95, 274.65, 274.75, 
    274.35, 274.05, 273.85, 273.65, 272.75, 272.85, 272.95, 273.35, 273.45, 
    273.75, 274.15, 274.75, 274.65, 275.25, 275.75, 275.25, 275.55, 275.35, 
    273.95, 275.95, 275.95, 276.75, 276.45, 275.75, 274.65, 275.65, 276.55, 
    276.45, 276.25, 275.85, 275.35, 275.85, 275.25, 276.05, 275.45, 275.35, 
    275.35, 274.95, 276.65, 276.25, 276.75, 276.25, 275.15, 275.15, 276.35, 
    275.75, 276.25, 275.25, 274.75, 274.65, 277.35, 278.45, 278.65, 278.65, 
    275.65, 276.25, 276.85, 276.35, 274.95, 278.95, 278.35, 278.55, 277.85, 
    275.25, 278.25, 275.25, 277.65, 274.75, 275.85, 274.05, 274.05, 274.55, 
    273.95, 273.55, 273.75, 274.45, 273.75, 273.85, 273.55, 273.55, 273.55, 
    273.65, 273.65, 273.45, 273.45, 273.55, 273.75, 273.85, 274.05, 273.95, 
    274.15, 274.35, 274.25, 274.65, 274.55, 274.25, 274.45, 274.35, 274.15, 
    273.85, 273.75, 273.65, 273.65, 273.65, 273.65, 273.75, 273.75, 273.75, 
    273.55, 273.65, 273.85, 273.95, 273.95, 274.15, 274.35, 274.05, 273.65, 
    273.65, 273.65, 273.65, 273.55, 273.35, 273.35, 273.25, 273.25, 273.25, 
    273.35, 273.45, 273.45, 273.45, 273.45, 273.45, 273.55, 273.65, 273.85, 
    274.55, 275.05, 275.85, 276.45, 275.85, 274.85, 275.35, 274.65, 275.15, 
    275.95, 276.45, 276.25, 276.15, 275.95, 275.95, 275.75, 275.65, 275.45, 
    275.45, 275.45, 275.35, 275.35, 275.35, 275.25, 275.15, 275.15, 275.05, 
    275.35, 275.25, 274.85, 274.55, 274.75, 274.55, 274.35, 274.25, 274.15, 
    274.05, 273.65, 273.85, 274.05, 274.05, 274.45, 274.85, 274.85, 274.95, 
    275.15, 275.05, 275.25, 275.15, 274.95, 275.05, 274.95, 275.25, 275.75, 
    275.45, 275.25, 275.95, 275.85, 275.05, 275.25, 275.45, 275.45, 275.25, 
    274.95, 274.45, 274.05, 274.15, 274.15, 273.65, 273.35, 273.75, 273.85, 
    273.85, 273.75, 274.05, 274.45, 274.45, 274.15, 274.15, 274.85, 274.75, 
    274.65, 275.05, 274.45, 273.45, 273.15, 274.05, 273.75, 273.45, 272.85, 
    272.65, 272.75, 273.15, 273.65, 273.95, 274.45, 275.05, 276.75, 274.35, 
    274.55, 274.75, 273.15, 273.15, 273.85, 274.25, 274.55, 274.75, 274.85, 
    274.95, 275.25, 275.25, 275.45, 275.45, 275.65, 275.85, 276.25, 276.05, 
    275.55, 274.95, 274.65, 274.85, 275.15, 275.25, 275.35, 275.15, 275.15, 
    275.35, 275.05, 275.55, 275.05, 275.05, 274.85, 275.45, 275.05, 275.25, 
    275.25, 276.35, 275.75, 276.65, 275.55, 275.95, 276.95, 275.45, 276.45, 
    276.45, 275.85, 275.95, 276.55, 277.35, 278.05, 278.15, 277.15, 277.85, 
    277.75, 277.75, 278.35, 277.85, 277.55, 278.05, 278.85, 279.35, 279.75, 
    280.05, 279.15, 279.45, 279.65, 279.25, 279.75, 280.55, 280.55, 279.85, 
    279.35, 279.95, 279.55, 279.95, 280.25, 280.25, 280.25, 280.05, 279.75, 
    279.45, 278.95, 279.25, 279.55, 279.75, 279.95, 279.85, 279.95, 280.25, 
    280.85, 281.55, 281.75, 281.45, 281.35, 281.35, 281.25, 281.15, 281.05, 
    281.05, 280.95, 280.35, 280.85, 280.85, 280.65, 280.05, 280.35, 279.85, 
    279.55, 279.95, 280.25, 280.65, 281.15, 281.55, 282.05, 282.45, 281.85, 
    281.45, 282.15, 282.85, 283.35, 282.95, 281.45, 282.85, 282.25, 279.65, 
    280.45, 280.85, 281.15, 281.45, 281.65, 278.35, 277.85, 278.35, 278.75, 
    278.85, 278.95, 279.15, 279.25, 279.45, 279.75, 280.35, 280.85, 281.35, 
    281.85, 282.25, 282.35, 281.35, 280.25, 280.85, 280.55, 282.05, 282.85, 
    282.45, 281.95, 282.85, 282.55, 282.35, 281.85, 280.55, 279.05, 277.35, 
    278.05, 278.05, 278.05, 278.25, 277.95, 279.35, 278.05, 278.25, 278.35, 
    277.35, 277.15, 276.95, 276.75, 276.55, 276.35, 276.05, 275.85, 275.85, 
    275.65, 275.35, 275.45, 276.05, 275.75, 275.55, 275.95, 276.45, 276.85, 
    277.05, 277.85, 277.25, 276.55, 276.55, 276.95, 276.95, 276.95, 276.95, 
    277.05, 277.15, 277.35, 277.35, 277.15, 276.95, 276.75, 276.45, 276.75, 
    277.15, 277.75, 277.75, 277.75, 277.75, 277.35, 277.65, 277.95, 278.05, 
    278.35, 278.85, 279.05, 278.95, 279.15, 279.15, 280.15, 279.55, 279.75, 
    279.55, 279.45, 279.05, 278.65, 278.15, 277.15, 277.05, 276.25, 276.15, 
    276.25, 276.25, 276.75, 276.65, 276.85, 276.85, 277.75, 277.55, 277.55, 
    277.65, 277.55, 277.35, 277.55, 277.45, 277.25, 278.25, 277.85, 278.15, 
    278.35, 277.45, 277.05, 276.65, 277.25, 276.85, 276.45, 276.15, 276.15, 
    276.45, 276.95, 277.05, 276.95, 276.95, 277.45, 277.35, 277.25, 277.15, 
    277.05, 277.05, 276.15, 278.35, 278.65, 278.25, 277.65, 277.35, 277.35, 
    277.55, 277.65, 277.45, 277.25, 277.45, 279.05, 278.25, 279.05, 278.15, 
    278.35, 277.75, 277.85, 278.75, 278.25, 277.65, 278.25, 278.05, 277.35, 
    277.35, 277.45, 277.35, 277.75, 278.05, 277.35, 277.25, 277.45, 277.85, 
    278.75, 278.75, 278.35, 278.45, 278.45, 278.35, 278.35, 278.55, 279.05, 
    278.75, 279.15, 279.25, 278.35, 276.85, 276.75, 278.15, 277.15, 276.35, 
    276.15, 276.75, 276.95, 277.05, 277.05, 277.05, 277.05, 277.45, 277.35, 
    277.45, 277.35, 277.25, 277.25, 277.25, 277.25, 276.85, 276.95, 276.75, 
    276.75, 276.35, 276.25, 276.15, 275.75, 275.95, 275.55, 275.45, 275.55, 
    275.85, 275.95, 276.25, 276.15, 275.85, 274.95, 276.35, 276.25, 276.25, 
    276.55, 276.45, 276.65, 276.45, 276.85, 276.75, 276.65, 276.35, 276.35, 
    276.25, 276.45, 276.75, 277.35, 277.55, 277.55, 277.45, 277.55, 277.45, 
    277.25, 277.25, 277.15, 277.25, 276.75, 276.75, 276.95, 277.65, 277.85, 
    278.25, 276.75, 276.85, 276.75, 277.25, 275.85, 276.75, 276.45, 276.25, 
    276.15, 276.25, 276.25, 275.95, 276.25, 276.35, 276.85, 276.75, 276.45, 
    276.25, 276.35, 276.55, 276.65, 276.25, 275.75, 275.75, 275.85, 275.75, 
    275.35, 275.25, 275.25, 274.85, 274.45, 274.45, 274.95, 275.25, 275.35, 
    275.25, 275.35, 275.25, 275.25, 275.25, 274.85, 274.05, 274.05, 274.05, 
    274.05, 275.05, 274.95, 274.95, 274.85, 274.55, 274.45, 274.15, 273.65, 
    273.15, 272.85, 272.55, 272.45, 272.45, 272.55, 272.65, 272.75, 272.75, 
    272.85, 273.55, 274.25, 274.25, 274.25, 274.25, 274.45, 274.15, 274.45, 
    274.25, 274.15, 274.05, 274.05, 274.05, 274.15, 274.05, 274.05, 274.05, 
    274.05, 273.45, 273.65, 273.75, 274.05, 274.25, 274.35, 274.75, 275.05, 
    275.25, 275.45, 275.95, 276.35, 276.65, 276.85, 277.05, 277.05, 276.85, 
    277.15, 278.25, 276.55, 277.25, 277.45, 276.95, 277.25, 276.75, 275.85, 
    276.55, 276.55, 276.25, 277.55, 277.95, 278.65, 278.15, 277.25, 276.65, 
    276.25, 276.35, 276.65, 276.65, 276.55, 276.15, 276.25, 275.85, 275.55, 
    275.85, 275.65, 276.25, 275.85, 275.85, 275.75, 275.55, 275.35, 275.65, 
    275.65, 275.65, 275.85, 275.65, 275.85, 275.65, 275.35, 275.95, 275.95, 
    275.75, 275.45, 275.75, 276.55, 277.25, 277.45, 277.55, 276.75, 276.65, 
    277.15, 276.55, 275.65, 276.25, 275.85, 276.95, 276.25, 277.55, 275.65, 
    278.05, 277.45, 277.75, 277.55, 277.45, 277.15, 277.15, 277.65, 277.15, 
    276.45, 276.35, 276.55, 277.05, 276.65, 276.45, 276.35, 276.15, 275.75, 
    275.75, 275.95, 276.05, 275.45, 275.35, 275.45, 275.35, 275.15, 275.35, 
    275.55, 275.15, 275.35, 275.45, 275.35, 275.25, 274.75, 274.55, 274.45, 
    274.35, 274.15, 273.95, 273.85, 273.65, 273.75, 273.55, 273.85, 273.45, 
    273.45, 273.25, 273.45, 273.65, 273.95, 273.75, 273.75, 273.75, 273.85, 
    273.95, 274.25, 273.85, 273.55, 273.35, 273.05, 272.95, 272.85, 272.65, 
    272.55, 272.65, 272.85, 273.15, 272.75, 272.65, 272.75, 272.75, 273.05, 
    272.95, 273.15, 274.05, 273.95, 274.05, 274.35, 274.05, 274.25, 274.05, 
    273.85, 273.75, 273.25, 272.55, 272.25, 272.15, 271.65, 271.45, 271.65, 
    271.35, 271.55, 272.25, 271.95, 272.35, 272.95, 272.65, 272.95, 273.35, 
    273.45, 273.75, 274.25, 274.35, 274.15, 274.35, 274.25, 274.15, 273.95, 
    274.05, 274.25, 274.15, 274.25, 273.65, 273.75, 274.25, 274.15, 274.65, 
    274.85, 274.95, 274.95, 275.15, 275.05, 275.15, 275.45, 275.55, 274.35, 
    274.95, 274.05, 273.55, 273.65, 273.35, 273.55, 272.75, 272.35, 271.75, 
    271.15, 271.85, 271.85, 272.15, 271.75, 271.75, 271.25, 271.35, 272.15, 
    273.15, 273.05, 273.05, 273.55, 273.35, 273.05, 272.55, 272.15, 272.35, 
    272.85, 273.25, 273.35, 273.25, 273.05, 272.75, 272.45, 272.15, 272.35, 
    272.05, 272.05, 271.95, 271.65, 271.55, 271.75, 272.05, 272.35, 272.25, 
    272.35, 272.45, 272.75, 272.65, 272.25, 272.55, 272.45, 272.45, 272.55, 
    272.75, 272.75, 272.75, 272.65, 272.55, 272.55, 272.65, 272.75, 272.95, 
    272.75, 272.75, 272.95, 272.95, 272.95, 273.05, 272.95, 272.95, 272.95, 
    273.05, 273.15, 272.95, 273.05, 272.85, 272.95, 273.05, 273.15, 273.25, 
    273.25, 273.25, 273.25, 272.85, 272.85, 272.15, 271.95, 272.45, 272.85, 
    273.25, 273.75, 273.65, 273.85, 274.15, 274.35, 273.95, 273.85, 273.75, 
    273.65, 273.45, 273.15, 272.95, 272.75, 272.75, 272.95, 272.95, 273.05, 
    273.15, 273.35, 273.55, 273.75, 273.75, 274.15, 274.15, 274.25, 274.95, 
    275.15, 274.95, 275.35, 275.45, 275.35, 275.45, 275.35, 275.05, 274.65, 
    273.85, 273.65, 272.15, 271.65, 271.45, 271.55, 271.55, 271.35, 271.25, 
    271.25, 271.15, 271.25, 270.95, 271.45, 271.25, 271.25, 271.45, 271.75, 
    271.85, 272.15, 271.75, 271.55, 271.25, 271.05, 270.55, 270.45, 269.65, 
    270.05, 270.05, 270.25, 271.05, 271.25, 271.85, 272.05, 272.15, 272.35, 
    272.55, 272.75, 272.95, 273.15, 273.15, 273.15, 273.15, 273.15, 273.35, 
    273.35, 273.35, 273.15, 273.15, 272.95, 273.15, 273.05, 273.05, 272.85, 
    272.65, 272.65, 272.55, 272.65, 272.65, 272.65, 272.75, 273.25, 273.15, 
    272.95, 272.65, 272.65, 272.45, 272.15, 271.65, 271.55, 271.25, 270.95, 
    271.05, 271.05, 270.95, 270.95, 271.45, 271.35, 271.55, 271.45, 271.35, 
    271.15, 271.25, 271.05, 270.95, 270.85, 271.05, 270.95, 271.15, 271.15, 
    271.35, 271.55, 271.65, 271.85, 271.85, 271.95, 271.95, 272.05, 272.05, 
    272.15, 271.75, 271.55, 271.75, 271.95, 272.05, 272.05, 272.25, 272.35, 
    272.45, 272.65, 272.75, 272.95, 273.05, 272.95, 272.75, 272.45, 272.45, 
    272.55, 272.55, 272.75, 272.85, 272.45, 272.05, 271.95, 272.05, 272.25, 
    272.35, 272.45, 272.25, 271.85, 271.55, 271.75, 271.65, 271.45, 271.05, 
    271.05, 270.95, 270.95, 270.85, 271.05, 271.05, 270.95, 270.65, 270.55, 
    270.25, 270.25, 270.45, 270.55, 270.45, 270.55, 270.45, 269.75, 269.45, 
    269.35, 269.35, 269.35, 269.55, 269.45, 269.65, 270.05, 270.65, 271.25, 
    271.65, 271.85, 272.05, 272.35, 272.75, 272.55, 271.75, 271.55, 272.25, 
    272.75, 272.85, 273.05, 272.95, 273.15, 273.35, 273.35, 273.45, 273.65, 
    273.75, 273.65, 273.65, 273.45, 273.25, 273.25, 273.65, 273.55, 273.45, 
    273.65, 273.65, 273.35, 273.35, 273.05, 272.55, 271.95, 271.45, 271.95, 
    272.75, 272.95, 273.55, 273.95, 273.85, 273.35, 273.65, 273.75, 273.75, 
    273.95, 273.85, 273.65, 273.95, 274.15, 274.45, 274.45, 274.55, 275.05, 
    274.65, 274.75, 274.85, 274.85, 274.65, 274.35, 273.85, 274.15, 274.05, 
    274.15, 274.25, 273.95, 274.15, 274.15, 274.05, 274.55, 274.55, 274.05, 
    273.85, 274.15, 273.95, 273.45, 273.75, 273.75, 273.65, 273.65, 273.65, 
    273.45, 273.45, 273.35, 273.05, 272.95, 272.65, 272.55, 272.55, 272.45, 
    272.45, 272.35, 272.35, 272.45, 272.55, 272.65, 272.75, 272.75, 272.35, 
    272.05, 271.45, 270.95, 271.05, 271.65, 271.45, 271.25, 271.05, 271.25, 
    271.55, 271.55, 271.45, 271.45, 271.55, 271.85, 271.95, 272.45, 272.95, 
    273.35, 273.35, 273.35, 273.55, 273.65, 273.35, 272.95, 273.25, 273.55, 
    273.65, 273.75, 274.05, 273.75, 273.25, 272.15, 271.25, 270.65, 270.55, 
    270.15, 269.95, 270.05, 270.05, 270.25, 270.35, 270.55, 270.85, 270.65, 
    270.25, 270.25, 270.55, 270.85, 271.05, 271.15, 271.35, 271.75, 271.65, 
    271.75, 272.05, 271.85, 272.35, 272.55, 272.75, 272.85, 273.15, 273.05, 
    273.15, 273.35, 273.55, 274.25, 274.35, 274.25, 274.05, 274.05, 274.05, 
    273.95, 273.85, 273.65, 273.25, 273.25, 273.35, 273.35, 273.35, 273.55, 
    273.75, 274.05, 274.25, 274.15, 274.25, 274.15, 274.45, 274.75, 275.95, 
    275.75, 275.85, 275.95, 274.35, 273.85, 273.95, 274.45, 274.35, 276.35, 
    274.65, 275.25, 275.85, 275.95, 275.95, 275.75, 276.05, 275.75, 277.25, 
    277.25, 276.65, 276.25, 276.25, 275.85, 276.15, 275.85, 276.65, 276.15, 
    275.75, 275.15, 275.15, 275.35, 275.65, 275.35, 275.05, 274.95, 275.05, 
    275.05, 275.05, 275.05, 274.75, 274.55, 274.55, 274.45, 274.05, 273.75, 
    273.05, 272.45, 272.05, 271.85, 271.75, 271.55, 271.45, 271.35, 271.25, 
    270.85, 270.75, 270.35, 270.35, 270.25, 270.05, 269.85, 269.65, 269.05, 
    268.75, 268.85, 268.15, 268.85, 269.05, 269.15, 268.95, 269.55, 269.65, 
    270.05, 270.85, 271.15, 271.05, 271.15, 271.35, 270.85, 270.95, 270.55, 
    270.25, 270.25, 270.65, 270.55, 271.05, 271.15, 271.25, 271.45, 271.55, 
    271.65, 271.75, 271.85, 271.85, 271.55, 271.55, 271.05, 271.35, 272.55, 
    274.25, 274.15, 273.25, 272.25, 271.45, 271.15, 271.15, 271.65, 272.25, 
    272.15, 272.95, 272.85, 273.15, 273.25, 273.65, 274.45, 273.65, 273.35, 
    272.85, 273.65, 273.45, 273.35, 273.25, 273.25, 272.35, 271.45, 270.75, 
    270.65, 271.05, 272.45, 272.35, 271.05, 270.75, 271.35, 271.85, 271.55, 
    271.65, 272.05, 270.75, 270.25, 269.85, 270.25, 270.15, 270.75, 270.85, 
    270.95, 271.25, 271.35, 271.55, 271.55, 271.65, 271.95, 272.05, 272.25, 
    272.45, 272.45, 272.65, 272.75, 272.95, 273.25, 273.25, 273.05, 273.05, 
    273.05, 273.15, 273.15, 273.35, 273.45, 273.55, 273.45, 273.45, 272.85, 
    272.65, 272.65, 271.65, 271.55, 270.95, 270.25, 269.95, 269.65, 270.45, 
    270.15, 270.95, 271.65, 273.25, 273.35, 273.45, 272.55, 272.15, 272.05, 
    271.85, 272.25, 272.65, 272.65, 272.55, 272.25, 272.05, 271.75, 271.85, 
    271.95, 271.95, 271.85, 271.85, 271.85, 272.05, 271.95, 271.75, 271.55, 
    272.35, 272.65, 272.95, 273.05, 273.05, 273.25, 273.35, 273.65, 274.15, 
    274.15, 274.05, 274.25, 274.35, 274.35, 274.05, 273.95, 274.05, 274.05, 
    274.05, 274.05, 274.05, 274.05, 273.95, 273.85, 274.05, 273.85, 274.15, 
    274.05, 274.25, 274.35, 274.45, 274.55, 274.45, 274.45, 274.25, 274.45, 
    274.45, 273.85, 273.55, 273.25, 273.15, 273.45, 272.55, 272.35, 272.25, 
    272.15, 271.95, 271.65, 271.35, 271.15, 270.85, 271.95, 271.65, 271.15, 
    271.15, 271.25, 271.35, 271.45, 271.65, 271.35, 271.15, 271.55, 271.65, 
    271.75, 272.35, 272.75, 272.55, 272.35, 272.35, 272.45, 272.45, 272.55, 
    272.75, 272.75, 272.95, 272.65, 272.95, 273.05, 273.15, 272.85, 272.95, 
    273.35, 273.95, 273.65, 273.65, 273.75, 273.75, 273.45, 272.55, 272.65, 
    272.55, 272.45, 272.25, 272.05, 271.95, 271.75, 271.65, 271.55, 271.35, 
    271.15, 270.65, 270.45, 270.05, 269.75, 269.65, 269.75, 269.55, 269.65, 
    269.25, 269.05, 269.25, 269.15, 268.85, 268.55, 268.25, 268.15, 267.75, 
    267.45, 267.15, 266.85, 266.65, 266.45, 266.45, 266.45, 266.55, 266.55, 
    266.55, 266.65, 266.65, 267.15, 267.55, 267.85, 267.65, 267.95, 268.25, 
    268.55, 268.85, 269.25, 269.85, 270.35, 270.95, 271.55, 271.95, 271.95, 
    271.85, 272.05, 272.35, 272.75, 272.65, 272.85, 273.25, 272.35, 272.15, 
    272.25, 273.05, 273.85, 274.15, 273.95, 274.05, 273.65, 273.45, 273.35, 
    273.65, 274.25, 274.45, 274.05, 274.35, 274.75, 274.65, 274.05, 274.25, 
    274.25, 274.55, 274.75, 274.45, 274.05, 274.05, 273.45, 273.55, 273.75, 
    273.75, 275.55, 274.25, 274.65, 275.15, 275.05, 275.35, 276.35, 275.85, 
    275.95, 275.45, 275.55, 275.45, 275.45, 275.45, 275.45, 275.25, 275.25, 
    275.35, 275.35, 275.05, 274.15, 273.75, 273.55, 273.35, 272.25, 271.95, 
    271.95, 271.85, 271.75, 271.45, 271.25, 271.25, 271.15, 271.05, 271.15, 
    270.95, 270.95, 271.15, 271.35, 271.75, 271.75, 271.65, 271.35, 271.25, 
    270.75, 270.75, 271.15, 270.85, 270.35, 269.85, 269.35, 269.25, 268.75, 
    269.15, 268.85, 268.55, 268.45, 268.25, 268.15, 267.95, 267.85, 267.75, 
    267.85, 267.75, 267.65, 268.15, 268.15, 268.25, 268.25, 268.25, 268.35, 
    268.45, 268.55, 268.65, 268.75, 268.85, 268.85, 268.35, 268.35, 268.15, 
    267.75, 267.85, 268.05, 268.05, 268.05, 267.95, 267.85, 267.85, 267.95, 
    267.85, 267.25, 266.95, 266.75, 266.75, 266.75, 266.75, 266.65, 266.45, 
    266.15, 265.95, 265.75, 266.45, 266.25, 266.05, 265.95, 265.85, 265.55, 
    265.45, 265.45, 265.45, 265.55, 265.75, 266.05, 269.45, 269.95, 270.75, 
    271.25, 271.65, 271.75, 271.85, 271.95, 271.95, 271.95, 271.95, 272.15, 
    271.55, 271.45, 271.35, 271.35, 271.25, 271.25, 271.25, 271.35, 271.55, 
    271.75, 271.85, 271.85, 271.45, 271.25, 270.75, 269.75, 269.25, 268.85, 
    268.45, 268.85, 268.95, 268.85, 269.25, 269.35, 269.35, 269.25, 269.65, 
    269.55, 269.35, 268.75, 268.55, 268.05, 266.85, 266.65, 266.15, 265.65, 
    265.55, 266.05, 266.35, 266.25, 266.55, 266.95, 266.65, 266.45, 266.85, 
    267.15, 268.25, 269.45, 269.25, 270.25, 269.65, 270.15, 270.45, 270.95, 
    271.15, 271.75, 272.15, 272.05, 272.05, 272.05, 271.85, 271.65, 271.45, 
    272.25, 271.95, 272.15, 272.05, 271.35, 271.85, 272.25, 272.25, 272.15, 
    271.95, 272.05, 272.05, 272.35, 271.25, 271.85, 271.75, 272.05, 272.05, 
    272.95, 272.85, 273.05, 272.95, 273.35, 273.35, 273.15, 273.65, 273.95, 
    273.85, 273.65, 273.55, 273.45, 273.15, 273.25, 273.15, 273.25, 272.45, 
    272.25, 272.45, 272.95, 271.95, 273.25, 273.65, 273.75, 274.45, 274.55, 
    273.85, 273.75, 273.65, 273.55, 273.45, 273.75, 273.65, 273.75, 273.85, 
    273.65, 273.65, 273.55, 273.35, 273.25, 273.25, 273.45, 273.75, 273.95, 
    273.85, 273.75, 273.75, 273.85, 273.45, 273.65, 273.45, 273.55, 273.35, 
    273.15, 273.35, 273.15, 273.05, 273.05, 272.95, 272.85, 272.45, 272.35, 
    272.45, 272.15, 273.25, 274.15, 274.15, 273.95, 273.75, 273.85, 273.65, 
    273.45, 273.35, 273.35, 273.35, 273.15, 273.15, 273.15, 273.45, 273.85, 
    274.05, 274.35, 274.25, 274.05, 273.85, 274.05, 273.85, 273.95, 273.95, 
    273.85, 274.15, 274.35, 273.95, 274.05, 273.65, 274.05, 274.05, 273.75, 
    274.15, 273.85, 273.65, 273.95, 273.75, 273.45, 273.45, 273.45, 273.35, 
    273.55, 273.15, 272.75, 273.25, 272.35, 272.15, 272.05, 271.85, 272.55, 
    272.65, 272.95, 272.85, 273.05, 272.95, 272.65, 272.65, 272.65, 272.85, 
    272.95, 272.85, 272.65, 272.45, 272.75, 272.65, 272.75, 272.85, 272.05, 
    271.55, 271.65, 272.85, 272.55, 272.25, 272.25, 272.25, 272.95, 273.05, 
    273.25, 273.15, 272.95, 272.65, 272.65, 272.35, 272.35, 272.25, 272.75, 
    272.55, 272.55, 272.05, 271.35, 271.85, 272.05, 272.25, 272.65, 272.55, 
    272.65, 272.25, 272.55, 272.85, 272.65, 272.45, 272.25, 272.35, 272.15, 
    272.25, 272.55, 273.15, 273.45, 273.45, 273.35, 273.25, 273.25, 273.35, 
    273.35, 273.65, 273.85, 273.85, 273.95, 274.05, 274.05, 274.15, 274.25, 
    274.05, 274.25, 274.65, 274.75, 274.75, 274.65, 274.55, 274.25, 274.35, 
    274.15, 274.05, 273.95, 273.85, 273.75, 273.75, 273.55, 273.55, 273.55, 
    273.55, 273.45, 273.05, 272.95, 272.65, 272.65, 272.75, 272.85, 273.15, 
    273.15, 273.25, 273.15, 273.25, 273.35, 273.55, 273.75, 273.55, 273.55, 
    273.55, 273.55, 273.45, 273.45, 273.45, 273.25, 273.05, 272.45, 272.75, 
    272.85, 272.65, 272.55, 272.45, 272.45, 272.25, 272.15, 272.45, 272.15, 
    272.25, 272.35, 272.35, 272.05, 271.85, 272.05, 272.05, 271.75, 272.25, 
    272.05, 272.05, 271.75, 271.95, 272.15, 272.35, 272.45, 272.55, 272.55, 
    272.85, 272.75, 272.65, 272.85, 272.95, 272.95, 272.85, 272.75, 272.75, 
    272.75, 272.55, 272.35, 272.75, 272.45, 271.85, 272.05, 271.75, 271.65, 
    270.75, 269.85, 268.75, 267.95, 267.15, 266.55, 265.95, 265.75, 265.55, 
    265.05, 265.65, 265.75, 266.05, 266.15, 266.05, 266.35, 266.45, 266.45, 
    266.35, 266.45, 266.75, 267.05, 267.65, 267.75, 267.75, 267.45, 267.55, 
    267.35, 267.55, 267.65, 266.85, 266.25, 264.95, 263.95, 263.95, 262.15, 
    264.05, 263.75, 264.75, 264.25, 264.95, 265.35, 265.45, 265.85, 264.95, 
    264.85, 265.35, 265.15, 266.55, 265.95, 266.85, 266.65, 267.05, 266.05, 
    267.55, 267.05, 266.25, 266.45, 267.85, 268.15, 268.45, 268.25, 267.95, 
    268.15, 268.85, 268.45, 268.55, 268.25, 267.55, 267.35, 267.65, 267.35, 
    267.35, 267.25, 267.25, 267.15, 267.05, 267.15, 266.85, 266.85, 266.85, 
    266.85, 266.75, 267.15, 267.05, 267.05, 267.25, 267.35, 267.35, 267.55, 
    267.45, 267.75, 267.75, 267.85, 267.85, 267.95, 268.05, 267.95, 268.35, 
    268.05, 268.45, 268.45, 268.65, 268.75, 268.85, 269.05, 269.05, 269.65, 
    270.05, 270.05, 270.25, 270.85, 271.65, 272.55, 271.65, 272.55, 272.45, 
    272.45, 272.45, 272.75, 272.35, 272.35, 272.15, 272.45, 272.45, 272.75, 
    272.75, 272.75, 272.85, 272.85, 272.95, 272.85, 272.95, 273.15, 273.45, 
    273.45, 273.75, 273.65, 273.95, 274.15, 274.05, 273.85, 273.35, 273.05, 
    272.25, 271.75, 271.25, 270.85, 270.15, 269.65, 269.25, 268.65, 268.45, 
    268.35, 268.25, 267.85, 267.45, 267.05, 266.85, 266.55, 266.05, 266.05, 
    265.85, 265.55, 265.65, 265.65, 265.55, 265.45, 265.45, 265.35, 265.25, 
    265.25, 265.15, 265.05, 264.85, 264.75, 264.95, 264.95, 264.65, 265.25, 
    265.15, 264.55, 263.55, 263.65, 264.05, 263.85, 263.65, 263.25, 262.95, 
    264.25, 263.95, 264.65, 265.75, 265.55, 265.55, 265.15, 264.95, 264.95, 
    264.45, 264.05, 263.75, 263.85, 263.55, 262.85, 263.05, 262.55, 262.55, 
    262.85, 262.95, 262.95, 262.45, 262.75, 263.05, 262.85, 262.75, 262.95, 
    263.05, 263.15, 262.95, 263.15, 263.05, 263.05, 263.05, 262.75, 262.65, 
    262.95, 262.85, 263.15, 263.15, 263.45, 263.75, 263.55, 263.75, 263.85, 
    263.75, 263.75, 264.05, 263.95, 263.95, 264.05, 263.95, 264.15, 264.05, 
    264.05, 264.15, 263.55, 263.25, 263.45, 263.55, 263.35, 263.35, 263.85, 
    264.95, 265.45, 265.65, 266.05, 266.45, 266.65, 266.95, 267.35, 267.55, 
    267.55, 267.65, 267.75, 268.05, 268.35, 268.75, 269.15, 269.55, 269.85, 
    269.95, 269.95, 270.05, 270.25, 270.45, 270.65, 270.75, 270.85, 271.25, 
    271.65, 271.85, 272.05, 272.05, 272.05, 272.15, 271.85, 271.85, 271.95, 
    272.65, 272.95, 272.85, 272.95, 273.05, 273.05, 272.55, 271.65, 271.35, 
    270.95, 271.55, 272.95, 273.05, 273.65, 273.45, 273.65, 273.55, 273.35, 
    273.35, 273.15, 273.05, 273.15, 273.15, 273.05, 273.05, 273.05, 273.05, 
    272.95, 272.95, 272.65, 272.95, 273.15, 272.85, 272.25, 272.35, 272.65, 
    272.65, 272.65, 273.25, 273.35, 273.35, 273.65, 273.65, 273.65, 273.65, 
    273.15, 273.15, 272.65, 272.45, 272.35, 272.05, 272.05, 271.45, 270.65, 
    269.25, 268.55, 268.35, 268.25, 267.95, 267.35, 267.15, 267.05, 266.85, 
    266.95, 266.95, 266.85, 266.95, 266.85, 266.85, 266.85, 266.95, 266.85, 
    266.85, 266.65, 266.65, 266.55, 266.55, 266.55, 266.65, 266.65, 266.55, 
    266.55, 266.35, 266.35, 266.15, 265.95, 265.65, 265.25, 264.95, 264.75, 
    264.45, 264.15, 263.95, 263.75, 263.75, 263.45, 262.85, 262.25, 262.35, 
    261.95, 261.35, 261.35, 260.75, 260.45, 260.45, 260.45, 259.85, 260.05, 
    259.65, 259.75, 259.55, 259.35, 259.35, 259.65, 259.85, 259.85, 259.35, 
    259.05, 260.35, 263.25, 262.45, 262.85, 262.15, 261.95, 262.25, 263.25, 
    263.25, 263.85, 263.85, 263.75, 263.75, 263.55, 263.35, 262.75, 263.05, 
    263.95, 264.45, 265.65, 265.95, 266.25, 266.45, 266.45, 266.55, 265.75, 
    264.95, 265.35, 263.95, 264.95, 266.55, 266.75, 267.15, 267.25, 267.35, 
    267.55, 267.55, 267.45, 267.25, 267.55, 267.55, 267.65, 267.25, 267.65, 
    268.05, 268.35, 269.05, 269.05, 269.15, 269.95, 270.65, 271.55, 271.95, 
    271.75, 271.45, 271.25, 271.05, 270.95, 270.85, 271.25, 271.45, 271.75, 
    271.75, 271.75, 271.25, 271.25, 272.15, 272.25, 272.25, 272.65, 272.95, 
    273.15, 273.15, 273.15, 273.15, 273.25, 273.35, 273.35, 273.25, 273.25, 
    273.05, 272.95, 272.95, 272.95, 272.85, 272.55, 272.45, 272.65, 272.65, 
    272.95, 273.05, 272.95, 272.55, 272.35, 272.35, 272.05, 272.05, 271.95, 
    272.25, 272.55, 272.75, 272.95, 272.75, 273.05, 273.15, 272.85, 272.95, 
    272.85, 272.95, 273.05, 273.15, 273.05, 272.95, 272.95, 272.95, 272.95, 
    273.05, 272.95, 272.95, 273.05, 273.15, 272.95, 272.95, 272.85, 272.95, 
    272.85, 273.05, 272.85, 273.05, 273.05, 272.95, 272.95, 272.95, 272.85, 
    272.85, 272.65, 272.75, 272.85, 273.15, 273.25, 273.15, 273.25, 273.25, 
    273.05, 272.85, 272.85, 272.95, 273.05, 273.15, 273.05, 272.95, 272.95, 
    273.05, 272.95, 272.95, 272.85, 272.85, 272.85, 272.75, 272.75, 272.65, 
    272.65, 272.75, 272.75, 272.65, 272.75, 272.55, 272.45, 272.15, 272.05, 
    271.45, 271.55, 271.75, 272.05, 272.25, 272.15, 271.75, 271.65, 271.65, 
    271.85, 271.95, 272.25, 271.95, 270.25, 269.95, 270.15, 270.65, 271.75, 
    271.25, 270.65, 271.65, 271.35, 271.25, 270.85, 270.95, 270.95, 270.55, 
    270.75, 270.65, 270.25, 270.25, 270.05, 269.95, 270.35, 270.45, 270.35, 
    270.55, 270.65, 270.75, 270.15, 270.15, 270.05, 270.25, 269.05, 270.15, 
    269.75, 269.95, 270.05, 270.05, 269.85, 269.95, 270.15, 269.65, 270.05, 
    270.05, 270.35, 270.25, 270.65, 270.85, 271.15, 271.35, 271.45, 271.55, 
    271.55, 271.75, 271.95, 272.15, 272.45, 272.65, 272.85, 272.95, 273.05, 
    273.35, 273.35, 273.25, 273.15, 273.05, 272.65, 272.55, 272.85, 273.15, 
    273.45, 273.15, 273.35, 272.75, 272.85, 272.75, 272.25, 271.85, 271.45, 
    271.35, 271.65, 271.95, 272.15, 272.35, 272.65, 272.65, 272.85, 272.55, 
    272.45, 272.45, 272.55, 272.55, 272.75, 272.45, 272.25, 272.25, 272.05, 
    271.95, 271.95, 271.75, 271.65, 271.25, 271.25, 271.55, 271.55, 271.55, 
    271.55, 271.25, 270.95, 271.45, 271.75, 271.85, 271.95, 271.85, 271.65, 
    270.75, 270.85, 270.25, 271.45, 269.35, 268.75, 267.85, 267.15, 266.75, 
    266.45, 266.15, 265.75, 265.95, 265.85, 265.85, 265.45, 265.35, 265.05, 
    264.95, 265.05, 265.05, 265.35, 265.25, 265.15, 265.25, 265.05, 265.35, 
    265.05, 265.35, 265.15, 265.25, 265.45, 265.85, 265.75, 265.95, 265.85, 
    265.85, 265.75, 265.65, 265.75, 265.75, 265.75, 266.35, 266.75, 267.45, 
    268.05, 268.45, 269.25, 270.05, 270.55, 270.55, 270.25, 270.25, 270.45, 
    269.95, 269.55, 269.55, 270.15, 270.05, 270.05, 269.15, 269.05, 268.55, 
    268.25, 267.95, 268.15, 268.05, 267.85, 267.85, 267.65, 267.35, 267.55, 
    267.45, 267.35, 267.15, 267.25, 267.15, 267.35, 267.25, 267.55, 267.65, 
    267.75, 268.05, 267.95, 268.15, 267.85, 268.05, 267.95, 267.85, 267.55, 
    267.25, 267.35, 267.45, 267.35, 267.25, 266.85, 266.65, 266.75, 266.65, 
    266.45, 266.35, 267.05, 267.85, 268.45, 268.95, 269.95, 269.35, 269.25, 
    268.55, 268.95, 269.35, 269.55, 269.75, 270.25, 269.95, 270.65, 267.95, 
    266.85, 265.85, 265.45, 265.75, 265.45, 265.85, 265.65, 265.05, 264.65, 
    265.05, 264.95, 264.55, 264.45, 263.85, 262.65, 261.55, 261.65, 262.55, 
    262.95, 265.35, 264.95, 264.45, 263.75, 266.05, 265.65, 265.85, 264.55, 
    263.95, 265.35, 267.95, 267.65, 267.65, 267.25, 267.25, 267.45, 267.05, 
    266.95, 267.25, 268.15, 268.75, 268.85, 268.95, 268.85, 267.75, 265.95, 
    266.95, 267.05, 267.35, 268.65, 268.55, 268.75, 269.15, 268.75, 269.55, 
    269.45, 269.65, 269.55, 269.15, 269.45, 269.15, 269.15, 268.75, 269.05, 
    269.05, 269.25, 269.25, 269.25, 269.05, 268.95, 269.15, 269.65, 269.55, 
    269.45, 269.55, 269.65, 269.65, 269.95, 269.95, 269.55, 268.95, 268.85, 
    268.85, 269.15, 269.05, 269.45, 268.85, 268.55, 268.35, 268.45, 268.15, 
    267.85, 267.95, 268.15, 268.05, 268.15, 268.25, 268.45, 268.65, 268.65, 
    268.45, 268.15, 268.25, 268.05, 268.15, 268.45, 268.55, 268.65, 268.55, 
    268.45, 268.05, 267.85, 267.85, 267.55, 266.95, 266.95, 267.05, 267.35, 
    267.05, 267.25, 266.65, 266.85, 265.95, 265.95, 265.65, 265.85, 265.25, 
    265.55, 265.15, 264.85, 265.15, 264.85, 264.85, 264.85, 264.95, 265.25, 
    265.15, 265.15, 264.95, 265.25, 264.05, 264.95, 264.35, 264.55, 264.55, 
    264.65, 265.05, 264.95, 264.65, 264.35, 264.15, 264.25, 264.25, 264.65, 
    265.35, 264.75, 265.45, 265.45, 265.35, 265.35, 265.45, 265.85, 265.95, 
    265.85, 265.55, 265.85, 266.25, 266.75, 266.95, 266.95, 267.35, 267.65, 
    267.85, 267.95, 268.25, 268.75, 269.05, 269.05, 268.85, 268.65, 268.45, 
    268.55, 268.55, 268.45, 268.65, 268.35, 268.35, 268.35, 268.45, 268.35, 
    268.85, 269.15, 269.15, 268.95, 268.85, 268.85, 268.75, 268.35, 268.15, 
    268.05, 268.05, 268.05, 268.15, 268.05, 268.15, 268.25, 268.45, 268.65, 
    268.65, 268.45, 268.95, 269.45, 269.95, 270.35, 270.65, 270.95, 271.05, 
    271.05, 271.35, 271.45, 271.55, 271.55, 271.55, 271.55, 271.45, 271.35, 
    271.35, 271.35, 271.45, 271.55, 271.55, 271.55, 271.55, 271.65, 271.45, 
    271.45, 271.25, 271.15, 271.15, 271.15, 271.25, 271.35, 271.25, 271.15, 
    271.05, 271.05, 271.05, 271.05, 271.15, 271.25, 271.35, 271.55, 271.75, 
    271.85, 271.85, 271.95, 272.25, 272.45, 272.45, 272.45, 272.35, 272.25, 
    272.25, 272.15, 272.15, 272.25, 272.15, 272.25, 272.05, 271.95, 271.95, 
    271.95, 271.95, 271.95, 271.95, 272.15, 272.35, 272.45, 272.55, 272.55, 
    272.45, 272.45, 272.25, 272.25, 272.25, 271.95, 271.95, 271.75, 271.65, 
    271.65, 271.85, 271.75, 271.65, 271.55, 271.55, 271.65, 271.95, 272.05, 
    272.15, 271.95, 272.05, 271.65, 271.35, 271.35, 271.05, 270.75, 270.45, 
    269.85, 269.75, 269.65, 269.25, 268.95, 268.55, 268.05, 267.85, 268.05, 
    267.85, 267.45, 267.55, 267.05, 266.75, 266.55, 266.75, 266.65, 266.95, 
    267.45, 267.45, 267.65, 267.75, 267.65, 267.65, 268.05, 269.85, 269.95, 
    269.55, 268.85, 268.35, 267.85, 267.55, 267.55, 267.75, 267.35, 266.75, 
    266.65, 266.45, 266.55, 266.85, 266.95, 266.95, 266.55, 266.55, 266.45, 
    266.15, 266.75, 267.15, 267.25, 267.05, 266.75, 266.35, 265.95, 265.45, 
    265.35, 265.15, 265.15, 264.95, 264.65, 264.35, 263.25, 264.25, 264.05, 
    263.75, 263.75, 264.05, 263.85, 263.85, 263.45, 263.45, 263.35, 263.35, 
    262.85, 262.95, 263.05, 262.45, 262.45, 262.35, 261.85, 261.85, 261.15, 
    260.35, 261.25, 261.15, 260.95, 260.75, 262.65, 259.85, 260.65, 259.35, 
    261.15, 260.25, 261.55, 260.75, 261.15, 261.65, 261.35, 261.25, 260.85, 
    261.05, 261.15, 261.15, 261.15, 261.05, 261.25, 260.95, 261.15, 261.15, 
    261.15, 261.05, 260.55, 259.85, 260.45, 260.55, 259.75, 261.15, 261.55, 
    261.55, 262.55, 262.85, 262.65, 263.25, 264.45, 264.95, 265.15, 265.05, 
    264.95, 265.15, 265.25, 265.45, 265.15, 264.95, 264.95, 262.75, 262.45, 
    262.15, 260.75, 261.05, 261.05, 260.75, 260.75, 260.65, 261.75, 261.45, 
    260.95, 260.55, 260.45, 259.95, 260.15, 259.85, 259.85, 259.85, 259.85, 
    259.95, 259.95, 259.75, 260.05, 259.85, 259.75, 259.65, 259.65, 259.85, 
    259.85, 260.05, 259.85, 260.05, 259.65, 259.85, 259.95, 259.65, 259.65, 
    259.15, 259.15, 259.15, 259.25, 259.45, 259.55, 259.65, 259.95, 259.75, 
    259.65, 260.05, 260.85, 261.55, 262.25, 261.55, 260.65, 259.45, 260.55, 
    262.35, 263.25, 262.65, 262.55, 262.15, 261.75, 262.75, 260.15, 258.85, 
    259.35, 259.95, 259.85, 260.55, 259.55, 259.35, 259.05, 259.65, 259.95, 
    259.75, 258.55, 260.35, 260.75, 258.35, 259.05, 260.65, 261.05, 260.45, 
    260.05, 259.95, 258.65, 260.55, 259.85, 259.05, 258.25, 258.15, 258.05, 
    259.05, 260.35, 261.15, 260.55, 259.95, 260.25, 261.25, 261.35, 261.05, 
    260.75, 260.45, 260.35, 260.05, 260.15, 260.15, 260.05, 259.45, 259.05, 
    258.75, 258.25, 258.65, 257.95, 257.95, 257.65, 257.75, 257.35, 257.05, 
    257.15, 256.55, 255.95, 255.75, 255.75, 255.75, 255.65, 255.75, 255.55, 
    255.45, 255.45, 255.25, 255.45, 255.35, 255.05, 254.95, 254.45, 254.25, 
    254.65, 254.95, 254.65, 255.45, 255.15, 253.75, 254.95, 254.65, 255.15, 
    255.25, 255.05, 253.85, 255.65, 255.55, 256.55, 256.65, 258.45, 258.45, 
    259.25, 259.25, 259.25, 258.25, 257.95, 257.45, 256.85, 257.05, 257.05, 
    256.35, 256.45, 256.35, 256.55, 256.75, 256.75, 256.85, 256.95, 257.05, 
    257.35, 257.85, 257.85, 257.75, 258.55, 258.15, 258.55, 258.95, 259.45, 
    260.25, 260.35, 260.75, 261.25, 261.45, 261.85, 262.05, 262.45, 263.05, 
    263.45, 263.85, 263.85, 264.25, 264.85, 265.15, 265.55, 266.15, 266.75, 
    267.15, 267.35, 267.45, 267.65, 267.85, 268.15, 268.65, 269.15, 269.15, 
    269.25, 269.25, 269.15, 269.15, 269.65, 270.65, 270.25, 269.95, 269.75, 
    269.65, 269.05, 268.95, 269.85, 270.75, 271.25, 271.45, 271.55, 271.55, 
    271.25, 271.75, 271.65, 271.65, 271.45, 271.45, 271.35, 271.35, 271.45, 
    271.45, 271.15, 270.95, 271.15, 271.05, 270.85, 270.95, 270.75, 270.55, 
    270.25, 269.65, 269.35, 268.95, 268.65, 268.35, 268.05, 268.15, 268.05, 
    268.05, 268.05, 267.85, 267.65, 267.45, 267.25, 267.15, 266.95, 266.85, 
    266.45, 265.75, 264.35, 264.15, 263.55, 263.05, 262.75, 262.65, 262.55, 
    262.75, 261.75, 261.65, 261.95, 261.65, 261.35, 261.05, 260.75, 260.45, 
    260.25, 259.95, 259.75, 259.45, 259.25, 259.05, 258.75, 258.65, 258.65, 
    258.75, 258.85, 259.05, 258.95, 259.25, 259.25, 259.05, 259.05, 258.95, 
    258.85, 258.65, 258.75, 259.25, 259.75, 260.25, 261.15, 261.85, 262.55, 
    263.45, 264.55, 266.05, 267.75, 269.25, 270.15, 270.55, 270.75, 270.75, 
    270.55, 270.55, 270.65, 270.65, 270.75, 270.65, 270.05, 268.95, 267.45, 
    265.75, 263.75, 261.25, 260.95, 260.15, 259.75, 259.45, 259.55, 259.75, 
    259.55, 259.25, 259.15, 260.35, 259.15, 259.25, 259.65, 259.65, 259.95, 
    260.15, 260.35, 260.55, 260.95, 261.25, 261.55, 261.65, 261.85, 261.75, 
    261.25, 260.65, 260.45, 259.75, 259.35, 259.25, 259.15, 259.15, 259.45, 
    259.75, 259.05, 258.35, 257.55, 257.15, 256.45, 256.05, 255.75, 255.05, 
    254.85, 254.55, 254.35, 254.45, 254.25, 254.25, 254.65, 255.05, 255.45, 
    255.95, 256.25, 256.45, 256.55, 256.65, 256.75, 256.85, 256.95, 257.45, 
    257.45, 257.15, 257.15, 257.25, 257.25, 257.15, 257.15, 257.25, 257.55, 
    257.95, 258.35, 258.65, 258.75, 258.55, 258.25, 258.05, 258.05, 257.75, 
    258.25, 258.75, 259.15, 259.45, 260.25, 261.15, 261.65, 262.15, 262.85, 
    263.55, 264.35, 264.15, 264.25, 264.55, 264.95, 265.25, 265.85, 265.55, 
    265.95, 267.25, 267.65, 268.15, 269.65, 269.45, 269.75, 269.95, 269.65, 
    269.35, 269.65, 270.15, 270.65, 270.75, 270.85, 272.05, 272.65, 273.05, 
    273.35, 273.45, 273.65, 273.05, 273.15, 273.25, 272.75, 272.85, 272.85, 
    272.85, 272.65, 272.55, 272.45, 272.15, 272.05, 272.35, 272.55, 272.75, 
    272.55, 272.45, 272.45, 272.55, 272.65, 272.75, 272.95, 273.05, 272.85, 
    272.45, 272.15, 272.05, 272.05, 271.95, 271.35, 271.25, 266.75, 272.05, 
    271.95, 272.55, 272.85, 272.65, 272.55, 273.05, 273.35, 273.55, 272.75, 
    272.95, 271.85, 272.25, 272.55, 272.75, 273.05, 273.25, 273.75, 273.15, 
    273.75, 273.75, 273.65, 272.85, 272.95, 273.45, 274.05, 274.15, 273.75, 
    273.55, 273.25, 272.45, 272.15, 272.65, 273.25, 273.35, 273.35, 273.05, 
    272.75, 273.05, 274.05, 273.25, 273.15, 273.05, 272.95, 272.85, 272.75, 
    272.95, 273.15, 273.15, 272.85, 272.85, 272.65, 272.25, 271.85, 271.35, 
    271.15, 271.45, 271.65, 271.75, 272.25, 273.05, 273.55, 271.35, 272.25, 
    271.95, 272.45, 271.75, 272.15, 272.95, 272.75, 272.45, 272.95, 272.75, 
    272.75, 272.75, 272.85, 273.15, 273.15, 273.05, 273.05, 273.05, 272.95, 
    272.85, 272.65, 272.45, 272.35, 272.25, 272.15, 272.05, 271.95, 271.75, 
    271.55, 271.25, 271.25, 271.35, 270.45, 270.35, 270.55, 270.65, 271.45, 
    270.65, 269.75, 269.45, 268.35, 267.55, 267.35, 267.25, 267.05, 266.85, 
    266.65, 266.45, 266.35, 265.15, 265.45, 265.85, 266.35, 266.05, 266.75, 
    267.45, 267.55, 268.35, 268.65, 268.45, 268.55, 268.55, 268.65, 268.75, 
    269.05, 268.85, 268.45, 268.25, 268.05, 267.95, 267.65, 267.45, 267.55, 
    267.65, 267.75, 266.25, 267.85, 268.15, 268.05, 267.55, 267.75, 267.05, 
    266.35, 265.85, 265.95, 265.85, 265.55, 265.35, 265.55, 265.65, 264.45, 
    263.45, 261.85, 262.25, 262.35, 262.15, 262.25, 261.65, 261.55, 260.95, 
    260.65, 261.15, 260.75, 260.75, 260.85, 260.95, 260.95, 261.35, 261.15, 
    261.25, 261.25, 261.25, 261.35, 261.35, 261.05, 260.65, 260.45, 258.55, 
    259.05, 258.65, 257.75, 257.15, 257.95, 257.35, 257.05, 256.75, 256.55, 
    256.85, 257.95, 259.25, 260.35, 259.85, 258.85, 258.65, 258.85, 259.15, 
    259.55, 259.95, 261.15, 262.05, 261.65, 261.05, 260.55, 260.05, 259.65, 
    259.55, 260.05, 259.85, 259.85, 260.35, 260.95, 260.45, 259.95, 260.65, 
    261.35, 261.15, 261.75, 262.25, 262.25, 262.05, 262.15, 262.55, 262.75, 
    263.05, 263.45, 263.55, 263.65, 263.95, 264.55, 264.45, 264.35, 264.85, 
    264.75, 264.65, 264.65, 264.75, 264.85, 264.95, 265.35, 264.85, 264.95, 
    264.85, 264.75, 265.15, 265.05, 265.15, 265.05, 264.85, 264.75, 264.75, 
    264.85, 264.95, 264.65, 265.45, 264.65, 265.15, 264.05, 262.75, 262.65, 
    262.45, 262.85, 262.65, 262.65, 262.95, 262.65, 262.55, 262.35, 263.15, 
    263.05, 263.45, 263.45, 263.65, 263.85, 264.25, 264.45, 264.05, 264.05, 
    263.45, 263.95, 264.95, 265.05, 264.95, 264.55, 262.25, 262.25, 261.65, 
    261.05, 260.65, 261.95, 263.85, 266.25, 266.05, 265.95, 266.05, 265.75, 
    265.55, 265.55, 265.25, 264.95, 265.05, 264.55, 264.15, 264.05, 263.35, 
    262.95, 262.55, 262.35, 262.35, 262.35, 262.45, 262.75, 263.15, 263.25, 
    263.95, 264.65, 264.95, 264.95, 265.35, 265.25, 264.55, 264.25, 264.05, 
    263.95, 263.95, 263.55, 263.95, 264.15, 265.05, 265.15, 264.75, 264.65, 
    264.05, 263.85, 263.05, 262.75, 262.55, 262.65, 262.95, 262.75, 262.95, 
    262.25, 262.85, 263.55, 264.05, 264.75, 264.45, 264.45, 264.05, 263.55, 
    263.35, 262.95, 263.35, 263.45, 262.05, 262.05, 261.35, 262.15, 264.35, 
    264.75, 264.15, 262.85, 262.55, 261.45, 261.25, 261.35, 261.75, 261.45, 
    261.95, 262.15, 263.35, 264.15, 264.95, 265.25, 266.15, 266.35, 267.15, 
    266.85, 266.85, 266.95, 266.85, 266.55, 266.55, 266.75, 266.65, 266.85, 
    267.75, 267.45, 267.45, 267.55, 267.75, 268.65, 269.05, 270.05, 270.05, 
    270.05, 269.95, 269.85, 269.85, 269.65, 269.35, 269.55, 269.75, 270.05, 
    270.25, 269.85, 269.65, 269.95, 270.35, 270.55, 270.55, 270.55, 270.35, 
    270.35, 270.15, 269.95, 269.45, 269.15, 269.35, 269.75, 269.55, 268.75, 
    267.95, 267.95, 268.55, 268.75, 267.75, 267.25, 267.25, 267.45, 267.45, 
    267.95, 268.25, 269.05, 269.55, 269.75, 269.55, 269.35, 268.85, 268.85, 
    268.65, 268.75, 268.15, 267.95, 267.75, 267.45, 268.05, 268.05, 268.05, 
    267.95, 267.85, 268.15, 267.55, 267.05, 267.55, 267.95, 267.45, 267.65, 
    267.35, 267.35, 267.15, 267.05, 266.35, 265.45, 265.35, 265.45, 265.75, 
    265.65, 265.85, 265.75, 266.25, 266.05, 265.85, 266.05, 266.45, 266.45, 
    266.35, 267.35, 267.35, 267.25, 266.35, 268.05, 268.55, 268.55, 266.85, 
    267.05, 267.05, 267.25, 267.95, 267.15, 266.55, 265.75, 266.05, 267.55, 
    268.05, 267.85, 267.95, 266.85, 267.15, 266.95, 266.35, 266.85, 267.05, 
    267.55, 267.35, 265.75, 264.35, 264.55, 264.45, 265.45, 262.95, 263.95, 
    263.85, 263.95, 264.95, 265.95, 266.15, 265.85, 266.35, 266.95, 267.45, 
    267.95, 268.65, 268.75, 268.75, 268.65, 268.35, 268.05, 266.15, 267.45, 
    266.65, 267.35, 267.35, 266.95, 266.85, 266.75, 266.45, 266.05, 265.95, 
    266.35, 265.85, 266.65, 267.25, 266.75, 267.45, 268.65, 269.05, 269.05, 
    268.45, 268.35, 266.95, 267.05, 267.15, 267.35, 267.65, 267.45, 267.95, 
    268.05, 267.85, 267.75, 267.85, 268.35, 268.25, 268.25, 268.35, 268.65, 
    269.45, 269.95, 270.85, 271.05, 270.85, 270.65, 271.25, 271.55, 271.65, 
    271.95, 272.25, 272.25, 272.25, 271.85, 271.85, 271.65, 271.55, 271.55, 
    271.55, 271.55, 271.35, 271.45, 271.55, 271.55, 271.55, 271.55, 271.55, 
    271.35, 271.35, 270.85, 271.15, 271.15, 270.85, 271.05, 270.75, 270.85, 
    270.45, 270.25, 270.15, 270.05, 269.85, 269.35, 269.05, 269.75, 269.25, 
    269.15, 268.75, 268.55, 268.95, 269.15, 268.95, 268.85, 268.95, 268.85, 
    268.75, 268.65, 268.35, 268.35, 268.25, 268.35, 268.45, 268.35, 268.05, 
    268.25, 268.15, 267.55, 267.65, 267.65, 267.65, 267.05, 267.25, 267.15, 
    266.95, 267.05, 266.85, 266.85, 266.85, 266.75, 266.55, 266.95, 266.45, 
    266.75, 266.65, 267.25, 266.75, 266.25, 266.15, 266.15, 266.25, 266.35, 
    266.35, 266.25, 265.55, 265.25, 264.95, 263.85, 263.05, 263.65, 263.45, 
    263.75, 263.55, 263.25, 263.25, 263.45, 263.35, 263.15, 263.45, 263.45, 
    263.55, 264.25, 264.65, 264.65, 264.35, 264.45, 264.25, 264.45, 264.85, 
    265.15, 265.55, 265.85, 266.05, 266.65, 267.05, 267.65, 268.75, 269.35, 
    269.35, 269.55, 269.85, 270.15, 270.35, 270.25, 270.25, 269.95, 269.55, 
    269.65, 269.65, 269.55, 269.25, 269.55, 269.85, 270.05, 270.15, 270.75, 
    270.55, 269.95, 269.45, 268.45, 268.45, 268.55, 268.05, 267.65, 267.75, 
    267.95, 267.95, 267.75, 267.75, 267.75, 267.55, 267.25, 266.95, 267.25, 
    267.35, 267.55, 267.65, 267.55, 267.75, 267.95, 268.05, 268.25, 268.95, 
    269.05, 268.65, 268.75, 268.35, 268.35, 268.85, 269.15, 268.85, 269.05, 
    269.05, 269.25, 269.15, 269.15, 269.35, 269.35, 269.15, 269.25, 268.95, 
    268.95, 268.75, 268.55, 268.55, 268.75, 269.15, 269.35, 269.25, 268.85, 
    268.45, 267.85, 267.45, 267.35, 266.95, 266.85, 266.45, 266.45, 265.45, 
    265.65, 266.55, 266.75, 266.85, 267.15, 267.35, 267.55, 267.45, 266.15, 
    265.15, 264.95, 264.75, 264.65, 264.65, 264.35, 264.15, 263.65, 263.95, 
    263.95, 263.45, 263.25, 263.45, 263.25, 263.35, 262.85, 262.25, 261.75, 
    261.45, 261.15, 260.25, 260.15, 260.15, 260.15, 260.45, 260.75, 261.05, 
    261.45, 262.05, 262.45, 262.95, 263.05, 263.55, 264.05, 264.15, 264.15, 
    263.85, 263.85, 263.65, 263.55, 263.55, 263.05, 263.25, 262.85, 262.05, 
    261.55, 261.25, 261.65, 263.05, 260.55, 262.45, 263.55, 264.15, 262.65, 
    264.65, 264.95, 264.75, 264.45, 264.55, 264.65, 264.55, 264.45, 264.45, 
    264.15, 263.25, 263.15, 263.45, 263.35, 263.55, 263.55, 264.05, 263.95, 
    263.65, 263.75, 264.05, 264.05, 264.25, 264.45, 264.05, 263.15, 263.25, 
    262.75, 261.75, 261.15, 260.85, 260.95, 260.95, 260.95, 261.05, 260.45, 
    260.05, 259.75, 260.55, 260.65, 260.85, 261.15, 261.55, 261.85, 261.25, 
    261.25, 260.95, 259.85, 259.85, 260.35, 260.55, 260.55, 261.05, 260.95, 
    260.95, 260.85, 260.75, 260.45, 261.05, 260.85, 260.25, 260.35, 260.65, 
    260.05, 259.85, 259.15, 258.95, 258.05, 258.55, 259.15, 259.45, 258.55, 
    258.65, 257.85, 258.65, 259.35, 259.05, 258.65, 258.35, 258.65, 258.75, 
    258.75, 258.65, 258.35, 258.65, 258.35, 258.55, 258.95, 258.65, 258.35, 
    258.75, 257.35, 258.25, 256.15, 256.25, 258.95, 259.45, 260.65, 261.05, 
    260.65, 259.75, 260.35, 260.65, 260.75, 261.05, 260.65, 260.75, 261.95, 
    263.15, 265.15, 266.15, 266.15, 266.25, 265.85, 266.15, 266.55, 266.95, 
    266.75, 266.85, 266.85, 266.95, 267.25, 267.35, 267.65, 267.85, 268.25, 
    268.45, 268.75, 269.15, 269.35, 269.85, 270.05, 269.85, 269.85, 269.95, 
    270.05, 270.05, 270.15, 270.25, 270.25, 270.25, 270.25, 270.15, 270.15, 
    270.25, 270.55, 269.95, 269.45, 269.55, 269.35, 269.05, 268.95, 268.55, 
    268.35, 267.65, 267.35, 266.85, 266.55, 266.25, 266.25, 266.45, 266.35, 
    266.45, 266.35, 266.35, 266.35, 266.05, 265.85, 265.15, 265.45, 265.45, 
    265.45, 265.25, 265.75, 265.95, 265.85, 265.75, 265.45, 265.05, 265.05, 
    264.65, 264.75, 264.95, 264.85, 264.75, 264.85, 264.65, 264.35, 263.95, 
    263.35, 263.15, 263.75, 264.05, 264.45, 264.55, 264.65, 264.75, 264.85, 
    264.85, 264.65, 264.85, 264.85, 264.65, 264.65, 264.65, 264.55, 264.85, 
    264.85, 264.75, 265.25, 265.35, 265.55, 264.85, 265.25, 265.15, 265.85, 
    266.55, 266.65, 266.65, 266.25, 265.95, 265.45, 265.35, 264.95, 264.75, 
    264.85, 264.85, 264.65, 264.65, 264.45, 264.05, 264.55, 261.45, 263.95, 
    264.45, 264.55, 264.75, 265.35, 265.75, 266.55, 266.55, 266.85, 267.05, 
    267.25, 267.85, 267.95, 267.25, 267.75, 268.05, 268.45, 268.55, 268.55, 
    267.75, 267.75, 267.15, 267.35, 267.65, 267.35, 267.55, 268.05, 268.25, 
    268.25, 268.45, 268.75, 268.85, 269.05, 269.15, 269.45, 269.75, 269.85, 
    269.95, 269.95, 270.15, 270.15, 270.15, 269.95, 269.85, 269.85, 269.85, 
    269.75, 269.75, 269.55, 269.65, 269.65, 269.65, 269.85, 269.85, 269.95, 
    270.05, 269.95, 269.65, 269.35, 269.45, 269.55, 269.65, 269.85, 269.75, 
    269.65, 269.75, 269.55, 269.55, 269.45, 269.35, 269.75, 269.25, 269.55, 
    269.65, 269.35, 268.85, 268.95, 268.65, 268.85, 268.75, 268.85, 269.25, 
    269.25, 268.75, 268.65, 268.55, 268.65, 269.15, 269.55, 269.95, 270.55, 
    270.25, 270.05, 269.95, 269.55, 269.35, 268.95, 268.85, 268.15, 268.15, 
    268.35, 268.55, 269.25, 269.55, 269.65, 270.15, 270.25, 270.25, 270.55, 
    271.05, 270.65, 270.55, 270.35, 270.45, 270.25, 269.45, 269.95, 270.05, 
    270.15, 270.95, 271.45, 271.75, 272.15, 271.35, 270.35, 270.35, 270.95, 
    271.05, 271.15, 271.45, 271.55, 271.65, 271.55, 271.55, 271.65, 271.55, 
    271.45, 271.05, 270.95, 271.05, 271.15, 271.05, 270.55, 270.95, 270.55, 
    270.45, 270.05, 270.75, 271.15, 271.55, 271.55, 271.25, 271.05, 270.85, 
    271.05, 271.45, 271.35, 271.35, 271.15, 270.85, 270.35, 269.95, 270.05, 
    269.85, 269.95, 270.35, 270.25, 269.35, 269.45, 269.45, 268.15, 268.75, 
    267.75, 267.75, 267.45, 267.65, 267.75, 267.75, 267.95, 268.95, 269.95, 
    270.05, 270.65, 271.05, 271.55, 271.45, 271.25, 271.15, 271.25, 271.25, 
    271.55, 271.55, 271.55, 271.65, 271.95, 272.05, 272.15, 272.05, 271.95, 
    272.05, 272.05, 272.05, 272.05, 272.05, 272.05, 272.15, 272.45, 272.35, 
    272.25, 272.15, 272.05, 271.95, 272.05, 272.15, 271.25, 270.65, 271.05, 
    270.95, 271.35, 271.35, 271.65, 271.55, 271.05, 270.75, 270.95, 271.35, 
    271.45, 271.35, 271.35, 271.45, 271.45, 271.55, 271.45, 271.35, 271.35, 
    271.25, 270.95, 270.85, 271.05, 271.55, 270.85, 271.05, 271.35, 270.85, 
    271.15, 270.65, 271.25, 270.65, 271.45, 271.55, 270.95, 270.75, 270.25, 
    270.45, 270.15, 269.95, 269.55, 269.05, 268.65, 268.25, 268.15, 268.25, 
    268.25, 268.75, 269.05, 269.15, 269.35, 269.15, 268.75, 268.95, 269.35, 
    269.25, 268.75, 268.05, 268.55, 268.45, 267.85, 266.85, 267.55, 267.85, 
    267.95, 265.05, 264.95, 265.45, 264.55, 264.35, 264.75, 263.85, 264.75, 
    265.85, 266.05, 265.65, 265.65, 266.15, 266.45, 265.75, 264.75, 265.05, 
    265.45, 265.45, 264.95, 264.45, 264.45, 264.45, 264.85, 264.55, 264.45, 
    265.95, 266.35, 265.65, 266.15, 265.85, 265.45, 265.55, 266.05, 266.05, 
    266.55, 265.75, 265.65, 265.95, 265.65, 265.85, 265.35, 265.55, 266.25, 
    266.25, 266.35, 265.55, 266.55, 266.85, 265.55, 264.65, 264.15, 264.25, 
    264.25, 265.25, 265.65, 266.15, 266.75, 265.85, 265.05, 265.45, 263.35, 
    262.95, 263.05, 262.75, 262.45, 260.95, 263.55, 262.55, 262.55, 263.75, 
    263.25, 263.25, 264.25, 264.15, 264.95, 263.75, 264.25, 263.65, 263.25, 
    262.75, 262.95, 261.75, 261.55, 261.05, 261.95, 263.35, 262.85, 262.65, 
    263.45, 263.95, 264.75, 264.65, 264.75, 264.15, 263.85, 263.75, 263.25, 
    264.05, 264.55, 264.95, 265.55, 266.05, 266.55, 266.45, 265.55, 266.45, 
    267.15, 265.95, 266.95, 266.85, 267.15, 267.45, 267.55, 267.45, 267.25, 
    267.35, 267.35, 268.05, 267.95, 268.25, 268.65, 269.15, 269.25, 269.65, 
    270.05, 270.45, 270.65, 270.55, 270.45, 270.35, 270.55, 270.95, 271.35, 
    271.65, 271.85, 272.15, 272.15, 272.05, 272.05, 272.05, 272.05, 272.15, 
    272.05, 272.05, 272.05, 272.05, 271.85, 271.85, 271.75, 271.75, 271.65, 
    271.55, 271.65, 271.55, 271.55, 271.55, 271.55, 271.65, 271.55, 271.55, 
    271.55, 271.55, 271.65, 271.65, 271.65, 271.65, 271.85, 271.95, 271.95, 
    271.75, 271.85, 271.95, 271.65, 271.65, 271.35, 271.45, 271.35, 271.15, 
    271.15, 271.25, 271.45, 271.35, 270.85, 270.65, 270.75, 271.35, 271.15, 
    271.05, 271.45, 271.45, 271.45, 271.35, 271.25, 271.45, 271.75, 271.65, 
    271.75, 271.65, 271.35, 271.05, 271.05, 271.05, 270.85, 270.65, 270.15, 
    269.65, 269.95, 268.85, 268.85, 268.35, 269.15, 269.45, 269.55, 269.15, 
    269.25, 269.45, 269.95, 270.65, 269.15, 269.15, 268.95, 270.15, 270.05, 
    269.65, 269.15, 269.75, 269.85, 269.65, 269.95, 270.25, 270.15, 269.65, 
    269.15, 268.65, 268.25, 267.75, 267.55, 267.25, 267.35, 268.65, 268.95, 
    268.95, 268.25, 267.65, 267.85, 267.95, 268.25, 268.15, 268.25, 268.55, 
    268.95, 268.65, 269.65, 269.45, 269.55, 268.85, 269.05, 269.15, 268.65, 
    266.45, 266.15, 266.25, 267.75, 268.05, 268.45, 268.55, 268.55, 268.95, 
    269.05, 269.15, 269.65, 270.25, 270.05, 270.25, 270.15, 270.35, 269.55, 
    269.95, 269.75, 269.65, 269.45, 269.35, 269.25, 268.75, 269.25, 269.25, 
    269.05, 268.75, 268.45, 268.35, 268.25, 268.45, 267.35, 267.55, 266.65, 
    267.55, 268.75, 269.25, 268.85, 268.85, 268.65, 268.55, 268.75, 269.15, 
    269.55, 270.25, 270.75, 270.85, 270.55, 270.45, 270.25, 269.95, 270.05, 
    270.15, 270.35, 270.45, 270.75, 271.05, 271.05, 271.05, 270.95, 270.55, 
    269.45, 269.75, 269.05, 268.85, 268.85, 269.65, 269.25, 267.65, 268.95, 
    268.55, 267.55, 267.75, 268.45, 268.65, 268.05, 268.35, 268.75, 268.45, 
    268.25, 267.35, 266.35, 266.75, 266.45, 266.25, 267.55, 268.55, 268.55, 
    268.85, 268.75, 268.85, 269.55, 269.85, 270.55, 270.85, 271.05, 271.45, 
    271.85, 271.95, 272.25, 272.15, 272.15, 272.25, 272.05, 271.95, 272.25, 
    272.35, 272.35, 272.25, 272.15, 271.15, 271.85, 271.25, 270.85, 270.75, 
    270.15, 269.85, 268.95, 268.85, 269.85, 270.65, 271.35, 271.35, 271.45, 
    271.55, 271.25, 271.45, 272.45, 272.45, 272.45, 272.45, 272.55, 272.35, 
    272.25, 271.55, 271.95, 272.45, 272.55, 272.75, 272.65, 272.35, 272.35, 
    272.75, 272.75, 272.65, 272.45, 271.65, 271.55, 270.85, 271.35, 271.35, 
    270.85, 269.95, 268.15, 268.05, 267.25, 266.55, 265.95, 265.45, 265.15, 
    264.75, 264.55, 264.45, 264.25, 264.25, 264.15, 263.65, 263.55, 263.55, 
    264.45, 265.15, 265.25, 265.75, 265.85, 266.05, 266.35, 266.55, 266.45, 
    266.05, 265.55, 264.75, 264.75, 263.75, 263.25, 262.85, 262.35, 262.35, 
    262.45, 262.25, 261.55, 261.65, 261.45, 261.15, 260.55, 260.55, 260.85, 
    260.65, 260.55, 260.55, 260.45, 260.95, 260.75, 260.55, 260.25, 259.45, 
    259.05, 259.05, 258.65, 258.85, 259.15, 259.25, 259.35, 259.75, 259.45, 
    259.35, 259.15, 259.05, 259.15, 259.55, 259.25, 259.65, 259.65, 259.45, 
    259.65, 259.95, 260.15, 259.85, 259.85, 259.55, 259.75, 260.05, 259.95, 
    259.95, 260.05, 259.85, 259.85, 259.65, 260.25, 260.35, 260.55, 261.25, 
    261.95, 261.65, 262.35, 262.25, 262.25, 261.95, 261.85, 261.65, 261.55, 
    261.75, 262.25, 261.75, 261.65, 261.95, 262.15, 261.75, 261.95, 262.25, 
    262.35, 262.45, 262.25, 263.05, 262.75, 262.45, 263.25, 262.95, 262.95, 
    262.95, 262.45, 262.65, 262.85, 262.35, 262.55, 261.95, 261.15, 260.85, 
    260.55, 260.75, 260.65, 260.45, 260.55, 260.75, 258.45, 257.95, 256.55, 
    256.35, 256.65, 257.25, 256.95, 257.25, 257.95, 254.95, 256.55, 257.35, 
    257.45, 257.95, 258.25, 258.05, 258.45, 259.45, 259.85, 260.35, 260.95, 
    260.75, 260.75, 260.85, 261.45, 262.05, 262.05, 262.15, 261.65, 261.45, 
    261.35, 261.35, 261.25, 261.15, 261.15, 261.15, 261.15, 260.85, 261.05, 
    260.75, 260.65, 260.55, 260.75, 260.75, 260.85, 260.95, 260.75, 260.55, 
    260.45, 260.15, 260.15, 260.15, 259.85, 260.05, 259.95, 259.85, 259.75, 
    259.75, 259.95, 260.15, 260.25, 260.25, 260.55, 260.85, 261.05, 261.15, 
    261.45, 261.55, 260.55, 260.95, 262.05, 260.55, 259.25, 259.25, 258.95, 
    259.45, 258.35, 256.95, 258.45, 258.25, 258.15, 258.15, 257.85, 258.75, 
    259.25, 259.85, 259.65, 260.45, 260.45, 260.95, 261.55, 261.55, 261.45, 
    261.95, 262.25, 262.45, 261.25, 260.75, 261.05, 260.55, 260.65, 260.05, 
    260.15, 258.45, 258.95, 259.35, 259.25, 258.85, 259.15, 258.35, 258.55, 
    258.25, 259.15, 258.55, 257.75, 259.55, 258.95, 259.45, 259.95, 260.25, 
    260.25, 259.05, 259.95, 259.65, 258.55, 258.55, 259.35, 258.05, 258.05, 
    258.25, 260.05, 260.75, 261.95, 263.05, 263.55, 263.95, 265.25, 267.65, 
    267.25, 267.35, 267.35, 267.75, 267.75, 267.95, 267.95, 268.35, 268.45, 
    268.25, 268.95, 269.15, 268.95, 268.75, 268.25, 268.25, 268.25, 268.15, 
    268.25, 268.25, 268.25, 268.15, 268.15, 267.85, 267.95, 267.95, 266.85, 
    267.75, 268.35, 268.15, 267.55, 267.85, 266.85, 266.45, 267.35, 267.25, 
    267.35, 267.35, 266.65, 267.05, 265.85, 266.35, 265.55, 266.05, 266.05, 
    265.05, 264.65, 264.75, 265.85, 265.95, 266.65, 267.25, 268.45, 268.25, 
    268.45, 268.45, 269.05, 269.15, 269.55, 269.45, 269.25, 269.45, 269.65, 
    269.85, 269.75, 269.75, 269.75, 269.85, 270.25, 270.65, 270.75, 270.95, 
    270.85, 270.85, 271.05, 271.05, 271.05, 271.25, 271.35, 271.45, 271.45, 
    271.35, 271.05, 270.95, 270.85, 270.85, 270.65, 270.45, 270.45, 270.45, 
    270.05, 269.75, 269.85, 269.95, 269.85, 270.05, 270.15, 270.15, 270.05, 
    270.05, 270.05, 270.25, 269.35, 269.05, 268.85, 267.55, 267.05, 268.15, 
    268.65, 268.05, 268.85, 268.35, 267.35, 267.35, 267.05, 267.15, 268.15, 
    267.75, 266.95, 266.95, 267.15, 267.85, 268.15, 267.45, 267.25, 267.25, 
    267.95, 267.15, 266.45, 266.55, 266.55, 265.95, 266.75, 266.45, 266.65, 
    266.25, 266.05, 265.65, 265.55, 265.65, 265.55, 265.45, 265.35, 265.25, 
    265.15, 264.85, 264.85, 264.55, 264.35, 263.95, 263.55, 263.05, 262.15, 
    261.95, 261.95, 262.15, 261.85, 261.85, 261.65, 261.25, 261.15, 260.75, 
    260.55, 260.55, 260.75, 260.75, 261.05, 261.65, 261.85, 262.05, 262.15, 
    262.05, 261.45, 260.85, 261.75, 263.45, 263.35, 263.45, 263.45, 263.25, 
    263.15, 263.15, 262.95, 261.25, 261.25, 261.95, 262.55, 262.35, 261.65, 
    262.05, 261.95, 261.25, 261.45, 262.85, 262.75, 263.15, 262.05, 262.65, 
    262.85, 263.25, 262.45, 262.45, 261.95, 261.75, 261.45, 262.55, 262.65, 
    262.25, 262.75, 263.75, 264.15, 263.95, 264.95, 265.25, 265.85, 266.15, 
    266.15, 266.75, 267.35, 267.55, 267.75, 267.95, 269.05, 269.25, 269.45, 
    269.35, 269.35, 268.95, 269.55, 269.35, 269.15, 269.25, 268.35, 268.75, 
    268.15, 268.35, 268.25, 267.95, 267.75, 267.95, 268.05, 267.65, 268.05, 
    267.75, 267.65, 267.35, 267.65, 268.25, 268.05, 267.55, 266.95, 266.95, 
    266.65, 265.95, 266.05, 266.25, 265.65, 265.65, 265.25, 265.15, 265.05, 
    265.25, 265.55, 265.65, 265.95, 266.55, 267.85, 268.05, 268.65, 268.65, 
    268.35, 268.25, 268.95, 268.35, 268.25, 268.15, 268.45, 268.55, 268.95, 
    268.75, 268.55, 268.25, 268.25, 268.15, 268.35, 267.85, 268.45, 267.95, 
    268.75, 269.35, 268.25, 267.95, 267.45, 268.15, 267.35, 266.65, 267.15, 
    267.45, 267.45, 267.95, 268.25, 268.55, 269.05, 269.55, 270.05, 269.55, 
    270.25, 270.25, 270.35, 270.45, 270.45, 270.35, 270.35, 270.15, 270.15, 
    270.05, 270.25, 270.25, 270.25, 269.65, 269.55, 269.45, 269.35, 268.75, 
    268.25, 267.25, 267.25, 267.95, 266.55, 266.45, 265.95, 265.85, 265.95, 
    265.75, 265.15, 265.75, 266.65, 266.25, 267.15, 267.15, 266.35, 266.65, 
    266.75, 267.25, 267.15, 267.55, 267.95, 267.65, 268.05, 268.05, 268.25, 
    267.75, 268.25, 268.45, 268.35, 268.25, 267.65, 268.35, 267.95, 268.05, 
    267.65, 267.65, 267.75, 267.95, 268.05, 267.85, 267.95, 267.75, 267.65, 
    267.65, 267.25, 267.15, 265.25, 264.35, 263.85, 262.85, 262.75, 261.65, 
    261.85, 260.65, 259.85, 259.55, 259.35, 259.15, 259.35, 259.85, 260.15, 
    260.25, 259.85, 259.35, 258.05, 256.95, 255.55, 255.45, 255.35, 254.45, 
    254.15, 254.15, 254.75, 255.05, 255.45, 255.85, 255.95, 256.35, 256.55, 
    256.85, 257.15, 257.95, 258.65, 259.25, 259.85, 260.45, 261.25, 261.55, 
    261.85, 262.65, 263.15, 264.05, 264.05, 263.55, 263.05, 262.85, 261.85, 
    261.25, 260.75, 260.45, 260.15, 259.95, 260.05, 259.35, 258.45, 258.25, 
    258.65, 258.55, 258.75, 258.75, 258.85, 258.85, 259.05, 258.95, 259.25, 
    259.35, 259.45, 259.55, 259.75, 260.05, 260.15, 260.15, 260.25, 260.45, 
    261.35, 260.55, 261.05, 261.35, 261.75, 262.15, 261.75, 260.95, 260.65, 
    260.85, 261.05, 261.15, 261.25, 261.35, 261.65, 261.15, 261.35, 261.25, 
    261.05, 260.45, 260.55, 260.25, 260.55, 260.25, 259.85, 259.35, 258.65, 
    258.75, 259.05, 258.75, 259.05, 259.65, 259.85, 259.85, 259.85, 259.55, 
    259.65, 259.75, 260.05, 259.75, 259.45, 259.55, 258.95, 259.35, 259.75, 
    259.45, 258.75, 259.15, 259.15, 259.65, 259.65, 260.05, 260.75, 260.95, 
    261.15, 262.05, 262.45, 263.05, 262.85, 263.05, 263.15, 262.75, 262.35, 
    260.95, 260.95, 262.25, 262.35, 262.35, 261.65, 261.75, 262.05, 262.15, 
    262.25, 262.35, 263.05, 262.95, 262.75, 262.65, 262.65, 262.85, 263.25, 
    263.45, 263.25, 262.85, 262.25, 261.85, 262.15, 261.15, 260.05, 260.15, 
    260.45, 259.75, 259.75, 259.65, 259.55, 259.35, 259.25, 258.95, 258.95, 
    259.65, 259.15, 259.35, 258.95, 259.45, 259.35, 260.55, 260.95, 261.65, 
    261.95, 261.65, 262.15, 261.55, 261.55, 262.55, 262.85, 262.65, 262.25, 
    261.15, 260.15, 259.75, 259.45, 259.65, 259.45, 258.65, 258.85, 259.45, 
    260.45, 260.95, 260.55, 261.15, 261.75, 262.15, 263.05, 264.05, 264.75, 
    265.95, 266.45, 268.75, 268.55, 267.65, 267.35, 267.55, 267.35, 267.75, 
    267.85, 268.25, 268.65, 269.15, 269.65, 270.15, 270.65, 270.85, 271.15, 
    271.15, 271.05, 271.05, 271.15, 270.65, 269.65, 269.65, 269.45, 269.15, 
    269.35, 269.25, 268.85, 268.55, 268.45, 268.55, 268.25, 268.25, 268.15, 
    268.05, 267.95, 268.05, 267.35, 265.85, 265.35, 264.95, 264.95, 264.55, 
    264.45, 264.05, 263.65, 263.55, 263.25, 263.05, 262.55, 262.65, 262.45, 
    262.05, 261.95, 261.85, 261.65, 261.65, 261.75, 261.95, 261.45, 261.55, 
    261.45, 261.35, 260.85, 260.65, 260.75, 260.45, 260.55, 260.65, 260.65, 
    260.75, 260.85, 260.85, 260.75, 260.85, 260.85, 261.05, 260.75, 261.15, 
    260.35, 262.05, 262.05, 261.95, 262.05, 262.15, 262.45, 262.35, 263.05, 
    263.35, 263.85, 264.35, 264.85, 265.25, 265.35, 265.65, 265.95, 266.25, 
    266.25, 266.35, 266.65, 266.75, 267.15, 266.85, 266.75, 266.95, 266.45, 
    266.35, 266.35, 266.65, 267.05, 267.45, 265.85, 267.15, 268.35, 268.15, 
    267.55, 265.85, 264.85, 264.75, 264.75, 264.15, 264.05, 264.45, 264.15, 
    263.95, 264.35, 264.45, 263.75, 264.05, 264.45, 264.55, 264.65, 264.55, 
    264.65, 264.45, 264.35, 264.25, 263.75, 263.85, 263.65, 264.05, 263.75, 
    263.15, 262.85, 262.75, 262.25, 261.85, 261.95, 261.65, 261.65, 261.15, 
    261.15, 261.15, 260.55, 260.15, 260.45, 260.55, 260.85, 260.95, 260.85, 
    260.65, 260.85, 260.85, 260.35, 259.25, 258.95, 258.45, 258.25, 258.05, 
    257.95, 260.15, 257.65, 257.65, 257.95, 256.85, 256.95, 257.45, 257.85, 
    259.25, 260.95, 262.35, 263.35, 264.45, 265.45, 265.35, 265.05, 265.65, 
    265.85, 265.95, 266.15, 266.15, 265.35, 263.85, 263.75, 263.55, 264.45, 
    264.65, 264.75, 264.35, 264.25, 264.85, 266.05, 266.45, 267.15, 267.35, 
    268.05, 268.45, 268.45, 267.65, 268.05, 268.45, 268.45, 266.95, 267.55, 
    266.85, 266.85, 266.85, 266.05, 265.45, 266.25, 265.85, 265.25, 265.15, 
    265.35, 265.45, 266.15, 265.85, 266.15, 266.95, 267.25, 269.05, 269.55, 
    268.05, 268.05, 268.25, 267.35, 267.25, 267.05, 266.65, 266.55, 267.15, 
    266.45, 265.95, 265.15, 264.05, 264.45, 264.05, 264.75, 264.65, 264.85, 
    264.95, 265.05, 265.05, 265.25, 265.25, 265.35, 265.55, 265.75, 265.95, 
    266.55, 267.15, 268.55, 267.75, 268.85, 268.95, 269.55, 270.05, 269.55, 
    269.55, 267.65, 266.85, 265.65, 266.05, 267.55, 267.75, 267.85, 268.45, 
    269.55, 270.45, 270.35, 271.25, 271.45, 272.55, 272.65, 271.45, 269.85, 
    268.55, 268.35, 268.45, 268.45, 268.25, 268.55, 269.05, 269.25, 269.45, 
    270.55, 270.75, 270.15, 271.55, 270.45, 270.65, 271.15, 271.75, 272.25, 
    272.75, 272.15, 270.75, 269.85, 268.45, 268.35, 267.95, 267.95, 268.05, 
    267.35, 267.75, 267.15, 266.25, 265.65, 265.05, 265.45, 265.25, 264.35, 
    264.05, 263.65, 263.65, 263.55, 263.35, 263.15, 262.95, 262.25, 262.45, 
    262.05, 262.25, 261.95, 261.45, 261.15, 261.35, 260.65, 260.35, 260.45, 
    259.45, 260.25, 259.65, 259.15, 259.45, 260.45, 260.55, 261.05, 261.25, 
    261.55, 262.15, 261.85, 261.85, 262.45, 262.15, 262.15, 261.85, 261.55, 
    261.15, 261.05, 261.05, 260.85, 261.15, 261.05, 260.85, 260.75, 260.75, 
    260.25, 258.95, 260.65, 260.45, 261.05, 260.65, 261.55, 262.35, 262.25, 
    262.75, 262.75, 263.25, 263.35, 263.65, 263.75, 263.25, 263.55, 264.15, 
    264.15, 264.05, 263.45, 263.05, 262.75, 262.65, 262.75, 264.05, 263.55, 
    263.85, 264.05, 264.35, 264.75, 264.55, 264.65, 264.95, 263.95, 264.05, 
    264.45, 264.55, 264.45, 264.65, 264.35, 264.25, 264.75, 265.15, 265.15, 
    265.55, 265.65, 265.55, 265.25, 265.45, 265.65, 266.75, 266.95, 267.05, 
    267.15, 267.15, 267.15, 267.15, 267.15, 267.25, 266.75, 266.85, 266.45, 
    266.25, 265.75, 265.55, 265.95, 266.05, 266.25, 266.15, 266.45, 266.85, 
    267.15, 267.05, 267.25, 267.85, 268.55, 269.35, 270.15, 269.65, 269.55, 
    269.25, 268.65, 268.25, 268.15, 267.75, 267.95, 268.95, 269.65, 269.85, 
    269.85, 270.25, 270.65, 271.05, 270.65, 270.95, 271.15, 271.35, 271.35, 
    271.25, 271.25, 271.25, 271.25, 271.05, 270.85, 270.65, 270.55, 270.35, 
    269.95, 270.05, 269.75, 269.45, 268.85, 268.75, 268.65, 268.85, 269.15, 
    269.15, 268.95, 269.05, 269.25, 269.35, 269.65, 269.85, 269.85, 269.85, 
    270.15, 270.25, 270.15, 270.15, 270.05, 269.45, 269.55, 269.55, 269.25, 
    269.05, 268.95, 268.75, 268.65, 268.55, 268.65, 268.45, 268.75, 268.85, 
    268.95, 268.75, 268.75, 268.65, 268.35, 268.75, 268.85, 269.25, 269.65, 
    269.85, 269.85, 269.85, 269.65, 269.65, 269.45, 269.55, 269.55, 269.55, 
    269.75, 269.85, 269.95, 270.15, 270.25, 270.35, 270.65, 270.65, 270.55, 
    270.25, 270.35, 270.25, 270.35, 270.45, 270.35, 270.35, 270.05, 269.85, 
    269.65, 269.35, 269.25, 269.15, 268.95, 269.05, 269.35, 269.35, 269.35, 
    269.45, 269.85, 270.15, 270.35, 270.85, 271.05, 271.05, 271.25, 271.65, 
    271.85, 272.05, 272.15, 272.25, 272.35, 272.35, 272.45, 272.35, 272.15, 
    271.95, 271.45, 271.25, 271.35, 271.45, 271.45, 271.45, 271.35, 271.35, 
    271.45, 271.65, 271.65, 271.55, 271.55, 271.25, 271.25, 271.35, 271.15, 
    271.15, 271.15, 271.25, 271.35, 271.25, 271.25, 271.15, 271.05, 270.95, 
    270.95, 270.95, 270.95, 270.95, 271.05, 271.05, 271.05, 270.95, 271.05, 
    271.05, 271.15, 271.25, 271.45, 271.35, 271.35, 271.35, 271.65, 271.65, 
    271.55, 271.75, 271.75, 271.65, 271.55, 271.55, 271.45, 271.55, 271.35, 
    271.25, 271.15, 271.25, 271.55, 271.75, 271.95, 272.05, 272.25, 272.25, 
    272.25, 272.55, 272.45, 272.75, 272.95, 272.95, 272.95, 273.25, 272.95, 
    273.15, 272.65, 271.95, 271.95, 271.55, 271.95, 271.85, 271.85, 271.95, 
    271.75, 271.85, 272.25, 272.55, 272.85, 272.55, 272.05, 271.95, 271.75, 
    271.15, 270.75, 271.35, 270.85, 270.75, 270.45, 270.85, 270.65, 270.75, 
    270.75, 270.75, 271.65, 271.35, 271.05, 270.65, 270.35, 269.65, 271.05, 
    269.85, 269.05, 269.85, 270.45, 272.95, 269.85, 269.65, 269.75, 269.55, 
    269.35, 268.95, 268.95, 268.85, 269.05, 268.95, 269.05, 268.95, 269.05, 
    269.05, 268.95, 268.95, 268.95, 268.95, 268.95, 269.15, 269.25, 269.05, 
    269.05, 269.05, 269.35, 269.25, 269.35, 269.15, 269.15, 269.05, 268.75, 
    268.55, 268.55, 268.35, 268.25, 268.15, 268.25, 268.35, 268.65, 268.55, 
    268.75, 268.85, 268.85, 269.25, 269.25, 269.15, 269.35, 269.45, 269.55, 
    269.65, 269.25, 269.35, 269.35, 268.95, 268.85, 268.75, 268.85, 268.85, 
    268.85, 268.25, 268.45, 268.15, 268.05, 268.75, 268.95, 269.15, 269.05, 
    269.75, 269.55, 269.25, 269.05, 269.15, 269.05, 269.45, 268.55, 268.45, 
    268.65, 268.55, 268.75, 269.15, 268.75, 269.35, 269.55, 269.65, 269.75, 
    269.45, 269.55, 269.65, 269.55, 269.45, 269.45, 269.05, 269.05, 268.85, 
    269.45, 270.15, 270.65, 271.15, 271.75, 272.15, 273.35, 272.05, 271.55, 
    271.45, 271.35, 271.25, 271.25, 270.75, 270.95, 270.75, 271.45, 270.65, 
    270.65, 271.35, 272.25, 271.25, 271.75, 272.45, 272.25, 272.25, 272.35, 
    272.35, 272.25, 272.35, 272.55, 272.75, 272.65, 272.35, 271.95, 271.35, 
    271.75, 271.75, 272.35, 271.95, 272.45, 273.25, 272.95, 273.05, 273.35, 
    273.55, 273.55, 273.65, 274.85, 274.35, 274.75, 274.25, 273.75, 272.75, 
    272.65, 272.65, 272.95, 272.45, 272.55, 272.35, 272.15, 272.15, 271.95, 
    272.05, 272.15, 272.25, 272.45, 272.35, 272.65, 272.85, 272.45, 272.35, 
    272.25, 272.35, 272.85, 273.15, 272.95, 272.25, 272.05, 272.05, 272.05, 
    272.05, 271.95, 271.95, 271.85, 271.85, 271.95, 271.65, 271.55, 271.25, 
    271.25, 272.15, 272.45, 272.75, 272.25, 272.25, 272.65, 272.15, 271.55, 
    271.85, 272.85, 272.15, 272.35, 272.05, 271.45, 271.25, 271.05, 270.75, 
    270.85, 271.05, 271.25, 271.15, 271.45, 271.25, 271.05, 270.65, 270.85, 
    271.45, 271.55, 271.35, 271.75, 272.05, 272.55, 272.65, 271.95, 271.55, 
    271.25, 270.95, 270.85, 270.65, 270.55, 270.55, 270.35, 270.35, 270.35, 
    270.35, 270.35, 270.15, 270.05, 270.15, 270.25, 270.45, 270.55, 270.75, 
    271.05, 271.25, 271.45, 271.35, 271.55, 271.55, 271.65, 271.95, 272.25, 
    272.85, 273.25, 273.35, 273.35, 273.15, 272.95, 272.65, 272.35, 272.25, 
    272.15, 272.15, 272.05, 272.85, 272.85, 273.05, 272.85, 272.75, 272.65, 
    272.35, 272.65, 272.55, 272.65, 272.65, 272.35, 272.05, 271.15, 271.75, 
    271.95, 271.85, 271.95, 271.95, 272.15, 272.15, 272.25, 272.45, 272.65, 
    272.15, 272.05, 272.15, 271.95, 272.25, 272.05, 272.25, 272.35, 272.45, 
    272.45, 272.45, 272.65, 272.75, 272.75, 272.95, 272.95, 273.15, 272.75, 
    272.45, 272.55, 272.35, 272.45, 272.45, 272.65, 272.45, 271.15, 270.95, 
    270.95, 271.15, 271.35, 271.75, 271.85, 271.75, 271.95, 272.05, 272.05, 
    272.15, 272.15, 272.15, 272.35, 272.65, 272.45, 272.45, 272.45, 272.25, 
    272.35, 272.15, 271.85, 272.25, 272.55, 272.65, 272.65, 272.75, 272.85, 
    272.75, 272.95, 272.85, 272.75, 272.85, 272.85, 272.65, 272.75, 272.65, 
    272.35, 273.15, 273.25, 274.25, 274.05, 273.05, 272.65, 272.15, 271.95, 
    272.15, 271.05, 271.25, 271.45, 271.35, 271.65, 271.35, 271.35, 271.55, 
    271.95, 271.75, 271.45, 271.15, 271.15, 271.05, 271.05, 270.85, 270.75, 
    270.35, 269.95, 269.95, 269.75, 270.15, 269.95, 270.05, 270.25, 270.45, 
    270.55, 270.25, 269.95, 269.75, 269.55, 269.65, 269.35, 269.15, 269.65, 
    269.85, 269.85, 270.25, 270.25, 270.25, 270.55, 270.25, 270.25, 270.45, 
    270.35, 270.55, 270.75, 270.75, 270.85, 271.05, 271.05, 270.95, 270.85, 
    270.85, 270.85, 270.65, 270.55, 270.65, 270.55, 270.25, 270.25, 270.35, 
    270.25, 270.15, 270.15, 269.75, 269.95, 269.95, 269.75, 269.45, 269.65, 
    269.65, 269.55, 269.65, 269.95, 269.95, 270.15, 270.25, 270.35, 270.65, 
    270.65, 270.75, 270.75, 270.65, 270.55, 270.45, 270.55, 270.55, 270.45, 
    270.55, 270.55, 270.45, 270.45, 270.45, 270.55, 270.55, 270.75, 270.65, 
    270.85, 270.95, 270.85, 270.75, 270.75, 270.75, 270.55, 269.65, 268.95, 
    268.95, 268.95, 269.35, 268.95, 269.65, 270.35, 270.35, 270.15, 270.05, 
    269.75, 269.55, 269.75, 269.95, 270.15, 270.25, 270.55, 270.85, 270.75, 
    270.55, 271.05, 270.65, 271.45, 271.55, 271.95, 271.95, 270.75, 271.75, 
    271.75, 271.75, 272.05, 272.15, 272.15, 272.25, 272.25, 272.15, 272.35, 
    272.35, 272.35, 272.05, 272.05, 272.65, 271.75, 271.65, 271.85, 271.95, 
    272.05, 271.65, 271.15, 271.05, 271.05, 271.75, 271.65, 271.65, 271.65, 
    271.65, 271.75, 271.55, 271.45, 271.35, 271.35, 271.25, 271.45, 271.65, 
    271.65, 271.75, 271.75, 272.15, 272.15, 272.15, 271.95, 271.55, 271.55, 
    271.45, 271.75, 271.85, 271.75, 271.85, 271.85, 271.95, 272.05, 272.15, 
    272.35, 272.15, 272.45, 272.45, 272.45, 272.65, 273.35, 272.55, 272.65, 
    272.75, 272.65, 273.05, 272.65, 272.65, 272.55, 272.45, 272.65, 272.45, 
    272.45, 272.35, 273.05, 272.45, 272.35, 272.35, 272.35, 272.55, 273.15, 
    273.05, 272.35, 272.25, 272.45, 272.65, 272.75, 272.85, 272.85, 272.95, 
    273.25, 272.65, 273.05, 272.85, 272.65, 273.55, 272.35, 272.05, 270.95, 
    271.85, 271.95, 271.35, 271.55, 270.35, 271.85, 271.85, 271.35, 271.05, 
    271.15, 271.65, 270.75, 270.55, 270.95, 271.05, 270.95, 271.15, 271.05, 
    271.25, 271.65, 271.25, 271.25, 270.95, 271.15, 271.25, 271.35, 271.65, 
    271.25, 271.25, 271.35, 271.65, 271.65, 271.85, 273.55, 273.05, 272.65, 
    272.65, 272.65, 272.75, 272.15, 272.75, 272.55, 272.45, 272.75, 272.55, 
    272.75, 272.55, 272.45, 272.95, 272.65, 272.55, 272.75, 272.65, 272.75, 
    272.85, 273.45, 273.15, 273.35, 273.25, 273.05, 273.15, 273.45, 273.65, 
    273.65, 273.25, 273.35, 272.95, 272.95, 273.25, 273.25, 273.35, 274.15, 
    273.35, 272.45, 273.05, 273.05, 272.95, 272.55, 272.75, 272.55, 272.45, 
    272.05, 271.95, 271.85, 271.25, 271.65, 271.65, 270.85, 271.25, 271.35, 
    271.35, 271.75, 271.35, 271.75, 272.65, 272.25, 272.65, 272.25, 272.75, 
    272.65, 273.45, 272.45, 272.55, 273.45, 274.75, 275.15, 274.45, 274.65, 
    274.35, 274.35, 274.45, 274.35, 274.05, 273.95, 273.95, 274.65, 273.75, 
    273.75, 273.15, 273.75, 273.75, 273.65, 273.95, 273.35, 273.75, 274.75, 
    274.55, 274.35, 274.25, 274.05, 274.65, 274.55, 274.15, 274.25, 274.05, 
    274.85, 274.85, 274.65, 275.05, 274.65, 274.85, 274.25, 274.25, 274.05, 
    273.35, 273.75, 273.75, 273.65, 273.95, 274.05, 274.55, 274.25, 274.15, 
    274.05, 273.35, 273.05, 273.45, 273.45, 273.35, 273.55, 273.85, 273.45, 
    272.75, 272.65, 272.65, 272.95, 273.05, 272.95, 272.95, 273.15, 273.15, 
    273.05, 273.15, 273.55, 273.95, 273.85, 273.65, 273.55, 273.95, 274.45, 
    274.45, 274.65, 273.75, 274.35, 274.65, 275.05, 275.15, 274.25, 273.55, 
    273.45, 273.35, 272.75, 272.85, 272.75, 272.75, 272.85, 272.85, 273.75, 
    272.85, 272.95, 273.05, 273.05, 274.05, 273.15, 273.05, 272.95, 273.05, 
    273.15, 273.05, 272.95, 272.85, 272.95, 273.35, 272.95, 273.05, 272.95, 
    272.95, 273.05, 273.15, 274.05, 273.35, 273.25, 273.55, 273.75, 273.65, 
    274.15, 274.35, 274.35, 274.45, 274.75, 275.25, 276.25, 276.25, 275.65, 
    276.25, 276.35, 275.75, 276.25, 275.55, 276.25, 275.65, 275.85, 275.45, 
    275.55, 277.15, 275.45, 275.55, 276.35, 276.95, 277.25, 275.65, 274.25, 
    274.15, 273.75, 275.25, 273.55, 273.65, 273.75, 273.85, 275.25, 273.65, 
    273.75, 273.45, 273.45, 274.95, 273.75, 273.95, 274.45, 274.65, 273.75, 
    274.65, 274.65, 274.65, 275.05, 275.25, 274.95, 274.85, 275.45, 275.35, 
    274.85, 275.05, 274.75, 274.85, 274.55, 274.15, 273.95, 273.55, 273.35, 
    273.15, 273.25, 273.55, 273.45, 273.15, 273.35, 273.55, 273.55, 273.45, 
    272.85, 273.15, 273.65, 273.75, 274.45, 274.65, 275.05, 275.35, 275.65, 
    275.05, 275.15, 274.75, 274.15, 273.85, 274.25, 274.05, 274.35, 274.75, 
    273.95, 274.05, 274.25, 274.55, 274.75, 275.25, 275.65, 275.95, 276.95, 
    276.25, 276.05, 276.25, 275.25, 275.45, 275.75, 275.55, 276.75, 275.95, 
    275.65, 275.45, 275.15, 274.45, 274.75, 274.65, 275.95, 275.15, 275.45, 
    275.15, 275.55, 275.55, 274.45, 274.55, 275.15, 275.55, 275.45, 275.65, 
    275.45, 274.65, 274.75, 274.75, 275.15, 274.65, 275.25, 275.65, 274.65, 
    275.15, 275.65, 276.05, 275.95, 275.65, 275.45, 275.25, 275.15, 274.55, 
    274.35, 274.25, 274.15, 273.95, 273.55, 273.65, 273.45, 273.35, 273.25, 
    273.35, 273.35, 273.55, 273.65, 273.65, 273.35, 274.05, 274.35, 274.55, 
    274.65, 274.65, 274.45, 274.55, 274.85, 275.35, 276.05, 276.25, 276.25, 
    276.25, 276.45, 275.75, 275.15, 275.35, 275.25, 276.25, 276.25, 275.85, 
    275.25, 274.95, 274.25, 274.35, 274.35, 274.15, 273.85, 273.85, 273.55, 
    273.35, 272.85, 272.75, 273.15, 273.55, 273.95, 273.95, 274.15, 274.15, 
    274.15, 274.65, 274.15, 273.95, 273.95, 274.25, 273.95, 274.15, 274.25, 
    274.75, 274.45, 274.75, 275.05, 275.05, 275.05, 274.95, 274.75, 274.65, 
    274.75, 274.95, 274.45, 274.45, 274.75, 274.95, 274.65, 274.55, 274.95, 
    274.65, 274.55, 274.25, 274.05, 273.85, 273.55, 273.55, 273.65, 273.65, 
    273.75, 273.85, 273.35, 274.05, 274.35, 274.55, 274.65, 274.35, 274.35, 
    274.45, 274.55, 274.35, 274.45, 274.35, 274.35, 274.35, 273.65, 273.45, 
    273.55, 273.65, 273.75, 273.95, 274.15, 274.05, 273.85, 274.75, 274.95, 
    274.55, 274.25, 275.05, 275.95, 276.15, 277.65, 274.45, 274.45, 274.65, 
    273.75, 273.75, 274.55, 274.25, 274.45, 274.45, 274.55, 274.05, 274.15, 
    274.45, 274.65, 275.45, 275.45, 275.45, 275.85, 275.65, 275.45, 275.15, 
    275.35, 275.45, 275.35, 275.65, 275.85, 275.65, 275.55, 275.65, 276.95, 
    276.65, 275.65, 273.85, 274.75, 275.35, 274.75, 274.55, 274.55, 274.75, 
    275.25, 275.35, 275.05, 275.15, 275.35, 275.35, 275.75, 275.65, 275.85, 
    276.25, 276.35, 276.15, 275.75, 275.65, 275.35, 275.15, 274.85, 275.05, 
    274.65, 274.45, 276.15, 276.55, 277.65, 275.95, 276.15, 275.95, 275.75, 
    276.05, 276.15, 276.15, 276.35, 275.65, 275.55, 275.15, 274.85, 274.85, 
    274.35, 274.45, 274.05, 273.95, 273.75, 273.35, 273.65, 273.75, 273.55, 
    273.15, 273.55, 273.75, 273.85, 274.25, 274.35, 274.75, 274.75, 274.85, 
    274.65, 274.55, 274.35, 274.75, 274.55, 274.95, 274.65, 274.75, 275.15, 
    275.35, 275.25, 274.55, 273.95, 273.95, 273.65, 272.95, 272.95, 273.05, 
    273.15, 273.35, 273.65, 273.85, 274.45, 274.55, 274.75, 274.95, 275.75, 
    275.85, 275.85, 275.65, 275.25, 275.75, 275.85, 275.75, 275.85, 275.75, 
    275.45, 275.45, 275.05, 274.95, 274.95, 275.65, 275.65, 275.65, 275.75, 
    276.65, 275.85, 276.55, 277.75, 277.55, 276.55, 277.55, 277.75, 277.75, 
    277.55, 277.25, 277.65, 275.75, 275.35, 275.75, 275.15, 274.15, 274.35, 
    274.55, 274.55, 274.95, 275.15, 275.25, 275.45, 274.95, 275.55, 275.55, 
    275.35, 276.15, 276.25, 276.65, 276.45, 276.45, 276.55, 276.65, 276.55, 
    276.45, 276.35, 277.45, 276.65, 275.85, 276.35, 276.25, 276.15, 276.65, 
    275.65, 275.25, 274.75, 274.25, 275.85, 275.15, 275.15, 276.15, 274.85, 
    275.25, 274.55, 273.95, 273.95, 274.05, 274.25, 273.75, 274.35, 273.95, 
    273.95, 275.35, 273.85, 273.85, 273.35, 272.95, 272.85, 273.55, 273.55, 
    273.45, 273.45, 273.65, 274.35, 275.25, 275.15, 275.35, 275.35, 276.75, 
    274.55, 274.45, 275.55, 276.05, 276.35, 276.45, 275.75, 276.05, 275.65, 
    276.15, 275.15, 275.65, 274.45, 275.15, 274.35, 275.05, 276.25, 275.75, 
    275.55, 274.85, 274.65, 274.85, 274.85, 274.45, 274.65, 274.85, 274.95, 
    274.85, 274.95, 275.15, 275.05, 275.25, 275.15, 275.25, 275.15, 275.25, 
    275.05, 275.15, 275.55, 275.65, 278.05, 276.95, 278.05, 276.05, 274.95, 
    275.55, 275.65, 275.55, 276.55, 275.75, 277.35, 276.95, 277.35, 276.15, 
    276.35, 275.15, 275.45, 275.85, 275.65, 275.85, 275.45, 276.25, 275.75, 
    276.15, 276.55, 275.95, 278.15, 276.25, 276.75, 277.15, 278.05, 278.15, 
    277.95, 277.85, 277.25, 276.85, 276.85, 276.65, 276.25, 276.05, 275.75, 
    275.35, 275.85, 275.85, 275.75, 275.55, 275.95, 276.05, 275.75, 275.55, 
    275.65, 275.65, 276.15, 276.55, 276.75, 278.25, 277.65, 278.75, 279.45, 
    276.45, 278.35, 280.65, 279.35, 277.25, 279.55, 279.25, 280.55, 280.65, 
    280.65, 279.25, 279.15, 280.05, 281.75, 279.05, 280.75, 280.45, 280.65, 
    281.85, 282.05, 282.55, 281.55, 282.05, 282.35, 280.75, 282.05, 281.45, 
    281.85, 281.45, 280.65, 281.35, 277.65, 277.65, 279.35, 279.05, 277.05, 
    277.05, 277.15, 277.65, 277.85, 278.35, 278.35, 277.95, 277.15, 276.45, 
    277.35, 278.85, 276.65, 275.65, 277.35, 276.05, 276.05, 276.05, 275.95, 
    276.05, 275.75, 275.55, 275.65, 277.05, 278.05, 275.35, 275.65, 276.25, 
    276.95, 277.65, 278.15, 277.05, 278.15, 276.85, 277.45, 276.55, 276.85, 
    276.75, 276.55, 275.95, 276.25, 276.95, 276.35, 275.95, 276.65, 276.75, 
    278.15, 277.65, 276.75, 276.65, 276.35, 277.85, 279.35, 276.45, 277.45, 
    277.75, 278.35, 279.05, 277.35, 277.25, 278.75, 278.25, 277.75, 277.95, 
    277.25, 278.25, 277.55, 277.55, 277.25, 277.75, 277.75, 277.45, 277.05, 
    276.75, 276.45, 276.55, 276.35, 277.25, 277.15, 277.15, 280.35, 280.75, 
    280.15, 278.95, 279.75, 278.85, 278.55, 277.75, 277.75, 276.55, 277.15, 
    276.85, 276.55, 276.55, 276.35, 276.35, 276.35, 276.45, 276.45, 276.45, 
    276.35, 276.35, 276.35, 276.75, 276.85, 276.45, 276.55, 276.65, 277.35, 
    277.65, 277.35, 277.25, 276.85, 277.65, 277.55, 276.75, 277.25, 277.15, 
    276.65, 276.45, 276.55, 276.65, 276.45, 276.05, 275.75, 275.75, 275.65, 
    275.65, 275.45, 275.55, 275.45, 275.45, 275.45, 275.25, 275.15, 275.05, 
    275.25, 275.45, 275.65, 275.45, 275.35, 275.05, 274.95, 275.05, 275.15, 
    275.25, 275.15, 275.15, 275.15, 275.05, 275.05, 275.05, 275.15, 274.95, 
    274.95, 275.35, 275.45, 275.25, 275.05, 275.05, 274.85, 275.05, 275.85, 
    275.25, 275.05, 274.75, 274.65, 275.75, 275.25, 275.45, 276.85, 277.85, 
    278.35, 278.45, 278.25, 278.25, 277.55, 277.55, 276.85, 277.25, 277.45, 
    276.65, 277.85, 277.65, 277.65, 277.85, 277.55, 277.15, 277.05, 277.05, 
    276.15, 276.45, 277.05, 276.85, 277.45, 277.45, 277.15, 277.25, 278.25, 
    277.85, 277.85, 278.35, 277.15, 277.85, 276.95, 276.55, 276.25, 276.75, 
    276.35, 275.95, 275.85, 275.35, 274.85, 274.65, 274.55, 274.35, 274.25, 
    274.35, 274.35, 274.35, 274.35, 274.35, 274.55, 274.45, 274.45, 274.35, 
    274.45, 274.45, 274.45, 274.25, 274.25, 274.45, 274.35, 274.45, 274.55, 
    274.25, 274.35, 274.35, 274.35, 274.45, 274.35, 274.35, 274.35, 274.35, 
    274.45, 274.35, 273.95, 273.65, 273.85, 273.55, 273.35, 273.35, 273.35, 
    273.25, 273.15, 273.15, 273.05, 272.85, 272.55, 274.15, 274.65, 274.35, 
    274.35, 274.15, 273.95, 274.15, 274.25, 274.55, 274.65, 274.65, 274.75, 
    275.35, 275.25, 275.25, 274.55, 274.45, 275.05, 275.25, 275.05, 275.35, 
    275.15, 275.05, 274.85, 274.95, 274.65, 274.85, 275.45, 276.05, 276.25, 
    276.05, 276.15, 276.25, 275.85, 276.45, 276.15, 275.85, 275.65, 275.85, 
    276.25, 276.65, 276.85, 276.75, 276.85, 276.55, 276.55, 276.45, 276.55, 
    276.25, 276.15, 276.05, 275.95, 275.85, 275.75, 275.95, 276.05, 276.15, 
    276.25, 276.05, 276.25, 275.75, 275.55, 275.35, 275.15, 274.25, 274.05, 
    274.35, 274.25, 274.15, 274.25, 273.95, 273.95, 274.15, 274.05, 273.95, 
    273.85, 273.85, 273.85, 274.15, 274.05, 273.45, 274.75, 273.75, 274.15, 
    273.55, 273.45, 273.75, 273.85, 273.85, 274.55, 274.85, 274.75, 274.75, 
    274.55, 274.85, 274.95, 274.75, 274.75, 274.65, 274.65, 274.55, 274.65, 
    274.55, 275.05, 274.65, 274.85, 275.05, 274.95, 275.05, 274.85, 275.15, 
    274.65, 274.75, 275.05, 275.05, 274.85, 275.05, 274.75, 274.25, 274.05, 
    273.05, 273.15, 273.45, 273.65, 273.95, 274.15, 274.15, 274.15, 274.35, 
    274.95, 274.95, 274.75, 274.65, 274.75, 274.85, 275.25, 274.95, 275.05, 
    274.65, 274.65, 274.65, 274.95, 274.55, 274.35, 274.55, 274.25, 274.05, 
    273.65, 274.35, 274.65, 274.85, 274.95, 275.15, 275.25, 275.75, 275.95, 
    276.15, 277.25, 277.25, 277.65, 277.75, 278.45, 277.45, 278.75, 277.75, 
    277.65, 277.25, 277.05, 277.65, 277.85, 277.45, 277.05, 275.75, 276.15, 
    276.75, 277.45, 277.65, 277.75, 277.25, 277.15, 276.65, 276.95, 276.15, 
    275.95, 275.85, 276.45, 276.05, 275.75, 275.55, 275.55, 275.35, 275.15, 
    275.05, 274.85, 274.45, 274.55, 274.65, 274.65, 275.35, 275.65, 276.05, 
    276.35, 276.15, 276.65, 276.75, 277.15, 277.15, 276.95, 276.85, 277.95, 
    277.25, 277.35, 277.25, 277.35, 275.15, 275.65, 273.85, 274.25, 274.55, 
    273.85, 273.45, 274.35, 275.05, 274.65, 274.25, 275.35, 275.25, 275.05, 
    276.65, 275.65, 276.45, 276.75, 276.95, 276.65, 276.55, 276.65, 276.75, 
    276.85, 276.35, 275.75, 275.85, 275.15, 275.15, 275.25, 275.25, 275.15, 
    274.95, 275.35, 274.65, 274.75, 274.35, 274.25, 273.95, 273.55, 273.45, 
    273.15, 273.45, 273.15, 272.95, 273.25, 273.65, 273.75, 273.85, 273.95, 
    274.45, 274.75, 274.75, 274.35, 274.75, 275.15, 275.25, 275.25, 275.75, 
    275.75, 275.55, 275.85, 275.95, 276.35, 276.95, 276.45, 276.15, 276.05, 
    276.35, 276.35, 276.25, 275.85, 275.95, 276.25, 276.25, 276.25, 276.35, 
    276.45, 276.35, 276.45, 276.25, 276.35, 276.65, 276.85, 277.45, 277.55, 
    277.45, 277.25, 277.65, 276.85, 276.95, 276.45, 275.65, 275.35, 275.15, 
    275.05, 274.85, 274.55, 274.75, 274.85, 274.95, 274.75, 274.85, 274.95, 
    275.15, 275.05, 275.55, 275.15, 275.35, 275.75, 275.65, 275.25, 274.95, 
    274.75, 274.75, 274.15, 273.95, 273.45, 272.85, 272.55, 272.25, 272.15, 
    271.65, 271.75, 271.95, 271.75, 272.05, 272.05, 272.15, 272.65, 272.85, 
    273.35, 272.85, 272.65, 273.15, 273.25, 273.05, 273.35, 273.35, 272.95, 
    272.85, 272.85, 272.85, 272.75, 272.35, 272.65, 272.95, 273.25, 273.15, 
    273.15, 273.85, 274.05, 273.45, 273.95, 274.25, 274.35, 274.55, 274.45, 
    274.55, 274.55, 273.45, 273.65, 274.05, 273.95, 273.65, 273.25, 272.75, 
    273.55, 273.55, 273.65, 273.55, 273.65, 273.85, 273.95, 273.95, 274.05, 
    274.35, 274.55, 274.45, 275.35, 274.75, 274.75, 274.75, 275.05, 275.05, 
    274.75, 275.65, 275.25, 275.25, 275.35, 275.55, 275.45, 275.55, 275.35, 
    275.45, 274.75, 274.35, 273.65, 274.25, 273.75, 274.05, 274.15, 274.45, 
    274.35, 274.05, 274.95, 275.15, 274.25, 274.95, 274.45, 273.25, 273.45, 
    271.85, 271.75, 271.85, 270.95, 270.75, 271.05, 271.85, 273.15, 274.55, 
    275.05, 275.95, 276.05, 276.15, 276.35, 276.15, 276.05, 275.85, 276.05, 
    276.05, 276.15, 276.15, 276.15, 276.45, 276.25, 276.65, 276.55, 276.25, 
    276.15, 273.65, 273.15, 273.55, 274.55, 275.15, 275.15, 274.95, 274.95, 
    274.85, 275.05, 275.15, 275.65, 275.85, 275.95, 275.85, 276.15, 276.15, 
    276.25, 276.25, 276.25, 275.85, 275.75, 275.65, 275.45, 275.85, 275.85, 
    275.55, 275.95, 275.95, 276.05, 275.95, 276.75, 276.45, 276.25, 276.95, 
    276.65, 277.75, 278.35, 277.45, 277.75, 277.55, 277.55, 277.35, 277.25, 
    277.55, 277.25, 277.35, 277.35, 277.25, 276.45, 276.95, 276.05, 275.05, 
    274.55, 274.35, 274.55, 274.65, 274.75, 275.75, 275.25, 275.25, 275.95, 
    276.55, 276.75, 276.55, 276.85, 277.05, 276.95, 277.65, 277.25, 276.85, 
    276.85, 277.05, 276.85, 276.65, 276.45, 275.95, 275.95, 276.45, 277.95, 
    277.75, 277.05, 277.05, 276.65, 276.75, 276.45, 276.55, 276.95, 276.45, 
    278.95, 277.85, 278.15, 278.25, 278.85, 278.25, 277.85, 278.15, 277.85, 
    277.65, 277.25, 277.35, 277.45, 277.45, 277.75, 277.95, 277.25, 276.65, 
    277.25, 278.55, 279.75, 278.45, 279.55, 280.95, 280.65, 280.55, 281.65, 
    277.55, 279.25, 278.45, 278.65, 277.95, 277.75, 277.15, 277.25, 276.25, 
    276.35, 276.65, 277.35, 277.15, 276.75, 277.35, 277.75, 278.75, 276.95, 
    277.45, 279.65, 278.25, 277.35, 276.95, 276.45, 276.85, 277.75, 278.05, 
    277.65, 277.05, 276.45, 276.65, 277.25, 277.75, 277.25, 276.95, 276.75, 
    275.85, 275.55, 276.55, 276.15, 276.05, 276.35, 276.75, 277.15, 276.75, 
    276.15, 276.15, 275.25, 274.65, 273.75, 273.25, 272.55, 272.75, 272.65, 
    272.55, 272.85, 273.05, 273.15, 273.25, 273.45, 273.15, 272.75, 272.75, 
    272.75, 272.75, 273.05, 273.25, 273.85, 274.05, 274.25, 274.75, 275.15, 
    275.35, 275.55, 275.45, 274.55, 274.55, 273.55, 273.45, 273.05, 272.65, 
    272.15, 271.95, 272.55, 272.25, 272.75, 272.75, 272.45, 272.35, 272.85, 
    272.65, 272.45, 272.05, 272.35, 271.95, 271.95, 272.05, 272.05, 272.05, 
    272.35, 272.55, 272.85, 273.05, 273.15, 273.45, 273.85, 273.85, 273.95, 
    274.15, 274.45, 274.75, 274.55, 274.85, 274.85, 274.85, 274.75, 274.55, 
    274.05, 274.55, 275.05, 274.25, 273.75, 273.45, 273.35, 273.05, 272.95, 
    273.15, 272.95, 272.85, 272.85, 272.75, 272.65, 272.25, 272.45, 272.65, 
    272.75, 272.95, 272.95, 273.15, 272.95, 272.75, 272.65, 271.95, 271.15, 
    271.85, 271.85, 271.35, 271.75, 271.55, 271.65, 271.95, 271.75, 271.85, 
    271.75, 271.55, 272.05, 272.15, 271.85, 271.95, 271.95, 272.25, 272.05, 
    271.55, 272.05, 271.45, 271.25, 271.05, 271.35, 271.05, 270.55, 270.25, 
    269.95, 270.35, 271.35, 271.35, 271.55, 272.05, 272.25, 272.25, 272.35, 
    272.35, 272.15, 272.15, 272.05, 272.15, 272.05, 272.35, 272.65, 272.65, 
    272.65, 272.85, 273.05, 272.55, 272.25, 272.25, 272.25, 272.05, 271.05, 
    272.05, 271.95, 271.95, 272.05, 272.25, 272.25, 272.35, 272.45, 272.35, 
    272.25, 272.35, 272.45, 272.45, 272.55, 272.65, 272.55, 272.65, 272.75, 
    272.75, 272.65, 272.75, 272.85, 273.05, 273.15, 273.25, 273.15, 273.05, 
    273.05, 272.95, 272.85, 272.95, 272.95, 272.95, 273.05, 273.15, 273.15, 
    272.95, 272.85, 272.55, 272.55, 271.65, 272.55, 273.15, 273.15, 273.65, 
    273.45, 272.95, 271.55, 271.35, 272.75, 272.15, 272.05, 272.35, 272.35, 
    272.25, 271.35, 271.55, 271.45, 271.45, 271.35, 271.15, 271.15, 271.05, 
    270.95, 272.65, 272.45, 272.25, 272.05, 271.95, 272.35, 272.55, 272.35, 
    272.65, 272.95, 273.05, 273.15, 273.35, 273.25, 272.45, 272.45, 273.85, 
    273.85, 273.85, 273.25, 274.05, 274.35, 274.15, 274.35, 272.95, 274.75, 
    275.05, 274.75, 274.45, 274.15, 274.05, 274.25, 273.75, 273.85, 274.35, 
    274.15, 274.45, 274.65, 274.55, 274.75, 274.75, 275.05, 275.35, 276.05, 
    276.65, 275.85, 274.75, 274.75, 274.25, 274.25, 274.15, 273.95, 273.75, 
    273.85, 273.75, 273.65, 273.65, 273.45, 273.35, 273.05, 273.25, 273.35, 
    273.35, 272.95, 272.85, 272.95, 273.15, 273.25, 273.35, 273.45, 273.45, 
    273.45, 273.45, 273.45, 273.55, 273.65, 273.85, 273.95, 273.85, 273.45, 
    273.65, 272.95, 272.85, 272.95, 273.15, 274.15, 274.45, 274.45, 274.35, 
    274.25, 274.65, 275.55, 275.15, 274.95, 274.45, 274.35, 273.55, 273.45, 
    273.15, 272.55, 272.35, 272.05, 272.25, 272.15, 271.95, 272.15, 272.55, 
    272.95, 271.95, 271.95, 272.25, 272.65, 272.75, 272.95, 273.35, 272.95, 
    272.65, 273.15, 272.45, 272.95, 272.45, 272.35, 271.95, 272.55, 272.25, 
    271.55, 272.55, 272.55, 272.45, 273.25, 271.45, 271.05, 271.25, 272.05, 
    272.15, 271.25, 270.85, 270.55, 270.85, 270.95, 270.95, 270.85, 270.45, 
    270.25, 270.05, 269.65, 269.15, 268.55, 269.35, 271.05, 271.55, 271.75, 
    271.75, 271.85, 271.25, 271.25, 271.75, 272.45, 272.45, 272.85, 272.75, 
    273.15, 273.25, 273.45, 273.75, 273.85, 274.05, 273.85, 273.45, 273.95, 
    273.75, 273.45, 273.75, 273.75, 273.75, 273.85, 274.05, 274.15, 274.25, 
    274.35, 274.35, 274.25, 274.15, 274.25, 274.25, 274.65, 275.05, 275.15, 
    275.15, 275.05, 274.95, 275.05, 274.45, 274.05, 273.85, 273.75, 273.95, 
    274.25, 273.05, 271.05, 270.85, 270.65, 270.45, 270.35, 270.15, 270.05, 
    269.85, 269.05, 269.95, 270.25, 270.65, 270.65, 270.55, 271.15, 271.05, 
    270.45, 270.75, 270.95, 270.15, 270.25, 271.15, 270.85, 270.45, 270.35, 
    269.95, 270.15, 270.35, 270.25, 270.05, 270.35, 270.35, 270.55, 270.55, 
    269.75, 271.95, 272.05, 271.65, 271.65, 271.45, 271.45, 271.45, 271.35, 
    270.65, 270.85, 270.25, 270.25, 269.95, 270.25, 270.15, 269.65, 269.45, 
    268.75, 268.95, 269.05, 268.95, 270.65, 269.55, 269.85, 270.95, 271.05, 
    270.85, 270.25, 270.65, 270.15, 270.85, 274.25, 271.15, 269.55, 271.35, 
    273.05, 271.55, 271.25, 271.05, 272.05, 272.35, 272.35, 272.55, 272.75, 
    272.85, 273.05, 273.35, 273.95, 274.15, 274.45, 274.15, 275.55, 275.95, 
    276.95, 276.75, 276.05, 276.65, 277.25, 277.05, 275.85, 275.75, 274.25, 
    274.35, 273.85, 274.05, 274.05, 273.25, 274.75, 275.15, 274.75, 273.75, 
    273.65, 273.35, 273.15, 273.75, 273.45, 274.95, 274.05, 274.15, 273.25, 
    273.25, 273.65, 273.35, 273.35, 273.35, 273.35, 273.35, 273.35, 273.35, 
    273.65, 273.55, 273.55, 273.65, 273.75, 273.75, 273.65, 274.05, 274.35, 
    274.95, 274.65, 274.55, 274.35, 274.15, 274.15, 274.05, 273.95, 273.85, 
    274.15, 274.35, 274.55, 274.75, 275.15, 275.05, 275.15, 275.35, 275.55, 
    275.95, 276.05, 276.05, 276.05, 275.95, 276.05, 276.15, 276.05, 275.85, 
    275.85, 275.85, 275.65, 275.75, 275.65, 275.35, 275.95, 275.35, 275.35, 
    275.45, 274.95, 275.05, 275.45, 275.55, 275.45, 275.85, 275.15, 274.95, 
    274.85, 274.65, 274.25, 273.55, 273.25, 273.05, 273.15, 273.25, 273.15, 
    272.95, 272.75, 272.75, 272.65, 272.45, 272.25, 272.25, 271.85, 270.85, 
    270.35, 269.95, 269.95, 270.25, 270.45, 270.45, 270.95, 271.05, 271.15, 
    272.15, 271.65, 271.65, 271.75, 271.55, 271.95, 272.15, 272.95, 273.15, 
    273.05, 273.35, 273.75, 274.05, 274.15, 274.35, 274.35, 274.45, 274.35, 
    274.65, 274.75, 275.05, 275.05, 275.05, 275.25, 275.85, 276.15, 276.15, 
    276.25, 276.35, 276.25, 276.05, 275.85, 275.85, 275.85, 275.65, 275.85, 
    275.75, 275.85, 275.65, 275.65, 275.45, 275.75, 275.55, 275.75, 275.65, 
    275.75, 275.45, 275.25, 275.85, 275.95, 275.65, 275.35, 275.75, 275.65, 
    276.05, 276.65, 276.45, 276.85, 277.05, 276.85, 276.65, 276.45, 276.45, 
    276.25, 276.45, 276.85, 275.95, 275.65, 275.35, 276.45, 276.75, 275.25, 
    274.45, 273.45, 273.15, 273.35, 273.35, 273.05, 272.95, 272.85, 272.75, 
    272.65, 272.55, 272.45, 272.25, 272.05, 272.35, 271.95, 271.75, 271.55, 
    271.35, 271.45, 271.45, 271.15, 271.35, 271.25, 271.25, 271.25, 271.15, 
    271.35, 271.45, 271.45, 271.65, 271.75, 271.85, 271.75, 272.15, 272.35, 
    272.55, 272.95, 273.05, 273.15, 273.45, 273.65, 274.05, 274.15, 274.05, 
    274.35, 274.45, 274.95, 276.05, 275.65, 275.45, 275.45, 274.75, 274.95, 
    275.55, 275.55, 275.55, 275.25, 274.95, 274.85, 273.25, 272.95, 272.35, 
    272.05, 272.15, 272.25, 272.05, 272.15, 272.45, 274.05, 274.95, 274.65, 
    274.75, 274.75, 274.15, 273.85, 273.55, 274.55, 273.75, 273.65, 273.45, 
    272.65, 272.15, 272.15, 271.95, 272.05, 272.15, 272.25, 272.45, 272.55, 
    272.65, 272.95, 272.75, 272.65, 272.95, 273.15, 273.55, 273.55, 273.45, 
    273.45, 273.45, 273.35, 273.35, 273.45, 273.35, 273.25, 272.95, 273.25, 
    273.55, 273.15, 272.95, 272.55, 273.45, 272.45, 271.95, 270.95, 271.75, 
    272.15, 272.15, 272.65, 272.85, 272.95, 273.05, 273.15, 273.35, 273.65, 
    273.95, 274.35, 274.35, 274.75, 274.25, 273.85, 273.35, 273.05, 272.95, 
    272.35, 271.95, 272.15, 272.05, 272.45, 272.85, 273.25, 273.85, 273.45, 
    273.35, 273.55, 273.65, 273.65, 273.45, 273.65, 273.75, 273.15, 273.75, 
    273.85, 271.85, 272.35, 273.45, 274.15, 274.45, 274.55, 274.25, 274.55, 
    274.75, 274.25, 274.45, 274.55, 274.65, 274.75, 274.85, 274.85, 274.85, 
    274.75, 274.65, 274.45, 274.35, 273.75, 274.05, 274.05, 274.25, 274.55, 
    274.95, 274.95, 274.95, 274.85, 274.75, 274.75, 274.95, 274.85, 275.05, 
    275.75, 275.85, 275.95, 275.75, 275.55, 275.25, 274.35, 275.35, 275.45, 
    275.15, 274.95, 274.95, 275.05, 275.25, 275.15, 275.05, 275.15, 274.75, 
    274.75, 274.95, 274.75, 274.35, 274.05, 273.75, 273.75, 273.95, 273.75, 
    273.75, 273.35, 272.75, 272.45, 272.75, 273.45, 273.45, 273.45, 273.65, 
    275.05, 275.65, 277.25, 276.05, 274.55, 273.65, 273.15, 272.55, 272.35, 
    271.95, 271.65, 271.25, 271.15, 271.15, 270.95, 270.85, 270.45, 270.35, 
    270.35, 270.55, 270.55, 270.65, 270.55, 270.85, 270.85, 270.95, 271.15, 
    271.35, 271.55, 271.75, 271.75, 272.05, 272.55, 273.55, 274.95, 275.05, 
    275.45, 275.45, 276.15, 276.15, 276.55, 276.25, 276.05, 275.75, 275.95, 
    276.25, 276.25, 276.05, 275.95, 275.85, 275.65, 275.45, 275.05, 274.95, 
    275.45, 275.35, 275.75, 275.45, 276.35, 276.45, 276.45, 276.25, 276.05, 
    276.15, 276.25, 275.95, 275.85, 275.45, 275.45, 275.45, 275.55, 275.65, 
    275.55, 275.45, 275.55, 275.45, 275.35, 275.45, 275.55, 275.75, 275.45, 
    275.55, 275.65, 275.55, 275.35, 275.45, 275.35, 275.45, 275.95, 275.85, 
    276.15, 275.95, 275.65, 275.65, 275.85, 275.95, 276.15, 275.75, 275.85, 
    275.85, 276.05, 275.75, 276.05, 274.25, 273.75, 273.35, 272.95, 272.55, 
    272.25, 272.25, 271.85, 271.85, 271.75, 271.75, 271.75, 271.55, 271.55, 
    271.65, 271.55, 271.65, 271.55, 271.55, 271.15, 271.05, 271.05, 271.05, 
    271.05, 271.05, 271.25, 271.95, 272.05, 272.25, 272.15, 272.05, 272.05, 
    272.25, 272.75, 273.05, 273.25, 273.15, 273.25, 273.05, 273.35, 273.45, 
    273.75, 274.05, 274.35, 274.15, 273.95, 273.95, 274.75, 274.95, 274.75, 
    273.65, 274.35, 274.55, 275.05, 274.95, 274.75, 274.95, 274.95, 275.05, 
    275.35, 275.35, 275.35, 275.25, 274.95, 275.15, 276.35, 276.35, 274.85, 
    274.35, 273.35, 272.55, 271.45, 271.15, 270.95, 270.85, 270.95, 270.55, 
    270.85, 271.15, 271.05, 271.05, 271.25, 270.25, 269.75, 270.05, 270.35, 
    270.45, 271.05, 272.45, 272.65, 272.75, 273.05, 273.45, 273.65, 273.95, 
    274.05, 274.35, 275.05, 275.15, 274.65, 275.55, 275.55, 275.65, 275.65, 
    276.45, 276.15, 275.75, 275.45, 275.25, 275.05, 274.85, 275.65, 275.45, 
    273.95, 272.65, 270.85, 270.75, 271.05, 271.05, 271.15, 271.25, 271.55, 
    271.25, 271.55, 271.35, 271.45, 271.65, 271.65, 271.55, 271.85, 271.85, 
    271.65, 271.65, 271.55, 271.45, 272.25, 272.85, 273.45, 273.85, 274.05, 
    273.95, 273.55, 273.15, 272.95, 272.85, 272.75, 272.55, 272.55, 272.85, 
    272.95, 272.45, 271.95, 272.35, 271.65, 271.95, 272.95, 273.05, 273.25, 
    273.35, 272.95, 273.15, 272.85, 272.55, 272.35, 273.05, 273.25, 273.35, 
    275.25, 275.75, 275.35, 275.05, 274.85, 274.65, 274.45, 275.05, 275.55, 
    275.45, 276.25, 276.05, 275.95, 275.65, 275.65, 275.65, 274.65, 274.85, 
    274.75, 273.45, 273.25, 272.05, 271.15, 271.05, 271.35, 271.85, 271.75, 
    271.45, 271.35, 271.45, 270.95, 271.05, 271.25, 272.05, 272.55, 271.65, 
    271.35, 271.35, 271.45, 271.85, 272.05, 272.35, 271.95, 271.95, 271.65, 
    271.55, 270.95, 270.25, 270.45, 270.45, 270.75, 270.85, 271.05, 270.95, 
    270.55, 270.75, 269.75, 269.45, 268.95, 268.55, 268.75, 268.35, 267.85, 
    267.85, 267.95, 267.95, 268.15, 268.15, 268.05, 268.15, 268.45, 268.35, 
    268.45, 268.55, 268.65, 268.85, 268.75, 268.75, 269.05, 269.65, 269.85, 
    270.25, 270.05, 271.05, 271.75, 271.65, 271.75, 271.85, 271.75, 272.05, 
    272.15, 272.15, 272.25, 272.25, 272.25, 271.75, 271.65, 271.75, 272.05, 
    271.75, 272.25, 272.35, 272.15, 272.35, 272.65, 272.95, 273.05, 273.15, 
    273.45, 273.55, 274.15, 274.55, 274.65, 274.95, 274.95, 274.95, 275.25, 
    275.35, 275.35, 275.45, 275.05, 274.45, 274.55, 274.35, 274.15, 274.65, 
    274.05, 274.25, 274.25, 272.95, 272.15, 270.45, 269.65, 270.25, 269.65, 
    269.95, 269.75, 269.95, 270.05, 270.15, 270.15, 269.75, 269.75, 269.15, 
    268.85, 269.25, 269.35, 269.15, 269.15, 269.15, 269.35, 269.25, 269.25, 
    269.05, 269.05, 268.95, 268.75, 268.85, 268.85, 268.75, 268.95, 268.85, 
    269.35, 269.45, 269.65, 269.85, 270.15, 270.15, 270.25, 269.85, 270.55, 
    271.85, 271.55, 271.75, 271.75, 271.85, 272.05, 272.05, 272.05, 272.05, 
    271.95, 271.65, 270.65, 270.45, 270.45, 270.55, 270.35, 270.95, 271.25, 
    271.65, 272.75, 272.55, 272.65, 272.75, 272.45, 272.55, 272.65, 272.75, 
    272.75, 272.25, 271.75, 270.65, 271.05, 271.85, 272.35, 272.95, 273.55, 
    274.25, 274.05, 274.55, 274.25, 274.15, 273.75, 273.85, 273.65, 274.05, 
    273.65, 274.05, 274.05, 274.35, 274.75, 274.75, 274.45, 274.95, 274.25, 
    273.85, 273.85, 274.25, 273.95, 273.95, 274.65, 274.95, 274.75, 274.55, 
    274.45, 274.55, 274.45, 274.35, 274.35, 274.25, 274.15, 275.05, 274.75, 
    274.85, 274.95, 275.15, 275.75, 274.85, 275.25, 275.35, 275.25, 274.85, 
    275.05, 275.05, 275.05, 274.25, 275.05, 274.75, 274.95, 275.15, 275.45, 
    275.75, 275.65, 275.65, 276.05, 275.85, 275.55, 275.25, 275.35, 275.25, 
    275.35, 275.55, 275.65, 275.35, 275.25, 274.75, 274.85, 274.75, 275.85, 
    274.75, 274.25, 274.25, 273.85, 272.65, 272.25, 272.35, 272.25, 272.15, 
    271.85, 271.75, 271.25, 270.85, 270.15, 269.75, 269.15, 268.65, 268.35, 
    267.95, 267.55, 267.15, 266.75, 266.35, 266.35, 265.95, 265.95, 265.65, 
    265.65, 265.55, 265.65, 265.55, 265.15, 264.75, 265.05, 265.15, 264.95, 
    265.65, 266.15, 266.85, 267.85, 268.35, 268.95, 269.45, 269.85, 270.55, 
    271.05, 271.45, 271.95, 272.25, 272.45, 273.25, 273.35, 273.25, 273.65, 
    273.95, 274.25, 274.65, 275.45, 273.85, 274.85, 273.95, 274.15, 274.65, 
    275.05, 274.35, 274.05, 273.85, 273.95, 274.25, 274.05, 273.65, 273.65, 
    272.95, 274.45, 275.45, 275.55, 275.75, 275.95, 274.15, 274.35, 273.75, 
    273.15, 273.05, 272.95, 273.85, 273.65, 274.05, 274.15, 274.05, 273.25, 
    273.55, 273.45, 273.95, 274.15, 274.15, 273.95, 274.05, 274.15, 274.35, 
    274.65, 275.05, 273.65, 273.95, 273.85, 273.95, 273.65, 273.15, 273.05, 
    273.05, 273.05, 273.05, 272.85, 272.75, 272.55, 272.15, 272.05, 272.45, 
    272.45, 271.35, 272.75, 273.15, 273.25, 274.15, 274.65, 275.15, 274.95, 
    275.65, 275.15, 275.15, 275.05, 274.65, 274.35, 274.35, 274.35, 274.55, 
    274.95, 274.95, 275.15, 274.85, 274.25, 274.35, 274.15, 273.95, 274.05, 
    274.05, 274.15, 274.15, 274.45, 274.45, 274.35, 274.45, 274.45, 274.25, 
    274.35, 274.35, 274.25, 274.25, 274.65, 274.75, 274.75, 274.95, 274.45, 
    274.25, 274.55, 274.45, 273.55, 273.35, 273.45, 272.95, 272.85, 272.25, 
    272.55, 272.65, 272.65, 272.35, 272.15, 271.45, 271.35, 271.35, 271.15, 
    271.15, 271.25, 271.25, 271.05, 270.95, 271.05, 270.95, 270.65, 270.55, 
    270.55, 270.15, 270.35, 270.65, 270.65, 270.55, 270.55, 270.15, 269.55, 
    269.35, 269.75, 269.15, 270.35, 270.05, 269.75, 269.25, 268.85, 268.55, 
    268.25, 267.45, 266.75, 266.35, 266.05, 266.05, 265.85, 265.95, 266.25, 
    266.45, 266.75, 266.85, 266.85, 266.85, 266.45, 266.55, 266.55, 266.75, 
    266.15, 265.95, 266.25, 267.05, 267.55, 267.75, 268.05, 268.15, 268.05, 
    268.15, 267.85, 267.05, 266.35, 266.45, 266.15, 265.35, 264.95, 266.75, 
    267.05, 267.15, 267.25, 266.65, 266.25, 265.65, 266.25, 266.45, 265.85, 
    266.45, 267.05, 266.95, 266.85, 266.85, 267.35, 267.25, 267.75, 267.55, 
    267.15, 267.75, 268.05, 267.65, 267.75, 267.85, 267.75, 268.35, 268.05, 
    268.35, 268.05, 268.55, 268.15, 269.65, 269.05, 268.95, 268.55, 268.25, 
    268.15, 268.25, 269.35, 269.95, 269.45, 269.85, 270.15, 271.05, 270.55, 
    270.35, 270.85, 271.65, 271.75, 271.25, 270.45, 270.85, 270.35, 269.85, 
    270.15, 271.15, 271.75, 271.35, 271.15, 271.35, 271.55, 271.55, 271.55, 
    271.55, 271.15, 271.05, 271.75, 272.15, 272.35, 271.95, 272.05, 272.05, 
    271.95, 271.95, 271.95, 271.85, 271.85, 271.75, 271.95, 272.15, 271.85, 
    272.15, 272.15, 271.95, 272.15, 272.05, 271.75, 272.25, 271.95, 272.15, 
    271.35, 271.85, 272.25, 272.45, 272.85, 272.55, 272.85, 272.55, 272.75, 
    272.45, 272.75, 272.65, 272.45, 272.15, 271.95, 270.85, 269.85, 269.35, 
    269.15, 269.15, 268.95, 268.75, 268.75, 268.65, 268.75, 268.75, 268.85, 
    268.65, 268.85, 268.75, 268.15, 267.95, 267.85, 268.15, 268.25, 268.45, 
    268.75, 269.35, 269.65, 270.15, 270.85, 271.15, 271.35, 271.75, 272.25, 
    272.55, 272.65, 272.65, 272.75, 272.55, 272.65, 272.55, 272.55, 272.85, 
    272.95, 272.95, 273.05, 272.95, 272.85, 272.45, 272.45, 272.65, 272.85, 
    273.05, 273.45, 273.75, 273.85, 274.15, 274.05, 274.15, 274.35, 274.45, 
    274.65, 274.85, 274.95, 274.95, 274.75, 273.85, 274.75, 274.95, 275.05, 
    275.15, 275.35, 275.25, 275.25, 275.25, 275.35, 276.15, 275.95, 275.05, 
    274.05, 274.15, 273.75, 273.25, 272.55, 271.85, 271.55, 271.45, 271.35, 
    271.35, 271.55, 271.65, 271.35, 271.25, 271.45, 271.25, 271.25, 271.05, 
    270.95, 270.95, 271.15, 271.05, 271.25, 271.35, 271.25, 271.25, 271.25, 
    271.25, 271.35, 271.55, 271.65, 271.45, 271.15, 271.25, 271.45, 271.65, 
    271.85, 272.05, 272.25, 272.45, 272.45, 272.55, 272.25, 272.25, 272.35, 
    272.25, 272.15, 272.05, 272.75, 273.05, 273.35, 273.95, 273.95, 274.25, 
    274.05, 273.55, 273.95, 274.05, 274.25, 273.75, 273.25, 273.55, 273.85, 
    273.25, 273.45, 273.45, 273.45, 273.45, 273.75, 273.25, 273.75, 273.15, 
    272.85, 272.85, 272.85, 272.85, 272.85, 272.65, 272.95, 273.05, 272.95, 
    272.95, 272.85, 272.65, 272.45, 272.15, 272.55, 272.55, 272.85, 272.95, 
    272.95, 273.25, 273.25, 273.15, 273.25, 273.35, 273.25, 273.25, 273.25, 
    273.35, 273.35, 273.35, 273.35, 273.25, 273.25, 273.15, 273.15, 273.35, 
    273.35, 273.25, 273.15, 273.25, 273.15, 273.25, 273.25, 273.15, 273.25, 
    273.15, 273.05, 273.15, 272.95, 272.95, 272.95, 272.95, 273.35, 273.35, 
    273.15, 272.95, 272.95, 272.85, 272.95, 272.75, 272.65, 271.95, 271.75, 
    271.95, 272.15, 272.35, 272.35, 272.75, 272.95, 273.05, 273.45, 273.45, 
    273.55, 273.55, 273.55, 273.55, 273.45, 274.25, 273.85, 274.05, 274.45, 
    274.75, 274.65, 274.35, 274.35, 274.05, 273.75, 273.55, 273.25, 273.75, 
    274.25, 274.55, 274.55, 274.25, 274.35, 274.45, 274.35, 274.45, 274.35, 
    274.25, 274.45, 274.45, 274.55, 274.45, 274.45, 274.25, 274.25, 274.35, 
    274.15, 274.25, 274.05, 273.85, 273.65, 273.35, 273.55, 274.05, 274.05, 
    273.85, 273.95, 273.75, 273.85, 273.95, 273.95, 274.05, 274.15, 274.25, 
    274.25, 274.35, 274.45, 274.45, 274.55, 274.65, 274.75, 275.15, 275.35, 
    275.25, 275.05, 274.85, 274.65, 274.45, 274.65, 274.45, 274.65, 274.55, 
    274.55, 274.15, 274.45, 274.15, 274.55, 274.85, 273.95, 273.65, 273.65, 
    273.85, 273.75, 273.65, 273.35, 273.65, 274.05, 273.75, 273.65, 273.75, 
    273.75, 273.55, 273.55, 273.55, 273.55, 273.35, 273.35, 273.25, 273.15, 
    273.15, 273.05, 273.05, 273.25, 273.25, 273.15, 273.05, 272.95, 272.85, 
    272.75, 272.75, 272.45, 272.55, 272.35, 272.05, 272.15, 272.05, 271.55, 
    271.65, 271.15, 271.35, 271.25, 270.95, 271.65, 271.75, 271.35, 270.65, 
    270.65, 270.45, 271.15, 271.45, 271.75, 271.85, 272.05, 272.35, 272.45, 
    271.35, 271.45, 271.55, 271.85, 272.05, 272.45, 272.55, 272.85, 272.65, 
    272.75, 272.45, 272.55, 272.65, 272.85, 272.65, 272.45, 272.65, 272.35, 
    272.35, 272.25, 272.25, 272.45, 272.15, 272.25, 271.65, 271.45, 271.65, 
    271.75, 271.55, 271.15, 271.05, 270.55, 269.35, 268.45, 267.35, 268.05, 
    269.15, 269.95, 269.65, 269.65, 269.65, 270.05, 269.35, 269.15, 269.65, 
    269.15, 269.95, 269.55, 270.15, 269.75, 268.45, 269.75, 270.45, 270.55, 
    270.55, 271.05, 270.85, 270.65, 271.05, 271.05, 270.75, 270.75, 270.45, 
    270.85, 270.75, 270.35, 269.65, 270.15, 269.95, 269.95, 270.25, 269.95, 
    269.95, 269.95, 267.75, 267.45, 267.75, 268.85, 268.15, 267.55, 267.55, 
    267.75, 268.45, 267.05, 267.45, 265.85, 266.35, 265.65, 266.05, 265.85, 
    266.25, 267.15, 267.55, 267.75, 268.45, 268.55, 268.65, 269.95, 269.15, 
    269.65, 270.45, 270.25, 268.65, 268.05, 267.65, 264.35, 266.45, 266.25, 
    266.25, 266.75, 267.75, 267.25, 267.95, 267.45, 267.65, 267.65, 267.45, 
    267.65, 268.45, 267.45, 266.65, 265.85, 266.55, 266.55, 266.95, 267.45, 
    267.25, 266.15, 265.95, 266.55, 266.35, 266.05, 265.55, 265.75, 264.95, 
    263.55, 263.15, 264.85, 264.45, 264.45, 263.55, 263.55, 263.95, 263.95, 
    264.35, 264.45, 264.45, 264.75, 264.45, 264.45, 263.05, 264.85, 265.15, 
    265.45, 265.55, 264.95, 264.65, 263.95, 265.05, 265.45, 263.85, 263.05, 
    263.25, 263.55, 263.25, 264.15, 264.95, 265.95, 266.75, 267.05, 267.45, 
    266.65, 265.15, 264.35, 263.85, 263.65, 264.05, 263.85, 265.75, 264.85, 
    266.05, 265.55, 266.25, 265.15, 265.35, 264.25, 265.25, 266.35, 267.15, 
    267.05, 266.95, 266.75, 266.65, 265.55, 264.15, 263.15, 264.05, 265.25, 
    264.65, 264.85, 264.25, 264.45, 264.05, 264.45, 265.65, 265.95, 264.35, 
    264.85, 263.95, 265.05, 266.25, 266.25, 266.05, 266.35, 266.25, 265.55, 
    265.35, 265.45, 265.25, 265.85, 265.85, 266.55, 265.65, 265.05, 266.35, 
    266.75, 265.85, 265.85, 265.75, 265.85, 265.85, 265.85, 264.95, 264.85, 
    265.35, 263.35, 262.75, 264.85, 265.95, 266.55, 267.15, 266.75, 266.35, 
    265.85, 265.05, 263.85, 263.45, 263.65, 264.95, 264.75, 263.45, 263.25, 
    262.25, 262.25, 262.55, 261.95, 261.45, 261.85, 261.05, 261.95, 262.05, 
    261.45, 261.25, 261.25, 261.85, 260.65, 261.45, 260.85, 261.45, 261.75, 
    261.75, 261.85, 261.95, 261.75, 261.15, 260.45, 259.75, 258.95, 258.35, 
    258.35, 258.25, 258.85, 260.05, 261.75, 261.75, 262.25, 263.05, 264.05, 
    264.75, 265.45, 265.95, 266.25, 266.35, 266.45, 267.75, 267.85, 267.75, 
    267.95, 267.65, 267.75, 268.15, 268.35, 268.45, 268.25, 268.25, 267.05, 
    268.65, 268.95, 269.35, 269.45, 269.25, 270.05, 269.95, 270.15, 270.45, 
    270.15, 270.75, 270.75, 270.85, 270.85, 270.95, 270.75, 270.95, 270.85, 
    271.05, 271.05, 270.85, 271.25, 271.05, 271.25, 271.05, 270.95, 270.95, 
    270.35, 269.45, 267.25, 266.65, 265.85, 264.95, 264.65, 263.95, 263.15, 
    262.65, 262.15, 262.15, 262.35, 262.25, 262.05, 261.75, 261.65, 261.75, 
    262.15, 262.65, 262.95, 263.15, 263.35, 263.75, 264.35, 264.85, 265.15, 
    264.85, 264.45, 264.15, 263.05, 262.85, 263.25, 263.75, 264.35, 263.45, 
    262.45, 262.45, 261.75, 261.65, 261.15, 260.55, 259.65, 260.25, 259.95, 
    259.85, 257.15, 257.25, 257.45, 257.65, 258.05, 258.35, 258.55, 258.85, 
    259.25, 259.35, 259.45, 259.75, 259.85, 259.75, 259.95, 259.85, 259.75, 
    259.85, 259.95, 259.85, 259.95, 259.95, 259.85, 259.75, 258.65, 258.55, 
    258.35, 258.35, 257.95, 257.75, 257.75, 257.85, 257.85, 258.05, 258.05, 
    258.15, 258.55, 258.45, 258.55, 258.45, 258.35, 258.35, 258.35, 258.55, 
    258.85, 259.05, 259.25, 259.45, 259.85, 260.45, 261.35, 262.75, 264.15, 
    264.05, 264.45, 264.45, 263.95, 263.45, 263.05, 262.75, 263.35, 262.85, 
    261.75, 260.55, 261.45, 262.75, 263.15, 262.85, 262.65, 262.75, 263.05, 
    263.15, 263.25, 263.35, 263.35, 263.35, 263.45, 263.65, 263.75, 263.75, 
    263.95, 264.15, 264.35, 264.55, 263.75, 263.85, 263.85, 263.85, 263.65, 
    263.45, 263.15, 262.85, 262.65, 262.45, 262.35, 262.25, 263.05, 263.15, 
    262.95, 262.65, 262.65, 262.65, 262.65, 262.65, 262.75, 262.95, 263.05, 
    262.95, 262.75, 262.85, 262.85, 262.75, 262.65, 262.55, 262.35, 262.25, 
    262.25, 262.35, 262.65, 262.95, 262.85, 263.25, 263.45, 263.55, 263.55, 
    263.55, 263.55, 263.45, 263.35, 263.15, 263.15, 263.15, 263.15, 263.25, 
    263.25, 263.15, 263.15, 263.15, 263.15, 263.05, 262.85, 262.55, 262.35, 
    262.25, 261.75, 261.65, 261.65, 261.55, 261.55, 261.45, 261.25, 261.25, 
    261.25, 261.35, 261.35, 261.55, 261.65, 261.35, 261.15, 260.95, 260.75, 
    260.45, 260.15, 259.95, 259.65, 259.45, 259.15, 259.15, 258.95, 258.75, 
    258.55, 258.35, 258.05, 257.85, 257.75, 257.85, 258.05, 258.05, 257.95, 
    257.85, 256.85, 256.95, 257.25, 257.95, 258.45, 259.05, 259.35, 259.55, 
    259.95, 260.35, 260.75, 261.05, 262.55, 262.95, 263.45, 263.95, 264.35, 
    264.65, 264.95, 265.15, 265.55, 266.05, 266.85, 267.65, 267.65, 268.05, 
    268.45, 268.75, 268.95, 269.15, 269.35, 270.65, 270.65, 270.95, 270.75, 
    271.25, 271.15, 270.95, 271.25, 271.25, 271.25, 271.35, 271.55, 271.75, 
    271.85, 271.95, 271.85, 271.75, 271.85, 271.85, 271.75, 271.55, 272.05, 
    271.95, 270.05, 268.45, 268.95, 268.35, 267.85, 267.35, 266.55, 266.05, 
    265.25, 265.05, 264.85, 265.45, 266.25, 265.65, 266.05, 267.65, 266.85, 
    267.05, 267.95, 268.55, 269.15, 269.15, 269.85, 270.35, 270.65, 270.95, 
    270.95, 271.15, 271.35, 271.35, 271.15, 270.55, 270.35, 270.65, 270.45, 
    269.95, 270.05, 270.25, 270.15, 270.05, 271.55, 271.25, 271.65, 270.25, 
    270.55, 270.15, 270.95, 271.25, 271.35, 271.65, 271.45, 271.55, 271.35, 
    271.45, 271.65, 271.85, 271.95, 271.85, 271.95, 271.95, 271.95, 271.95, 
    271.95, 271.85, 271.95, 272.15, 272.45, 272.25, 272.25, 272.45, 272.25, 
    272.35, 272.35, 272.25, 272.25, 271.95, 272.15, 271.95, 271.85, 271.35, 
    271.25, 271.25, 271.15, 271.05, 271.25, 271.75, 270.85, 270.55, 269.15, 
    269.75, 270.35, 270.25, 270.15, 270.05, 270.15, 270.25, 270.15, 270.35, 
    270.15, 270.35, 270.85, 271.05, 271.25, 271.25, 271.65, 272.25, 272.45, 
    272.55, 272.45, 272.45, 272.25, 271.85, 272.25, 272.35, 272.35, 272.45, 
    272.25, 272.25, 272.15, 272.15, 271.95, 271.95, 271.45, 271.05, 270.35, 
    269.85, 269.05, 268.65, 270.65, 269.75, 270.75, 271.05, 269.35, 269.95, 
    271.15, 271.35, 271.55, 272.05, 271.95, 272.05, 272.25, 272.65, 272.55, 
    272.85, 272.65, 272.95, 273.05, 273.35, 273.35, 273.35, 273.25, 273.35, 
    272.95, 272.95, 273.05, 272.95, 272.95, 273.05, 272.95, 273.05, 272.75, 
    272.85, 273.25, 272.75, 273.05, 272.35, 272.35, 273.45, 273.85, 273.55, 
    273.55, 272.95, 272.55, 272.15, 273.05, 271.65, 271.15, 271.45, 272.05, 
    271.55, 271.85, 271.85, 271.65, 271.65, 271.75, 271.65, 271.55, 271.55, 
    271.55, 271.35, 271.35, 271.25, 271.15, 271.35, 271.45, 271.55, 271.55, 
    271.35, 271.25, 271.05, 270.95, 271.65, 271.15, 270.35, 269.55, 269.55, 
    270.25, 269.95, 269.45, 270.45, 270.75, 269.85, 271.05, 270.55, 270.25, 
    270.05, 269.15, 270.15, 270.55, 271.15, 270.95, 271.45, 270.65, 271.15, 
    271.05, 271.35, 271.55, 270.75, 270.75, 270.65, 270.55, 269.75, 270.15, 
    270.35, 270.45, 270.75, 271.25, 271.75, 271.55, 271.15, 272.05, 271.15, 
    271.15, 271.05, 270.75, 270.55, 270.35, 270.95, 271.15, 271.35, 271.35, 
    271.15, 271.25, 270.95, 270.85, 270.75, 271.35, 271.05, 270.45, 269.65, 
    269.35, 269.55, 270.25, 270.95, 271.15, 271.35, 271.35, 271.15, 270.35, 
    269.65, 268.75, 268.25, 267.65, 267.05, 266.75, 266.15, 265.95, 265.75, 
    264.95, 265.05, 264.95, 264.55, 263.85, 262.65, 263.15, 261.95, 261.55, 
    262.85, 262.95, 263.35, 263.45, 263.75, 263.45, 263.55, 263.95, 264.15, 
    265.05, 264.25, 263.85, 264.15, 263.35, 263.75, 261.75, 262.05, 260.95, 
    261.35, 262.05, 262.95, 263.05, 262.65, 261.85, 263.05, 262.65, 262.95, 
    263.55, 263.05, 262.65, 262.05, 262.25, 262.35, 262.35, 262.85, 262.75, 
    263.05, 263.55, 263.05, 263.45, 263.45, 263.65, 264.05, 264.25, 264.05, 
    264.55, 264.55, 264.75, 265.15, 264.75, 264.45, 264.75, 264.25, 264.35, 
    263.85, 263.55, 262.75, 262.55, 262.55, 262.35, 262.45, 262.35, 262.65, 
    262.55, 262.85, 263.05, 263.05, 263.05, 262.75, 262.55, 262.05, 261.85, 
    261.85, 261.85, 262.15, 262.05, 262.05, 262.15, 261.85, 261.85, 261.95, 
    262.05, 261.85, 261.45, 261.65, 261.85, 261.95, 262.15, 261.75, 262.15, 
    262.15, 261.85, 261.85, 261.75, 261.65, 261.85, 262.15, 261.25, 262.05, 
    261.45, 261.75, 261.45, 261.45, 261.35, 261.15, 261.55, 261.55, 261.85, 
    261.65, 261.75, 261.75, 261.85, 262.15, 262.15, 262.45, 262.85, 262.65, 
    263.05, 263.05, 263.35, 263.25, 263.45, 264.05, 264.05, 264.65, 264.75, 
    264.75, 264.55, 264.95, 265.65, 265.55, 265.45, 264.75, 265.65, 265.65, 
    264.25, 264.65, 264.45, 264.75, 265.15, 263.85, 265.15, 265.55, 266.35, 
    266.15, 266.75, 267.05, 266.65, 267.65, 266.75, 266.85, 266.75, 266.15, 
    266.45, 267.75, 267.75, 267.75, 267.75, 267.75, 267.75, 267.75, 267.75, 
    267.95, 267.75, 268.15, 268.05, 268.35, 267.75, 268.25, 268.15, 268.15, 
    268.25, 268.65, 268.65, 268.55, 268.45, 268.55, 268.85, 269.15, 268.95, 
    269.25, 269.45, 269.65, 269.65, 269.65, 269.35, 269.55, 269.65, 269.75, 
    269.55, 269.35, 269.65, 269.35, 269.45, 269.35, 269.35, 269.25, 269.55, 
    270.15, 270.25, 270.05, 268.75, 268.75, 268.85, 268.85, 268.85, 267.95, 
    265.05, 264.55, 265.35, 266.05, 266.65, 265.35, 266.25, 267.75, 267.95, 
    270.65, 271.35, 271.25, 271.15, 271.25, 270.95, 271.05, 271.45, 271.25, 
    270.95, 271.05, 270.85, 270.95, 270.45, 270.85, 270.55, 269.45, 268.65, 
    270.15, 269.35, 269.95, 269.15, 268.45, 267.95, 267.85, 268.05, 267.85, 
    268.05, 267.45, 267.75, 267.45, 266.75, 266.65, 266.85, 266.85, 266.45, 
    266.05, 265.85, 265.15, 265.55, 265.65, 265.75, 265.65, 265.25, 265.25, 
    265.25, 265.55, 265.25, 265.35, 265.25, 265.05, 264.45, 264.05, 264.15, 
    264.05, 263.85, 263.55, 263.15, 263.25, 263.05, 262.25, 262.75, 262.55, 
    262.45, 262.15, 261.05, 260.95, 261.25, 261.75, 261.45, 260.85, 261.05, 
    261.75, 261.95, 261.75, 260.95, 261.25, 261.15, 261.05, 261.55, 261.95, 
    261.95, 261.65, 261.45, 260.75, 260.75, 260.75, 260.95, 260.25, 260.05, 
    259.55, 259.55, 259.85, 259.85, 260.05, 260.75, 260.55, 261.15, 261.55, 
    261.75, 261.45, 261.55, 261.75, 262.15, 262.35, 262.85, 263.35, 263.65, 
    263.95, 264.65, 264.75, 265.05, 265.65, 266.05, 265.45, 264.85, 264.85, 
    264.55, 264.45, 264.45, 263.95, 264.15, 263.95, 264.05, 263.95, 264.05, 
    264.15, 264.05, 264.05, 264.35, 264.45, 264.05, 264.25, 264.45, 264.05, 
    264.25, 263.85, 263.65, 263.55, 263.55, 263.55, 262.75, 262.65, 263.65, 
    263.65, 263.55, 263.65, 263.65, 261.75, 262.75, 263.25, 263.45, 263.85, 
    263.75, 263.85, 263.85, 263.95, 263.25, 263.05, 262.65, 262.35, 263.05, 
    264.05, 263.05, 262.45, 263.85, 262.45, 263.85, 264.95, 263.15, 263.75, 
    264.05, 264.25, 263.65, 263.35, 263.55, 264.75, 264.55, 265.35, 264.95, 
    265.25, 265.85, 264.35, 266.55, 268.35, 268.25, 267.75, 267.45, 267.65, 
    267.35, 267.05, 266.85, 266.75, 266.65, 266.35, 266.55, 266.55, 266.25, 
    266.15, 266.15, 265.95, 265.95, 265.95, 264.55, 264.75, 263.75, 265.35, 
    264.35, 264.15, 262.95, 264.15, 264.35, 265.75, 266.15, 266.25, 265.85, 
    265.45, 265.65, 265.85, 265.85, 266.25, 266.55, 266.75, 267.05, 267.35, 
    267.15, 267.65, 268.05, 268.25, 268.15, 268.35, 268.75, 268.55, 268.15, 
    267.75, 268.15, 268.25, 268.65, 268.75, 268.85, 268.85, 268.95, 268.95, 
    269.55, 269.85, 270.25, 270.45, 270.55, 270.65, 269.65, 269.85, 269.65, 
    269.45, 269.25, 268.85, 269.15, 269.25, 269.05, 268.95, 268.75, 268.95, 
    269.25, 269.75, 270.15, 271.05, 271.05, 271.15, 271.55, 271.55, 271.55, 
    270.95, 271.05, 271.45, 271.65, 271.95, 272.15, 272.05, 272.05, 272.05, 
    272.05, 271.65, 271.55, 271.75, 271.75, 271.95, 271.45, 271.75, 271.45, 
    271.65, 271.65, 271.25, 271.05, 271.25, 270.35, 269.15, 268.15, 267.65, 
    267.05, 264.85, 262.25, 261.25, 260.45, 260.15, 259.25, 259.15, 259.05, 
    259.55, 259.25, 260.45, 261.35, 261.05, 260.75, 260.95, 260.85, 260.85, 
    261.05, 260.95, 260.45, 260.25, 260.25, 260.15, 259.85, 260.15, 259.95, 
    259.85, 260.15, 260.25, 260.25, 260.55, 261.15, 261.35, 261.05, 261.55, 
    261.55, 261.45, 262.65, 262.45, 263.65, 263.05, 263.15, 262.75, 261.85, 
    261.65, 261.25, 261.35, 260.85, 260.75, 261.75, 262.15, 262.55, 263.65, 
    264.05, 264.25, 263.85, 264.45, 264.45, 264.95, 264.25, 263.15, 262.95, 
    261.15, 260.45, 260.45, 260.85, 261.05, 261.75, 261.45, 260.75, 260.55, 
    260.55, 261.15, 261.25, 261.35, 261.65, 261.65, 262.25, 262.85, 264.25, 
    266.45, 268.25, 268.15, 268.05, 267.65, 267.95, 266.95, 266.95, 266.85, 
    266.55, 266.25, 266.45, 266.55, 266.25, 267.95, 265.75, 264.95, 264.65, 
    264.05, 263.45, 264.35, 265.25, 266.35, 265.45, 265.55, 265.45, 266.05, 
    265.85, 265.95, 265.75, 264.95, 263.95, 263.65, 264.25, 264.45, 262.15, 
    262.95, 262.65, 262.65, 262.85, 262.65, 262.85, 263.25, 263.95, 265.35, 
    265.65, 265.65, 265.95, 266.35, 266.35, 266.55, 266.65, 266.45, 266.35, 
    266.55, 267.35, 267.25, 267.15, 267.45, 266.85, 267.15, 267.35, 266.85, 
    267.45, 268.05, 268.15, 268.25, 268.75, 269.25, 269.35, 269.75, 269.85, 
    270.15, 270.35, 270.55, 270.15, 270.35, 270.75, 271.05, 271.15, 271.35, 
    271.55, 271.65, 271.55, 271.65, 268.55, 267.65, 265.95, 265.05, 263.65, 
    263.45, 263.15, 264.15, 263.65, 262.65, 263.05, 263.55, 263.15, 263.05, 
    262.65, 262.35, 262.25, 261.95, 261.45, 261.45, 260.75, 261.05, 261.35, 
    261.85, 261.15, 260.95, 260.95, 260.45, 260.45, 260.05, 259.75, 260.05, 
    259.75, 259.45, 259.05, 259.15, 258.65, 258.85, 258.25, 258.45, 258.65, 
    258.65, 258.45, 258.45, 258.65, 258.85, 259.15, 259.15, 258.85, 258.45, 
    258.75, 258.65, 258.55, 258.95, 258.85, 258.85, 259.15, 258.75, 258.75, 
    258.95, 259.05, 259.05, 258.65, 258.85, 258.55, 258.05, 257.95, 258.15, 
    258.25, 258.55, 257.95, 257.65, 257.15, 257.35, 257.15, 257.85, 258.95, 
    259.95, 261.25, 261.65, 262.35, 262.45, 262.95, 262.45, 262.05, 261.85, 
    262.15, 261.95, 261.75, 262.05, 261.55, 261.05, 260.55, 260.15, 259.95, 
    258.85, 259.45, 258.15, 257.85, 257.85, 258.25, 257.55, 257.65, 257.45, 
    256.85, 257.05, 256.85, 257.55, 257.55, 257.55, 257.55, 257.75, 257.85, 
    257.85, 257.85, 257.75, 257.55, 257.35, 256.95, 256.85, 256.85, 256.55, 
    256.65, 256.85, 256.35, 255.95, 255.75, 255.65, 255.45, 255.55, 255.95, 
    256.25, 256.85, 257.15, 257.45, 257.95, 258.65, 259.05, 259.25, 259.95, 
    259.15, 257.95, 257.65, 257.65, 256.85, 257.65, 258.15, 258.55, 260.55, 
    260.65, 261.15, 261.85, 261.45, 260.15, 260.45, 260.35, 261.15, 262.35, 
    261.85, 261.85, 261.95, 261.65, 262.15, 261.85, 261.75, 261.15, 261.05, 
    261.15, 261.05, 261.25, 261.95, 261.55, 261.15, 261.15, 261.25, 261.25, 
    261.15, 260.85, 260.45, 260.55, 261.15, 260.75, 260.65, 261.15, 260.95, 
    261.05, 261.65, 260.95, 260.75, 261.05, 260.95, 261.15, 261.15, 260.95, 
    260.85, 261.35, 262.05, 262.25, 262.45, 262.45, 264.25, 264.45, 264.55, 
    264.45, 264.65, 264.75, 264.95, 265.45, 265.55, 265.75, 265.95, 266.25, 
    266.85, 267.55, 267.55, 267.85, 268.45, 268.55, 268.45, 268.15, 268.55, 
    267.95, 268.15, 268.45, 268.75, 269.25, 269.65, 269.75, 269.55, 269.65, 
    269.85, 270.25, 270.15, 270.25, 270.35, 270.35, 270.45, 270.25, 270.35, 
    270.45, 270.05, 270.25, 270.45, 270.65, 270.85, 270.85, 270.95, 271.15, 
    271.25, 271.35, 271.45, 271.55, 271.45, 271.45, 271.55, 271.45, 271.05, 
    271.25, 269.85, 269.05, 269.15, 269.45, 269.15, 268.75, 268.35, 269.15, 
    269.35, 269.05, 268.65, 268.95, 269.05, 269.05, 269.55, 269.95, 270.35, 
    270.25, 270.75, 270.85, 270.75, 270.85, 270.85, 270.75, 270.85, 271.35, 
    271.25, 271.85, 271.85, 272.45, 272.55, 272.55, 272.55, 272.05, 273.45, 
    272.95, 272.55, 271.95, 271.55, 271.25, 271.45, 271.25, 272.05, 272.55, 
    271.55, 271.15, 271.05, 271.65, 273.55, 273.45, 273.15, 273.05, 271.95, 
    271.55, 272.05, 273.05, 273.25, 272.95, 273.45, 272.95, 273.45, 273.05, 
    273.15, 272.95, 272.75, 272.95, 272.85, 273.45, 273.75, 273.75, 273.25, 
    272.95, 273.15, 272.95, 272.95, 272.65, 272.75, 272.75, 272.55, 272.35, 
    271.55, 271.25, 270.65, 269.85, 269.25, 269.05, 269.15, 269.85, 269.05, 
    269.05, 268.45, 268.35, 268.35, 268.15, 268.35, 268.65, 268.75, 269.15, 
    269.85, 270.55, 271.55, 272.35, 273.45, 272.75, 272.25, 272.05, 272.45, 
    272.95, 272.65, 271.45, 272.35, 273.15, 274.05, 273.95, 274.25, 273.65, 
    274.75, 272.35, 271.85, 272.95, 272.85, 273.95, 273.15, 274.05, 274.35, 
    274.05, 274.95, 274.85, 273.95, 273.45, 273.25, 273.05, 272.95, 272.65, 
    272.45, 272.25, 272.15, 272.75, 271.95, 271.65, 271.75, 272.05, 271.65, 
    271.85, 270.85, 270.45, 271.15, 271.25, 270.25, 270.65, 271.35, 271.95, 
    271.95, 272.65, 272.75, 272.95, 273.05, 273.35, 273.55, 273.25, 273.25, 
    273.15, 272.55, 272.55, 271.65, 273.15, 272.15, 272.65, 272.35, 272.05, 
    271.85, 271.95, 271.55, 271.65, 272.45, 272.65, 271.75, 272.45, 272.15, 
    272.05, 271.95, 271.85, 271.65, 271.65, 271.35, 271.35, 271.15, 270.95, 
    270.45, 269.85, 269.45, 270.55, 269.75, 270.55, 269.35, 268.35, 267.85, 
    267.45, 269.05, 268.75, 267.55, 266.25, 265.35, 264.65, 263.75, 263.25, 
    262.65, 262.55, 262.45, 262.45, 262.05, 261.75, 261.85, 261.65, 261.55, 
    261.55, 261.45, 261.05, 260.45, 260.35, 259.85, 259.55, 259.95, 259.45, 
    258.95, 259.05, 259.05, 258.05, 258.55, 258.55, 258.15, 257.35, 257.75, 
    257.75, 258.15, 258.65, 258.75, 259.45, 260.15, 260.05, 260.15, 260.15, 
    260.55, 261.25, 261.25, 261.45, 261.15, 261.45, 262.05, 262.05, 261.45, 
    261.15, 261.25, 260.75, 260.45, 259.85, 259.85, 259.55, 259.15, 258.95, 
    258.75, 258.35, 258.15, 258.05, 257.35, 257.05, 256.95, 256.45, 256.45, 
    256.15, 255.65, 255.65, 254.75, 254.65, 254.55, 254.55, 254.35, 254.35, 
    254.35, 254.15, 253.85, 254.15, 253.75, 253.45, 252.95, 253.35, 253.45, 
    253.55, 253.95, 254.45, 254.45, 254.25, 254.45, 254.55, 254.75, 254.45, 
    254.55, 254.05, 254.05, 253.85, 253.45, 253.55, 252.95, 253.05, 253.05, 
    252.75, 253.35, 252.75, 252.45, 252.65, 253.45, 253.45, 253.35, 253.35, 
    253.25, 253.65, 253.85, 253.85, 253.55, 253.65, 253.35, 253.95, 253.95, 
    253.65, 253.65, 253.75, 253.55, 253.75, 253.95, 254.05, 253.85, 253.55, 
    253.95, 253.85, 254.05, 254.05, 253.95, 254.25, 254.25, 254.35, 254.65, 
    254.15, 253.35, 253.55, 253.85, 254.15, 254.95, 255.75, 255.35, 255.35, 
    255.75, 255.65, 256.65, 256.85, 258.65, 258.95, 258.85, 258.65, 258.85, 
    259.15, 259.05, 259.05, 258.85, 258.85, 258.65, 258.35, 258.35, 258.45, 
    258.75, 258.85, 258.45, 258.55, 259.35, 259.95, 260.95, 261.45, 262.15, 
    262.35, 263.05, 262.45, 261.85, 261.55, 261.75, 262.25, 262.95, 264.15, 
    264.75, 264.75, 264.85, 264.75, 264.45, 264.25, 264.45, 264.05, 262.45, 
    261.55, 260.55, 259.55, 259.15, 258.75, 258.45, 258.15, 257.85, 257.35, 
    257.35, 256.85, 256.55, 256.55, 256.75, 256.55, 256.45, 257.45, 257.15, 
    257.65, 257.45, 257.65, 257.85, 257.75, 258.25, 258.25, 258.55, 259.05, 
    258.75, 258.85, 259.15, 259.25, 259.25, 260.25, 260.45, 260.85, 260.85, 
    260.45, 258.35, 257.75, 257.35, 257.15, 257.25, 256.95, 256.95, 256.85, 
    257.35, 257.65, 256.85, 256.95, 256.95, 257.25, 258.65, 259.65, 261.05, 
    261.75, 261.15, 260.85, 260.45, 260.25, 260.55, 260.25, 260.15, 260.25, 
    260.55, 260.65, 260.65, 260.65, 260.65, 260.75, 260.85, 260.75, 261.45, 
    262.15, 262.75, 263.45, 263.75, 264.65, 265.45, 266.15, 266.35, 266.45, 
    266.55, 266.65, 266.65, 266.65, 266.55, 266.35, 265.95, 266.35, 266.25, 
    266.15, 266.35, 266.15, 266.15, 265.85, 265.85, 265.65, 265.55, 265.55, 
    265.75, 265.75, 265.35, 265.45, 265.65, 265.35, 264.95, 264.85, 264.65, 
    264.15, 263.55, 262.95, 262.55, 262.45, 261.95, 262.15, 262.15, 262.35, 
    262.15, 262.15, 262.05, 261.55, 261.95, 261.85, 261.55, 262.15, 262.25, 
    262.35, 263.05, 263.25, 262.85, 263.15, 263.85, 264.45, 264.95, 264.75, 
    264.75, 264.25, 264.25, 263.85, 263.65, 263.05, 263.35, 264.05, 264.45, 
    264.85, 265.05, 267.55, 267.25, 266.85, 266.25, 265.45, 264.85, 264.55, 
    264.35, 264.75, 264.95, 265.55, 265.45, 265.05, 264.55, 264.55, 264.95, 
    264.55, 264.05, 264.25, 263.75, 264.15, 264.15, 262.85, 261.95, 261.25, 
    261.95, 261.85, 261.55, 261.45, 261.75, 263.25, 263.15, 262.25, 262.85, 
    262.75, 263.35, 264.85, 264.75, 264.25, 262.95, 263.35, 263.45, 264.45, 
    265.25, 265.65, 265.45, 265.45, 265.85, 266.05, 266.25, 265.85, 265.65, 
    266.05, 266.35, 266.45, 266.25, 266.15, 266.15, 265.85, 266.05, 265.55, 
    266.15, 266.25, 266.25, 266.05, 265.95, 266.05, 265.95, 265.75, 265.85, 
    265.25, 264.45, 264.55, 265.55, 265.55, 265.35, 263.95, 264.35, 263.55, 
    263.85, 264.05, 264.55, 264.45, 265.05, 264.45, 264.15, 264.25, 264.25, 
    264.25, 263.75, 263.25, 262.55, 263.35, 262.45, 263.95, 263.95, 264.15, 
    264.15, 262.75, 260.45, 262.25, 262.25, 261.75, 261.75, 262.45, 263.05, 
    262.85, 262.75, 262.95, 263.05, 260.55, 262.45, 262.75, 262.25, 262.05, 
    262.15, 262.25, 262.45, 262.85, 262.25, 261.95, 261.95, 262.75, 262.05, 
    262.25, 262.45, 262.25, 261.95, 262.85, 262.45, 262.55, 263.05, 262.45, 
    262.35, 261.65, 261.65, 261.85, 261.25, 261.15, 260.65, 260.55, 260.55, 
    260.65, 261.05, 261.45, 261.55, 262.05, 262.65, 263.15, 263.85, 264.45, 
    264.95, 265.55, 266.55, 266.55, 263.75, 262.15, 260.15, 259.35, 258.25, 
    258.05, 256.95, 256.85, 256.65, 256.75, 256.65, 256.35, 256.55, 256.25, 
    256.45, 256.25, 256.15, 255.95, 256.15, 256.05, 256.05, 256.25, 256.35, 
    256.55, 256.65, 256.75, 256.85, 256.65, 256.65, 256.75, 256.65, 256.15, 
    256.55, 256.65, 256.65, 256.65, 257.05, 256.65, 256.85, 256.75, 256.75, 
    257.25, 256.85, 256.95, 256.95, 257.15, 257.35, 257.35, 256.45, 256.35, 
    256.85, 256.85, 256.55, 257.35, 258.35, 259.35, 259.25, 259.65, 260.05, 
    260.15, 260.25, 260.35, 260.65, 260.65, 260.45, 260.65, 260.85, 260.85, 
    260.85, 261.35, 261.85, 262.05, 261.65, 261.95, 261.65, 261.95, 262.45, 
    262.85, 260.85, 261.25, 261.25, 260.45, 259.65, 259.15, 258.45, 257.95, 
    257.55, 257.25, 256.75, 256.95, 256.85, 256.95, 257.25, 257.25, 257.25, 
    257.35, 257.05, 256.95, 256.75, 256.65, 256.55, 257.05, 256.95, 257.65, 
    258.45, 258.15, 257.85, 257.35, 257.05, 257.25, 257.05, 257.25, 256.85, 
    256.45, 255.95, 256.05, 256.25, 256.45, 256.65, 256.85, 257.15, 257.75, 
    258.05, 258.35, 258.85, 259.55, 261.65, 263.35, 265.05, 263.05, 260.85, 
    259.05, 257.65, 256.75, 255.55, 254.65, 253.85, 253.85, 253.75, 254.05, 
    255.35, 256.65, 259.05, 259.55, 259.35, 259.35, 258.75, 258.55, 257.95, 
    257.35, 256.65, 256.45, 256.45, 256.65, 256.85, 256.45, 255.65, 256.15, 
    256.95, 257.55, 259.55, 259.15, 258.45, 257.75, 257.45, 257.25, 257.05, 
    256.05, 255.95, 255.65, 254.85, 254.45, 253.65, 254.05, 254.05, 254.45, 
    254.15, 254.15, 254.45, 255.55, 257.05, 258.75, 261.15, 261.55, 262.05, 
    262.15, 262.55, 263.75, 264.65, 265.75, 266.25, 266.95, 267.15, 264.05, 
    261.85, 261.15, 260.75, 259.95, 259.65, 258.65, 256.85, 256.55, 256.45, 
    256.05, 255.85, 255.85, 256.75, 256.75, 258.65, 259.35, 261.15, 260.95, 
    261.15, 261.55, 262.15, 262.35, 263.85, 264.05, 265.35, 266.15, 266.45, 
    266.95, 268.05, 268.45, 268.95, 270.45, 270.95, 271.25, 271.15, 271.15, 
    271.55, 271.45, 271.05, 271.55, 271.15, 271.75, 271.95, 271.75, 272.05, 
    271.95, 268.85, 268.05, 267.35, 266.85, 266.55, 265.95, 265.45, 265.15, 
    264.95, 264.55, 264.35, 263.95, 263.65, 263.05, 262.45, 261.65, 261.15, 
    260.55, 260.45, 259.95, 259.85, 259.65, 259.55, 259.35, 259.15, 258.85, 
    258.65, 258.35, 258.45, 258.15, 258.25, 260.65, 258.15, 258.15, 258.05, 
    258.05, 258.35, 258.15, 258.05, 257.55, 257.35, 257.25, 257.25, 256.95, 
    256.95, 256.65, 255.95, 255.35, 255.05, 254.85, 254.35, 254.35, 253.55, 
    252.95, 252.55, 252.05, 251.65, 250.85, 250.35, 249.95, 249.65, 249.25, 
    249.25, 249.15, 249.25, 249.45, 249.75, 249.65, 250.05, 250.45, 250.15, 
    250.35, 250.65, 250.75, 250.65, 250.85, 250.85, 250.75, 250.65, 250.55, 
    250.55, 250.85, 250.95, 250.95, 250.85, 250.75, 250.55, 250.65, 250.85, 
    251.25, 251.35, 251.45, 251.75, 251.85, 251.85, 252.35, 252.65, 252.55, 
    252.35, 251.85, 251.55, 252.15, 252.05, 251.85, 251.85, 251.95, 251.85, 
    251.75, 251.55, 250.65, 251.55, 251.55, 251.45, 251.35, 251.15, 251.25, 
    251.15, 251.45, 251.35, 251.05, 250.95, 250.85, 250.65, 250.45, 250.45, 
    251.05, 251.25, 251.55, 251.65, 251.55, 252.05, 252.45, 252.25, 252.05, 
    251.95, 251.75, 251.35, 251.25, 251.25, 251.65, 252.05, 251.95, 252.25, 
    252.45, 252.35, 252.25, 251.95, 252.45, 252.05, 250.85, 251.35, 250.65, 
    250.85, 251.55, 250.65, 249.75, 251.35, 251.45, 254.65, 252.95, 253.25, 
    252.45, 253.25, 253.95, 253.65, 253.65, 255.15, 256.65, 257.95, 257.85, 
    257.95, 257.95, 256.75, 257.05, 257.95, 258.15, 258.65, 259.15, 259.35, 
    259.75, 260.15, 260.25, 260.45, 260.55, 260.95, 261.25, 261.45, 262.75, 
    263.25, 264.65, 266.05, 267.85, 269.15, 270.35, 269.85, 267.55, 265.75, 
    264.45, 263.95, 263.65, 261.75, 260.35, 259.15, 258.45, 257.75, 257.65, 
    256.65, 255.75, 255.55, 254.95, 255.15, 254.95, 255.85, 255.75, 255.45, 
    255.25, 255.55, 255.65, 256.05, 255.65, 255.35, 255.35, 254.85, 254.45, 
    253.95, 252.45, 251.15, 250.45, 249.75, 249.85, 250.35, 251.25, 251.75, 
    252.05, 252.55, 253.35, 253.75, 254.25, 253.85, 253.55, 253.35, 253.15, 
    253.25, 253.15, 252.55, 251.95, 251.65, 251.95, 251.55, 251.55, 251.05, 
    251.15, 252.15, 252.95, 252.35, 251.85, 251.05, 250.85, 250.85, 251.05, 
    251.15, 251.25, 251.15, 250.65, 250.65, 250.75, 250.85, 250.75, 249.65, 
    249.55, 249.55, 249.55, 249.15, 248.85, 248.25, 248.15, 247.75, 247.45, 
    247.45, 247.35, 247.05, 247.35, 247.75, 248.35, 249.15, 249.75, 250.45, 
    251.25, 251.75, 252.15, 252.55, 252.65, 252.15, 252.25, 251.95, 251.25, 
    251.25, 251.45, 251.15, 251.15, 250.25, 249.95, 249.55, 248.75, 248.25, 
    247.65, 247.55, 247.55, 247.55, 247.55, 247.65, 247.75, 247.65, 247.55, 
    247.85, 247.85, 248.05, 248.45, 248.75, 249.25, 249.45, 249.25, 248.95, 
    248.25, 247.55, 247.15, 246.95, 246.65, 246.85, 246.95, 247.35, 247.65, 
    248.15, 248.75, 249.45, 250.85, 250.65, 250.65, 250.15, 249.45, 248.55, 
    247.45, 246.85, 247.15, 247.45, 247.75, 247.65, 247.45, 247.45, 247.05, 
    247.95, 248.25, 248.35, 249.25, 250.35, 249.85, 249.45, 249.45, 249.75, 
    250.15, 251.75, 252.15, 252.45, 252.55, 252.15, 252.35, 252.25, 251.95, 
    252.25, 252.85, 252.95, 252.95, 252.55, 252.45, 252.25, 251.85, 251.55, 
    251.25, 251.15, 250.95, 250.85, 250.85, 250.65, 250.45, 250.65, 250.65, 
    250.75, 250.45, 250.35, 249.85, 249.85, 249.85, 249.55, 249.15, 249.05, 
    248.75, 247.75, 248.45, 248.35, 247.65, 247.55, 248.05, 248.25, 248.15, 
    248.35, 248.15, 248.85, 248.95, 249.15, 249.35, 249.25, 249.35, 249.25, 
    249.25, 248.45, 248.35, 249.55, 249.05, 249.55, 249.35, 249.95, 251.35, 
    251.35, 251.25, 251.65, 251.95, 252.35, 252.65, 252.75, 253.95, 254.25, 
    254.35, 254.35, 254.65, 254.25, 253.25, 253.75, 253.35, 253.05, 252.85, 
    253.35, 252.05, 252.85, 254.35, 253.45, 255.25, 255.75, 255.75, 255.45, 
    254.25, 255.25, 254.05, 253.95, 253.75, 254.45, 254.35, 253.55, 254.65, 
    253.25, 254.05, 255.45, 253.25, 252.95, 251.65, 250.35, 250.15, 251.05, 
    249.75, 250.45, 250.75, 250.65, 250.65, 250.65, 250.25, 250.05, 250.35, 
    250.65, 251.15, 251.75, 252.05, 252.45, 253.75, 254.35, 253.85, 254.25, 
    259.25, 259.95, 260.35, 259.75, 259.35, 259.25, 259.45, 259.45, 258.75, 
    259.65, 259.65, 259.75, 260.15, 260.35, 259.95, 258.85, 257.55, 256.65, 
    256.35, 258.95, 260.85, 262.05, 262.05, 263.15, 262.45, 261.55, 261.15, 
    261.55, 260.45, 259.65, 259.55, 260.75, 259.85, 260.25, 260.35, 260.65, 
    260.55, 260.15, 260.25, 260.35, 260.45, 260.45, 260.35, 260.65, 260.95, 
    261.15, 260.85, 261.05, 260.75, 260.25, 260.35, 261.25, 260.15, 259.85, 
    260.05, 259.95, 259.85, 260.25, 259.15, 258.55, 258.15, 257.65, 257.65, 
    257.85, 257.25, 257.75, 258.15, 258.35, 257.85, 257.55, 257.85, 257.45, 
    257.75, 258.35, 258.95, 259.25, 259.35, 259.25, 259.55, 258.75, 261.25, 
    258.85, 260.95, 262.25, 261.75, 263.65, 264.65, 264.95, 265.35, 265.65, 
    265.95, 266.25, 265.75, 265.65, 265.45, 265.55, 265.65, 265.65, 265.55, 
    265.15, 264.55, 264.85, 265.45, 265.95, 265.85, 265.45, 265.65, 265.25, 
    265.75, 266.05, 265.55, 265.85, 266.15, 266.35, 266.65, 266.55, 266.15, 
    265.35, 265.25, 265.65, 266.05, 265.45, 264.95, 264.45, 264.05, 263.75, 
    263.65, 263.25, 263.15, 262.55, 263.35, 263.15, 264.05, 263.15, 264.45, 
    264.75, 264.15, 264.15, 264.45, 264.35, 264.35, 263.45, 262.25, 263.75, 
    261.55, 260.75, 260.15, 260.85, 260.35, 260.35, 259.85, 259.85, 259.15, 
    259.05, 261.65, 262.05, 262.15, 259.95, 261.55, 262.55, 261.45, 263.25, 
    264.95, 263.85, 263.45, 264.15, 264.55, 264.55, 264.95, 265.05, 264.65, 
    263.85, 263.85, 264.55, 264.15, 263.35, 262.25, 261.35, 260.45, 258.85, 
    261.55, 260.35, 260.75, 261.95, 264.65, 263.75, 264.15, 262.35, 262.25, 
    263.15, 263.85, 262.85, 263.95, 262.15, 262.85, 262.25, 260.35, 259.05, 
    258.45, 257.05, 256.45, 256.35, 256.35, 256.45, 257.55, 258.45, 259.05, 
    259.35, 259.55, 259.95, 260.35, 260.75, 262.15, 260.85, 261.05, 262.45, 
    263.05, 263.95, 264.35, 264.45, 263.35, 259.55, 257.05, 255.55, 254.15, 
    253.15, 252.05, 251.75, 250.85, 251.05, 252.15, 250.75, 249.75, 251.05, 
    250.75, 251.15, 251.15, 251.35, 252.05, 252.25, 252.95, 252.65, 252.25, 
    251.75, 251.75, 251.15, 252.45, 253.35, 253.95, 254.05, 254.35, 253.85, 
    253.35, 252.85, 252.85, 253.65, 254.05, 254.25, 254.65, 254.75, 255.05, 
    255.45, 255.75, 256.05, 256.05, 256.25, 256.25, 256.25, 255.95, 256.65, 
    256.75, 256.85, 257.25, 256.85, 257.25, 257.45, 257.55, 257.55, 257.55, 
    257.65, 257.55, 257.85, 257.85, 257.85, 257.95, 257.95, 258.05, 257.65, 
    257.55, 257.45, 257.25, 257.05, 257.45, 257.15, 257.45, 256.95, 256.85, 
    257.65, 258.25, 258.35, 257.45, 258.65, 258.45, 259.85, 260.05, 260.25, 
    260.55, 260.55, 261.05, 261.35, 263.65, 263.65, 263.25, 262.75, 262.25, 
    261.85, 261.95, 262.45, 262.05, 261.75, 261.65, 261.75, 262.55, 261.85, 
    261.95, 262.55, 262.35, 262.35, 261.95, 262.55, 262.85, 262.35, 263.15, 
    263.25, 262.95, 263.25, 262.75, 262.45, 262.15, 261.75, 261.15, 261.55, 
    261.15, 261.15, 262.15, 262.35, 262.05, 261.95, 262.25, 262.45, 263.05, 
    263.95, 263.25, 263.55, 263.85, 263.15, 263.75, 263.55, 263.35, 264.65, 
    265.35, 265.75, 265.65, 265.85, 265.65, 265.55, 264.95, 264.75, 264.55, 
    264.45, 264.05, 264.15, 264.25, 264.05, 264.05, 264.55, 264.85, 265.45, 
    265.65, 264.85, 264.65, 264.75, 264.95, 264.95, 265.75, 266.05, 266.05, 
    265.75, 266.65, 267.05, 266.35, 266.15, 265.55, 265.25, 264.65, 264.65, 
    263.15, 263.85, 262.25, 263.95, 264.65, 265.05, 265.75, 265.95, 265.85, 
    265.95, 266.35, 265.95, 265.05, 263.75, 261.85, 260.35, 260.55, 260.55, 
    261.15, 261.65, 260.65, 261.35, 260.25, 260.25, 259.45, 259.95, 259.95, 
    260.75, 260.25, 260.05, 260.05, 260.15, 260.35, 260.05, 259.75, 258.75, 
    258.15, 258.45, 259.25, 259.05, 259.45, 259.85, 259.85, 260.15, 260.25, 
    260.35, 260.55, 260.45, 260.35, 260.45, 260.35, 260.25, 260.05, 259.85, 
    260.45, 261.15, 260.05, 260.65, 261.45, 260.35, 261.05, 261.15, 261.55, 
    261.05, 260.75, 260.45, 260.25, 260.45, 260.65, 260.75, 260.55, 260.45, 
    260.55, 261.35, 261.15, 260.55, 260.25, 260.25, 260.25, 260.35, 260.35, 
    260.15, 260.15, 259.85, 259.75, 259.95, 259.55, 259.45, 258.85, 259.05, 
    259.15, 258.95, 258.65, 258.45, 258.55, 258.65, 258.55, 258.65, 258.55, 
    258.65, 258.55, 258.45, 258.85, 259.05, 259.45, 259.35, 260.05, 259.65, 
    259.55, 259.75, 259.25, 258.55, 258.15, 258.45, 258.15, 257.95, 257.85, 
    258.05, 258.25, 257.75, 257.25, 257.45, 258.15, 259.25, 259.85, 260.15, 
    260.35, 260.45, 260.55, 260.65, 260.45, 260.35, 260.05, 259.85, 260.05, 
    260.25, 260.45, 260.55, 260.95, 261.05, 261.15, 261.65, 262.35, 262.95, 
    263.45, 260.95, 257.25, 256.25, 256.55, 257.15, 257.75, 257.45, 257.35, 
    257.35, 257.35, 257.05, 256.45, 255.85, 255.25, 254.95, 255.05, 255.05, 
    256.25, 256.55, 257.25, 257.75, 257.85, 259.25, 259.95, 260.75, 261.15, 
    261.75, 262.25, 263.35, 264.35, 265.35, 266.55, 267.35, 268.05, 268.65, 
    268.15, 268.65, 268.45, 267.95, 267.85, 267.85, 267.75, 268.05, 268.45, 
    269.05, 266.25, 265.35, 263.65, 262.15, 261.25, 260.95, 260.15, 259.35, 
    258.95, 258.35, 257.85, 257.65, 257.05, 256.65, 256.35, 256.15, 256.25, 
    256.15, 255.95, 255.85, 257.05, 258.05, 258.65, 258.95, 259.05, 258.65, 
    258.45, 258.65, 258.95, 259.35, 259.55, 259.75, 259.85, 260.15, 260.25, 
    259.85, 259.75, 259.85, 260.15, 260.85, 261.25, 261.65, 262.05, 262.25, 
    262.45, 262.35, 262.45, 261.95, 261.75, 261.85, 262.15, 262.55, 263.05, 
    263.05, 263.05, 263.25, 263.25, 263.35, 263.25, 262.75, 262.35, 262.05, 
    261.85, 261.65, 261.75, 262.25, 262.85, 262.85, 262.95, 263.35, 262.85, 
    262.05, 261.05, 259.95, 260.05, 259.65, 259.85, 260.15, 260.35, 260.55, 
    260.55, 260.65, 260.25, 260.25, 260.15, 259.75, 259.55, 259.25, 258.75, 
    258.15, 257.95, 257.65, 257.55, 257.45, 257.55, 257.65, 257.65, 257.75, 
    257.95, 258.15, 258.65, 258.75, 260.35, 261.55, 260.65, 260.95, 261.55, 
    261.55, 262.65, 263.55, 264.35, 264.75, 265.15, 265.55, 265.75, 266.15, 
    266.15, 266.15, 266.35, 266.65, 266.95, 267.35, 267.95, 267.95, 268.15, 
    268.45, 268.35, 266.75, 265.75, 265.35, 263.85, 262.75, 261.95, 260.95, 
    260.85, 260.45, 260.55, 260.65, 260.75, 260.65, 260.05, 258.45, 258.05, 
    258.25, 258.35, 259.05, 259.45, 259.95, 259.95, 259.05, 258.75, 258.85, 
    259.15, 259.15, 259.25, 259.75, 259.85, 259.55, 259.25, 258.55, 258.65, 
    258.75, 258.65, 258.25, 258.15, 258.35, 258.35, 257.75, 258.25, 258.75, 
    259.25, 259.65, 259.85, 260.15, 261.15, 261.55, 261.65, 261.65, 261.15, 
    260.15, 260.65, 260.65, 261.15, 261.45, 261.55, 261.55, 261.55, 261.25, 
    261.15, 261.15, 260.75, 260.75, 260.65, 260.65, 260.55, 260.55, 260.95, 
    260.95, 261.05, 261.05, 261.05, 260.85, 260.85, 260.65, 260.65, 260.55, 
    260.45, 260.25, 260.25, 260.05, 259.65, 259.65, 259.55, 259.35, 259.45, 
    259.45, 259.05, 258.95, 258.85, 258.75, 258.55, 258.75, 258.65, 258.55, 
    258.35, 258.15, 258.25, 258.25, 258.35, 258.35, 258.35, 258.35, 258.25, 
    258.45, 258.85, 259.05, 259.05, 259.05, 259.15, 259.05, 259.75, 259.85, 
    259.85, 259.95, 259.65, 259.75, 259.65, 259.85, 259.45, 259.35, 258.35, 
    258.45, 258.65, 258.75, 258.85, 258.95, 259.05, 259.15, 259.35, 259.65, 
    259.85, 259.65, 259.85, 260.15, 259.75, 259.75, 259.95, 260.25, 260.75, 
    261.45, 260.85, 260.35, 260.15, 260.05, 259.75, 259.85, 259.65, 259.55, 
    259.05, 259.05, 259.45, 259.95, 258.75, 258.45, 258.95, 258.95, 258.05, 
    259.05, 258.15, 259.05, 258.85, 259.05, 259.45, 260.15, 261.25, 261.15, 
    261.15, 261.75, 261.45, 261.55, 261.35, 261.65, 261.15, 260.55, 260.65, 
    260.45, 260.25, 260.55, 260.75, 261.45, 261.25, 262.55, 262.45, 263.45, 
    262.25, 261.25, 262.05, 261.75, 262.55, 261.85, 261.45, 261.15, 261.25, 
    260.85, 260.85, 260.45, 260.25, 260.45, 260.65, 261.05, 260.95, 261.25, 
    261.25, 261.75, 262.05, 261.85, 262.05, 262.15, 262.45, 262.15, 262.25, 
    262.35, 262.35, 262.25, 262.05, 262.15, 262.75, 263.65, 263.35, 262.55, 
    262.35, 262.65, 261.95, 262.85, 262.75, 263.25, 263.35, 263.45, 263.75, 
    264.25, 264.75, 264.85, 265.55, 266.45, 266.45, 267.35, 268.25, 268.05, 
    268.65, 268.85, 269.35, 269.15, 268.45, 268.55, 268.35, 267.95, 267.85, 
    267.35, 267.15, 266.65, 266.45, 266.25, 266.55, 266.95, 267.85, 268.65, 
    268.55, 269.45, 269.75, 270.05, 270.65, 271.05, 270.95, 270.65, 269.05, 
    266.55, 264.45, 262.65, 261.15, 260.65, 260.35, 260.05, 260.05, 259.95, 
    259.95, 261.05, 261.35, 261.15, 260.95, 260.75, 260.95, 261.35, 261.65, 
    261.75, 261.75, 261.55, 261.65, 261.55, 261.75, 261.55, 261.45, 260.75, 
    260.55, 260.55, 260.75, 261.05, 261.55, 261.15, 262.15, 262.35, 262.75, 
    263.25, 263.35, 263.65, 262.95, 261.25, 260.85, 261.05, 260.75, 260.75, 
    260.85, 260.65, 260.75, 260.75, 260.75, 260.55, 260.35, 260.15, 260.25, 
    260.05, 259.75, 259.75, 259.05, 259.15, 259.15, 259.35, 259.45, 259.35, 
    259.65, 259.65, 259.95, 260.25, 260.45, 260.95, 261.25, 261.05, 261.25, 
    261.15, 261.05, 261.05, 260.35, 260.65, 260.75, 260.45, 260.05, 260.35, 
    260.35, 259.85, 259.65, 259.65, 259.75, 259.85, 260.05, 259.95, 260.25, 
    260.75, 260.85, 260.75, 260.95, 261.15, 261.25, 260.75, 261.15, 260.35, 
    260.75, 260.45, 259.15, 260.05, 258.95, 259.55, 259.85, 259.65, 259.95, 
    260.15, 260.15, 261.45, 260.85, 261.55, 262.35, 262.25, 262.25, 262.25, 
    262.05, 262.05, 262.45, 262.65, 262.75, 262.45, 262.75, 263.45, 263.55, 
    263.65, 264.55, 264.95, 265.25, 265.35, 265.25, 265.25, 265.65, 266.05, 
    266.35, 266.95, 267.35, 267.55, 268.05, 268.35, 269.35, 269.65, 270.05, 
    270.05, 270.05, 270.25, 270.35, 270.25, 270.55, 270.65, 270.65, 270.75, 
    271.05, 268.05, 266.95, 266.55, 266.35, 266.45, 266.15, 266.15, 265.85, 
    265.75, 265.75, 265.25, 264.85, 264.75, 264.35, 264.35, 264.55, 265.05, 
    265.45, 265.85, 266.05, 265.95, 265.85, 266.15, 264.55, 264.75, 264.95, 
    265.15, 265.25, 265.35, 265.95, 266.25, 266.55, 266.85, 266.65, 266.75, 
    266.75, 266.75, 266.85, 266.85, 266.85, 266.85, 267.25, 266.95, 267.35, 
    266.45, 267.25, 266.15, 265.75, 265.65, 265.75, 265.55, 265.55, 265.95, 
    265.95, 266.05, 266.45, 267.15, 267.55, 267.55, 267.65, 268.35, 268.55, 
    267.75, 267.05, 265.85, 265.45, 265.35, 264.55, 263.25, 263.45, 264.45, 
    264.05, 263.15, 262.25, 262.05, 262.15, 262.75, 263.15, 263.55, 264.25, 
    264.45, 263.75, 264.05, 264.05, 264.05, 264.35, 264.25, 264.25, 264.35, 
    264.15, 264.55, 263.95, 263.85, 263.75, 263.95, 264.05, 264.05, 264.15, 
    264.05, 263.95, 264.15, 265.05, 265.45, 265.65, 265.85, 265.85, 265.95, 
    265.95, 266.25, 265.95, 265.95, 265.85, 265.65, 265.85, 265.85, 266.05, 
    265.75, 265.15, 265.05, 264.45, 264.85, 265.15, 266.55, 267.05, 268.55, 
    266.55, 266.65, 267.25, 266.55, 267.55, 267.65, 267.75, 267.35, 267.25, 
    267.45, 267.15, 267.05, 266.75, 266.65, 266.45, 266.55, 266.55, 266.35, 
    266.45, 266.35, 266.45, 266.65, 266.85, 267.05, 266.85, 266.95, 267.15, 
    267.15, 266.95, 266.65, 266.15, 265.85, 265.55, 265.65, 265.55, 265.25, 
    265.05, 264.55, 264.75, 264.75, 264.35, 264.95, 266.25, 267.65, 268.45, 
    268.65, 268.85, 269.05, 269.55, 269.95, 270.45, 270.45, 269.95, 270.05, 
    269.85, 269.95, 270.05, 270.25, 270.25, 270.35, 270.75, 270.85, 270.95, 
    271.05, 271.05, 271.05, 271.05, 271.05, 271.25, 271.45, 271.45, 271.65, 
    272.55, 271.75, 272.25, 272.05, 272.35, 272.65, 272.75, 272.95, 272.95, 
    272.85, 272.85, 272.95, 273.15, 273.15, 273.15, 272.45, 271.85, 269.95, 
    269.65, 271.45, 270.55, 269.25, 269.65, 269.85, 269.75, 269.15, 269.85, 
    270.95, 270.95, 271.75, 271.95, 272.25, 271.25, 271.25, 271.35, 271.45, 
    271.25, 271.25, 271.25, 270.55, 269.75, 269.55, 269.95, 270.15, 270.15, 
    270.15, 270.35, 270.65, 271.05, 271.25, 272.15, 272.65, 272.65, 272.85, 
    273.35, 272.75, 272.35, 272.85, 271.55, 271.35, 271.35, 270.95, 270.55, 
    270.35, 270.05, 269.95, 269.45, 269.95, 269.25, 269.15, 268.75, 270.15, 
    268.85, 268.85, 269.05, 269.85, 270.15, 270.95, 270.95, 270.55, 270.05, 
    270.05, 270.05, 269.55, 269.65, 269.65, 269.45, 269.15, 269.15, 269.25, 
    268.65, 268.55, 268.15, 268.35, 268.25, 268.15, 268.25, 267.95, 267.85, 
    268.45, 268.65, 268.65, 268.75, 268.65, 268.75, 268.95, 268.75, 268.55, 
    268.75, 268.75, 268.35, 268.25, 267.65, 267.55, 267.65, 267.85, 267.65, 
    267.75, 267.95, 268.35, 269.05, 269.65, 269.95, 270.05, 269.55, 269.35, 
    269.55, 268.75, 269.05, 269.65, 268.95, 268.85, 268.75, 268.15, 267.75, 
    267.25, 266.85, 266.85, 267.05, 267.25, 267.15, 267.15, 266.55, 266.55, 
    266.75, 267.05, 267.85, 268.95, 269.95, 269.15, 269.35, 269.45, 270.05, 
    269.45, 269.85, 268.85, 269.15, 268.95, 268.45, 268.15, 269.95, 271.55, 
    269.95, 271.15, 270.45, 271.05, 271.25, 271.65, 272.05, 271.35, 271.45, 
    271.45, 271.85, 271.65, 271.85, 272.05, 271.95, 271.45, 271.25, 271.15, 
    271.15, 271.25, 271.15, 271.05, 271.25, 271.55, 271.65, 271.65, 271.75, 
    272.45, 272.25, 272.15, 272.55, 272.65, 272.85, 273.15, 272.55, 272.65, 
    272.85, 272.55, 272.75, 272.95, 273.25, 272.45, 272.45, 272.35, 272.35, 
    272.35, 272.45, 272.45, 272.45, 272.45, 272.65, 272.55, 271.95, 272.55, 
    271.75, 271.95, 271.25, 270.65, 270.15, 269.45, 269.75, 270.05, 270.35, 
    270.05, 269.85, 269.75, 269.35, 269.35, 269.25, 269.05, 268.85, 268.35, 
    268.15, 267.45, 267.15, 266.75, 266.65, 267.05, 267.15, 266.95, 267.25, 
    267.55, 268.05, 268.75, 268.55, 269.05, 269.35, 269.15, 269.55, 269.25, 
    269.75, 269.45, 269.75, 271.05, 271.25, 271.15, 271.55, 271.65, 271.85, 
    271.95, 271.95, 272.15, 272.25, 272.15, 271.75, 271.65, 271.75, 271.55, 
    271.35, 271.25, 271.25, 271.35, 270.95, 271.15, 271.15, 271.35, 270.95, 
    271.45, 272.55, 273.15, 274.65, 275.15, 274.85, 273.85, 273.35, 272.75, 
    272.45, 272.75, 272.55, 272.75, 272.85, 272.85, 273.05, 272.95, 272.95, 
    273.05, 272.75, 272.55, 272.55, 272.25, 272.25, 272.35, 272.55, 272.35, 
    272.45, 272.25, 272.35, 272.35, 272.45, 272.55, 272.45, 272.45, 272.85, 
    273.15, 272.75, 272.85, 272.75, 272.55, 271.85, 271.75, 271.15, 270.15, 
    269.55, 269.45, 269.35, 269.25, 269.35, 269.45, 269.45, 269.45, 269.35, 
    269.55, 269.55, 269.45, 269.15, 269.25, 269.35, 269.25, 269.55, 269.65, 
    269.85, 269.75, 269.65, 269.85, 270.15, 270.45, 270.45, 270.55, 270.55, 
    270.45, 270.45, 270.35, 270.55, 270.85, 270.95, 271.15, 271.45, 271.95, 
    272.45, 272.45, 272.35, 272.45, 272.65, 273.15, 273.75, 273.75, 273.05, 
    274.15, 272.05, 271.85, 271.55, 272.05, 272.55, 272.35, 272.15, 271.95, 
    271.75, 271.75, 271.45, 271.55, 271.25, 271.25, 271.45, 271.55, 271.75, 
    271.65, 271.85, 271.95, 271.65, 271.65, 271.45, 271.45, 271.45, 271.45, 
    271.25, 271.25, 271.05, 270.75, 270.75, 270.75, 270.75, 270.55, 270.55, 
    270.55, 270.55, 270.55, 270.55, 271.15, 271.05, 270.95, 271.15, 270.95, 
    270.95, 270.95, 271.05, 270.95, 270.85, 270.75, 270.65, 270.75, 270.75, 
    270.95, 270.75, 270.55, 270.45, 270.55, 270.85, 270.75, 271.05, 271.25, 
    271.35, 271.55, 271.65, 272.35, 272.35, 271.95, 272.35, 272.55, 272.65, 
    272.65, 272.35, 272.25, 272.15, 272.25, 271.95, 271.55, 271.05, 270.85, 
    270.35, 270.35, 270.05, 270.65, 270.75, 270.65, 270.95, 270.75, 271.35, 
    270.95, 271.15, 271.35, 271.55, 271.85, 271.85, 271.65, 271.95, 272.45, 
    272.45, 272.45, 272.55, 272.45, 272.55, 272.35, 272.25, 272.25, 272.35, 
    272.15, 272.55, 272.85, 272.95, 273.15, 273.45, 273.75, 274.05, 274.25, 
    274.75, 275.15, 275.15, 275.15, 274.85, 274.05, 273.25, 272.85, 273.15, 
    272.75, 272.65, 272.25, 272.05, 272.25, 272.35, 272.55, 272.65, 272.85, 
    273.05, 273.25, 273.25, 273.35, 273.55, 273.45, 273.45, 273.45, 273.55, 
    273.25, 273.15, 273.05, 272.95, 272.65, 272.45, 272.65, 272.05, 272.35, 
    272.15, 271.65, 272.05, 272.25, 272.25, 272.15, 272.45, 272.65, 272.25, 
    272.55, 273.05, 272.65, 272.95, 272.75, 272.55, 272.65, 272.65, 272.55, 
    272.55, 272.65, 272.55, 272.65, 272.65, 272.65, 272.65, 272.95, 273.15, 
    273.05, 273.15, 273.35, 273.45, 273.35, 273.45, 273.65, 273.45, 273.15, 
    273.05, 273.15, 273.15, 273.15, 273.15, 273.05, 272.95, 272.85, 272.95, 
    273.05, 272.75, 272.65, 272.45, 272.75, 272.65, 272.75, 272.65, 272.55, 
    272.95, 272.95, 273.15, 273.45, 273.85, 273.65, 273.85, 273.55, 273.25, 
    273.05, 273.15, 273.15, 273.35, 273.15, 273.05, 272.85, 272.85, 272.75, 
    272.85, 272.75, 272.65, 272.65, 272.75, 272.85, 273.25, 273.55, 273.45, 
    273.45, 273.15, 273.25, 273.65, 273.15, 273.95, 273.45, 273.25, 273.25, 
    273.15, 273.15, 273.15, 273.25, 272.65, 272.45, 272.45, 272.45, 272.45, 
    272.45, 272.55, 272.65, 272.65, 272.85, 272.35, 272.35, 272.15, 272.35, 
    273.35, 274.05, 274.15, 274.55, 273.75, 272.75, 272.75, 272.55, 272.55, 
    272.45, 272.85, 272.75, 273.05, 273.25, 273.85, 274.05, 273.85, 273.95, 
    273.95, 273.95, 274.05, 273.95, 274.35, 274.75, 274.05, 274.35, 274.05, 
    273.85, 273.85, 273.85, 273.55, 273.25, 273.15, 272.95, 272.85, 272.65, 
    272.45, 272.45, 272.15, 272.35, 272.75, 272.75, 272.95, 273.05, 273.35, 
    273.45, 273.45, 273.25, 273.35, 273.05, 273.05, 273.35, 273.55, 273.65, 
    273.85, 273.85, 274.05, 273.95, 274.05, 273.95, 273.75, 273.55, 273.45, 
    273.45, 273.35, 273.65, 273.45, 273.95, 273.65, 273.55, 273.75, 273.65, 
    273.55, 273.45, 273.75, 273.75, 273.85, 273.95, 273.75, 273.25, 273.35, 
    273.45, 273.45, 273.55, 273.65, 273.65, 273.65, 273.65, 273.75, 273.95, 
    274.15, 274.25, 274.45, 273.95, 273.85, 273.75, 273.85, 273.65, 273.55, 
    273.65, 273.45, 273.35, 272.95, 272.35, 272.85, 272.85, 272.85, 272.75, 
    272.45, 272.45, 272.45, 272.35, 272.35, 272.15, 272.15, 272.15, 271.95, 
    271.95, 271.85, 271.85, 271.85, 271.95, 272.15, 271.25, 272.35, 272.25, 
    272.35, 272.65, 272.85, 272.75, 272.55, 272.35, 272.25, 272.15, 272.35, 
    272.45, 272.25, 272.35, 272.25, 272.35, 272.25, 272.35, 272.55, 272.75, 
    272.95, 272.75, 272.65, 272.55, 272.45, 272.45, 272.55, 271.95, 271.25, 
    270.75, 270.35, 269.85, 269.15, 269.65, 269.45, 269.35, 269.75, 270.05, 
    269.95, 270.05, 270.45, 271.15, 271.75, 271.95, 271.85, 272.05, 271.25, 
    271.25, 270.65, 270.05, 269.75, 269.65, 269.45, 269.25, 269.25, 269.15, 
    269.05, 269.35, 270.45, 270.15, 269.75, 270.35, 270.55, 270.95, 271.75, 
    272.15, 272.55, 271.85, 272.65, 272.15, 271.65, 271.45, 271.95, 271.95, 
    272.45, 271.95, 272.25, 272.55, 272.05, 272.55, 272.25, 272.15, 272.25, 
    272.25, 272.35, 272.05, 272.05, 272.85, 273.95, 273.65, 272.65, 273.35, 
    273.45, 273.45, 273.45, 273.45, 273.35, 273.35, 273.55, 273.35, 273.15, 
    273.25, 273.25, 272.95, 272.85, 272.65, 272.65, 272.65, 272.65, 272.75, 
    272.85, 272.95, 273.05, 273.15, 273.15, 273.25, 273.55, 273.85, 272.35, 
    272.55, 272.75, 272.55, 273.05, 273.55, 273.85, 274.05, 274.75, 274.25, 
    274.85, 274.95, 275.05, 274.95, 274.35, 274.05, 274.05, 274.55, 273.35, 
    274.35, 274.35, 275.15, 276.35, 276.85, 276.75, 274.75, 275.15, 275.65, 
    276.45, 275.05, 276.05, 276.75, 275.35, 276.55, 276.65, 277.05, 275.45, 
    275.75, 277.25, 275.95, 276.55, 275.55, 274.25, 274.85, 274.55, 274.15, 
    274.35, 274.85, 275.45, 276.75, 277.45, 277.25, 277.35, 276.85, 276.15, 
    275.65, 275.45, 275.25, 274.95, 274.25, 274.25, 273.15, 273.15, 273.35, 
    273.55, 273.35, 273.25, 273.25, 273.35, 273.35, 273.35, 273.35, 273.25, 
    273.15, 273.15, 273.45, 273.15, 273.25, 273.15, 272.85, 272.65, 272.75, 
    272.85, 272.85, 272.95, 272.95, 272.85, 272.85, 272.75, 272.95, 273.05, 
    273.25, 273.75, 273.65, 273.25, 273.65, 273.55, 273.45, 273.05, 272.85, 
    272.35, 272.45, 271.85, 271.95, 272.15, 271.95, 271.75, 272.85, 273.45, 
    274.05, 273.95, 274.55, 274.95, 275.25, 275.65, 275.65, 275.45, 275.85, 
    274.95, 274.95, 274.95, 274.55, 274.75, 274.75, 274.95, 275.45, 275.55, 
    275.75, 276.95, 276.95, 275.45, 275.35, 274.95, 275.15, 276.15, 276.55, 
    276.15, 276.15, 275.65, 275.85, 275.75, 275.35, 275.15, 275.15, 274.45, 
    272.75, 272.25, 272.65, 273.85, 273.85, 273.85, 273.45, 272.85, 272.25, 
    272.25, 273.95, 273.75, 274.25, 274.35, 274.85, 274.65, 274.45, 274.45, 
    274.55, 274.75, 274.85, 274.85, 274.95, 274.95, 274.75, 274.35, 274.05, 
    273.75, 273.35, 273.15, 272.85, 272.65, 272.25, 272.35, 271.75, 271.75, 
    271.65, 271.85, 272.15, 272.35, 272.75, 273.05, 273.75, 274.95, 273.95, 
    276.55, 275.75, 275.55, 275.15, 275.65, 274.35, 274.75, 275.65, 275.85, 
    275.85, 275.45, 275.65, 275.05, 274.85, 274.15, 273.65, 273.65, 274.25, 
    274.35, 274.45, 275.65, 275.35, 275.45, 274.95, 274.85, 274.55, 274.45, 
    275.85, 274.55, 275.05, 274.75, 274.95, 274.95, 274.75, 274.55, 274.65, 
    275.25, 275.75, 276.15, 276.45, 276.45, 276.05, 278.35, 276.55, 278.35, 
    280.25, 280.55, 277.05, 279.75, 277.95, 279.35, 279.45, 279.05, 277.85, 
    277.45, 277.95, 276.65, 277.85, 274.55, 273.65, 275.35, 275.25, 276.15, 
    276.15, 273.95, 273.85, 274.45, 276.25, 276.65, 277.15, 275.45, 276.25, 
    275.95, 274.95, 274.75, 275.65, 275.25, 275.15, 274.55, 274.95, 274.45, 
    273.55, 273.25, 273.85, 273.95, 274.35, 274.75, 274.95, 274.95, 275.05, 
    274.35, 274.95, 275.15, 275.25, 275.15, 276.85, 278.25, 279.05, 279.25, 
    278.25, 276.85, 275.65, 275.25, 274.75, 275.75, 276.25, 275.55, 275.65, 
    275.45, 275.55, 275.25, 275.25, 274.75, 275.05, 275.35, 275.85, 276.65, 
    275.15, 276.25, 275.85, 276.35, 278.75, 281.35, 275.85, 275.55, 274.15, 
    276.85, 276.65, 274.35, 274.05, 274.55, 274.75, 275.55, 274.45, 277.25, 
    278.25, 277.35, 277.35, 277.75, 276.55, 277.25, 277.05, 276.85, 276.95, 
    277.35, 278.15, 278.15, 277.55, 274.25, 274.95, 275.15, 274.75, 274.35, 
    274.25, 274.25, 274.05, 273.75, 273.45, 273.45, 273.95, 274.85, 275.55, 
    273.85, 274.35, 275.05, 275.95, 275.85, 275.65, 275.75, 275.75, 275.95, 
    276.45, 275.75, 275.25, 274.95, 274.65, 274.65, 274.95, 275.15, 274.95, 
    275.05, 275.15, 275.35, 275.35, 275.55, 275.45, 274.85, 274.85, 275.45, 
    274.95, 274.65, 276.65, 277.35, 277.35, 277.25, 277.25, 277.25, 277.25, 
    277.15, 275.95, 276.25, 275.85, 275.15, 274.85, 274.55, 274.85, 275.75, 
    275.85, 275.85, 275.25, 276.15, 275.95, 275.55, 275.45, 275.25, 274.85, 
    273.95, 273.75, 273.65, 276.25, 276.45, 275.35, 276.55, 277.55, 277.75, 
    277.55, 277.15, 277.35, 277.55, 277.25, 277.25, 276.95, 276.55, 276.35, 
    276.05, 276.35, 276.65, 276.95, 275.95, 274.55, 274.55, 274.85, 275.65, 
    276.75, 276.15, 276.15, 275.95, 275.75, 276.45, 276.45, 276.65, 277.05, 
    277.45, 275.05, 277.05, 276.45, 276.65, 276.15, 276.25, 275.65, 276.35, 
    276.15, 276.55, 277.35, 276.05, 276.95, 277.45, 278.05, 278.55, 279.05, 
    278.95, 277.05, 276.85, 276.75, 275.25, 274.25, 274.15, 273.35, 273.75, 
    273.55, 275.45, 274.75, 274.35, 272.95, 272.35, 272.55, 272.65, 273.65, 
    272.95, 272.15, 272.25, 272.25, 271.75, 271.45, 271.35, 271.45, 271.45, 
    271.25, 270.75, 270.55, 270.35, 269.85, 269.85, 269.75, 270.55, 271.05, 
    271.75, 272.65, 272.55, 273.25, 273.75, 276.55, 277.95, 274.25, 274.15, 
    274.85, 272.55, 272.15, 272.35, 272.25, 272.75, 271.75, 271.65, 271.65, 
    271.85, 271.85, 272.05, 271.95, 272.25, 272.25, 272.05, 272.65, 273.75, 
    274.95, 274.75, 273.65, 274.25, 274.05, 273.95, 273.25, 272.75, 273.15, 
    273.45, 273.45, 274.25, 274.55, 274.65, 274.15, 274.85, 274.05, 273.35, 
    274.05, 274.75, 273.15, 273.55, 274.65, 273.75, 273.75, 273.35, 273.25, 
    273.55, 273.15, 273.15, 273.35, 272.75, 272.75, 272.85, 272.95, 272.95, 
    272.95, 272.85, 272.65, 272.95, 272.85, 272.65, 272.45, 272.35, 272.15, 
    272.15, 272.05, 271.95, 271.65, 271.55, 271.65, 271.75, 272.25, 272.65, 
    272.45, 272.45, 272.05, 271.65, 271.25, 271.05, 270.75, 270.85, 270.75, 
    270.95, 271.15, 270.85, 270.45, 270.55, 270.75, 271.35, 271.75, 271.95, 
    272.15, 272.25, 272.05, 272.15, 272.15, 272.25, 272.35, 272.15, 272.25, 
    272.25, 272.35, 272.45, 272.45, 272.25, 272.25, 272.05, 271.85, 271.85, 
    271.95, 271.95, 272.05, 271.95, 271.95, 271.85, 271.95, 271.95, 272.05, 
    272.15, 272.25, 272.35, 272.55, 272.45, 272.45, 272.55, 272.35, 271.75, 
    271.55, 271.55, 271.85, 271.65, 271.65, 272.05, 272.05, 272.25, 273.05, 
    273.35, 274.35, 276.75, 275.15, 274.75, 274.85, 275.05, 275.25, 275.95, 
    275.15, 274.65, 274.35, 274.05, 275.35, 275.55, 275.15, 274.95, 274.65, 
    274.65, 274.95, 275.35, 274.75, 274.75, 274.35, 273.85, 273.35, 273.05, 
    272.95, 272.85, 272.95, 272.75, 272.55, 272.35, 272.15, 271.75, 271.55, 
    271.65, 271.55, 271.45, 271.15, 271.25, 270.65, 270.15, 271.05, 272.55, 
    272.35, 271.95, 273.15, 274.15, 275.45, 273.45, 274.85, 276.75, 275.45, 
    276.55, 275.85, 277.35, 276.95, 276.65, 275.85, 275.75, 275.05, 276.65, 
    275.45, 276.35, 276.65, 276.65, 275.75, 275.35, 275.75, 276.45, 276.75, 
    275.15, 275.05, 274.35, 273.25, 273.15, 274.05, 274.55, 274.25, 274.35, 
    274.25, 274.55, 274.35, 273.95, 273.55, 273.65, 273.25, 273.35, 273.35, 
    272.55, 271.95, 271.75, 271.45, 271.65, 271.65, 271.85, 272.65, 272.45, 
    272.95, 273.05, 273.45, 274.45, 276.25, 276.75, 275.75, 274.55, 274.25, 
    272.35, 271.85, 271.75, 271.95, 271.85, 271.45, 270.55, 270.25, 270.15, 
    270.55, 270.35, 270.65, 271.15, 271.05, 271.05, 271.65, 271.25, 271.65, 
    271.65, 272.15, 272.55, 272.55, 273.25, 273.45, 273.45, 273.75, 274.15, 
    274.55, 274.25, 274.25, 274.25, 274.15, 274.05, 274.05, 274.95, 275.05, 
    275.55, 275.65, 276.65, 276.65, 277.05, 276.95, 276.25, 276.65, 276.15, 
    276.45, 276.25, 275.55, 275.05, 276.15, 275.65, 275.05, 275.15, 275.15, 
    275.35, 275.55, 275.35, 275.35, 276.15, 275.55, 275.25, 275.35, 275.05, 
    274.75, 274.75, 274.45, 274.35, 274.65, 274.05, 274.35, 274.45, 274.35, 
    274.25, 274.35, 274.85, 273.85, 274.05, 274.25, 273.85, 274.35, 274.45, 
    274.55, 273.85, 274.55, 274.95, 275.85, 273.85, 275.75, 275.15, 275.85, 
    276.45, 276.35, 275.85, 275.75, 276.25, 275.65, 275.25, 276.15, 276.85, 
    274.55, 274.55, 274.25, 274.55, 275.05, 275.05, 275.05, 275.35, 275.35, 
    275.65, 275.45, 275.25, 275.25, 275.25, 275.15, 275.25, 275.05, 275.15, 
    274.95, 275.15, 275.15, 275.35, 275.25, 275.25, 275.35, 275.55, 275.05, 
    275.15, 274.55, 274.65, 274.95, 274.25, 274.05, 273.95, 274.05, 274.35, 
    274.25, 274.15, 274.15, 274.45, 274.15, 274.25, 274.15, 273.95, 273.55, 
    273.45, 273.35, 273.25, 273.95, 274.65, 274.25, 274.45, 275.05, 274.95, 
    274.95, 275.15, 275.25, 274.85, 274.75, 274.55, 274.55, 274.55, 274.75, 
    274.55, 274.55, 274.35, 274.05, 273.65, 273.75, 273.75, 273.65, 273.85, 
    273.75, 273.95, 273.95, 273.45, 273.25, 272.85, 272.75, 272.45, 272.65, 
    272.95, 273.05, 273.75, 273.75, 273.45, 273.35, 273.35, 273.05, 272.95, 
    272.85, 273.05, 273.15, 273.05, 273.15, 273.35, 273.25, 273.05, 272.75, 
    273.35, 273.75, 274.15, 274.05, 274.15, 274.15, 274.55, 274.35, 274.55, 
    274.15, 273.85, 273.55, 273.65, 273.55, 273.45, 273.25, 273.35, 273.45, 
    273.65, 273.85, 274.45, 272.25, 273.25, 272.45, 272.55, 272.85, 272.85, 
    272.45, 272.65, 272.35, 272.35, 272.05, 271.85, 271.95, 271.75, 271.45, 
    271.75, 271.55, 271.55, 271.75, 271.85, 271.95, 271.95, 272.05, 272.05, 
    272.05, 272.05, 271.95, 271.95, 271.75, 271.15, 271.15, 271.05, 271.05, 
    270.75, 270.35, 270.65, 270.65, 270.95, 271.15, 271.15, 270.95, 270.75, 
    271.35, 271.25, 271.15, 271.25, 271.55, 271.85, 272.15, 271.95, 271.85, 
    272.05, 272.25, 272.35, 272.45, 272.55, 272.45, 272.55, 272.65, 272.75, 
    272.95, 272.75, 272.85, 272.45, 272.55, 272.55, 272.45, 272.15, 272.15, 
    271.95, 271.95, 271.85, 271.75, 271.45, 271.45, 271.15, 271.05, 270.95, 
    271.05, 271.15, 271.15, 271.25, 271.25, 271.35, 271.45, 271.55, 271.65, 
    271.75, 271.85, 271.95, 272.15, 272.25, 272.45, 272.25, 272.25, 272.05, 
    271.85, 271.75, 271.55, 271.75, 271.75, 271.75, 271.85, 271.55, 271.65, 
    271.75, 271.85, 271.95, 271.95, 272.25, 272.45, 272.45, 272.85, 272.45, 
    272.45, 272.35, 272.35, 272.45, 272.55, 272.75, 272.45, 272.05, 271.55, 
    271.75, 271.65, 271.55, 271.35, 271.25, 270.85, 270.65, 270.45, 270.45, 
    270.95, 270.95, 270.95, 270.65, 270.85, 270.65, 270.65, 271.05, 271.15, 
    271.05, 271.35, 271.45, 271.55, 271.75, 271.95, 272.05, 272.25, 272.05, 
    271.65, 271.75, 271.95, 272.25, 272.55, 272.65, 272.85, 272.95, 273.35, 
    273.25, 273.35, 273.25, 273.35, 273.45, 273.45, 273.55, 273.05, 272.65, 
    272.45, 273.05, 272.25, 271.95, 271.65, 271.85, 271.95, 271.75, 271.65, 
    271.55, 271.55, 271.65, 271.25, 270.05, 269.75, 269.75, 269.45, 269.55, 
    269.45, 269.35, 269.15, 269.55, 269.75, 270.05, 269.55, 269.45, 269.15, 
    269.05, 268.85, 268.75, 268.85, 268.85, 269.15, 268.85, 269.65, 270.15, 
    271.95, 272.75, 273.25, 273.45, 273.15, 272.65, 272.25, 272.45, 272.85, 
    273.25, 272.75, 273.15, 273.65, 273.85, 273.35, 273.85, 274.15, 273.75, 
    273.35, 273.15, 273.15, 272.35, 272.25, 272.25, 273.25, 273.85, 273.15, 
    275.75, 275.75, 275.35, 273.95, 273.95, 274.05, 273.95, 274.35, 275.05, 
    274.75, 274.15, 274.25, 274.15, 274.55, 273.75, 274.35, 274.55, 275.25, 
    275.25, 274.95, 275.15, 275.35, 275.55, 275.25, 275.15, 275.25, 275.25, 
    275.05, 275.05, 275.05, 274.95, 275.35, 274.95, 274.65, 274.45, 274.15, 
    274.05, 273.95, 273.85, 273.75, 273.45, 273.55, 273.35, 273.75, 273.65, 
    273.15, 272.95, 273.45, 273.65, 273.65, 273.85, 275.05, 273.65, 273.55, 
    273.35, 272.65, 272.45, 272.05, 272.35, 271.85, 272.45, 272.15, 272.25, 
    272.75, 272.85, 272.75, 273.05, 272.75, 273.35, 273.45, 273.45, 273.95, 
    273.75, 274.05, 274.45, 272.45, 272.05, 271.65, 271.75, 271.55, 272.35, 
    272.75, 272.95, 273.25, 273.35, 273.75, 274.35, 274.25, 274.35, 274.35, 
    274.45, 274.35, 274.25, 274.55, 274.35, 274.45, 274.35, 274.15, 274.35, 
    274.15, 274.65, 275.15, 275.05, 275.45, 275.65, 276.25, 275.75, 275.65, 
    276.45, 275.15, 274.45, 275.25, 276.15, 276.55, 275.85, 275.25, 275.35, 
    275.85, 275.15, 275.05, 274.95, 274.95, 274.85, 275.05, 275.15, 275.15, 
    275.45, 275.15, 275.45, 275.95, 276.25, 276.55, 276.75, 277.25, 276.75, 
    276.15, 275.55, 275.35, 275.25, 275.75, 275.25, 275.55, 275.75, 275.75, 
    275.65, 276.05, 276.25, 275.65, 275.25, 273.45, 273.25, 273.35, 272.75, 
    272.45, 272.05, 271.75, 271.35, 270.95, 270.55, 270.45, 270.35, 270.35, 
    270.15, 270.05, 269.85, 269.85, 269.65, 269.55, 269.45, 269.45, 269.45, 
    269.55, 269.55, 269.55, 269.65, 270.05, 269.95, 270.65, 270.25, 269.45, 
    269.25, 269.65, 269.35, 269.05, 268.95, 268.75, 268.65, 268.55, 268.75, 
    268.25, 268.45, 268.15, 268.45, 268.15, 268.35, 269.45, 271.95, 271.45, 
    271.05, 271.85, 271.55, 271.95, 271.35, 271.05, 270.65, 271.25, 270.95, 
    271.05, 271.55, 272.05, 272.25, 272.65, 272.95, 273.05, 273.35, 273.35, 
    272.75, 273.65, 273.55, 273.55, 273.75, 273.75, 273.25, 273.15, 273.95, 
    273.75, 274.05, 274.35, 274.15, 274.15, 274.05, 274.15, 274.25, 274.15, 
    274.55, 274.35, 274.55, 274.35, 274.55, 274.95, 275.05, 274.85, 274.85, 
    275.05, 275.55, 275.85, 275.45, 275.15, 275.15, 274.95, 274.95, 274.85, 
    274.45, 274.45, 274.35, 274.35, 274.65, 275.15, 274.95, 274.85, 274.95, 
    274.75, 274.45, 274.35, 273.85, 274.05, 274.25, 274.15, 274.05, 274.05, 
    273.95, 273.65, 272.95, 272.65, 272.45, 272.45, 272.35, 272.15, 272.35, 
    271.95, 271.75, 272.05, 271.95, 271.55, 271.35, 271.15, 271.15, 271.05, 
    271.05, 271.25, 271.15, 271.15, 270.95, 270.85, 270.65, 269.95, 269.25, 
    269.75, 269.85, 270.05, 270.25, 269.95, 269.95, 269.85, 269.65, 270.35, 
    270.95, 271.65, 271.55, 270.45, 271.25, 270.85, 271.15, 271.25, 271.35, 
    270.85, 271.15, 271.25, 271.55, 271.75, 271.75, 272.55, 272.55, 272.35, 
    272.25, 272.25, 272.55, 272.45, 272.45, 272.25, 272.45, 272.55, 272.55, 
    272.75, 272.75, 273.05, 272.95, 273.35, 273.55, 273.65, 273.65, 273.65, 
    273.65, 273.75, 273.65, 273.55, 273.65, 273.65, 273.65, 273.75, 273.85, 
    273.75, 273.85, 274.35, 274.25, 274.25, 274.45, 275.25, 275.35, 275.35, 
    275.25, 274.95, 275.05, 275.15, 275.05, 274.95, 274.85, 274.65, 274.45, 
    274.65, 274.35, 274.35, 273.75, 274.55, 274.45, 274.95, 273.05, 273.65, 
    272.75, 272.25, 272.15, 272.65, 272.75, 273.35, 273.65, 274.05, 274.55, 
    274.75, 274.65, 274.75, 275.05, 275.55, 275.25, 274.75, 274.95, 274.75, 
    274.75, 274.75, 274.25, 273.95, 273.75, 274.75, 274.65, 275.05, 274.75, 
    274.95, 274.95, 275.15, 275.35, 275.15, 274.85, 275.25, 275.35, 275.35, 
    275.25, 275.15, 275.55, 274.85, 274.25, 274.25, 274.35, 274.35, 274.35, 
    274.45, 274.45, 274.35, 274.35, 274.25, 274.25, 274.25, 274.25, 274.25, 
    274.35, 274.05, 273.55, 273.55, 273.85, 273.55, 273.45, 273.55, 273.85, 
    273.55, 273.25, 273.25, 273.15, 273.35, 273.05, 272.85, 273.05, 273.05, 
    272.55, 272.75, 272.75, 272.85, 272.55, 272.55, 272.25, 272.45, 272.25, 
    272.25, 272.45, 272.45, 272.55, 272.45, 272.25, 272.45, 272.45, 271.85, 
    271.65, 271.85, 272.45, 272.95, 272.75, 272.65, 272.45, 272.95, 272.95, 
    273.35, 273.35, 273.45, 273.75, 273.45, 273.35, 273.85, 273.45, 273.85, 
    272.95, 272.95, 272.95, 272.45, 272.05, 271.65, 271.55, 271.65, 271.15, 
    272.05, 271.35, 270.85, 270.55, 270.55, 270.35, 270.55, 270.55, 270.15, 
    269.85, 269.45, 269.65, 269.15, 268.85, 269.55, 269.25, 269.05, 269.05, 
    268.85, 268.35, 268.35, 267.85, 268.15, 268.05, 267.95, 268.15, 268.35, 
    268.65, 268.65, 268.75, 268.65, 268.75, 268.85, 268.75, 269.25, 269.15, 
    268.75, 268.55, 268.65, 269.05, 269.45, 269.85, 270.05, 270.45, 270.55, 
    270.85, 271.15, 271.55, 271.35, 271.45, 271.75, 271.55, 271.75, 271.95, 
    272.05, 272.05, 271.95, 272.25, 272.25, 272.45, 272.35, 272.25, 272.05, 
    271.95, 272.35, 272.15, 272.45, 272.45, 272.45, 272.55, 272.75, 272.75, 
    272.85, 272.95, 272.85, 272.85, 272.95, 273.15, 273.45, 273.85, 273.65, 
    273.45, 272.95, 273.05, 272.85, 273.05, 273.85, 274.35, 274.55, 275.65, 
    273.15, 272.95, 273.15, 273.05, 272.55, 272.65, 272.15, 272.45, 272.95, 
    273.05, 273.15, 273.85, 274.45, 274.95, 274.85, 275.05, 274.85, 274.65, 
    274.65, 274.55, 274.35, 274.85, 274.95, 274.85, 275.35, 275.25, 274.95, 
    275.45, 275.15, 274.95, 275.35, 275.05, 274.85, 274.85, 274.65, 274.65, 
    273.75, 273.25, 272.75, 271.55, 270.85, 270.45, 271.05, 270.65, 271.15, 
    271.25, 271.35, 271.35, 271.25, 271.15, 271.05, 270.75, 270.95, 270.75, 
    270.95, 271.15, 271.25, 271.05, 271.05, 271.15, 271.15, 271.25, 271.45, 
    271.35, 271.55, 271.35, 271.35, 271.35, 271.25, 271.35, 271.35, 271.35, 
    271.55, 271.35, 271.25, 271.15, 271.15, 271.55, 271.45, 271.55, 271.35, 
    271.25, 271.25, 271.45, 271.65, 271.95, 272.15, 271.55, 271.45, 271.55, 
    270.95, 271.15, 270.55, 270.35, 270.45, 270.25, 269.95, 269.85, 269.65, 
    270.35, 270.85, 271.35, 271.25, 271.45, 271.55, 271.55, 271.75, 271.85, 
    271.95, 272.15, 272.15, 271.95, 271.65, 272.15, 272.25, 272.15, 272.15, 
    272.15, 272.15, 272.25, 272.15, 272.15, 272.15, 272.45, 272.45, 272.15, 
    272.45, 272.65, 273.15, 273.05, 273.65, 273.45, 273.85, 273.85, 274.45, 
    273.85, 273.85, 273.55, 274.25, 273.95, 272.95, 272.35, 273.05, 273.85, 
    274.35, 274.35, 273.85, 273.25, 272.65, 272.25, 272.25, 272.15, 271.95, 
    271.65, 271.45, 271.15, 270.95, 270.65, 270.15, 269.85, 269.75, 269.65, 
    269.75, 270.05, 269.75, 269.85, 270.05, 270.25, 270.65, 271.15, 271.05, 
    271.15, 271.35, 271.05, 271.75, 271.75, 272.15, 272.85, 273.35, 273.35, 
    273.65, 273.95, 274.25, 274.85, 274.75, 274.25, 275.25, 275.35, 275.95, 
    275.95, 276.25, 276.45, 275.75, 275.75, 276.95, 276.95, 276.65, 275.25, 
    275.65, 276.25, 276.15, 275.75, 276.15, 276.45, 276.35, 276.25, 276.75, 
    277.55, 278.25, 274.85, 275.95, 274.95, 275.05, 274.85, 275.05, 275.25, 
    274.55, 275.85, 275.05, 275.85, 274.95, 275.05, 274.75, 274.65, 274.45, 
    274.05, 274.05, 274.35, 273.75, 273.95, 273.65, 273.65, 273.25, 273.05, 
    272.85, 272.75, 272.85, 272.85, 272.25, 272.45, 272.65, 272.95, 273.25, 
    273.15, 273.45, 274.05, 274.25, 274.85, 275.75, 275.55, 275.75, 275.15, 
    276.25, 277.45, 276.85, 277.25, 278.85, 278.05, 278.55, 277.15, 276.05, 
    276.65, 277.55, 276.95, 277.55, 277.55, 277.45, 277.05, 277.35, 277.15, 
    277.45, 277.65, 278.15, 280.65, 277.95, 278.45, 277.55, 277.75, 277.55, 
    277.05, 276.55, 276.15, 276.25, 276.95, 276.45, 275.45, 276.65, 275.95, 
    276.45, 275.15, 274.05, 272.55, 272.85, 272.65, 272.55, 272.15, 272.25, 
    276.65, 274.95, 272.75, 272.45, 272.55, 272.75, 272.65, 272.25, 272.05, 
    271.65, 271.65, 271.45, 271.65, 271.85, 272.05, 274.75, 276.65, 274.45, 
    273.65, 274.65, 275.05, 275.75, 276.95, 278.05, 276.25, 276.05, 277.95, 
    278.55, 279.25, 279.25, 278.55, 276.15, 273.35, 273.95, 274.55, 273.45, 
    273.95, 273.45, 275.95, 274.65, 275.55, 273.85, 274.25, 273.55, 273.75, 
    274.35, 274.15, 273.35, 272.35, 272.05, 272.15, 272.65, 273.05, 273.85, 
    274.45, 274.55, 274.75, 275.05, 275.15, 275.15, 274.85, 274.85, 274.65, 
    274.45, 274.35, 274.25, 274.25, 274.25, 274.45, 274.15, 274.25, 274.55, 
    274.55, 275.05, 274.85, 274.85, 274.95, 274.85, 274.35, 274.35, 274.55, 
    274.55, 274.55, 274.75, 274.85, 274.95, 275.05, 275.15, 275.45, 275.65, 
    276.05, 273.95, 274.55, 273.75, 273.45, 273.25, 273.15, 273.05, 273.05, 
    273.55, 273.35, 273.35, 273.95, 272.75, 272.75, 272.45, 272.35, 273.05, 
    273.55, 272.75, 273.65, 273.45, 272.75, 272.25, 272.05, 271.55, 271.05, 
    271.15, 271.25, 271.15, 271.25, 271.05, 270.95, 270.65, 270.15, 269.25, 
    268.65, 268.45, 268.05, 267.65, 267.35, 267.55, 267.45, 267.35, 267.45, 
    267.45, 267.25, 267.45, 267.45, 267.35, 267.25, 267.05, 267.25, 267.45, 
    267.55, 267.85, 268.15, 268.35, 268.35, 268.25, 268.25, 267.85, 268.15, 
    268.65, 268.75, 268.85, 268.85, 268.75, 268.25, 267.15, 267.45, 268.55, 
    267.95, 268.75, 268.55, 268.15, 268.25, 268.35, 268.65, 268.65, 268.85, 
    268.95, 268.85, 268.95, 269.05, 268.95, 269.05, 268.95, 268.95, 269.15, 
    269.05, 269.15, 269.25, 269.15, 269.25, 269.25, 269.25, 269.35, 269.25, 
    269.15, 269.05, 268.85, 267.85, 267.45, 268.05, 267.85, 268.05, 267.25, 
    267.75, 267.35, 267.55, 267.65, 267.85, 267.75, 267.85, 267.85, 267.75, 
    268.05, 268.35, 268.45, 268.55, 268.75, 268.85, 268.95, 268.85, 268.65, 
    268.55, 268.45, 268.35, 268.65, 268.85, 268.65, 268.75, 268.95, 269.35, 
    269.85, 270.55, 270.85, 272.15, 272.35, 272.25, 272.35, 272.45, 272.15, 
    271.45, 271.25, 271.35, 271.65, 271.45, 271.55, 272.45, 272.55, 272.35, 
    272.45, 272.55, 272.45, 272.85, 272.75, 272.95, 273.15, 273.25, 273.25, 
    273.75, 273.55, 273.65, 273.95, 274.15, 274.55, 274.35, 275.75, 273.45, 
    273.55, 275.95, 274.65, 274.15, 274.35, 274.15, 273.45, 273.05, 273.25, 
    272.65, 272.65, 272.55, 272.45, 272.75, 272.15, 272.35, 272.85, 272.85, 
    272.85, 272.95, 273.25, 273.25, 273.15, 273.05, 272.95, 272.95, 273.05, 
    273.05, 272.85, 272.55, 272.75, 273.15, 272.95, 272.85, 272.55, 272.45, 
    272.45, 272.15, 272.05, 272.25, 272.35, 271.95, 272.15, 271.85, 272.15, 
    272.15, 272.15, 272.15, 272.15, 272.05, 271.95, 272.15, 272.05, 272.05, 
    272.05, 271.95, 272.15, 272.25, 272.15, 272.15, 272.05, 272.15, 272.05, 
    272.05, 272.05, 272.15, 272.55, 272.55, 272.05, 272.35, 272.25, 272.35, 
    272.45, 272.15, 272.15, 272.15, 272.25, 272.25, 272.25, 272.25, 272.25, 
    272.05, 271.65, 271.45, 271.65, 271.35, 271.65, 271.75, 271.95, 271.95, 
    272.05, 272.05, 272.25, 272.35, 272.25, 272.15, 272.05, 272.15, 272.05, 
    272.25, 272.25, 272.45, 272.75, 272.95, 272.85, 272.85, 272.75, 272.65, 
    272.55, 272.45, 272.35, 272.45, 272.45, 272.55, 272.55, 272.45, 272.25, 
    272.25, 272.05, 272.05, 272.05, 271.85, 271.85, 271.85, 271.75, 271.65, 
    271.85, 272.05, 272.35, 272.65, 272.55, 272.65, 272.55, 272.65, 272.55, 
    272.45, 272.35, 272.05, 271.95, 271.95, 271.95, 272.05, 272.15, 272.15, 
    271.95, 271.95, 271.85, 271.95, 271.95, 271.75, 271.65, 271.55, 271.55, 
    271.65, 271.65, 271.65, 271.55, 271.35, 271.05, 271.05, 270.95, 270.65, 
    270.65, 270.55, 270.25, 270.35, 270.35, 270.35, 270.25, 270.35, 270.45, 
    270.35, 270.25, 270.15, 270.45, 270.05, 269.75, 269.55, 269.45, 269.35, 
    268.85, 268.75, 268.25, 267.45, 267.85, 267.95, 267.55, 268.05, 267.25, 
    268.15, 265.15, 266.35, 266.95, 266.55, 265.85, 265.95, 266.15, 266.25, 
    266.15, 266.55, 266.65, 267.35, 268.15, 268.35, 268.55, 268.25, 267.85, 
    267.75, 267.95, 268.05, 267.75, 267.25, 267.05, 267.05, 267.25, 267.25, 
    267.05, 266.85, 266.75, 266.75, 266.75, 266.95, 266.45, 266.45, 266.05, 
    265.95, 266.15, 265.85, 265.45, 265.35, 265.35, 265.15, 265.05, 264.75, 
    264.45, 264.25, 264.35, 264.45, 264.45, 265.05, 265.35, 265.35, 265.35, 
    265.45, 265.55, 265.55, 265.55, 265.65, 265.75, 265.75, 266.05, 266.15, 
    266.35, 266.35, 266.55, 266.85, 267.15, 267.25, 267.95, 268.05, 268.65, 
    269.15, 269.75, 270.05, 270.15, 270.75, 270.75, 271.15, 271.25, 271.45, 
    271.55, 271.65, 271.75, 271.65, 271.55, 271.65, 271.75, 272.25, 272.55, 
    272.75, 273.25, 274.85, 273.95, 273.65, 273.35, 273.35, 273.75, 274.65, 
    274.45, 274.35, 275.05, 275.25, 274.95, 274.25, 273.75, 272.75, 272.05, 
    271.85, 271.45, 270.95, 270.55, 270.25, 269.65, 269.05, 268.85, 268.45, 
    268.05, 268.15, 267.75, 267.65, 267.45, 267.85, 267.85, 267.65, 267.65, 
    267.55, 267.45, 267.25, 267.15, 267.05, 267.05, 266.85, 266.65, 266.25, 
    266.15, 266.05, 265.85, 265.65, 265.45, 265.25, 265.25, 265.15, 265.15, 
    265.05, 264.85, 264.75, 264.55, 264.65, 264.55, 264.65, 264.55, 264.55, 
    264.45, 264.75, 264.75, 264.75, 264.95, 264.85, 264.45, 264.45, 264.35, 
    264.65, 264.75, 264.75, 264.95, 265.05, 264.75, 264.35, 264.65, 264.35, 
    264.15, 264.15, 264.65, 264.85, 265.55, 266.15, 266.35, 266.95, 267.05, 
    267.35, 267.35, 266.95, 266.65, 266.45, 266.35, 266.75, 266.85, 267.05, 
    267.15, 267.15, 267.25, 267.25, 267.15, 266.85, 267.05, 266.95, 266.85, 
    267.25, 267.05, 266.95, 267.25, 267.25, 267.65, 267.45, 267.15, 266.45, 
    266.85, 266.25, 265.55, 265.25, 265.05, 265.05, 264.95, 265.05, 265.45, 
    266.05, 266.45, 266.85, 266.65, 266.45, 266.05, 265.95, 265.85, 265.65, 
    265.45, 265.15, 265.25, 265.55, 266.35, 267.05, 267.55, 267.95, 268.05, 
    267.85, 267.45, 266.85, 266.75, 266.75, 266.65, 266.35, 266.25, 266.25, 
    266.55, 266.75, 267.05, 267.65, 268.15, 268.55, 269.75, 270.35, 271.95, 
    271.95, 271.65, 271.55, 271.25, 270.95, 270.85, 270.85, 270.75, 270.75, 
    270.75, 270.75, 270.75, 270.85, 271.05, 271.05, 271.15, 271.05, 270.85, 
    270.45, 270.15, 269.85, 269.65, 269.55, 270.05, 270.65, 270.85, 270.75, 
    270.55, 270.35, 270.25, 270.55, 270.95, 270.95, 270.45, 270.05, 270.65, 
    271.45, 271.05, 270.95, 270.75, 270.55, 271.05, 270.85, 270.75, 270.45, 
    270.75, 270.75, 270.15, 270.35, 269.65, 270.25, 270.55, 269.95, 270.55, 
    270.65, 270.85, 270.75, 270.75, 270.75, 270.85, 270.75, 270.65, 270.65, 
    270.75, 270.85, 270.75, 270.45, 270.25, 270.15, 270.05, 270.05, 270.05, 
    269.95, 269.95, 269.95, 269.95, 270.05, 269.95, 269.75, 269.55, 269.45, 
    269.35, 268.85, 268.85, 269.05, 268.95, 268.75, 268.75, 268.35, 268.05, 
    268.05, 268.15, 268.25, 268.25, 268.55, 268.25, 268.35, 268.25, 268.05, 
    268.45, 268.45, 268.25, 268.75, 269.65, 270.15, 271.05, 271.15, 271.25, 
    271.15, 271.25, 270.85, 270.55, 270.35, 270.35, 270.35, 269.85, 269.45, 
    269.45, 269.65, 269.75, 269.85, 269.95, 269.75, 269.75, 269.85, 270.05, 
    270.25, 270.35, 270.45, 270.65, 270.95, 271.05, 270.95, 271.05, 270.95, 
    270.75, 270.25, 270.45, 270.15, 270.25, 269.65, 268.65, 268.55, 268.35, 
    268.65, 268.55, 268.65, 268.45, 268.35, 267.95, 267.95, 268.05, 268.65, 
    269.15, 269.35, 270.05, 270.45, 270.65, 270.75, 271.15, 271.05, 271.25, 
    270.95, 270.65, 270.35, 270.35, 270.35, 270.65, 270.55, 270.25, 270.35, 
    270.15, 270.95, 270.65, 269.75, 269.65, 269.55, 270.05, 270.45, 270.05, 
    270.05, 270.35, 270.15, 270.05, 269.75, 269.55, 269.35, 269.45, 269.75, 
    269.85, 269.55, 269.35, 269.35, 269.55, 269.25, 269.05, 268.95, 269.05, 
    269.25, 269.65, 269.05, 269.05, 268.85, 269.05, 269.05, 268.95, 268.55, 
    267.35, 267.45, 266.55, 266.65, 265.85, 266.25, 265.25, 265.15, 266.25, 
    267.05, 266.45, 265.95, 267.45, 267.35, 266.95, 266.85, 267.45, 268.05, 
    267.85, 267.75, 268.05, 268.25, 267.65, 267.25, 266.45, 266.85, 266.25, 
    266.15, 265.65, 265.05, 265.45, 265.75, 265.25, 265.55, 265.25, 265.05, 
    265.05, 265.25, 265.95, 265.85, 266.75, 267.75, 267.05, 266.95, 267.75, 
    267.35, 267.65, 268.75, 268.55, 268.85, 269.05, 268.75, 268.65, 268.65, 
    268.75, 268.95, 268.95, 268.75, 268.95, 268.45, 268.45, 268.45, 268.85, 
    269.15, 269.25, 269.65, 270.25, 270.75, 271.65, 271.45, 271.15, 270.55, 
    269.55, 269.55, 268.85, 269.75, 269.35, 269.35, 269.15, 268.85, 268.35, 
    268.25, 268.35, 268.45, 268.55, 268.15, 268.25, 268.35, 268.25, 268.25, 
    268.25, 267.85, 267.75, 267.85, 268.05, 268.05, 268.25, 268.35, 268.55, 
    268.65, 268.65, 269.05, 269.15, 269.25, 269.25, 269.55, 269.45, 269.55, 
    269.25, 269.45, 269.65, 269.75, 269.75, 269.65, 269.75, 270.25, 270.35, 
    270.55, 270.55, 270.65, 270.75, 270.85, 270.95, 271.25, 271.45, 271.75, 
    272.05, 272.35, 272.45, 272.15, 272.25, 272.25, 272.15, 272.25, 272.05, 
    272.05, 272.25, 272.45, 272.45, 272.55, 272.45, 272.65, 272.45, 271.75, 
    272.05, 271.85, 272.25, 272.25, 272.35, 272.25, 272.55, 272.65, 272.55, 
    272.75, 272.45, 272.65, 271.95, 271.95, 271.95, 272.35, 271.65, 272.05, 
    272.95, 272.25, 271.75, 272.75, 272.85, 273.35, 273.45, 273.45, 273.15, 
    273.05, 273.45, 273.45, 273.25, 273.25, 273.35, 273.35, 273.15, 272.85, 
    272.45, 272.35, 272.25, 272.25, 272.15, 271.65, 271.55, 271.55, 271.45, 
    270.75, 271.15, 270.85, 270.45, 270.35, 270.95, 271.75, 272.45, 272.65, 
    272.65, 272.45, 272.35, 271.95, 271.75, 271.55, 271.35, 271.05, 270.65, 
    270.25, 269.75, 269.85, 269.85, 269.15, 269.35, 269.25, 268.75, 269.45, 
    269.35, 269.05, 269.05, 268.85, 268.85, 268.45, 268.45, 268.15, 268.05, 
    267.95, 267.95, 267.75, 268.05, 267.75, 267.75, 267.75, 267.75, 267.65, 
    267.75, 267.45, 267.35, 267.45, 267.75, 267.65, 267.75, 267.95, 268.25, 
    268.35, 268.05, 268.75, 268.55, 268.95, 268.85, 268.65, 268.45, 268.55, 
    268.55, 268.85, 268.75, 268.65, 268.45, 268.25, 268.25, 268.15, 267.95, 
    268.05, 268.25, 268.25, 268.25, 268.25, 267.95, 267.95, 267.95, 267.85, 
    267.65, 267.15, 267.65, 267.35, 266.85, 266.45, 266.65, 266.45, 266.25, 
    266.05, 264.65, 265.35, 266.25, 266.15, 266.05, 265.25, 265.25, 265.15, 
    264.65, 264.65, 263.85, 263.15, 262.95, 263.45, 263.85, 265.35, 265.75, 
    264.75, 265.55, 265.55, 265.75, 264.65, 265.35, 264.45, 264.65, 265.15, 
    266.25, 266.65, 265.65, 264.65, 263.85, 263.65, 263.55, 264.25, 263.55, 
    263.75, 264.05, 264.85, 265.75, 265.55, 264.85, 265.45, 265.35, 265.15, 
    266.15, 267.55, 267.45, 267.05, 266.35, 265.95, 265.95, 265.35, 265.35, 
    264.65, 264.85, 263.75, 263.15, 263.75, 263.35, 263.25, 264.85, 265.15, 
    263.85, 263.65, 264.45, 265.65, 266.35, 266.85, 266.45, 267.15, 265.45, 
    266.65, 266.35, 265.45, 265.25, 265.45, 265.45, 264.85, 265.25, 264.55, 
    265.05, 264.65, 265.35, 265.55, 265.05, 265.55, 264.55, 265.35, 264.15, 
    265.45, 265.45, 265.95, 265.65, 265.85, 266.45, 266.55, 266.95, 267.55, 
    267.45, 266.85, 266.55, 266.35, 266.25, 266.35, 265.95, 265.65, 265.25, 
    265.65, 265.45, 265.55, 265.45, 265.75, 265.45, 265.85, 265.65, 265.45, 
    265.65, 264.85, 265.25, 265.45, 265.45, 265.15, 265.05, 265.05, 265.15, 
    264.85, 264.95, 265.05, 265.05, 265.15, 265.25, 264.95, 264.95, 265.25, 
    264.65, 264.75, 264.95, 264.85, 264.55, 264.55, 264.25, 264.25, 264.25, 
    264.15, 264.05, 264.15, 264.55, 264.95, 265.25, 265.65, 265.75, 266.05, 
    266.15, 266.35, 266.45, 266.55, 266.45, 266.55, 266.75, 266.75, 266.85, 
    266.85, 266.85, 266.85, 266.85, 266.85, 266.75, 266.65, 266.65, 266.65, 
    266.65, 266.75, 266.85, 267.15, 267.25, 267.35, 267.25, 267.55, 267.25, 
    267.45, 267.65, 267.75, 268.15, 268.95, 269.65, 269.55, 269.25, 269.25, 
    268.05, 266.35, 266.95, 265.45, 264.95, 263.85, 264.95, 265.25, 265.25, 
    264.95, 264.35, 264.05, 263.65, 262.95, 262.65, 262.05, 261.35, 261.75, 
    260.25, 260.65, 261.65, 262.95, 262.15, 261.45, 260.55, 259.45, 258.65, 
    258.25, 258.15, 258.25, 259.25, 260.15, 259.45, 258.75, 259.45, 260.95, 
    262.75, 267.25, 267.75, 267.15, 265.55, 265.25, 264.75, 263.55, 263.15, 
    262.85, 262.45, 262.35, 261.95, 261.05, 260.25, 259.15, 259.15, 259.05, 
    258.75, 258.25, 257.25, 257.95, 257.55, 257.35, 256.55, 256.35, 256.55, 
    257.25, 257.75, 258.45, 257.75, 258.75, 258.05, 259.95, 258.05, 259.05, 
    258.95, 257.65, 258.25, 259.25, 260.05, 260.75, 260.85, 260.75, 261.65, 
    261.85, 262.75, 263.15, 263.65, 264.05, 263.55, 262.95, 262.25, 261.65, 
    261.75, 260.95, 260.65, 260.75, 260.75, 260.85, 260.15, 260.75, 260.45, 
    260.95, 261.45, 262.25, 263.05, 262.85, 262.95, 261.65, 262.25, 262.25, 
    262.05, 262.55, 263.05, 263.45, 263.55, 263.55, 263.65, 263.95, 264.35, 
    264.95, 266.15, 268.95, 269.75, 269.85, 269.95, 271.05, 271.65, 271.85, 
    272.05, 272.15, 271.75, 271.65, 271.55, 271.45, 271.05, 270.55, 270.35, 
    270.55, 270.75, 270.95, 271.35, 271.25, 271.35, 271.45, 271.65, 271.85, 
    272.15, 272.05, 272.25, 272.05, 271.95, 271.65, 271.65, 271.35, 271.35, 
    271.15, 271.15, 271.05, 270.75, 270.75, 270.65, 270.45, 270.25, 270.15, 
    270.05, 269.65, 269.05, 269.15, 269.15, 269.25, 269.35, 269.55, 269.15, 
    269.65, 269.85, 269.75, 269.85, 270.25, 269.85, 269.45, 269.35, 268.95, 
    268.85, 268.75, 268.85, 268.95, 269.05, 268.75, 268.65, 268.65, 268.95, 
    268.85, 268.65, 268.15, 267.35, 266.65, 266.25, 265.95, 265.45, 266.05, 
    265.55, 265.15, 264.65, 265.65, 266.05, 266.55, 266.95, 267.75, 268.25, 
    268.15, 267.85, 267.05, 266.05, 265.75, 265.75, 265.75, 265.95, 265.65, 
    265.95, 266.55, 266.75, 266.65, 266.75, 266.55, 266.55, 266.65, 266.85, 
    266.45, 266.75, 266.75, 266.45, 266.35, 266.35, 266.05, 266.25, 266.35, 
    266.25, 266.35, 266.35, 266.35, 266.25, 266.35, 266.35, 266.25, 266.35, 
    266.15, 265.85, 266.05, 265.85, 266.05, 265.95, 265.65, 265.55, 265.45, 
    265.45, 265.45, 265.25, 265.25, 265.15, 265.45, 265.75, 265.95, 266.75, 
    266.35, 266.75, 266.65, 267.05, 267.05, 267.35, 267.45, 267.55, 267.45, 
    267.45, 267.25, 266.55, 266.85, 266.85, 266.95, 266.95, 266.45, 267.15, 
    267.05, 267.25, 267.45, 267.75, 267.95, 267.75, 268.05, 268.05, 268.35, 
    268.75, 268.25, 267.85, 268.05, 267.85, 267.75, 267.75, 267.55, 267.45, 
    267.25, 267.15, 267.25, 266.85, 266.55, 267.05, 267.05, 266.85, 266.65, 
    266.55, 266.45, 266.75, 266.05, 266.15, 265.85, 265.85, 265.65, 265.65, 
    265.55, 265.45, 265.45, 265.45, 264.65, 265.05, 265.25, 264.95, 265.15, 
    265.25, 265.45, 265.95, 266.15, 265.95, 265.75, 265.45, 265.85, 265.85, 
    265.85, 266.25, 266.25, 266.35, 266.35, 266.35, 266.35, 265.85, 265.55, 
    265.35, 265.05, 264.65, 264.05, 264.15, 264.05, 264.45, 264.25, 264.45, 
    265.05, 266.55, 266.95, 267.15, 267.05, 267.45, 267.35, 267.45, 267.45, 
    267.45, 266.95, 266.85, 266.95, 267.25, 267.55, 267.75, 267.35, 267.95, 
    267.95, 267.95, 267.85, 267.75, 268.95, 269.15, 268.55, 268.75, 268.65, 
    268.55, 267.95, 267.15, 266.65, 266.05, 265.55, 264.95, 264.05, 263.85, 
    263.85, 264.05, 264.95, 265.15, 265.35, 265.65, 266.55, 268.05, 268.35, 
    269.15, 269.45, 269.75, 270.15, 270.65, 270.35, 270.55, 271.55, 272.25, 
    272.35, 272.15, 272.35, 271.95, 271.95, 271.55, 271.15, 271.05, 270.45, 
    270.35, 269.55, 267.95, 266.45, 265.05, 264.15, 263.45, 262.95, 261.55, 
    261.95, 261.35, 260.45, 260.85, 260.95, 260.85, 260.95, 260.85, 260.95, 
    260.65, 260.35, 260.45, 260.35, 260.45, 260.45, 260.15, 260.25, 259.95, 
    259.85, 259.95, 259.95, 260.55, 260.35, 259.75, 259.45, 258.35, 257.85, 
    257.65, 257.75, 258.05, 260.55, 261.05, 261.05, 261.05, 261.45, 260.65, 
    261.15, 261.05, 260.65, 260.75, 260.95, 260.65, 260.45, 260.15, 259.95, 
    260.25, 260.15, 260.05, 259.65, 259.35, 259.15, 258.95, 258.85, 258.85, 
    258.95, 258.75, 258.85, 259.15, 259.45, 259.45, 259.35, 259.45, 259.55, 
    259.35, 260.45, 260.65, 261.55, 261.45, 261.45, 261.35, 262.45, 262.75, 
    263.15, 263.25, 263.65, 263.85, 263.95, 264.15, 264.95, 265.85, 265.75, 
    267.25, 267.55, 267.55, 268.05, 269.05, 269.25, 269.75, 270.55, 271.25, 
    271.25, 271.15, 271.35, 271.35, 271.55, 271.25, 271.25, 271.25, 271.15, 
    271.05, 270.95, 271.05, 270.95, 270.95, 270.85, 269.25, 268.55, 268.15, 
    266.95, 266.85, 266.55, 265.05, 264.95, 266.65, 266.65, 265.95, 266.25, 
    266.05, 267.15, 267.65, 267.95, 268.75, 269.25, 268.35, 269.25, 269.45, 
    269.15, 268.65, 268.85, 268.75, 270.15, 270.65, 271.05, 271.25, 271.25, 
    271.45, 271.45, 271.35, 271.15, 270.95, 270.95, 271.15, 271.15, 271.35, 
    271.35, 271.55, 272.05, 272.05, 272.15, 272.15, 272.05, 272.15, 272.05, 
    271.95, 271.95, 271.95, 271.85, 271.65, 271.75, 271.75, 271.65, 271.55, 
    271.75, 271.15, 271.35, 271.35, 271.35, 271.15, 271.15, 271.05, 271.15, 
    271.15, 271.55, 271.55, 271.35, 271.45, 271.55, 271.55, 271.55, 271.55, 
    271.45, 271.35, 271.55, 271.35, 271.25, 271.35, 271.55, 271.75, 271.85, 
    271.75, 271.65, 271.55, 270.55, 271.25, 270.65, 270.95, 271.45, 271.45, 
    271.65, 271.75, 271.95, 271.95, 271.95, 271.85, 271.65, 271.65, 272.15, 
    271.85, 272.05, 272.05, 272.05, 271.95, 271.85, 271.95, 271.85, 271.65, 
    271.75, 271.85, 271.65, 271.55, 271.45, 271.35, 271.05, 270.55, 270.25, 
    269.55, 269.65, 269.75, 269.35, 268.95, 268.55, 268.95, 268.85, 268.05, 
    267.95, 267.85, 267.45, 267.25, 266.65, 266.35, 266.05, 265.85, 265.45, 
    265.15, 265.45, 265.05, 265.25, 265.25, 264.95, 265.25, 265.05, 264.95, 
    265.45, 265.85, 266.35, 266.75, 267.15, 267.35, 267.75, 268.15, 268.75, 
    268.95, 269.65, 269.65, 269.05, 268.45, 267.85, 267.25, 264.75, 263.75, 
    263.45, 263.05, 262.75, 262.95, 262.55, 263.95, 264.55, 264.35, 264.25, 
    263.65, 263.35, 262.95, 263.15, 261.95, 262.35, 262.05, 263.05, 263.55, 
    263.25, 263.05, 264.85, 265.75, 266.45, 266.55, 266.65, 264.55, 262.75, 
    262.45, 262.55, 263.45, 263.65, 264.05, 262.65, 261.05, 259.75, 257.65, 
    256.45, 255.35, 254.75, 253.75, 253.15, 253.45, 252.65, 253.05, 252.65, 
    252.15, 252.35, 252.55, 253.65, 255.05, 255.05, 255.35, 255.75, 256.05, 
    256.05, 255.85, 256.35, 258.25, 259.05, 259.55, 261.35, 262.45, 264.35, 
    263.85, 263.65, 263.45, 263.15, 263.15, 262.35, 262.55, 262.95, 262.05, 
    262.25, 261.45, 261.25, 262.45, 262.85, 261.45, 262.05, 261.55, 261.15, 
    260.95, 261.25, 259.55, 258.05, 257.35, 256.65, 256.55, 254.95, 256.25, 
    257.05, 256.55, 256.45, 256.85, 256.65, 256.45, 256.85, 257.05, 257.15, 
    257.15, 257.45, 257.35, 257.45, 257.65, 257.25, 257.55, 257.65, 257.95, 
    258.15, 258.45, 258.65, 259.05, 259.35, 259.15, 259.05, 258.45, 258.05, 
    258.15, 257.95, 257.95, 256.95, 257.55, 258.15, 258.15, 258.65, 258.45, 
    258.05, 258.25, 257.95, 258.05, 257.75, 257.65, 257.95, 257.55, 257.55, 
    257.25, 256.85, 256.45, 256.25, 256.35, 256.05, 255.85, 255.95, 255.95, 
    255.85, 255.45, 255.45, 255.15, 254.45, 253.85, 253.55, 253.95, 254.45, 
    254.35, 253.35, 254.95, 256.25, 256.25, 253.75, 254.25, 254.55, 254.85, 
    254.85, 256.05, 255.95, 256.65, 256.25, 256.55, 255.95, 257.05, 256.35, 
    257.05, 257.15, 257.65, 258.95, 258.75, 259.15, 259.45, 259.55, 259.15, 
    259.65, 260.45, 259.75, 260.85, 260.05, 260.55, 260.55, 259.35, 257.95, 
    259.25, 256.15, 256.95, 255.75, 255.85, 255.95, 255.75, 255.55, 256.55, 
    256.35, 256.45, 256.05, 256.25, 255.95, 256.05, 255.95, 255.85, 255.95, 
    255.55, 255.45, 255.85, 256.35, 256.35, 256.15, 256.35, 256.65, 256.95, 
    256.65, 256.95, 257.05, 256.95, 256.65, 256.35, 256.15, 256.55, 256.25, 
    256.35, 256.15, 255.35, 254.65, 254.65, 254.95, 255.05, 254.35, 253.85, 
    253.85, 253.75, 253.45, 252.75, 251.95, 252.05, 251.85, 252.05, 253.05, 
    252.05, 251.35, 251.75, 251.95, 251.35, 251.35, 251.15, 251.25, 251.65, 
    251.35, 251.95, 253.45, 254.05, 254.45, 254.85, 255.05, 255.45, 255.25, 
    255.15, 255.55, 255.45, 254.45, 254.55, 254.45, 253.55, 254.55, 254.35, 
    255.35, 255.45, 254.85, 255.25, 254.65, 254.45, 255.35, 256.45, 258.35, 
    258.35, 257.35, 258.25, 258.75, 258.85, 259.85, 259.75, 260.35, 262.45, 
    262.95, 263.05, 263.05, 263.55, 265.25, 264.85, 264.85, 264.95, 264.65, 
    263.95, 264.05, 263.35, 263.35, 263.25, 263.15, 262.95, 263.15, 263.75, 
    264.15, 263.95, 263.55, 261.75, 264.75, 266.45, 267.05, 267.55, 267.75, 
    267.85, 267.75, 267.65, 268.05, 267.95, 268.25, 268.65, 268.85, 268.75, 
    269.45, 269.45, 269.05, 269.35, 269.25, 269.05, 269.05, 268.95, 269.25, 
    269.15, 268.85, 269.15, 269.05, 269.15, 268.85, 269.05, 268.95, 268.45, 
    268.45, 268.45, 268.05, 268.15, 268.45, 268.55, 267.75, 267.35, 267.45, 
    267.45, 267.35, 267.35, 267.35, 267.05, 267.35, 267.55, 267.65, 267.85, 
    268.05, 268.15, 268.25, 268.35, 268.45, 268.25, 268.25, 268.05, 268.05, 
    268.05, 267.95, 267.75, 267.65, 267.55, 267.25, 266.75, 266.75, 266.85, 
    267.35, 267.55, 268.15, 268.05, 268.35, 268.45, 268.55, 268.55, 268.75, 
    269.05, 269.45, 269.65, 269.95, 270.05, 270.25, 270.25, 270.15, 270.15, 
    269.95, 269.75, 269.25, 268.85, 268.85, 269.25, 268.25, 269.05, 269.25, 
    269.65, 269.85, 269.05, 268.05, 270.05, 270.35, 270.55, 270.35, 269.25, 
    269.05, 269.15, 269.25, 269.15, 269.15, 268.75, 269.55, 270.95, 270.95, 
    270.75, 270.55, 270.35, 270.35, 269.25, 268.55, 268.65, 268.75, 270.05, 
    268.75, 268.55, 267.55, 266.95, 267.75, 268.05, 268.25, 269.05, 269.25, 
    269.85, 269.95, 271.25, 271.45, 270.65, 270.35, 270.65, 270.45, 270.35, 
    270.25, 270.35, 270.55, 270.05, 270.45, 271.15, 271.55, 272.15, 272.65, 
    272.95, 273.05, 273.05, 272.75, 273.25, 273.45, 273.65, 273.75, 273.75, 
    273.75, 273.65, 273.05, 272.75, 272.35, 272.35, 272.25, 271.35, 271.05, 
    271.05, 271.45, 270.95, 270.15, 269.95, 269.45, 268.75, 268.95, 268.85, 
    268.35, 267.85, 268.35, 267.35, 267.65, 267.35, 267.55, 267.55, 267.25, 
    267.45, 267.15, 268.05, 267.35, 268.25, 267.95, 268.45, 268.55, 268.75, 
    269.15, 269.85, 270.05, 269.85, 270.75, 270.65, 270.65, 270.05, 270.35, 
    270.95, 271.25, 271.55, 271.55, 272.25, 271.75, 271.95, 271.95, 272.25, 
    272.85, 272.25, 272.95, 272.45, 271.75, 271.65, 271.75, 271.85, 271.75, 
    271.75, 271.35, 271.35, 270.75, 270.35, 270.05, 270.15, 270.25, 270.25, 
    270.05, 269.65, 269.25, 268.95, 268.75, 268.45, 268.35, 268.15, 267.75, 
    267.45, 267.45, 267.65, 267.65, 267.55, 266.45, 265.65, 266.05, 265.75, 
    265.85, 266.15, 265.85, 265.45, 265.35, 265.45, 265.45, 265.25, 265.55, 
    265.85, 266.55, 267.15, 268.25, 269.15, 269.65, 269.25, 269.45, 268.65, 
    268.45, 268.25, 268.35, 268.65, 269.05, 269.55, 269.95, 270.75, 271.35, 
    271.55, 271.55, 271.85, 271.95, 271.45, 271.25, 271.35, 271.75, 271.15, 
    271.05, 271.15, 271.05, 270.55, 270.95, 271.05, 270.85, 270.05, 269.75, 
    269.15, 269.15, 269.25, 269.15, 270.05, 270.05, 269.55, 269.05, 268.45, 
    266.95, 265.95, 266.55, 267.75, 268.15, 268.25, 268.05, 268.05, 268.15, 
    268.35, 268.75, 269.45, 269.65, 269.85, 270.05, 270.45, 270.35, 270.55, 
    270.25, 270.15, 270.15, 270.65, 271.35, 271.45, 270.55, 270.55, 270.95, 
    270.35, 269.55, 267.85, 267.95, 267.85, 268.45, 268.65, 268.65, 268.95, 
    268.75, 268.95, 270.05, 270.05, 270.75, 270.65, 270.55, 269.65, 269.45, 
    269.45, 270.15, 270.55, 270.75, 271.15, 271.05, 271.45, 271.15, 271.05, 
    271.15, 271.25, 271.25, 271.05, 270.85, 270.65, 270.75, 270.55, 271.25, 
    270.45, 270.55, 270.65, 270.25, 270.35, 270.65, 270.45, 270.55, 270.35, 
    270.25, 270.25, 269.65, 269.45, 269.75, 269.75, 269.25, 269.15, 269.65, 
    270.15, 270.35, 270.35, 270.15, 269.95, 270.05, 269.85, 269.75, 269.85, 
    269.75, 269.75, 269.65, 269.75, 269.65, 269.55, 269.35, 269.35, 268.65, 
    268.75, 268.25, 268.05, 267.95, 267.65, 267.55, 267.65, 267.05, 267.25, 
    266.75, 267.75, 268.45, 268.65, 268.05, 267.65, 267.45, 267.75, 267.75, 
    267.05, 266.85, 266.75, 266.35, 265.25, 265.35, 265.65, 265.55, 265.05, 
    264.85, 265.05, 264.85, 264.95, 263.95, 263.25, 262.85, 263.25, 262.35, 
    262.35, 261.95, 261.65, 261.55, 261.05, 262.95, 262.15, 262.15, 261.15, 
    259.05, 257.25, 255.05, 254.25, 256.15, 257.65, 258.15, 257.75, 257.45, 
    257.35, 257.75, 257.95, 258.05, 257.75, 258.35, 258.15, 257.65, 257.65, 
    257.25, 257.65, 257.45, 258.15, 258.05, 258.45, 259.15, 259.15, 258.85, 
    260.65, 262.55, 261.15, 261.25, 261.15, 261.15, 261.45, 261.85, 261.75, 
    261.25, 262.15, 261.55, 257.65, 257.35, 255.65, 255.05, 256.85, 256.45, 
    255.95, 256.25, 256.35, 256.25, 255.15, 255.35, 256.65, 255.85, 255.05, 
    255.35, 256.25, 257.15, 257.65, 257.45, 255.35, 255.65, 255.35, 255.95, 
    256.15, 256.05, 255.85, 255.75, 255.75, 255.45, 255.65, 255.15, 254.85, 
    254.55, 254.25, 254.65, 253.15, 253.25, 254.05, 253.95, 253.45, 253.25, 
    254.35, 253.45, 252.55, 252.55, 252.05, 252.75, 252.95, 253.05, 253.35, 
    252.95, 253.25, 253.95, 253.85, 253.65, 253.35, 253.85, 254.45, 254.15, 
    254.25, 253.65, 253.85, 254.05, 254.05, 253.75, 253.85, 253.85, 253.85, 
    253.35, 252.35, 251.15, 251.45, 251.85, 251.15, 250.55, 251.05, 251.35, 
    251.85, 251.35, 250.85, 251.35, 251.85, 252.25, 252.35, 252.05, 253.25, 
    253.35, 253.45, 252.95, 252.75, 252.65, 253.25, 253.25, 251.25, 251.75, 
    251.65, 251.75, 251.05, 251.15, 251.25, 251.15, 250.65, 251.35, 251.65, 
    251.65, 251.95, 251.65, 252.25, 252.25, 252.05, 251.95, 252.15, 251.95, 
    252.45, 253.15, 253.45, 252.75, 252.95, 252.95, 252.95, 253.05, 253.75, 
    253.85, 253.75, 253.75, 253.25, 253.65, 254.05, 253.95, 253.85, 253.65, 
    253.35, 253.85, 253.45, 254.05, 254.45, 254.85, 254.75, 254.95, 254.75, 
    254.55, 254.75, 255.15, 255.85, 256.45, 256.65, 256.75, 256.85, 257.45, 
    258.35, 259.15, 259.35, 260.15, 260.85, 261.25, 261.75, 261.65, 260.55, 
    265.95, 261.95, 262.35, 262.65, 262.35, 262.85, 263.65, 263.55, 265.85, 
    264.65, 265.45, 264.95, 266.55, 266.95, 267.35, 267.75, 268.25, 267.75, 
    268.75, 268.35, 267.95, 268.45, 268.85, 269.65, 269.55, 269.65, 269.95, 
    270.45, 270.85, 270.95, 270.95, 270.95, 270.95, 271.25, 271.25, 271.35, 
    271.55, 271.75, 271.05, 270.25, 270.95, 271.15, 271.15, 271.35, 271.65, 
    271.85, 272.15, 272.25, 272.55, 272.95, 273.75, 273.75, 273.05, 272.75, 
    272.65, 272.65, 272.45, 272.25, 272.15, 271.65, 270.75, 270.45, 269.95, 
    268.75, 267.75, 267.85, 267.85, 267.75, 267.75, 267.45, 267.35, 267.55, 
    267.05, 266.55, 266.65, 266.55, 265.95, 266.55, 265.85, 265.65, 265.95, 
    265.95, 265.15, 264.95, 264.45, 265.05, 265.85, 266.75, 267.55, 267.95, 
    267.85, 267.15, 266.05, 266.35, 266.35, 266.35, 266.45, 266.45, 266.65, 
    266.75, 267.15, 267.55, 267.65, 267.85, 268.25, 269.05, 270.15, 270.55, 
    270.75, 270.75, 270.95, 271.05, 270.85, 270.95, 270.75, 270.85, 270.85, 
    270.55, 270.25, 269.65, 269.25, 269.05, 268.65, 268.85, 269.25, 268.95, 
    268.85, 268.05, 267.25, 267.15, 266.75, 267.25, 267.85, 269.05, 269.05, 
    269.05, 268.55, 269.45, 269.25, 269.15, 268.85, 268.35, 267.65, 267.35, 
    266.45, 265.45, 265.45, 265.45, 266.45, 266.15, 266.35, 266.25, 266.75, 
    268.25, 267.95, 267.95, 268.95, 269.45, 269.65, 269.75, 269.45, 269.05, 
    268.85, 268.25, 268.45, 269.45, 270.65, 270.85, 271.45, 270.95, 269.85, 
    269.75, 271.35, 271.75, 272.05, 271.85, 271.45, 271.75, 271.75, 271.65, 
    271.55, 271.75, 271.95, 272.15, 272.05, 271.85, 271.75, 271.65, 271.75, 
    271.85, 271.75, 271.35, 271.15, 271.05, 270.85, 270.85, 270.75, 270.55, 
    270.15, 270.15, 269.85, 270.95, 270.75, 270.65, 270.45, 270.45, 269.55, 
    269.65, 270.85, 270.65, 269.95, 270.25, 269.95, 269.65, 269.55, 269.25, 
    269.05, 268.25, 268.45, 268.65, 268.55, 268.85, 268.85, 268.95, 268.75, 
    268.55, 268.75, 268.75, 268.75, 268.75, 268.45, 268.15, 268.15, 268.35, 
    268.25, 268.55, 268.75, 268.65, 268.25, 268.25, 268.05, 267.85, 268.05, 
    267.75, 267.75, 267.75, 267.85, 267.95, 267.55, 267.95, 268.15, 267.85, 
    267.65, 267.65, 267.35, 266.75, 266.65, 266.65, 266.55, 266.45, 266.65, 
    266.35, 265.05, 265.05, 266.35, 267.05, 267.15, 267.45, 267.75, 267.45, 
    266.05, 265.05, 266.25, 266.45, 264.65, 264.75, 264.45, 264.65, 264.95, 
    264.55, 264.35, 263.45, 261.85, 262.85, 261.75, 262.85, 264.15, 262.85, 
    263.05, 263.45, 263.25, 263.65, 262.95, 262.85, 261.65, 263.35, 262.95, 
    262.75, 261.25, 262.95, 262.95, 262.45, 261.55, 261.05, 262.45, 260.75, 
    260.75, 261.75, 262.55, 262.45, 262.95, 263.55, 263.65, 263.65, 263.65, 
    263.45, 263.35, 263.25, 263.15, 263.45, 263.65, 263.55, 263.55, 263.25, 
    264.05, 263.55, 262.95, 262.45, 261.85, 261.35, 260.85, 260.05, 260.25, 
    260.35, 260.15, 260.45, 259.55, 257.95, 258.05, 258.45, 258.35, 258.35, 
    258.55, 258.15, 258.55, 258.65, 258.45, 258.75, 258.85, 259.55, 260.15, 
    260.35, 260.55, 259.75, 259.25, 259.55, 258.95, 259.15, 259.15, 259.25, 
    259.55, 260.15, 260.55, 260.85, 261.05, 261.05, 261.05, 260.85, 260.85, 
    260.75, 260.65, 260.65, 260.55, 261.15, 261.15, 261.25, 260.85, 260.75, 
    260.85, 261.05, 261.25, 261.15, 261.25, 261.15, 261.15, 261.45, 261.35, 
    260.75, 260.65, 260.95, 261.35, 261.35, 261.25, 261.45, 261.75, 261.95, 
    262.05, 261.75, 260.75, 260.55, 259.35, 258.75, 258.35, 258.05, 257.65, 
    257.85, 257.55, 257.15, 256.65, 256.35, 255.75, 256.25, 257.05, 257.85, 
    258.25, 258.15, 258.25, 257.95, 257.55, 258.15, 257.35, 257.25, 257.05, 
    256.75, 256.05, 255.65, 255.45, 255.35, 255.75, 254.15, 255.15, 255.05, 
    254.85, 254.65, 255.05, 255.65, 255.25, 255.25, 255.45, 255.85, 255.45, 
    256.05, 256.85, 257.05, 257.25, 258.25, 257.95, 258.35, 259.25, 258.45, 
    259.85, 259.45, 259.75, 260.15, 260.05, 260.15, 260.15, 260.85, 260.95, 
    261.35, 261.65, 262.45, 262.45, 262.45, 263.25, 264.05, 262.75, 262.55, 
    262.55, 263.35, 263.55, 264.45, 264.45, 264.35, 264.35, 264.45, 263.65, 
    263.55, 263.05, 263.15, 262.85, 262.95, 263.05, 263.25, 263.75, 263.75, 
    264.65, 263.85, 264.25, 264.65, 265.15, 264.75, 264.85, 265.25, 265.55, 
    265.25, 265.05, 264.85, 264.85, 265.65, 266.25, 266.55, 266.85, 267.25, 
    267.45, 267.95, 268.45, 268.65, 269.05, 268.55, 268.85, 268.65, 268.35, 
    267.95, 267.85, 267.85, 267.55, 267.85, 267.75, 267.55, 267.65, 267.65, 
    267.95, 267.75, 267.65, 267.65, 267.65, 267.85, 267.75, 267.85, 268.05, 
    267.95, 268.15, 268.05, 268.25, 268.45, 268.65, 269.05, 269.55, 269.65, 
    269.85, 269.55, 269.45, 269.35, 269.25, 269.65, 269.75, 270.25, 270.55, 
    270.55, 270.45, 270.55, 270.75, 271.15, 271.65, 271.65, 271.85, 271.85, 
    271.75, 272.25, 272.85, 273.15, 271.75, 272.05, 271.95, 272.95, 272.95, 
    273.05, 272.95, 272.75, 273.25, 272.45, 273.15, 272.85, 272.75, 272.65, 
    272.65, 272.55, 272.35, 271.05, 270.15, 269.65, 268.55, 268.05, 267.35, 
    266.85, 265.95, 264.85, 264.05, 263.75, 263.45, 263.65, 263.05, 262.95, 
    262.55, 262.35, 261.85, 261.65, 260.75, 261.35, 261.65, 261.35, 261.35, 
    261.55, 260.95, 261.35, 261.55, 261.55, 261.45, 261.55, 261.55, 261.45, 
    261.75, 261.45, 261.25, 261.15, 261.15, 260.25, 260.15, 259.95, 260.05, 
    260.05, 259.95, 259.55, 259.55, 259.55, 259.85, 259.65, 260.55, 260.45, 
    260.45, 260.75, 260.85, 260.85, 261.45, 260.95, 261.05, 261.25, 261.25, 
    261.35, 261.45, 261.85, 261.45, 261.45, 261.55, 261.85, 261.75, 261.75, 
    261.65, 261.65, 261.75, 261.65, 261.65, 261.35, 260.75, 260.35, 260.65, 
    261.15, 260.55, 261.05, 260.55, 260.95, 261.05, 260.75, 261.35, 259.95, 
    261.05, 259.85, 259.35, 258.85, 259.65, 259.75, 261.05, 261.75, 261.55, 
    262.15, 262.25, 261.85, 261.95, 261.95, 261.25, 261.15, 260.95, 260.05, 
    259.25, 259.45, 259.15, 258.45, 259.15, 259.95, 259.65, 259.25, 260.55, 
    259.95, 258.75, 259.35, 259.25, 259.75, 258.45, 259.55, 259.45, 259.25, 
    259.65, 259.95, 260.55, 260.45, 260.15, 260.25, 260.65, 259.25, 259.45, 
    258.85, 258.65, 258.35, 258.15, 259.95, 261.25, 261.35, 260.95, 260.65, 
    259.85, 259.15, 258.95, 258.65, 259.25, 259.35, 258.75, 259.15, 257.75, 
    258.95, 258.45, 257.95, 258.25, 256.75, 256.95, 256.05, 257.95, 256.25, 
    258.15, 257.75, 257.65, 257.75, 257.45, 257.55, 257.15, 257.25, 256.35, 
    255.75, 255.35, 255.15, 256.65, 256.95, 257.35, 257.95, 258.35, 258.35, 
    258.15, 257.95, 257.45, 257.25, 257.45, 257.35, 257.45, 257.35, 257.25, 
    257.15, 256.95, 256.75, 256.45, 256.55, 257.15, 257.55, 257.95, 258.15, 
    257.95, 257.75, 257.35, 256.95, 256.75, 257.15, 257.05, 257.05, 256.85, 
    256.55, 256.45, 256.35, 256.35, 256.15, 255.95, 256.05, 256.05, 256.15, 
    256.25, 256.25, 256.35, 256.55, 256.45, 256.45, 256.65, 256.35, 256.45, 
    256.35, 256.25, 256.25, 256.15, 256.15, 256.05, 256.05, 256.05, 256.25, 
    255.95, 255.85, 256.15, 256.25, 256.25, 255.85, 255.25, 254.85, 254.15, 
    254.45, 254.15, 253.85, 253.95, 253.85, 254.05, 254.25, 254.45, 254.35, 
    254.05, 253.65, 254.25, 253.75, 253.35, 254.05, 254.35, 253.25, 252.45, 
    252.65, 252.15, 252.95, 253.55, 253.75, 254.85, 255.15, 256.65, 258.35, 
    259.25, 259.05, 259.85, 260.25, 259.55, 258.85, 258.55, 258.45, 257.35, 
    256.95, 256.55, 256.85, 257.25, 255.95, 255.95, 255.45, 255.65, 256.65, 
    257.35, 258.25, 258.65, 258.35, 259.95, 260.95, 261.75, 262.25, 259.75, 
    258.35, 257.45, 256.85, 256.45, 255.25, 255.85, 255.75, 255.45, 256.35, 
    257.15, 257.25, 257.35, 258.05, 258.35, 258.75, 259.05, 259.05, 260.55, 
    260.95, 261.55, 262.05, 259.25, 258.95, 259.95, 260.35, 260.25, 259.55, 
    259.55, 258.95, 258.45, 257.55, 257.65, 257.65, 258.05, 257.85, 257.65, 
    257.45, 257.25, 257.75, 257.65, 257.55, 256.65, 255.95, 255.95, 256.05, 
    255.95, 255.85, 255.95, 256.65, 256.45, 256.55, 256.25, 255.55, 256.05, 
    254.85, 255.75, 255.05, 254.45, 254.25, 252.45, 252.25, 251.85, 251.95, 
    250.75, 251.45, 251.85, 252.05, 253.25, 253.75, 256.05, 254.65, 255.45, 
    256.15, 256.75, 257.45, 256.65, 256.95, 257.45, 257.85, 257.05, 257.55, 
    257.35, 257.55, 258.75, 259.25, 260.45, 260.95, 261.25, 262.05, 262.45, 
    262.15, 262.15, 261.85, 261.85, 261.25, 261.85, 261.65, 260.95, 260.65, 
    260.95, 260.95, 261.35, 259.95, 259.55, 259.25, 258.95, 258.95, 257.15, 
    256.55, 256.75, 257.15, 259.55, 259.95, 260.85, 261.25, 260.95, 260.45, 
    260.65, 260.85, 261.65, 261.15, 261.75, 262.05, 262.45, 262.65, 262.65, 
    263.05, 263.05, 263.45, 263.75, 264.05, 264.85, 265.35, 265.45, 266.25, 
    266.25, 266.35, 266.55, 266.45, 266.35, 266.35, 266.45, 266.15, 265.95, 
    265.75, 265.05, 264.95, 264.65, 263.85, 263.05, 262.55, 262.75, 263.05, 
    263.05, 262.45, 262.15, 261.95, 261.85, 261.75, 261.55, 260.95, 260.05, 
    258.65, 257.95, 257.45, 257.35, 256.85, 256.05, 255.55, 255.05, 254.75, 
    254.85, 254.45, 254.25, 253.95, 253.95, 253.95, 254.05, 253.65, 253.65, 
    253.75, 254.05, 254.35, 254.55, 255.15, 255.25, 253.95, 254.55, 254.05, 
    253.35, 253.65, 252.75, 253.05, 253.05, 254.05, 252.85, 252.25, 251.65, 
    251.85, 250.95, 252.55, 250.95, 251.35, 251.75, 253.25, 253.35, 253.45, 
    253.35, 253.35, 253.35, 252.75, 253.45, 253.65, 252.95, 253.15, 253.05, 
    253.05, 252.35, 251.95, 252.15, 251.55, 251.45, 251.95, 251.15, 251.85, 
    250.45, 250.35, 249.55, 249.35, 248.65, 249.35, 249.55, 250.75, 250.85, 
    252.05, 253.35, 253.35, 253.85, 254.25, 254.05, 254.65, 254.15, 255.85, 
    256.25, 256.65, 256.75, 256.95, 257.15, 257.05, 257.25, 257.25, 257.55, 
    257.25, 256.65, 255.15, 253.75, 250.85, 251.65, 252.55, 253.55, 254.55, 
    255.85, 258.05, 257.95, 256.95, 256.65, 255.75, 256.25, 254.25, 253.95, 
    253.55, 253.15, 252.85, 253.75, 254.15, 255.95, 256.55, 255.05, 252.55, 
    252.05, 251.15, 251.65, 251.25, 251.25, 251.55, 252.35, 251.55, 251.75, 
    253.15, 253.55, 252.95, 253.45, 253.65, 253.95, 254.05, 254.05, 254.65, 
    254.95, 256.05, 255.15, 255.25, 254.65, 254.45, 254.85, 254.55, 254.65, 
    255.15, 255.25, 255.95, 255.65, 256.15, 256.35, 256.45, 256.45, 256.05, 
    255.25, 254.75, 253.75, 253.35, 252.95, 253.05, 252.95, 253.45, 253.75, 
    254.05, 254.25, 254.25, 255.05, 255.35, 255.55, 256.05, 256.95, 257.45, 
    257.55, 258.05, 258.65, 259.35, 259.65, 260.55, 260.65, 260.55, 260.45, 
    259.05, 258.05, 258.15, 257.25, 257.05, 256.95, 257.35, 257.75, 258.05, 
    258.35, 258.55, 258.95, 259.15, 259.45, 259.65, 259.65, 260.15, 260.65, 
    260.25, 259.75, 258.85, 258.15, 257.45, 257.35, 257.95, 257.85, 257.95, 
    258.15, 258.05, 258.05, 258.55, 258.65, 258.55, 258.75, 258.95, 259.15, 
    259.35, 259.55, 260.15, 260.45, 260.55, 260.75, 260.65, 260.75, 260.45, 
    260.15, 260.05, 260.05, 260.25, 260.35, 260.45, 260.55, 260.65, 260.35, 
    259.45, 259.05, 259.25, 259.15, 258.95, 258.75, 258.95, 259.15, 259.05, 
    259.65, 259.55, 259.75, 259.35, 259.35, 258.85, 258.65, 258.75, 259.15, 
    258.35, 257.65, 258.45, 258.65, 256.25, 258.75, 258.45, 258.05, 258.25, 
    257.85, 257.05, 258.15, 258.65, 258.85, 258.95, 258.95, 258.85, 258.75, 
    258.75, 258.65, 258.95, 259.05, 258.55, 258.25, 258.15, 258.35, 258.65, 
    257.75, 257.15, 256.95, 256.85, 256.85, 256.95, 257.25, 257.65, 257.75, 
    257.45, 257.35, 257.15, 256.95, 256.95, 257.35, 257.65, 257.85, 257.15, 
    257.25, 252.55, 255.65, 255.65, 255.25, 255.65, 255.75, 255.45, 255.35, 
    255.35, 253.85, 252.15, 257.15, 254.45, 254.85, 254.95, 255.05, 255.65, 
    256.15, 256.25, 256.25, 257.65, 255.95, 256.05, 257.05, 256.25, 256.15, 
    254.55, 253.65, 253.85, 254.25, 254.85, 254.05, 254.55, 253.85, 254.05, 
    254.25, 254.95, 255.65, 255.85, 255.75, 255.85, 255.75, 256.05, 256.65, 
    256.45, 257.15, 257.45, 256.65, 256.05, 256.35, 255.55, 254.85, 255.05, 
    254.85, 255.45, 255.85, 255.85, 255.05, 254.95, 255.35, 254.95, 255.45, 
    256.45, 256.85, 257.15, 257.85, 257.25, 257.75, 257.65, 256.65, 256.55, 
    256.15, 255.55, 255.95, 255.45, 255.35, 254.85, 254.95, 254.85, 254.45, 
    255.55, 254.35, 254.55, 255.55, 254.95, 254.65, 255.65, 256.45, 256.25, 
    256.45, 256.55, 256.15, 256.05, 256.55, 255.45, 256.05, 256.45, 257.55, 
    256.35, 255.35, 256.05, 255.25, 254.55, 254.55, 255.35, 255.85, 252.85, 
    255.25, 256.25, 256.15, 256.55, 256.25, 255.45, 255.75, 256.15, 254.95, 
    255.35, 254.85, 254.85, 254.55, 253.55, 253.05, 252.95, 253.35, 253.15, 
    253.05, 252.55, 252.65, 252.55, 252.45, 252.65, 253.15, 253.75, 253.55, 
    253.35, 254.65, 253.75, 254.25, 254.75, 254.05, 254.05, 254.25, 253.85, 
    253.05, 252.75, 252.85, 252.95, 252.15, 251.95, 252.85, 252.35, 252.65, 
    252.85, 252.75, 252.95, 254.05, 253.95, 256.15, 254.95, 255.35, 255.45, 
    255.35, 255.65, 254.65, 255.65, 254.65, 254.75, 254.95, 254.25, 253.25, 
    252.95, 254.15, 253.25, 252.95, 252.75, 251.95, 251.75, 252.05, 252.15, 
    252.85, 252.35, 252.95, 253.05, 254.95, 255.55, 255.65, 255.85, 255.95, 
    255.95, 255.25, 255.15, 254.55, 254.55, 253.75, 254.15, 253.95, 253.75, 
    253.15, 254.05, 255.05, 256.35, 256.85, 257.15, 257.55, 258.75, 259.45, 
    260.45, 261.65, 264.35, 263.05, 261.85, 262.35, 261.85, 261.45, 260.95, 
    260.65, 260.25, 259.95, 260.05, 260.35, 259.95, 260.15, 260.45, 260.35, 
    260.45, 261.85, 262.45, 263.05, 262.95, 263.05, 265.45, 264.35, 264.05, 
    264.45, 264.65, 263.65, 263.45, 263.65, 263.45, 263.85, 263.05, 264.05, 
    264.85, 264.45, 265.55, 266.05, 266.85, 267.15, 267.15, 267.55, 267.75, 
    268.15, 267.25, 267.55, 266.15, 265.95, 265.15, 265.85, 263.75, 262.35, 
    261.45, 261.25, 260.35, 260.75, 260.35, 259.85, 259.15, 258.95, 259.15, 
    258.85, 259.25, 259.45, 259.35, 259.35, 259.15, 259.95, 261.45, 260.85, 
    260.35, 260.95, 261.05, 260.95, 260.85, 260.15, 260.95, 260.35, 260.85, 
    260.75, 261.45, 260.55, 261.15, 262.25, 261.95, 262.85, 262.95, 263.45, 
    263.65, 264.05, 263.95, 264.15, 264.45, 264.85, 265.45, 266.15, 265.95, 
    266.95, 267.55, 267.85, 268.05, 267.85, 267.65, 267.65, 267.35, 267.65, 
    268.15, 268.25, 268.55, 268.95, 268.95, 268.75, 268.75, 268.15, 267.05, 
    266.75, 265.95, 265.85, 265.95, 266.25, 266.15, 266.15, 266.25, 265.95, 
    266.65, 265.25, 264.45, 263.75, 262.95, 262.55, 261.85, 261.25, 260.65, 
    260.05, 259.65, 259.15, 259.45, 259.45, 259.15, 259.75, 259.75, 259.95, 
    260.45, 260.55, 260.55, 260.75, 260.75, 260.65, 260.45, 259.65, 259.35, 
    258.45, 259.05, 258.95, 258.85, 259.65, 260.35, 260.45, 259.65, 258.45, 
    257.75, 257.65, 257.15, 257.75, 259.65, 259.05, 262.05, 260.35, 260.65, 
    260.35, 260.55, 260.45, 259.15, 258.75, 258.05, 258.35, 258.75, 258.95, 
    259.65, 259.65, 259.05, 259.65, 260.15, 260.95, 261.15, 261.35, 261.65, 
    262.25, 262.55, 262.85, 263.05, 263.45, 264.15, 264.65, 265.05, 265.45, 
    265.75, 266.15, 266.35, 266.45, 266.45, 266.45, 266.25, 266.05, 266.65, 
    267.15, 268.05, 267.35, 267.85, 268.65, 268.45, 267.95, 267.55, 266.75, 
    265.95, 265.25, 264.85, 264.65, 264.55, 264.85, 265.95, 264.15, 262.95, 
    260.35, 259.75, 259.55, 259.25, 259.35, 260.65, 260.45, 260.25, 260.35, 
    260.35, 260.75, 261.15, 261.15, 261.65, 261.65, 261.35, 261.15, 261.55, 
    261.75, 261.75, 261.85, 261.95, 261.95, 262.15, 262.35, 262.65, 262.85, 
    263.05, 262.55, 262.05, 261.45, 261.15, 261.85, 261.55, 261.55, 261.65, 
    261.85, 261.95, 262.05, 262.45, 263.05, 263.35, 263.05, 263.55, 263.55, 
    263.35, 263.15, 263.05, 263.25, 263.35, 263.25, 262.95, 262.45, 262.85, 
    262.65, 261.95, 261.55, 261.15, 261.05, 260.45, 259.65, 258.95, 260.75, 
    261.15, 261.35, 261.15, 261.45, 261.35, 261.55, 261.45, 261.05, 260.05, 
    259.75, 259.25, 258.25, 258.45, 259.25, 258.15, 258.45, 258.45, 259.85, 
    260.45, 260.85, 261.85, 262.35, 262.15, 262.15, 262.05, 262.15, 261.65, 
    261.35, 261.65, 261.65, 261.75, 261.95, 261.75, 261.95, 261.55, 261.45, 
    261.45, 261.35, 261.25, 261.55, 261.65, 261.65, 261.65, 261.45, 261.85, 
    261.75, 261.65, 261.65, 260.95, 260.95, 261.05, 261.25, 261.15, 261.05, 
    261.35, 261.75, 262.05, 262.15, 262.35, 262.65, 262.75, 262.85, 262.35, 
    261.15, 258.95, 257.55, 257.05, 256.65, 256.55, 256.85, 257.15, 256.85, 
    257.85, 259.05, 259.35, 259.05, 259.25, 259.05, 259.45, 259.05, 258.15, 
    256.95, 256.55, 255.15, 255.35, 255.85, 255.25, 255.25, 254.95, 255.75, 
    256.05, 256.15, 256.35, 257.65, 258.15, 257.95, 259.85, 258.35, 257.95, 
    257.15, 257.55, 257.45, 257.05, 256.65, 256.85, 256.45, 256.45, 255.45, 
    255.95, 254.85, 253.85, 254.05, 253.05, 252.85, 253.65, 254.05, 254.25, 
    255.35, 255.65, 255.75, 256.35, 256.55, 256.55, 256.95, 256.75, 256.65, 
    257.05, 256.95, 257.15, 256.95, 257.25, 256.85, 256.65, 256.45, 255.95, 
    256.15, 256.15, 256.45, 256.55, 256.75, 257.25, 258.05, 258.75, 258.95, 
    259.55, 259.85, 260.15, 260.15, 260.25, 260.05, 259.75, 260.45, 258.05, 
    258.15, 257.95, 258.65, 258.15, 256.95, 255.85, 256.55, 258.35, 257.95, 
    258.45, 258.55, 257.85, 259.35, 260.95, 259.95, 260.85, 262.15, 261.65, 
    263.15, 262.75, 262.05, 261.85, 261.55, 261.35, 261.55, 260.65, 260.45, 
    260.45, 260.15, 259.85, 259.65, 259.65, 259.55, 259.45, 258.95, 258.55, 
    257.95, 258.75, 259.15, 259.85, 260.65, 261.05, 261.25, 261.15, 261.45, 
    261.55, 261.75, 261.65, 261.95, 261.55, 261.65, 262.15, 262.25, 261.95, 
    262.95, 263.35, 264.15, 264.15, 264.65, 265.15, 265.55, 266.15, 267.05, 
    266.75, 266.65, 268.15, 268.35, 269.75, 266.65, 266.55, 265.75, 264.55, 
    264.35, 264.65, 264.85, 264.55, 264.25, 264.55, 264.45, 262.45, 262.95, 
    263.55, 261.15, 260.95, 259.35, 258.85, 260.05, 259.85, 257.65, 257.65, 
    257.85, 257.85, 258.15, 258.15, 258.25, 258.65, 258.55, 257.95, 257.75, 
    258.55, 258.55, 258.75, 259.05, 258.25, 258.35, 258.55, 258.75, 258.45, 
    258.05, 257.75, 257.85, 257.95, 258.15, 258.35, 258.35, 258.55, 258.75, 
    258.15, 258.15, 258.05, 257.45, 257.95, 257.85, 256.95, 256.45, 258.75, 
    259.05, 259.95, 260.55, 260.45, 261.25, 261.65, 261.55, 262.25, 262.55, 
    264.05, 264.25, 264.95, 265.75, 266.05, 266.35, 266.25, 266.25, 266.55, 
    266.75, 266.95, 266.95, 265.85, 265.25, 265.05, 265.25, 265.55, 266.35, 
    267.05, 267.15, 267.35, 267.85, 268.55, 269.15, 269.15, 269.65, 270.35, 
    270.75, 270.75, 271.05, 271.15, 270.85, 270.95, 271.35, 271.45, 271.95, 
    271.85, 271.75, 271.45, 271.25, 270.85, 270.95, 270.65, 270.45, 270.15, 
    270.35, 270.45, 270.85, 271.05, 271.45, 271.75, 272.05, 272.45, 272.95, 
    273.15, 273.35, 273.35, 273.55, 273.75, 273.55, 273.35, 273.15, 273.05, 
    272.85, 272.65, 273.05, 273.25, 273.05, 273.15, 273.25, 273.55, 274.05, 
    274.15, 273.65, 273.25, 272.95, 272.95, 272.65, 272.85, 272.85, 273.05, 
    273.25, 273.15, 273.55, 273.45, 273.35, 273.45, 273.65, 273.45, 273.45, 
    273.35, 273.35, 273.35, 273.35, 273.35, 273.45, 273.35, 273.45, 273.45, 
    273.45, 273.55, 273.45, 273.65, 273.35, 273.15, 272.95, 272.95, 272.85, 
    272.85, 272.65, 272.65, 272.55, 272.45, 272.55, 272.65, 272.75, 272.85, 
    273.05, 273.15, 273.25, 274.15, 272.95, 272.65, 272.65, 272.65, 272.65, 
    272.25, 271.95, 271.95, 272.45, 271.95, 270.65, 270.65, 271.45, 271.25, 
    271.75, 270.35, 270.95, 271.75, 272.15, 272.35, 272.25, 272.85, 272.65, 
    272.55, 272.65, 272.75, 272.75, 273.25, 273.55, 273.35, 273.55, 272.95, 
    273.35, 273.15, 273.15, 272.75, 272.45, 272.85, 272.35, 272.15, 271.95, 
    272.15, 271.95, 271.95, 272.25, 273.05, 273.45, 272.95, 273.05, 273.65, 
    274.45, 274.35, 273.35, 272.75, 272.55, 271.65, 270.95, 271.05, 271.25, 
    271.05, 270.75, 270.35, 270.15, 270.05, 270.05, 270.15, 270.35, 270.35, 
    270.65, 270.95, 270.95, 271.25, 271.15, 271.25, 271.25, 271.35, 271.45, 
    271.65, 271.75, 271.85, 271.95, 272.05, 272.15, 272.25, 271.95, 271.95, 
    271.95, 271.75, 271.45, 271.75, 271.85, 271.85, 271.85, 272.15, 272.35, 
    272.85, 272.75, 273.45, 273.75, 273.65, 271.95, 272.65, 272.25, 271.75, 
    271.75, 271.35, 271.15, 271.05, 270.75, 270.85, 271.25, 271.35, 271.45, 
    271.25, 271.25, 271.35, 271.15, 270.85, 270.75, 270.65, 270.75, 270.65, 
    270.75, 270.75, 270.85, 270.95, 270.95, 270.85, 270.75, 270.85, 270.15, 
    270.55, 270.45, 270.05, 270.05, 269.75, 269.55, 269.55, 269.15, 269.15, 
    269.05, 269.45, 269.45, 268.85, 268.75, 268.75, 268.95, 269.15, 269.25, 
    269.25, 269.35, 269.35, 269.55, 269.65, 269.55, 269.75, 269.65, 269.75, 
    269.65, 269.75, 269.85, 269.55, 268.75, 268.85, 268.15, 268.55, 268.95, 
    268.55, 269.05, 268.85, 268.95, 269.25, 269.45, 268.85, 268.45, 268.25, 
    268.05, 267.95, 268.05, 267.85, 267.25, 267.45, 267.55, 268.25, 268.55, 
    268.85, 269.45, 269.45, 269.75, 269.85, 270.25, 270.45, 270.65, 270.75, 
    270.85, 271.25, 271.05, 270.85, 270.85, 270.75, 270.95, 270.55, 270.55, 
    270.35, 270.15, 269.95, 269.85, 269.65, 269.65, 269.65, 269.85, 270.05, 
    269.75, 269.75, 269.75, 269.85, 269.95, 270.15, 270.45, 270.15, 270.35, 
    270.25, 270.15, 270.05, 270.05, 270.05, 270.25, 270.25, 269.95, 269.75, 
    269.75, 269.65, 269.55, 269.55, 269.65, 269.85, 269.65, 269.75, 270.05, 
    270.05, 269.75, 269.75, 269.45, 269.25, 269.05, 269.05, 269.25, 269.45, 
    269.55, 269.75, 269.95, 270.25, 270.55, 270.95, 271.25, 271.45, 271.55, 
    271.75, 271.85, 271.95, 272.05, 272.35, 272.45, 272.65, 272.65, 272.65, 
    272.75, 272.85, 273.25, 272.95, 272.55, 272.15, 272.25, 272.55, 272.75, 
    272.85, 272.75, 272.65, 272.55, 272.25, 272.05, 272.05, 271.95, 272.15, 
    272.55, 272.65, 272.35, 272.55, 272.55, 272.65, 272.85, 272.45, 272.25, 
    271.85, 271.75, 271.75, 271.85, 271.75, 271.85, 271.95, 271.95, 271.75, 
    271.55, 271.45, 271.55, 271.75, 271.75, 271.55, 271.55, 271.95, 271.85, 
    271.95, 271.75, 271.45, 271.85, 271.35, 271.15, 270.85, 270.95, 270.85, 
    270.65, 270.45, 270.35, 270.35, 270.35, 270.25, 270.15, 270.15, 270.15, 
    269.75, 269.85, 269.85, 270.15, 270.15, 269.65, 269.35, 269.05, 268.75, 
    268.65, 268.75, 268.55, 268.75, 268.55, 268.45, 268.35, 268.25, 268.95, 
    268.45, 268.35, 268.25, 268.35, 268.35, 269.15, 269.05, 269.05, 268.85, 
    268.95, 268.95, 269.15, 269.25, 269.95, 270.65, 270.95, 270.55, 270.55, 
    270.55, 270.45, 270.25, 270.15, 270.05, 269.95, 269.85, 269.85, 269.95, 
    270.05, 270.15, 269.95, 269.75, 270.15, 270.45, 270.65, 270.75, 270.75, 
    270.75, 270.75, 271.35, 271.55, 271.35, 271.05, 270.15, 270.25, 270.35, 
    270.45, 270.25, 270.05, 270.15, 270.15, 270.15, 270.15, 270.15, 270.05, 
    269.65, 269.75, 270.05, 270.45, 270.55, 270.65, 270.65, 270.95, 271.35, 
    271.25, 271.35, 271.95, 271.85, 271.95, 271.95, 271.95, 272.15, 272.75, 
    273.35, 272.85, 273.35, 273.25, 273.75, 273.85, 274.05, 274.15, 274.45, 
    274.55, 273.15, 272.05, 271.95, 271.45, 271.35, 271.25, 270.95, 271.25, 
    270.95, 271.15, 271.15, 270.95, 270.75, 270.65, 270.45, 270.25, 270.15, 
    270.05, 269.95, 270.05, 270.05, 270.15, 270.25, 270.45, 270.45, 270.55, 
    270.25, 270.05, 270.25, 270.05, 269.85, 269.85, 270.05, 270.55, 270.35, 
    270.75, 270.55, 270.55, 270.45, 270.05, 270.25, 269.95, 270.15, 270.35, 
    270.25, 270.25, 270.25, 270.35, 270.65, 270.75, 270.55, 271.15, 271.05, 
    271.35, 271.85, 272.25, 272.25, 272.15, 272.05, 272.05, 271.95, 270.95, 
    270.85, 270.85, 269.85, 271.55, 271.35, 271.75, 271.95, 271.25, 271.15, 
    271.45, 271.55, 272.15, 272.15, 272.25, 272.15, 272.45, 272.15, 272.15, 
    272.05, 271.55, 271.15, 270.85, 270.55, 270.15, 269.65, 269.75, 269.55, 
    270.15, 269.45, 269.35, 269.05, 269.35, 269.45, 269.75, 269.65, 269.85, 
    270.15, 270.15, 270.15, 270.35, 269.95, 270.75, 269.55, 269.35, 270.15, 
    269.25, 269.45, 268.85, 269.25, 268.65, 268.85, 268.75, 269.25, 269.25, 
    269.15, 269.15, 269.95, 270.25, 271.15, 270.15, 270.75, 270.75, 272.05, 
    271.85, 271.15, 271.05, 271.15, 271.65, 271.45, 271.65, 271.25, 271.25, 
    271.15, 271.05, 271.15, 271.15, 271.25, 271.45, 271.15, 271.15, 271.45, 
    271.75, 271.05, 271.25, 271.15, 271.45, 271.75, 271.75, 271.45, 271.45, 
    271.15, 270.95, 270.95, 270.85, 270.85, 270.85, 270.85, 271.05, 271.05, 
    271.25, 271.25, 271.35, 271.55, 271.55, 271.55, 271.65, 271.75, 271.85, 
    272.15, 272.25, 272.15, 271.85, 271.75, 271.85, 271.95, 272.35, 272.45, 
    272.75, 272.75, 272.65, 272.55, 272.45, 272.15, 272.05, 272.25, 272.25, 
    272.15, 272.15, 272.15, 272.25, 272.25, 272.25, 272.15, 272.05, 272.05, 
    271.95, 271.85, 271.75, 271.65, 271.75, 271.55, 271.25, 271.05, 270.85, 
    270.95, 271.25, 271.55, 272.15, 272.45, 272.35, 272.45, 272.35, 272.35, 
    272.45, 272.55, 272.65, 272.45, 272.65, 272.45, 272.35, 272.45, 272.35, 
    272.75, 272.65, 272.65, 272.75, 272.55, 272.25, 272.15, 272.25, 272.15, 
    272.05, 271.95, 271.95, 271.95, 271.75, 271.95, 271.55, 272.25, 271.75, 
    271.35, 271.15, 270.95, 271.05, 270.35, 270.15, 270.55, 270.95, 270.75, 
    270.35, 270.25, 270.05, 269.85, 269.95, 270.05, 270.15, 270.25, 269.85, 
    269.65, 269.95, 270.05, 269.45, 269.85, 270.35, 270.35, 269.95, 269.75, 
    269.75, 269.95, 269.85, 270.15, 270.35, 270.65, 270.55, 270.45, 270.65, 
    270.85, 271.15, 271.25, 271.25, 271.15, 271.25, 271.35, 271.35, 271.35, 
    271.35, 271.55, 271.75, 272.05, 271.95, 271.95, 271.95, 272.05, 272.15, 
    272.75, 272.65, 272.35, 272.25, 272.25, 272.05, 271.95, 271.85, 271.95, 
    271.55, 271.55, 271.35, 271.55, 271.75, 271.85, 272.15, 272.15, 272.25, 
    272.15, 272.15, 272.05, 272.05, 271.65, 271.45, 271.35, 271.55, 271.65, 
    271.75, 271.65, 271.65, 271.65, 271.75, 271.65, 271.45, 271.45, 271.45, 
    271.35, 271.45, 271.35, 271.45, 271.45, 271.65, 271.75, 271.85, 271.95, 
    271.85, 271.85, 271.75, 271.75, 271.85, 271.85, 271.85, 271.85, 271.55, 
    271.65, 271.65, 271.85, 271.85, 271.95, 271.75, 271.85, 271.95, 272.05, 
    271.75, 272.25, 272.05, 272.05, 271.95, 271.85, 271.95, 271.55, 271.75, 
    271.75, 271.65, 271.45, 271.45, 271.35, 271.25, 271.25, 271.25, 271.05, 
    271.35, 271.25, 271.15, 270.85, 270.65, 270.85, 270.85, 270.75, 270.85, 
    270.65, 270.55, 270.15, 270.15, 270.45, 270.45, 270.65, 270.65, 271.05, 
    270.95, 270.65, 270.65, 270.15, 270.35, 270.35, 270.05, 270.15, 269.95, 
    270.25, 270.15, 270.35, 270.35, 270.25, 270.15, 270.05, 270.05, 269.95, 
    270.05, 270.05, 270.25, 270.55, 270.55, 270.55, 270.55, 270.55, 270.55, 
    270.65, 270.65, 270.75, 270.85, 271.15, 271.55, 271.45, 271.85, 272.65, 
    270.95, 271.75, 273.05, 272.65, 272.35, 272.05, 272.05, 271.75, 271.85, 
    271.85, 271.75, 271.75, 272.05, 271.95, 271.75, 273.15, 271.95, 272.85, 
    273.15, 273.55, 273.65, 272.65, 273.15, 273.35, 273.25, 274.25, 274.55, 
    273.85, 273.85, 273.45, 273.45, 273.75, 273.35, 273.35, 273.15, 272.85, 
    272.65, 272.55, 273.05, 272.65, 272.75, 272.85, 272.15, 272.05, 272.05, 
    272.15, 272.15, 272.25, 272.35, 272.45, 272.65, 272.55, 272.65, 272.95, 
    272.95, 273.05, 272.95, 271.75, 271.75, 272.05, 272.85, 273.35, 273.35, 
    273.05, 272.75, 272.85, 272.45, 272.45, 271.85, 271.15, 271.05, 271.35, 
    271.15, 271.55, 272.25, 273.05, 273.65, 273.95, 273.35, 273.95, 274.95, 
    274.15, 274.65, 272.75, 274.65, 274.85, 274.75, 274.45, 274.35, 274.75, 
    274.55, 273.85, 274.15, 273.65, 273.85, 273.55, 274.05, 273.95, 273.75, 
    273.65, 273.55, 273.55, 274.45, 274.35, 274.05, 274.05, 273.95, 273.65, 
    273.55, 273.45, 273.15, 273.05, 273.15, 273.15, 273.35, 273.55, 274.45, 
    274.55, 274.55, 274.35, 275.75, 275.25, 275.15, 275.15, 274.75, 274.35, 
    274.05, 274.05, 273.95, 273.85, 273.45, 273.15, 272.95, 273.05, 273.05, 
    273.15, 273.15, 273.25, 273.85, 273.35, 273.75, 273.75, 273.15, 273.75, 
    275.25, 274.65, 275.55, 274.75, 274.55, 274.15, 273.75, 274.05, 273.95, 
    274.55, 275.25, 274.95, 274.15, 274.65, 274.85, 275.05, 275.15, 274.75, 
    274.35, 274.25, 274.45, 274.35, 274.95, 275.05, 274.85, 274.25, 274.45, 
    274.85, 275.15, 275.25, 274.95, 275.05, 274.95, 274.55, 274.35, 274.15, 
    273.75, 273.65, 273.25, 273.05, 273.15, 273.15, 273.15, 273.45, 273.55, 
    273.75, 273.95, 273.95, 273.95, 273.95, 274.35, 274.05, 274.85, 274.45, 
    274.45, 274.05, 274.05, 273.75, 273.35, 273.15, 273.25, 273.25, 273.55, 
    273.75, 274.15, 274.15, 273.75, 274.15, 273.95, 274.05, 273.95, 273.65, 
    273.85, 273.45, 274.85, 276.45, 274.05, 274.35, 274.75, 274.55, 274.15, 
    274.25, 274.35, 273.85, 273.65, 274.15, 274.05, 274.05, 273.75, 273.85, 
    274.25, 273.65, 273.05, 273.45, 273.45, 273.45, 273.55, 273.95, 273.45, 
    273.95, 274.55, 275.05, 274.45, 274.75, 275.25, 275.85, 275.35, 274.55, 
    274.75, 274.65, 274.45, 274.45, 274.35, 274.15, 273.95, 274.25, 274.65, 
    273.85, 273.55, 273.55, 274.05, 272.85, 272.05, 272.05, 272.35, 271.35, 
    271.85, 272.45, 273.55, 276.05, 274.55, 278.25, 278.85, 273.55, 274.45, 
    273.55, 273.95, 272.45, 273.85, 272.15, 274.55, 273.35, 273.55, 273.75, 
    273.15, 278.15, 275.75, 274.35, 274.35, 274.25, 274.25, 274.65, 274.55, 
    274.65, 274.55, 274.45, 275.05, 274.65, 274.35, 274.65, 274.15, 275.45, 
    276.75, 275.25, 275.75, 273.95, 276.75, 274.45, 275.05, 275.15, 275.15, 
    275.25, 275.35, 274.05, 275.45, 274.75, 274.45, 275.25, 274.05, 274.05, 
    274.25, 274.45, 272.95, 273.75, 274.45, 273.95, 273.25, 273.35, 273.35, 
    273.25, 273.35, 273.55, 273.85, 274.05, 273.95, 274.25, 274.35, 274.45, 
    274.25, 274.25, 274.35, 274.85, 275.25, 275.25, 275.35, 275.35, 275.05, 
    274.35, 275.25, 274.55, 274.65, 273.55, 273.65, 273.55, 273.45, 273.55, 
    273.65, 273.45, 273.55, 274.05, 273.55, 273.35, 273.35, 273.35, 273.35, 
    273.15, 273.15, 273.15, 273.15, 273.15, 273.15, 273.05, 273.15, 273.15, 
    273.05, 273.05, 273.05, 273.05, 273.05, 272.95, 272.95, 272.95, 272.95, 
    272.95, 273.05, 273.05, 272.95, 272.95, 273.05, 273.05, 273.05, 273.05, 
    272.95, 272.95, 272.85, 272.95, 272.95, 272.95, 272.95, 273.05, 272.95, 
    272.85, 272.85, 272.95, 272.95, 272.95, 272.95, 272.95, 273.05, 273.05, 
    273.05, 272.95, 272.95, 273.05, 273.05, 273.05, 272.95, 272.95, 272.85, 
    272.85, 272.85, 272.85, 272.85, 272.85, 272.95, 272.95, 272.85, 272.85, 
    272.75, 272.75, 272.75, 272.95, 272.95, 273.15, 273.15, 273.25, 273.25, 
    273.15, 273.25, 273.15, 273.15, 273.15, 272.95, 273.15, 273.05, 273.15, 
    273.15, 273.45, 273.65, 273.95, 273.85, 273.75, 274.05, 274.05, 274.25, 
    274.45, 274.25, 274.15, 274.05, 273.95, 273.65, 273.35, 273.35, 273.35, 
    273.15, 272.85, 272.85, 273.05, 273.15, 272.65, 272.85, 272.95, 272.95, 
    272.85, 272.85, 272.95, 272.95, 273.15, 273.05, 272.75, 272.85, 272.95, 
    272.85, 273.25, 273.55, 273.65, 273.45, 273.35, 273.35, 273.15, 273.05, 
    273.15, 272.75, 272.75, 272.85, 272.65, 272.45, 272.55, 272.65, 272.65, 
    272.45, 272.65, 272.75, 272.85, 272.85, 272.75, 272.85, 272.75, 272.85, 
    272.85, 272.75, 272.75, 272.75, 272.85, 272.75, 272.55, 272.45, 272.85, 
    272.85, 273.05, 273.25, 273.15, 273.65, 274.35, 274.95, 275.15, 275.25, 
    275.45, 275.55, 275.45, 274.75, 273.45, 272.95, 272.35, 272.35, 272.45, 
    272.25, 272.25, 272.45, 273.25, 273.45, 273.15, 273.25, 273.55, 273.85, 
    274.05, 274.35, 274.05, 274.75, 275.45, 274.85, 274.65, 275.25, 275.85, 
    275.55, 275.45, 275.55, 275.75, 276.35, 276.25, 276.25, 276.05, 276.65, 
    276.45, 276.65, 276.45, 275.95, 276.95, 276.75, 277.05, 277.55, 276.15, 
    275.85, 277.65, 275.65, 275.85, 275.85, 276.55, 277.15, 276.85, 279.15, 
    278.85, 277.95, 277.15, 278.35, 277.35, 276.55, 276.15, 275.45, 274.95, 
    274.35, 275.55, 275.45, 275.25, 275.45, 275.35, 274.75, 274.45, 274.25, 
    274.25, 274.85, 276.05, 275.35, 275.65, 275.55, 275.25, 274.85, 274.75, 
    274.95, 274.75, 275.65, 276.05, 275.65, 275.65, 275.75, 276.15, 276.75, 
    276.25, 276.45, 275.65, 275.55, 275.25, 275.55, 275.65, 275.65, 275.35, 
    275.35, 275.45, 275.45, 275.65, 275.45, 275.15, 274.85, 275.05, 274.95, 
    274.95, 274.85, 274.75, 274.65, 274.95, 274.85, 275.05, 275.15, 275.55, 
    275.55, 276.05, 275.85, 275.45, 275.55, 275.55, 276.05, 277.05, 276.15, 
    275.45, 275.75, 276.45, 278.05, 276.45, 276.45, 276.85, 275.95, 275.65, 
    275.25, 275.25, 275.55, 275.65, 275.35, 275.35, 276.05, 276.45, 276.15, 
    276.65, 276.55, 276.15, 275.75, 276.35, 276.95, 277.05, 276.85, 276.05, 
    275.75, 276.25, 276.35, 276.35, 276.15, 275.65, 276.15, 276.45, 276.15, 
    276.85, 276.55, 277.55, 276.25, 277.45, 277.15, 276.95, 276.85, 277.35, 
    276.45, 276.85, 278.15, 278.75, 278.35, 276.75, 277.05, 276.65, 277.45, 
    276.95, 276.05, 277.15, 278.15, 277.55, 277.75, 277.45, 277.15, 277.15, 
    277.35, 277.25, 277.05, 277.05, 277.05, 276.35, 276.05, 276.85, 277.25, 
    277.25, 276.45, 276.45, 275.95, 275.45, 274.95, 275.05, 275.15, 274.95, 
    274.55, 274.85, 275.25, 275.75, 276.45, 276.45, 276.35, 275.75, 275.95, 
    276.85, 276.15, 275.35, 275.15, 275.35, 275.45, 275.35, 275.35, 275.75, 
    274.95, 275.25, 275.15, 275.35, 274.95, 274.95, 275.45, 275.95, 276.15, 
    275.95, 276.75, 276.25, 276.05, 275.85, 275.85, 275.35, 275.35, 275.35, 
    275.15, 275.15, 275.35, 275.45, 276.15, 275.05, 274.95, 274.25, 274.65, 
    275.05, 275.05, 274.65, 273.45, 272.95, 272.65, 272.45, 272.85, 272.75, 
    273.95, 274.45, 275.05, 274.65, 276.25, 277.55, 276.55, 276.15, 275.55, 
    276.35, 276.15, 275.85, 275.85, 275.35, 274.55, 273.95, 273.95, 274.75, 
    274.95, 275.05, 275.15, 275.25, 275.55, 276.15, 275.45, 275.35, 275.55, 
    275.75, 275.55, 275.05, 275.05, 274.95, 274.85, 274.35, 274.55, 274.55, 
    274.35, 273.25, 273.15, 273.35, 273.25, 273.35, 273.75, 273.75, 273.75, 
    273.65, 273.25, 273.35, 273.35, 273.85, 273.85, 273.85, 273.85, 274.05, 
    273.95, 274.65, 275.05, 275.15, 274.85, 274.75, 274.85, 274.75, 274.95, 
    274.05, 275.15, 275.25, 275.15, 275.25, 272.55, 272.65, 275.15, 275.45, 
    275.35, 275.85, 276.15, 276.25, 276.45, 275.55, 275.85, 273.95, 274.85, 
    275.35, 274.85, 274.65, 275.05, 275.25, 275.25, 275.05, 275.05, 274.95, 
    275.05, 275.15, 275.25, 275.15, 275.25, 275.65, 275.45, 275.85, 275.85, 
    276.05, 276.45, 276.45, 277.85, 278.35, 278.35, 278.25, 277.85, 277.35, 
    276.95, 276.85, 275.85, 276.35, 276.15, 276.05, 276.05, 276.55, 277.35, 
    277.15, 276.55, 276.35, 275.65, 276.05, 276.45, 276.35, 276.05, 276.15, 
    276.35, 276.65, 276.75, 276.85, 276.65, 276.55, 276.55, 276.55, 276.45, 
    276.65, 276.65, 276.45, 276.05, 276.15, 276.05, 276.45, 276.25, 276.25, 
    276.15, 275.85, 275.05, 275.35, 275.25, 275.15, 275.65, 276.85, 276.15, 
    276.45, 276.25, 275.65, 275.45, 275.75, 276.15, 275.85, 276.05, 274.45, 
    273.45, 274.05, 273.65, 273.75, 273.95, 273.55, 273.35, 273.95, 274.05, 
    274.15, 276.65, 276.05, 276.75, 275.05, 276.45, 276.95, 277.35, 275.85, 
    276.15, 275.45, 275.05, 275.35, 275.15, 275.25, 275.85, 277.15, 275.95, 
    276.35, 275.75, 275.95, 276.85, 276.15, 275.55, 276.25, 275.95, 275.35, 
    275.85, 275.65, 276.35, 276.35, 276.35, 276.65, 277.35, 276.15, 276.15, 
    275.45, 275.25, 278.35, 275.45, 275.55, 275.65, 276.55, 275.65, 276.55, 
    276.25, 275.95, 275.75, 275.35, 275.65, 275.75, 275.65, 275.85, 275.45, 
    275.75, 275.95, 275.85, 276.15, 276.15, 275.85, 276.15, 275.95, 276.25, 
    276.15, 276.15, 276.05, 275.65, 275.55, 275.25, 275.05, 275.25, 275.65, 
    275.55, 276.25, 277.15, 277.85, 278.15, 277.15, 277.35, 277.95, 277.45, 
    277.85, 277.25, 276.15, 276.55, 275.85, 275.95, 276.45, 276.65, 277.35, 
    276.65, 276.65, 275.95, 276.15, 277.45, 277.15, 277.45, 277.65, 277.05, 
    276.85, 277.05, 276.25, 276.15, 276.55, 276.65, 276.45, 276.35, 276.45, 
    276.45, 276.85, 277.25, 277.05, 276.65, 275.75, 276.25, 276.75, 276.15, 
    275.75, 276.35, 276.55, 276.55, 276.45, 275.85, 276.45, 276.25, 276.15, 
    275.95, 276.15, 275.85, 276.65, 276.95, 277.05, 277.85, 277.45, 277.05, 
    277.65, 277.25, 277.35, 277.15, 277.25, 277.35, 277.65, 278.05, 279.25, 
    278.95, 278.05, 276.65, 275.85, 276.15, 275.85, 276.45, 278.55, 280.15, 
    278.65, 278.65, 277.85, 277.35, 277.85, 277.65, 278.05, 277.85, 277.35, 
    276.95, 277.15, 277.45, 277.55, 276.65, 277.45, 276.65, 275.75, 275.75, 
    275.55, 275.55, 275.85, 276.35, 275.05, 274.15, 273.95, 274.35, 274.05, 
    273.85, 274.15, 274.45, 274.75, 275.05, 275.25, 275.65, 275.55, 275.05, 
    275.25, 274.85, 274.75, 274.75, 275.55, 276.45, 277.55, 276.85, 278.25, 
    276.45, 275.25, 274.75, 274.65, 275.25, 275.95, 275.15, 275.45, 275.45, 
    275.25, 274.85, 275.05, 275.05, 275.55, 275.55, 275.75, 275.65, 275.75, 
    275.55, 275.55, 275.95, 276.45, 276.55, 276.45, 276.65, 277.05, 277.35, 
    277.65, 277.75, 277.85, 277.75, 277.95, 277.35, 277.05, 277.05, 276.85, 
    279.15, 280.65, 276.45, 277.55, 277.45, 278.45, 279.55, 279.45, 278.45, 
    277.15, 277.95, 277.65, 278.35, 279.15, 278.15, 278.15, 277.65, 278.15, 
    277.25, 276.65, 276.25, 275.05, 274.45, 274.35, 274.45, 274.55, 274.35, 
    274.15, 274.45, 274.85, 274.45, 274.95, 274.25, 274.35, 274.35, 274.35, 
    274.45, 274.15, 274.15, 274.05, 274.05, 273.85, 273.85, 273.75, 273.65, 
    273.75, 273.75, 273.75, 273.95, 273.85, 273.85, 274.15, 274.25, 274.55, 
    274.35, 274.85, 275.05, 275.25, 275.35, 275.15, 275.25, 275.15, 275.05, 
    275.35, 274.45, 274.65, 274.65, 274.35, 273.65, 273.85, 273.75, 273.75, 
    273.75, 274.05, 274.25, 274.55, 274.85, 275.35, 275.25, 275.35, 275.65, 
    276.05, 275.85, 275.65, 276.15, 275.65, 275.15, 275.15, 275.15, 274.95, 
    275.45, 277.45, 277.45, 275.95, 275.85, 275.75, 275.95, 276.55, 276.85, 
    276.75, 276.65, 276.45, 276.65, 275.65, 275.95, 275.45, 275.35, 275.85, 
    275.45, 274.95, 277.65, 276.65, 274.25, 274.05, 274.45, 274.55, 274.55, 
    274.55, 273.95, 274.15, 273.95, 274.05, 274.45, 274.55, 275.05, 275.05, 
    275.55, 275.65, 275.45, 275.05, 274.85, 274.65, 274.55, 274.85, 274.75, 
    274.75, 274.65, 274.35, 273.95, 274.05, 274.25, 274.35, 274.25, 274.25, 
    274.25, 274.45, 274.15, 274.25, 274.35, 274.35, 274.45, 274.25, 274.55, 
    274.45, 274.45, 274.65, 274.55, 274.45, 274.05, 274.55, 275.05, 274.75, 
    275.05, 275.15, 274.75, 274.85, 274.75, 274.95, 274.95, 275.35, 275.15, 
    274.95, 275.35, 275.65, 275.25, 275.05, 274.55, 275.45, 274.95, 274.95, 
    275.05, 274.75, 274.65, 274.55, 274.35, 274.15, 274.05, 273.65, 273.55, 
    273.25, 274.35, 274.25, 274.05, 273.95, 274.05, 274.25, 274.55, 274.35, 
    274.75, 274.75, 274.65, 274.25, 274.45, 274.85, 274.65, 274.25, 274.05, 
    274.85, 273.65, 272.85, 272.55, 272.55, 272.95, 272.75, 272.85, 272.45, 
    273.05, 272.75, 272.25, 273.65, 274.35, 275.15, 274.95, 274.85, 274.95, 
    274.85, 274.45, 274.75, 274.55, 274.25, 274.25, 274.15, 274.15, 274.15, 
    274.35, 274.25, 274.25, 274.35, 274.45, 274.35, 274.35, 274.35, 274.35, 
    274.35, 274.35, 274.45, 274.65, 274.75, 274.75, 274.85, 274.75, 274.65, 
    274.55, 274.65, 274.75, 274.65, 274.25, 274.05, 274.55, 274.85, 274.95, 
    275.05, 274.85, 274.85, 274.65, 274.55, 274.45, 274.35, 274.45, 274.65, 
    274.75, 274.75, 274.65, 274.45, 274.55, 274.65, 274.55, 274.45, 274.15, 
    274.45, 274.05, 273.85, 273.95, 273.65, 273.85, 274.25, 273.75, 273.55, 
    273.25, 273.25, 273.35, 273.45, 273.35, 273.35, 273.45, 273.45, 273.55, 
    273.55, 273.65, 273.45, 273.55, 273.55, 273.55, 273.45, 273.35, 273.25, 
    273.25, 273.35, 273.25, 273.25, 273.45, 273.75, 273.65, 273.85, 274.05, 
    273.95, 273.95, 274.05, 274.15, 274.05, 274.15, 274.95, 275.35, 275.55, 
    275.65, 275.35, 275.85, 275.85, 275.85, 275.45, 274.95, 275.15, 275.35, 
    275.15, 274.75, 274.35, 274.65, 274.55, 274.35, 276.05, 275.45, 275.55, 
    276.05, 276.15, 276.15, 275.95, 275.55, 275.55, 276.75, 278.55, 278.05, 
    277.25, 276.85, 276.85, 276.15, 274.45, 275.95, 275.15, 275.35, 273.95, 
    273.25, 273.25, 272.65, 273.25, 273.15, 274.35, 274.75, 274.55, 275.35, 
    274.75, 274.75, 274.95, 274.75, 274.95, 275.55, 274.85, 275.05, 274.45, 
    274.25, 274.45, 273.85, 273.75, 273.25, 273.45, 273.55, 273.75, 274.15, 
    274.25, 274.25, 274.15, 274.25, 273.65, 274.25, 274.25, 273.65, 274.05, 
    273.65, 273.35, 274.05, 274.55, 275.15, 275.25, 275.45, 275.25, 274.95, 
    274.25, 274.35, 274.45, 274.65, 274.65, 274.75, 274.95, 275.25, 275.55, 
    275.65, 276.05, 276.05, 276.15, 276.35, 275.65, 275.65, 275.75, 276.45, 
    276.25, 276.35, 276.85, 276.05, 276.75, 276.35, 276.35, 276.15, 275.85, 
    275.95, 275.85, 276.45, 276.55, 276.65, 276.35, 275.85, 276.05, 276.05, 
    276.05, 276.05, 275.95, 276.15, 275.95, 275.75, 275.75, 275.85, 276.15, 
    275.95, 276.05, 276.05, 275.65, 276.25, 276.35, 276.45, 276.35, 276.25, 
    277.35, 276.85, 276.95, 276.85, 276.75, 276.45, 276.35, 276.75, 276.65, 
    276.55, 276.85, 277.85, 277.65, 278.05, 277.35, 275.65, 275.15, 274.85, 
    274.65, 274.65, 274.65, 274.65, 274.45, 274.55, 274.75, 274.55, 274.55, 
    274.45, 274.35, 274.35, 274.35, 274.05, 274.05, 274.05, 274.05, 274.05, 
    274.05, 274.25, 274.25, 274.05, 274.25, 274.25, 274.35, 274.35, 274.55, 
    274.75, 274.75, 274.75, 274.75, 274.95, 274.75, 274.75, 274.75, 274.65, 
    274.75, 274.75, 274.75, 274.75, 274.95, 274.75, 274.75, 274.85, 275.05, 
    274.75, 274.85, 274.75, 274.45, 274.95, 275.05, 274.95, 275.25, 275.85, 
    275.85, 275.95, 276.15, 275.85, 276.25, 276.15, 275.35, 275.55, 274.95, 
    274.55, 274.15, 274.05, 273.75, 274.35, 274.25, 274.05, 274.35, 274.05, 
    274.05, 274.05, 274.05, 274.15, 274.15, 274.35, 274.35, 274.35, 274.35, 
    274.45, 274.35, 274.45, 274.35, 273.75, 273.65, 273.75, 273.85, 273.95, 
    273.95, 273.95, 274.25, 274.35, 274.35, 274.25, 273.65, 273.55, 273.65, 
    273.85, 273.85, 274.05, 273.95, 274.25, 274.45, 274.35, 274.45, 274.55, 
    274.65, 274.75, 275.05, 275.05, 274.95, 274.55, 274.55, 274.35, 274.35, 
    274.05, 274.55, 274.45, 273.95, 273.65, 273.65, 273.35, 273.45, 273.65, 
    273.75, 273.45, 273.55, 273.55, 273.75, 273.85, 273.85, 274.05, 273.95, 
    273.95, 273.95, 273.95, 273.75, 273.45, 273.65, 274.05, 274.15, 274.25, 
    274.25, 274.25, 274.15, 274.25, 274.35, 274.65, 274.45, 274.35, 274.45, 
    274.55, 274.75, 275.15, 275.05, 275.25, 276.85, 275.95, 275.45, 274.35, 
    274.75, 274.65, 274.55, 274.15, 273.65, 272.85, 274.25, 274.15, 273.95, 
    274.05, 274.25, 274.15, 274.35, 274.65, 275.25, 274.55, 274.35, 273.95, 
    273.75, 273.95, 273.55, 273.55, 273.55, 273.95, 273.75, 274.05, 274.15, 
    274.15, 274.45, 274.25, 274.35, 273.85, 274.05, 274.55, 274.75, 274.65, 
    274.65, 274.55, 275.05, 275.25, 275.55, 275.75, 275.85, 275.95, 275.95, 
    275.95, 275.95, 275.95, 275.85, 275.75, 275.65, 275.75, 275.75, 275.55, 
    275.25, 275.35, 275.55, 275.85, 275.75, 275.65, 275.65, 275.55, 275.95, 
    276.25, 275.95, 277.05, 276.25, 276.65, 276.95, 278.35, 278.45, 278.45, 
    278.35, 276.35, 276.65, 276.55, 276.25, 276.55, 276.75, 276.95, 276.85, 
    277.95, 277.65, 276.75, 276.45, 275.65, 275.75, 276.15, 276.45, 276.35, 
    276.55, 275.05, 275.55, 275.15, 275.25, 275.65, 275.55, 275.65, 275.95, 
    275.75, 275.45, 275.45, 275.45, 275.35, 275.35, 275.25, 274.85, 274.95, 
    275.15, 275.05, 274.95, 274.95, 274.95, 275.05, 275.15, 276.25, 276.25, 
    276.55, 275.95, 275.55, 275.45, 275.35, 275.15, 275.15, 275.05, 275.25, 
    275.65, 275.85, 276.95, 276.45, 276.15, 275.65, 275.65, 275.35, 275.15, 
    275.85, 275.75, 277.85, 275.55, 276.25, 276.05, 276.35, 276.05, 276.25, 
    275.95, 276.05, 275.75, 275.65, 275.25, 274.45, 274.35, 274.95, 275.05, 
    275.35, 275.75, 276.15, 276.05, 275.95, 276.05, 275.45, 275.45, 275.95, 
    275.55, 275.35, 274.75, 274.95, 275.45, 275.55, 275.05, 274.75, 274.45, 
    274.15, 274.05, 273.95, 273.95, 273.65, 274.05, 273.85, 272.75, 273.25, 
    273.85, 273.35, 273.85, 274.35, 275.05, 275.35, 275.55, 275.25, 275.05, 
    275.15, 275.25, 274.95, 275.25, 275.35, 275.55, 275.05, 275.45, 275.45, 
    275.05, 275.05, 275.05, 274.95, 275.05, 275.55, 274.95, 275.25, 275.15, 
    275.35, 275.55, 275.45, 275.75, 275.65, 275.75, 275.65, 275.75, 275.55, 
    275.25, 275.65, 275.35, 275.65, 275.85, 275.75, 275.95, 275.85, 275.65, 
    275.65, 275.55, 275.35, 274.85, 274.45, 274.75, 274.65, 274.65, 274.75, 
    274.85, 274.65, 273.65, 273.45, 273.35, 273.15, 273.35, 273.45, 273.65, 
    273.55, 273.65, 273.95, 273.85, 274.05, 274.05, 273.55, 273.85, 273.55, 
    273.15, 273.35, 273.85, 274.05, 273.95, 273.95, 274.45, 275.35, 274.95, 
    274.55, 274.45, 274.35, 274.35, 273.95, 273.65, 274.25, 274.35, 274.45, 
    274.55, 274.75, 274.85, 274.75, 274.45, 274.35, 274.45, 274.85, 275.35, 
    275.35, 274.95, 274.95, 275.15, 275.15, 275.15, 274.95, 274.45, 274.75, 
    274.95, 274.75, 274.45, 274.45, 274.25, 274.35, 274.65, 274.75, 274.75, 
    274.75, 274.35, 273.95, 274.25, 274.85, 275.55, 275.75, 275.55, 276.05, 
    276.25, 275.75, 275.75, 275.85, 275.15, 275.05, 274.95, 274.75, 274.65, 
    274.25, 274.25, 273.75, 273.25, 272.65, 272.35, 272.15, 272.05, 271.75, 
    271.55, 271.45, 271.55, 271.35, 271.25, 271.55, 271.75, 272.15, 272.05, 
    272.45, 273.45, 272.55, 272.65, 272.55, 272.15, 271.85, 271.55, 270.95, 
    271.85, 271.55, 271.65, 270.95, 271.95, 271.65, 271.05, 271.65, 272.05, 
    272.35, 272.55, 272.45, 272.25, 272.45, 272.75, 272.35, 272.45, 272.65, 
    272.65, 272.75, 272.75, 272.55, 272.85, 272.85, 272.85, 272.75, 272.95, 
    272.85, 272.35, 272.45, 272.65, 272.65, 272.75, 272.95, 273.15, 272.75, 
    272.05, 271.75, 271.95, 271.55, 271.55, 271.65, 271.55, 271.65, 271.55, 
    271.75, 271.95, 272.35, 272.65, 272.95, 273.25, 273.45, 273.55, 273.65, 
    273.85, 274.15, 274.25, 274.25, 274.35, 274.25, 274.05, 274.25, 273.95, 
    273.35, 273.15, 271.85, 271.95, 271.45, 271.45, 270.85, 270.35, 270.25, 
    270.95, 271.45, 271.95, 272.05, 272.25, 272.65, 272.65, 272.65, 272.95, 
    272.95, 272.75, 272.65, 272.35, 272.35, 272.35, 272.55, 272.35, 272.15, 
    272.35, 272.45, 272.35, 271.95, 272.05, 272.05, 272.05, 271.95, 271.85, 
    271.85, 271.85, 271.75, 271.95, 271.95, 272.45, 272.75, 272.95, 273.05, 
    273.35, 273.65, 273.55, 273.55, 273.65, 274.15, 273.95, 274.15, 274.25, 
    274.15, 274.15, 274.45, 274.55, 274.55, 274.45, 274.55, 274.65, 274.45, 
    274.55, 274.45, 274.55, 274.65, 274.65, 274.65, 274.55, 274.15, 273.65, 
    274.15, 273.85, 273.65, 273.65, 273.65, 273.55, 273.55, 273.15, 273.45, 
    273.45, 273.45, 273.35, 273.15, 272.85, 272.55, 272.55, 272.35, 272.35, 
    272.35, 272.35, 272.05, 272.15, 272.25, 271.95, 271.35, 271.65, 271.65, 
    271.65, 271.35, 271.55, 271.55, 271.35, 271.55, 271.25, 271.05, 271.35, 
    271.05, 271.15, 271.35, 271.35, 271.55, 271.95, 272.05, 271.95, 272.15, 
    272.15, 271.95, 272.15, 271.85, 271.85, 271.65, 270.95, 271.05, 270.75, 
    271.15, 271.55, 271.75, 271.85, 271.95, 271.95, 272.05, 271.85, 271.75, 
    271.95, 271.95, 271.85, 271.75, 271.95, 271.75, 271.45, 272.25, 272.15, 
    271.95, 271.95, 271.75, 271.55, 271.35, 271.55, 271.25, 271.55, 271.75, 
    271.75, 271.75, 271.85, 271.55, 271.75, 271.55, 270.85, 271.35, 271.45, 
    271.55, 271.65, 271.65, 271.45, 271.25, 271.55, 271.65, 271.75, 271.55, 
    271.25, 271.45, 270.65, 270.45, 270.65, 272.05, 271.85, 271.95, 272.05, 
    272.15, 271.95, 272.15, 272.25, 272.05, 272.35, 272.15, 272.05, 272.05, 
    271.75, 272.05, 272.05, 271.05, 271.75, 271.85, 271.55, 271.35, 271.75, 
    271.95, 272.15, 272.35, 272.05, 273.15, 272.75, 273.05, 272.75, 272.65, 
    272.55, 272.45, 272.15, 272.15, 272.15, 272.45, 272.55, 272.15, 272.15, 
    272.15, 272.35, 271.75, 271.55, 271.75, 271.65, 271.45, 271.35, 271.55, 
    272.05, 272.45, 272.05, 272.35, 272.75, 273.05, 273.15, 273.45, 273.45, 
    273.35, 273.45, 273.35, 273.25, 273.35, 273.45, 273.65, 273.85, 273.95, 
    273.85, 273.95, 274.05, 274.05, 274.25, 274.35, 274.45, 274.45, 274.45, 
    274.65, 276.25, 275.45, 276.05, 275.05, 275.15, 275.05, 275.95, 276.35, 
    276.05, 275.55, 275.05, 275.65, 276.25, 274.55, 275.45, 274.25, 274.25, 
    274.05, 273.95, 274.85, 274.75, 274.85, 275.15, 275.15, 275.05, 274.95, 
    274.95, 274.85, 274.85, 274.75, 274.75, 274.75, 274.65, 274.55, 274.45, 
    274.45, 274.65, 274.55, 274.65, 275.05, 274.35, 273.95, 273.95, 273.95, 
    274.15, 273.95, 273.85, 273.75, 273.65, 273.35, 273.05, 272.85, 272.85, 
    272.85, 272.25, 272.65, 272.55, 272.45, 271.95, 271.95, 272.05, 271.85, 
    271.65, 271.55, 271.65, 271.65, 271.55, 271.35, 271.05, 271.05, 271.05, 
    271.15, 271.25, 271.15, 271.25, 271.05, 271.15, 271.15, 271.45, 271.25, 
    271.05, 270.95, 270.95, 270.85, 270.85, 270.75, 270.75, 270.55, 270.55, 
    270.45, 270.35, 270.05, 270.15, 270.05, 270.25, 270.35, 270.65, 270.65, 
    270.75, 270.95, 271.15, 271.25, 271.45, 271.55, 269.95, 270.45, 269.75, 
    268.75, 270.65, 270.35, 270.85, 270.75, 270.95, 270.45, 271.35, 271.05, 
    270.75, 271.65, 271.55, 271.75, 271.95, 270.15, 269.85, 270.25, 271.45, 
    271.45, 270.55, 270.35, 269.95, 269.65, 270.05, 270.25, 270.05, 269.65, 
    269.95, 270.15, 270.35, 270.05, 270.35, 270.05, 269.85, 269.05, 269.25, 
    270.05, 271.85, 271.75, 272.05, 272.05, 271.85, 271.75, 271.75, 271.55, 
    271.05, 270.95, 270.95, 270.85, 271.45, 271.35, 270.95, 271.05, 270.55, 
    269.75, 270.05, 269.45, 269.85, 270.15, 270.65, 270.75, 270.25, 270.55, 
    270.65, 270.75, 270.95, 271.05, 271.25, 271.55, 272.05, 272.55, 273.05, 
    273.05, 273.15, 273.05, 273.15, 273.15, 273.05, 273.05, 272.95, 272.95, 
    273.05, 273.05, 272.95, 272.95, 272.85, 272.85, 272.85, 272.85, 272.95, 
    272.85, 272.25, 272.25, 273.15, 272.95, 273.05, 273.15, 273.15, 273.05, 
    273.15, 273.15, 273.25, 273.15, 273.25, 273.35, 273.35, 273.35, 273.15, 
    273.05, 273.45, 273.35, 273.35, 273.35, 273.35, 272.85, 272.85, 272.85, 
    272.85, 272.75, 272.95, 272.85, 272.75, 272.65, 272.25, 272.55, 272.75, 
    272.65, 272.55, 272.25, 272.25, 272.05, 272.15, 271.95, 272.15, 271.85, 
    271.65, 271.45, 271.55, 271.85, 271.35, 271.65, 271.65, 271.55, 271.35, 
    271.55, 271.05, 271.25, 271.85, 271.75, 271.65, 271.35, 270.95, 270.85, 
    270.35, 270.25, 270.65, 270.75, 270.95, 270.95, 270.85, 270.55, 270.45, 
    270.65, 270.75, 270.75, 270.45, 270.45, 270.15, 270.05, 270.05, 270.15, 
    270.45, 270.65, 270.55, 270.75, 270.65, 271.15, 270.95, 271.15, 271.15, 
    270.85, 271.45, 271.75, 271.55, 271.75, 271.85, 271.65, 271.75, 271.35, 
    270.95, 271.15, 271.25, 271.05, 271.05, 271.05, 271.25, 271.15, 271.05, 
    271.35, 271.35, 271.65, 271.25, 271.45, 271.85, 271.75, 271.55, 271.85, 
    272.45, 272.75, 272.95, 272.95, 272.95, 272.95, 273.05, 272.95, 272.75, 
    272.45, 272.15, 271.75, 271.45, 271.35, 271.05, 270.75, 270.55, 270.45, 
    270.35, 270.25, 270.25, 270.45, 270.25, 269.85, 270.35, 270.45, 270.75, 
    270.35, 270.75, 270.75, 270.65, 270.65, 270.65, 270.55, 270.55, 270.45, 
    270.45, 270.35, 270.55, 270.45, 270.05, 270.05, 271.05, 270.95, 271.15, 
    271.05, 271.35, 271.35, 271.35, 271.45, 271.45, 271.25, 270.95, 269.65, 
    269.55, 270.65, 270.55, 270.55, 270.65, 270.65, 271.15, 270.15, 270.35, 
    270.25, 270.25, 268.75, 269.15, 270.25, 270.65, 269.65, 268.75, 268.95, 
    269.15, 269.65, 270.35, 270.15, 270.05, 269.65, 269.35, 269.35, 268.95, 
    269.15, 269.05, 268.95, 269.05, 268.85, 269.15, 268.85, 269.35, 269.55, 
    269.45, 269.45, 269.45, 269.35, 269.15, 269.25, 269.35, 269.35, 269.35, 
    269.55, 269.45, 269.55, 269.35, 269.55, 269.55, 269.75, 269.85, 270.05, 
    270.05, 270.15, 270.25, 270.35, 268.25, 269.45, 270.15, 270.45, 271.25, 
    270.25, 270.85, 270.85, 272.05, 271.75, 272.25, 272.65, 272.35, 272.65, 
    272.75, 273.05, 273.25, 273.25, 272.95, 272.95, 271.95, 271.95, 270.95, 
    270.15, 270.65, 269.75, 270.45, 270.65, 270.85, 270.05, 271.05, 271.05, 
    271.45, 272.45, 272.95, 272.95, 273.35, 273.85, 273.95, 273.65, 273.35, 
    273.85, 274.05, 273.85, 273.85, 273.85, 273.85, 273.65, 273.65, 273.55, 
    273.45, 273.55, 273.65, 273.45, 273.75, 273.65, 273.85, 273.75, 274.15, 
    274.25, 274.25, 274.25, 274.25, 274.15, 274.05, 274.15, 274.15, 274.15, 
    274.05, 274.25, 274.25, 274.35, 274.35, 274.25, 274.35, 274.45, 274.45, 
    274.25, 274.15, 274.05, 274.05, 274.15, 274.25, 274.05, 273.75, 273.65, 
    273.55, 274.15, 274.35, 274.05, 274.15, 274.35, 274.25, 274.05, 273.75, 
    273.75, 273.45, 273.35, 273.25, 273.15, 272.95, 272.95, 272.95, 272.85, 
    272.55, 272.25, 272.15, 272.05, 272.05, 271.95, 271.95, 272.05, 272.05, 
    271.85, 271.45, 271.55, 271.95, 271.95, 271.85, 272.15, 271.85, 271.65, 
    271.15, 270.95, 270.85, 270.45, 270.25, 270.35, 270.95, 271.15, 271.05, 
    270.85, 270.95, 270.95, 271.05, 271.55, 271.25, 271.45, 271.45, 271.85, 
    272.05, 272.35, 272.45, 272.55, 272.55, 272.25, 272.35, 271.75, 271.75, 
    271.65, 271.85, 271.15, 271.45, 271.55, 271.75, 272.15, 272.05, 272.25, 
    272.75, 272.65, 272.45, 272.35, 272.55, 272.25, 272.05, 271.55, 271.25, 
    271.25, 271.55, 271.75, 271.65, 271.05, 271.25, 271.05, 270.75, 270.85, 
    271.05, 271.45, 271.45, 272.15, 272.05, 272.05, 272.15, 272.05, 271.85, 
    271.45, 270.35, 270.85, 271.15, 271.05, 270.55, 270.65, 270.65, 270.95, 
    271.85, 270.55, 270.85, 270.65, 270.45, 270.45, 269.95, 270.15, 268.65, 
    269.25, 270.15, 270.85, 271.35, 271.15, 271.25, 271.25, 271.25, 271.35, 
    271.55, 271.55, 272.25, 271.95, 271.85, 271.45, 271.25, 271.65, 271.85, 
    271.85, 272.05, 272.05, 272.05, 272.15, 272.15, 272.35, 272.65, 272.65, 
    272.55, 272.45, 272.25, 272.65, 272.55, 272.45, 272.65, 272.95, 272.95, 
    273.25, 273.55, 273.85, 273.85, 273.95, 273.95, 274.15, 274.15, 274.15, 
    274.05, 273.95, 273.95, 273.95, 273.85, 273.75, 273.75, 273.65, 273.55, 
    273.55, 273.75, 273.85, 273.95, 273.85, 273.75, 273.75, 273.65, 273.55, 
    273.35, 273.35, 273.25, 273.05, 272.45, 272.45, 272.75, 272.75, 272.25, 
    272.05, 272.15, 271.45, 271.25, 271.25, 270.85, 270.95, 271.05, 271.25, 
    271.05, 270.95, 271.35, 270.65, 271.15, 270.35, 269.05, 270.45, 269.85, 
    270.05, 270.85, 271.05, 270.85, 270.65, 270.95, 270.55, 270.35, 270.35, 
    270.35, 269.95, 269.15, 268.15, 267.85, 268.45, 268.65, 268.45, 269.65, 
    269.75, 268.35, 268.55, 268.35, 268.05, 267.25, 267.25, 267.25, 267.15, 
    266.65, 266.15, 267.15, 267.25, 267.15, 267.65, 267.35, 266.65, 267.75, 
    269.35, 269.25, 269.05, 268.85, 268.25, 268.25, 268.15, 267.65, 267.25, 
    265.95, 266.45, 267.55, 266.55, 265.95, 267.35, 266.95, 266.55, 267.15, 
    266.05, 266.95, 267.05, 267.25, 267.25, 266.85, 266.55, 266.45, 266.15, 
    266.15, 266.05, 266.25, 266.35, 266.05, 265.15, 265.15, 265.45, 265.65, 
    265.65, 265.65, 265.75, 265.75, 265.95, 265.75, 265.75, 265.95, 265.85, 
    266.55, 266.85, 266.35, 266.45, 266.35, 266.15, 266.15, 265.85, 265.75, 
    265.85, 265.85, 265.75, 265.95, 265.75, 265.75, 265.85, 265.85, 265.95, 
    265.85, 265.65, 265.85, 266.05, 265.75, 265.25, 264.85, 265.35, 265.65, 
    265.45, 265.65, 265.85, 265.95, 266.35, 266.45, 267.45, 269.05, 268.75, 
    268.55, 269.35, 269.35, 269.45, 269.65, 269.85, 269.65, 269.55, 270.05, 
    270.55, 271.45, 272.25, 272.65, 272.75, 272.75, 272.85, 272.85, 272.85, 
    272.95, 272.85, 272.85, 272.65, 272.65, 272.35, 272.45, 272.25, 272.95, 
    272.55, 271.65, 272.05, 272.45, 272.85, 272.95, 272.55, 271.85, 271.35, 
    271.15, 270.85, 270.45, 270.15, 269.85, 269.45, 269.15, 268.95, 269.05, 
    269.05, 269.15, 269.25, 268.95, 268.75, 269.15, 269.35, 269.35, 269.65, 
    270.25, 270.45, 270.75, 271.05, 271.25, 271.35, 271.35, 271.35, 271.25, 
    271.05, 271.25, 271.45, 271.55, 271.65, 271.75, 271.85, 272.05, 272.35, 
    272.75, 272.25, 271.95, 272.15, 272.75, 269.25, 268.65, 268.25, 267.75, 
    267.45, 266.75, 266.65, 266.65, 266.75, 266.25, 266.15, 265.95, 266.05, 
    266.35, 265.75, 266.25, 266.75, 266.75, 266.35, 266.35, 266.55, 267.05, 
    267.05, 267.25, 267.45, 267.45, 266.65, 265.85, 265.35, 265.45, 265.15, 
    264.85, 265.55, 265.45, 265.55, 265.55, 265.95, 265.85, 265.85, 266.05, 
    266.15, 266.15, 266.25, 266.15, 266.15, 265.95, 265.85, 266.15, 265.55, 
    265.45, 265.35, 265.45, 265.35, 265.85, 265.85, 266.45, 266.65, 267.15, 
    267.65, 267.75, 267.65, 267.75, 267.95, 267.65, 267.95, 267.95, 267.85, 
    267.45, 267.85, 268.55, 268.75, 268.85, 268.85, 268.75, 268.65, 268.35, 
    267.05, 268.05, 269.55, 269.55, 269.45, 269.25, 269.45, 269.25, 269.45, 
    268.75, 269.15, 269.55, 269.15, 269.25, 269.65, 269.35, 269.35, 269.65, 
    269.45, 269.55, 269.35, 269.45, 269.05, 268.85, 268.35, 268.25, 268.05, 
    267.65, 267.35, 266.75, 266.35, 266.55, 265.85, 266.55, 266.65, 267.25, 
    266.55, 265.85, 267.55, 267.45, 266.05, 267.15, 267.35, 267.05, 266.85, 
    266.55, 266.55, 266.35, 266.15, 265.95, 265.55, 265.55, 265.65, 265.15, 
    265.55, 265.45, 265.65, 266.55, 266.35, 266.05, 265.75, 265.65, 265.55, 
    265.85, 265.65, 265.75, 266.15, 266.05, 266.25, 266.25, 266.45, 266.65, 
    266.75, 266.45, 266.85, 266.85, 266.15, 265.65, 265.95, 266.65, 266.85, 
    266.75, 266.45, 266.45, 266.55, 266.45, 266.85, 266.65, 266.75, 266.85, 
    267.05, 267.15, 267.05, 267.25, 267.25, 267.35, 267.55, 267.35, 267.95, 
    267.85, 268.15, 268.75, 269.05, 269.15, 269.45, 270.05, 270.35, 270.55, 
    271.05, 271.15, 271.45, 271.85, 272.15, 272.35, 272.55, 272.65, 272.65, 
    272.65, 272.55, 272.55, 272.45, 272.35, 272.45, 272.65, 272.95, 273.05, 
    273.25, 273.35, 273.35, 273.35, 273.45, 273.35, 273.35, 273.05, 273.15, 
    273.15, 273.35, 273.35, 273.25, 273.35, 273.25, 273.25, 273.35, 273.45, 
    273.45, 273.45, 273.35, 273.35, 272.95, 272.15, 271.95, 272.85, 272.55, 
    272.25, 272.45, 272.25, 272.15, 272.45, 272.65, 272.75, 272.85, 272.85, 
    272.75, 272.85, 272.25, 272.05, 271.65, 271.35, 270.85, 270.25, 270.45, 
    271.15, 271.45, 271.25, 271.15, 271.25, 271.05, 271.25, 271.35, 271.25, 
    271.05, 270.25, 269.65, 268.65, 268.05, 267.95, 268.05, 267.75, 267.45, 
    267.45, 267.45, 267.25, 267.55, 267.15, 267.05, 267.15, 267.45, 267.55, 
    267.85, 269.35, 268.95, 268.85, 269.25, 269.85, 269.35, 270.25, 270.85, 
    269.45, 269.35, 269.05, 268.35, 267.65, 267.15, 266.45, 266.15, 265.45, 
    265.55, 265.45, 264.85, 264.55, 264.25, 264.35, 264.15, 263.75, 263.25, 
    263.05, 263.25, 263.05, 263.35, 262.95, 262.85, 262.95, 263.05, 263.45, 
    263.75, 264.05, 263.95, 264.05, 264.15, 263.35, 264.45, 265.65, 266.05, 
    266.15, 266.85, 268.55, 268.95, 270.35, 270.35, 270.65, 270.85, 270.95, 
    270.35, 270.75, 270.95, 271.05, 270.85, 271.65, 271.65, 270.95, 270.95, 
    266.85, 265.95, 264.95, 264.75, 263.25, 263.05, 263.85, 264.05, 263.45, 
    263.15, 262.65, 261.75, 261.15, 260.65, 261.05, 260.95, 261.15, 261.45, 
    261.65, 261.75, 262.35, 262.55, 262.45, 262.35, 262.55, 262.35, 261.95, 
    262.15, 262.35, 262.35, 262.55, 262.95, 262.35, 262.55, 262.65, 262.45, 
    262.35, 262.65, 262.65, 262.75, 263.05, 263.15, 263.75, 264.35, 265.25, 
    266.55, 267.45, 267.95, 268.55, 267.95, 268.55, 268.85, 268.55, 269.05, 
    269.15, 269.35, 268.65, 269.75, 270.45, 270.55, 270.55, 271.25, 271.05, 
    271.85, 271.15, 271.05, 271.35, 271.85, 271.75, 271.95, 272.25, 272.45, 
    272.65, 273.05, 273.25, 273.55, 273.55, 273.55, 273.35, 273.35, 273.45, 
    273.45, 273.25, 274.05, 274.15, 273.95, 273.75, 274.05, 273.15, 273.15, 
    273.15, 272.25, 272.45, 273.05, 272.55, 271.35, 270.65, 271.75, 271.85, 
    271.85, 272.15, 271.75, 271.75, 271.25, 270.35, 270.95, 270.85, 268.95, 
    267.55, 265.85, 264.55, 265.05, 264.45, 263.25, 262.85, 262.25, 262.25, 
    262.25, 262.45, 262.05, 262.25, 262.05, 261.85, 261.65, 261.25, 261.15, 
    260.65, 260.15, 260.35, 259.95, 260.35, 260.35, 260.55, 260.65, 260.55, 
    261.05, 260.75, 261.35, 261.45, 261.05, 261.05, 261.45, 261.45, 261.85, 
    262.05, 262.25, 262.35, 262.65, 262.85, 262.75, 262.65, 262.65, 262.45, 
    262.15, 262.25, 262.05, 262.45, 262.25, 262.85, 263.05, 262.85, 263.25, 
    263.55, 263.45, 263.75, 263.95, 263.95, 264.25, 264.15, 264.35, 264.05, 
    264.25, 264.85, 264.45, 264.15, 263.35, 263.35, 263.45, 263.45, 263.35, 
    263.25, 263.35, 264.05, 264.75, 265.05, 264.95, 264.95, 265.25, 265.05, 
    264.75, 264.65, 264.35, 264.55, 264.35, 264.25, 264.15, 264.35, 264.05, 
    263.85, 263.85, 263.85, 264.25, 263.95, 264.05, 264.25, 263.75, 263.45, 
    263.65, 263.35, 262.65, 263.65, 263.95, 263.85, 264.25, 264.55, 263.65, 
    263.55, 263.35, 263.35, 263.75, 263.45, 263.85, 264.05, 263.25, 263.45, 
    264.35, 263.75, 263.95, 264.35, 264.55, 264.65, 265.55, 266.35, 266.25, 
    266.25, 265.75, 265.95, 265.65, 265.55, 263.55, 262.75, 263.45, 263.95, 
    263.35, 262.85, 263.65, 263.15, 262.75, 262.85, 263.15, 262.45, 263.45, 
    264.35, 264.45, 264.65, 262.75, 263.85, 262.85, 261.25, 262.85, 264.45, 
    264.85, 264.95, 264.45, 264.15, 263.95, 264.95, 264.35, 264.85, 264.75, 
    264.75, 264.75, 265.05, 265.45, 265.35, 265.65, 265.55, 265.45, 265.25, 
    264.35, 264.15, 264.85, 264.35, 264.45, 264.05, 263.75, 264.25, 264.35, 
    264.75, 263.25, 264.05, 264.25, 265.95, 266.65, 267.05, 267.55, 267.95, 
    268.05, 267.65, 267.75, 268.15, 268.65, 269.15, 269.05, 269.15, 269.35, 
    269.65, 270.15, 270.55, 270.65, 270.85, 270.75, 270.55, 270.35, 270.35, 
    270.45, 270.35, 269.65, 269.05, 269.45, 269.75, 269.55, 269.25, 269.25, 
    269.35, 269.35, 269.55, 269.15, 268.65, 268.25, 267.55, 268.15, 267.95, 
    267.85, 268.05, 267.45, 267.35, 267.75, 268.05, 268.25, 267.85, 267.55, 
    266.55, 267.45, 266.95, 266.85, 266.95, 266.45, 266.65, 266.55, 266.45, 
    266.95, 267.15, 267.25, 267.15, 266.95, 267.05, 267.05, 267.15, 266.75, 
    266.55, 266.35, 266.35, 266.35, 266.05, 266.05, 266.15, 266.25, 265.95, 
    265.45, 265.85, 265.35, 265.45, 265.75, 265.85, 265.75, 265.95, 265.85, 
    265.75, 265.65, 265.45, 265.45, 265.25, 265.15, 265.05, 265.35, 265.65, 
    265.65, 265.55, 265.55, 265.65, 265.65, 265.65, 265.35, 265.35, 265.45, 
    265.35, 265.45, 265.55, 265.75, 265.95, 266.15, 266.15, 266.15, 266.35, 
    266.75, 266.85, 266.75, 266.95, 266.95, 267.05, 267.05, 266.85, 266.95, 
    266.75, 266.55, 266.95, 267.05, 267.05, 267.15, 267.45, 267.75, 268.15, 
    268.55, 268.45, 268.35, 268.15, 268.05, 267.75, 267.85, 268.25, 267.95, 
    267.75, 267.85, 267.85, 267.75, 267.45, 267.65, 267.75, 268.05, 268.65, 
    269.45, 269.55, 269.85, 270.35, 270.65, 271.45, 271.75, 272.35, 272.55, 
    272.65, 272.85, 272.45, 272.15, 272.05, 271.95, 271.95, 272.05, 271.85, 
    272.15, 272.45, 272.35, 272.35, 272.15, 272.15, 272.15, 272.25, 272.65, 
    272.75, 272.85, 273.45, 274.65, 273.35, 273.95, 273.75, 273.55, 273.75, 
    272.85, 273.05, 272.95, 272.95, 272.75, 272.85, 272.85, 272.95, 272.95, 
    272.95, 272.85, 272.65, 272.75, 272.75, 272.75, 272.75, 272.65, 272.75, 
    272.75, 272.65, 272.45, 272.35, 271.15, 271.45, 271.65, 271.85, 271.65, 
    272.15, 272.25, 271.85, 272.25, 272.15, 272.45, 272.65, 272.85, 272.75, 
    272.65, 272.85, 272.75, 272.55, 272.35, 272.45, 272.75, 272.45, 272.25, 
    272.25, 272.05, 271.85, 271.85, 271.75, 271.75, 271.85, 271.85, 271.65, 
    271.55, 271.45, 271.45, 271.45, 271.55, 271.35, 271.35, 271.25, 271.35, 
    271.25, 271.45, 271.45, 270.95, 270.85, 270.75, 270.55, 270.55, 270.25, 
    270.05, 269.85, 269.45, 269.35, 269.25, 268.25, 268.85, 268.55, 268.65, 
    267.35, 267.95, 268.05, 268.55, 268.55, 269.25, 269.65, 269.55, 269.85, 
    269.35, 269.55, 270.15, 270.55, 271.05, 271.45, 271.35, 270.95, 270.85, 
    271.05, 270.95, 270.65, 270.45, 270.35, 270.05, 270.05, 269.65, 269.05, 
    269.05, 270.75, 268.45, 268.35, 268.15, 267.85, 267.85, 267.35, 266.85, 
    266.35, 265.95, 265.55, 265.55, 265.05, 264.25, 264.15, 262.95, 262.25, 
    262.35, 261.15, 260.55, 260.15, 260.25, 259.75, 260.75, 260.65, 262.35, 
    262.75, 262.75, 263.25, 263.85, 263.85, 264.35, 262.85, 264.15, 264.05, 
    264.45, 264.35, 263.65, 263.85, 262.95, 264.65, 265.55, 265.65, 265.85, 
    266.25, 266.55, 267.05, 266.95, 266.95, 264.85, 263.35, 262.55, 261.55, 
    259.95, 259.75, 259.95, 258.95, 258.15, 258.45, 258.75, 259.95, 260.85, 
    260.15, 260.45, 260.45, 260.95, 261.25, 261.65, 262.05, 262.65, 263.45, 
    263.65, 263.85, 264.05, 264.65, 267.45, 268.05, 268.35, 267.85, 267.25, 
    267.85, 268.25, 268.25, 269.05, 269.25, 269.35, 269.35, 269.35, 269.15, 
    269.05, 268.95, 268.65, 268.45, 268.05, 268.65, 268.25, 267.95, 267.85, 
    267.95, 267.95, 267.85, 268.25, 268.15, 268.25, 268.15, 268.35, 268.35, 
    267.65, 267.15, 266.75, 266.65, 266.95, 267.25, 266.95, 266.75, 267.25, 
    269.05, 269.15, 269.45, 270.15, 270.65, 270.35, 270.95, 271.25, 271.25, 
    271.25, 270.75, 270.15, 269.65, 268.25, 269.15, 269.65, 270.45, 270.65, 
    270.85, 271.15, 271.25, 271.05, 271.35, 271.65, 271.95, 272.55, 271.55, 
    272.25, 271.05, 269.55, 270.35, 270.75, 271.15, 272.05, 272.05, 272.15, 
    270.15, 268.35, 266.55, 265.95, 265.25, 265.05, 264.35, 263.85, 263.35, 
    262.95, 262.75, 262.95, 262.95, 262.85, 262.75, 263.05, 262.85, 263.05, 
    263.05, 263.05, 263.15, 263.45, 263.55, 263.35, 263.25, 262.75, 262.85, 
    262.55, 262.25, 262.05, 262.15, 262.45, 262.15, 261.75, 261.85, 261.95, 
    261.75, 262.15, 262.55, 262.55, 262.85, 263.05, 262.95, 263.05, 263.25, 
    263.25, 262.65, 262.85, 262.75, 262.85, 262.85, 262.65, 262.95, 262.85, 
    263.35, 263.25, 263.25, 263.45, 263.65, 263.35, 262.45, 263.85, 263.65, 
    263.65, 263.15, 263.25, 264.35, 265.15, 265.35, 266.45, 267.55, 268.35, 
    269.25, 270.15, 270.95, 271.55, 271.85, 272.15, 272.35, 272.25, 272.35, 
    272.55, 272.65, 272.55, 271.75, 271.25, 270.25, 269.95, 269.65, 268.65, 
    267.85, 267.35, 267.05, 266.35, 266.55, 266.45, 266.45, 265.45, 265.55, 
    265.15, 265.95, 265.95, 265.55, 265.55, 265.45, 265.45, 265.45, 265.25, 
    265.15, 265.15, 265.35, 265.25, 264.85, 264.85, 264.75, 265.15, 265.35, 
    265.45, 265.55, 265.85, 266.65, 267.15, 268.05, 269.15, 269.75, 270.55, 
    271.05, 271.25, 271.45, 271.25, 271.15, 271.35, 271.55, 271.85, 271.95, 
    271.65, 271.35, 271.95, 272.15, 272.15, 271.95, 272.15, 271.75, 271.95, 
    272.05, 271.85, 271.45, 271.75, 269.35, 269.05, 268.95, 268.95, 269.45, 
    270.15, 269.75, 269.45, 269.05, 268.75, 269.15, 269.45, 269.55, 270.25, 
    270.75, 271.65, 272.25, 272.25, 271.65, 271.25, 270.75, 268.75, 267.25, 
    266.85, 266.65, 265.65, 265.05, 264.15, 263.15, 261.95, 260.85, 260.35, 
    259.55, 258.55, 257.95, 257.15, 257.15, 256.55, 256.05, 256.15, 256.35, 
    256.15, 256.65, 256.95, 257.15, 257.05, 257.15, 257.75, 257.95, 258.15, 
    258.35, 258.35, 260.45, 260.85, 261.05, 261.85, 261.95, 261.75, 262.45, 
    259.95, 259.25, 258.85, 258.75, 258.35, 258.15, 258.15, 258.05, 258.05, 
    258.35, 258.35, 258.45, 258.65, 258.65, 258.85, 258.65, 258.85, 259.25, 
    259.05, 258.95, 259.05, 259.35, 259.55, 259.55, 259.55, 259.75, 259.95, 
    260.25, 260.45, 260.35, 260.75, 260.55, 260.75, 260.95, 260.85, 260.95, 
    261.15, 261.25, 258.05, 261.25, 261.15, 261.35, 261.65, 261.75, 261.45, 
    261.65, 261.35, 260.85, 260.55, 259.95, 259.15, 258.15, 257.55, 257.05, 
    256.25, 256.35, 255.75, 255.65, 255.55, 255.45, 255.55, 254.95, 254.05, 
    253.95, 254.15, 253.75, 254.05, 253.85, 254.05, 254.35, 254.65, 254.25, 
    254.55, 254.45, 253.95, 253.95, 253.75, 253.45, 253.55, 253.55, 254.65, 
    254.85, 254.85, 255.55, 255.65, 255.25, 254.85, 254.75, 254.65, 254.55, 
    254.65, 254.05, 254.25, 253.75, 253.15, 252.35, 252.15, 252.35, 252.25, 
    253.15, 254.15, 253.85, 253.75, 254.05, 254.45, 254.65, 254.15, 254.55, 
    254.25, 254.45, 254.35, 253.95, 254.15, 254.75, 254.55, 254.75, 254.55, 
    254.25, 253.85, 254.35, 256.15, 256.95, 257.45, 256.65, 257.45, 257.35, 
    257.55, 257.95, 257.95, 258.45, 258.55, 258.35, 258.75, 257.85, 257.55, 
    257.65, 257.45, 257.35, 257.25, 257.05, 257.35, 257.05, 258.35, 256.55, 
    256.45, 256.85, 257.15, 257.25, 257.45, 258.05, 257.75, 257.25, 256.75, 
    256.45, 256.45, 256.35, 256.15, 256.45, 256.45, 256.85, 256.95, 256.85, 
    256.15, 256.15, 256.55, 256.85, 256.35, 256.05, 256.05, 256.25, 256.35, 
    255.85, 256.05, 256.15, 255.95, 255.75, 255.25, 254.95, 254.85, 254.95, 
    254.85, 254.75, 254.85, 255.25, 254.95, 254.85, 254.35, 254.75, 254.45, 
    254.65, 255.65, 256.45, 255.95, 256.05, 256.35, 257.05, 255.95, 254.55, 
    253.85, 253.65, 253.85, 254.15, 253.85, 254.25, 254.05, 254.15, 253.75, 
    253.95, 254.05, 254.25, 254.75, 255.25, 255.15, 255.45, 255.55, 255.25, 
    255.65, 255.95, 255.85, 256.55, 256.55, 256.35, 255.85, 256.05, 256.65, 
    257.85, 257.35, 258.45, 260.25, 261.35, 262.05, 262.65, 263.45, 263.75, 
    264.45, 265.25, 265.75, 266.05, 266.55, 266.95, 267.25, 267.25, 267.75, 
    267.95, 268.25, 268.25, 268.15, 268.35, 268.45, 268.55, 268.55, 268.85, 
    268.75, 268.05, 267.35, 266.65, 265.35, 265.45, 265.15, 264.25, 262.75, 
    260.75, 259.85, 263.45, 259.15, 258.65, 258.55, 258.35, 258.05, 257.75, 
    257.85, 258.15, 258.15, 258.15, 257.85, 257.65, 258.25, 258.55, 258.05, 
    258.25, 261.25, 258.85, 258.95, 258.55, 259.15, 259.45, 259.45, 258.65, 
    258.55, 256.85, 256.35, 260.05, 259.65, 259.35, 260.25, 260.65, 259.85, 
    260.15, 260.75, 260.35, 260.75, 260.35, 260.25, 260.35, 260.35, 260.15, 
    260.95, 260.25, 260.35, 260.65, 260.55, 260.35, 260.15, 259.95, 260.35, 
    260.75, 261.05, 261.55, 261.95, 262.25, 262.55, 262.65, 262.75, 262.35, 
    262.15, 261.75, 262.35, 261.35, 260.95, 261.25, 261.15, 261.35, 261.25, 
    261.25, 260.95, 260.75, 260.75, 260.65, 260.85, 261.05, 260.65, 260.75, 
    259.85, 258.95, 259.05, 259.25, 259.25, 259.65, 260.35, 258.85, 259.15, 
    259.65, 259.85, 260.15, 260.05, 260.25, 260.55, 260.45, 260.35, 260.45, 
    260.45, 260.65, 260.65, 260.65, 260.95, 260.85, 261.15, 261.35, 261.55, 
    262.15, 263.05, 263.55, 263.15, 263.45, 263.55, 263.55, 263.55, 263.35, 
    263.45, 263.75, 264.15, 264.15, 264.15, 264.45, 265.25, 265.05, 264.85, 
    264.55, 264.35, 264.15, 264.05, 264.05, 263.95, 263.15, 262.75, 262.45, 
    261.85, 261.55, 260.85, 260.15, 260.05, 259.95, 259.85, 259.45, 259.15, 
    259.15, 258.95, 258.75, 258.35, 258.05, 258.05, 257.95, 257.85, 257.45, 
    257.25, 256.95, 256.05, 255.65, 254.85, 254.65, 254.65, 254.55, 254.55, 
    254.65, 254.95, 255.35, 255.45, 255.65, 256.15, 255.85, 255.95, 256.05, 
    255.85, 256.35, 256.55, 256.45, 256.45, 256.45, 256.45, 256.55, 256.15, 
    256.25, 256.25, 256.75, 257.05, 257.15, 257.15, 257.55, 257.35, 257.05, 
    256.75, 256.75, 257.15, 256.75, 258.55, 259.05, 259.25, 259.35, 259.05, 
    259.25, 259.95, 260.25, 260.35, 260.65, 261.35, 260.45, 260.95, 261.05, 
    261.75, 261.15, 261.25, 261.35, 261.45, 261.65, 261.75, 261.05, 261.35, 
    260.35, 260.65, 260.35, 259.65, 259.05, 258.95, 259.15, 260.25, 260.25, 
    260.85, 261.15, 261.15, 259.65, 258.95, 257.35, 256.45, 255.95, 256.45, 
    256.75, 256.95, 256.65, 255.55, 255.85, 255.55, 254.35, 255.45, 257.05, 
    258.75, 257.75, 258.45, 258.05, 258.45, 257.65, 256.95, 257.25, 256.25, 
    256.55, 256.45, 256.05, 256.65, 257.35, 257.75, 258.15, 257.95, 257.65, 
    257.65, 256.15, 256.45, 256.25, 256.55, 256.55, 256.85, 257.25, 256.15, 
    257.55, 256.05, 255.15, 254.55, 254.65, 255.35, 254.85, 254.45, 254.75, 
    255.05, 254.75, 254.75, 255.45, 255.85, 255.35, 255.15, 254.95, 254.85, 
    253.95, 254.65, 255.25, 255.35, 254.45, 254.65, 255.45, 254.95, 253.95, 
    253.85, 253.45, 253.15, 252.65, 252.55, 252.65, 253.05, 253.65, 252.65, 
    253.25, 252.85, 251.95, 251.75, 252.25, 254.25, 254.05, 253.45, 252.25, 
    251.85, 251.95, 251.85, 251.95, 253.25, 252.95, 252.15, 252.45, 252.85, 
    253.55, 254.75, 253.25, 252.95, 251.85, 252.05, 252.95, 251.85, 251.55, 
    251.25, 251.05, 250.15, 249.55, 250.65, 250.85, 248.85, 249.15, 248.35, 
    248.45, 248.75, 248.85, 249.15, 249.25, 249.45, 249.75, 249.95, 250.35, 
    249.85, 250.55, 249.95, 250.75, 250.85, 251.05, 251.45, 252.15, 252.35, 
    252.15, 252.35, 252.25, 252.65, 252.95, 253.15, 252.65, 253.05, 253.15, 
    253.45, 253.95, 253.95, 252.25, 251.95, 251.75, 252.15, 252.35, 252.15, 
    251.85, 251.25, 251.45, 250.85, 250.85, 251.55, 252.05, 252.25, 252.15, 
    252.15, 252.15, 252.25, 251.25, 251.25, 251.15, 250.75, 250.15, 250.65, 
    250.25, 250.15, 249.95, 249.45, 249.85, 249.85, 249.85, 249.75, 249.85, 
    250.75, 251.05, 251.45, 252.45, 253.55, 254.15, 254.55, 253.95, 253.15, 
    253.45, 253.35, 253.25, 253.45, 254.05, 253.85, 253.85, 253.35, 252.55, 
    253.15, 253.65, 253.85, 253.35, 253.05, 253.65, 254.65, 254.15, 254.85, 
    253.65, 254.65, 256.45, 257.15, 256.65, 256.45, 256.45, 256.25, 257.65, 
    257.85, 258.05, 257.25, 257.05, 257.35, 257.75, 257.85, 257.75, 257.65, 
    257.95, 258.15, 258.15, 257.75, 258.05, 257.65, 258.05, 257.85, 257.65, 
    258.35, 258.05, 258.65, 259.55, 260.15, 260.35, 260.35, 260.75, 261.25, 
    261.65, 262.25, 262.95, 263.75, 264.25, 264.55, 265.15, 265.85, 266.25, 
    266.65, 266.55, 266.45, 266.55, 266.65, 266.95, 267.25, 267.15, 267.25, 
    266.65, 267.35, 267.35, 266.75, 266.45, 267.05, 266.55, 265.25, 265.65, 
    265.35, 264.85, 264.55, 263.45, 263.25, 262.75, 262.35, 261.75, 261.75, 
    262.25, 262.35, 263.35, 263.15, 263.75, 263.85, 263.75, 259.85, 263.85, 
    264.05, 263.45, 263.45, 265.05, 263.35, 263.35, 263.05, 263.75, 264.05, 
    263.65, 264.15, 263.25, 262.65, 262.55, 263.25, 264.15, 263.45, 262.95, 
    263.95, 264.45, 264.45, 264.55, 264.95, 264.95, 265.75, 266.45, 266.75, 
    266.75, 267.15, 267.15, 268.05, 268.05, 267.55, 267.55, 267.45, 267.15, 
    267.65, 266.95, 267.45, 266.75, 266.65, 266.65, 266.35, 266.75, 267.05, 
    267.75, 267.45, 267.15, 267.35, 267.25, 267.45, 266.75, 265.95, 266.35, 
    265.75, 266.05, 266.45, 266.85, 267.45, 267.95, 267.65, 267.75, 267.05, 
    267.25, 267.35, 267.65, 267.85, 267.55, 267.45, 267.25, 266.65, 266.65, 
    266.25, 266.05, 265.45, 265.45, 265.25, 263.95, 263.65, 263.95, 265.65, 
    266.65, 266.85, 267.05, 267.15, 267.35, 267.05, 267.05, 267.15, 267.35, 
    267.35, 267.35, 267.45, 267.55, 267.65, 267.55, 267.75, 267.85, 267.75, 
    267.55, 267.65, 267.65, 267.75, 268.05, 268.15, 268.05, 268.25, 268.55, 
    268.65, 268.55, 268.55, 268.65, 268.95, 268.55, 268.45, 268.95, 269.15, 
    269.05, 268.95, 268.65, 268.75, 268.75, 269.05, 268.85, 268.85, 268.95, 
    269.05, 269.25, 269.45, 269.45, 269.55, 269.65, 269.75, 269.75, 269.85, 
    269.75, 269.65, 269.75, 269.65, 269.75, 269.75, 269.55, 269.55, 269.55, 
    269.55, 269.55, 269.55, 269.45, 269.65, 269.75, 269.65, 269.65, 269.55, 
    269.65, 269.75, 269.65, 269.65, 269.15, 269.55, 269.25, 269.55, 269.45, 
    269.45, 269.45, 269.25, 269.25, 269.25, 268.35, 268.75, 268.05, 268.55, 
    267.85, 267.95, 268.65, 268.55, 268.75, 268.75, 268.75, 268.35, 268.55, 
    268.75, 268.85, 268.45, 268.55, 268.35, 268.35, 268.35, 268.05, 267.75, 
    268.15, 268.05, 268.15, 268.45, 268.45, 267.85, 268.15, 268.45, 268.65, 
    268.95, 269.15, 269.15, 269.35, 269.35, 269.55, 269.75, 269.65, 269.85, 
    269.85, 269.95, 270.15, 270.35, 270.35, 270.25, 270.35, 270.55, 270.35, 
    270.45, 270.55, 270.65, 270.65, 270.65, 270.55, 270.45, 270.55, 270.55, 
    270.85, 270.65, 270.55, 270.55, 270.85, 270.85, 270.65, 270.45, 270.75, 
    270.65, 270.75, 270.65, 270.55, 270.65, 270.55, 270.55, 270.45, 270.45, 
    270.35, 270.15, 269.95, 269.95, 269.75, 269.55, 269.55, 269.45, 269.35, 
    269.25, 269.25, 269.15, 269.15, 268.85, 268.75, 267.85, 267.85, 268.05, 
    268.15, 268.15, 267.55, 267.35, 266.95, 266.75, 267.35, 267.65, 267.45, 
    266.95, 267.05, 268.25, 266.55, 266.65, 266.75, 267.35, 266.05, 267.05, 
    267.35, 267.05, 266.15, 266.85, 267.25, 266.65, 267.05, 267.15, 267.25, 
    267.15, 267.45, 267.05, 267.65, 266.85, 266.15, 266.65, 266.55, 266.75, 
    267.15, 267.25, 267.35, 266.45, 267.25, 266.85, 266.65, 266.25, 266.05, 
    266.05, 265.85, 265.95, 265.75, 265.05, 264.75, 265.65, 265.45, 265.35, 
    265.45, 265.05, 264.75, 264.75, 264.25, 263.85, 263.45, 263.55, 263.75, 
    263.15, 262.75, 262.75, 263.15, 263.45, 263.65, 263.45, 263.25, 263.95, 
    263.95, 263.75, 263.35, 263.45, 263.45, 263.45, 263.15, 263.35, 263.65, 
    263.65, 263.25, 262.95, 262.85, 262.85, 262.65, 262.45, 262.35, 262.45, 
    262.55, 262.95, 262.75, 262.85, 262.95, 263.05, 263.05, 263.05, 262.35, 
    262.45, 262.45, 262.45, 263.25, 263.25, 263.55, 263.95, 264.35, 264.35, 
    264.65, 265.05, 264.65, 264.55, 265.25, 266.05, 266.15, 267.35, 266.95, 
    266.55, 266.35, 266.95, 266.65, 266.15, 265.95, 265.75, 266.15, 268.05, 
    268.45, 268.45, 268.25, 265.85, 264.95, 264.25, 263.75, 262.95, 262.35, 
    261.65, 261.25, 260.65, 259.75, 258.95, 258.45, 258.05, 257.65, 256.95, 
    256.35, 256.05, 255.95, 256.05, 256.05, 256.45, 256.45, 256.55, 256.35, 
    256.05, 255.55, 255.25, 255.75, 256.65, 256.85, 257.55, 258.25, 259.45, 
    260.85, 260.95, 260.15, 259.85, 259.95, 259.75, 259.15, 259.15, 259.45, 
    259.95, 260.35, 260.55, 261.15, 260.35, 261.15, 260.85, 261.35, 261.05, 
    260.95, 261.15, 260.85, 259.95, 259.55, 260.25, 261.05, 262.05, 262.15, 
    262.25, 261.95, 261.95, 261.55, 261.95, 262.25, 262.45, 263.05, 263.65, 
    263.95, 264.25, 264.05, 263.85, 263.65, 263.25, 262.15, 260.25, 260.05, 
    259.45, 259.55, 259.15, 258.45, 257.85, 257.25, 257.15, 256.35, 257.35, 
    257.45, 256.45, 255.65, 254.65, 253.75, 253.35, 253.65, 253.55, 252.55, 
    251.35, 250.95, 250.85, 251.55, 251.25, 251.55, 251.95, 251.25, 251.35, 
    251.65, 252.15, 253.15, 254.05, 253.45, 254.15, 254.45, 254.95, 255.25, 
    256.55, 253.95, 251.85, 249.45, 248.25, 247.95, 247.45, 247.35, 247.25, 
    246.65, 245.05, 245.75, 245.55, 245.65, 245.45, 244.85, 244.45, 243.55, 
    243.25, 243.25, 243.45, 243.55, 243.45, 242.75, 241.45, 240.15, 239.55, 
    239.45, 239.45, 239.55, 239.95, 239.95, 240.15, 241.05, 241.35, 241.85, 
    243.05, 243.25, 243.95, 244.65, 245.25, 245.05, 245.15, 245.15, 245.35, 
    245.65, 245.65, 245.95, 246.25, 246.25, 245.95, 245.55, 245.85, 246.15, 
    246.25, 246.85, 246.95, 245.85, 244.35, 244.25, 244.55, 244.75, 245.35, 
    245.75, 246.05, 246.15, 246.35, 246.85, 247.05, 247.15, 247.35, 247.95, 
    248.45, 249.05, 250.35, 249.85, 249.55, 249.15, 249.15, 249.25, 248.65, 
    248.55, 248.15, 248.05, 248.35, 248.05, 247.65, 247.75, 247.85, 248.35, 
    248.75, 251.95, 253.05, 254.35, 254.85, 255.55, 256.15, 256.25, 255.95, 
    255.35, 252.55, 251.85, 251.95, 251.85, 251.65, 251.75, 251.95, 251.95, 
    252.45, 253.55, 255.05, 255.75, 256.35, 256.05, 256.15, 256.95, 257.05, 
    256.65, 256.65, 256.55, 256.55, 256.35, 255.85, 255.55, 255.65, 255.45, 
    255.55, 255.05, 254.65, 254.35, 254.45, 255.75, 256.05, 256.15, 255.25, 
    255.45, 256.15, 257.25, 257.25, 257.95, 257.85, 258.85, 259.75, 260.95, 
    261.75, 262.15, 262.75, 264.35, 265.65, 266.45, 267.45, 268.45, 269.05, 
    269.35, 269.15, 267.75, 266.45, 264.95, 264.55, 263.75, 263.55, 263.95, 
    263.45, 263.25, 263.15, 264.45, 264.55, 265.05, 264.75, 264.05, 264.65, 
    264.25, 263.65, 264.05, 263.75, 263.75, 263.65, 261.55, 260.65, 261.05, 
    261.15, 261.35, 260.25, 259.45, 258.85, 258.25, 258.45, 257.15, 255.95, 
    256.65, 256.85, 257.55, 256.35, 256.65, 255.45, 255.55, 255.25, 256.15, 
    256.45, 255.35, 256.35, 256.85, 256.65, 256.05, 255.95, 256.25, 256.55, 
    256.15, 255.55, 256.75, 254.85, 253.55, 251.05, 249.15, 247.25, 246.05, 
    245.65, 245.25, 244.55, 243.75, 243.45, 243.55, 243.25, 243.75, 244.25, 
    244.55, 244.95, 245.15, 245.25, 246.25, 246.55, 247.05, 247.25, 247.65, 
    247.45, 247.95, 247.75, 247.75, 247.45, 248.65, 250.25, 250.55, 251.25, 
    250.65, 250.95, 252.05, 251.35, 251.35, 251.25, 251.35, 251.65, 251.65, 
    251.45, 251.05, 251.55, 251.55, 251.55, 249.65, 249.35, 248.95, 248.75, 
    248.35, 248.05, 247.75, 248.25, 248.05, 248.45, 248.45, 248.05, 247.85, 
    248.35, 248.55, 248.35, 248.45, 248.05, 248.25, 248.35, 248.45, 248.65, 
    248.65, 248.65, 249.85, 249.75, 249.65, 249.45, 248.95, 248.75, 248.65, 
    249.45, 249.65, 249.35, 249.75, 249.95, 249.85, 249.45, 249.65, 249.85, 
    249.45, 249.05, 248.75, 248.55, 248.25, 248.15, 248.15, 248.15, 247.55, 
    247.55, 247.65, 247.45, 247.65, 247.15, 247.75, 247.45, 248.15, 247.95, 
    248.05, 248.95, 249.35, 249.05, 248.75, 249.65, 249.65, 249.05, 248.95, 
    249.65, 248.75, 250.45, 250.65, 252.45, 252.05, 252.65, 252.05, 251.65, 
    251.65, 251.15, 250.65, 250.05, 249.45, 248.95, 248.65, 248.65, 248.15, 
    247.75, 248.25, 248.25, 248.15, 248.55, 249.15 ;

 air_pressure_at_sea_level_qnh = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 99880, 99820, 99780, 99780, 100290, 
    100380, 100460, 100460, 100410, 100440, 100490, 100660, 100760, 101010, 
    101020, 101080, 101070, 100960, 100940, 100960, 100920, 100790, 100760, 
    100920, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    100730, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    100830, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    101180, 101190, 101250, 101280, 101310, 101310, 101310, 101300, 101270, 
    101240, 101200, 101210, 101160, 101110, 101140, 101120, 101120, 101100, 
    101070, 101050, 101030, 101010, 101000, 100990, 100990, 101020, 101050, 
    101120, 101140, 101160, 101150, 101150, 101150, 101160, 101200, 101240, 
    101240, 101240, 101270, 101300, 101390, _, _, _, _, _, _, _, _, _, 
    101560, 101600, 101640, 101690, 101750, 101770, 101780, 101820, 101800, 
    101840, 101920, 101950, 102020, 102110, 102190, 102240, 102310, 102350, 
    102410, 102440, 102460, 102470, 102480, 102500, _, 102650, 102690, 
    102780, 102820, 102890, 102870, 102920, 102950, 102950, 102960, 103010, 
    103040, 103100, 103100, 103130, 103140, 103160, 103180, 103160, 103170, 
    103150, 103180, 103200, 103250, 103280, 103300, 103300, 103290, 103300, 
    103310, 103320, 103330, 103370, 103410, 103440, 103480, 103490, 103520, 
    103520, 103540, 103570, 103620, 103660, 103710, 103740, 103770, 103810, 
    103840, 103900, 103940, 103960, 103960, 103960, 103960, 103990, 103980, 
    103980, 103990, 103990, 103930, 103900, 103970, 103980, 103940, 103920, 
    103880, 103820, 103790, 103630, 103650, 103610, 103630, 103640, 103650, 
    103640, 103620, 103620, 103630, 103640, 103650, 103660, 103670, 103670, 
    103670, 103660, 103690, 103660, 103640, 103630, 103650, 103680, 103690, 
    103680, 103710, 103730, 103740, 103770, 103760, 103770, 103810, 103820, 
    103850, 103840, 103860, 103850, 103840, 103790, 103790, 103790, 103800, 
    103790, 103770, 103750, 103750, 103730, 103720, 103730, 103740, 103740, 
    103760, 103760, 103770, 103760, 103760, 103780, 103790, 103810, 103830, 
    103820, 103820, 103850, 103880, 103890, 103940, 103960, 104010, 104010, 
    104000, 104030, 104020, 104040, 104030, 104040, _, 104090, 104110, 
    104140, 104130, 104110, 104100, 104080, 104040, 104000, 103970, 103940, 
    103910, 103880, 103840, 103790, 103760, 103720, 103670, 103630, 103590, 
    103560, 103510, 103450, 103380, 103350, 103310, 103290, 103230, 103180, 
    103130, 103070, 103060, 103030, 103000, 102970, 102950, 102960, 102910, 
    102900, 102860, 102830, 102780, 102770, 102730, 102690, 102680, 102660, 
    102700, 102700, 102680, 102690, 102690, 102680, 102650, 102630, 102600, 
    102590, 102580, 102570, 102560, 102590, 102590, 102590, 102560, 102530, 
    102500, 102460, 102460, 102460, 102460, 102460, 102460, 102460, 102470, 
    102460, 102420, 102430, 102400, 102380, 102340, 102330, 102310, 102300, 
    102280, 102290, 102270, 102220, 102200, 102170, 102140, 102110, 102110, 
    102100, 102050, 102030, 102030, 102030, 102020, 102020, 101970, 101920, 
    101850, 101780, 101720, 101670, 101640, 101590, 101540, 101510, 101490, 
    101480, 101440, 101430, 101400, 101370, 101350, 101360, 101360, 101380, 
    101410, 101390, 101370, 101380, 101410, 101390, 101370, 101360, 101330, 
    101320, 101280, 101270, 101270, 101240, 101190, 101170, 101100, 101060, 
    101020, 101000, 100990, 100970, 100990, 100980, 100990, 101050, 101080, 
    101150, 101140, 101160, 101160, 101210, 101240, 101280, 101300, 101320, 
    101360, 101380, 101410, 101440, 101470, 101470, 101510, 101460, 101530, 
    101550, 101560, 101620, 101670, 101740, 101800, 101800, 101830, 101870, 
    101910, 101950, 101980, 102060, 102130, 102210, 102280, 102370, 102370, 
    102430, 102470, 102540, 102590, 102640, 102710, 102790, 102890, 102970, 
    103030, 103100, 103150, 103190, 103220, 103260, 103310, 103370, 103410, 
    103470, 103500, 103520, 103570, 103600, 103600, 103600, 103560, 103490, 
    103400, 103390, 103330, 103240, 103160, 103060, 102920, 102840, 102680, 
    102500, 102380, 102320, 102290, 102290, 102300, 102320, 102340, 102330, 
    102340, 102320, 102330, 102340, 102310, 102290, 102340, 102390, 102380, 
    102400, 102460, 102510, 102550, 102610, 102680, 102710, 102760, 102800, 
    102780, 102810, 102830, 102880, 102870, 102880, 102920, 102960, 102960, 
    102970, 103010, 103010, 103010, 102990, 103030, 103010, 103090, 103130, 
    103210, 103250, 103310, 103350, 103410, 103430, 103440, 103430, 103450, 
    103480, 103480, 103490, 103500, 103500, 103500, 103500, 103470, 103420, 
    103370, 103380, 103340, 103280, 103220, 103190, 103150, 103120, 103090, 
    103060, 102990, 102920, 102860, 102730, 102680, 102660, 102600, 102540, 
    102490, 102470, 102400, 102360, 102300, 102280, 102250, 102220, 102190, 
    102150, 102130, 102090, 102100, 102100, 102080, 102040, 102010, 102010, 
    101960, 101920, 101890, 101890, 101870, 101870, 101890, 101870, 101870, 
    101860, 101870, 101900, 101910, 101940, 101950, 101980, 101980, 102020, 
    102060, 102100, 102100, 102120, 102140, 102140, 102110, 102060, 102040, 
    101990, 101930, 101890, 101850, 101770, 101650, 101540, 101430, 101420, 
    101380, 101300, 101230, 101190, 101130, 101040, 100940, 100860, 100830, 
    100750, 100630, 100560, 100500, 100430, 100360, 100300, 100270, 100260, 
    100240, 100230, 100220, 100230, 100230, 100230, 100200, 100170, 100120, 
    100140, 100170, 100210, 100280, 100300, 100420, 100670, 100790, 100950, 
    101070, 101230, 101340, 101430, 101590, 101680, 101790, 101870, 101970, 
    102020, 102050, 102090, 102110, 102150, 102160, 102200, 102260, 102310, 
    102370, 102440, 102490, 102540, 102620, 102670, 102760, 102830, 102900, 
    102950, 103000, 103060, 103100, 103160, 103200, 103220, 103240, 103230, 
    103250, 103230, 103220, 103160, 103060, 102990, 102910, 102810, 102680, 
    102570, 102430, 102260, 102070, 101840, 101690, 101520, 101350, 101150, 
    101140, 101100, 101060, 101090, 101170, 101230, 101220, _, 101400, 
    101540, 101700, 101830, 102010, 102150, 102280, 102410, 102470, 102530, 
    102660, 102710, 102780, 102840, 102890, 102910, 102940, 102960, 102940, 
    102930, 102930, 102960, 102970, 102980, 103000, 103040, 103040, 103060, 
    103110, 103140, 103160, 103190, 103180, 103210, 103240, 103200, 103080, 
    103070, 102920, 102840, 102720, 102560, 102410, 102230, 101910, 101610, 
    101370, 101170, 100980, 100730, 100350, 100170, 100100, 100040, 99990, 
    99940, 99840, 99780, 99710, 99620, 99570, 99540, 99560, 99510, 99460, 
    99370, 99290, 99250, 99240, 99270, 99270, 99290, 99370, 99710, 100000, 
    100240, 100530, 100730, 100930, 101150, 101270, 101320, 101380, 101710, 
    101900, 101840, 102000, 102140, 102240, 102280, 102330, 102330, 102320, 
    102360, 102340, 102320, 102290, 102230, 102170, 102120, 102050, 101980, 
    101880, 101750, 101630, 101480, 101330, 101150, 101000, 100820, 100680, 
    100590, 100510, 100440, 100390, 100270, 100190, 100090, 99990, 99900, 
    99790, 99680, 99570, 99490, 99420, 99380, 99340, 99320, 99290, 99260, 
    99260, 99240, 99290, 99300, 99310, 99310, 99370, 99420, 99450, 99470, 
    99470, 99470, 99460, 99430, 99440, 99420, 99410, 99420, 99460, 99460, 
    99490, 99540, 99510, 99510, 99540, 99500, 99470, 99430, 99360, 99300, 
    99280, 99300, 99300, 99250, 99180, 99110, 99020, 98940, 98720, 98490, 
    98320, 97810, 97690, 97640, 97560, 97450, 97460, 97490, 97720, 97980, 
    98360, 98550, 98700, 98880, 99000, 99100, 99170, 99200, 99210, 99250, 
    99300, 99320, 99350, 99390, 99430, 99430, 99510, 99570, 99620, 99650, 
    99640, 99670, 99710, 99780, 99850, 99900, 99950, 100010, 100070, 100120, 
    100190, 100250, 100320, 100370, 100410, 100510, 100550, 100600, 100670, 
    100750, 100750, 100790, 100800, 100790, 100620, 100590, 100610, 100630, 
    100620, 100640, 100660, 100700, 100720, 100790, 100830, 100840, 100810, 
    100780, 100800, 100790, 100800, 100780, 100820, 100770, 100810, 100790, 
    100790, 100770, 100770, 100730, 100720, 100710, 100660, 100850, 100890, 
    100920, 100980, 101030, 101080, 101110, 101150, 101180, 101170, 101170, 
    101190, 101180, 101190, 101170, 101190, 101180, 101220, 101210, 101210, 
    101180, 101110, 101090, 101100, 101110, 101110, 101150, 101130, 101130, 
    101130, 101140, 101140, 101150, 101180, 101180, 101180, 101200, 101220, 
    101190, 101160, 101140, 101170, 101100, 101110, 101130, 101130, 101080, 
    101080, 101020, 100990, 100970, 100970, 100930, 100950, 100930, 100890, 
    100890, 100910, 100920, 100900, 100870, 100890, 100840, 100810, 100820, 
    100770, 100740, 100730, 100720, 100710, 100690, 100700, 100740, 100720, 
    100760, 100740, 100740, 100740, 100720, 100680, 100690, 100670, 100620, 
    100580, 100530, 100490, 100450, 100490, 100480, 100500, 100460, 100380, 
    100390, 100380, 100300, 100270, 100260, 100200, 100110, 100020, 99960, 
    100000, 99940, 99910, 99840, 99880, 99870, 99880, 99920, 99880, 99930, 
    99970, 100060, 100060, 100090, 100130, 100210, 100270, 100280, 100320, 
    100330, 100360, 100400, 100460, 100450, 100430, 100470, 100490, 100530, 
    _, 100600, 100630, 100650, 100680, 100730, 100770, 100810, 100840, 
    100860, 100850, 100890, 100900, 100970, 100980, 101040, 101090, 101150, 
    101200, 101270, 101330, 101360, 101400, 101460, 101500, 101560, 101610, 
    101640, 101670, 101730, 101790, 101850, 101900, 101910, 101940, 101970, 
    101960, 101970, 101960, 101910, 101890, 101890, 101860, 101830, 101780, 
    101740, 101670, 101610, 101550, 101450, 101310, 101180, 101090, 101000, 
    100900, 100790, 100730, 100640, 100510, 100370, 100300, 100220, 100150, 
    100070, 99980, 99920, 99790, 99720, 99630, 99560, 99510, 99460, 99380, 
    99300, 99240, 99190, 99180, 99120, 99090, 99080, 99120, 99190, 99250, 
    99300, 99350, 99370, 99410, 99430, 99430, 99450, 99470, 99470, 99460, 
    99450, 99450, 99500, 99540, 99540, 99550, 99530, 99550, 99570, 99610, 
    99680, 99770, 99820, 99870, 99960, 100050, 100110, 100170, 100210, 
    100270, 100340, 100400, 100470, 100530, 100580, 100650, 100690, 100750, 
    100780, 100820, 100850, 100930, 101000, 101040, 101090, 101130, 101140, 
    101180, 101180, 101190, 101210, 101190, 101150, 101110, 101080, 101030, 
    101050, 101040, 101010, 100980, 100950, 100890, 100880, 100820, 100770, 
    100750, 100680, 100620, 100580, 100560, 100430, 100300, 100220, 100100, 
    100020, 99940, 99850, 99810, 99760, 99730, 99680, 99580, 99430, 99310, 
    99150, 99000, 98920, 98760, 98710, 98700, 98760, 98810, 98880, 98950, 
    99030, 99090, 99130, 99150, 99230, 99280, 99340, 99500, 99630, 99800, 
    99990, 100120, 100210, 100230, 100290, 100310, 100370, 100410, 100460, 
    100490, 100520, 100560, 100580, 100560, 100530, 100550, 100580, 100560, 
    100600, 100620, 100650, 100690, 100680, 100710, 100710, 100730, 100590, 
    100680, 100700, _, 100820, 100910, 100880, 100870, 100920, 100970, 
    101020, 101080, 101130, 101120, 101170, 101210, 101260, 101310, 101380, 
    101420, 101470, 101540, 101580, 101630, 101700, 101750, 101790, 101830, 
    101860, 101900, 101930, 101960, 101990, 102040, 102110, 102140, 102170, 
    102190, 102200, 102220, 102240, 102260, 102280, 102280, 102280, 102270, 
    102270, 102280, 102280, 102290, 102300, 102290, 102280, 102230, 102230, 
    102200, 102210, 102210, 102210, 102210, 102200, 102190, 102150, 102100, 
    102080, 102070, 102050, 102020, 101990, 101930, 101890, 101850, 101820, 
    101780, 101730, 101680, 101630, 101550, 101460, 101400, 101310, 101320, 
    101210, 101210, 101180, 101140, 101080, 101020, 100990, 100890, 100850, 
    100830, 100720, 100750, 100710, 100680, 100630, 100620, 100580, 100650, 
    100650, 100680, 100700, 100710, 100690, 100590, 100570, 100460, 100470, 
    100450, 100420, 100410, 100430, 100420, 100530, 100480, 100510, 100580, 
    100630, 100590, 100600, 100640, 100600, 100660, 100720, 100710, 100700, 
    100720, 100660, 100680, 100630, 100530, 100540, 100620, 100730, 100770, 
    100870, 100970, 101110, 101130, 101260, 101340, 101470, 101520, 101580, 
    101650, 101680, 101730, 101740, 101750, 101760, 101780, 101800, 101800, 
    101810, 101830, 101860, 101840, 101830, 101830, 101810, 101820, 101800, 
    101750, 101700, 101710, 101670, 101560, 101530, 101440, 101380, 101310, 
    101200, 101090, 101020, 100910, 100810, 100730, 100690, 100570, 100500, 
    100390, 100300, 100210, 100160, 100060, 100040, 100020, 99990, 100100, 
    100120, 100210, 100270, 100290, 100330, 100460, 100520, 100560, 100740, 
    100730, 100740, 100760, 100810, 100890, 100910, 100930, 100950, 101010, 
    101060, 101070, 101100, 101170, 101170, 101190, 101240, 101250, 101250, 
    101200, 101220, 101210, 101240, 101210, 101200, 101210, 101260, 101260, 
    101230, 101230, 101260, 101250, 101230, 101210, 101240, 101240, 101250, 
    101240, 101280, 101270, 101300, 101380, 101500, 101560, 101710, 101720, 
    101810, 101830, 101980, 102000, 101990, 101990, 102180, 102310, 102330, 
    102390, 102410, 102420, 102410, 102380, 102390, 102400, 102390, 102340, 
    102280, 102320, 102290, 102270, 102250, 102170, 102150, 102100, 102090, 
    102040, 101980, 101910, 101850, 101770, 101690, 101620, 101550, 101500, 
    101500, 101520, 101550, 101560, 101530, 101580, 101580, 101560, 101540, 
    101510, 101480, 101450, 101400, 101370, 101330, 101300, 101280, 101260, 
    101240, 101220, 101160, 101130, 101130, 101150, 101150, 101140, 101130, 
    101130, 101130, 101160, 101150, 101130, 101120, 101110, 101090, 101080, 
    101100, 101090, 101090, 101040, 101030, 101020, 101080, 101090, 101070, 
    101060, 101030, 101020, 101000, 100990, 100970, 100930, 100910, 100870, 
    100870, 100860, 100870, 100870, 100850, 100840, 100860, 100860, 100860, 
    100860, 100850, 100860, 100880, 100890, 100880, 100880, 100860, 100850, 
    100830, 100850, 100810, 100810, 100800, 100800, 100800, 100800, 100810, 
    100780, 100760, 100770, 100750, 100740, 100750, 100760, 100780, 100760, 
    100770, 100790, 100810, 100830, 100840, 100860, 100860, 100870, 100900, 
    100910, 100910, 100920, 100960, 100960, 100970, 100970, 100970, 100980, 
    100960, 100980, 100960, 100950, 100940, 100950, 100970, 101000, 101010, 
    101010, 101000, 101010, 101000, 100980, 100970, 100970, 100960, 100940, 
    100910, 100890, 100870, 100840, 100840, 100790, 100780, 100730, 100670, 
    100630, 100580, 100550, 100500, 100500, 100460, 100590, 100410, 100480, 
    100550, 100530, 100500, 100470, 100440, 100420, 100420, 100340, 100300, 
    100260, 100230, 100270, 100280, 100330, 100220, 100250, 100280, 100320, 
    100440, 100510, 100560, 100560, 100570, 100570, 100600, 100610, 100620, 
    100630, 100670, 100680, 100670, 100670, 100660, 100650, 100560, 100580, 
    100590, 100650, 100610, 100600, 100630, 100650, 100640, 100640, 100640, 
    100630, 100610, 100600, 100590, 100590, 100580, 100580, 100570, 100540, 
    100560, 100560, 100560, 100520, 100510, 100500, 100500, 100460, 100450, 
    100500, 100500, 100520, 100530, 100510, 100500, 100600, 100530, 100540, 
    100540, 100520, 100520, 100490, 100480, 100480, 100460, 100410, 100360, 
    100330, 100230, 100320, 100400, 100380, 100360, 100350, 100370, 100300, 
    100380, 100340, 100270, 100280, 100310, 100300, 100260, 100260, 100240, 
    100250, 100250, 100280, 100310, 100330, 100330, 100330, 100340, 100360, 
    100380, 100390, 100440, 100440, 100440, 100480, 100490, 100520, 100470, 
    100460, 100470, 100500, 100500, 100520, 100530, 100560, 100600, 100620, 
    100640, 100680, 100710, 100700, 100700, 100690, 100770, 100840, 100880, 
    100930, 100970, 101030, 101070, 101130, 101170, 101180, 101220, 101260, 
    101300, 101340, 101380, 101410, 101460, 101490, 101510, 101550, 101590, 
    101620, 101640, 101660, 101690, 101720, 101740, 101750, 101760, 101780, 
    101810, 101820, 101820, 101810, 101810, 101800, 101820, 101810, 101790, 
    101790, 101750, 101740, 101740, 101730, 101690, 101670, 101660, 101670, 
    101640, 101640, 101610, 101600, 101600, 101600, 101590, 101590, 101600, 
    101600, 101600, 101560, 101530, 101560, 101530, 101520, 101500, 101490, 
    101490, 101500, 101490, 101490, 101460, 101450, 101440, 101450, 101450, 
    101430, 101420, 101430, 101460, 101450, 101440, 101430, 101400, 101400, 
    101410, 101400, 101410, 101420, 101380, 101400, 101380, 101360, 101360, 
    101310, 101280, 101300, 101300, 101260, 101240, 101230, 101210, 101220, 
    101190, 101190, 101190, 101180, 101170, 101170, 101170, 101150, 101130, 
    101080, 101080, 101090, 101100, 101130, 101130, 101130, 101150, 101140, 
    101150, 101190, 101180, 101190, 101230, 101250, 101270, 101290, 101290, 
    101260, 101200, 101090, 101040, 100930, 100880, 100850, 100760, 100680, 
    100770, 100810, 100870, 100900, 100920, 101000, 101090, 101150, 101240, 
    101350, 101410, 101530, 101560, 101580, 101650, 101660, 101660, 101660, 
    101690, 101690, 101680, 101640, 101660, 101660, 101660, 101660, 101740, 
    101780, 101870, 101990, 102010, 102050, 102110, 102150, 102190, 102220, 
    102250, 102260, 102290, 102310, 102330, 102350, 102380, 102390, 102420, 
    102430, 102440, 102420, 102410, 102370, 102350, 102340, 102290, 102280, 
    102200, 102160, 102110, 102060, 102040, 102080, 102080, 102040, 102060, 
    102060, 102070, 102050, 102040, 102020, 102010, 101990, 101980, 101970, 
    101960, 101930, 101930, 101900, 101880, 101830, 101760, 101730, 101610, 
    101530, 101450, 101420, 101360, 101320, 101260, 101210, 101100, 101040, 
    100950, 100870, 100770, 100670, 100600, 100520, 100480, 100450, 100470, 
    100420, 100390, 100360, 100360, 100370, 100450, 100520, 100590, 100640, 
    100700, 100740, 100770, 100830, 100850, 100910, 100880, 100890, 100970, 
    101060, 101160, 101230, 101310, 101370, 101490, 101560, 101630, 101700, 
    101760, 101850, 101880, 101930, 101950, 102000, 102050, 102080, 102100, 
    102130, 102150, 102130, 102130, 102120, 102110, 102110, 102090, 102080, 
    102110, 102110, 102060, 102030, 102020, 101960, 101950, 101910, 101860, 
    101870, 101860, 101820, 101790, 101780, 101740, 101700, 101650, 101600, 
    101580, 101530, 101490, 101500, 101530, 101580, 101610, 101610, 101750, 
    101860, 101940, 102020, 102050, 102060, 102120, 102210, 102270, 102310, 
    102320, 102330, 102450, 102520, 102610, 102650, 102650, 102740, 102740, 
    102760, 102760, 102730, 102710, 102660, 102600, 102550, 102500, 102360, 
    102310, 102250, 102180, 102120, 102050, 102000, 101980, 101970, 102030, 
    102060, 102100, 102160, 102240, 102290, 102320, 102310, 102330, 102330, 
    102330, 102300, 102250, 102220, 102170, 102120, 102080, 102020, 101960, 
    101910, 101860, 101790, 101730, 101680, 101600, 101550, 101510, 101470, 
    101450, 101450, 101480, 101530, 101560, 101590, 101660, 101620, 101730, 
    101770, 101790, 101840, 101870, 101900, 101910, 101960, 101990, 102010, 
    102050, 102060, 102130, 102180, 102180, 102250, 102260, 102260, 102330, 
    102400, 102400, 102430, 102520, 102510, 102520, 102510, 102510, 102500, 
    102560, 102550, 102480, 102410, 102430, 102460, 102460, 102400, 102390, 
    102350, 102300, 102270, 102210, 102200, 102120, 102090, 102070, 102020, 
    101990, 101950, 101880, 101800, 101740, 101680, 101620, 101530, 101460, 
    101420, 101400, 101390, 101390, 101350, 101390, 101400, 101450, 101430, 
    101420, 101380, 101380, 101360, 101350, 101340, 101330, 101340, 101340, 
    101360, 101310, 101280, 101230, 101210, 101170, 101140, 101180, 101150, 
    101180, 101280, 101310, 101310, 101370, 101440, 101500, 101520, 101530, 
    101610, 101710, 101750, 101790, 101820, 101820, 101820, 101790, 101800, 
    101790, 101750, 101700, 101690, 101630, 101570, 101540, 101520, 101470, 
    101420, 101370, 101320, 101270, 101250, 101220, 101190, 101160, 101160, 
    101160, 101160, 101190, 101240, 101270, 101310, 101360, 101390, 101430, 
    101470, 101520, 101620, 101700, 101770, 101830, 101910, 102000, 102050, 
    102120, 102180, 102210, 102250, 102300, 102340, 102390, 102420, 102460, 
    102490, 102480, 102500, 102500, 102510, 102490, 102480, 102460, 102490, 
    102500, 102540, 102530, 102540, 102550, 102550, 102550, 102520, 102510, 
    102500, 102480, 102490, 102510, 102520, 102500, 102500, 102480, 102460, 
    102440, 102420, 102380, 102350, 102310, 102310, 102300, 102290, 102260, 
    102280, 102250, 102250, 102240, 102250, 102230, 102220, 102230, 102230, 
    102220, 102200, 102200, 102190, 102120, 102150, 102160, 102150, 102140, 
    102130, 102160, 102160, 102180, 102170, _, 102160, 102140, 102130, 
    102120, 102110, 102070, 102050, 102050, 102050, _, 102010, 101970, 
    101960, 101930, 101910, 101890, 101870, 101840, 101840, 101850, 101840, 
    101860, 101840, 101830, 101850, 101840, 101820, 101790, 101790, 101770, 
    101760, 101750, 101700, 101700, _, 101650, 101650, 101630, 101630, 
    101630, 101610, 101570, 101570, 101600, 101660, 101750, 101820, 101880, 
    101910, 101950, 101910, 101940, 101890, 101950, 101920, 101820, 101800, 
    101800, 101820, 101810, 101790, 101710, 101690, 101680, 101640, 101610, 
    _, 101550, 101630, 101660, 101740, 101680, 101710, 101700, 101670, 
    101670, 101720, 101630, 101640, 101760, 101750, 101680, _, 101710, 
    101790, 101840, 101890, 101970, 102040, 102140, 102160, 102180, 102250, 
    102370, 102480, 102530, 102590, 102690, 102760, 102830, 102860, 102890, 
    102910, 102910, 102960, 103000, 102950, 102890, 102850, 102870, 102850, 
    102790, 102780, 102800, 102800, 102830, 102810, 102770, 102800, 102740, 
    102660, 102640, 102620, 102610, 102550, 102560, 102530, 102530, 102580, 
    102560, 102530, 102530, 102530, 102510, 102520, 102510, 102550, 102560, 
    102570, 102590, 102630, 102650, 102700, 102700, 102730, 102760, 102740, 
    102740, 102740, 102760, 102790, 102800, 102830, 102830, 102820, 102840, 
    102830, 102790, 102720, 102710, 102610, 102600, 102580, 102500, 102430, 
    102350, 102270, 102220, 102130, 102160, 102070, 102160, 102110, 102060, 
    102010, 102030, 102010, 101990, 102000, 101930, 101940, 101940, 101970, 
    102020, 102060, 102040, 102040, 102000, 102090, 102160, 102210, 102210, 
    102200, 102190, 102250, 102220, 102180, 102180, 102180, 102160, 102170, 
    102130, 102080, 102150, 102160, 102130, 102220, 102190, 102260, 102320, 
    102370, 102400, 102450, 102520, 102570, 102580, 102610, 102620, 102640, 
    102660, 102660, 102630, 102680, 102690, 102700, 102720, 102720, 102730, 
    102680, 102680, 102650, 102630, 102580, 102600, 102630, 102570, 102470, 
    102470, 102600, 102500, 102580, 102580, 102540, 102540, 102460, 102350, 
    102360, 102350, 102320, 102380, 102330, 102360, 102340, 102300, 102270, 
    102270, 102290, 102330, 102290, 102290, 102280, 102320, 102290, 102290, 
    102240, 102200, 102190, 102150, 102100, 102030, 101990, 101900, 101830, 
    101770, 101720, 101690, 101650, 101600, 101530, 101550, 101540, 101490, 
    101440, 101440, 101430, 101390, 101330, 101320, 101270, 101240, 101200, 
    101170, 101160, 101140, 101130, 101060, 101060, 101050, 100980, 100960, 
    100920, 100880, 100820, 100750, 100690, 100680, 100620, 100570, 100560, 
    100560, 100530, 100490, 100470, 100450, 100450, 100450, 100460, 100480, 
    100510, 100530, 100580, 100620, 100670, 100710, 100780, 100840, 100890, 
    100940, 101010, 101070, 101120, 101180, 101250, 101300, 101350, 101390, 
    101450, 101480, 101520, 101530, 101530, 101520, 101580, 101590, 101630, 
    101670, 101680, 101750, 101730, 101760, 101810, 101850, 101910, 101830, 
    101830, 101860, 101920, 101950, 101960, 101970, 101980, 102000, 102110, 
    102200, 102290, 102370, 102480, 102540, 102660, 102710, 102770, 102830, 
    102890, 102940, 103030, 103090, 103160, 103250, 103310, 103330, 103400, 
    103490, 103540, 103590, 103620, 103640, 103660, 103740, 103810, 103880, 
    103980, 104090, 104150, 104220, 104240, 104330, 104410, 104480, 104540, 
    104600, 104620, 104670, 104700, 104720, 104750, 104840, 104880, 104910, 
    104890, 104950, 104950, 104980, 105020, 105070, 105090, 105140, 105110, 
    105140, 105140, 105140, 105250, 105020, 105050, 105080, 104950, 104990, 
    105100, 105130, 105190, 105270, 105300, 105320, 105330, 105370, 105400, 
    105390, 105410, 105400, 105420, 105470, 105520, 105590, 105660, 105700, 
    105750, 105780, 105790, 105830, 105880, 105890, 105910, 105930, 105920, 
    105950, 105970, 106010, 106010, 106000, 106010, 106000, 106000, 105970, 
    105930, 105900, 105870, 105830, 105780, 105720, 105650, 105600, 105520, 
    105450, 105370, 105290, 105190, 105120, 105060, 105020, 104970, 104960, 
    104880, 104790, 104680, 104710, 104550, 104460, 104320, 104270, 104220, 
    104170, 104210, 104130, 104120, 104060, 103980, 103850, 103790, 103750, 
    103690, 103590, 103460, 103430, 103400, 103360, 103330, 103320, 103320, 
    103300, 103280, 103280, 103270, 103260, 103240, 103270, 103270, 103290, 
    103260, 103270, 103220, 103220, 103240, 103210, 103180, 103160, 103210, 
    103230, 103190, 103200, 103190, 103210, 103210, 103180, 103150, 103130, 
    103090, 103050, 103020, 103010, 103000, 102990, 102970, 102960, 102960, 
    102930, 102930, 102920, 102930, 102930, 102940, 103000, 103020, 103060, 
    103060, 103060, 103080, 103090, 103110, 103120, 103120, 103120, 103130, 
    103140, 103140, 103120, 103100, 103100, 103080, 103060, 103020, 103010, 
    102920, 102870, 102920, 102850, 102770, 102730, 102610, 102560, 102540, 
    102560, 102600, 102590, 102590, 102540, 102550, 102570, 102580, 102580, 
    102570, 102570, 102430, 102390, 102430, 102490, 102530, 102530, 102520, 
    102590, 102580, 102600, 102590, 102520, 102430, 102210, 102160, 102090, 
    102150, 102110, 102080, 102150, 102190, 102160, 102150, 102190, 102180, 
    102280, 102280, 102170, 102150, 102170, 102220, 102280, 102250, 102310, 
    102300, 102350, 102380, 102370, 102350, 102340, 102310, 102230, 102170, 
    102190, 102220, 102250, 102220, 102240, 102180, 102240, 102280, 102290, 
    102270, 102300, 102330, 102350, 102370, 102360, 102350, 102340, 102320, 
    102300, 102280, 102270, 102260, 102260, 102230, 102230, 102210, 102180, 
    102150, 102150, 102120, 102080, 102060, 102050, 102050, 102030, 102010, 
    102000, 101970, 101970, 101910, 101860, 101810, 101780, 101750, 101680, 
    101620, 101560, 101520, 101480, 101450, 101450, 101430, 101400, 101390, 
    101360, 101340, 101310, 101290, 101250, 101210, 101150, 101140, 101110, 
    101040, 100960, 100930, 100870, 100830, 100740, 100640, 100630, 100620, 
    100610, 100550, 100510, 100480, 100430, 100410, 100360, 100320, 100300, 
    100260, 100220, 100180, 100190, 100180, 100130, 100060, 100080, 100080, 
    100090, 100110, 100140, 100140, 100140, 100080, 100110, 100150, 100170, 
    100180, 100160, 100130, 100170, 100200, 100230, 100230, 100210, 100170, 
    100170, 100200, 100210, 100190, 100210, 100180, 100290, 100330, 100420, 
    100510, 100600, 100690, 100820, 100910, 100980, 101060, 101130, 101230, 
    101280, 101310, 101350, 101400, 101440, 101450, 101470, 101570, 101620, 
    101620, 101660, 101620, 101600, 101800, 101820, 101860, 101800, 101840, 
    101830, 101910, 101910, 101890, 101900, 101910, 101870, 101880, 101840, 
    101810, 101810, 101790, 101650, 101760, 101730, 101710, 101690, 101760, 
    101810, 101760, 101770, 101790, 101850, 101960, 101990, 102040, 102090, 
    102060, 101990, 102020, 102060, 102040, 102110, 102120, 102130, 102200, 
    102230, 102250, 102240, 102290, 102290, 102340, 102380, 102430, 102440, 
    102460, 102440, 102320, 102440, 102480, 102530, 102500, 102470, 102390, 
    102310, 102280, 102310, 102390, 102390, 102400, 102400, 102340, 102380, 
    102420, 102490, 102530, 102560, 102540, 102550, 102560, 102530, 102540, 
    102560, 102490, 102500, 102470, 102410, 102400, 102400, 102370, 102320, 
    102230, 102210, 102170, 102110, 102070, 102000, 102010, 101980, 101920, 
    101830, 101790, 101720, 101730, 101750, 101770, 101680, 101680, 101620, 
    101590, 101610, 101660, 101630, 101610, 101570, 101560, 101550, 101480, 
    101500, 101440, 101560, 101520, 101500, 101500, 101480, 101430, 101450, 
    101430, 101350, 101320, 101290, 101260, 101220, 101160, 101120, 101090, 
    101020, 101030, 101000, 100990, 100970, 100990, 100960, 100980, 100960, 
    100920, 100910, 100910, 100900, 100870, 100840, 100830, 100830, 100820, 
    100830, 100780, 100780, 100770, 100770, 100780, 100720, 100720, 100720, 
    100690, 100710, 100740, 100740, 100710, 100710, 100690, 100650, 100630, 
    100640, 100620, 100600, 100590, 100600, 100610, 100560, 100560, 100540, 
    100520, 100510, 100470, 100490, 100500, 100460, 100460, 100450, 100450, 
    100470, 100480, 100460, 100530, 100540, 100530, 100600, 100580, 100580, 
    100620, 100640, 100710, 100760, 100740, 100790, 100870, 100910, 100920, 
    100930, 100970, 101030, 101060, 101110, 101080, 100940, 101270, 101330, 
    101330, 101320, _, 101410, 101400, 101450, 101450, 101500, 101550, 
    101590, 101600, 101610, 101640, 101660, 101640, 101650, 101640, 101640, 
    101650, 101670, 101670, 101680, 101660, 101630, 101630, 101620, 101620, 
    101590, 101570, 101570, 101560, 101560, 101540, 101560, 101560, 101550, 
    101520, 101500, 101510, 101500, 101500, 101480, 101470, 101470, 101490, 
    101500, 101510, 101510, 101500, 101490, 101500, 101470, 101460, 101480, 
    101470, 101460, 101460, 101420, 101400, 101370, 101330, 101300, 101260, 
    101250, 101210, 101180, 101150, 101080, 101060, 101010, 100990, 100950, 
    100920, 100870, 100860, 100850, 100820, 100830, 100790, 100800, 100810, 
    100810, 100790, 100800, 100780, 100770, 100770, 100770, 100800, 100810, 
    100800, 100840, 100850, 100850, 100870, 100850, 100840, 100840, 100810, 
    100810, 100840, 100900, 100930, 100980, 101020, 101060, 101090, 101130, 
    101170, 101200, 101220, 101230, 101250, 101270, 101320, 101340, 101370, 
    101380, 101410, 101410, 101410, 101410, 101410, 101380, 101370, 101370, 
    101360, 101360, 101330, 101280, 101240, 101240, 101210, 101170, 101100, 
    101070, 101040, 100980, 100940, 100920, 100870, 100830, 100760, 100770, 
    100750, 100730, 100650, 100610, 100620, 100570, 100580, 100560, 100520, 
    100490, 100480, 100480, 100440, 100440, 100390, 100400, 100440, 100460, 
    100460, 100450, 100450, 100440, 100420, 100440, 100470, 100450, 100480, 
    100500, 100490, 100480, 100510, 100510, 100520, 100540, 100540, 100540, 
    100560, 100570, 100580, 100560, 100580, 100610, 100610, 100640, 100640, 
    100670, 100690, 100710, 100720, 100730, 100790, 100810, 100840, 100870, 
    100970, 101000, 100960, 101000, 101010, 101030, 101040, 101080, 101120, 
    101130, 101200, 101220, 101250, 101290, 101330, 101350, 101410, 101460, 
    101470, 101510, 101540, 101600, 101580, 101620, 101660, 101670, 101680, 
    101680, 101740, 101740, 101790, 101820, 101870, 101870, 101930, 101960, 
    101990, 102020, 102060, 102100, 102090, 102080, 102050, 102030, 102000, 
    101970, 101930, 101890, 101860, 101810, 101740, 101680, 101650, 101580, 
    101490, 101420, 101300, 101220, 101050, 100960, 100910, 100850, 100810, 
    100740, 100690, 100660, 100580, 100550, 100520, 100510, 100480, 100480, 
    100430, 100340, 100300, 100280, 100180, 100080, 100040, 99990, 99940, 
    99880, 99830, 99780, 99730, 99710, 99670, 99640, 99590, 99590, 99530, 
    99540, 99560, 99580, 99610, 99670, 99740, 99800, 99820, 99840, 99860, 
    99870, 99830, 99830, 99820, 99780, 99750, 99740, 99730, 99730, 99690, 
    99670, 99620, 99570, 99540, 99540, 99510, 99530, 99560, 99590, 99630, 
    99660, 99700, 99720, 99770, 99820, 99850, 99840, 99870, 99860, 99910, 
    99930, 99950, 99950, 99980, 99960, 99970, 99990, 100030, 100070, 100080, 
    100110, 100120, 100150, 100180, 100230, 100250, 100290, 100350, 100380, 
    100440, 100470, 100480, 100510, 100530, 100560, 100550, 100560, 100590, 
    100590, 100580, 100580, 100580, 100580, 100560, 100530, 100510, 100490, 
    100490, 100480, 100480, 100460, 100470, 100470, 100480, 100530, 100570, 
    100590, 100590, 100640, 100680, 100720, 100770, 100790, 100850, 100910, 
    100940, 101000, 101060, 101060, 101070, 101140, 101170, 101220, 101240, 
    101300, 101330, 101380, 101410, 101440, 101460, 101450, 101460, 101470, 
    101410, 101430, 101420, 101420, 101380, 101260, 101260, 101270, 101230, 
    101090, 100990, 100860, 100810, 100860, 100870, 100840, 100790, 100770, 
    100730, 100700, 100690, 100670, 100610, 100610, 100580, 100560, 100590, 
    100620, 100680, 100730, 100790, 100830, 100860, 100890, 100900, 100920, 
    100940, 100960, 100960, 100990, 101080, 101120, 101120, 101140, 101170, 
    101180, 101210, 101240, 101250, 101280, 101310, 101340, 101370, 101400, 
    101420, 101430, 101440, 101430, 101440, 101450, 101480, _, 101520, 
    101550, 101560, 101570, 101580, 101600, 101580, 101610, 101570, 101580, 
    101580, 101580, 101580, 101580, 101580, 101540, 101510, 101470, 101430, 
    101380, 101330, 101250, 101230, 101180, 101150, 101110, 101080, 101070, 
    101000, 100960, 100960, 100920, 100900, 100880, 100880, 100910, 100900, 
    100890, 100890, 100880, 100860, 100840, 100810, 100770, 100720, 100680, 
    100630, 100600, 100550, 100490, 100450, 100400, 100360, 100320, 100280, 
    100240, 100210, 100200, 100200, 100190, 100220, 100240, 100260, 100280, 
    100290, 100300, 100330, 100340, 100350, 100360, 100370, 100400, 100430, 
    100460, 100470, 100490, 100530, 100540, 100560, 100560, 100600, 100640, 
    100680, 100710, 100760, 100840, 100890, 100940, 101000, 101020, 101030, 
    101050, 101080, 101110, 101170, 101190, 101220, 101250, 101290, 101300, 
    101330, 101350, 101350, 101360, 101380, 101360, 101370, 101400, 101450, 
    101450, 101510, 101530, 101540, 101540, 101540, 101530, 101570, 101610, 
    101610, 101610, 101610, 101630, 101660, 101690, 101680, 101660, 101630, 
    101630, 101620, 101600, 101600, 101600, 101590, 101580, 101600, 101610, 
    101600, 101590, 101580, 101550, 101520, 101500, 101480, 101470, 101450, 
    101430, 101420, 101390, 101370, 101360, 101340, 101320, 101300, 101270, 
    101250, 101220, 101200, 101190, 101160, 101160, 101130, 101110, 101080, 
    101050, 101010, 101010, 100990, 100980, 100960, 100960, 100980, 101000, 
    101030, 101040, 101060, 101080, 101090, 101120, 101140, 101180, 101210, 
    101250, 101290, 101310, 101340, 101360, 101390, 101400, 101410, 101420, 
    101440, 101450, 101460, 101480, 101510, 101520, 101540, 101520, 101550, 
    101560, 101580, 101600, 101600, 101620, 101630, 101660, 101680, 101700, 
    101710, 101690, 101680, 101680, 101680, 101660, 101640, 101640, 101640, 
    101620, 101610, 101580, 101580, 101560, 101540, 101510, 101480, 101450, 
    101410, 101390, 101330, 101300, 101290, 101270, 101240, 101170, 101150, 
    101100, 101060, 101040, 101020, 100980, 100940, 100930, 100940, 100980, 
    100970, 100970, 101000, 100990, 101020, 101050, 101060, 101110, 101160, 
    101190, 101240, 101290, 101340, 101380, 101400, 101440, 101480, 101500, 
    101590, 101650, 101700, 101750, 101790, 101820, 101860, 101880, 101930, 
    101970, 102000, 102030, 102060, 102090, 102130, 102150, 102200, 102240, 
    102240, 102270, 102290, 102300, 102330, 102370, 102390, 102420, 102480, 
    102510, 102540, 102570, 102600, 102650, 102710, 102760, 102780, 102820, 
    102850, 102890, 102910, 102950, 102980, 102980, 102990, 102990, 102990, 
    102970, 102970, 102970, 102950, 102970, 102960, 102970, 102940, 102920, 
    102920, 102910, 102920, 102900, 102880, 102880, 102870, 102860, 102860, 
    102860, 102850, 102810, 102820, 102830, 102820, 102800, 102800, 102800, 
    102790, 102770, 102760, 102740, 102740, 102730, 102730, 102700, 102690, 
    102700, 102690, 102700, 102680, 102690, 102700, 102710, 102710, 102730, 
    102730, 102730, 102740, 102760, 102790, 102790, 102800, 102820, 102840, 
    102860, 102870, 102900, 102920, 102950, 102970, 103010, 103040, 103050, 
    103090, 103120, 103150, 103180, 103220, 103270, 103270, 103280, 103310, 
    103330, 103350, 103370, 103390, 103380, 103410, 103410, 103410, 103420, 
    103410, 103410, 103400, 103390, 103380, 103330, 103260, 103210, 103140, 
    103110, 103090, 103040, 102990, 102910, 102900, 102840, 102780, 102660, 
    102570, 102510, 102440, 102370, 102260, 102160, 102040, 101930, 101860, 
    101780, 101660, 101550, 101460, 101400, 101370, 101260, 101160, 101150, 
    101100, 101080, 101080, 101170, 101130, 101160, 101190, 101220, 101230, 
    101280, 101350, 101390, 101460, 101490, 101530, 101570, 101640, 101690, 
    101720, 101780, 101840, 101900, 101940, 101980, 102060, 102090, 102090, 
    102140, 102170, 102190, 102230, 102260, 102290, 102310, 102350, 102330, 
    102340, 102380, 102380, 102350, 102340, 102340, 102320, 102320, 102300, 
    102290, 102260, 102260, 102270, 102280, 102240, 102210, 102210, 102210, 
    102200, 102160, 102170, 102150, 102140, 102100, 102100, 102070, 102040, 
    102020, 101990, 101990, 101980, 101990, 102010, 102070, 102130, 102170, 
    102180, 102200, 102230, 102270, 102310, 102330, 102360, 102360, 102410, 
    102440, 102460, 102490, 102490, 102500, 102500, 102510, 102510, 102520, 
    102540, 102540, 102560, 102590, 102620, 102640, 102660, 102680, 102690, 
    102690, 102670, 102660, 102650, 102670, 102680, 102690, 102690, 102700, 
    102680, 102660, 102650, 102630, 102590, 102570, 102530, 102490, 102430, 
    102360, 102290, 102210, 102150, 102030, 101960, 101850, 101750, 101670, 
    101550, 101470, 101410, 101330, 101250, 101210, 101140, 101070, 101030, 
    100960, 100910, 100830, 100730, 100670, 100590, 100520, 100430, 100330, 
    100280, 100170, 100060, 99970, 99880, 99880, 99830, 99850, 99810, 99900, 
    99940, 99970, 100070, 100120, 100250, 100390, 100530, 100620, 100730, 
    100860, 100970, 101050, 101160, 101220, 101300, 101360, 101410, 101440, 
    101470, 101510, 101500, 101520, 101520, 101540, 101570, 101580, 101560, 
    101540, 101540, 101560, 101560, 101560, 101590, 101600, 101680, 101740, 
    101770, 101770, 101790, 101800, 101800, 101800, 101810, 101800, 101810, 
    101830, 101770, 101850, 101870, 101870, 101890, 101890, 101880, 101880, 
    101890, 101900, 101920, 101940, 101960, 101970, 101980, 101970, 101980, 
    101980, 101960, 101940, 101910, 101920, 101900, 101910, 101920, 101930, 
    101930, 101950, 101970, 102000, 102010, 102030, 102050, 102080, 102120, 
    102170, 102210, 102270, 102290, 102310, 102330, 102350, 102360, 102350, 
    102380, 102390, 102380, 102410, 102410, 102430, 102410, 102380, 102320, 
    102280, 102210, 102080, 101970, 101820, 101800, 101660, 101660, 101670, 
    101690, 101750, 101880, 101950, 101980, 102020, 102110, 102150, 102220, 
    102230, 102270, 102300, 102270, 102280, 102230, 102200, 102180, 102150, 
    102080, 102030, 102010, 102020, 101980, 101910, 101870, 101840, 101780, 
    101730, 101660, 101630, 101570, 101540, 101520, 101540, 101550, 101570, 
    101560, 101560, 101570, 101550, 101580, 101560, 101580, 101610, 101640, 
    101670, 101700, 101750, 101790, 101820, 101850, 101900, 101890, 101950, 
    101970, 102000, 102000, 102060, 102110, 102150, 102190, 102210, 102230, 
    102250, 102270, 102310, 102310, 102370, 102420, 102470, 102510, 102540, 
    102620, 102640, 102670, 102720, 102730, 102760, 102780, 102810, 102800, 
    102810, 102850, 102850, 102840, 102850, 102850, 102850, 102810, 102830, 
    102800, 102790, 102770, 102780, 102800, 102820, 102800, 102760, 102740, 
    102700, 102680, 102640, 102610, 102590, 102570, 102570, 102560, 102540, 
    102490, 102450, 102410, 102340, 102270, 102250, 102200, 102090, 102000, 
    101980, 102000, 101950, 101890, 101820, 101800, 101740, 101740, 101710, 
    101660, 101660, 101630, 101590, 101550, 101560, 101510, 101390, 101330, 
    101270, 101180, 101160, 101100, 101150, 101160, 101180, 101290, 101350, 
    101410, 101470, 101490, 101500, 101460, 101470, 101450, 101500, 101540, 
    101620, 101630, 101660, 101730, 101780, 101710, 101730, 101650, 101550, 
    101540, 101460, 101350, 101270, 101170, 101060, 101030, 101000, 100970, 
    100930, 100880, 100860, 100830, 100780, 100760, 100720, 100700, 100790, 
    100780, 100810, 100850, 100880, 100900, 100920, 100950, 100970, 100990, 
    101010, 101040, 101080, 101100, 101120, 101150, 101150, 101220, 101180, 
    101130, 101090, 101110, 101090, 101090, 101020, 101000, 100890, 100810, 
    100700, 100580, 100470, 100340, 100230, 100210, 100240, 100260, 100320, 
    100400, 100500, 100650, 100780, 100900, 100990, 101070, 101110, 101170, 
    101180, 101190, 101250, 101280, 101240, 101210, 101190, 101140, 101050, 
    101070, 101110, 101120, 101190, 101210, 101300, 101340, 101360, 101400, 
    101430, 101420, 101400, 101370, 101320, 101270, 101240, 101210, 101150, 
    101060, 100970, 100920, 100840, 100780, 100720, 100670, 100610, 100570, 
    100530, 100480, 100480, 100500, 100500, 100470, 100450, 100460, 100480, 
    100540, 100600, 100660, 100700, 100750, 100740, 100730, 100700, 100690, 
    100670, 100680, 100640, 100600, 100590, 100570, 100550, 100550, 100560, 
    100520, 100490, 100470, 100440, 100440, 100450, 100470, 100490, 100460, 
    100500, 100570, 100630, 100590, 100570, 100590, 100610, 100770, 100780, 
    100800, 100790, 100760, 100800, 100870, 100900, 100920, 100930, 100960, 
    100960, 100910, 100910, 100870, 100850, 100810, 100790, 100760, 100720, 
    100700, 100670, 100630, 100600, 100550, 100530, 100500, 100470, 100460, 
    100420, 100450, 100430, 100440, 100410, 100410, 100430, 100480, 100480, 
    100500, 100470, 100490, 100510, 100500, 100450, 100400, 100380, 100370, 
    100380, 100340, 100320, 100320, 100320, 100290, 100250, 100230, 100210, 
    100150, 100110, 100060, 100020, 100010, 99990, 99940, 99850, 99800, 
    99740, 99720, 99710, 99700, 99660, 99590, 99540, 99500, 99480, 99480, 
    99490, 99480, 99490, 99490, 99460, 99410, 99440, 99470, 99490, 99460, 
    99440, 99440, 99440, 99450, 99440, 99480, 99440, 99510, 99520, 99580, 
    99600, 99650, 99710, 99730, 99770, 99780, 99810, 99840, 99860, 99900, 
    99960, 99970, 100000, 100040, 100060, 100070, 100050, 100060, 100080, 
    100110, 100140, 100140, 100140, 100140, 100140, 100150, 100140, 100170, 
    100190, 100200, 100210, 100220, 100230, 100230, 100230, 100250, 100270, 
    100280, 100290, 100290, 100300, 100300, 100310, 100320, 100310, 100280, 
    100250, 100230, 100190, 100160, 100130, 100120, 100100, 100100, 100100, 
    100110, 100130, 100140, 100150, 100150, 100150, 100150, 100140, 100140, 
    100150, 100150, 100170, 100200, 100250, 100260, 100310, 100340, 100370, 
    100410, 100450, 100470, 100500, 100550, 100580, 100630, 100680, 100710, 
    100750, 100770, 100800, 100820, 100820, 100840, 100840, 100840, 100810, 
    100800, 100800, 100810, 100810, 100800, 100780, 100810, 100820, 100800, 
    100830, 100860, 100870, 100920, 100950, 100990, 101020, 101060, 101070, 
    101100, 101120, 101150, 101150, 101140, 101140, 101110, 101110, 101110, 
    101060, 101030, 101020, 101000, 100990, 100980, 100930, 100940, 100950, 
    100980, 100980, 101000, 101000, 100990, 101020, 101020, 101040, 101030, 
    101030, 101070, 101070, 101070, 101070, 101090, 101100, 101110, 101120, 
    101130, 101150, 101150, _, 101180, 101170, 101190, 101190, 101190, 
    101200, 101200, 101180, 101180, 101170, 101190, 101230, 101230, 101230, 
    101240, _, 101250, 101250, 101260, 101260, 101260, 101250, 101250, 
    101250, 101260, 101240, 101280, 101280, 101290, _, 101280, 101270, 
    101240, 101180, 101140, 101100, 101030, 100950, 100910, 100840, 100670, 
    100500, 100350, 100270, 100200, 100150, 100080, 100030, 99990, 99930, 
    99940, 99920, 99840, 99810, 99780, 99740, 99720, 99680, 99690, 99660, 
    99650, 99620, 99630, 99660, 99650, 99650, 99660, 99660, 99670, 99690, 
    99650, 99640, 99610, 99650, 99700, 99830, 99980, 100110, 100230, 100360, 
    100470, 100640, 100820, _, _, _, _, _, 101330, 101390, 101420, 101470, 
    101520, 101560, 101570, 101610, 101660, 101670, 101690, 101700, 101690, 
    101690, 101680, 101640, 101570, 101520, 101480, 101430, 101360, 101360, 
    101330, 101300, 101270, 101240, 101220, 101220, 101200, 101180, 101150, 
    101150, 101120, 101130, 101130, 101130, 101120, 101130, _, 101140, 
    101120, 101120, 101090, 101100, 101070, 101090, 101080, 101080, 101060, 
    101040, 101030, 101050, 101030, 101020, 101030, 101030, 101030, 101040, 
    101030, 101070, 101070, 101090, 101090, 101100, 101110, 101130, 101110, 
    101130, 101160, 101210, 101210, 101190, 101190, 101200, 101200, 101270, 
    101290, 101240, 101170, 101160, 101170, 101240, 101310, 101350, 101370, 
    _, 101460, 101550, 101570, 101600, 101610, 101660, 101690, 101700, 
    101750, 101790, 101760, 101740, 101730, 101700, 101690, 101650, 101580, 
    101540, 101460, 101390, 101310, 101230, 101250, 101190, 101140, 101080, 
    101060, 101040, 100990, 100990, 101050, 101110, 101090, 101180, 101170, 
    101150, 101150, 101240, 101220, 101190, 101210, 101220, 101250, 101200, 
    101200, 101190, 101100, 101100, 101010, 100890, 100830, 100730, 100630, 
    100630, 100600, 100550, 100510, 100550, 100590, 100580, 100580, 100600, 
    100650, 100660, 100700, 100720, 100730, 100820, 100850, 100930, 100970, 
    100960, 100960, 100940, 100960, 100980, 100930, 100910, 100870, 100890, 
    100870, 100860, 100810, 100800, 100780, 100770, 100790, 100840, 100890, 
    100940, 100980, 101060, 101140, 101220, 101270, 101290, 101310, 101340, 
    101370, 101390, 101410, 101450, 101460, 101500, 101540, 101550, 101570, 
    101570, 101570, 101570, 101580, 101580, 101590, 101580, 101500, 101540, 
    101580, 101540, 101530, 101510, 101550, 101470, 101450, 101430, 101410, 
    101360, 101360, 101350, 101310, 101280, 101280, 101240, 101170, 101090, 
    101060, 101010, 101000, 100930, 100930, 100910, 100840, 100550, 100450, 
    100510, 100460, 100480, 100470, 100380, 100330, 100300, 100330, 100300, 
    100280, 100310, 100370, 100370, 100400, 100420, 100430, 100470, 100470, 
    100440, 100470, 100520, 100550, 100590, 100630, 100650, 100680, 100700, 
    100730, 100770, 100780, _, 100830, 100860, 100890, 100910, 100980, 
    100980, 100970, 101010, 101040, 101050, 101030, 101040, 101000, 101010, 
    101030, 101050, 101050, 101080, 101080, 101060, 101040, 100980, 101000, 
    101030, 101020, 100990, 100990, 100960, _, 100970, 101000, 101000, 
    101010, 100980, 100950, 100920, 100930, 100940, 100940, 100950, 100940, 
    100870, 100800, 100740, 100670, 100640, 100610, 100570, 100550, 100530, 
    100530, 100530, 100520, 100530, 100570, 100560, 100570, 100530, 100520, 
    100500, 100490, 100470, 100450, 100450, 100400, 100340, 100310, 100230, 
    100170, 100150, 100100, 100030, 99960, 99930, 99900, 99870, 99830, 99800, 
    99780, 99750, 99740, 99740, 99700, 99670, 99650, 99650, 99670, 99660, 
    99650, 99660, 99650, 99630, 99620, 99610, 99610, 99610, 99610, 99590, 
    99590, 99570, 99570, 99550, 99530, 99560, 99600, 99650, 99670, 99700, 
    99730, 99770, 99800, 99790, 99820, _, 99910, 99910, 99930, 99910, 99870, 
    99850, 99920, 99960, 99990, 100030, 100050, 100070, 100050, 100040, 
    100040, 100050, 100050, 100060, 100040, 100050, 100110, 100120, 100130, 
    100180, 100240, 100290, 100370, 100430, 100470, 100520, 100610, 100660, 
    100710, 100780, 100820, 100900, 100980, 101030, 101080, 101110, 101150, 
    101200, 101260, 101290, 101350, 101400, 101450, 101480, 101510, 101540, 
    101550, 101560, 101580, 101590, 101590, 101570, 101550, 101540, 101540, 
    101560, 101550, 101530, 101480, 101480, 101450, 101430, 101420, 101400, 
    101380, 101350, 101350, 101320, 101320, 101300, 101260, 101230, 101180, 
    101180, 101120, 101110, 101110, 101100, 101100, 101130, 101080, 101050, 
    101020, 101000, 100950, 100880, 100750, 100670, 100650, 100570, 100420, 
    100300, _, 100230, 100170, _, 100120, 100050, 99980, 99930, 99970, 99900, 
    99900, 99960, 99940, 99860, 99820, 99790, 99760, 99730, 99690, 99700, 
    99660, 99660, 99700, 99670, 99640, 99630, 99640, 99620, 99600, 99590, 
    99560, 99550, 99550, 99550, 99570, 99550, 99560, 99580, 99580, 99580, 
    99600, 99600, 99650, 99680, 99710, 99760, 99790, 99840, 99870, 99920, 
    99960, 100000, 100050, 100080, 100140, 100160, 100210, 100250, 100290, 
    100320, 100340, 100360, 100370, 100380, 100380, 100380, 100400, 100430, 
    100450, 100460, 100510, 100550, 100620, 100680, 100740, 100790, 100820, 
    100880, 100950, 101000, 101060, 101070, 101120, 101170, 101210, 101220, 
    101240, 101260, 101310, 101350, 101370, 101420, 101450, _, 101530, 
    101580, 101600, 101630, 101670, 101680, 101720, 101760, 101740, 101790, 
    101850, 101890, 101900, 101940, 102000, 102010, 102010, 102040, 102050, 
    102050, _, _, 102150, 102170, 102180, 102210, 102190, 102200, 102160, 
    102170, 102170, 102130, 102100, 102070, 102020, 102000, 102080, 102040, 
    101800, 101760, 101800, 101730, 101700, 101440, 101420, 101270, 101070, 
    100900, 100870, 100800, 100800, 100720, 100550, 100500, 100410, 100440, 
    100400, 100400, 100350, 100470, 100470, 100480, 100440, 100330, 100220, 
    100100, 100000, 99930, 99880, 99910, 99980, 100130, 100260, 100380, 
    100490, 100580, 100600, 100650, 100680, 100700, 100810, 100880, 100920, 
    100960, _, 101060, 101090, 101100, 101120, 101120, 101140, 101170, 
    101160, _, 101190, 101210, 101240, 101230, 101220, 101210, 101200, 
    101190, 101200, 101200, 101220, 101210, 101210, 101210, 101230, 101230, 
    101240, 101230, 101270, 101270, 101300, 101320, 101350, 101360, 101420, 
    101480, 101520, 101560, 101590, 101620, 101620, 101650, 101670, 101670, 
    101670, 101680, 101690, 101680, 101680, 101720, 101710, 101720, 101720, 
    101730, 101720, 101740, 101750, 101750, 101790, 101800, 101790, 101810, 
    101820, 101800, 101800, 101780, 101770, 101740, 101750, 101750, 101760, 
    101730, 101710, 101710, 101690, 101680, 101670, 101630, 101590, 101570, 
    101570, 101550, 101540, 101540, 101510, 101510, 101510, 101480, 101460, 
    101440, 101420, 101430, 101430, 101430, 101420, 101420, 101400, 101400, 
    101400, 101390, 101370, 101360, 101350, 101350, 101360, 101360, 101350, 
    101340, 101360, 101370, 101370, 101340, 101340, 101320, 101310, 101260, 
    101230, 101210, 101200, 101200, 101170, 101160, 101160, 101140, 101140, 
    101120, 101110, 101110, 101120, 101100, 101100, 101130, 101130, 101120, 
    101140, 101130, 101140, 101140, 101140, 101140, 101160, 101170, 101200, 
    101190, 101180, 101190, 101220, 101220, 101240, 101260, 101260, 101270, 
    101310, 101330, 101360, 101370, 101390, 101400, 101420, 101440, 101440, 
    101470, 101460, 101460, 101470, 101450, 101470, 101450, 101450, 101450, 
    101450, 101420, 101400, 101360, 101370, 101380, 101360, 101400, 101430, 
    101470, 101500, 101530, 101560, 101540, 101560, 101590, 101600, 101610, 
    101620, 101610, 101630, 101630, 101630, 101620, 101600, 101610, 101610, 
    101590, 101560, 101600, 101590, 101580, 101600, 101610, 101620, 101620, 
    101610, 101640, 101640, 101660, 101650, 101690, 101720, 101730, 101760, 
    101750, 101740, 101740, 101740, 101750, 101730, 101740, 101720, 101690, 
    101650, 101580, 101560, 101540, 101510, 101470, 101470, 101440, 101400, 
    101430, 101400, 101380, 101380, 101380, 101370, 101350, 101380, 101380, 
    101340, 101360, 101310, 101250, 101200, 101130, 101140, 101150, 101110, 
    101120, 101010, 100970, 100960, 100790, 100710, 100600, 100570, 100360, 
    100350, 100400, 100370, 100350, 100460, 100470, 100460, 100430, 100450, 
    100450, 100460, 100520, 100540, 100600, 100650, 100690, 100760, 100830, 
    100860, 100910, 100970, 100990, 101050, 101100, 101150, 101190, 101240, 
    101290, 101330, 101350, 101370, 101400, 101470, 101500, 101520, 101560, 
    101610, 101650, 101670, 101690, 101740, 101740, 101760, 101770, 101770, 
    101760, 101750, 101770, 101770, 101750, 101760, 101750, 101770, 101750, 
    101760, 101760, 101720, 101740, 101740, 101750, 101750, 101740, 101800, 
    101800, 101780, 101750, 101760, 101750, 101750, 101770, 101760, 101750, 
    101750, 101750, 101740, 101750, 101760, 101750, 101740, 101720, 101670, 
    101690, 101670, 101650, 101630, 101630, 101640, 101630, 101620, 101650, 
    101630, 101640, 101650, 101620, 101650, 101700, 101680, 101700, 101710, 
    101740, 101790, 101870, 101870, 101870, 101870, 101880, 101890, 101890, 
    101890, 101910, 101920, 101910, 101890, 101880, 101840, 101840, 101810, 
    101790, 101740, 101730, 101700, 101680, 101650, 101610, 101580, 101550, 
    101520, 101480, 101460, 101420, 101390, 101380, 101340, 101280, 101250, 
    101200, 101160, 101120, 101060, 100970, 100910, 100840, 100780, 100690, 
    100600, 100550, 100550, 100540, 100520, 100520, 100530, 100540, 100540, 
    100560, 100590, 100720, 100740, 100820, 100860, 100900, 100980, 101020, 
    101050, 101090, 101080, 101090, 101040, 101030, 101050, 101030, 100990, 
    100990, 100970, 100940, 100920, 100900, 100880, 100830, 100780, 100770, 
    100750, 100730, 100720, 100710, 100680, 100670, 100670, 100650, 100630, 
    100610, 100590, 100550, 100510, 100480, 100470, 100460, 100420, 100350, 
    100290, 100220, 100110, 100040, 100020, 99960, 99900, 99850, 99810, 
    99790, 99800, 99840, 99850, 99910, 99930, 99940, 99990, 100010, 100060, 
    100080, 100090, 100130, 100110, 100090, 100090, 100070, 100050, 100020, 
    100010, 100000, 100000, 99980, 99990, 100030, 100030, 100030, 99990, 
    99970, 99920, 99840, 99800, 99770, 99730, 99660, 99610, 99560, 99530, 
    99520, 99500, 99470, 99450, 99420, 99420, 99440, 99460, 99530, 99540, 
    99560, 99610, 99610, 99580, 99580, 99610, 99600, 99560, 99570, 99530, 
    99520, 99530, 99520, 99490, 99530, 99550, 99570, 99610, 99660, 99690, 
    99740, 99810, 99840, 99870, 99900, 99950, 99960, 99970, 99980, 99990, 
    99970, 99960, 99970, 99970, 99940, 99920, 99910, 99940, 99950, 99980, 
    100020, 100100, 100170, 100250, 100300, 100380, 100430, 100520, 100590, 
    100640, 100700, 100720, 100720, 100710, 100670, 100570, 100480, 100420, 
    100320, 100210, 100130, 100020, 99990, 99920, 99940, 99950, 99960, 99980, 
    100050, 100080, 100190, 100250, 100330, 100390, 100430, 100450, 100490, 
    100520, 100520, 100540, 100530, 100550, 100530, 100550, 100520, 100490, 
    100460, 100470, 100460, 100430, 100450, 100450, 100460, 100460, 100510, 
    100520, 100530, 100550, 100560, 100570, 100600, 100620, 100650, 100650, 
    100650, 100650, 100660, 100680, 100680, 100670, 100680, 100720, 100700, 
    100710, 100730, 100740, 100760, 100780, 100810, 100850, 100850, 100890, 
    100910, 100970, 101000, 101030, 101060, 101050, 101110, 101120, 101120, 
    101160, 101200, 101210, 101250, 101290, 101310, 101320, 101350, 101350, 
    101350, 101400, 101430, 101440, 101450, 101450, 101460, 101440, 101440, 
    101390, 101370, 101310, 101270, 101190, 101130, 101100, 101060, 101020, 
    101000, 100960, 100950, 100950, 100930, 100910, 100910, 100920, 100940, 
    100960, 100950, 100960, 100960, 100920, 100880, 100830, 100810, 100830, 
    100750, 100750, 100730, 100740, 100700, 100710, 100710, 100700, 100640, 
    100570, 100560, 100490, 100390, 100290, 100260, 100240, 100210, 100240, 
    100230, 100210, 100180, 100140, 100070, 100020, 99920, 99770, 99740, 
    99770, 99840, 99960, 100050, 100090, 100140, 100210, 100280, 100330, 
    100410, 100420, 100440, 100500, 100520, 100580, 100600, 100630, 100690, 
    100670, 100660, 100650, 100660, 100640, 100590, 100560, 100570, 100600, 
    100610, 100590, 100570, 100640, 100630, 100640, 100640, 100650, 100660, 
    100650, 100680, 100720, 100740, 100750, 100780, 100780, 100790, 100790, 
    100790, 100780, 100800, 100780, 100770, 100770, 100790, 100790, 100830, 
    100830, 100850, 100850, 100830, 100840, 100850, 100850, 100860, 100870, 
    100890, 100880, 100840, 100820, 100800, 100740, 100730, 100690, 100690, 
    100720, 100710, 100720, 100730, 100770, 100800, 100850, 100920, 100950, 
    101010, 101080, 101150, 101210, 101280, 101340, 101390, 101440, 101470, 
    101520, 101560, 101610, 101690, 101720, 101760, 101810, 101830, 101830, 
    101880, 101940, 101960, 101990, 102020, 102020, 102010, 102020, 102030, 
    102050, 102060, 102060, 102030, 102000, 101960, 101900, 101860, 101810, 
    101790, 101750, 101720, 101680, 101630, 101590, 101540, 101430, 101370, 
    101310, 101230, 101180, 101140, 101070, 101000, 100950, 100930, 100880, 
    100860, 100810, 100730, 100710, 100620, 100580, 100510, 100510, 100410, 
    100420, 100400, 100370, 100330, 100300, 100280, 100250, 100240, 100260, 
    100250, 100240, 100270, 100270, 100280, 100270, 100260, 100290, 100290, 
    100350, 100350, 100330, 100350, 100350, 100350, 100350, 100330, 100320, 
    100270, 100210, 100170, 100150, 100130, 100090, 100120, 100150, 100140, 
    100130, 100080, 100080, 100110, 100120, 100130, 100110, 100100, 100070, 
    100070, 100010, 99950, 99910, 99860, 99800, 99720, 99660, 99600, 99490, 
    99490, 99480, 99480, 99420, 99280, 99200, 99210, 99150, 99120, 99070, 
    99050, 99030, 99000, 98890, 98920, 98930, 98960, 98980, 98980, 99060, 
    99100, 99180, 99210, 99300, 99320, 99350, 99440, 99510, 99560, 99600, 
    99690, 99810, 99930, 100050, 100100, 100170, 100260, 100310, 100360, 
    100430, 100470, 100490, 100530, 100570, 100600, 100610, 100680, 100730, 
    100760, 100750, 100750, 100810, 100840, 100890, 100910, 100920, 100970, 
    101010, 101030, 101010, 101030, 101050, 101100, 101180, 101210, 101190, 
    101200, 101210, 101240, 101260, 101240, 101240, 101230, 101230, 101250, 
    101300, 101330, 101350, 101350, 101390, 101400, 101400, 101390, 101400, 
    101410, 101390, 101380, 101370, 101390, 101400, 101400, 101400, 101410, 
    101410, 101420, 101390, 101380, 101390, 101400, 101390, 101410, 101420, 
    101440, 101440, 101460, 101490, 101520, 101520, 101530, 101530, 101530, 
    101530, 101520, 101500, 101520, 101520, 101540, 101540, 101530, 101510, 
    101490, 101480, 101500, 101500, 101520, 101530, 101540, 101550, 101560, 
    101560, 101550, 101540, 101540, 101530, 101520, 101460, 101460, 101440, 
    101410, 101390, 101360, 101330, 101310, 101290, 101260, 101250, 101250, 
    101210, 101210, 101180, 101160, 101130, 101130, 101140, 101120, 101110, 
    101060, 101030, 101000, 100970, 100940, 100960, 100930, 100900, 100850, 
    100860, 100790, 100750, 100680, 100680, 100610, 100610, 100560, 100530, 
    100460, 100400, 100340, 100270, 100180, 100170, 100140, 100130, 100080, 
    100080, 100060, 100030, 100010, 99980, 99930, 99880, 99870, 99870, 99840, 
    99820, 99810, 99830, 99850, 99860, 99870, 99860, 99880, 99870, 99900, 
    99910, 99900, 99920, 99940, 99960, 99960, 99970, 99990, 99980, 99960, 
    99910, 99830, 99780, 99750, 99700, 99670, 99610, 99640, 99620, 99630, 
    99680, 99760, 99820, 99910, 100000, 100080, 100180, 100250, 100330, 
    100370, 100380, 100420, 100400, 100390, 100370, 100360, 100300, 100290, 
    100270, 100260, 100230, 100190, 100190, 100210, 100240, 100250, 100330, 
    100350, 100400, 100500, 100550, 100610, 100660, 100680, 100730, 100770, 
    100780, 100800, 100790, 100790, 100740, 100710, 100670, 100680, 100670, 
    100640, 100660, 100670, 100720, 100740, 100820, 100900, 100930, 100990, 
    101070, 101160, 101200, 101270, 101330, 101350, 101360, 101400, 101440, 
    101420, 101410, 101560, 101640, 101670, 101700, 101700, 101710, 101780, 
    101810, 101820, 101830, 101850, 101820, 101790, 101730, 101700, 101680, 
    101610, 101570, 101530, 101460, 101400, 101300, 101240, 101130, 101030, 
    101000, 100930, 100900, 100780, 100740, 100680, 100580, 100540, 100290, 
    100230, 100220, 100220, 100220, 100220, 100200, 100220, 100210, 100220, 
    100250, 100220, 100290, 100290, 100340, 100440, 100440, 100510, 100570, 
    100650, 100680, 100770, 100870, 100920, 100980, 101040, 101130, 101130, 
    101130, 101190, 101250, 101300, 101330, 101350, 101420, 101450, 101460, 
    101480, 101500, 101510, 101550, 101540, 101570, 101600, 101620, 101630, 
    101650, 101680, 101620, 101610, 101630, 101560, 101520, 101450, 101410, 
    101360, 101250, 101190, 101160, 101060, 101020, 100930, 100860, 100800, 
    100700, 100710, 100670, 100680, 100660, 100690, 100690, 100690, 100730, 
    100750, 100740, 100780, 100780, 100820, 100830, 100850, 100840, 100830, 
    100810, 100770, 100740, 100700, 100700, 100680, 100690, 100700, 100720, 
    100750, 100760, 100810, 100820, 100890, 100910, 100940, 100940, 100940, 
    100950, 100970, 101010, 101010, 101020, 101050, 101090, 101150, 101190, 
    101230, 101280, 101320, 101370, 101430, 101510, 101560, 101610, 101640, 
    101700, 101750, 101780, 101810, 101880, 101910, 101930, 101930, 101970, 
    101980, 102010, 102020, 102030, 102020, 102010, 101990, 101980, 101940, 
    101920, 101880, 101820, 101770, 101750, 101720, 101660, 101640, 101620, 
    101550, 101520, 101490, 101460, 101460, 101450, 101480, 101510, 101520, 
    101530, 101530, 101560, 101560, 101570, 101560, 101540, 101550, 101550, 
    101600, 101620, 101620, 101650, 101620, 101590, 101560, 101560, 101590, 
    101590, 101620, 101630, 101670, 101690, 101710, 101760, 101760, 101800, 
    101840, 101890, 101920, 101960, 102010, 102040, 102070, 102120, 102140, 
    102180, 102210, 102230, 102260, 102300, 102310, 102340, 102360, 102400, 
    102430, 102440, 102460, 102450, 102470, 102500, 102520, 102520, 102540, 
    102560, 102550, 102570, 102580, 102600, 102610, 102640, 102650, 102680, 
    102710, 102710, 102740, 102780, 102790, 102780, 102790, 102720, 102690, 
    102760, 102740, 102780, 102770, 102820, 102850, 102870, 102880, 102900, 
    102910, 102930, 102970, _, 103010, 103040, 103040, 103070, 103070, 
    103070, 103090, 103090, 103120, 103130, 103140, 103160, 103160, 103170, 
    103180, 103180, 103190, 103180, 103190, 103190, 103200, 103190, 103220, 
    103230, 103250, 103260, 103270, 103280, 103310, 103320, 103320, 103340, 
    103350, 103380, 103390, 103400, _, 103400, 103430, 103430, 103440, 
    103440, 103460, 103450, 103470, 103480, 103490, 103510, 103510, 103520, 
    103500, 103490, _, 103500, 103500, 103490, 103480, 103470, 103470, 
    103500, 103480, 103480, 103470, 103470, 103470, 103430, 103430, 103450, 
    _, 103480, _, 103470, 103470, 103440, 103420, 103420, 103410, 103390, 
    103400, 103380, 103370, 103350, _, 103360, 103350, 103330, 103330, 
    103330, 103330, 103330, 103320, 103300, 103310, 103320, 103340, 103350, 
    103370, 103370, 103340, 103320, 103320, 103310, 103320, 103320, 103300, 
    103300, 103280, 103270, 103260, 103240, 103230, 103230, 103260, 103250, 
    103250, 103230, 103230, 103240, 103260, 103280, 103280, 103290, 103280, 
    103270, 103260, 103280, 103280, 103290, 103270, 103280, 103280, 103290, 
    103280, 103270, 103260, 103260, 103270, 103250, 103260, 103250, 103260, 
    103280, 103270, 103280, 103310, 103310, 103300, 103290, 103270, 103240, 
    103230, 103240, 103230, 103220, 103230, 103240, 103230, 103210, 103210, 
    103210, 103190, 103160, 103150, 103140, 103130, 103120, 103110, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    102780, 102740, 102720, 102690, 102670, 102640, 102630, 102610, 102560, 
    102540, 102550, 102510, 102510, 102490, 102470, 102430, 102400, 102380, 
    102350, 102340, 102350, 102340, 102320, 102310, 102270, 102220, 102140, 
    102070, 102020, 101950, 101890, 101780, 101670, 101610, 101480, 101380, 
    101320, 101200, 101090, 100990, 100870, 100740, 100590, 100500, 100400, 
    100280, 100170, 100060, 99920, 99780, 99700, 99610, 99540, 99490, 99430, 
    99380, 99310, 99230, 99170, 99120, _, 99090, 99190, 99290, 99400, 99470, 
    99570, 99660, 99720, 99740, 99750, 99700, 99640, 99570, 99480, 99420, 
    99340, 99230, 99070, 98900, 98650, 98350, 98080, 98040, 97970, 98010, 
    98010, 98200, 98330, 98480, 98620, 98740, 98830, 98850, 98850, 98800, 
    98790, 98800, 98870, 98940, 98980, 99040, 99080, 99130, 99160, 99140, 
    99140, 99160, 99240, 99290, 99340, 99350, 99400, 99440, 99480, 99520, 
    99570, 99600, 99640, 99650, 99730, 99750, 99790, 99860, 99880, 99920, 
    99950, 99980, 100020, 100050, 100070, 100100, _, 100140, 100230, 100300, 
    100390, 100410, 100500, 100580, 100650, 100720, 100780, 100840, 100890, 
    100920, 100950, 100960, 101000, 101030, 101060, 101090, 101110, 101150, 
    101200, 101240, 101250, 101310, _, 101340, 101360, 101380, 101410, 
    101430, 101470, 101490, 101530, 101530, 101560, 101570, 101590, 101610, 
    101630, 101630, 101660, 101660, 101680, 101710, 101730, 101770, 101780, 
    101790, 101810, 101840, 101850, 101870, 101860, 101880, 101910, 101940, 
    101960, 101990, 102000, 102000, 102000, 102000, 102000, 102000, 102010, 
    102010, 102000, 101990, 102000, 101990, 101960, 101950, 101930, 101910, 
    101910, 101880, 101870, 101870, 101890, 101890, 101890, 101870, 101840, 
    101830, 101800, 101780, 101740, 101710, 101690, 101670, 101640, 101600, 
    101580, 101550, 101530, 101500, 101480, 101450, 101430, 101400, 101380, 
    101380, 101360, 101330, 101310, 101270, 101230, 101180, 101160, 101120, 
    101090, 101070, 101030, 101000, 100960, 100910, 100860, 100800, _, 
    100670, 100540, 100430, 100300, 100210, 100190, 100140, 100140, 100110, 
    100100, 100070, 100040, 100010, 99980, 99930, 99900, 99820, 99820, 99790, 
    99740, 99710, 99660, 99580, 99530, 99520, 99510, 99470, 99480, 99500, 
    99560, 99600, 99630, 99640, 99690, 99800, 99830, 99820, 99880, 99920, 
    99970, 99990, 100020, 100050, 100100, 100120, 100180, 100220, 100220, 
    100230, 100310, 100340, 100340, 100340, 100350, 100360, 100360, 100380, 
    100430, 100480, 100530, 100610, 100720, 100820, 100930, 101020, 101130, 
    101270, 101430, 101570, 101700, 101830, 101900, 101970, 102030, 102080, 
    102130, 102150, 102170, 102190, 102200, 102200, 102210, 102220, 102200, 
    102200, 102170, 102150, 102120, 102090, 102080, 102050, 102030, 102010, 
    _, 101970, 101940, _, 101890, 101860, 101830, 101810, 101780, 101770, 
    101800, 101790, 101760, 101720, 101740, 101720, 101690, 101690, 101670, 
    101660, 101640, 101640, 101670, 101690, 101710, 101730, 101750, 101740, 
    101760, 101770, 101790, 101780, 101790, 101820, 101850, 101890, 101890, 
    101910, 101930, 101920, 101940, 101920, 101920, 101920, 101910, 101910, 
    101890, 101880, 101850, 101810, 101780, 101740, 101710, 101670, 101630, 
    101590, 101490, 101470, 101430, 101380, 101320, 101270, 101210, 101140, 
    101070, 101000, 100930, 100890, 100840, 100790, 100760, 100720, 100690, 
    100650, 100660, _, 100680, 100680, 100690, 100690, 100700, 100730, 
    100760, 100790, 100830, 100870, 100890, 100900, 100900, 100920, 100930, 
    100950, 100970, 101000, 101050, 101070, 101090, 101110, 101150, 101150, 
    101160, 101190, 101210, 101260, 101310, 101320, 101360, 101430, 101490, 
    101530, 101560, 101600, 101620, 101660, 101670, 101680, 101690, 101710, 
    101730, 101750, 101760, 101750, 101740, 101720, 101720, 101710, 101710, 
    101720, 101720, 101740, 101780, 101790, 101810, _, 101810, 101790, 
    101790, 101810, 101810, 101810, 101820, 101830, 101830, 101830, 101830, 
    101820, 101810, _, 101790, 101760, 101730, 101700, 101680, 101660, 
    101660, 101640, 101620, 101580, 101530, 101500, 101470, 101430, 101390, 
    101370, 101330, 101280, 101240, 101220, 101180, 101120, 101060, 101010, 
    100950, 100910, 100860, 100780, 100710, 100630, 100540, 100430, 100300, 
    100200, 100100, 100120, 100130, 100170, 100150, 100140, 100150, 100150, 
    100110, 100120, 100100, 100080, 100040, 100010, 99990, _, 100000, 99970, 
    99950, 99900, 99840, 99800, 99730, _, 99610, 99620, 99610, 99610, 99650, 
    99710, 99750, 99790, 99830, 99910, 99950, 99980, 100000, 100010, 100040, 
    100050, 100050, 100060, 100090, 100090, 100120, 100130, 100150, 100150, 
    100120, 100110, 100070, 100050, _, 100020, 100000, 99970, 99970, 99930, 
    99900, 99850, 99800, 99770, 99730, 99760, 99760, 99710, 99680, 99680, 
    99680, 99700, 99720, 99740, 99740, 99730, 99710, 99720, 99700, 99660, 
    99680, 99670, 99700, 99690, 99690, 99670, 99660, 99640, 99620, 99600, 
    99570, 99560, 99540, 99550, 99580, 99590, 99600, 99610, 99570, 99560, _, 
    _, _, 99630, 99620, 99620, 99600, 99600, 99600, 99610, 99640, 99660, 
    99650, 99650, 99680, 99690, 99700, 99740, 99760, 99790, 99820, 99820, 
    99820, 99830, 99870, 99930, 99960, 99990, 100010, 100040, 100100, 100150, 
    100190, 100210, 100250, 100260, 100270, 100280, 100290, 100310, 100310, 
    100330, 100380, 100420, 100470, 100500, 100510, 100530, 100540, 100550, 
    100540, 100550, 100570, 100570, 100590, 100600, 100600, 100610, 100600, 
    100580, 100600, 100580, 100600, 100580, 100610, 100610, 100630, 100630, 
    100630, 100650, 100660, 100680, 100650, 100650, 100660, 100660, 100680, 
    100690, 100710, 100730, 100740, 100740, 100760, 100770, 100770, 100770, 
    100780, 100780, 100810, 100820, 100850, 100870, 100870, 100890, 100870, 
    100860, 100870, 100870, 100880, 100900, 100880, 100880, 100890, 100900, 
    100890, 100890, 100890, 100870, 100850, 100850, 100820, 100810, 100790, 
    100780, 100790, 100780, 100770, 100760, 100750, 100710, 100710, 100700, 
    100670, 100660, 100660, 100650, 100650, 100650, 100680, 100710, 100730, 
    100740, 100760, 100750, 100750, 100790, 100760, 100800, 100820, 100850, 
    100870, 100890, 100910, 100940, 100950, 100930, 100950, 100970, 100970, 
    101020, 101050, _, 101110, 101120, 101140, 101160, 101180, 101190, 
    101190, 101200, 101190, 101210, 101240, 101270, 101290, 101310, 101310, 
    101330, 101310, 101300, 101270, 101250, 101250, 101230, 101240, 101200, 
    101200, 101170, 101140, 101120, 101130, 101100, 101060, _, 100960, 
    100940, 100930, 100920, 100870, 100790, 100770, 100720, 100640, 100540, 
    100340, 100330, 100180, 100110, 100080, 100010, 99860, _, 99560, 99390, 
    99290, 99210, 99060, 98940, 98820, 98670, 98630, 98630, 98670, 98640, 
    98620, 98600, 98580, 98520, 98500, 98470, 98460, 98440, 98440, _, 98460, 
    98490, 98530, 98620, 98670, 98710, 98840, 98960, 99080, 99230, 99370, 
    99440, 99470, 99630, 99640, 99700, 99790, 99860, 99940, 99960, 99960, 
    99950, 99710, 99710, 99690, 99570, 99440, 99500, 99380, 99360, 99340, 
    99200, 99000, 98900, 98830, 98860, 98760, 98780, 98700, 98570, 98470, 
    98380, 98270, 98170, 98070, 98010, 97930, 97900, 97840, _, 97830, 97790, 
    97720, 97670, 97600, 97550, 97550, 97600, 97660, 97770, 97850, 97890, 
    97920, 97950, 97990, 98020, 98050, 98050, 98090, 98090, 98090, _, 98080, 
    98050, 98040, 98050, 98050, 98050, 98080, 98100, 98120, 98120, 98120, 
    98130, 98100, 98090, 98070, 98060, 98040, 98010, 97990, 97960, 97940, 
    97960, 97970, 97980, 98010, 98050, 98080, 98060, 98130, 98200, 98230, 
    98300, 98320, 98430, 98520, 98610, 98690, 98820, 98890, 98990, 99100, 
    99230, 99300, 99400, 99520, 99620, 99740, 99820, 99900, 99940, 100000, 
    100050, 100090, 100100, 100150, 100180, 100200, 100210, 100210, 100180, 
    100230, 100210, 100180, 100150, 100100, 100060, 100000, 99930, 99980, 
    99920, 99870, 99860, 99850, 99790, 99770, 99730, 99700, 99670, 99620, 
    99620, 99650, 99680, 99690, 99690, 99690, 99670, 99650, 99610, 99590, 
    99560, 99530, 99500, 99460, 99450, 99410, 99370, 99310, 99260, 99190, 
    99110, 98950, 98930, 98830, 98750, 98700, 98660, 98670, 98660, 98680, 
    98720, 98760, 98780, 98810, 98820, 98820, 98780, 98830, 98850, 98950, 
    98990, 99000, 99050, 99050, 99060, 99040, 99030, 99010, 99000, 98990, 
    99000, 99020, 99060, 99060, 99060, 99040, 98960, 98920, 98870, 98800, 
    98750, 98710, 98680, 98640, 98630, 98640, 98670, 98650, 98600, 98630, 
    98730, 98790, 98890, 99000, 99100, 99180, 99230, 99330, 99380, 99450, 
    99480, 99570, 99620, 99720, 99750, 99790, 99840, 99900, 99950, 99970, 
    99990, 100050, 100100, 100120, 100160, 100180, 100230, 100230, 100260, 
    100350, 100360, 100390, 100460, 100500, 100550, 100530, 100560, 100540, 
    100520, 100480, 100430, 100360, 100290, 100260, 100130, 100040, 99930, 
    99790, 99660, 99520, 99380, 99230, 99040, 98830, 98630, 98370, 98090, 
    97820, 97500, 97320, 97140, 96930, 96790, 96690, 96610, 96600, 96630, 
    96660, 96660, 96660, 96650, 96660, 96660, 96690, 96700, 96720, 96760, 
    96870, 96940, 97000, 97040, 97070, 97100, 97100, 97110, 97100, 97070, 
    97020, 97000, 96960, 96840, 96850, 96800, 96770, 96740, 96750, 96750, 
    96750, 96810, 96740, 96690, 96700, 96740, 96860, 97030, 97190, 97340, 
    97500, 97590, 97710, 97820, 97880, 97970, 98050, 98100, 98170, 98190, 
    98200, 98230, 98280, 98300, 98360, 98410, 98490, 98540, 98600, 98640, 
    98700, 98690, 98720, 98710, 98730, 98730, 98730, 98760, 98760, 98760, 
    98770, 98780, 98790, 98770, 98760, 98750, 98730, 98710, 98710, 98720, 
    98730, 98760, 98800, 98820, 98860, 98900, 98900, 98920, 98950, 98970, 
    99010, 99080, 99130, 99180, 99240, 99320, 99350, 99370, 99390, 99410, 
    99440, 99470, 99480, 99480, 99470, 99480, 99490, 99480, 99480, 99470, 
    99480, 99490, 99530, 99550, 99570, 99600, 99610, 99620, 99670, 99720, 
    99750, 99770, 99800, 99840, 99870, 99910, 99940, 99960, 99990, 100030, 
    100090, 100130, 100140, 100170, 100200, 100230, 100240, 100270, 100270, 
    100280, 100280, 100260, 100190, 100200, 100190, 100140, 100080, 100060, 
    100020, 99980, 99950, 99910, 99860, 99840, 99860, 99880, 99860, 99860, 
    99830, 99800, 99730, 99740, 99710, 99640, 99560, 99490, 99440, 99380, 
    99360, 99330, 99290, 99240, 99220, 99180, 99070, 98980, 98860, 98740, 
    98650, 98620, 98580, 98630, 98660, 98700, 98760, 98790, 98790, 98730, 
    98800, 98870, 98970, 99040, 99090, 99170, 99210, 99200, 99220, 99280, 
    99350, 99390, 99440, 99470, 99500, 99540, 99590, 99620, 99640, 99650, 
    99700, 99750, 99810, 99840, 99860, 99870, 99920, 99950, 99970, 100030, 
    100040, 100020, 100030, 100070, 100080, 100120, 100120, 100140, 100150, 
    100150, 100160, 100200, 100230, 100230, 100220, 100240, 100260, 100290, 
    100280, 100290, 100290, 100270, 100290, 100290, 100310, 100290, 100250, 
    100230, 100220, 100190, 100190, 100150, 100150, 100150, 100140, 100120, 
    100110, 100080, 100060, 100040, 100000, 99980, 99970, 99980, 99990, 
    99980, 99990, 99980, 99950, 99920, 99880, 99850, 99840, 99800, 99800, 
    99760, 99770, 99770, 99760, 99780, 99770, 99780, 99790, 99790, 99800, 
    99810, 99830, 99870, 99910, 99930, 99950, 99980, 99990, 100000, 100020, 
    100060, 100070, 100090, 100110, 100140, 100210, 100190, 100200, 100180, 
    100170, 100150, 100120, 100110, 100090, 100090, 100080, 100030, 100020, 
    99990, 99930, 99880, 99830, 99780, 99720, 99660, 99590, 99480, 99400, 
    99360, 99310, 99240, 99170, 99090, 99000, 98930, 98890, 98830, 98780, 
    98750, 98700, 98650, 98600, 98590, 98570, 98540, 98530, 98520, 98500, 
    98480, 98460, 98410, 98430, 98450, 98460, 98480, 98500, 98490, 98510, 
    98510, 98550, 98580, 98600, 98610, 98620, 98620, 98600, 98650, 98670, 
    98680, 98690, 98710, 98770, 98840, 98900, 98930, 98980, 99020, 99060, 
    99070, 99100, 99130, 99130, 99120, 99110, 99130, 99140, 99160, 99130, 
    99130, 99200, 99210, 99210, 99240, 99240, 99240, 99260, 99260, 99270, 
    99270, 99280, 99280, 99270, 99310, 99290, 99260, 99260, 99280, 99260, 
    99270, 99270, 99250, 99220, 99220, 99180, 99150, 99090, 99050, 99010, 
    98980, 98930, 98910, 98880, 98860, 98840, 98810, 98790, 98780, 98770, 
    98790, 98790, 98800, 98790, 98840, 98850, 98870, 98890, 98910, 98950, 
    98980, 99020, 99060, 99070, 99090, 99120, 99160, 99180, 99200, 99240, 
    99250, 99280, 99340, 99350, 99370, 99400, 99430, 99450, 99460, 99470, 
    99510, 99530, 99560, 99550, 99580, 99600, 99630, 99620, 99630, 99650, 
    99700, 99690, 99680, 99690, 99720, 99730, 99780, 99830, 99760, 99840, 
    99870, 99920, 99950, 99980, 100070, 100080, 100100, 100130, 100180, 
    100220, 100240, 100260, 100300, 100340, 100320, 100300, 100310, 100330, 
    100380, 100390, 100400, 100440, 100460, 100420, 100390, 100370, 100400, 
    100370, 100370, 100370, 100370, 100350, 100350, 100360, 100350, 100320, 
    100330, 100320, 100310, 100300, 100290, 100320, 100320, 100330, 100310, 
    100330, 100310, 100310, 100300, 100290, 100310, 100280, 100280, 100280, 
    100310, 100330, 100310, 100350, 100320, 100310, 100320, 100310, 100380, 
    100360, 100370, 100390, 100360, 100360, 100300, 100330, 100390, 100390, 
    100420, 100450, 100470, 100510, 100530, 100530, 100560, 100600, 100640, 
    100680, 100700, 100750, 100810, 100850, 100860, 100890, 100910, 100960, 
    101000, 101050, 101050, 101090, 101110, 101160, 101170, 101160, 101200, 
    101200, 101230, 101190, 101160, 101180, 101200, 101170, 101190, 101160, 
    101180, 101190, 101200, 101220, 101180, 101190, 101240, 101250, 101260, 
    101270, 101300, 101300, 101290, 101320, 101340, 101300, 101290, 101270, 
    101220, 101200, 101220, 101160, 101110, 101060, 100980, 100910, 100820, 
    100730, 100650, 100530, 100400, 100310, 100210, 100020, 99910, 99780, 
    99700, 99580, 99550, 99400, 99340, 99290, 99300, 99270, 99240, 99230, 
    99210, 99180, 99170, 99110, 99150, 99200, 99230, 99350, 99410, 99560, 
    99590, 99590, 99650, 99700, 99720, 99770, 99800, 99900, 100000, 100090, 
    100180, 100250, 100310, 100340, 100400, 100460, 100530, 100570, 100600, 
    100640, 100650, 100670, 100740, 100790, 100820, 100820, 100850, 100910, 
    100920, 100960, 100980, 100950, 100940, 100970, 100980, 100990, 101000, 
    100970, 100930, 100880, 100790, 100720, 100650, 100600, 100530, 100440, 
    100440, 100350, 100290, 100230, 100120, 100090, 100060, 100010, 100020, 
    100000, 100030, 99990, 100000, 100020, 100050, 100050, 100070, 100110, 
    100120, 100100, 100080, 100080, 100060, 100050, 100070, 100090, 100110, 
    100120, 100090, 100060, 100040, 100000, 99980, 99940, 99840, 99820, 
    99730, 99660, 99590, 99550, 99470, 99410, 99370, 99290, 99250, 99250, 
    99200, 99130, 99200, 99250, 99300, 99340, 99320, 99270, 99250, 99250, 
    99250, 99260, 99220, 99170, 99050, 98960, 98870, 98810, 98760, 98720, 
    98700, 98620, 98620, 98660, 98700, 98600, 98650, 98660, 98640, 98630, 
    98590, 98540, 98490, 98480, 98550, 98590, 98590, 98590, 98600, 98620, 
    98720, 98750, 98810, 98860, 98900, 98980, 99100, 99190, 99270, 99370, 
    99480, 99560, 99700, 99810, 99900, 99980, 100080, 100160, 100260, 100320, 
    100350, 100410, 100450, 100500, 100550, 100570, 100600, 100590, 100590, 
    100590, 100590, 100580, 100600, 100590, 100600, 100600, 100630, 100600, 
    100610, 100620, 100600, 100610, 100610, 100600, 100600, 100610, 100610, 
    100600, 100590, 100610, 100600, 100600, 100600, 100610, 100620, 100610, 
    100600, 100600, 100630, 100630, 100650, 100640, 100640, 100650, 100640, 
    100660, 100660, 100650, 100630, 100620, 100680, 100660, 100660, 100660, 
    100660, 100670, 100690, 100700, 100670, 100660, 100650, 100680, 100660, 
    100650, 100670, 100680, 100670, 100700, 100700, 100700, 100720, 100750, 
    100740, 100770, 100790, 100800, 100840, 100860, 100890, 100920, 100940, 
    100950, 100940, 101040, 101130, 101160, 101170, 101230, 101200, 101130, 
    101250, 101370, 101410, 101420, 101390, 101370, 101340, 101300, 101400, 
    101430, 101450, 101500, 101480, 101540, 101560, 101540, 101500, 101540, 
    101560, 101570, 101580, 101620, 101610, 101570, 101540, 101560, 101560, 
    101610, 101610, 101600, 101600, 101600, 101600, 101650, 101640, 101600, 
    101590, 101650, 101630, 101620, 101610, 101640, 101660, 101670, 101800, 
    101830, 101870, 101860, 101920, 101900, 101920, 101900, 101840, 101790, 
    101980, 101990, 101980, 102030, 102030, 102010, 102000, 102010, 102010, 
    101950, 101920, 101830, 101850, 101900, 101940, 101940, 101950, 101930, 
    101920, 101860, 101770, 101770, 101790, 101780, 101760, 101730, 101710, 
    101680, 101680, 101660, 101610, 101550, 101500, 101420, 101300, 101270, 
    101270, 101260, 101310, 101250, 101240, 101220, 101210, 101140, 101100, 
    101060, 101030, 100960, 100960, 100930, 100940, 100950, 100960, 100970, 
    100930, 100910, 100920, 100920, 100940, 100960, 100970, 100980, 100990, 
    101020, 101080, 101110, 101070, 101090, 101090, 101060, 101060, 101040, 
    101040, 101050, 101070, 101090, 101070, 101080, 101090, 101110, 101080, 
    100960, 100980, 100980, 100950, 100980, 101020, 101030, 101060, 101030, 
    101030, 101010, 101000, 101040, 101040, 101030, 101060, 101040, 101070, 
    101080, 101120, 101140, 101150, 101170, 101200, 101210, 101230, 101230, 
    101250, 101270, 101280, 101320, 101360, 101400, 101420, 101420, 101440, 
    101440, 101460, 101510, 101480, 101460, 101480, 101510, 101530, 101610, 
    101610, 101640, 101680, 101730, 101770, 101800, 101820, 101860, 101890, 
    101920, 101960, 102030, 102060, 102060, 102060, 102070, 102110, 102090, 
    102090, 102130, 102140, 102140, 102150, 102200, 102170, 102180, 102190, 
    102160, 102160, 102150, 102190, 102170, 102150, 102140, 102170, 102190, 
    102210, 102210, 102170, 102180, 102170, 102170, 102160, 102150, 102160, 
    102160, 102180, 102180, 102180, 102160, 102180, 102140, 102130, 102110, 
    102090, 102090, 102110, 102100, 102090, 102110, 102120, 102100, 102060, 
    102000, 101960, 101860, 101840, 101840, 101830, 101810, 101780, 101770, 
    101820, 101790, 101810, 101810, 101830, 101850, 101870, 101890, 101910, 
    101940, 101980, 102000, 102000, 102000, 101990, 101970, 101970, 101960, 
    101930, 101910, 101910, 101910, 101900, 101880, 101850, 101850, 101790, 
    101760, 101760, 101760, 101760, 101780, 101810, 101850, 101860, 101890, 
    101890, 101920, 101900, 101910, 101910, 101910, 101900, 101900, 101890, 
    101920, 101920, 101920, 101960, 101950, 101940, 101930, 101920, 101920, 
    101930, 101930, 101930, 101960, 101980, 102010, 102050, 102020, 102000, 
    102020, 102020, 102030, 102030, 102040, 102050, 102070, 102080, 102130, 
    102150, 102150, 102130, 102130, 102140, 102160, 102170, 102180, 102190, 
    102230, 102270, 102310, 102310, 102320, 102340, 102350, 102350, 102360, 
    102370, 102380, 102400, 102410, 102440, 102440, 102440, 102430, 102450, 
    102460, 102460, 102480, 102510, 102490, 102520, 102540, 102580, 102590, 
    102610, 102600, 102620, 102640, 102650, 102660, 102670, 102660, 102660, 
    102700, 102710, 102730, 102720, 102740, 102740, 102760, 102730, 102760, 
    102770, 102770, 102810, 102810, 102850, 102880, 102910, 102910, 102900, 
    102910, 102880, 102860, 102870, 102850, 102880, 102790, 102790, 102810, 
    102840, 102840, 102780, 102740, 102770, 102710, 102690, 102920, 102770, 
    102800, 102790, 102810, 102810, 102790, 102740, 102720, 102680, 102620, 
    102580, 102600, 102590, 102580, 102560, 102530, 102500, 102490, 102460, 
    102420, 102390, 102310, 102300, 102290, 102290, 102260, 102200, 102210, 
    102140, 102110, 102060, 102000, 101830, 101810, 101790, 101690, 101530, 
    101450, 101410, 101380, 101290, 101160, 101100, 101040, 100970, 100890, 
    100850, 100830, 100810, 100830, 100810, 100790, 100790, 100790, 100780, 
    100770, 100780, 100800, 100780, 100790, 100810, 100820, 100860, 100880, 
    100820, 100810, 100870, 100820, 100800, 100800, 100790, 100800, 100810, 
    100800, 100820, 100830, 100820, 100790, 100800, 100810, 100800, 100800, 
    100820, 100820, 100840, 100880, 100870, 100890, 100890, 100930, 100940, 
    100970, 100980, 100990, 101000, 101040, 101060, 101130, 101150, 101190, 
    101220, 101240, 101260, 101310, 101330, 101380, 101410, 101440, 101470, 
    101510, 101570, 101610, 101630, 101640, 101670, 101690, 101720, 101730, 
    101750, 101760, 101760, 101780, 101820, 101830, 101820, 101790, 101780, 
    101760, 101750, 101740, 101710, 101700, 101700, 101750, 101790, 101900, 
    101970, 102010, 102070, 102130, 102220, 102310, 102390, 102450, 102460, 
    102520, 102540, 102580, 102590, 102600, 102580, 102560, 102580, 102550, 
    102520, 102490, 102490, 102450, 102440, 102410, 102340, 102260, 102200, 
    102150, 102090, 102030, 101960, 101930, 101930, 101920, 101930, 101950, 
    101930, 101920, 101930, 101900, 101880, 101870, 101880, 101880, 101860, 
    101850, 101860, 101850, 101850, 101850, 101820, 101780, 101730, 101720, 
    101700, 101660, 101640, 101660, 101650, 101670, 101670, 101640, 101610, 
    101530, 101460, 101410, 101340, 101310, 101270, 101220, 101170, 101130, 
    101110, 101100, 101120, 101090, 101090, 101080, 101070, 101050, 101080, 
    101080, 101100, 101120, 101110, 101120, 101100, 101070, 101080, 101080, 
    101050, 101010, 101020, 101000, 101000, 100980, 101000, 101020, 101000, 
    100980, 100950, 100920, 100880, 100840, 100780, 100770, 100750, 100730, 
    100750, 100740, 100730, 100820, 100890, 100970, 101010, 101080, 101130, 
    101140, 101210, 101250, 101330, 101350, 101360, 101380, 101380, 101400, 
    101450, 101480, 101560, 101590, 101600, 101650, 101700, 101680, 101760, 
    101830, 101860, 101880, 101900, 102010, 102040, 102050, 102120, 102160, 
    102180, 102230, 102240, 102250, 102250, 102260, 102260, 102260, 102260, 
    102270, 102280, 102290, 102260, 102220, 102180, 102150, 102080, 101970, 
    101890, 101800, 101690, 101640, 101560, 101460, 101380, 101280, 101230, 
    101190, 101130, 101080, 101080, 101100, 101120, 101100, 101080, 101100, 
    101120, 101190, 101250, 101320, 101430, 101520, 101600, 101660, 101700, 
    101740, 101780, 101820, 101830, 101850, 101850, 101840, 101820, 101750, 
    101720, 101660, 101620, 101610, 101550, 101510, 101470, 101400, 101330, 
    101270, 101190, 101090, 101000, 100940, 100880, 100810, 100740, 100710, 
    100680, 100640, 100640, 100660, 100630, 100630, 100630, 100670, 100700, 
    100740, 100800, 100850, 100910, 100940, 100990, 101000, 101050, 101140, 
    101180, 101240, 101290, 101360, 101390, 101410, 101450, 101490, 101530, 
    101560, 101590, 101630, 101650, 101670, 101690, 101740, 101750, 101760, 
    101770, 101800, 101810, 101780, 101760, 101790, 101740, 101710, 101710, 
    101730, 101740, 101780, 101810, 101820, 101800, 101830, 101850, 101880, 
    101900, 101930, 101980, 102050, 102100, 102170, 102230, 102290, 102360, 
    102430, 102460, 102550, 102590, 102650, 102710, 102740, 102810, 102840, 
    102950, 103020, 103030, 103040, 103070, 103100, 103140, 103140, 103130, 
    103170, 103220, 103220, 103200, 103200, 103200, 103200, 103190, 103250, 
    103340, 103390, 103430, 103490, 103540, 103580, 103590, 103610, 103630, 
    103650, 103650, 103630, 103590, 103620, 103630, 103620, 103610, 103610, 
    103570, 103540, 103510, 103490, 103460, 103430, 103420, 103420, 103400, 
    103390, 103380, 103340, 103310, 103300, 103270, 103230, 103200, 103150, 
    103120, 103100, 103080, 103070, 103080, 103060, 103010, 102980, 102920, 
    102890, 102820, 102790, 102740, 102690, 102650, 102620, 102570, 102520, 
    102460, 102400, 102330, 102250, 102170, 102090, 102000, 101950, 101880, 
    101830, 101800, 101740, 101660, 101600, 101520, 101440, 101390, 101320, 
    101270, 101210, 101150, 101160, 101150, 101150, 101140, 101120, 101110, 
    101140, 101120, 101140, 101130, 101140, 101160, 101220, 101280, 101320, 
    101370, 101400, 101440, 101480, 101490, 101510, 101520, 101570, 101620, 
    101660, 101720, 101750, 101790, 101800, 101860, 101870, 101870, 101850, 
    101880, 101850, 101880, 101890, 101910, 101950, 101960, 101980, 102000, 
    102000, 102030, 102010, 102050, 102060, 102070, 102070, 102100, 102130, 
    102160, 102170, 102190, 102200, 102210, 102210, 102220, 102220, 102230, 
    102270, 102300, 102310, 102300, 102290, 102270, 102280, 102290, 102280, 
    102290, 102320, 102330, 102360, 102360, 102360, 102340, 102320, 102290, 
    102250, 102230, 102210, 102190, 102180, 102180, 102200, 102220, 102220, 
    102200, 102170, 102070, 102070, 102010, 101970, 101960, 101940, 101920, 
    101880, 101840, 101830, 101790, 101740, 101680, 101610, 101560, 101490, 
    101430, 101370, 101310, 101250, 101200, 101160, 101090, 101030, 100970, 
    100910, 100830, 100750, 100680, 100610, 100530, 100520, 100490, 100430, 
    100380, 100350, 100310, 100290, 100270, 100240, 100250, 100250, 100260, 
    100300, 100340, 100380, 100410, 100450, 100470, 100500, 100520, 100540, 
    100570, 100590, 100640, 100660, 100710, 100740, 100750, 100770, 100800, 
    100820, 100850, 100870, 100870, 100880, 100920, 100950, 100970, 101020, 
    101050, 101080, 101080, 101110, 101120, 101140, 101140, 101150, 101170, 
    101200, 101240, 101260, 101300, 101310, 101310, 101310, 101350, 101380, 
    101380, 101390, 101410, 101440, 101460, 101460, 101450, 101460, 101450, 
    101470, 101460, 101470, 101460, 101430, 101400, 101390, 101390, 101380, 
    101420, 101400, 101370, 101350, 101320, 101270, 101230, 101240, 101210, 
    101190, 101220, 101240, 101230, 101230, 101220, 101200, 101180, 101100, 
    101090, 101090, 101030, 100990, 100950, 100940, 100970, 100970, 100970, 
    100950, 100940, 100930, 100910, 100890, 100860, 100840, 100780, 100680, 
    100750, 100760, 100750, 100730, 100690, 100660, 100650, 100620, 100590, 
    100580, 100560, 100530, 100500, 100470, 100430, 100400, 100360, 100330, 
    100320, 100300, 100300, 100290, 100300, 100320, 100300, 100310, 100300, 
    100300, 100280, 100270, 100220, 100210, 100160, 100130, 100150, 100150, 
    100100, 99970, 99920, 99870, 99810, 99720, 99640, 99620, 99570, 99540, 
    99530, 99520, 99500, 99480, 99440, 99380, 99330, 99250, 99190, 99150, 
    99170, 99200, 99220, 99230, 99230, 99210, 99190, 99170, 99160, 99180, 
    99190, 99230, 99370, 99390, 99470, 99580, 99610, 99630, 99720, 99800, 
    99920, 99960, 100030, 100110, 100160, 100230, 100320, 100360, 100430, 
    100450, 100530, 100590, 100650, 100710, 100760, 100820, 100860, 100940, 
    101010, 101070, 101130, 101190, 101200, 101250, 101290, 101260, 101300, 
    101350, 101430, 101460, 101510, 101580, 101600, 101610, 101630, 101650, 
    101670, 101670, 101660, 101630, 101650, 101640, 101680, 101700, 101720, 
    101720, 101720, 101710, 101650, 101630, 101570, 101500, 101560, 101540, 
    101470, 101540, 101560, 101610, 101560, 101540, 101490, 101490, 101510, 
    101520, 101520, 101520, 101510, 101530, 101500, 101450, 101400, 101380, 
    101320, 101200, 101130, 101080, 101130, 101160, 101130, 101100, 101110, 
    101050, 101040, 101030, 101010, 100950, 100880, 100760, 100740, 100750, 
    100770, 100820, 100850, 100820, 100830, 100820, 100810, 100760, 100760, 
    100740, 100670, 100600, 100570, 100590, 100590, 100570, 100550, 100510, 
    100510, 100470, 100410, 100350, 100310, 100280, 100220, 100200, 100240, 
    100180, 100120, 100120, 100130, 100140, 100160, 100190, 100220, 100220, 
    100270, 100280, 100290, 100350, 100410, 100480, 100560, 100660, 100730, 
    100830, 100910, 101000, 101090, 101170, 101270, 101360, 101420, 101460, 
    101500, 101570, 101600, 101640, 101670, 101700, 101730, 101760, 101850, 
    101890, 101920, 101970, 102000, 102020, 102030, 102020, 102050, 102090, 
    102120, 102160, 102180, 102200, 102220, 102220, 102240, 102240, 102250, 
    102240, 102250, 102240, 102220, 102220, 102210, 102190, 102200, 102190, 
    102180, 102170, 102150, 102120, 102090, 102080, 102050, 102040, 102010, 
    101950, 101910, 101880, 101820, 101770, 101700, 101680, 101640, 101610, 
    101560, 101540, 101470, 101430, 101400, 101380, 101340, 101290, 101240, 
    101180, 101160, 101130, 101120, 101090, 101090, 101060, 101020, 100990, 
    100950, 100920, 100900, 100850, 100820, 100770, 100690, 100670, 100620, 
    100600, 100580, 100560, 100510, 100490, 100440, 100440, 100420, 100420, 
    100440, 100450, 100440, 100420, 100390, 100390, 100370, 100380, 100370, 
    100360, 100370, 100410, 100460, 100500, 100500, 100500, 100500, 100500, 
    100490, 100460, 100430, 100390, 100350, 100350, 100370, 100350, 100350, 
    100330, 100330, 100320, 100310, 100270, 100240, 100230, 100220, 100210, 
    100190, 100170, 100130, 100110, 100070, 100040, 100000, 99980, 99960, 
    99920, 99880, 99870, 99840, 99800, 99800, 99770, 99730, 99680, 99620, 
    99640, 99630, 99590, 99530, 99510, 99540, 99550, 99550, 99500, 99540, 
    99510, 99510, 99510, 99490, 99430, 99390, 99390, 99420, 99440, 99470, 
    99460, 99510, 99540, 99560, 99650, 99690, 99700, 99720, 99680, 99690, 
    99680, 99670, 99720, 99740, 99770, 99800, 99810, 99870, 99880, 99900, 
    99880, 99930, 99950, 99880, 99910, 99990, 100030, 100060, 100110, 100120, 
    100150, 100190, 100220, 100210, 100310, 100410, 100510, 100520, 100540, 
    100530, 100580, 100680, 100780, 100860, 100940, 101000, 101030, 101080, 
    101260, 101270, 101300, 101350, 101390, 101400, 101450, 101460, 101460, 
    101460, 101470, 101470, 101440, 101400, 101360, 101300, 101230, 101170, 
    101130, 101100, 101070, 101060, 101030, 101050, 101020, 100990, 100970, 
    100920, 100880, 100860, 100840, 100830, 100810, 100820, 100830, 100860, 
    100820, 100780, 100780, 100770, 100840, 100780, 100830, 100830, 100750, 
    100700, 100790, 100850, 100820, 100800, 100830, 100910, 100970, 101000, 
    101010, 101050, 101100, 101140, 101170, 101200, 101300, 101380, 101390, 
    101420, 101410, 101440, 101420, 101410, 101440, 101470, 101570, 101620, 
    101640, 101670, 101700, 101700, 101740, 101780, 101790, 101780, 101830, 
    101840, 101830, 101830, 101820, 101850, 101860, 101840, 101850, 101850, 
    101840, 101810, 101780, 101790, 101780, 101710, 101660, 101610, 101570, 
    101490, 101430, 101340, 101260, 101150, 101130, 101080, 101020, 100950, 
    100890, 100810, 100720, 100620, 100470, 100350, 100230, 100130, 100020, 
    99870, 99750, 99630, 99570, 99490, 99440, 99530, 99440, 99380, 99340, 
    99300, 99260, 99240, 99270, 99320, 99330, 99420, 99490, 99560, 99620, 
    99670, 99720, 99800, 99850, 99990, 100110, 100220, 100290, 100390, 
    100460, 100560, 100640, 100660, 100660, 100740, 100760, 100820, 100870, 
    100910, 100920, 100950, 100980, 100980, 100980, 100980, 100960, 100940, 
    100880, 100830, 100810, 100820, 100880, 100920, 100930, 101030, 101030, 
    101020, 101010, 101000, 101000, 101000, 101020, 101010, 101000, 100960, 
    100930, 100880, 100850, 100800, 100730, 100660, 100600, 100540, 100450, 
    100350, 100280, 100180, 100130, 100010, 99880, 99720, 99610, 99480, 
    99390, 99330, 99220, 99100, 99000, 98920, 98880, 98890, 98860, 98780, 
    98720, 98690, 98670, 98640, 98600, 98540, 98550, 98540, 98550, 98530, 
    98510, 98490, 98460, 98470, 98490, 98530, 98560, 98610, 98620, 98650, 
    98660, 98670, 98690, 98790, 98830, 98840, 98890, 98950, 98930, 98970, 
    98970, 99000, 99050, 99050, 99110, 99150, 99190, 99190, 99240, 99230, 
    99250, 99250, 99260, 99280, 99290, 99280, 99260, 99240, 99220, 99220, 
    99240, 99250, 99250, 99240, 99250, 99240, 99220, 99220, 99200, 99160, 
    99120, 99090, 99110, 99100, 99100, 99090, 99080, 99060, 99060, 99040, 
    99040, 99000, 98980, 98980, 99000, 99080, 99160, 99210, 99220, 99230, 
    99250, 99310, 99340, 99410, 99410, 99480, 99490, 99490, 99560, 99660, 
    99670, 99690, 99730, 99770, 99750, 99800, 99810, 99830, 99840, 99880, 
    99880, 99870, 99900, 99910, 99870, 99870, 99830, 99780, 99740, 99710, 
    99740, 99740, 99680, 99670, 99680, 99730, 99760, 99760, 99800, 99830, 
    99860, 99880, 99950, 100020, 100080, 100130, 100190, 100230, 100280, 
    100340, 100380, 100430, 100400, 100400, 100460, 100510, 100570, 100580, 
    100610, 100730, 100800, 100840, 100800, 100770, 100790, 100830, 100840, 
    100870, 100880, 100880, 100850, 100840, 100800, 100770, 100750, 100700, 
    100660, 100620, 100610, 100620, 100610, 100580, 100550, 100510, 100480, 
    100460, 100430, 100430, 100420, 100450, 100490, 100530, 100570, 100590, 
    100610, 100620, 100620, 100620, 100630, 100630, 100580, 100570, 100560, 
    100590, 100560, 100560, 100560, 100560, 100530, 100510, 100480, 100480, 
    100470, 100460, 100430, 100490, 100520, 100560, 100560, 100560, 100570, 
    100570, 100550, 100550, 100560, 100560, 100560, 100540, 100550, 100560, 
    100570, 100570, 100570, 100530, 100540, 100520, 100490, 100450, 100430, 
    100410, 100400, 100470, 100460, 100450, 100440, 100440, 100380, 100410, 
    100290, 100200, 100160, 100140, 99970, 99970, 99820, 99860, 99830, 99780, 
    99650, 99570, 99530, 99530, 99540, 99550, 99510, 99380, 99320, 99300, 
    99340, 99410, 99510, 99550, 99550, 99550, 99540, 99540, 99580, 99550, 
    99530, 99500, 99480, 99480, 99460, 99490, 99460, 99480, 99510, 99510, 
    99530, 99540, 99530, 99570, 99570, 99600, 99600, 99600, 99620, 99630, 
    99640, 99650, 99660, 99680, 99740, 99790, 99820, 99810, 99800, 99820, 
    99870, 99930, 99950, 99980, 100020, 100070, 100090, 100110, 100130, 
    100170, 100210, 100200, 100170, 100200, 100240, 100240, 100230, 100230, 
    100230, 100240, 100230, 100240, 100240, 100200, 100210, 100200, 100180, 
    100180, 100160, 100150, 100130, 100130, 100120, 100080, 100070, 100030, 
    99990, 99950, 99910, 99870, 99820, 99750, 99710, 99650, 99610, 99560, 
    99520, 99440, 99400, 99330, 99270, 99270, 99240, 99200, 99170, 99140, 
    99100, 99070, 99040, 98970, 98950, 98930, 98910, 98890, 98900, 98890, 
    98880, 98850, 98840, 98840, 98810, 98800, 98790, 98800, 98820, 98830, 
    98850, 98860, 98890, 98890, 98910, 98950, 98960, 98980, 99000, 99030, 
    99050, 99070, 99110, 99130, 99180, 99230, 99260, 99280, 99300, 99320, 
    99350, 99400, 99450, 99480, 99520, 99540, 99550, 99570, 99550, 99520, 
    99500, 99460, 99440, 99430, 99410, 99400, 99370, 99350, 99320, 99280, 
    99280, 99250, 99230, 99200, 99180, 99180, 99200, 99230, 99250, 99260, 
    99290, 99320, 99360, 99400, 99460, 99480, 99530, 99580, 99620, 99690, 
    99740, 99770, 99880, 99950, 100010, 100060, 100120, 100180, 100290, 
    100380, 100450, 100530, 100610, 100690, 100720, 100820, 100890, 100940, 
    101000, 101040, 101060, 101080, 101130, 101130, 101120, 101130, 101210, 
    101250, 101250, 101290, 101340, 101360, 101380, 101400, 101390, 101430, 
    101450, 101430, 101400, 101410, 101380, 101410, 101410, 101410, 101540, 
    101590, 101660, 101740, 101840, 101910, 101990, 102070, 102100, 102150, 
    102220, 102280, 102310, 102400, 102410, 102410, 102440, 102440, 102380, 
    102420, 102380, 102270, 102140, 101970, 101840, 101780, 101690, 101430, 
    101270, 101110, 100910, 100730, 100550, 100420, 100300, 100190, 100140, 
    100160, 100140, 100140, 100120, 100060, 99980, 99910, 99810, 99660, 
    99540, 99460, 99440, 99430, 99430, 99360, 99220, 99310, 99450, 99510, 
    99640, 99690, 99750, 99830, 99950, 100050, 100090, 100150, 100180, 
    100310, 100340, 100370, 100400, 100430, 100450, 100510, 100530, 100500, 
    100510, 100500, 100510, 100640, 100730, 100790, 100810, 100930, 101010, 
    101000, 100990, 100940, 100980, 101010, 100960, 100910, 100860, 100830, 
    100830, 100830, 100810, 100780, 100800, 100810, 100850, 100900, 100930, 
    100900, 100930, 100920, 100890, 100880, 100850, 100830, 100830, 100800, 
    100830, 100870, 100870, 100880, 100880, 100880, 100910, 100940, 100890, 
    100850, 100820, 100800, 100820, 100860, 100880, 100870, 100870, 100860, 
    100780, 100750, 100750, 100680, 100660, 100630, 100540, 100550, 100500, 
    100400, 100360, 100320, 100300, 100230, 100150, 100080, 100040, 100000, 
    99980, 99950, 99920, 99880, 99870, 99900, 99920, 99940, 99930, 99920, 
    99900, 99860, 99870, 99930, 99970, 99950, 99950, 99940, 99990, 99980, 
    100010, 100010, 100010, 99990, 100020, 100050, 100070, 100090, 100120, 
    100090, 100110, 100140, 100140, 100130, 100150, 100170, 100160, 100150, 
    100150, 100110, 100080, 100090, 100090, 100050, 100010, 100010, 99970, 
    99940, 99900, 99880, 99860, 99860, 99820, 99790, 99760, 99730, 99710, 
    99680, 99640, 99610, 99580, 99570, 99550, 99530, 99500, 99460, 99410, 
    99400, 99370, 99340, 99300, 99290, 99280, 99270, 99270, 99260, 99280, 
    99310, 99330, 99360, 99360, 99370, 99420, 99460, 99490, 99530, 99550, 
    99590, 99640, 99670, 99680, 99720, 99740, 99740, 99720, 99720, 99740, 
    99740, 99760, 99790, 99800, 99860, 99910, 100040, 100120, 100120, 100200, 
    100270, 100360, 100440, 100520, 100640, 100720, 100810, 100860, 100930, 
    100980, 101020, 101070, 101120, 101180, 101230, 101310, 101350, 101380, 
    101430, 101480, 101570, 101620, 101650, 101680, 101680, 101700, 101730, 
    101770, 101830, 101850, 101890, 101930, 101950, 101960, 102030, 102050, 
    102070, 102090, 102110, 102140, 102170, 102180, 102190, 102190, 102210, 
    102250, 102230, 102220, 102240, 102210, 102230, 102230, 102210, 102190, 
    102150, 102110, 102040, 102010, 101940, 101890, 101820, 101750, 101720, 
    101670, 101590, 101500, 101450, 101400, 101360, 101320, 101260, 101220, 
    101180, 101190, 101230, 101230, 101230, 101220, 101220, 101220, 101210, 
    101150, 101080, 101020, 100950, 100890, 100770, 100720, 100620, 100560, 
    100460, 100380, 100340, 100260, 100220, 100180, 100130, 100100, 100040, 
    99970, 99920, 99830, 99770, 99730, 99660, 99630, 99590, 99580, 99600, 
    99520, 99520, 99510, 99530, 99590, 99610, 99680, 99670, 99610, 99640, 
    99590, 99660, 99680, 99690, 99700, 99680, 99690, 99670, 99680, 99690, 
    99670, 99660, 99630, 99620, 99600, 99580, 99590, 99570, 99570, 99540, 
    99530, 99530, 99530, 99530, 99540, 99560, 99580, 99580, 99600, 99640, 
    99670, 99730, 99760, 99780, 99840, 99870, 99940, 99980, 99960, 100030, 
    100110, 100150, 100180, 100240, 100240, 100220, 100240, 100260, 100310, 
    100310, 100340, 100350, 100360, 100380, 100420, 100430, 100410, 100400, 
    100390, 100400, 100390, 100400, 100390, 100400, 100380, 100370, 100350, 
    100330, 100330, 100320, 100330, 100330, 100330, 100320, 100310, 100300, 
    100270, 100230, 100190, 100140, 100070, 100010, 99940, 99930, 99930, 
    99960, 99960, 99970, 100010, 100060, 100090, 100120, 100150, 100190, 
    100200, 100250, 100320, 100380, 100450, 100530, 100600, 100630, 100660, 
    100680, 100680, 100660, 100650, 100640, 100650, 100640, 100670, 100680, 
    100700, 100720, 100690, 100680, 100670, 100640, 100620, 100590, 100550, 
    100490, 100460, 100430, 100390, 100330, 100250, 100140, 100010, 99810, 
    99580, 99350, 99180, 98970, 98780, 98640, 98450, 98270, 98120, 97940, 
    97740, 97540, 97340, 97110, 96890, 96660, 96430, 96310, 96220, 96130, 
    96120, 96120, 96160, 96210, 96410, 96580, 96790, 96940, 97100, 97170, 
    97330, 97510, 97780, 97980, 98000, 98100, 98240, 98450, 98540, 98600, 
    98680, 98790, 98870, 98960, 99010, 99060, 99040, 99050, 99050, 99030, 
    99020, 98990, 98940, 98920, 98880, 98830, 98820, 98780, 98700, 98670, 
    98610, 98610, 98560, 98580, 98560, 98550, 98550, 98580, 98620, 98620, 
    98670, 98690, 98790, 98800, 98880, 98990, 99030, 99100, 99180, 99270, 
    99380, 99560, 99620, 99670, 99730, 99810, 99950, 100010, 100050, 100080, 
    100180, 100250, 100320, 100380, 100430, 100430, 100460, 100490, 100510, 
    100520, 100570, 100610, 100600, 100550, 100560, 100550, 100550, 100510, 
    100480, 100420, 100410, 100410, 100400, 100390, 100400, 100360, 100320, 
    100340, 100320, 100280, 100260, 100230, 100240, 100220, 100220, 100240, 
    100270, 100310, 100340, 100360, 100430, 100480, 100510, 100540, 100600, 
    100640, 100740, 100840, 100900, 101000, 101090, 101140, 101190, 101250, 
    101280, 101330, 101370, 101410, 101440, 101490, 101530, 101570, 101600, 
    101610, 101660, 101680, 101700, 101700, 101740, 101790, 101820, 101830, 
    101860, 101860, 101890, 101850, 101850, 101850, 101880, 101890, 101880, 
    101870, 101850, 101880, 101920, 101920, 101910, 101930, 101900, 101880, 
    101890, 101920, 101930, 101940, 101960, 101990, 102010, 102030, 102060, 
    102110, 102170, 102190, 102150, 102140, 102130, 102140, 102150, 102190, 
    102220, 102210, 102230, 102230, 102220, 102230, 102230, 102220, 102230, 
    102240, 102250, 102190, 102170, 102170, 102180, 102150, 102110, 102110, 
    102130, 102110, 102060, 102000, 102000, 102010, 101970, 101940, 101880, 
    101810, 101810, 101800, 101790, 101790, 101760, 101810, 101840, 101840, 
    101820, 101810, 101800, 101800, 101790, 101900, 101830, 101730, 101710, 
    101620, 101640, 101610, 101610, 101570, 101520, 101520, 101440, 101400, 
    101390, 101400, 101380, 101400, 101390, 101410, 101400, 101430, 101460, 
    101490, 101520, 101540, 101570, 101620, 101660, 101710, 101760, 101850, 
    101910, 102000, 102070, 102120, 102180, 102220, 102260, 102290, 102330, 
    102370, 102400, 102430, 102450, 102470, 102490, 102480, 102450, 102410, 
    102360, 102290, 102270, 102230, 102170, 102150, 102080, 102030, 101940, 
    101930, 101950, 101870, 101910, 101960, 101980, 101930, 101980, 102030, 
    102060, 102070, 102070, 102070, 102050, 102040, 102030, 102010, 102020, 
    102010, 102020, 102000, 101990, 101970, 101980, 101970, 101980, 101980, 
    101970, 101950, 101930, 101950, 101950, 101950, 101940, 101940, 101930, 
    101920, 101940, 101950, 101960, 101960, 101970, 101980, 102000, 101990, 
    102010, 102020, 102010, 102000, 102000, 101980, 101970, 101970, 101990, 
    101990, 102000, 102020, 102030, 102050, 102040, 102070, 102090, 102110, 
    102160, 102180, 102200, 102230, 102270, 102310, 102340, 102350, 102380, 
    102390, 102400, 102420, 102420, 102430, 102470, 102480, 102500, 102520, 
    102530, 102540, 102510, 102510, 102510, 102490, 102490, 102480, 102480, 
    102470, 102460, 102470, 102470, 102470, 102440, 102400, 102380, 102360, 
    102340, 102360, 102340, 102330, 102330, 102360, 102350, 102340, 102310, 
    102280, 102270, 102260, 102250, 102180, 102170, 102180, 102160, 102170, 
    102150, 102130, 102120, 102100, 102110, 102090, 102080, 102060, 102060, 
    102070, 102070, 102070, 102090, 102090, 102080, 102120, 102120, 102130, 
    102150, 102140, 102150, 102140, 102150, 102140, 102170, 102190, 102210, 
    102210, 102220, 102220, 102230, 102240, 102290, 102260, 102300, 102340, 
    102350, 102350, 102390, 102400, 102420, 102420, 102450, 102450, 102480, 
    102470, 102470, 102440, 102440, 102440, 102450, 102490, 102480, 102460, 
    102530, 102490, 102550, 102550, 102570, 102620, 102630, 102640, 102620, 
    102610, 102610, 102600, 102570, 102570, 102530, 102540, 102530, 102500, 
    102500, 102460, 102450, 102430, 102420, 102400, 102350, 102330, 102310, 
    102280, 102190, 102140, 102110, 102060, 101990, 101940, 101900, 101840, 
    101780, 101740, 101670, 101600, 101520, 101410, 101300, 101210, 101110, 
    100990, 100870, 100790, 100870, 100990, 101050, 101070, 101040, 101080, 
    101170, 101170, 101200, 101210, 101260, 101310, 101300, 101310, 101290, 
    101290, 101280, 101270, 101250, 101250, 101220, 101200, 101180, 101160, 
    101130, 101110, 101080, 101080, 101060, 101030, 101020, 100990, 100970, 
    100940, 100920, 100870, 100850, 100840, 100830, 100820, 100800, 100790, 
    100770, 100750, 100780, 100770, 100770, 100770, 100770, 100770, 100790, 
    100780, 100790, 100810, 100800, 100790, 100830, 100820, 100790, 100810, 
    100810, 100810, 100820, 100810, 100810, 100820, 100800, 100810, 100790, 
    100770, 100760, 100740, 100730, 100730, 100730, 100730, 100720, 100720, 
    100720, 100700, 100700, 100700, 100700, 100680, 100660, 100640, 100640, 
    100640, 100640, 100640, 100640, 100630, 100610, 100570, 100540, 100510, 
    100520, 100530, 100540, 100550, 100550, 100610, 100640, 100700, 100770, 
    100820, 100850, 100850, 100920, 100960, 101000, 101030, 101060, 101080, 
    101080, 101090, 101100, 101120, 101140, 101140, 101150, 101160, 101180, 
    101200, 101230, 101230, 101250, 101280, 101280, 101270, 101270, 101250, 
    101260, 101270, 101260, 101260, 101270, 101280, 101260, 101260, 101260, 
    101250, 101230, 101210, 101180, 101160, 101160, 101150, 101120, 101100, 
    101120, 101120, 101100, 101110, 101140, 101140, 101180, 101240, 101270, 
    101270, 101280, 101290, 101270, 101270, 101280, 101260, 101260, 101260, 
    101240, 101240, 101250, 101250, 101250, 101260, 101260, 101290, 101310, 
    101340, 101360, 101360, 101350, 101330, 101300, 101280, 101250, 101220, 
    101180, 101130, 101110, 101070, 101030, 101010, 100970, 100930, 100890, 
    100840, 100810, 100790, 100730, 100710, 100690, 100670, 100640, 100610, 
    100570, 100540, 100490, 100420, 100320, 100220, 100120, 100040, 99940, 
    99800, 99720, 99630, 99590, 99500, 99380, 99360, 99310, 99270, 99230, 
    99220, 99190, 99210, 99210, 99220, 99250, 99230, 99290, 99340, 99390, 
    99410, 99470, 99530, 99620, 99750, 99880, 99990, 100080, 100110, 100200, 
    100290, 100340, 100410, 100490, 100600, 100680, 100730, 100810, 100890, 
    100950, 100990, 101050, 101130, 101190, 101270, 101330, 101350, 101380, 
    101400, 101410, 101420, 101460, 101480, 101510, 101550, 101580, 101600, 
    101630, 101620, 101620, 101570, 101530, 101470, 101410, 101360, 101330, 
    101300, 101270, 101230, 101200, 101170, 101130, 101110, 101110, 101090, 
    101060, 101070, 101080, 101100, 101110, 101090, 101060, 101030, 100990, 
    100960, 100920, 100880, 100840, 100800, 100750, 100690, 100640, 100560, 
    100540, 100490, 100440, 100370, 100330, 100280, 100200, 100130, 100060, 
    100020, 100040, 100040, 100080, 100110, 100180, 100210, 100250, 100280, 
    100330, 100390, 100470, 100570, 100630, 100670, 100710, 100730, 100820, 
    100880, 100940, 100990, 101070, 101100, 101140, 101180, 101240, 101330, 
    101380, 101450, 101490, 101520, 101560, 101570, 101600, 101660, 101720, 
    101770, 101800, 101850, 101900, 101940, 102000, 102010, 102050, 102060, 
    102030, 102040, 102090, 102140, 102200, 102250, 102290, 102340, 102380, 
    102400, 102430, 102460, 102460, 102500, 102520, 102510, 102520, 102500, 
    102500, 102560, 102660, 102590, 102600, 102600, 102640, 102650, 102670, 
    102650, 102650, 102640, 102630, 102600, 102600, 102590, 102630, 102650, 
    102610, 102600, 102620, 102570, 102650, 102660, 102680, 102640, 102600, 
    102560, 102570, 102580, 102600, 102620, 102620, 102630, 102650, 102700, 
    102770, 102720, 102800, 102840, 102880, 102900, 102930, 102940, 102940, 
    102970, 103000, 103040, 103080, 103100, 103120, 103180, 103230, 103250, 
    103270, 103270, 103270, 103300, 103310, 103310, 103310, 103310, 103330, 
    103310, 103300, 103290, 103290, 103280, 103250, 103220, 103240, 103210, 
    103210, 103210, 103190, 103190, 103180, 103160, 103100, 103090, 103090, 
    103080, 103050, 103040, 103010, 102960, 102930, 102870, 102770, 102690, 
    102630, 102540, 102470, 102410, 102390, 102350, 102310, 102300, 102290, 
    102300, 102310, 102330, 102350, 102340, 102340, 102370, 102400, 102370, 
    102400, 102410, 102400, 102370, 102390, 102350, 102300, 102280, 102270, 
    102240, 102250, 102240, 102240, 102240, 102220, 102220, 102200, 102210, 
    102210, 102210, 102200, 102200, 102210, 102230, 102250, 102250, 102250, 
    102250, 102230, 102210, 102200, 102140, 102120, 102120, 102100, 102090, 
    102040, 102000, 101990, 101940, 101920, 101880, 101860, 101810, 101790, 
    101800, 101800, 101790, 101790, 101790, 101780, 101780, 101780, 101760, 
    101730, 101690, 101660, 101660, 101660, 101630, 101590, 101570, 101550, 
    101530, 101500, 101460, 101440, 101450, 101460, 101460, 101480, 101480, 
    101490, 101480, 101450, 101440, 101440, 101450, 101400, 101390, 101380, 
    101390, 101430, 101450, 101490, 101490, 101510, 101500, 101520, 101500, 
    101490, 101510, 101500, 101510, 101560, 101600, 101620, 101620, 101650, 
    101650, 101660, 101640, 101620, 101640, 101660, 101670, 101680, 101700, 
    101710, 101720, 101740, 101780, 101790, 101790, 101800, 101800, 101800, 
    101800, 101810, 101840, 101860, 101840, 101830, 101800, 101770, 101730, 
    101690, 101660, 101620, 101570, 101540, 101500, 101490, 101440, 101400, 
    101380, 101360, 101340, 101350, 101330, 101340, 101370, 101400, 101410, 
    101420, 101440, 101480, 101510, 101550, 101570, 101610, 101670, 101710, 
    101760, 101830, 101900, 101980, 102040, 102080, 102140, 102170, 102200, 
    102240, 102310, 102380, 102430, 102490, 102530, 102580, 102620, 102660, 
    102690, 102710, 102710, 102710, 102700, 102690, 102690, 102710, 102720, 
    102690, 102680, 102670, 102650, 102660, 102630, 102620, 102610, 102610, 
    102600, 102590, 102580, 102560, 102530, 102490, 102460, 102430, 102390, 
    102360, 102320, 102250, 102210, 102170, 102160, 102120, 102080, 102040, 
    102000, 101960, 101920, 101880, 101870, 101860, 101860, 101850, 101850, 
    101860, 101850, 101840, 101870, 101870, 101880, 101880, 101860, 101860, 
    101860, 101890, 101900, 101910, 101900, 101920, 101930, 101930, 101930, 
    101930, 101930, 101950, 101990, 102000, 102000, 101990, 101990, 102010, 
    102000, 101980, 101950, 101910, 101870, 101830, 101800, 101760, 101700, 
    101680, 101630, 101620, 101580, 101550, 101500, 101460, 101420, 101400, 
    101420, 101420, 101420, 101400, 101380, 101350, 101330, 101330, 101310, 
    101320, 101340, 101380, 101470, 101530, 101590, 101670, 101710, 101740, 
    101760, 101820, 101860, 101920, 101980, 102030, 102100, 102170, 102240, 
    102260, 102320, 102370, 102400, 102420, 102440, 102450, 102470, 102480, 
    102470, 102500, 102500, 102490, 102480, 102460, 102420, 102410, 102390, 
    102340, 102290, 102250, 102210, 102170, 102120, 102050, 102020, 101950, 
    101910, 101830, 101770, 101690, 101630, 101560, 101510, 101480, 101450, 
    101430, 101400, 101400, 101400, 101430, 101460, 101470, 101470, 101480, 
    101510, 101530, 101570, 101580, 101610, 101620, 101630, 101620, 101620, 
    101610, 101570, 101550, 101520, 101520, 101510, 101490, 101460, 101430, 
    101390, 101380, 101350, 101340, 101330, 101320, 101350, 101350, 101390, 
    101420, 101440, 101450, 101470, 101500, 101490, 101480, 101470, 101470, 
    101490, 101490, 101490, 101470, 101420, 101380, 101340, 101290, 101260, 
    101220, 101190, 101160, 101130, 101100, 101120, 101110, 101080, 101030, 
    100980, 100910, 100840, 100770, 100720, 100660, 100600, 100560, 100500, 
    100470, 100420, 100410, 100390, 100390, 100370, 100330, 100300, 100270, 
    100240, 100220, 100180, 100150, 100120, 100080, 100040, 100000, 99950, 
    99900, 99830, 99810, 99810, 99830, 99840, 99870, 99900, 99960, 100010, 
    100040, 100160, 100250, 100320, 100400, 100390, 100340, 100360, 100390, 
    100490, 100550, 100620, 100690, 100800, 100930, 101010, 101060, 101170, 
    101270, 101330, 101350, 101370, 101380, 101470, 101530, 101550, 101590, 
    101610, 101570, 101600, 101590, 101610, 101590, 101610, 101550, 101550, 
    101530, 101510, 101490, 101440, 101430, 101390, 101360, 101290, 101300, 
    101260, 101220, 101170, 101150, 101130, 101140, 101130, 101130, 101150, 
    101160, 101170, 101190, 101240, 101260, 101280, 101290, 101280, 101280, 
    101300, 101360, 101350, 101320, 101330, 101330, 101330, 101300, 101260, 
    101230, 101200, 101150, 101100, 101080, 101050, 101010, 100990, 101000, 
    100970, 100920, 100900, 100860, 100810, 100780, 100790, 100760, 100690, 
    100710, 100710, 100710, 100700, 100680, 100660, 100670, 100680, 100680, 
    100670, 100700, 100720, 100770, 100810, 100900, 100980, 101060, 101120, 
    101180, 101260, 101340, 101390, 101430, 101490, 101490, 101580, 101660, 
    101700, 101740, 101780, 101800, 101790, 101850, 101860, 101850, 101870, 
    101900, 101920, 101950, 101970, 101970, 101950, 101920, 101900, 101920, 
    101920, 101900, 101930, 101950, 101930, 101900, 101880, 101830, 101830, 
    101830, 101810, 101810, 101800, 101770, 101760, 101750, 101730, 101730, 
    101740, 101760, 101790, 101800, 101800, 101790, 101830, 101840, 101850, 
    101870, 101910, 101940, 101980, 102010, 102040, 102070, 102070, 102080, 
    102080, 102100, 102120, 102190, 102210, 102270, 102300, 102320, 102350, 
    102340, 102330, 102350, 102370, 102370, 102400, 102390, 102390, 102380, 
    102380, 102380, 102370, 102330, 102320, 102320, 102310, 102290, 102290, 
    102310, 102320, 102300, 102330, 102310, 102310, 102290, 102310, 102300, 
    102300, 102300, 102310, 102320, 102330, 102340, 102340, 102340, 102340, 
    102350, 102360, 102380, 102370, 102370, 102390, 102410, 102420, 102440, 
    102440, 102450, 102450, 102450, 102430, 102420, 102430, 102420, 102400, 
    102380, 102360, 102350, 102330, 102330, 102310, 102320, 102310, 102300, 
    102290, 102290, 102300, 102300, 102290, 102270, 102280, 102280, 102260, 
    102260, 102260, 102250, 102240, 102240, 102210, 102190, 102160, 102150, 
    102130, 102110, 102100, 102110, 102090, 102070, 102080, 102070, 102030, 
    102030, 102060, 102060, 102060, 102050, 102050, 102070, 102080, 102080, 
    102070, 102060, 102050, 102040, 102030, 102030, 102030, 102000, 102000, 
    102010, 102010, 102000, 102000, 102030, 102030, 102020, 102040, 102040, 
    102040, 102030, 102030, 102030, 102040, 102020, 102000, 101980, 101980, 
    101990, 101980, 101970, 101960, 101930, 101940, 101940, 101920, 101920, 
    101920, 101900, 101890, 101890, 101900, 101890, 101880, 101870, 101860, 
    101860, 101830, 101810, 101800, 101760, 101750, 101730, 101730, 101710, 
    101670, 101650, 101630, 101610, 101580, 101550, 101520, 101490, 101470, 
    101470, 101460, 101450, 101450, 101420, 101410, 101390, 101380, 101360, 
    101350, 101330, 101320, 101320, 101320, 101310, 101300, 101280, 101230, 
    101210, 101190, 101230, 101190, 101160, 101130, 101120, 101120, 101140, 
    101110, 101060, 101050, 101040, 101030, 101010, 100990, 101010, 101020, 
    101020, 101020, 101000, 101000, 101010, 101050, 101070, 101090, 101110, 
    101120, 101140, 101160, 101190, 101230, 101240, 101250, 101280, 101300, 
    101290, 101320, 101350, 101360, 101370, 101390, 101420, 101460, 101480, 
    101510, 101540, 101560, 101560, 101620, 101680, 101710, 101740, 101760, 
    101790, 101850, 101870, 101890, 101940, 101950, 101980, 102000, 102000, 
    102000, 102000, 102010, 102010, 102030, 102010, 102010, 102010, 102000, 
    101990, 101970, 101960, 101930, 101920, 101940, 101930, 101930, 101950, 
    101940, 101930, 101900, 101880, 101880, 101880, 101840, 101800, 101780, 
    101790, 101760, 101740, 101730, 101710, 101690, 101670, 101640, 101610, 
    101610, 101590, 101600, 101610, 101600, 101610, 101610, 101610, 101620, 
    101640, 101640, 101660, 101660, 101700, 101730, 101760, 101790, 101820, 
    101830, 101850, 101860, 101870, 101890, 101910, 101920, 101940, 101950, 
    101980, 102020, 102070, 102110, 102110, 102110, 102140, 102150, 102150, 
    102160, 102160, 102160, 102170, 102170, 102190, 102200, 102200, 102160, 
    102160, 102160, 102150, 102140, 102120, 102130, 102140, 102150, 102160, 
    102140, 102150, 102150, 102120, 102140, 102130, 102120, 102090, 102090, 
    102080, 102120, 102120, 102130, 102150, 102160, 102180, 102180, 102200, 
    102240, 102280, 102330, 102390, 102440, 102500, 102510, 102550, 102560, 
    102580, 102560, 102590, 102580, 102620, 102650, 102630, 102660, 102670, 
    102690, 102680, 102690, 102710, 102710, 102770, 102760, 102790, 102820, 
    102830, 102850, 102900, 102910, 102900, 102960, 102980, 102940, 102920, 
    102950, 102950, 102920, 102950, 102920, 102900, 102840, 102820, 102770, 
    102710, 102610, 102590, 102540, 102440, 102380, 102320, 102280, 102230, 
    102180, 102110, 102020, 101970, 101960, 101940, 101910, 101850, 101860, 
    101800, 101820, 101810, 101800, 101810, 101800, 101780, 101790, 101750, 
    101710, 101710, 101690, 101670, 101640, 101600, 101530, 101430, 101330, 
    101310, 101220, 101050, 100920, 100840, 100760, 100700, 100630, 100610, 
    100590, 100550, 100560, 100520, 100550, 100580, 100640, 100720, 100760, 
    100710, 100770, 100770, 100780, 100750, 100790, 100780, 100760, 100740, 
    100710, 100670, 100650, 100610, 100610, 100570, 100560, 100530, 100530, 
    100540, 100510, 100540, 100570, 100620, 100630, 100640, 100680, 100710, 
    100730, 100770, 100790, 100820, 100860, 100900, 100910, 100890, 100910, 
    100910, 100930, 100940, 100960, 100980, 101020, 101050, 101050, 101070, 
    101080, 101090, 101080, 101080, 101140, 101180, 101160, 101220, 101250, 
    101290, 101300, 101290, 101320, 101330, 101330, 101320, 101320, 101350, 
    101350, 101340, 101360, 101400, 101400, 101390, 101380, 101440, 101440, 
    101490, 101490, 101510, 101560, 101570, 101560, 101550, 101580, 101650, 
    101670, 101700, 101700, 101700, 101730, 101810, 101860, 101910, 101970, 
    102030, 102080, 102100, 102140, 102180, 102190, 102230, 102300, 102310, 
    102360, 102380, 102410, 102430, 102420, 102410, 102410, 102390, 102370, 
    102380, 102340, 102340, 102310, 102290, 102270, 102220, 102200, 102160, 
    102150, 102100, 102100, 102120, 102130, 102160, 102170, 102160, 102100, 
    102070, 102010, 101950, 101930, 101880, 101860, 101810, 101780, 101750, 
    101730, 101680, 101650, 101600, 101560, 101520, 101470, 101450, 101410, 
    101380, 101380, 101380, 101390, 101380, 101390, 101410, 101380, 101370, 
    101350, 101350, 101350, 101350, 101370, 101380, 101370, 101350, 101400, 
    101410, 101440, 101440, 101480, 101530, 101520, 101570, 101610, 101630, 
    101660, 101690, 101730, 101750, 101760, 101760, 101770, 101770, 101800, 
    101800, 101830, 101840, 101840, 101830, 101840, 101830, 101840, 101820, 
    101830, 101820, 101820, 101850, 101860, 101820, 101830, 101810, 101790, 
    101720, 101730, 101720, 101680, 101610, 101550, 101500, 101500, 101460, 
    101390, 101410, 101430, 101440, 101450, 101450, 101480, 101440, 101470, 
    101490, 101530, 101510, 101510, 101500, 101480, 101470, 101460, 101460, 
    101460, 101460, 101460, 101470, 101480, 101470, 101460, 101450, 101440, 
    101400, 101380, 101370, 101360, 101360, 101340, 101320, 101320, 101330, 
    101340, 101380, 101370, 101380, 101390, 101390, 101420, 101460, 101530, 
    101570, 101630, 101680, 101720, 101720, 101760, 101830, 101860, 101860, 
    101900, 101950, 101980, 102040, 102080, 102130, 102150, 102150, 102160, 
    102150, 102130, 102090, 102080, 102050, 102020, 102000, 101940, 101890, 
    101850, 101800, 101710, 101650, 101570, 101500, 101390, 101300, 101220, 
    101170, 101120, 101060, 100970, 100920, 100880, 100850, 100800, 100750, 
    100710, 100690, 100660, 100630, 100600, 100590, 100560, 100490, 100440, 
    100410, 100380, 100340, 100260, 100220, 100240, 100220, 100230, 100250, 
    100280, 100310, 100290, 100280, 100260, 100350, 100380, 100390, 100420, 
    100460, 100490, 100510, 100590, 100600, 100660, 100740, 100790, 100840, 
    100860, 100890, 100900, 100980, 101040, 101060, 101110, 101130, 101130, 
    101180, 101190, 101200, 101180, 101170, 101180, 101180, 101200, 101200, 
    101210, 101240, 101210, 101210, 101210, 101190, 101200, 101190, 101190, 
    101190, 101170, 101190, 101180, 101160, 101140, 101130, 101110, 101120, 
    101080, 101050, 101050, 101060, 101060, 101070, 101080, 101070, 101060, 
    101040, 101050, 101050, 101070, 101080, 101080, 101090, 101110, 101120, 
    101160, 101180, 101210, 101210, 101200, 101200, 101220, 101220, 101230, 
    101260, 101260, 101270, 101270, 101260, 101260, 101260, 101270, 101270, 
    101290, 101290, 101290, 101300, 101330, 101360, 101380, 101400, 101410, 
    101430, 101430, 101430, 101450, 101450, 101450, 101440, 101460, 101460, 
    101470, 101480, 101480, 101470, 101470, 101480, 101470, 101470, 101470, 
    101470, 101480, 101500, 101520, 101520, 101510, 101500, 101480, 101470, 
    101450, 101420, 101390, 101380, 101350, 101330, 101290, 101250, 101230, 
    101220, 101200, 101160, 101140, 101100, 101040, 101000, 100960, 100930, 
    100900, 100860, 100820, 100780, 100740, 100690, 100670, 100630, 100580, 
    100520, 100500, 100490, 100440, 100410, 100380, 100350, 100320, 100270, 
    100230, 100200, 100200, 100190, 100190, 100190, 100190, 100160, 100140, 
    100140, 100120, 100120, 100110, 100100, 100080, 100090, 100080, 100080, 
    100070, 100070, 100070, 100050, 100020, 100010, 100020, 100020, 100020, 
    100010, 100030, 100030, 100030, 100020, 100010, 100010, 100020, 100020, 
    100010, 100000, 99990, 99970, 99960, 99930, 99920, 99910, 99910, 99880, 
    99880, 99900, 99920, 99970, 100000, 100040, _, _, 100180, 100240, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 101450, 101490, _, 
    101520, 101540, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    101630, 101600, 101570, 101560, 101560, _, _, _, 101490, _, 101500, 
    101490, 101520, 101540, 101520, 101530, _, _, _, 101520, 101490, 101510, 
    101520, 101550, 101600, 101650, 101710, 101790, 101830, 101820, 101870, 
    101920, 101920, 101930, 101970, 102070, 102070, 102120, 102160, 102190, 
    102240, 102270, 102280, 102260, 102230, _, _, _, 102270, 102290, 102290, 
    102330, 102320, 102290, 102280, 102220, 102230, 102220, 102140, 102140, 
    102110, 102070, 102030, _, _, _, _, 101760, 101650, 101600, 101560, 
    101480, 101420, 101370, 101350, 101340, 101360, 101290, 101260, 101190, 
    101180, 101170, _, _, _, _, _, _, 101230, 101260, 101280, _, 101360, _, 
    101440, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 102160, 102190, _, 
    102200, 102210, 102180, _, _, _, _, _, 102170, 102150, 102150, 102140, 
    102130, 102080, 102050, 102060, 102040, 102030, _, _, _, _, _, _, _, _, 
    101980, 101960, _, 101910, 101900, _, 101910, 101910, 101900, 101890, _, 
    _, 101830, 101800, _, _, 101710, 101700, 101680, 101650, 101620, _, 
    101550, 101530, _, _, _, _, 101360, 101350, 101310, 101290, 101260, 
    101230, 101210, 101210, 101220, 101180, _, _, 101120, 101140, 101140, 
    101120, _, 101120, _, _, _, _, _, _, _, 100990, 100980, 101000, 100990, 
    100970, 100940, 100900, 100900, 100910, 100910, 100880, 100870, 100880, 
    100870, 100860, 100850, 100860, 100850, 100850, 100840, 100840, 100800, 
    100780, 100810, 100820, 100810, 100810, 100800, 100770, 100760, 100740, 
    100740, 100740, 100730, 100730, 100720, 100720, 100740, 100740, 100710, 
    100640, 100650, 100650, 100650, 100660, 100640, 100670, 100710, 100760, 
    100760, 100840, 100880, 100910, 100960, 100990, 101020, 101040, 101070, 
    101020, 101020, 101030, 100980, 101030, 101070, 101060, 101060, 101050, 
    101040, 101020, 101010, 100990, 100970, 100960, 101030, 101050, 101060, 
    101030, 101050, 101090, 101090, 101080, 101100, 101040, 101050, 101050, 
    101050, 101040, 101030, 101010, 100960, 100900, 100840, 100830, 100780, 
    100770, 100780, 100760, 100760, 100760, 100770, 100760, 100720, 100700, 
    100690, 100670, 100650, 100620, 100590, 100580, 100550, 100560, 100560, 
    100540, 100510, 100510, 100480, 100500, 100530, 100560, 100590, 100610, 
    100610, 100530, 100510, 100520, _, _, 100640, 100640, _, _, _, _, _, _, 
    _, _, _, 100860, 100890, 100920, 100950, 101000, 101030, 101090, 101120, 
    101150, 101190, 101210, 101240, 101260, 101280, 101270, 101290, 101330, 
    _, _, _, _, _, _, _, 101360, 101310, _, _, 101310, 101290, 101290, 
    101340, _, 101310, 101280, 101270, 101260, _, 101200, 101180, 101180, 
    101180, _, _, 101080, 101090, 101090, 101090, 101040, 101010, 101000, 
    100960, _, 100910, 100880, 100830, 100820, _, 100750, 100710, 100670, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 99690, 99660, 99660, 99680, 99730, 
    99790, 99840, 99940, 99980, 100010, 100050, _, _, _, _, _, 100110, 
    100140, _, 100230, 100290, 100350, 100370, 100400, _, _, 100530, 100540, 
    100590, 100630, 100660, 100680, _, 100740, _, _, _, _, _, _, _, _, 
    100780, 100780, 100790, _, 100850, 100850, 100850, 100860, _, 100850, _, 
    _, 101080, 101140, 101170, 101190, 101250, 101290, 101300, 101340, _, _, 
    _, 101540, 101630, 101670, 101720, 101780, 101800, 101810, _, _, _, 
    101910, 101950, 101970, 102000, 102050, 102060, 102080, 102090, 102080, 
    _, _, 102090, 102100, 102120, 102130, 102120, 102120, 102130, 102120, 
    102100, _, 102080, 102080, 102090, 102080, 102080, 102100, 102110, 
    102130, _, 102150, 102150, 102130, 102120, 102120, 102140, 102140, 
    102140, _, _, _, _, _, 102060, 102050, 101960, 101930, 101850, 101850, 
    101820, 101840, 101830, 101800, 101820, _, _, 101720, _, 101680, 101660, 
    101630, 101610, 101550, 101510, 101470, _, 101380, 101330, 101260, 
    101220, 101160, 101140, 101110, 101110, _, 101090, 101060, 101020, 
    100980, 100910, 100840, 100760, 100670, _, 100550, 100510, _, 100400, 
    100360, _, _, 100260, 100250, 100240, _, 100260, 100290, 100310, 100360, 
    100410, 100480, 100490, 100500, 100520, 100510, 100490, 100500, 100510, 
    100520, 100510, 100540, 100580, 100580, 100600, 100620, 100660, 100690, 
    100750, 100750, 100770, 100810, 100850, 100920, 100970, 100980, 101000, 
    101030, 101010, 101020, 101010, 100990, 100940, 100850, 100840, 100790, 
    100740, 100690, 100660, 100620, 100590, 100560, 100540, 100560, 100590, 
    100610, 100610, 100610, 100610, 100630, 100640, 100620, 100620, 100600, 
    100590, 100560, 100570, 100570, 100560, 100620, 100650, 100610, 100630, 
    100610, 100600, 100610, 100610, _, 100590, 100590, 100570, 100570, 
    100570, 100590, 100620, 100650, 100660, 100700, 100730, 100770, 100820, 
    100860, 100940, 101020, 101080, 101090, 101130, 101100, 101210, 101310, 
    101320, 101370, 101440, 101480, _, 101530, 101580, 101620, 101670, 
    101670, 101690, 101700, 101700, 101710, _, _, _, 101700, 101710, 101720, 
    101710, 101700, 101680, 101670, 101680, _, _, _, 101610, 101610, 101620, 
    101610, 101600, 101570, 101560, 101530, 101510, _, _, _, _, _, _, _, _, 
    _, _, 101350, 101330, _, 101320, 101310, 101330, 101340, 101360, 101350, 
    _, _, _, _, _, _, _, _, 101320, 101340, 101350, 101350, 101330, 101330, 
    101330, 101300, _, _, 101280, 101290, 101280, 101300, 101310, 101300, 
    101310, 101310, _, _, _, _, _, _, 101190, 101180, 101140, 101140, 101110, 
    101080, 101040, 101000, _, _, _, _, _, 100730, 100700, 100640, 100580, 
    100510, 100440, 100360, _, _, _, _, 100010, 99970, 99930, 99880, 99840, 
    99810, 99790, 99770, 99760, _, _, _, _, _, _, 100030, 100070, 100140, 
    100190, 100300, 100410, 100430, 100480, _, _, _, _, 100760, 100780, 
    100820, 100860, 100860, 100880, 100880, 100910, _, 100970, 101040, 
    101040, 101050, 101070, 101080, 101070, 101070, _, _, 101020, 101000, 
    100970, 100950, 100920, 100880, 100820, 100730, _, _, 100560, 100510, 
    100450, 100430, 100380, 100340, 100270, 100190, _, 100010, 99940, 99870, 
    99860, 99840, 99790, 99790, 99760, _, _, _, _, _, _, 99800, 99810, _, 
    99860, 99880, _, 99920, 99950, 99960, 99970, 99970, 99960, 99920, 99910, 
    99920, 99910, 99900, _, _, _, _, _, _, _, _, 99910, 99900, 99900, 99900, 
    99880, 99870, 99870, 99860, _, 99780, 99790, 99750, 99760, 99780, 99810, 
    99840, 99850, _, _, _, _, 100170, 100240, 100330, 100430, 100470, 100550, 
    100660, 100730, _, 100890, 101020, 101070, 101130, 101180, 101210, 
    101220, 101230, _, _, _, 101080, 101040, 100980, 100890, 100790, 100680, 
    100580, 100460, _, _, _, 100070, 99950, 99860, 99770, 99650, 99480, 
    99340, 99150, 98950, _, _, _, 98410, 98370, 98370, 98310, 98320, 98340, 
    98340, 98380, _, 98470, 98560, 98610, 98760, 98900, 98980, 99140, 99270, 
    99360, 99430, 99480, 99580, 99630, 99730, 99790, _, _, _, 100150, 100240, 
    100330, 100440, 100550, 100710, 100830, 100950, _, 101160, 101300, 
    101440, 101540, 101590, 101670, 101690, 101720, 101730, 101750, _, _, _, 
    _, 101750, 101720, 101650, 101600, 101540, 101470, 101370, 101290, _, _, 
    _, 100990, 100920, 100850, 100770, 100670, 100610, 100500, 100480, _, _, 
    _, 100260, 100230, 100160, 100150, 100100, 100040, 99970, 99910, 99860, 
    _, _, _, 99590, 99560, 99500, 99440, 99370, 99390, 99430, 99430, _, _, _, 
    99410, 99390, 99380, 99340, 99320, 99280, 99250, 99220, _, _, _, 99210, 
    99280, 99320, 99360, 99370, 99350, 99380, 99460, _, _, _, _, _, _, _, _, 
    99370, 99350, 99310, 99280, 99270, 99260, 99240, 99240, _, _, 99280, 
    99320, 99350, 99400, 99430, 99480, 99530, 99590, _, _, _, _, _, _, _, _, 
    _, _, 100240, 100310, 100350, _, _, _, 100600, 100620, 100590, _, 100660, 
    _, _, 100750, _, 100790, _, _, _, 100860, 100870, 100880, 100880, _, _, 
    100920, _, _, 101000, 101050, _, 101200, 101280, _, _, _, _, _, _, _, _, 
    _, 101870, _, _, _, _, _, _, _, 102170, 102170, 102190, 102200, 102210, 
    102270, _, _, _, _, _, 102340, 102340, _, 102280, 102270, 102230, 102210, 
    102220, _, _, 102130, 102120, 102100, _, 102030, 102030, 102000, 102020, 
    _, _, 102030, 102020, 102020, 102020, 102010, 102020, 102000, _, 101930, 
    101920, 101920, 101920, 101840, 101850, 101770, 101710, _, 101700, _, 
    101580, 101580, 101570, 101550, 101550, 101540, 101520, 101470, 101420, 
    101400, 101370, 101360, 101340, 101340, _, _, 101310, 101300, _, _, 
    101280, 101240, 101210, 101200, _, _, 101130, 101130, 101110, 101070, 
    101030, 100970, 100920, 100840, 100780, _, _, _, 100450, 100390, 100330, 
    _, _, _, 99950, 99800, 99670, 99560, 99500, 99440, 99390, _, 99240, 
    99160, 99060, 98960, 98840, 98790, 98690, 98720, _, _, _, 98480, 98460, 
    98410, _, 98320, 98340, 98310, 98310, 98280, 98250, 98270, _, 98330, _, 
    98360, _, _, _, _, _, 98580, 98610, _, 98670, _, 98750, _, 98830, 98810, 
    _, 98920, 98940, 98980, 99010, _, _, _, _, _, _, 99180, _, 99200, _, 
    99240, _, 99340, _, _, _, 99570, 99630, 99630, 99710, 99760, 99810, 
    99920, 99980, _, 100070, 100100, 100140, _, 100310, 100360, 100390, 
    100460, _, _, 100610, 100630, 100660, 100700, 100740, 100780, 100830, _, 
    100910, _, _, _, 101050, 101100, 101130, 101170, 101180, 101200, 101230, 
    101210, _, _, 101210, _, _, 101160, 101230, 101290, _, 101330, _, _, _, 
    _, _, _, _, _, 101540, 101600, 101630, 101610, 101590, 101620, 101630, _, 
    101630, 101620, 101610, 101590, 101550, 101510, 101510, _, _, _, _, 
    101150, 101030, _, 100840, 100760, _, 100590, 100480, 100380, 100290, _, 
    100110, _, 100070, 100060, 100050, 100080, _, _, 100070, 100070, 100090, 
    _, _, _, 100410, 100540, 100650, 100760, 100850, 100990, 101160, 101320, 
    _, 101540, _, 101740, _, _, 102040, _, _, _, 102440, 102500, 102500, 
    102500, 102530, 102540, 102510, 102520, 102410, _, 102300, _, 102250, _, 
    102140, 102060, 101980, 101950, _, _, _, 101680, 101680, 101730, 101710, 
    101690, 101730, 101710, 101730, _, _, _, _, _, _, _, _, _, _, 101890, 
    101870, 101820, 101780, 101700, 101620, 101440, 101240, _, _, 100930, _, 
    100980, 101090, _, 101350, 101480, _, _, _, _, 101930, _, 102010, 102020, 
    102070, 102130, _, _, 102140, _, _, 102090, _, 102140, 102070, 102090, 
    102060, 102040, 102000, _, _, _, 102150, _, _, _, 102410, 102500, 102570, 
    102670, 102820, 102900, 102980, 103060, 103090, _, _, _, _, 103440, 
    103460, 103490, 103500, 103500, 103530, 103530, 103560, _, 103600, 
    103580, 103570, 103540, 103530, 103510, 103490, 103490, 103490, 103470, 
    103460, 103430, 103410, 103380, 103360, 103330, 103290, _, _, _, _, 
    103100, 103050, _, 102940, 102870, 102820, 102740, 102690, 102630, 
    102590, 102510, _, _, _, _, 102240, 102190, 102100, 102050, 101980, 
    101930, 101860, 101820, _, _, 101730, 101710, 101710, 101720, 101740, 
    101760, 101810, 101830, _, _, 101860, 101890, 101880, 101870, 101840, 
    101800, 101780, 101750, _, _, 101580, 101500, 101470, 101460, 101450, 
    101450, 101450, 101470, _, _, 101450, 101450, 101470, 101480, 101490, 
    101480, 101510, 101530, 101530, 101530, 101530, 101520, 101500, 101480, 
    101490, 101470, 101460, 101470, _, _, _, _, 101550, 101550, 101540, 
    101530, 101500, 101500, _, _, 101520, 101540, 101530, 101500, 101500, 
    101510, 101500, 101510, _, _, 101530, 101520, 101540, 101560, 101550, 
    101530, _, 101540, 101510, _, _, 101580, 101560, 101540, 101610, 101630, 
    101650, 101680, 101690, _, _, _, _, 101730, 101760, 101770, 101810, 
    101840, 101850, 101930, 101940, _, _, _, 101940, 101930, 101930, 101960, 
    101990, 102040, 102030, 102030, 102050, _, _, 102060, 102050, 102040, 
    101970, 101950, 101940, 101870, 101870, _, 101820, 101810, 101820, 
    101830, 101830, 101780, 101740, 101740, _, _, _, _, _, 101810, 101790, 
    101780, 101790, 101780, 101770, 101790, 101810, _, _, 101840, 101840, _, 
    101840, 101840, 101840, 101860, 101860, _, _, _, 101920, 101910, 101900, 
    101860, 101840, 101780, 101650, 101540, _, _, 101140, 100820, 100640, 
    100460, 100380, 100400, 100430, 100670, 100910, _, _, 101290, 101360, 
    101410, 101460, 101480, 101520, 101560, 101570, _, _, _, _, 101670, 
    101690, 101710, 101750, 101780, 101780, 101800, 101840, _, _, _, _, _, _, 
    _, _, _, 101910, 101890, 101860, 101830, 101800, 101800, 101790, 101730, 
    101730, 101730, 101730, 101720, 101690, 101700, 101700, 101690, _, _, _, 
    _, _, _, 101720, 101710, 101720, 101700, 101680, 101650, 101650, 101650, 
    _, _, 101650, 101670, 101690, 101690, 101720, 101720, 101710, 101740, _, 
    _, 101720, 101720, 101710, 101720, 101730, 101750, 101760, 101780, 
    101770, 101770, 101800, 101820, 101820, 101840, 101890, _, 101960, 
    101990, 102020, 102040, 102040, 102040, _, _, _, _, _, _, 102070, 102050, 
    102010, 101980, 101940, 101890, 101840, 101810, _, _, _, _, _, 101740, 
    101690, 101680, 101630, 101560, 101550, 101540, 101500, _, _, _, _, _, _, 
    _, _, _, 101240, 101220, 101190, 101180, 101160, 101160, 101160, 101200, 
    _, _, _, 101260, 101270, 101300, 101310, 101340, 101360, 101350, 101370, 
    _, _, _, _, 101180, 101130, 101070, 101040, 101010, 101040, 101030, 
    101020, _, _, 101020, 101030, 101060, 101040, 101080, 101150, 101150, 
    101160, _, _, _, _, 101060, 101030, 101020, 101000, 100980, 101000, 
    101010, _, _, _, 101070, 101110, 101110, 101100, 101130, 101170, 101170, 
    101220, _, _, _, 101340, 101360, 101350, 101320, 101280, 101260, 101220, 
    101170, _, _, 101080, 101060, 101050, 101000, 100950, 100890, 100840, 
    100790, _, _, _, 100620, 100560, 100500, 100420, 100390, 100350, 100300, 
    100290, _, _, _, _, 100250, 100260, 100340, 100360, 100370, 100350, 
    100280, 100320, _, _, _, _, _, 100550, 100600, 100630, 100690, _, 100750, 
    100770, 100800, 100820, 100870, 100940, 101020, 101080, 101140, 101180, 
    _, 101250, 101270, 101310, 101330, 101350, 101370, 101380, _, _, _, _, _, 
    _, _, _, 101470, 101460, 101460, 101480, 101470, 101480, 101500, 101500, 
    101500, 101480, 101480, 101470, 101450, 101430, 101440, 101430, 101430, 
    101440, 101430, 101420, 101430, 101430, 101410, 101410, 101400, 101400, 
    101410, 101450, 101470, 101500, 101550, 101580, 101620, 101630, 101640, 
    101660, 101670, 101690, 101700, 101720, 101730, 101760, 101770, 101780, 
    101780, 101790, 101810, 101830, 101830, 101810, 101800, 101810, 101820, 
    101810, 101800, 101800, 101780, 101740, 101700, 101670, 101620, 101590, 
    101540, 101490, 101440, 101480, 101480, 101490, 101490, 101500, 101440, 
    101420, 101480, 101470, 101450, 101450, 101460, 101410, 101440, 101460, 
    101380, 101430, 101430, 101420, 101390, 101370, 101310, 101290, 101250, 
    101180, 101170, 101130, 101070, 101010, 100980, 100890, 100870, 100830, 
    100790, 100740, 100700, 100660, 100610, 100550, 100530, 100540, 100470, 
    100420, 100370, 100360, 100320, 100290, 100210, 100260, 100270, 100240, 
    100170, 100140, 100100, 100060, 100010, 99980, 99980, 99950, 99950, 
    99930, 99980, 100010, 99980, 100010, 99990, 100050, 100050, 100060, 
    100100, 100160, 100330, 100360, 100370, 100420, 100400, 100410, 100510, 
    100420, 100470, 100530, 100560, 100550, 100510, 100560, 100580, 100600, 
    100610, 100590, 100610, 100570, 100540, 100520, 100480, 100480, 100440, 
    100420, 100350, 100310, 100270, 100190, 100150, 100110, 100040, 100010, 
    99960, 99930, 99900, 99870, 99870, 99910, 99910, 99910, 99920, 99900, 
    99910, 99930, 99960, 100020, 100100, 100190, 100320, 100380, 100470, 
    100550, 100620, 100650, 100730, 100740, 100810, 100850, 100910, 100960, 
    101020, 101070, 101080, 101070, 101110, 101150, 101180, 101170, 101180, 
    101220, 101240, 101270, 101290, 101310, 101300, 101300, 101320, 101320, 
    101270, 101320, 101290, 101250, 101270, 101250, 101240, 101230, 101210, 
    101130, 101090, 101070, 100980, 100920, 100820, 100680, 100600, 100500, 
    100350, 100180, 99880, 99680, 99590, 99600, 99410, 99310, 99060, 98860, 
    98790, 98730, 98640, 98450, 98410, 98410, 98380, 98450, 98440, 98400, 
    98340, 98470, 98660, 98770, 98910, 98970, 99010, 99060, 99190, 99260, 
    99330, 99410, 99480, 99630, 99720, 99800, 99840, 99880, 100100, 100090, 
    99980, 100110, 100160, 100230, 100270, 100290, 100290, 100270, 100250, 
    100230, 100250, 100280, 100200, 100230, 100270, 100280, 100280, 100310, 
    100340, 100380, 100400, 100440, 100480, 100480, 100510, 100560, 100560, 
    100570, 100580, 100620, 100620, 100660, 100700, 100750, 100740, 100750, 
    100770, 100750, 100760, 100820, 100850, 100850, 100930, 101000, 101110, 
    101170, 101230, 101250, 101280, 101270, 101310, 101370, 101400, 101410, 
    101470, 101490, 101500, 101520, 101570, 101620, 101650, 101660, 101700, 
    101740, 101770, 101790, 101840, 101920, 101970, 102000, 102000, 102030, 
    101980, 101940, 102060, 102090, 102050, 102030, 102100, 102110, 102110, 
    102120, 102180, 102170, 102210, 102280, 102310, 102300, 102250, 102200, 
    102220, 102240, 102280, 102300, 102280, 102280, 102310, 102410, 102400, 
    102390, 102350, 102320, 102330, 102450, 102510, 102570, 102600, 102600, 
    102620, 102660, 102670, 102670, 102630, 102640, 102680, 102670, 102660, 
    102650, 102710, 102800, 102720, 102680, 102650, 102600, 102630, 102580, 
    102550, 102500, 102440, 102350, 102240, 102150, 102010, 101890, 101700, 
    101520, 101330, 101170, 100960, 100850, 100690, 100520, 100350, 100270, 
    100180, 100150, 100230, 100170, 100180, 100190, 100180, 100150, 100160, 
    100140, 100170, 100190, 100190, 100160, 100240, 100330, 100470, 100570, 
    100700, 100890, 101030, 101060, 101060, 101050, 101040, 100990, 101030, 
    101010, 100990, 101030, 101060, 101060, 101090, 101160, 101180, 101250, 
    101230, 101200, 101160, 101150, 101050, 100980, 100930, 100860, 100770, 
    100730, 100620, 100590, 100500, 100410, 100410, 100350, 100350, 100290, 
    100290, 100220, 100230, 100210, 100150, 100150, 100250, 100270, 100210, 
    100160, 100200, 100170, 100150, 100200, 100190, 100160, 100150, 100200, 
    100230, 100250, 100230, 100250, 100230, 100260, 100340, 100490, 100510, 
    100610, 100650, 100710, 100730, 100730, 100770, 100790, 100830, 100830, 
    100880, 100910, 100940, 100970, 101010, 101070, 101140, 101210, 101280, 
    101350, 101410, 101400, 101490, 101560, 101630, 101690, 101700, 101760, 
    101700, 101710, 101730, 101760, 101800, 101860, 101890, 101950, 102020, 
    102050, 102110, 102090, 102140, 102080, 102210, 102180, 102180, 102150, 
    102120, 102120, 102130, 102130, 102110, 102100, 102010, 101940, 101830, 
    101830, 101740, 101680, 101630, 101620, 101560, 101600, 101570, 101620, 
    101560, 101550, 101590, 101540, 101620, 101620, 101650, 101700, 101670, 
    101640, 101620, 101650, 101630, 101600, 101510, 101400, 101400, 101290, 
    101110, 101080, 101090, 101040, 100950, 100920, 100870, 100850, 100810, 
    100800, 100760, 100770, 100750, 100750, 100770, 100770, 100770, 100730, 
    100660, 100640, 100620, 100650, 100610, 100560, 100590, 100570, 100530, 
    100480, 100420, 100380, 100300, 100190, 100070, 99960, 99840, 99720, 
    99620, 99550, 99430, 99390, 99480, 99470, 99610, 99780, 99960, 100070, 
    100170, 100250, 100320, 100350, 100360, 100390, 100430, 100450, 100450, 
    100530, 100530, 100530, 100610, 100630, 100690, 100730, 100750, 100850, 
    100880, 100920, 100930, 100940, 101010, 101070, 101120, 101130, 101140, 
    101160, 101230, 101310, 101320, 101340, 101330, 101320, 101310, 101310, 
    101350, 101330, 101370, 101360, 101360, 101420, 101410, 101380, 101420, 
    101410, 101370, 101340, 101320, 101290, 101310, 101320, 101280, 101280, 
    101240, 101190, 101130, 101100, 100990, 100950, 100880, 100740, 100580, 
    100490, 100440, 100370, 100330, 100220, 100180, 100130, 100070, 99990, 
    99960, 99940, 99870, 99850, 99800, 99740, 99710, 99660, 99600, 99590, 
    99520, 99480, 99500, 99490, 99490, 99480, 99520, 99570, 99620, 99660, 
    99690, 99720, 99730, 99720, 99720, 99710, 99710, 99710, 99740, 99710, 
    99730, 99770, 99740, 99770, 99830, 99920, 100050, 100200, 100340, 100530, 
    100700, 100870, 101000, 101120, 101270, 101400, 101550, 101680, 101790, 
    101890, 101970, 102060, 102130, 102340, 102420, 102480, 102590, 102700, 
    102840, 102900, 102920, 102970, 103030, 103080, 103140, 103170, 103190, 
    103220, 103240, 103290, 103330, 103330, 103330, 103370, 103410, 103400, 
    103400, 103390, 103380, 103350, 103310, 103290, 103290, 103280, 103220, 
    103200, 103160, 103170, 103100, 103040, 103000, 102980, 102940, 102910, 
    102900, 102890, 102880, 102910, 102910, 102940, 102960, 102980, 103000, 
    103020, 103030, 103040, 103060, 103060, 103110, 103110, 103160, 103160, 
    103140, 103210, 103190, 103200, 103150, 103130, 102970, 103020, 103110, 
    103160, 103150, 103140, 103060, 103000, 102900, 102800, 102740, 102720, 
    102710, 102590, 102420, 102260, 102300, 102280, 102470, 102280, 102320, 
    102250, 102260, 102190, 102170, 102080, 101970, 101770, 101810, 101870, 
    101770, 101860, 101840, 101820, 101930, 101940, 101850, 101900, 101930, 
    101920, 101940, 102010, 102060, 102090, 102130, 102150, 102140, 102160, 
    102150, 102100, 102060, 102000, 102000, 101940, 101870, 101840, 101780, 
    101720, 101650, 101630, 101620, 101560, 101510, 101500, 101470, 101490, 
    101460, 101450, 101410, 101320, 101300, 101280, 101290, 101270, 101270, 
    101250, 101240, 101190, 101170, 101150, 101100, 101020, 100950, 100910, 
    100820, 100740, 100700, 100580, 100500, 100420, 100260, 100100, 100140, 
    100020, 99920, 99710, 99560, 99370, 99250, 99160, 99000, 98860, 98700, 
    98480, 98420, 98050, 98180, 98060, 97900, 97770, 97470, 97370, 97340, 
    97290, 97330, 97210, 97100, 97260, 97390, 97430, 97470, 97520, 97580, 
    97630, 97700, 97710, 97770, 97810, 97850, 97770, 97870, 98260, 98400, 
    98400, 98420, 98460, 98530, 98510, 98560, 98660, 98700, 98750, 98790, 
    98810, 98800, 98840, 98900, 98850, 98910, 99000, 98940, 98990, 98960, 
    98930, 98890, 98800, 98750, 98630, 98520, 98510, 98380, 98370, 98320, 
    98280, 98260, 98220, 98190, 98220, 98230, 98300, 98400, 98510, 98580, 
    98600, 98640, 98620, 98670, 98720, 98750, 98770, 98840, 98890, 98910, 
    98950, 98970, 99010, 99050, 99070, 99100, 99110, 99130, 99150, 99180, 
    99220, 99230, 99260, 99270, 99300, 99350, 99390, 99430, 99470, 99480, 
    99500, 99520, 99560, 99590, 99610, 99640, 99660, 99710, 99720, 99730, 
    99720, 99720, 99730, 99690, 99680, 99630, 99570, 99520, 99450, 99350, 
    99300, 99170, 99080, 98990, 98870, 98680, 98490, 98290, 98120, 97970, 
    97850, 97740, 97680, 97540, 97450, 97450, 97390, 97330, 97250, 97240, 
    97210, 97160, 97160, 97150, 97170, 97180, 97190, 97210, 97260, 97270, 
    97300, 97370, 97430, 97510, 97580, 97640, 97680, 97760, 97800, 97830, 
    97860, 97890, 97930, 97950, 98020, 98030, 98050, 98100, 98130, 98130, 
    98200, 98200, 98180, 98190, 98180, 98260, 98320, 98400, 98420, 98500, 
    98550, 98580, 98640, 98640, 98670, 98690, 98710, 98760, 98800, 98870, 
    98910, 98960, 98960, 99000, 99070, 99080, 99130, 99170, 99210, 99210, 
    99200, 99180, 99190, 99060, 99080, 99090, 99100, 99110, 99090, 99100, 
    99110, 99080, 99110, 99070, 99110, 99120, 99120, 99100, 99090, 99060, 
    99010, 98950, 98930, 98900, 98900, 98890, 98920, 98880, 98840, 98810, 
    98700, 98640, 98580, 98490, 98440, 98380, 98320, 98310, 98330, 98320, 
    98270, 98270, 98260, 98220, 98160, 98140, 98160, 98130, 98090, 98050, 
    97990, 98010, 98030, 98050, 98090, 98080, 98080, 98100, 98110, 98150, 
    98190, 98250, 98300, 98350, 98390, 98360, 98320, 98280, 98280, 98360, 
    98440, 98500, 98560, 98640, 98730, 98840, 98890, 98950, 98970, 99010, 
    99070, 99080, 99180, 99200, 99230, 99270, 99300, 99330, 99340, 99340, 
    99330, 99310, 99310, 99250, 99240, 99210, 99210, 99220, 99240, 99220, 
    99230, 99210, 99230, 99240, 99260, 99260, 99270, 99300, 99310, 99310, 
    99300, 99300, 99340, 99320, 99310, 99300, 99290, 99300, 99300, 99280, 
    99300, 99300, 99340, 99340, 99380, 99340, 99390, 99430, 99460, 99510, 
    99540, 99550, 99550, 99640, 99670, 99770, 99790, 99820, 99830, 99870, 
    99930, 99960, 99990, 100060, 100040, 100090, 100120, 100170, 100210, 
    100210, 100220, 100210, 100210, 100250, 100280, 100340, 100370, 100380, 
    100390, 100390, 100390, 100390, 100410, 100440, 100470, 100480, 100500, 
    100480, 100550, 100530, 100540, 100590, 100590, 100530, 100520, 100540, 
    100530, 100510, 100490, 100440, 100410, 100380, 100420, 100450, 100490, 
    100460, 100390, 100420, 100440, 100500, 100470, 100450, 100460, 100440, 
    100440, 100480, 100470, 100460, 100450, 100440, 100430, 100460, 100530, 
    100550, 100580, 100580, 100590, 100670, 100700, 100720, 100730, 100720, 
    100700, 100730, 100750, 100740, 100760, 100780, 100790, 100790, 100840, 
    100840, 100830, 100840, 100820, 100850, 100850, 100880, 100920, 100920, 
    100900, 100900, 100940, 100930, 100940, 100990, 100980, 101000, 101020, 
    101030, 101040, 101070, 101130, 101110, 101160, 101160, 101210, 101190, 
    101250, 101260, 101300, 101300, 101300, 101350, 101380, 101440, 101490, 
    101500, 101490, 101480, 101460, 101500, 101500, 101500, 101500, 101520, 
    101510, 101520, 101520, 101450, 101510, 101490, 101470, 101520, 101550, 
    101560, 101620, 101650, 101720, 101770, 101800, 101870, 101870, 101860, 
    101880, 101860, 101890, 101900, 101890, 101910, 101950, 101980, 101990, 
    101960, 101950, 101940, 101950, 101950, 101960, 101940, 101930, 101940, 
    101970, 101990, 102010, 102020, 101980, 101940, 101930, 101910, 101860, 
    101880, 101870, 101850, 101850, 101880, 101910, 101890, 101920, 101920, 
    101910, 101860, 101850, 101880, 101830, 101840, 101850, 101860, 101840, 
    101820, 101790, 101760, 101730, 101710, 101690, 101670, 101600, 101500, 
    101480, 101480, 101480, 101460, 101360, 101310, 101220, 101180, 101160, 
    101100, 101090, 101070, 101110, 101100, 100930, 101050, 100930, 100690, 
    100600, 100560, 100500, 100510, 100470, 100490, 100420, 100360, 100260, 
    100250, 100300, 100300, 100290, 100270, 100100, 100010, 99830, 99700, 
    99640, 99530, 99530, 99500, 99410, 99280, 99160, 98990, 98900, 98870, 
    98810, 98760, 98770, 98750, 98740, 98730, 98700, 98590, 98450, 98430, 
    98510, 98500, 98550, 98620, 98740, 98810, 98730, 98840, 98900, 98910, 
    98950, 99000, 99060, 99140, 99120, 99160, 99180, 99140, 99130, 99160, 
    99150, 99130, 99110, 99160, 99150, 99120, 99130, 99150, 99190, 99200, 
    99170, 99150, 99140, 99060, 98980, 98940, 98890, 98870, 98860, 98830, 
    98790, 98790, 98740, 98710, 98680, 98670, 98620, 98590, 98600, 98610, 
    98610, 98580, 98590, 98640, 98750, 98820, 98830, 98850, 98880, 98930, 
    98950, 98990, 99020, 99100, 99130, 99160, 99130, 99190, 99240, 99350, 
    99470, 99570, 99640, 99750, 99790, 99910, 100050, 100150, 100250, 100350, 
    100420, 100490, 100550, 100600, 100650, 100740, 100790, 100860, 100920, 
    100990, 101080, 101120, 101200, 101250, 101310, 101360, 101370, 101400, 
    101420, 101470, 101520, 101580, 101600, 101670, 101700, 101730, 101750, 
    101760, 101780, 101790, 101810, 101840, 101860, 101850, 101870, 101890, 
    101870, 101840, 101850, 101830, 101820, 101770, 101760, 101750, 101750, 
    101770, 101750, 101750, 101730, 101730, 101750, 101740, 101760, 101750, 
    101730, 101740, 101720, 101690, 101700, 101690, 101650, 101600, 101580, 
    101540, 101500, 101430, 101410, 101380, 101330, 101300, 101260, 101210, 
    101190, 101140, 101050, 101000, 100960, 100900, 100820, 100780, 100760, 
    100700, 100620, 100570, 100540, 100480, 100410, 100340, 100320, 100290, 
    100270, 100270, 100280, 100260, 100250, 100230, 100200, 100160, 100100, 
    100060, 100040, 99980, 99950, 99930, 99820, 99750, 99710, 99640, 99590, 
    99540, 99460, 99420, 99400, 99460, 99520, 99630, 99730, 99810, 99880, 
    99940, 100000, 100060, 100060, 100080, 100100, 100160, 100200, 100240, 
    100300, 100330, 100360, 100390, 100400, 100420, 100460, 100460, 100500, 
    100530, 100540, 100550, 100560, 100570, 100570, 100620, 100630, 100640, 
    100640, 100670, 100660, 100710, 100730, 100730, 100760, 100740, 100750, 
    100750, 100750, 100740, 100710, 100680, 100670, 100640, 100630, 100620, 
    100630, 100620, 100620, 100600, 100590, 100610, 100640, 100670, 100690, 
    100700, 100740, 100800, 100860, 100910, 100990, 101040, 101070, 101070, 
    101160, 101160, 101150, 101160, 101130, 101180, 101220, 101260, 101270, 
    101320, 101280, 101290, 101280, 101270, 101270, 101270, 101270, 101250, 
    101250, 101230, 101210, 101200, 101170, 101130, 101090, 101060, 101010, 
    100970, 100940, 100910, 100920, 100900, 100840, 100800, 100750, 100670, 
    100600, 100550, 100550, 100510, 100520, 100510, 100520, 100550, 100590, 
    100530, 100610, 100560, 100590, 100630, 100630, 100630, 100670, 100720, 
    100750, 100860, 100780, 100870, 100890, 100870, 100860, 100860, 100900, 
    100910, 100910, 100940, 100990, 101000, 100980, 100990, 100980, 101000, 
    101010, 100930, 100900, 100940, 100980, 101000, 101030, 101000, 101020, 
    101040, 101020, 101010, 101010, 101000, 101020, 101020, 101020, 101030, 
    101030, 101010, 101000, 100980, 100980, 100970, 100950, 100930, 100950, 
    100920, 100920, 100940, 100940, 100990, 101010, 101030, 101060, 101090, 
    101080, 101090, 101080, 101090, 101120, 101130, 101170, 101170, 101200, 
    101240, 101250, 101260, 101280, 101270, 101300, 101310, 101300, 101340, 
    101380, 101380, 101390, 101370, 101370, 101370, 101390, 101420, 101380, 
    101400, 101390, 101370, 101380, 101450, 101440, 101410, 101410, 101450, 
    101420, 101390, 101360, 101340, 101370, 101390, 101430, 101420, 101460, 
    101470, 101460, 101500, 101530, 101530, 101550, 101560, 101560, 101560, 
    101590, 101610, 101600, 101560, 101530, 101480, 101440, 101400, 101290, 
    101290, 101250, 101180, 101150, 101130, 101080, 101050, 100980, 100910, 
    100880, 100850, 100820, 100790, 100770, 100780, 100820, 100910, 101020, 
    101090, 101160, 101250, 101230, 101350, 101360, 101270, 101330, 101260, 
    101140, 101160, 101040, 100950, 100830, 100680, 100540, 100430, 100360, 
    100270, 100120, 100080, 100060, 100070, 100070, 100020, 100130, 100070, 
    100120, 100220, 100230, 100260, 100330, 100470, 100530, 100600, 100760, 
    100850, 100930, 101060, 101160, 101270, 101420, 101470, 101560, 101770, 
    101920, 102000, 102050, 102120, 102200, 102260, 102350, 102300, 102360, 
    102380, 102370, 102400, 102370, 102400, 102360, 102330, 102220, 102150, 
    102100, 102050, 101960, 101890, 101820, 101720, 101610, 101550, 101420, 
    101300, 101140, 100930, 100770, 100530, 100430, 100300, 100240, 100200, 
    100170, 100140, 100060, 100040, 100030, 99980, 100010, 100030, 100050, 
    100010, 100030, 100020, 100040, 100040, 100040, 100020, 99970, 99960, 
    99930, 99920, 99920, 99930, 99950, 99970, 100020, 100080, 100120, 100160, 
    100200, 100230, 100250, 100280, 100260, 100280, 100320, 100330, 100400, 
    100410, 100470, 100480, 100520, 100530, 100550, 100560, 100580, 100600, 
    100610, 100640, 100670, 100710, 100760, 100800, 100820, 100840, 100890, 
    100940, 101010, 101020, 101060, 101090, 101140, 101170, 101220, 101270, 
    101310, 101330, 101360, 101390, 101420, 101460, 101480, 101520, 101550, 
    101600, 101630, 101650, 101650, 101680, 101700, 101590, 101670, 101700, 
    101660, 101610, 101640, 101610, 101620, 101640, 101650, 101630, 101630, 
    101600, 101640, 101590, 101620, 101640, 101690, 101650, 101700, 101740, 
    101710, 101680, 101670, 101730, 101860, 101880, 101890, 101880, 101910, 
    101930, 101940, 101910, 101870, 101870, 101900, 101900, 101890, 101840, 
    101830, 101800, 101760, 101750, 101760, 101720, 101670, 101660, 101650, 
    101690, 101690, 101690, 101660, 101690, 101690, 101680, 101740, 101720, 
    101740, 101750, 101780, 101750, 101730, 101740, 101730, 101680, 101690, 
    101680, 101640, 101540, 101550, 101530, 101470, 101430, 101410, 101370, 
    101370, 101420, 101450, 101480, 101520, 101520, 101550, 101590, 101620, 
    101630, 101690, 101720, 101720, 101750, 101800, 101850, 101900, 101950, 
    101980, 101970, 101980, 102000, 102050, 102060, 102070, 102070, 102100, 
    102120, 102140, 102160, 102140, 102150, 102160, 102190, 102200, 102180, 
    102200, 102210, 102230, 102260, 102270, 102280, 102250, 102240, 102240, 
    102210, 102210, 102230, 102210, 102210, 102220, 102250, 102270, 102270, 
    102290, 102270, 102270, 102310, 102320, 102320, 102330, 102360, 102380, 
    102430, 102470, 102510, 102530, 102550, 102560, 102580, 102600, 102650, 
    102690, 102700, 102730, 102790, 102820, 102830, 102840, 102810, 102820, 
    102830, 102840, 102850, 102820, 102830, 102850, 102910, 102920, 102900, 
    102950, 102910, 102930, 102930, 102930, 102920, 102910, 102950, 102930, 
    102880, 102930, 102930, 102970, 102870, 102850, 102910, 102850, 102860, 
    102840, 102810, 102870, 103000, 103010, 103020, 103020, 102990, 102980, 
    103020, 103030, 103040, 103030, 102930, 102930, 102960, 102960, 102930, 
    102880, 102830, 102820, 102770, 102730, _, 102700, _, _, 102620, 102560, 
    102490, 102490, 102330, 102180, 102050, 101990, 101900, 101770, 101680, 
    101630, 101600, 101580, 101490, 101390, 101330, 101280, 101270, 101260, 
    101230, 101190, 101180, 101180, 101150, 101120, 101050, 100980, 100820, 
    100680, 100530, 100320, 100130, 99950, 99770, 99650, 99530, 99410, 99290, 
    99210, 99090, 98980, 98850, 98690, 98550, 98390, 98270, 98100, 97950, 
    97870, 97790, 97700, 97630, 97550, 97460, 97400, 97460, 97470, 97530, 
    97620, 97710, 97790, 97840, 97880, 97910, 98040, 98090, 98120, 98120, 
    98100, 98120, 98130, 98160, 98180, 98190, 98200, 98210, 98190, _, 98150, 
    98130, _, _, 97960, _, 97910, 97850, 97760, _, 97670, _, 97550, 97480, 
    97450, 97410, 97390, _, 97410, 97400, 97420, 97420, 97460, 97500, 97530, 
    97600, 97690, 97800, 97920, 97960, _, 98140, _, 98200, 98240, 98280, 
    98350, 98380, 98400, 98420, 98430, 98440, 98410, 98420, 98410, 98400, 
    98400, 98400, 98430, 98430, 98450, 98450, 98460, 98490, 98470, 98490, 
    98480, 98450, 98440, 98420, 98400, 98380, 98350, 98350, 98320, 98310, 
    98300, 98250, 98200, 98170, 98110, 98100, 98050, 97960, 97930, 97900, 
    97860, 97830, 97830, 97820, 97810, 97810, 97820, 97810, 97810, 97830, 
    97870, 97920, 97980, 98030, 98060, 98080, 98110, 98160, 98190, 98220, 
    98260, 98260, 98280, 98320, 98380, 98430, 98480, 98510, 98540, 98560, 
    98590, 98630, 98640, 98680, 98720, 98750, 98790, 98830, 98860, 98880, 
    98880, 98890, 98920, 98920, 98910, 98920, 98870, 98880, 98880, 98900, 
    98900, 98900, 98860, 98820, 98800, 98800, 98800, 98810, 98780, 98810, 
    98810, 98800, 98830, 98810, 98770, 98770, 98740, 98750, 98830, 98830, 
    98830, 98840, 98850, 98870, 98870, 98850, 98870, 98860, 98850, 98880, 
    98900, 98950, 98980, 99020, 99050, 99080, 99140, 99180, 99220, 99290, 
    99350, 99420, 99490, 99520, 99540, 99590, 99670, 99700, 99770, 99840, 
    99880, 99930, 99990, 100040, 100090, 100120, 100160, 100220, 100300, 
    100340, 100410, 100460, 100490, 100510, 100590, 100640, 100670, 100720, 
    100760, 100810, 100840, 100890, 100950, 101010, 101110, 101200, 101340, 
    101430, 101510, 101620, 101620, 101710, 101820, 101860, 101830, 101800, 
    101730, 101630, 101490, 101380, 101160, 100990, 100740, 100460, 100210, 
    99920, 99690, 99480, 99150, 99000, 98710, 98640, 98470, 98410, 98320, 
    98300, 98310, 98310, 98310, 98350, 98350, 98300, 98260, 98190, 98180, 
    98130, 98090, 98130, 98160, 98220, 98260, 98250, 98250, 98230, 98250, 
    98300, 98330, 98350, 98430, 98520, 98570, 98620, 98580, 98580, 98610, 
    98560, 98480, 98380, 98300, 98250, 98270, 98180, 98140, 98070, 98020, 
    98010, 97960, 97880, 97880, 97940, 98010, 98070, 98080, 98190, 98330, 
    98410, 98540, 98560, 98580, 98600, 98640, 98650, 98670, 98690, 98750, 
    98750, 98790, 98810, 98840, 98880, 98890, 98900, 98900, 98890, 98880, 
    98880, 98880, 98890, 98870, 98890, 98910, 98890, 98890, 98890, 98890, 
    98890, 98850, 98820, 98780, 98800, 98820, 98810, 98790, 98800, 98770, 
    98770, 98770, 98790, 98780, 98770, 98760, 98740, 98740, 98760, 98780, 
    98780, 98780, 98770, 98780, 98750, 98760, 98760, 98760, 98750, 98740, 
    98740, 98720, 98690, 98710, 98670, 98670, 98650, 98610, 98630, 98660, 
    98670, 98710, 98730, 98750, 98760, 98750, 98750, 98760, 98770, 98760, 
    98750, 98760, 98770, 98770, 98790, 98810, 98800, 98800, 98780, 98790, 
    98770, 98710, 98670, 98620, 98550, 98510, 98440, 98350, 98290, 98130, 
    98090, 98090, 98090, 98130, 98220, 98320, 98430, 98540, 98650, 98770, 
    98870, 98960, 99040, 99120, 99220, 99300, 99360, 99440, 99530, 99620, 
    99700, 99790, 99880, 99960, 100020, 100100, 100160, 100210, 100260, 
    100330, 100370, 100440, 100490, 100550, 100590, 100620, 100620, 100680, 
    100670, 100730, 100750, 100720, 100810, 100830, 100860, 100850, 100950, 
    100940, 100960, 100960, 100960, 101010, 101030, 101000, 100970, 100930, 
    100870, 100770, 100700, 100490, 100500, 100480, 100490, 100470, 100410, 
    100370, 100320, 100280, 100270, 100240, 100190, 100200, 100080, 100040, 
    100000, 99980, 99940, 99870, 99800, 99770, 99730, 99710, 99690, 99700, 
    99730, 99770, 99820, 99830, 99810, 99840, 99870, 99900, 99930, 99960, 
    100030, 100090, 100170, 100200, 100270, 100340, 100410, 100460, 100540, 
    100570, 100650, 100760, 100850, 100960, 100960, 100990, 101010, 101040, 
    101060, 101080, 101170, 101200, 101240, 101320, 101320, 101290, 101350, 
    101350, 101410, 101330, 101340, 101340, 101360, 101330, 101300, 101260, 
    101260, 101220, 101200, 101160, 101110, 101070, 101000, 100990, 100970, 
    100960, 100940, 100890, 100870, 100850, 100870, 100810, 100770, 100790, 
    100770, 100740, 100720, 100700, 100680, 100720, 100700, 100680, 100660, 
    100670, 100620, 100550, 100580, 100630, 100560, 100550, 100540, 100470, 
    100490, 100470, 100510, 100570, 100580, 100550, 100510, 100510, 100530, 
    100580, 100580, 100590, 100600, 100600, 100590, 100600, 100630, 100610, 
    100650, 100690, 100690, 100710, 100710, 100740, 100740, 100770, 100670, 
    100630, 100580, 100490, 100540, 100320, 100440, 100410, 100340, 100350, 
    100400, 100170, 100210, 100140, 100200, 100240, 100180, 100130, 100080, 
    100020, 100020, 100060, 100050, 100030, 99980, 100020, 100000, 100000, 
    99970, 99980, 100050, 100080, 100100, 100130, 100160, 100220, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 101890, 101880, 101840, 101760, 101640, 
    101500, 101320, 101110, 100850, 100500, 100240, 99940, 99700, 99510, 
    99250, 99070, 99130, 99110, 99090, 99000, 98980, 98870, 98710, 98480, 
    98220, 97920, 97540, 97320, 97210, 97280, 97530, 97710, 97890, 98030, 
    98200, 98340, 98550, 98620, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 101440, 101450, 101490, 
    101530, 101570, 101610, 101650, 101730, 101760, 101800, 101830, 101860, 
    101880, 101890, 101940, 101960, 101980, 102020, 102050, 102090, 102120, 
    102120, 102110, 102080, 102070, 102120, 102050, 102060, 102080, 102070, 
    102090, 102070, 102040, 102040, 102030, 102050, 102010, 101970, 101950, 
    101960, 101960, 102010, 102010, 102070, 102070, 102030, 102070, 102070, 
    102090, 102060, 102060, 102060, 102080, 102100, 102150, 102150, 102100, 
    102080, 102060, 102090, 102080, 102080, 102090, 102070, 102010, 102020, 
    102050, 102080, 102100, 102090, 102090, 102090, 102060, 102010, 101990, 
    102000, 102000, 102000, 102020, 102010, 102010, 102010, 101990, 101990, 
    101980, 102010, 102020, 101990, 101970, 101940, 101910, 101910, 101930, 
    101920, 101910, 101860, 101790, 101780, 101750, 101680, 101680, 101650, 
    101600, 101550, 101550, 101510, 101450, 101410, _, 101370, _, _, 101320, 
    101340, 101370, 101390, 101390, 101410, _, 101410, 101400, _, 101420, 
    101440, _, 101410, 101420, _, _, _, _, 101450, 101410, 101420, 101430, _, 
    101460, 101450, 101490, 101470, 101530, 101510, 101510, 101540, 101520, 
    101490, 101560, 101570, 101540, 101560, 101570, 101590, 101600, 101590, 
    101590, 101540, 101500, 101540, 101500, 101500, 101470, 101430, 101430, 
    101460, 101480, 101540, 101520, 101490, 101450, 101510, 101560, 101560, 
    101550, 101550, 101570, 101560, 101560, 101540, 101550, 101530, 101540, 
    101530, 101530, 101550, 101590, 101570, 101590, 101560, 101480, 101450, 
    101440, 101410, 101340, 101280, 101210, 101150, 101110, 101070, 101000, 
    100870, 100830, 100790, 100660, 100540, 100480, 100420, 100320, 100260, 
    100230, 100180, 100100, 100020, 99900, 99860, 99840, 99800, 99790, 99740, 
    99740, 99770, 99800, 99830, 99880, 99910, 99940, 99960, 99970, 99920, 
    99960, 99970, 99960, 99930, 99930, 99900, 99850, _, _, _, 99610, 99550, 
    99480, 99430, 99380, 99310, 99260, 99230, 99230, 99210, 99180, 99150, 
    99140, 99120, 99090, 99060, 99060, 99100, 99110, 99090, 99080, 99080, 
    99100, 99100, 99070, 99060, 99060, 99070, 99120, 99160, 99220, 99280, 
    99360, 99490, 99680, 99730, 99770, 99850, 99900, 100010, 100090, 100160, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 100620, 100470, 100480, 100510, 100310, 100280, 100120, 100060, _, 
    100040, 99900, 99940, 99870, 99720, _, _, 99690, 99690, 99670, 99720, 
    99740, 99790, 99800, 99810, _, 99920, 100020, 100040, 100080, _, 100150, 
    100220, 100240, 100290, 100330, 100390, 100390, 100370, 100350, 100400, 
    100420, 100420, 100430, 100450, 100410, 100310, 100300, 100340, 100350, 
    100310, 100290, 100190, 100200, 100180, 100130, 100050, 99970, 99900, 
    99870, 99810, 99770, 99750, 99770, 99730, 99760, 99750, 99760, 99770, 
    99790, 99860, 99920, 99970, 100040, 100100, 100150, 100230, 100300, 
    100390, 100500, 100600, 100660, 100780, 100890, 100980, 101100, 101220, 
    101240, 101320, 101400, 101530, 101600, 101690, 101740, 101820, 101880, 
    101940, _, 101930, 101950, 101990, 102040, 102060, 102100, 102100, 
    102090, 102160, 102250, 102260, 102330, 102360, 102380, 102420, 102460, 
    102480, 102510, 102550, 102550, 102570, 102620, 102680, 102700, 102720, 
    102770, 102800, 102840, 102840, 102870, 102900, 102940, 102960, 103000, 
    103010, 103010, 103030, 103050, 103040, 103060, 103050, 103050, 103080, 
    103050, 103050, 103030, 103010, 103000, 102970, 102960, 102940, 102930, 
    102940, 102890, 102790, 102720, 102730, 102660, 102520, 102430, 102240, 
    102250, 102150, 101980, 101880, 101800, 101780, 101720, 101610, 101550, 
    101420, 101300, 101150, 101030, 100950, 100810, 100720, 100640, 100550, 
    100460, 100390, 100320, 100240, 100140, 100100, 100010, 99920, 99880, _, 
    99840, 99800, 99740, 99610, 99570, 99560, 99480, 99300, 99250, 99140, 
    99090, 99060, 98970, 98890, 98800, 98780, 98730, 98720, 98740, 98740, 
    98760, 98760, 98760, 98760, 98810, 98850, 98880, 98930, 98940, 99020, 
    99080, 99140, 99190, 99250, 99320, 99360, 99440, 99490, 99520, 99550, 
    99600, 99640, 99680, 99720, 99770, 99790, 99800, 99810, 99840, 99850, 
    99880, 99870, 99840, 99830, 99840, 99850, 99830, 99830, 99820, 99750, 
    99680, 99620, 99590, 99550, 99580, 99560, 99540, 99490, 99450, 99450, 
    99490, 99460, 99450, 99460, 99470, 99460, 99440, 99470, 99510, 99560, 
    99580, 99590, 99590, 99600, 99610, 99610, 99620, 99630, 99640, 99660, 
    99650, 99690, 99720, 99720, 99730, 99750, 99750, 99760, 99800, 99870, 
    99900, 99950, 100000, 100030, 100050, 100080, 100120, 100140, 100130, 
    100150, 100170, 100180, 100200, 100230, 100250, 100270, 100280, 100300, 
    100300, 100310, 100330, 100350, 100390, 100430, 100480, 100480, 100510, 
    100550, 100560, 100550, 100550, 100570, 100570, 100580, 100610, 100620, 
    100630, 100620, 100600, 100630, 100630, 100610, 100570, 100590, 100610, 
    100600, 100610, 100620, 100600, 100610, 100600, 100560, 100540, 100480, 
    100440, 100420, 100390, 100370, 100340, 100280, 100250, 100220, 100190, 
    100160, 100120, 100030, 100010, 99990, 100000, 100000, 100050, 100080, 
    100090, 100120, 100170, 100210, 100230, 100270, 100320, 100380, 100420, 
    100470, 100530, 100580, 100610, 100650, 100690, 100730, 100770, 100780, 
    100790, 100800, 100820, 100920, 100940, 100950, 100970, 100950, 100830, 
    100810, 100770, 100770, 100750, 100690, 100640, 100590, 100530, 100450, 
    100380, 100300, 100250, 100140, 100050, 99960, 99820, 99750, 99740, 
    99730, 99740, 99790, 99940, 100100, 100240, 100320, 100440, 100530, 
    100630, 100660, 100740, 100820, 100900, 100920, 101020, 101050, 101010, 
    100980, 100930, 100810, 100730, 100630, 100530, 100470, 100330, 100210, 
    100080, 99990, 99850, 99760, 99650, 99560, 99470, 99410, 99370, 99320, 
    99290, 99270, 99290, 99290, 99320, 99340, 99370, 99440, 99520, 99610, 
    99680, 99830, 99930, 100010, 100100, 100100, 100180, 100270, 100340, 
    100400, 100480, 100550, 100580, 100640, 100660, 100690, 100730, 100760, 
    100740, 100730, 100710, 100730, 100730, 100730, 100760, 100760, 100770, 
    100800, 100830, 100850, 100880, 100920, 100950, 100970, 101000, 101050, 
    101140, 101190, 101230, 101240, 101280, 101320, 101340, 101360, 101360, 
    101380, 101400, 101420, 101460, 101450, 101470, 101420, 101400, 101380, 
    101340, 101280, 101270, 101230, 101190, 101000, 100990, 100980, 100970, 
    100930, 100890, 100870, 100850, 100830, 100780, 100770, 100730, 100710, 
    100650, 100660, 100660, 100660, 100620, 100510, 100500, 100570, 100530, 
    100500, 100440, 100290, 100280, 100110, 100200, 100320, 100420, 100670, 
    100860, 100940, 101250, 101240, 101690, 101780, 101870, 102010, 102030, 
    102090, 102050, 102230, 102250, 102270, 102260, 102260, 102300, 102320, 
    102250, 102320, 102370, 102360, 102400, 102380, 102340, 102390, 102420, 
    102360, 102170, 101970, 102190, 102000, 101910, 101800, 101700, 101620, 
    101510, 101460, 101430, 101400, 101320, 101300, 101310, 101300, 101290, 
    101240, 101310, 101330, 101460, 101440, 101460, 101470, 101480, 101490, 
    101590, 101590, 101590, 101600, 101530, 101560, 101650, 101580, 101620, 
    101610, 101620, 101630, 101570, 101610, 101600, 101600, 101580, 101620, 
    101600, 101620, 101600, 101600, 101610, 101580, 101460, 101530, 101510, 
    101510, 101520, 101490, 101510, 101510, 101540, 101600, 101610, 101650, 
    101650, 101670, 101700, 101720, 101750, 101760, 101810, 101830, 101860, 
    101880, 101880, 101910, 101940, 101930, 101950, 101920, 101920, 101920, 
    101930, 101940, 101950, 101960, 101960, 101960, 101950, 101950, 101950, 
    101960, 101950, 101960, 101940, 101930, 101910, 101920, 101960, 102010, 
    102030, 102020, 102020, 102010, 102030, 102060, 102070, 102090, 102120, 
    102140, 102160, 102170, 102150, 102150, 102150, 102150, 102130, 102100, 
    102110, 102110, 102090, 102090, 102080, 102070, 102080, 102070, 102060, 
    102000, 101990, 101990, 101980, 101980, 101950, 101970, 101970, 101950, 
    101940, 101930, 101900, 101880, 101850, 101830, 101830, 101460, 101440, 
    101420, 101410, 101390, 101390, 101390, 101380, 101370, 101380, 101390, 
    101380, 101380, 101380, 101410, 101410, 101420, 101430, 101450, 101520, 
    101570, 101600, 101630, 101670, 101710, 101740, 101790, 101830, 101880, 
    101900, 101910, 101930, 101960, 102000, 102020, 102060, 102080, 102090, 
    102120, 102110, 102110, 102130, 102140, 102120, 102110, 102120, 102110, 
    102070, 102080, 102110, 102120, 102120, 102130, 102120, 102100, 102100, 
    102110, 102130, 102110, 102110, 102090, 102080, 102040, 102020, 102010, 
    102010, 102010, 101980, 101940, 101860, 101740, 101690, 101660, 101580, 
    101560, 101570, 101560, 101510, 101470, 101430, 101410, 101420, 101390, 
    101390, 101390, 101410, 101450, 101490, 101530, 101570, 101620, 101650, 
    101690, 101700, 101710, 101720, 101790, 101810, 101880, 101880, 101890, 
    101910, 101950, 101980, 101990, 102000, 102000, 102010, 102020, 102030, 
    102040, 102110, 102180, 102220, 102210, 102220, 102210, 102260, 102300, 
    102300, 102340, 102360, 102350, 102360, 102370, 102370, 102370, 102350, 
    102340, 102340, 102330, 102290, 102250, 102220, 102200, 102160, 102120, 
    102070, 102050, 101990, 101940, 101880, 101860, 101840, 101800, 101760, 
    101750, 101730, 101700, 101540, 101460, 101490, 101500, 101480, 101440, 
    101390, 101340, 101290, 101230, 101200, 101150, 101100, 101030, 100980, 
    100940, 100900, 100880, 100850, 100840, 100820, 100790, 100780, 100790, 
    100770, 100760, 100750, 100720, 100700, 100700, 100730, 100750, 100790, 
    100840, 100860, 100880, 100880, 100860, 100880, 100900, 100950, 100980, 
    101020, 101030, 101060, 101090, 101110, 101140, 101160, 101170, 101160, 
    101180, 101200, 101210, 101230, 101230, 101250, 101270, 101290, 101290, 
    101290, 101270, 101270, 101300, 101320, 101330, 101330, 101320, 101330, 
    101350, 101370, 101370, 101360, 101370, 101400, 101430, 101440, 101480, 
    101520, 101540, 101550, 101570, 101610, 101640, 101650, 101680, 101690, 
    101730, 101770, 101790, 101830, 101860, 101880, 101900, 101910, 101920, 
    101940, 101950, 101950, 101940, 101980, 101980, 101970, 101940, 101910, 
    101910, 101920, 101900, 101890, 101860, 101830, 101840, 101830, 101810, 
    101800, 101790, 101790, 101780, 101750, 101710, 101710, 101690, 101670, 
    101660, 101650, 101600, 101580, 101590, 101570, 101550, 101530, 101510, 
    101500, 101460, 101440, 101400, 101390, 101350, 101300, 101260, 101250, 
    101200, 101130, 101090, 101040, 100980, 100900, 100870, 100830, 100790, 
    100790, 100790, 100790, 100850, 100850, 100850, 100860, 100900, 101000, 
    101070, 101170, 101250, 101300, 101360, 101430, 101450, 101490, 101520, 
    101580, 101600, 101610, 101610, 101650, 101680, 101730, 101730, 101780, 
    101790, 101810, 101820, 101830, 101850, 101880, 101920, 101940, 101950, 
    101970, 101970, 101980, 101960, 101960, 101930, 101910, 101880, 101830, 
    101770, 101710, 101720, 101680, 101680, 101690, 101670, 101640, 101640, 
    101630, 101630, 101630, 101630, 101640, 101640, 101640, 101650, 101640, 
    101630, 101610, 101590, 101540, 101500, 101500, 101510, 101500, 101480, 
    101480, 101480, 101460, 101470, 101420, 101410, 101380, 101380, 101380, 
    101400, 101390, 101370, 101360, 101310, 101290, 101220, 101210, 101180, 
    101120, 101100, 101080, 101070, 101020, 101020, 100960, 100950, 100900, 
    100860, 100820, 100770, 100730, 100670, 100650, 100580, 100580, 100530, 
    100480, 100420, 100380, 100310, 100220, 100140, 100040, 99970, 99850, 
    99720, 99650, 99530, 99460, 99390, 99360, 99340, 99270, 99300, 99300, 
    99270, 99280, 99280, 99280, 99260, 99270, 99270, 99260, 99250, 99220, 
    99260, 99250, 99300, 99360, 99400, 99440, 99470, 99460, 99530, 99560, 
    99560, 99620, 99720, 99730, 99770, 99810, 99880, 99920, 99970, 100040, 
    100090, 100140, 100190, 100260, 100290, 100340, 100390, 100460, 100510, 
    100540, 100580, 100630, 100690, 100750, 100760, 101010, 101030, 101090, 
    101110, 101120, 101130, 101150, 101170, 101180, 101200, 101180, 101190, 
    101210, 101220, 101210, 101200, 101220, 101230, 101240, 101260, 101310, 
    101340, 101360, 101390, 101410, 101420, 101460, 101490, 101500, 101530, 
    101550, 101570, 101590, 101600, 101670, 101710, 101740, 101800, 101840, 
    101870, 101900, 101930, 101940, 101980, 102000, 102020, 102040, 102040, 
    102070, 102080, 102110, 102130, 102140, 102160, 102180, 102180, 102200, 
    102200, 102200, 102200, 102200, 102210, 102240, 102240, 102240, 102250, 
    102260, 102250, 102240, 102230, 102220, 102210, 102200, 102180, 102170, 
    102160, 102140, 102130, 102120, 102100, 102080, 102070, 102050, 102030, 
    102030, 102050, 102040, 102040, 102030, 102020, 101990, 101980, 101970, 
    101970, 101970, 101940, 101970, 101940, 101930, 101930, 101930, 101920, 
    101910, 101920, 101900, 101860, _, 101830, 101810, 101790, 101810, _, 
    101770, _, _, 101730, 101690, 101650, 101610, 101620, 101580, 101560, 
    101570, 101540, 101530, _, 101500, 101460, 101430, 101410, _, 101360, 
    101340, 101310, 101290, _, 101220, 101230, 101160, _, _, 101030, 100990, 
    100980, 100980, 100920, 100960, 100980, 100930, 100920, 100910, 100920, 
    100910, 100940, 100920, 100930, 100910, 100950, 100900, 100980, 101030, 
    101130, 101160, 101220, 101260, 101280, 101310, 101330, 101340, 101370, 
    101430, 101510, 101510, 101550, 101560, 101540, 101540, 101560, 101580, 
    101580, 101580, 101580, 101570, 101590, 101590, 101580, 101600, 101610, 
    101610, 101580, 101580, 101560, 101560, 101550, 101520, 101530, 101540, 
    101510, 101490, 101460, 101410, 101380, 101320, 101310, 101290, 101280, 
    101220, 101220, 101170, 101180, 101130, 101100, 101030, 100970, 100910, 
    100870, 100750, 100720, 100670, 100590, 100510, 100430, 100310, 100230, 
    100110, 100040, 99980, 99930, 99870, 99800, 99770, 99750, 99680, 99650, 
    99630, 99580, 99540, 99500, 99500, 99440, 99380, 99370, 99360, 99340, 
    99330, 99290, 99260, 99240, 99180, 99200, 99130, 99130, 99140, 99160, 
    99150, 99180, 99170, 99140, 99190, 99190, 99210, 99220, 99160, 99160, 
    99170, 99120, 99110, 99120, 99130, 99130, 99090, 99160, 99110, 99100, 
    99130, 99110, 99140, 99170, 99220, 99260, 99300, 99350, 99390, 99400, 
    99430, 99490, 99510, 99530, 99580, 99630, 99650, 99680, 99710, 99780, 
    99850, 99920, 99970, 100020, 100040, 100070, 100130, 100180, 100220, 
    100260, 100300, 100330, 100370, 100390, 100420, 100450, 100480, 100490, 
    100520, 100530, 100530, 100550, 100540, 100580, 100590, 100580, 100580, 
    100560, 100550, 100590, 100600, 100610, 100640, 100640, 100650, 100670, 
    100680, 100680, 100680, 100700, 100670, 100670, 100660, 100680, 100670, 
    100670, 100650, 100640, 100640, 100630, 100620, 100610, 100600, 100580, 
    100590, 100580, 100570, 100560, 100530, 100510, 100520, 100510, 100490, 
    100480, 100450, 100430, 100420, 100430, 100420, 100430, 100430, 100430, 
    100440, 100430, 100450, 100450, 100460, 100480, 100480, 100490, 100530, 
    100550, 100560, 100560, 100570, 100550, 100520, 100510, 100490, 100480, 
    100480, 100490, 100470, 100450, 100400, 100380, 100380, 100360, 100350, 
    100370, 100330, 100370, 100430, 100450, 100500, 100520, 100510, 100510, 
    100450, 100490, 100510, 100510, 100460, 100440, 100420, 100410, 100410, 
    100350, 100360, 100280, 100250, 100260, 100210, 100100, 100040, 100010, 
    99970, 99930, 99800, 99710, 99580, 99470, 99370, 99240, 99150, 99060, 
    99100, 99080, 99100, 99190, 99190, 99180, 99290, 99310, 99290, 99240, 
    99220, 99200, 99280, 99270, 99290, 99280, 99310, 99290, 99340, 99360, 
    99360, 99430, 99410, 99530, 99640, 99710, 99760, 99760, 99820, 99830, 
    99940, 99970, 100020, 100040, 100030, 100000, 99970, 99950, 99980, 99960, 
    99950, 99990, 100000, 100010, 100030, 100070, 100090, 100170, 100190, 
    100190, 100240, 100230, 100280, 100240, 100310, 100340, 100360, 100360, 
    100360, 100360, 100430, 100440, 100460, 100530, 100600, 100670, 100730, 
    100750, 100800, 100850, 100870, 100980, 100990, 100930, 101000, 101050, 
    101060, 101160, 101220, 101260, 101220, 101320, 101340, 101340, 101330, 
    101320, 101310, 101300, 101290, 101290, 101270, 101250, 101210, 101160, 
    101120, 101140, 101140, 101130, 101100, 101090, 101020, 100980, 100960, 
    100900, 100890, 100890, 100880, 100870, 100850, 100860, 100830, 100850, 
    100830, 100820, 100800, 100810, 100790, 100770, 100750, 100730, 100670, 
    100630, 100660, 100650, 100620, 100590, 100550, 100490, 100450, 100480, 
    100470, 100450, 100440, 100440, 100430, 100420, 100400, 100410, 100430, 
    100430, 100450, 100440, 100450, 100430, 100420, 100410, 100370, 100360, 
    100370, 100390, 100380, 100370, 100370, 100360, 100370, 100380, 100370, 
    100380, 100400, 100430, 100450, 100470, 100510, 100530, 100560, 100580, 
    100610, 100630, 100650, 100670, 100680, 100710, 100720, 100740, 100750, 
    100790, 100820, 100830, 100850, 100890, 100920, 100970, 100980, 101020, 
    101050, 101060, 101100, 101130, 101130, 101170, 101180, 101200, 101220, 
    101230, 101250, 101270, 101300, 101320, 101330, 101350, 101360, 101390, 
    101390, 101410, 101410, 101420, 101430, 101430, 101450, 101480, 101500, 
    101490, 101490, 101510, 101520, 101510, 101540, 101550, 101550, 101580, 
    101590, 101600, 101620, 101650, 101650, 101660, 101650, 101670, 101690, 
    101690, 101700, 101740, 101770, 101810, 101830, 101870, 101880, 101920, 
    101940, 101960, 101990, 102010, 102030, 102070, 102090, 102120, 102130, 
    102140, 102160, 102160, 102160, 102190, 102190, 102200, 102220, 102230, 
    102230, 102240, 102250, 102270, 102260, 102290, 102260, 102260, 102270, 
    102260, 102250, 102250, 102260, 102270, 102260, 102280, 102280, 102280, 
    102290, 102270, 102260, 102260, 102270, 102260, 102250, 102270, 102280, 
    102270, 102270, 102260, 102250, 102220, 102210, 102200, 102220, 102190, 
    102210, 102200, 102200, 102190, 102180, 102180, 102150, 102150, 102120, 
    102090, 102090, 102100, 102110, 102090, 102070, 102070, 102040, 102030, 
    102000, 102000, 101980, 101980, 101970, 101960, 101950, 101940, 101920, 
    101910, 101890, 101870, 101890, 101870, 101830, 101810, 101800, 101780, 
    101780, 101770, 101760, 101740, 101730, 101720, 101700, 101700, 101670, 
    101590, 101570, 101590, 101590, 101570, 101600, 101610, 101620, 101600, 
    101600, 101570, 101600, 101600, 101600, 101620, 101610, 101610, 101580, 
    101550, 101540, 101540, 101510, 101500, 101490, 101470, 101440, 101430, 
    101400, 101380, 101360, 101350, 101340, 101350, 101350, 101320, 101300, 
    101300, 101280, 101290, 101300, 101330, 101350, 101360, 101370, 101390, 
    101390, 101400, 101430, 101430, 101450, 101490, 101510, 101530, 101550, 
    101560, 101590, 101610, 101610, 101630, 101650, 101660, 101680, 101680, 
    101720, 101750, 101770, 101790, 101780, 101780, 101810, 101800, 101800, 
    101780, 101760, 101760, 101760, 101770, 101740, 101740, 101720, 101690, 
    101650, 101660, 101630, 101620, 101600, 101590, 101570, 101550, 101500, 
    101460, 101460, 101440, 101440, 101420, 101410, 101400, 101380, 101350, 
    101390, 101400, 101400, 101410, 101410, 101390, 101410, 101440, 101440, 
    101480, 101490, 101550, 101620, 101660, 101690, 101700, 101720, 101760, 
    101780, 101780, 101760, 101750, 101730, 101710, 101690, 101720, 101750, 
    101750, 101740, 101720, 101720, 101730, 101710, 101690, 101700, 101720, 
    101710, 101710, 101720, 101730, 101700, 101690, 101690, 101680, 101650, 
    101640, 101640, 101610, 101570, 101590, 101600, 101560, 101530, 101500, 
    101480, 101460, 101470, 101460, 101450, 101440, 101440, 101440, 101430, 
    101430, 101390, 101370, 101350, 101370, 101350, 101340, 101320, 101340, 
    101350, 101340, 101340, 101360, 101360, 101370, 101380, 101390, 101420, 
    101440, 101470, 101490, 101520, 101570, 101610, 101640, 101670, 101690, 
    101720, 101750, 101760, 101770, 101800, 101800, 101840, 101840, 101860, 
    101880, 101880, 101920, 101930, 101950, 102000, 102020, 102050, 102090, 
    102130, 102190, 102210, 102240, 102300, 102330, 102340, 102360, 102380, 
    102420, 102410, 102420, 102420, 102440, 102440, 102470, 102480, 102490, 
    102470, 102500, 102490, 102500, 102520, 102540, 102560, 102590, 102610, 
    102630, 102660, 102660, 102660, 102690, 102690, 102700, 102690, 102660, 
    102670, 102660, 102650, 102640, 102630, 102620, 102600, 102590, 102570, 
    102560, 102550, 102560, 102580, 102560, 102540, 102520, 102500, 102480, 
    102450, 102430, 102420, 102330, 102360, 102420, 102420, 102370, 102270, 
    102280, 102290, 102270, 102240, 102220, 102170, 102110, 102090, 102020, 
    102080, 102050, 102030, 102030, 102000, 102050, 102050, 102020, 102000, 
    102060, _, 102080, 102110, 102130, 102160, 102170, 102190, 102200, 
    102220, 102250, 102200, 102270, 102290, 102260, 102340, 102340, _, _, _, 
    102360, _, 102410, 102370, 102350, 102380, 102350, 102360, _, _, 102350, 
    _, 102310, 102290, 102270, 102240, 102200, _, 102230, _, 102200, _, _, 
    102270, 102320, 102330, 102290, _, 102300, _, 102330, 102350, 102340, _, 
    102370, 102340, 102360, _, 102360, 102370, 102310, _, 102380, 102370, _, 
    102380, 102400, 102360, 102330, 102350, 102360, 102300, 102320, 102290, 
    102290, _, _, _, _, 102250, 102250, _, 102250, 102210, 102230, 102210, 
    102240, 102220, 102260, 102300, 102300, 102290, 102310, 102330, 102300, 
    _, _, 102280, _, 102340, 102310, 102340, 102330, 102380, 102380, 102380, 
    102370, 102380, 102370, 102370, 102390, 102390, 102410, 102370, 102370, 
    102360, 102370, 102330, 102340, 102350, 102340, 102310, 102240, 102210, 
    102210, 102210, 102170, 102140, 102130, 102140, 102090, 102060, 102030, 
    102010, 102020, 102000, 101970, 101940, 101950, 101910, _, 101830, 
    101820, 101810, 101770, 101740, _, 101650, 101630, _, 101560, 101530, 
    101490, 101480, 101440, 101370, _, 101300, 101280, 101280, 101250, 
    101230, 101240, 101230, 101180, 101150, 101120, 101100, 101090, 101050, 
    101030, 101010, 101030, 101050, 101050, 101080, 101060, 101040, 101040, 
    101060, 101010, 100950, 100900, 100860, 100790, 100750, 100680, 100700, 
    100660, 100660, 100650, 100660, 100660, 100670, 100710, 100740, 100750, 
    100770, 100790, 100770, 100730, 100700, 100700, 100630, 100640, 100670, 
    100730, 100830, 100880, 100930, 100930, 100970, 100980, 101020, 101050, 
    101060, 101090, 101090, 101140, 101170, 101190, 101220, 101330, 101230, 
    _, 101310, 101340, 101340, 101370, 101410, 101390, 101420, 101470, 
    101480, 101440, 101480, 101600, 101600, 101620, 101620, 101660, 101630, 
    101640, 101640, 101610, 101560, 101520, 101490, 101520, 101520, 101500, 
    101510, 101490, 101490, 101500, 101540, 101530, 101560, 101570, 101570, 
    101600, 101630, 101630, 101610, 101620, 101620, 101630, 101650, 101660, 
    101700, 101700, 101700, 101680, 101710, 101730, 101750, 101750, 101750, 
    101750, 101750, 101750, 101770, 101780, 101780, 101780, 101790, 101800, 
    101770, 101760, 101730, 101700, 101690, 101760, 101780, 101800, 101820, 
    101810, 101800, 101780, 101770, 101770, 101750, 101750, 101770, 101760, 
    101750, 101810, 101810, 101820, 101830, 101800, 101770, 101750, 101720, 
    101690, 101660, 101680, 101710, 101690, 101680, 101670, 101650, 101640, 
    101620, 101590, 101560, 101560, 101560, 101520, 101520, 101560, 101530, 
    101550, 101540, 101520, 101500, 101500, 101470, 101450, 101420, 101400, 
    101410, 101380, 101350, 101320, 101270, 101350, 101320, 101270, 101220, 
    101160, 101090, 101060, 101020, 100960, 100900, 100820, 100800, 100710, 
    100650, 100630, 100580, 100530, 100490, 100470, 100410, 100440, 100390, 
    100380, 100350, 100310, 100280, 100290, 100300, 100330, 100340, 100370, 
    100400, 100420, 100430, 100420, _, 100410, 100350, _, _, 100270, _, _, 
    100200, 100190, _, 100110, 100070, 100070, _, _, 100000, 100050, 100060, 
    100110, 100160, 100180, 100230, 100280, _, 100370, 100410, 100450, 
    100500, 100570, _, 100680, 100700, _, 100770, 100820, 100860, 100890, 
    100940, 100940, 100990, 101010, 101020, 101040, 101080, 101080, 101110, 
    101110, 101140, 101130, 101160, _, 101200, 101240, 101260, 101300, _, 
    101400, 101450, 101500, 101550, 101610, 101660, _, 101760, 101790, _, 
    101870, _, _, 101970, 102010, _, 102050, 102080, 102130, 102150, 102170, 
    102200, 102240, 102290, 102320, 102340, 102350, _, 102340, 102350, _, 
    102410, 102410, 102460, 102420, 102410, 102490, 102520, 102520, _, _, 
    102520, _, 102490, 102500, 102480, 102490, 102480, _, 102480, 102470, 
    102440, _, _, 102410, _, 102360, 102340, 102320, 102320, 102290, 102270, 
    102240, 102190, 102110, 102000, 101990, 101960, 101960, 101930, 101860, 
    101870, 101920, 101900, 101860, 101850, 101830, 101870, 101870, 101900, 
    101870, _, 101890, 101930, 101950, 101970, 101960, 102020, 102050, 
    101990, 102010, 102050, 102090, 102150, 102160, 102180, 102190, 102210, 
    102230, 102310, 102300, 102330, 102360, 102380, 102380, 102360, 102470, 
    102450, 102420, _, 102490, _, _, 102480, _, 102440, 102460, _, 102400, _, 
    102340, 102390, _, 102410, _, 102400, 102430, 102420, _, _, _, _, _, _, 
    102390, 102360, 102340, _, 102390, 102350, 102370, _, 102340, 102340, 
    102430, _, _, 102400, _, 102400, 102420, 102400, 102400, 102410, 102430, 
    102430, 102450, 102430, 102460, 102470, 102460, _, 102450, _, 102470, 
    102470, 102480, _, 102460, 102440, _, _, _, 102400, _, _, _, _, _, 
    102400, 102400, 102400, 102400, 102370, 102360, 102340, 102320, _, 
    102310, 102310, 102320, 102310, 102280, _, 102280, 102250, 102250, _, 
    102260, 102260, 102280, 102290, 102310, _, 102330, 102320, _, _, _, 
    102330, _, _, 102240, 102260, 102300, 102310, 102290, 102250, _, 102260, 
    _, _, 102260, 102250, 102260, _, 102320, 102340, 102340, _, _, 102370, _, 
    102370, 102360, 102350, _, 102340, 102350, 102340, 102340, 102310, 
    102310, 102300, _, 102250, 102220, _, 102170, 102150, 102130, 102090, 
    102060, 102010, 101960, 101920, 101860, 101810, 101770, 101720, 101680, 
    101650, 101640, 101600, 101590, 101530, 101510, 101470, 101410, 101380, 
    101330, 101300, 101290, 101280, 101260, 101250, 101230, 101190, 101180, 
    101160, 101130, 101120, 101110, 101080, 101070, 101040, 101040, 101050, 
    101040, 101030, 101010, 101000, 100990, 100970, 100980, 100980, 100990, 
    101020, _, 101060, 101070, 101090, 101110, 101120, 101120, 101130, 
    101130, 101150, 101150, 101180, 101190, 101220, 101240, 101260, 101260, 
    _, 101280, 101280, 101290, 101320, 101360, 101380, 101400, 101420, 
    101430, 101420, 101430, 101440, 101420, 101410, 101410, 101360, 101340, 
    101350, 101370, 101360, 101370, 101350, 101360, 101350, 101360, 101360, 
    101360, 101350, 101370, 101380, 101390, 101410, 101410, 101430, 101430, 
    101420, 101420, 101450, 101430, 101440, 101460, 101470, 101470, 101500, 
    101500, 101500, 101500, 101510, 101510, 101510, 101500, 101510, 101540, 
    101560, 101580, 101590, 101600, 101620, 101630, 101640, 101650, 101650, 
    101680, 101690, 101700, 101730, 101730, 101750, 101770, 101780, 101770, 
    101780, 101790, 101810, 101830, 101810, 101830, 101840, 101840, 101840, 
    101850, 101870, 101850, 101850, 101840, 101830, 101810, 101790, 101790, 
    101770, 101760, 101740, 101720, 101690, 101650, 101610, 101580, 101550, 
    101520, 101490, 101470, 101470, 101460, 101450, 101410, 101410, 101400, 
    101380, 101350, 101330, 101340, 101320, 101300, 101280, 101260, 101250, 
    101230, 101230, 101220, 101220, 101210, 101210, 101220, 101220, 101230, 
    101250, 101260, 101290, 101320, 101340, 101360, 101380, 101400, 101430, 
    101450, 101470, 101490, 101520, 101570, 101620, 101670, 101700, 101740, 
    101770, 101790, 101810, 101840, 101900, 101990, 102030, 102070, 102150, 
    102220, 102270, 102310, 102360, 102380, 102400, 102420, 102470, 102520, 
    102580, 102610, 102640, 102680, 102700, 102710, 102720, 102730, 102720, 
    102730, 102780, 102800, 102810, 102800, 102830, 102860, 102850, 102830, 
    102830, 102840, 102820, 102790, 102760, 102730, 102720, 102700, 102690, 
    102660, 102630, 102610, 102600, 102560, 102550, 102520, 102460, 102470, 
    102480, 102490, 102500, 102520, 102510, 102490, 102510, 102480, 102440, 
    102460, 102430, 102400, 102390, 102380, 102320, 102290, 102270, 102240, 
    102200, 102140, 102050, 102020, 101930, 101870, 101850, 101790, 101730, 
    101680, 101590, 101540, 101510, 101400, 101330, 101230, 101170, 101130, 
    101070, 101050, 101050, 101030, 101030, 100990, 100960, 100940, 100910, 
    100940, 100930, 100940, 100970, 101000, 101010, 101080, 101150, 101230, 
    101230, 101240, 101210, 101190, 101160, 101130, 101140, 101140, 101130, 
    101160, 101180, 101170, 101140, 101120, 101090, 101080, 101070, 101070, 
    101080, 101050, 101020, 101020, 101000, 100980, 100950, 100920, 100920, 
    100910, 100900, 100920, 100960, 100990, 101020, 101020, 101050, 101060, 
    101060, 101070, 101070, 101080, 101100, 101070, 101090, 101110, 101110, 
    101110, 101110, 101100, 101110, 101130, 101140, 101160, 101200, 101230, 
    101280, 101320, 101410, 101480, 101530, 101560, 101600, 101620, 101640, 
    101670, 101650, 101720, 101780, 101840, 101890, 101950, 101960, 101980, 
    102050, 102120, 102200, 102220, 102240, 102290, 102340, 102380, 102420, 
    102450, 102490, 102540, 102550, 102550, 102580, 102610, 102630, 102670, 
    102710, 102760, 102770, 102780, 102830, 102840, 102850, 102870, 102880, 
    102900, 102880, 102880, 102870, 102850, 102820, 102820, 102770, 102710, 
    102630, 102560, 102520, 102440, 102390, 102360, 102330, 102300, 102240, 
    102180, 102130, 102090, 102030, 101980, 101940, 101910, 101880, 101850, 
    101830, 101810, 101790, 101770, 101790, 101780, 101790, 101800, 101800, 
    101800, 101790, 101830, 101860, 101870, 101900, 101930, 101960, 101970, 
    101990, 102010, 102030, 102030, 102040, 102050, 102050, 102050, 102050, 
    102020, 102000, 102000, 101970, 101950, 101930, 101910, 101870, 101870, 
    101860, 101860, 101830, 101800, 101770, 101740, 101700, 101660, 101630, 
    101610, 101580, 101570, 101570, 101600, 101580, 101550, 101500, 101500, 
    101480, 101450, 101420, 101470, 101450, 101420, 101390, 101420, 101420, 
    101400, 101400, 101360, 101430, 101410, 101390, 101430, 101420, 101440, 
    101470, 101460, 101470, 101500, 101520, 101540, 101550, 101560, 101560, 
    101570, 101570, 101600, 101620, 101640, 101660, 101680, 101710, 101740, 
    101740, 101740, 101750, 101760, 101750, 101750, 101750, 101750, 101770, 
    101780, 101800, 101800, 101820, 101830, 101830, 101830, 101830, 101830, 
    101850, 101870, 101880, 101880, 101890, 101890, 101880, 101870, 101850, 
    101840, 101810, 101810, 101760, 101750, 101740, 101700, 101650, 101590, 
    101530, 101470, 101420, 101370, 101390, 101320, 101270, 101260, 101210, 
    101170, 101150, 101130, 101090, 101080, 101080, 101070, 101110, 101110, 
    101130, 101160, 101190, 101220, 101270, 101290, 101320, 101350, 101340, 
    101350, 101370, 101370, 101380, 101390, 101390, 101380, 101370, 101350, 
    101360, 101360, 101350, 101310, 101280, 101260, 101270, 101260, 101240, 
    101210, 101210, 101200, 101180, 101180, 101160, 101160, 101160, 101150, 
    101160, 101170, 101170, 101190, 101210, 101210, 101220, 101210, 101210, 
    101170, 101180, 101150, 101170, 101210, 101230, 101210, 101230, 101300, 
    101300, 101310, 101330, 101350, 101360, 101410, 101450, 101490, 101520, 
    101520, 101510, 101530, 101570, 101590, 101580, 101570, 101550, 101540, 
    101520, 101520, 101520, 101520, 101490, 101500, 101500, 101460, 101440, 
    101450, 101380, 101330, 101340, 101310, 101340, 101340, 101320, 101310, 
    101300, 101240, 101220, 101200, 101100, 101130, 101020, 101030, 100980, 
    100950, 100960, 100900, 100860, 100880, 100820, 100770, 100830, 100850, 
    100820, 100810, 100820, 100840, 100810, 100780, 100830, 100830, 100800, 
    100770, 100760, 100700, 100670, 100650, 100520, 100480, 100480, 100460, 
    100390, 100400, 100320, 100280, 100260, 100280, 100260, 100190, 100190, 
    100190, 100170, 100170, 100190, 100190, 100190, 100170, 100160, 100150, 
    _, 100220, 100240, 100270, 100340, 100420, 100430, 100450, 100480, 
    100500, 100510, 100530, 100570, 100630, 100670, 100700, 100730, 100760, 
    100790, 100800, 100820, 100830, 100890, 100920, 100960, 100990, 101020, 
    101060, 101080, _, 101100, 101120, 101130, 101140, 101170, 101190, 
    101230, 101260, 101270, 101290, 101320, 101330, 101330, 101330, 101320, 
    101310, 101300, 101290, 101270, 101240, 101220, _, 101110, 101060, 
    101000, 100960, 100960, 100950, 100920, 100890, 100890, 100880, 100850, 
    100830, 100810, 100740, 100660, 100560, 100490, 100370, 100320, 100280, 
    100210, 100140, 100060, 99930, 99850, 99800, 99750, 99740, 99720, 99730, 
    99720, 99730, 99700, 99740, 99740, 99760, 99760, 99740, 99740, 99750, 
    99740, 99730, 99740, 99770, 99770, 99750, 99760, 99760, 99770, 99760, 
    99840, 99880, 99880, 99910, 100020, 100080, 100120, 100150, 100220, 
    100270, 100350, 100420, 100450, 100500, 100570, 100560, 100620, 100720, 
    100760, 100800, 100870, 100940, 101000, 101030, 101080, 101070, 101030, 
    101040, 101010, 101020, 100980, 100950, 100940, 100910, 100860, 100790, 
    100750, 100720, 100670, 100660, 100640, 100620, 100640, 100640, 100680, 
    100710, 100730, 100780, 100810, 100880, 100920, 100940, 100960, 100960, 
    100970, 100950, 100960, 100930, 100870, 100790, 100720, 100650, 100580, 
    100550, 100520, 100500, 100520, 100540, 100590, 100600, 100680, 100720, 
    100760, 100810, 100890, 100920, 100990, 101060, 101120, 101190, 101250, 
    101270, 101390, 101450, 101480, 101510, 101540, 101570, 101570, 101570, 
    101550, 101540, 101540, 101500, 101420, 101370, 101330, 101260, 101200, 
    101160, 101130, 101130, 101150, 101170, 101240, 101280, 101340, 101400, 
    101420, 101450, 101480, 101510, 101570, 101600, 101650, 101690, 101720, 
    101730, 101720, 101730, 101730, 101750, 101720, 101690, 101650, 101630, 
    101620, 101590, 101580, 101530, 101510, 101450, 101410, 101350, 101350, 
    101320, 101290, 101230, 101190, 101190, 101160, 101120, 101060, 101080, 
    101050, 101060, 101100, 101160, 101220, 101270, 101360, 101410, 101450, 
    101500, 101570, 101620, 101670, 101660, 101700, 101750, 101780, 101790, 
    101830, _, 101850, 101850, 101830, 101830, 101820, 101810, 101780, 
    101800, 101800, 101750, 101740, 101730, 101690, 101670, 101670, 101670, 
    101620, 101590, 101550, 101530, 101500, 101440, 101390, 101320, 101290, 
    101230, 101220, 101130, 101080, 101050, 101020, 101030, 101020, 101010, 
    101010, 101010, 100980, 101000, 101030, 101040, 101060, 101070, 101040, 
    101050, 101130, 101230, 101270, 101290, 101300, 101310, 101320, 101350, 
    101350, 101360, 101400, 101460, 101470, 101470, 101440, 101500, 101580, 
    101660, 101680, 101720, 101740, 101760, 101780, 101770, 101780, 101820, 
    101790, 101790, 101790, 101780, 101790, 101820, 101810, 101780, 101800, 
    101810, 101790, 101770, 101780, 101790, 101790, 101800, 101790, 101750, 
    101730, 101680, 101660, 101610, 101590, 101570, 101530, 101460, 101460, 
    101440, 101390, 101380, 101340, 101300, 101260, 101230, 101190, 101180, 
    101170, 101170, 101180, 101170, 101180, 101170, 101170, 101170, 101150, 
    101140, 101140, 101160, 101160, 101180, 101210, 101270, 101280, 101300, 
    101340, 101360, 101400, 101410, 101430, 101450, 101490, 101520, 101580, 
    101620, 101650, 101710, 101720, 101730, 101750, 101780, 101750, 101800, 
    101810, 101820, 101810, 101780, 101750, 101720, 101650, 101640, 101560, 
    101480, 101450, 101390, 101310, 101310, 101290, 101260, 101230, 101200, 
    101150, 101110, 101050, 101000, 100940, 100970, 100940, 100920, 100900, 
    100880, 100920, 100890, 100900, 100920, 100930, 100980, 101010, 101040, 
    101070, 101120, 101130, 101200, 101220, 101260, 101280, 101350, 101360, 
    101350, 101400, 101430, 101510, 101510, 101540, 101560, 101570, 101590, 
    101590, 101580, 101590, 101590, 101580, 101610, 101610, 101620, 101600, 
    101610, 101600, 101570, 101550, 101530, 101510, 101500, 101480, 101480, 
    _, 101430, 101430, _, 101380, 101380, 101360, 101360, 101350, 101360, 
    101360, 101380, 101390, 101400, 101420, 101440, 101450, 101470, 101470, 
    101490, 101530, 101540, 101560, _, _, _, _, _, _, _, 101800, 101830, 
    101890, 101920, 101950, 102000, 102050, 102110, 102140, 102170, 102210, 
    102240, 102250, 102290, 102320, 102350, 102380, 102410, 102450, 102490, 
    102520, 102570, 102590, 102610, 102650, 102700, 102740, 102770, 102770, 
    102820, 102870, 102890, 102910, 102940, 102950, 102960, 102960, 102950, 
    102950, 102950, 102910, 102860, 102800, 102770, 102740, 102710, 102660, 
    102630, 102610, 102540, 102490, 102440, 102340, 102280, 102180, 102140, 
    102060, 101990, 101950, 101870, 101830, 101740, 101670, 101560, 101490, 
    101390, 101260, 101110, 100940, 100780, 100730, 100720, 100740, 100740, 
    100710, 100570, 100410, 100290, 100220, 100120, 100000, 99890, 99710, 
    99390, 99120, 98740, 98360, 98170, 97920, 97620, 97390, 97210, 97080, 
    96920, 96780, 96640, 96480, 96350, 96240, 96140, 96030, 96000, 95980, 
    96030, 96080, 96130, 96190, 96340, 96450, 96610, 96830, 97040, 97170, 
    97340, 97440, 97560, 97660, 97730, 97820, 97930, 97990, 98120, 98200, 
    98250, 98330, 98400, 98460, 98550, 98600, 98670, 98710, 98770, 98840, 
    98880, 98910, 99030, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 102120, 
    102170, 102220, 102270, 102320, 102380, 102420, 102420, 102440, 102440, 
    102490, 102530, 102550, 102590, 102610, 102650, 102650, 102680, 102700, 
    102740, 102760, 102770, 102780, 102830, 102850, 102890, 102900, 102880, 
    102920, 102910, 102920, _, 102890, 102880, 102900, 102900, 102890, 
    102890, 102900, 102890, 102880, 102910, 102920, 102930, 102920, 102970, 
    103010, 103020, 103050, 103060, 103100, 103100, 103120, 103120, 103130, 
    103140, 103160, 103140, 103130, 103150, 103130, 103120, 103100, 103060, 
    103030, 103030, 102990, 102960, 102930, 102900, 102880, 102860, 102870, 
    102870, 102820, 102790, 102760, 102770, 102750, 102730, 102690, 102690, 
    102670, 102670, 102660, 102640, 102580, 102620, 102610, 102570, 102580, 
    102560, 102600, 102580, 102590, 102590, 102590, 102610, 102570, 102560, 
    102530, 102490, 102500, _, 102450, 102410, 102380, 102310, _, 102300, 
    102270, 102230, 102180, 102120, 102110, 102050, 102010, 102010, 102000, 
    101970, 101970, 101950, 101920, 101880, 101850, 101810, 101750, 101780, 
    101720, 101650, 101620, 101560, 101520, 101450, 101410, 101380, 101350, 
    101310, 101270, 101230, 101160, 101100, 101090, 101090, 101090, 101070, 
    101040, 101010, 100960, 100930, 100880, 100850, 100840, 100820, 100800, 
    100770, 100740, 100740, 100740, 100720, 100710, 100710, 100690, 100690, 
    100710, 100720, 100720, 100720, 100760, 100810, 100820, 100870, 100890, 
    100920, 100950, _, 101000, 101010, 101020, 101040, 101060, 101070, 
    101090, 101110, 101100, 101130, 101120, 101140, 101130, 101130, 101110, 
    101130, 101140, 101150, 101160, 101180, 101190, 101220, 101220, 101230, 
    101240, 101260, 101270, 101290, 101310, 101350, 101390, 101380, 101390, 
    101400, 101410, 101420, 101440, 101420, 101430, 101430, 101420, 101370, 
    101380, 101380, 101360, 101340, 101300, 101250, 101240, 101190, 101140, 
    101130, 101090, 101040, 101020, 100960, 100910, 100860, 100800, 100770, 
    100650, 100590, 100490, 100340, 100240, 100130, 100080, 99970, 99770, 
    99650, 99510, 99320, 99150, 98970, 98800, 98590, 98380, 98180, 98090, 
    98110, 98210, 98350, 98480, 98560, 98670, 98730, 98820, 98880, 98950, 
    98990, 99110, 99100, 99110, 99140, 99160, 99210, 99240, 99290, 99310, 
    99360, 99400, 99390, 99430, 99540, 99570, 99640, 99680, 99720, 99780, 
    99810, 99870, 99930, 99980, 100060, 100150, 100150, 100180, 100240, 
    100240, 100270, 100290, 100290, 100300, 100340, 100380, 100410, 100460, 
    100460, 100490, 100510, 100540, 100560, 100570, 100590, 100620, 100640, 
    100630, 100650, 100630, 100610, 100580, 100530, 100480, 100410, 100350, 
    _, _, 100140, 100090, 100010, 99910, 99810, _, 99600, 99470, _, 99290, 
    99240, 99200, 99180, 99170, 99160, 99150, 99100, 99060, 99060, 99060, 
    99060, 99080, 99130, 99230, 99330, 99420, 99500, 99610, 99700, 99800, 
    99860, 99910, 99970, 100030, 100120, 100170, 100200, 100270, 100330, 
    100400, 100470, 100530, 100570, 100610, 100630, 100670, 100710, 100730, 
    100750, 100770, 100780, 100800, 100810, 100840, 100840, 100830, 100830, 
    100830, 100830, 100820, 100840, 100810, 100770, 100730, 100720, 100700, 
    100660, 100620, 100570, 100550, 100520, 100500, 100460, 100430, 100410, 
    100400, 100370, 100350, 100300, 100300, 100270, 100240, 100240, 100240, 
    100230, 100220, 100200, 100170, 100190, 100200, 100190, 100210, 100180, 
    100190, 100200, 100200, 100160, 100170, 100190, 100190, 100200, 100190, 
    100210, 100210, 100220, 100230, 100260, 100250, 100280, 100320, 100330, 
    100360, 100380, 100420, 100400, 100410, 100400, _, 100380, 100380, 
    100320, 100270, 100240, 100200, 100150, 100080, 99940, 99830, 99690, 
    99670, 99550, 99400, 99340, 99250, 99280, 99280, 99250, 99190, 99080, 
    99020, 98980, 98890, 98820, 98720, 98660, 98570, 98490, 98330, 98120, 
    97880, 97820, 97690, 97700, 97650, 97610, 97620, 97590, 97570, 97500, 
    97460, 97410, 97400, 97380, 97380, 97440, 97510, 97580, 97680, 97800, 
    97920, 97980, 98120, 98180, 98170, 98300, 98280, 98390, 98540, 98750, 
    98920, 99000, 99100, 99270, 99420, 99550, 99610, 99670, 99760, 99860, 
    99970, 100010, 100090, 100160, 100210, 100250, 100310, 100350, 100380, 
    100410, 100470, 100480, 100510, 100540, 100560, 100590, 100610, 100630, 
    100660, 100670, 100650, 100630, 100640, 100610, 100600, 100580, 100570, 
    100580, 100590, 100620, 100600, 100630, 100630, 100620, 100630, 100650, 
    100710, 100750, 100780, 100830, 100870, 100890, 100950, 101010, 101060, 
    101120, 101170, 101210, 101260, 101280, 101290, 101330, 101380, 101400, 
    101430, 101440, 101480, 101520, 101560, 101570, 101600, 101640, 101660, 
    101680, 101710, 101730, 101720, 101740, 101780, 101750, 101760, 101760, 
    101770, 101770, 101800, 101780, 101800, 101760, 101760, 101720, 101710, 
    101670, 101580, 101490, 101420, 101390, 101310, 101330, 101310, 101220, 
    101190, 101170, 101160, 101160, 101090, 101100, 101080, 101110, 101100, 
    101110, 101090, 101080, 101040, 101010, 100980, 100920, 100900, 100870, 
    100830, 100790, 100710, 100700, 100690, 100660, 100590, 100540, 100510, 
    100420, 100370, 100280, 100210, 100090, 100100, 100030, 99980, 99880, 
    99840, 99750, 99630, 99550, 99470, 99380, 99300, 99180, 99050, 98990, 
    98960, 98940, 98910, 98880, 98820, 98820, 98770, 98740, 98740, 98730, 
    98720, _, 98710, 98700, 98690, 98720, 98680, 98680, 98710, 98720, 98710, 
    98740, 98770, 98770, 98770, 98730, 98760, 98790, 98810, 98850, 98850, 
    98870, 98880, 98910, 98930, 98960, 98980, 99050, 99100, 99150, 99220, 
    99290, 99350, 99390, 99430, 99550, 99580, 99600, 99660, 99710, 99750, 
    99760, 99740, 99740, 99730, 99720, 99700, 99660, 99650, 99640, 99560, 
    99550, 99520, 99510, 99500, 99480, 99440, 99400, 99380, 99390, _, 99440, 
    99490, 99510, 99540, 99590, 99640, 99700, 99770, 99830, 99860, 99920, 
    99980, 100030, 100100, 100200, 100290, 100400, 100480, 100560, 100620, 
    100660, 100730, 100800, 100860, 100890, 100920, 100980, 101000, 101010, 
    101020, 101040, 101000, 100950, 100900, 100910, 100990, 101100, 101140, 
    101150, 101160, 101150, 101120, 101110, 101150, 101200, 101240, 101300, 
    101360, 101400, 101400, 101370, 101320, 101320, 101300, 101290, 101270, 
    101260, 101240, 101250, 101220, 101200, 101180, 101140, 101130, 101110, 
    101100, 101090, 101100, 101100, 101080, 101070, 101040, 101080, 101050, 
    101020, 100990, 100940, 100910, 100850, 100770, 100700, 100650, 100580, 
    100550, 100540, 100540, 100570, 100570, 100530, 100510, 100490, 100490, 
    100420, 100380, 100390, 100370, 100290, 100220, 100190, 100140, 100090, 
    100010, 99920, 99850, 99780, 99730, 99670, 99610, 99560, 99530, 99450, 
    99350, 99310, 99320, 99380, 99430, 99440, 99500, 99510, 99520, 99600, 
    99600, 99590, 99590, 99610, 99640, 99620, 99750, 99770, 99800, 99850, 
    99840, 99860, 99870, 99900, 99900, 99950, 99980, 99960, 99970, 99970, 
    99970, 99990, 100030, 100060, 100090, 100110, 100120, 100100, 100110, 
    100140, 100160, 100180, 100190, 100180, 100210, 100260, 100270, 100300, 
    100290, 100320, 100330, 100380, 100400, 100450, 100490, 100540, 100550, 
    100620, 100730, 100820, 100870, 100930, 100990, 101050, 101110, _, 
    101190, 101200, 101290, 101330, 101380, 101450, 101500, 101530, 101590, 
    101670, 101730, 101770, 101840, 101890, 101930, 101980, 102050, 102110, 
    102170, 102200, 102240, 102310, 102380, 102410, 102470, 102510, 102540, 
    102600, 102630, 102670, 102710, 102730, 102760, 102810, 102830, 102840, 
    102830, 102850, 102860, 102880, 102890, 102900, 102900, _, 102870, 
    102870, 102840, 102830, 102820, 102770, 102750, 102710, 102660, 102620, 
    102580, 102520, 102460, 102390, 102310, 102210, 102140, 102050, 102010, 
    101970, 101940, 101900, 101860, 101820, 101770, 101690, 101640, _, 
    101510, 101480, 101430, 101380, 101340, 101260, 101140, 101090, 101050, 
    100970, 100860, 100770, 100640, 100500, 100410, 100320, 100210, 100140, 
    100010, 99970, 99890, 99860, 99810, 99770, 99740, 99730, 99730, 99710, 
    99740, 99780, 99800, 99820, 99820, 99830, 99890, 99920, 99900, 99870, 
    99880, 99870, 99890, 99870, 99840, _, 99700, _, 99590, 99550, 99520, 
    99510, 99480, 99420, 99400, 99340, 99300, 99250, 99180, 99100, 99050, 
    99080, 99060, 99040, 99050, 99090, 99130, 99140, 99180, 99190, 99190, 
    99200, 99210, _, 99220, 99240, 99250, 99290, 99310, 99340, 99340, 99330, 
    99330, 99320, 99320, 99370, 99450, 99500, 99550, 99590, 99650, 99680, 
    99710, 99720, 99740, 99760, 99830, 99880, 99920, 99960, 99990, 100000, 
    100060, 100070, 100070, 100090, 100100, 100100, 100080, 100060, 100060, 
    100020, 99990, 99950, 99940, 99900, 99840, _, 99650, 99570, 99460, 99350, 
    99220, 99080, 98980, 98820, 98690, 98580, 98520, 98440, 98370, 98300, 
    98250, 98200, 98150, 98080, 98030, 97980, 97960, 97950, 97940, 97880, 
    97930, 97970, 98050, 98080, 98160, 98230, 98310, 98380, 98530, 98680, 
    98780, 98870, 98970, 99050, 99150, 99230, 99300, 99370, 99460, 99530, 
    99600, 99630, 99670, 99700, 99720, 99760, 99780, 99800, 99830, 99860, 
    99840, 99840, 99830, 99830, 99830, 99780, 99730, 99680, 99610, 99440, 
    99310, 99260, 99190, 99150, 99110, 99060, 99030, 99000, 98940, 98890, _, 
    98750, 98680, 98540, 98400, 98470, 98460, 98450, 98470, 98490, 98520, 
    98550, 98590, 98600, 98600, 98570, 98580, 98560, 98560, 98510, _, 98510, 
    98530, 98570, 98600, 98640, 98730, 98820, 98920, 99020, 99090, 99130, 
    99170, 99210, 99250, 99250, 99260, 99250, 99230, 99250, 99220, 99320, 
    99330, 99320, 99270, 99250, 99340, 99470, 99580, 99670, 99690, 99760, 
    99800, 99810, 99820, 99840, 99840, 99870, 99910, 99910, 99920, 99930, 
    99930, 99950, 99960, 100000, 100040, 100030, 100030, 100040, 100040, 
    100030, 100040, 100000, 99990, 100010, 100020, 100010, 100020, 100000, 
    99970, 99950, 99900, 99870, 99840, 99820, 99770, 99730, 99730, 99710, 
    99670, 99670, _, 99610, 99580, 99530, 99470, _, 99390, 99320, 99260, 
    99230, 99200, 99180, _, 99130, 99100, 99100, 99080, 99050, 99080, 99150, 
    99150, 99190, 99250, 99310, 99330, 99350, 99390, 99420, 99420, 99440, 
    99460, 99450, 99490, 99530, 99550, 99580, 99580, 99590, 99610, 99600, 
    99600, 99590, 99580, 99610, 99630, 99660, 99680, 99700, 99700, 99700, 
    99680, 99710, 99710, 99720, 99720, 99750, 99720, 99700, 99670, 99700, 
    99720, 99720, 99730, 99720, 99690, 99640, 99640, 99600, 99600, 99580, 
    99580, 99570, _, 99400, 99370, 99400, 99340, 99290, 99260, 99240, 99250, 
    99250, 99290, 99330, _, 99340, 99400, 99420, 99510, 99520, 99600, 99670, 
    99720, 99780, 99860, 99950, 100030, 100070, 100120, 100180, _, 100250, 
    100280, 100290, 100330, 100310, _, 100450, 100520, 100520, 100510, _, 
    100570, _, 100720, 100750, 100770, _, _, 100840, 100850, 100870, 100880, 
    100910, 100910, _, _, 100900, _, 100920, 100900, 100900, 100920, 100930, 
    _, 100960, 100940, 100950, 100930, 100930, 100910, 100910, 100880, 
    100860, 100820, _, 100790, 100770, 100770, _, 100640, _, _, 100450, 
    100390, 100340, 100260, 100150, _, 99980, 99880, 99770, 99680, _, _, _, 
    99270, 99190, 99110, 98990, 98870, 98820, 98810, 98790, 98790, 98770, 
    98780, 98760, 98740, 98710, 98640, 98580, 98450, 98340, 98340, 98400, 
    98380, 98290, 98240, 98200, 98220, 98250, 98290, 98290, 98290, 98320, 
    98300, 98260, 98240, 98230, 98070, 98070, 98260, 98360, 98330, 98370, 
    98380, 98430, 98420, 98430, 98430, 98470, 98470, 98480, 98560, 98530, 
    98590, 98550, 98540, 98600, 98490, _, 98650, 98620, 98630, 98630, 98630, 
    98630, 98730, 98860, 98850, 98830, 98850, 98740, 98670, 98660, 98660, 
    98670, 98680, 98700, 98730, 98750, 98720, 98780, 98790, 98760, 98680, 
    98690, 98780, _, 98990, 99070, 99060, 99090, 99140, 99200, 99250, 99290, 
    99340, 99430, 99480, 99520, 99580, 99590, 99620, 99660, 99710, 99750, 
    99820, 99890, 99940, 99990, 100070, 100160, 100240, 100280, 100340, 
    100400, 100490, 100560, 100590, 100650, 100690, 100720, 100760, 100800, 
    100840, 100900, 100910, 100970, 100950, 100950, 100970, _, 100960, 
    100940, 100950, 100950, 100960, 100950, _, 100920, 100900, 100880, 
    100840, 100810, 100780, 100790, 100780, 100760, 100730, 100700, 100700, 
    100660, 100630, 100590, 100560, 100570, 100530, 100490, 100450, 100410, 
    100400, 100370, 100320, 100270, 100260, 100210, 100170, 100100, 99990, 
    99960, 99910, 99840, 99760, 99660, 99530, 99450, 99370, 99240, 99180, 
    99110, 99060, 98990, 98980, 98940, 98900, 98870, 98880, 98890, 98880, 
    98880, 98900, 98910, 98930, 99000, 99070, 99170, 99230, 99290, 99320, 
    99320, 99320, 99330, 99330, 99330, 99360, 99370, 99380, 99400, 99400, 
    99400, _, 99400, 99420, 99430, 99420, 99430, 99410, 99410, 99420, 99460, 
    99480, 99490, 99500, 99500, 99490, 99510, 99520, 99530, 99550, 99510, 
    99530, 99530, 99510, 99490, 99470, 99470, 99480, 99440, 99420, 99410, 
    99370, 99330, 99290, 99300, 99330, 99330, 99330, 99280, 99210, 99210, 
    99180, 99160, 99160, 99130, 99150, 99160, 99190, 99220, 99240, 99260, 
    99270, 99310, 99340, 99370, 99390, 99400, 99430, 99470, 99520, 99530, 
    99510, 99580, 99610, 99620, 99650, 99670, 99730, 99740, 99770, 99830, 
    99880, 99880, 99940, 99890, 99880, 99910, 99880, 99800, 99820, 99800, 
    99810, 99840, 99870, 99940, 99990, 100000, 100130, 100170, 100290, 
    100400, 100450, 100510, 100570, 100610, 100660, 100730, 100800, 100850, 
    100920, 100970, 101060, 101120, 101210, 101320, 101430, 101470, 101450, 
    101460, 101550, 101550, 101580, 101650, 101770, 101860, 101910, 101890, 
    101930, 101960, 102010, 102100, 102100, 102120, 102080, 102160, 102180, 
    102190, 102170, 102170, 102170, 102190, 102210, 102180, 102170, 102180, 
    102160, 102150, 102120, 102100, 102070, 101980, 101900, 101930, 101840, 
    101720, 101750, 101700, 101630, 101480, 101380, 101370, 101240, 101190, 
    101160, 101130, 101080, 101030, 100980, 100810, 100720, 100720, 100700, 
    100560, 100500, 100400, 100430, 100360, 100270, 100110, 100020, 100000, 
    99910, 99820, 99750, 99750, 99700, 99660, 99680, 99680, 99560, 99460, 
    99420, 99310, 99250, 99200, 99160, 99120, 98980, 98910, 98850, 98810, 
    98780, 98750, 98630, 98590, 98420, 98490, 98450, 98460, 98390, 98340, 
    98260, 98100, 98070, 98100, 98080, 98070, 98010, 97910, 97810, 97760, 
    97720, 97670, 97620, 97550, 97500, 97410, 97360, 97370, 97320, 97220, 
    97120, 97220, 97150, 97120, 97060, 97050, 97060, 97000, 96980, 96870, 
    96860, 96890, 96890, 96930, 96920, _, 96930, _, _, _, 97040, _, _, 97220, 
    _, 97390, 97500, 97570, 97680, 97780, _, _, 98100, 98140, 98240, 98290, 
    98360, _, _, 98560, 98610, _, _, 98810, _, _, _, 99100, 99130, 99190, _, 
    99250, _, 99360, 99410, 99430, _, _, _, _, 99500, 99450, 99440, 99390, _, 
    99250, 99110, 98970, 98790, _, 98620, _, _, 98430, 98380, 98330, 98290, 
    98260, 98260, _, 98180, _, 98070, 98000, _, _, 97800, 97710, 97650, 
    97600, 97590, 97590, 97590, 97640, 97640, 97680, _, 97650, 97660, 97710, 
    97610, 97620, 97610, 97600, 97550, 97530, 97500, 97440, 97390, 97360, 
    97340, 97330, 97360, 97360, _, 97440, 97540, 97570, 97610, 97680, 97720, 
    97740, 97800, 97800, 97900, 97930, 97990, 98000, 98060, _, 97990, 97970, 
    97920, _, 97880, 97900, 97890, 97920, _, 97970, 97970, 98030, _, _, 
    98270, _, 98490, 98580, 98640, 98830, 99030, 99210, _, _, 99700, 99810, 
    99910, _, 100190, 100280, _, _, 100640, 100780, _, 100880, 100970, 
    101060, 101060, _, 101020, 100990, _, 100930, _, 100870, _, 100970, 
    101020, 101080, 101150, 101250, 101300, 101370, 101420, 101480, 101530, 
    101590, _, 101660, 101700, 101750, 101730, 101720, _, 101660, 101610, 
    101560, 101510, _, 101370, 101310, 101290, 101230, 101190, 101150, 
    101110, 101060, 101030, 100980, 100980, 100890, _, 100720, 100580, _, 
    100490, 100480, 100480, 100410, 100460, 100350, 100230, 100240, _, _, 
    100320, 100310, _, 100480, 100590, 100590, 100630, _, _, 100650, 100670, 
    100670, _, 100650, 100630, 100660, 100430, 100360, 100110, 100080, 
    100110, 100080, 100050, 100460, 100590, _, 100760, _, _, 100970, 101010, 
    101080, 101130, 101120, 101090, 101090, _, _, _, 100830, 100820, _, 
    100520, 100570, 100540, _, 100610, _, 100660, _, 100760, 100880, 100870, 
    100860, 100870, _, _, 100890, 100830, _, 100710, _, _, _, 100540, _, _, 
    _, 101250, 101440, _, 101810, _, _, 102110, 102170, 102180, 102170, 
    102140, 102140, 102100, 102010, _, 101870, 101790, 101690, _, _, 101500, 
    101430, _, _, 101320, _, 101310, _, _, 101300, _, 101310, 101300, 101270, 
    _, _, 101240, 101220, 101200, 101180, 101170, 101200, 101240, 101280, 
    101350, 101420, 101510, 101590, 101620, 101710, _, 101830, _, 101950, _, 
    102040, 102090, 102120, _, 102200, 102220, 102240, _, 102240, 102230, 
    102210, _, _, _, _, _, _, _, 102090, 102090, 102060, 102050, 102030, 
    102020, 101970, 101960, 101950, 101940, 101920, 101950, 101940, 101930, 
    101920, 101930, 101900, 101920, 101950, 101940, 101980, 102020, 102030, 
    102070, 102070, 102140, 102160, 102220, 102280, 102310, 102310, 102340, 
    102370, 102390, 102420, 102460, 102470, 102450, 102450, 102440, 102420, 
    102410, 102380, 102350, 102330, 102310, 102290, 102260, 102280, 102290, 
    102290, 102290, 102320, 102320, 102310, 102310, 102300, 102300, 102320, 
    102330, 102330, 102350, 102370, 102360, 102350, 102370, 102360, 102350, 
    102370, 102380, 102380, 102400, 102410, 102420, 102430, 102440, 102440, 
    102450, 102450, 102440, 102430, 102450, 102440, 102450, 102450, 102440, 
    102420, 102400, 102400, 102400, 102410, 102420, 102410, 102410, 102410, 
    102410, 102420, 102410, 102390, 102410, 102400, 102390, 102380, 102370, 
    102370, 102370, 102390, 102410, 102460, 102460, 102480, 102490, 102510, 
    102530, 102540, 102550, 102570, 102590, 102630, 102660, 102710, 102740, 
    102760, 102800, 102830, 102850, 102880, 102910, 102920, 102970, 103030, 
    103080, 103100, 103140, 103170, 103230, 103250, 103270, 103310, 103330, 
    103340, 103380, 103420, 103450, 103480, 103490, 103490, 103500, 103510, 
    103510, 103500, 103490, 103490, 103460, 103450, 103430, 103380, 103350, 
    103300, 103220, 103190, 103150, 103090, 102990, 102900, 102760, 102640, 
    102550, 102440, 102320, 102190, 102040, 101940, 101820, 101720, 101640, 
    101580, 101540, 101530, 101530, 101530, 101500, 101490, 101440, 101390, 
    101360, 101310, 101260, 101210, 101130, 101080, 101010, 100970, 100910, 
    100900, 100900, 100900, 100890, 100870, 100870, 100840, 100810, 100810, 
    100850, 100910, 100920, 100900, 100900, 100910, 100940, 100990, 101010, 
    101030, 101060, 101070, 101090, 101130, 101150, 101120, 101030, 101010, 
    101050, 101140, 101230, 101310, 101430, 101530, 101630, 101730, 101800, 
    101840, 101870, 101930, 101990, 102020, 102060, 102070, 102090, 102130, 
    102170, 102180, 102200, 102240, 102240, 102230, 102180, 102230, 102260, 
    102280, 102340, 102370, 102390, 102420, 102460, 102450, 102450, 102490, 
    102500, 102520, 102540, 102540, 102520, 102500, 102490, 102480, 102460, 
    102430, 102400, 102400, 102420, 102420, 102380, 102380, 102340, 102230, 
    102280, 102310, 102250, 102230, 102190, 102180, 102110, 102070, 102080, 
    102080, 102080, 102070, 102050, 102000, 102070, 102040, 102020, 101930, 
    101910, 101900, 101880, 101840, 101810, 101790, 101780, 101810, 101840, 
    101870, 101870, 101850, 101860, 101860, 101870, 101860, 101830, 101830, 
    101840, 101840, 101830, 101790, 101780, 101750, 101720, 101700, 101680, 
    101660, 101650, 101630, 101600, 101570, 101540, 101490, 101440, 101400, 
    101370, 101330, 101290, 101250, 101230, 101180, 101160, 101120, 101090, 
    101050, 101030, 100980, 100950, 100910, 100890, 100870, 100840, 100810, 
    100800, 100810, 100800, 100780, 100750, 100720, 100710, 100690, 100660, 
    100650, 100640, 100640, 100640, 100640, 100640, 100660, 100650, 100670, 
    100680, 100660, 100680, 100670, 100650, 100660, 100660, 100660, 100640, 
    100570, 100480, 100400, 100310, 100310, 100350, 100350, 100360, 100350, 
    100330, 100350, 100340, 100310, 100270, 100240, 100200, 100180, 100140, 
    100110, 100060, 100010, 99990, 99950, 99940, 99940, 99960, 99990, 100020, 
    100060, 100110, 100150, 100190, 100200, 100260, 100300, 100300, 100310, 
    100310, 100270, 100270, 100270, 100280, 100290, 100270, 100350, 100410, 
    100490, 100510, 100560, 100650, 100670, 100720, 100740, 100820, 100840, 
    100840, 100880, 100950, 100990, 101000, 101010, 101030, 101070, 101080, 
    101110, 101130, 101130, 101160, 101200, 101210, 101260, 101280, 101310, 
    101310, 101310, 101350, 101370, 101390, 101400, 101460, 101470, 101500, 
    101560, 101620, 101600, 101570, 101600, 101620, 101580, 101610, 101640, 
    101640, 101630, 101670, 101680, 101690, 101750, 101740, 101740, 101780, 
    101780, 101800, 101840, 101840, 101840, 101870, 101860, 101860, 101860, 
    101820, 101770, 101730, 101680, 101640, 101590, 101500, 101480, 101420, 
    101370, 101320, 101290, 101250, 101190, 101140, 101070, 100980, 100890, 
    100800, 100700, 100640, 100530, 100460, 100380, 100260, 100150, 100020, 
    99890, 99750, 99630, 99610, 99570, 99530, 99490, 99450, 99410, 99380, 
    99330, 99370, 99340, 99290, 99230, 99220, 99190, 99180, 99190, 99160, 
    99140, 99130, 99110, 99130, 99120, 99070, 99020, 98980, 98950, 98950, 
    98970, 98960, 98910, 98870, 98790, 98780, 98750, 98640, 98590, 98530, 
    98520, 98360, 98470, 98280, 98150, 98010, 97970, 97910, 97910, 97910, 
    97890, 97930, 97970, 98010, 98070, 98100, 98110, 98170, 98230, 98290, 
    98330, 98380, 98380, 98400, 98420, 98480, 98590, 98620, 98670, 98690, 
    98680, 98720, 98770, 98810, 98860, 98940, 98990, 99040, 99000, 98990, 
    98990, 99020, 98980, 98960, 98990, 98990, 99080, 99170, 99200, 99240, 
    99270, 99280, 99230, 99160, 99120, 99100, 99050, 98990, 99010, 98990, 
    99000, 99050, 98970, 98960, 99010, 99090, 99130, 99200, 99190, 99230, 
    99230, 99240, 99270, 99290, 99250, 99200, 99310, 99460, 99530, 99490, 
    99420, 99400, 99350, 99380, 99490, 99540, 99630, 99650, 99670, 99700, 
    99720, 99750, 99780, 99800, 99790, 99810, 99740, 99760, 99800, 99800, 
    99790, 99830, 99880, 99870, 99910, 99890, 99930, 99600, 99560, 99670, 
    99860, 100080, 100110, 100130, 100170, 100170, 100190, 100190, 100170, 
    100150, 100170, 100200, 100250, 100320, 100370, 100380, 100400, 100370, 
    100430, 100510, 100580, 100540, 100630, 100680, 100700, 100730, 100700, 
    100560, 100630, 100750, 100760, 100800, 100730, 100700, 100680, 101080, 
    101390, 101420, 101450, 101470, 101470, 101410, 101460, 101380, 101520, 
    101550, 101490, 101470, 101500, 101550, 101510, 101460, 101440, 101380, 
    101350, 101320, 101220, 101240, 101210, 101180, 101160, 101140, 101100, 
    101070, 101020, 100970, 100940, 100870, 100800, 100740, 100760, 100760, 
    _, 100730, 100720, 100700, 100670, 100690, 100680, 100700, 100700, 
    100690, 100660, 100660, 100640, 100620, 100610, 100610, 100590, 100580, 
    100540, 100500, 100490, 100470, 100460, 100480, 100460, 100480, 100490, 
    100470, 100460, 100450, 100420, 100410, 100410, _, 100370, 100380, 
    100390, 100410, 100430, 100460, 100470, 100480, 100490, 100480, 100490, 
    100500, 100510, 100530, 100570, 100590, 100600, 100610, _, 100610, 
    100590, 100580, 100590, 100600, 100610, 100630, 100640, 100620, 100600, 
    100580, 100550, 100540, 100500, 100470, 100450, 100410, 100370, 100350, 
    100320, 100270, 100190, 100140, 100020, 99970, 99920, 99840, 99740, 
    99690, 99540, _, 99370, 99150, 99070, 99020, 98960, 98800, 98840, 98780, 
    98750, _, 98630, 98560, 98460, 98330, 98210, 98180, 98100, 97980, 97880, 
    97790, 97720, 97670, 97680, 97620, 97600, 97550, 97520, 97470, 97500, 
    97490, 97440, 97440, 97380, 97400, 97430, 97460, 97500, 97550, 97590, 
    97610, 97630, 97710, 97790, 97880, 97960, 98050, 98160, 98230, 98320, 
    98380, 98450, 98500, 98570, 98600, 98620, 98640, 98670, 98710, 98780, 
    98840, 98880, 98940, 98970, 99000, 99030, 99060, 99090, 99140, 99180, 
    99230, 99280, 99320, 99370, 99420, 99470, 99510, 99550, 99610, 99640, 
    99670, 99720, 99760, 99820, 99880, 99940, 99960, 99990, 100020, 100040, 
    100070, 100100, 100130, 100130, 100140, 100140, 100170, 100190, 100200, 
    100210, 100210, 100200, 100190, 100180, 100180, 100170, 100180, 100190, 
    100210, 100220, 100220, 100200, 100210, 100230, 100290, 100340, 100380, 
    100480, 100520, 100580, 100630, 100700, 100770, 100840, 100900, 100930, 
    100960, 100990, 101030, 101070, 101110, 101150, 101180, 101280, 101290, 
    101330, 101390, 101450, 101500, 101540, 101570, 101620, 101660, 101710, 
    101750, 101800, 101800, 101800, 101770, 101770, 101780, 101780, 101740, 
    101700, 101680, 101670, 101690, 101690, 101700, 101680, 101630, 101610, 
    101600, 101570, 101540, 101520, 101520, 101540, 101550, 101520, 101460, 
    101460, 101450, 101430, 101400, 101390, 101350, 101370, 101340, 101330, 
    101290, 101260, 101250, 101230, 101220, 101230, 101220, 101200, 101160, 
    101160, 101130, 101150, 101150, 101130, 101130, 101080, 101060, 101080, 
    101070, 101060, 101020, 101020, 100980, 100930, 100880, 100870, 100890, 
    100890, 100810, 100760, 100730, 100680, 100630, 100580, 100500, 100430, 
    100390, 100360, 100350, 100350, 100360, 100410, 100430, 100460, 100510, 
    100540, 100590, 100620, 100660, 100680, 100690, 100690, 100710, 100700, 
    100710, 100690, 100690, 100650, 100680, 100590, 100620, 100650, 100600, 
    100570, 100510, 100470, 100420, 100370, 100330, 100280, 100180, 100110, 
    100070, 100000, 99870, 99770, 99630, 99540, 99440, 99380, 99330, 99250, 
    99190, 99160, 99170, 99210, 99210, 99210, 99210, 99240, _, 99280, 99290, 
    99280, 99280, 99290, 99300, 99320, 99340, 99370, 99390, 99430, 99440, 
    99450, 99430, 99450, 99470, 99520, 99560, 99620, 99680, 99710, 99720, 
    99760, 99810, 99880, 99940, 100030, 100070, 100160, 100240, 100320, 
    100400, 100460, 100510, 100540, 100550, 100570, 100550, 100520, 100530, 
    100500, 100490, 100420, 100370, 100310, 100260, 100230, 100180, 100110, 
    100090, 100110, 100130, 100150, 100190, 100240, 100290, 100310, 100350, 
    100360, 100400, 100430, 100500, 100540, 100590, 100630, 100680, 100730, 
    100760, 100790, 100830, 100870, _, 100930, 100960, 100980, 101000, 
    101000, 101010, 101070, 101100, 101070, 101100, _, 101110, 101140, 
    101140, 101160, 101190, 101250, 101320, 101390, 101440, 101470, 101480, 
    101530, 101560, 101590, 101630, 101640, 101650, 101660, 101680, 101700, 
    101700, 101690, 101680, 101670, 101650, 101650, 101650, 101640, 101640, 
    101620, 101570, 101600, 101620, 101630, 101600, 101590, 101580, 101580, 
    101540, 101530, 101530, 101560, 101550, 101570, 101550, 101550, 101530, 
    101530, 101530, 101530, 101550, 101560, 101580, 101560, 101570, 101550, 
    101560, 101560, 101530, 101530, 101520, 101520, 101500, 101520, 101530, 
    101540, 101530, 101540, 101560, 101560, 101540, 101520, 101510, 101490, 
    101490, 101460, 101450, 101440, 101420, 101410, 101390, 101360, 101330, 
    101290, 101250, 101240, 101210, 101180, 101160, 101130, 101120, 101100, 
    101080, 101050, 101040, 101000, 100980, 100950, 100920, 100880, 100880, 
    100870, 100850, 100840, 100810, 100820, 100800, 100770, 100750, 100760, 
    100760, 100740, 100730, 100730, 100740, 100750, 100770, 100770, 100760, 
    100770, 100770, 100770, 100760, 100750, 100740, 100740, 100710, 100730, 
    100740, 100720, 100720, 100710, 100680, 100680, 100680, 100710, 100720, 
    100720, 100750, 100760, 100760, 100780, 100760, 100760, 100750, 100750, 
    100760, 100730, 100720, 100740, 100690, 100680, 100690, 100670, 100660, 
    100640, 100630, 100620, 100620, 100640, 100650, 100660, 100640, 100660, 
    100640, 100610, 100590, 100550, 100490, 100400, 100420, 100430, 100380, 
    100420, 100470, 100480, 100420, 100450, 100510, 100510, 100490, 100470, 
    100410, 100350, 100220, 100180, 100230, 100280, 100280, 100300, 100310, 
    100310, 100320, 100380, 100430, 100500, 100540, 100610, 100680, 100710, 
    100740, 100770, 100780, 100770, 100740, 100780, 100770, 100750, 100730, 
    100740, 100730, 100740, 100750, 100800, 100800, 100780, 100790, 100780, 
    100770, 100750, 100710, 100710, 100700, 100710, 100760, 100790, 100830, 
    100830, 100830, 100830, 100830, 100820, 100810, 100800, 100800, 100770, 
    100810, 100800, 100780, 100750, 100720, 100660, 100640, 100610, 100560, 
    100510, 100450, 100410, 100360, 100280, 100200, 100140, 100060, 100010, 
    99980, 99970, 99970, 99960, 100020, 100090, 100140, 100160, 100170, 
    100120, 100120, 100080, 100080, 100070, 100070, 100080, 100130, 100180, 
    100230, 100290, 100340, 100380, 100450, 100470, 100510, 100550, 100590, 
    100580, 100620, 100650, 100690, 100700, 100700, 100700, 100690, 100700, 
    100710, 100720, 100740, 100750, 100770, 100810, 100850, 100880, 100950, 
    100990, 101010, 101070, 101100, 101140, 101160, 101170, 101210, 101210, 
    101230, 101230, 101240, 101240, 101230, 101240, 101240, 101250, 101250, 
    101280, 101280, 101290, 101260, 101280, 101300, 101270, 101260, 101260, 
    101300, 101330, 101360, 101370, 101400, 101450, 101470, 101510, 101510, 
    101530, 101550, 101590, 101610, 101640, 101690, 101700, 101670, 101660, 
    101680, 101760, 101800, 101810, 101810, 101820, 101830, 101840, 101850, 
    101870, 101870, 101880, 101860, 101840, 101840, 101790, 101720, 101650, 
    101610, 101570, 101550, 101520, 101480, 101440, 101380, 101340, 101310, 
    101290, 101230, 101180, 101180, 101170, 101130, 101100, 101110, 101110, 
    101100, 101110, 101130, 101160, 101150, 101160, 101150, 101170, 101200, 
    101210, 101230, 101250, 101260, 101250, 101280, 101290, 101290, 101330, 
    101320, 101340, 101350, 101340, 101330, 101290, 101280, 101240, 101220, 
    101190, 101160, 101090, 101050, 101000, 100930, 100910, 100850, 100810, 
    100780, 100720, 100710, 100670, 100650, 100580, 100510, 100450, 100390, 
    100450, 100420, 100430, 100450, 100470, 100510, 100490, 100500, 100540, 
    100530, 100560, 100540, 100540, 100550, 100570, 100530, 100500, 100480, 
    100420, 100360, 100330, 100270, 100220, 100140, 100070, 99950, 99880, 
    99700, 99510, 99370, 99210, 99060, 98980, 98920, 98930, 98910, 98940, 
    98960, 98990, 98980, 99040, 99040, 99130, 99170, 99330, 99550, 99620, 
    99760, 99900, 100040, 100180, 100210, 100240, 100330, 100290, 100230, 
    100180, 100090, 99990, 99880, 99670, 99460, 99210, 98980, 98810, 98570, 
    98450, 98360, 98350, 98350, 98470, 98520, 98620, 98780, 98890, 98990, 
    99130, 99240, 99400, 99540, 99580, 99670, 99730, 99790, 99870, 99950, 
    99990, 100040, 100000, 100060, 100100, 100140, 100140, 100110, 100110, 
    100110, 100110, 100110, 100090, 100110, 100090, 100070, 100060, 100050, 
    100050, 100090, 100110, 100110, 100140, 100210, 100250, 100300, 100350, 
    100400, 100470, 100540, 100600, 100640, 100670, 100730, 100790, 100830, 
    100850, 100890, 100930, 100970, 101010, 101050, 101060, 101030, 101010, 
    101050, 100960, 100910, 100930, 100870, 100800, 100780, 100780, 100750, 
    100830, 100840, 100840, 100830, 100850, 100850, 100890, 100890, 100930, 
    100930, 100890, 100910, 100940, 100910, 100850, 100850, 100840, 100890, 
    100900, 100890, 100840, 100810, 100780, 100750, 100710, 100680, 100660, 
    100610, 100590, 100590, 100620, 100650, 100660, 100650, 100650, 100680, 
    100650, 100670, 100690, 100720, 100740, 100740, 100780, 100810, 100830, 
    100810, 100780, 100790, 100790, 100820, 100840, 100820, 100780, 100800, 
    100790, 100820, 100820, 100820, 100810, 100810, 100790, 100800, 100760, 
    100750, 100730, 100720, 100710, 100620, 100540, 100500, 100510, 100520, 
    100470, 100410, 100390, 100380, 100320, 100300, 100320, 100320, 100310, 
    100310, 100290, 100280, 100300, 100260, 100250, 100250, 100240, 100230, 
    100250, 100240, 100230, 100230, 100230, 100220, 100240, 100230, 100240, 
    100240, 100250, 100270, 100320, 100350, 100370, 100360, 100400, 100420, 
    100470, 100510, 100530, 100560, 100580, 100590, 100630, 100650, 100660, 
    100670, 100670, 100700, 100690, 100720, 100730, 100730, 100730, 100730, 
    100730, 100740, 100760, 100760, 100770, 100780, 100800, 100810, 100820, 
    100830, 100830, 100850, 100850, 100860, 100860, 100870, 100860, 100870, 
    100870, 100870, 100880, 100870, 100870, 100880, 100900, 100920, 100920, 
    100910, 100920, 100910, 100920, 100930, 100920, 100910, 100880, 100890, 
    100880, 100860, 100850, 100830, 100790, 100720, 100660, 100550, 100520, 
    100500, 100500, 100500, 100500, 100490, 100490, 100480, 100450, 100420, 
    100390, 100340, 100320, 100310, 100350, 100340, 100380, 100400, 100410, 
    100410, 100450, 100470, 100490, 100500, 100520, 100520, 100510, 100540, 
    100550, 100580, 100580, 100560, 100530, 100520, 100510, 100490, 100470, 
    100450, 100410, 100400, 100400, 100370, 100380, 100360, 100340, 100330, 
    100330, 100290, 100240, 100200, 100150, 100120, 100110, 100050, 99970, 
    99910, 99860, 99770, 99710, 99640, 99550, 99460, 99370, 99280, 99220, 
    99180, 99050, 98910, 98770, 98560, 98430, 98380, 98390, 98350, 98350, 
    98300, 98250, 98190, 98120, 98090, 98040, 98000, 97990, 98020, 98050, 
    98060, 97950, 97970, 98100, 98280, 98270, 98420, 98430, 98390, 98420, 
    98450, 98500, 98540, 98600, 98610, 98700, 98790, 98810, 98830, 98910, 
    99090, 99170, 99220, 99270, 99320, 99360, 99380, 99380, 99430, 99430, 
    99430, 99430, 99410, 99390, 99390, 99390, 99400, 99430, 99430, 99450, 
    99440, 99460, 99460, 99440, 99450, 99460, 99460, 99460, 99480, 99490, 
    99470, 99470, 99480, 99510, 99530, 99530, 99530, 99560, 99580, 99610, 
    99620, 99660, 99700, 99720, 99750, 99810, 99830, 99870, 99920, 99930, 
    99930, 99980, 100030, 100080, 100100, 100110, 100170, 100210, 100280, 
    100330, 100370, 100400, 100420, 100470, 100530, 100580, 100650, 100720, 
    100780, 100840, 100920, 100960, 101020, 101040, 101090, 101120, 101150, 
    101200, 101240, 101290, 101350, 101380, 101410, 101430, 101450, 101460, 
    101490, 101530, 101560, 101570, 101580, 101600, 101600, 101630, 101630, 
    101620, 101630, 101630, 101630, 101630, 101610, 101630, 101630, 101630, 
    101620, 101640, 101600, 101610, 101590, 101600, 101580, 101550, 101540, 
    101540, 101560, 101590, 101600, 101610, 101610, 101610, 101580, 101580, 
    101570, 101600, 101620, 101630, 101650, 101680, 101700, 101700, 101720, 
    101720, 101730, 101720, 101740, 101760, 101770, 101760, 101820, 101860, 
    101880, 101890, 101880, 101890, 101890, 101890, 101900, 101920, 101930, 
    101960, 101980, 102010, 102010, 102000, 101970, 101950, 101950, 101930, 
    101930, 101920, 101880, 101870, 101870, 101880, 101870, 101830, 101820, 
    101800, 101760, 101730, 101710, 101700, 101660, 101640, 101610, 101590, 
    101580, 101570, 101540, 101500, 101490, 101460, 101460, 101460, 101460, 
    101450, 101460, 101470, 101490, 101490, 101500, 101520, 101560, 101550, 
    101580, 101590, 101630, 101630, 101620, 101620, 101620, 101610, 101600, 
    101630, 101640, 101650, 101670, 101670, 101690, 101720, 101740, 101760, 
    101750, 101760, 101780, 101780, 101770, 101780, 101820, 101830, 101860, 
    101870, 101880, 101910, 101930, 101940, 101940, 101930, 101940, 101950, 
    101940, 101940, 101930, 101920, 101920, 101920, 101900, 101880, 101810, 
    101800, 101770, 101780, 101780, 101760, 101740, 101720, 101700, 101680, 
    101680, 101640, 101580, 101570, 101550, 101510, 101480, 101450, 101450, 
    101420, 101390, 101360, 101360, 101330, 101280, 101250, 101220, 101220, 
    101210, 101180, 101140, 101120, 101140, 101180, 101200, 101240, 101250, 
    101300, 101340, 101400, 101420, 101430, 101450, 101470, 101470, 101460, 
    101420, 101380, 101350, 101330, 101340, 101360, 101370, 101370, 101370, 
    101360, 101380, 101400, 101360, 101350, 101340, 101300, 101290, 101210, 
    101150, 101060, 101030, 101020, 100960, 100990, 100940, 100940, 100970, 
    101010, 101050, 101080, 101090, 101080, 101080, 101110, 101120, 101160, 
    101220, 101200, 101220, 101220, 101230, 101230, 101250, 101230, 101270, 
    101320, 101330, 101360, 101370, 101380, 101390, 101430, 101410, 101370, 
    101320, 101260, 101330, 101320, 101310, 101280, 101240, 101250, 101170, 
    101140, 101110, 101050, 100980, 100940, 100890, 100900, 100880, 100880, 
    100910, 100880, 100890, 100890, 100870, 100850, 100800, 100770, 100780, 
    100740, 100680, 100640, 100700, 100730, 100690, 100660, 100680, 100660, 
    100720, 100720, 100820, 100850, 100870, 100870, 100900, 100910, 100920, 
    100980, 100950, 100970, 100980, 100980, 101060, 101100, 101050, 101040, 
    101090, 101080, 101060, 101100, 101080, 101080, 101070, 101070, 101080, 
    101100, 101100, 101150, 101170, 101130, 101110, 101120, 101090, 101080, 
    101100, 101100, 101220, 101200, 101220, 101210, 101210, 101170, 101230, 
    101290, 101290, 101270, 101290, 101320, 101310, 101340, 101350, 101370, 
    101380, 101400, 101410, 101430, 101440, 101460, 101460, 101470, 101480, 
    101510, 101530, 101530, 101530, 101520, 101500, 101500, 101500, 101480, 
    101460, 101470, 101460, 101460, 101450, 101440, 101430, 101430, 101410, 
    101400, 101390, 101380, 101350, 101340, 101330, 101300, 101280, 101260, 
    101240, 101230, 101230, 101200, 101160, 101140, 101110, 101080, 101060, 
    101020, 100990, 100920, 100840, 100780, 100670, 100610, 100540, 100450, 
    100380, 100320, 100260, 100140, 100090, 100030, 99990, 99910, 99860, 
    99820, 99740, 99640, 99600, 99610, 99590, 99590, 99590, 99600, 99610, 
    99620, 99630, 99650, 99650, 99650, 99680, 99700, 99710, 99730, 99750, 
    99770, 99780, 99800, 99830, 99850, 99880, 99890, 99920, 99960, 100010, 
    100030, 100060, 100090, 100170, 100230, 100260, 100370, 100490, 100530, 
    100610, 100660, 100700, 100740, 100780, 100810, 100860, 100910, 100980, 
    101070, 101110, 101150, 101210, 101240, 101320, 101390, 101460, 101530, 
    101600, 101670, 101750, 101790, 101860, 101880, 101910, 101950, 101990, 
    102020, 102060, 102100, 102130, 102140, 102110, 102120, 102120, 102120, 
    102090, 102080, 102090, 102050, 102050, 102010, 101940, 101900, 101870, 
    101820, 101810, 101810, 101810, 101760, 101750, 101740, 101720, _, 
    101720, 101730, 101720, 101700, 101690, 101640, 101610, 101570, 101560, 
    101540, _, 101460, 101420, _, 101340, 101290, 101240, 101240, 101200, 
    101170, 101110, 101100, 101110, 101090, 101070, 101110, 101150, 101160, 
    101180, 101200, 101220, 101250, 101310, 101380, 101450, 101500, 101570, 
    101630, 101670, 101710, 101760, 101780, 101820, 101840, 101870, 101900, 
    101940, 101960, 101980, 101980, 101930, 101960, 102020, 102040, 101990, 
    102000, 102010, 102060, 102120, 102170, 102240, 102290, 102390, 102430, 
    102480, 102570, 102650, 102740, 102860, 102990, 103110, _, 103280, 
    103350, 103440, 103500, 103590, 103660, 103730, 103810, 103850, 103920, 
    _, 103980, 104010, 104060, 104090, 104090, 104080, 104100, 104120, 
    104140, 104140, 104180, 104160, 104130, 104110, 104080, 104030, 104020, 
    103990, 103930, 103900, 103820, 103860, 103750, 103810, 103780, 103760, 
    103760, 103750, 103730, 103720, 103700, 103680, 103680, 103650, 103630, 
    _, 103600, 103590, 103560, 103530, 103470, 103400, 103350, 103300, 
    103260, 103230, 103200, 103170, 103120, 103080, 103060, 103020, 102970, 
    102990, 102980, 102970, 102980, 103000, 103010, 103040, _, 103140, 
    103160, 103190, 103230, 103240, 103280, 103280, 103330, 103360, 103390, 
    103430, 103460, 103490, 103500, 103490, 103500, 103510, 103470, 103450, 
    103400, 103380, 103340, 103300, _, 103250, 103240, 103270, 103260, 
    103240, 103240, 103220, 103230, 103210, 103190, 103190, 103180, 103150, 
    103110, 103100, 103070, 103030, 102970, 102920, 102840, 102770, 102700, 
    102650, 102550, 102450, 102340, 102270, 102190, 102140, 102040, 101930, 
    101890, 101850, 101840, 101760, 101730, 101700, 101650, 101620, 101610, 
    101620, 101640, 101620, 101640, 101650, 101650, 101680, 101680, 101720, 
    101710, 101730, 101800, 101840, 101850, 101890, 101890, 101950, 101960, 
    102020, 102080, 102100, 102130, 102180, 102210, 102250, 102270, 102310, 
    102320, 102350, 102380, 102420, 102470, 102510, 102540, 102560, 102580, 
    102600, 102610, 102610, 102630, 102650, 102690, 102730, 102750, 102760, 
    102790, 102810, 102830, 102830, 102840, 102830, 102840, 102840, 102850, 
    102870, 102890, 102890, 102900, 102910, 102890, 102890, 102880, 102890, 
    102870, 102860, 102870, 102880, 102890, 102900, 102890, 102900, 102890, 
    102900, 102890, 102860, 102860, 102890, 102850, 102850, 102850, 102860, 
    102870, 102860, 102860, 102850, 102840, 102840, 102850, 102860, 102880, 
    102900, 102910, 102920, 102920, 102930, 102930, 102910, 102900, 102910, 
    102900, 102880, 102860, 102860, _, 102840, 102850, 102850, 102800, 
    102780, 102750, 102730, 102710, 102690, 102680, 102690, 102690, 102690, 
    102660, 102620, 102610, 102600, 102560, 102560, 102550, 102520, 102530, 
    102480, 102470, 102490, 102460, 102430, 102400, 102380, 102380, 102370, 
    102340, 102300, 102290, 102280, 102300, 102340, 102330, 102320, 102310, 
    102220, 102190, 102180, 102170, 102150, 102170, 102130, 102120, 102100, 
    102060, 102040, 102010, 101990, 101970, 101960, 101980, 101980, 102040, 
    102070, _, 102140, 102050, 102070, 102090, 102100, 102100, 102100, 
    102180, 102160, 102100, 102120, 102180, 102210, 102190, 102190, 102180, 
    102180, 102180, 102180, 102200, 102210, 102210, 102230, 102200, 102230, 
    102230, 102240, 102240, 102240, 102230, 102220, 102210, 102170, 102160, 
    102140, 102120, 102110, 102120, 102120, 102110, 102100, 102090, 102100, 
    102100, 102090, 102100, 102110, 102130, 102130, 102160, 102150, 102150, 
    102170, 102150, 102160, 102150, 102140, 102150, 102150, 102150, 102160, 
    102170, 102170, 102180, 102180, 102180, 102180, 102180, 102200, 102200, 
    102190, 102180, 102200, 102210, 102220, 102190, 102140, 102140, 102130, 
    102090, 102030, 102030, 102020, 101970, 101930, 101900, 101830, 101810, 
    101780, 101750, 101700, 101640, 101650, 101650, 101670, 101690, 101710, 
    101720, 101790, 101810, 101840, 101890, 101950, 101970, 102000, 102000, 
    102000, 102030, 102060, 102090, 102110, 102110, 102130, 102160, 102180, 
    102160, 102150, 102170, 102190, 102190, 102170, 102180, 102160, 102170, 
    102150, 102130, 102110, 102110, 102080, 102080, 102040, 102040, 101990, 
    101960, 101930, 101930, 101880, 101860, 101820, 101770, 101740, 101690, 
    101660, 101630, 101620, 101590, 101540, 101530, 101460, 101400, 101350, 
    101300, 101230, 101150, 101060, 100980, 100950, 100860, 100750, 100620, 
    100590, 100550, 100540, 100550, 100540, 100540, 100500, 100510, 100540, 
    100580, 100580, 100570, 100570, 100540, 100560, 100530, 100540, 100550, 
    100540, 100580, 100590, 100570, 100520, 100500, 100510, 100460, 100400, 
    100370, 100350, 100310, 100210, 100180, 100250, 100170, 100130, 100080, 
    100130, 100120, 100150, 100200, 100200, 100180, 100170, 100190, 100200, 
    100210, 100210, 100210, 100220, 100220, 100230, 100250, 100270, 100290, 
    100320, 100330, 100350, 100370, 100350, 100350, 100350, 100360, 100350, 
    100360, 100340, 100330, 100330, 100300, 100290, 100270, 100260, 100240, 
    100200, 100170, 100150, 100110, 100090, 100080, 100060, 100050, 100040, 
    100010, 99980, 99960, 99930, 99910, 99890, 99870, 99840, 99830, 99800, 
    99790, 99770, 99760, 99750, 99740, 99730, 99720, 99740, 99720, 99730, 
    99740, 99760, 99790, 99820, 99840, 99850, 99880, 99900, 99920, 99960, 
    99960, 100000, 100030, 100060, 100100, 100150, 100180, 100200, 100220, 
    100250, 100260, 100280, 100320, 100330, 100370, 100400, 100420, 100450, 
    100470, 100460, 100470, 100490, 100520, 100550, 100580, 100570, 100570, 
    100570, 100560, 100630, 100700, 100730, 100790, 100880, 100930, 101020, 
    101120, 101140, 101220, 101300, 101360, 101420, 101490, 101530, 101560, 
    101590, 101610, 101650, 101640, 101650, 101670, 101680, 101700, 101730, 
    101760, 101800, 101840, 101860, 101890, 101900, 101930, 101960, 101990, 
    102030, 102040, 102080, 102110, 102120, 102120, 102130, 102130, 102120, 
    102110, 102110, 102090, 102100, 102090, 102080, 102090, 102060, 102040, 
    102010, 101970, 101940, 101920, 101910, 101900, 101900, 101900, 101900, 
    101890, 101890, 101920, 101890, 101880, 101860, 101860, 101840, 101880, 
    101900, 101870, 101840, 101790, 101740, 101730, 101750, 101750, 101700, 
    101800, 101810, 101810, 101790, 101760, 101720, 101620, 101560, 101470, 
    101540, 101490, 101480, 101530, 101590, 101550, 101560, 101600, 101650, 
    101620, 101620, 101590, 101620, 101670, 101640, 101640, 101640, 101590, 
    101600, 101580, 101570, 101580, 101560, 101570, 101580, 101580, 101610, 
    101600, 101630, 101640, 101650, 101620, 101620, 101630, 101620, 101650, 
    101660, 101690, 101680, 101690, 101710, 101740, 101750, 101760, 101770, 
    101780, 101800, 101820, 101810, 101830, 101820, 101800, 101810, 101790, 
    101790, 101810, 101800, 101790, 101760, 101760, 101760, 101770, 101700, 
    101730, 101700, 101660, 101610, 101570, 101520, 101430, 101390, 101290, 
    101230, 101120, 101010, 100940, 100840, 100760, 100730, 100690, 100720, 
    100640, 100600, 100550, 100520, 100460, 100450, 100380, 100360, 100350, 
    100400, 100450, 100480, 100530, 100580, 100640, 100700, 100780, 100870, 
    100990, 101110, 101190, 101310, 101440, 101600, 101770, 101950, 102080, 
    102210, 102340, 102440, 102540, 102650, 102760, 102860, 102930, 102990, 
    103090, 103130, 103180, 103250, 103300, 103310, 103330, 103360, 103380, 
    103380, 103390, 103400, 103410, 103380, 103380, 103350, 103320, 103300, 
    103260, 103230, 103210, 103190, 103180, 103180, 103140, 103130, 103110, 
    103060, 103010, 102960, 102910, 102870, 102820, 102780, 102730, 102680, 
    102630, 102610, 102550, 102480, 102420, 102360, 102320, 102250, 102190, 
    102120, 102070, 102020, 101980, 101940, 101890, 101840, 101780, 101720, 
    101700, 101650, 101590, 101580, 101550, 101540, 101490, 101470, 101450, 
    101440, 101420, 101430, 101510, 101560, 101650, 101700, 101760, 101880, 
    101950, 102010, 102070, 102070, 102100, 102130, 102130, 102120, 102100, 
    102100, 102090, 102080, 102050, 102030, 102000, 101930, 101860, 101780, 
    101730, 101670, 101610, 101540, 101490, 101420, 101370, 101320, 101270, 
    101230, 101200, 101120, 101080, 101040, 100990, 100930, 100870, 100800, 
    100800, 100830, 100800, 100830, 100830, 100810, 100810, 100860, 100880, 
    100920, 100940, 100950, 100970, 100970, 100990, 100990, 101000, 100970, 
    100950, 100990, 100960, 100970, 100990, 101020, 101030, 101040, 101020, 
    101050, 101030, 101040, 101030, 100980, 100940, 100990, 101090, 101130, 
    101170, 101260, 101320, 101360, 101390, 101440, 101430, 101480, 101530, 
    101630, 101700, 101710, 101720, 101780, 101810, 101820, 101840, 101860, 
    101890, 101910, 101900, 101920, 101980, 102000, 102020, 102050, 102060, 
    102050, 102050, 102030, 102050, 102040, 102010, 102030, 101990, 101980, 
    101960, 101960, 101930, 101910, 101900, 101870, 101820, 101800, 101790, 
    101740, 101720, 101690, 101650, 101600, 101540, 101490, 101470, 101410, 
    101340, 101300, 101260, 101220, 101200, 101140, 101100, 101060, 101020, 
    100990, 100960, 101030, 100920, 100930, 100930, 100940, 100930, 100940, 
    100940, 100970, 100970, 100940, 100930, 100920, 100960, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 101160, 101160, 101140, 101150, 101160, 
    101180, 101230, 101230, 101250, 101240, 101220, 101200, 101160, 101100, 
    101070, 101030, 101000, 100950, 100910, 100860, 100820, 100810, 100790, 
    100760, 100780, 100790, 100800, 100800, 100790, 100790, 100780, 100780, 
    100790, 100820, 100810, 100800, 100800, 100820, 100810, 100800, 100800, 
    _, _, _, _, 100740, _, 100660, _, 100540, 100490, 100410, 100380, _, 
    100290, _, 100140, 100060, _, 100060, _, _, 100150, _, _, 100180, _, 
    100210, 100240, 100300, 100370, 100400, _, 100480, 100550, 100590, 
    100630, 100630, _, _, 100700, _, 100750, 100770, 100780, 100820, 100830, 
    100840, _, _, 100880, 100890, _, 100910, 100960, _, 100990, 100990, 
    101010, 101010, _, _, _, _, 101080, _, 101130, _, 101170, 101170, _, _, 
    101240, _, 101280, _, 101310, _, 101400, 101430, _, 101490, 101520, 
    101560, 101570, _, 101650, 101670, 101710, 101760, _, 101840, 101890, _, 
    101940, _, 101990, 102000, 102050, 102070, 102090, 102120, 102160, 
    102190, 102220, 102230, 102230, 102260, 102260, _, 102280, 102280, 
    102270, 102240, 102220, _, 102170, _, _, 102090, 102000, 101950, 101860, 
    101770, 101700, _, 101480, _, 101440, 101370, _, 101130, _, 101000, 
    100910, 100880, 100870, _, 101010, 100820, _, 100950, _, 100980, 101000, 
    101020, _, _, 101040, _, 101080, 101120, _, 101110, 101110, 101110, 
    101110, _, 101100, 101100, 101150, 101230, _, 101270, 101270, 101310, 
    101350, 101330, 101320, 101290, 101280, 101210, 101180, 101170, 101160, 
    101150, 101150, 101150, 101160, 101170, 101170, 101190, 101210, 101220, 
    101250, 101270, 101270, 101260, 101310, _, 101300, 101310, 101290, 
    101310, _, 101300, 101280, 101280, 101270, _, 101260, 101230, 101180, 
    101130, _, 101020, 100960, _, 100760, _, 100620, 100570, 100490, 100380, 
    _, 100270, 100220, 100170, 100110, _, 100070, 100070, 100070, 100080, _, 
    100110, 100100, 100100, 100100, _, 100120, 100140, 100140, 100130, _, _, 
    100120, 100110, 100080, 100050, 100020, _, 100000, 100000, 100000, 
    100000, 100000, 100020, 100060, 100090, 100100, 100140, _, _, 100250, 
    100230, _, 100260, 100290, 100280, 100300, _, 100300, 100350, 100320, 
    100340, _, 100370, 100410, 100420, 100500, _, 100600, 100660, 100690, 
    100740, _, 100800, 100790, 100840, 100820, _, 100800, 100820, 100870, 
    100890, _, 100900, 100900, 100900, 100900, 100900, 100870, 100880, _, 
    100910, _, 100930, 100930, 100940, 100900, _, 100910, 100890, 100870, 
    100860, 100840, 100820, _, 100790, 100750, 100720, 100700, 100640, 
    100630, 100600, 100580, 100580, 100560, 100560, 100570, 100550, 100540, 
    _, 100500, 100460, 100420, 100420, 100460, 100480, 100520, 100550, 
    100620, 100630, 100660, 100650, 100680, 100710, 100730, 100720, 100710, 
    100720, 100700, 100730, 100770, 100790, 100790, 100790, 100810, 100850, 
    100860, 100860, 100890, 100910, 100950, 100970, 101000, 101040, 101080, 
    101120, 101160, 101200, 101240, 101280, 101320, 101350, 101410, 101460, 
    101490, 101530, 101580, 101600, 101620, 101640, 101650, 101670, 101690, 
    101720, 101740, 101770, 101760, 101770, 101770, 101770, 101790, 101770, 
    101780, 101780, 101770, 101780, 101780, 101790, 101760, 101720, 101730, 
    101690, 101650, 101590, 101570, 101550, 101480, 101430, 101360, 101330, 
    101290, 101250, 101180, 101140, 101100, 101050, 101010, 100950, 100920, 
    100890, 100860, 100840, 100840, 100840, 100840, 100860, 100830, 100870, 
    100860, 100870, 100890, 100940, 100980, 100980, 100990, 101020, 101040, 
    101030, 101050, 101040, 101060, 101050, 101070, 101130, 101140, 101170, 
    101220, 101240, 101270, 101310, 101340, 101360, 101370, 101410, 101400, 
    101440, 101460, 101480, 101480, 101510, 101510, 101530, 101530, 101540, 
    101550, 101570, 101580, 101590, 101610, 101630, 101620, 101660, 101670, 
    101680, 101690, 101710, 101730, 101740, 101740, 101770, 101780, 101800, 
    101800, 101810, 101800, 101800, 101830, 101800, 101790, 101780, 101770, 
    101760, 101770, 101760, 101730, 101730, 101720, 101720, 101700, 101680, 
    101650, 101640, 101620, 101600, 101590, 101580, 101570, 101550, 101530, 
    101510, 101490, 101450, 101430, 101420, 101410, 101410, 101450, 101420, 
    101410, 101420, 101440, 101460, 101450, 101460, 101480, 101480, 101490, 
    101500, 101510, 101550, 101540, 101530, 101520, 101530, 101530, 101520, 
    101510, 101500, 101510, 101520, 101530, 101540, 101540, 101550, 101540, 
    101540, 101520, 101510, 101490, 101470, 101460, 101440, 101430, 101380, 
    101350, 101340, 101310, 101270, 101220, 101140, 101100, 100990, 101060, 
    101000, 100970, 100910, 100900, 100870, _, 100860, _, _, _, _, _, _, _, 
    _, _, _, 99860, _, _, _, _, _, _, _, _, _, 99150, 99190, 99310, 99410, 
    99470, 99600, 99660, 99770, 99850, 99950, 100040, 100120, 100250, 100350, 
    100480, 100550, 100620, 100690, 100750, 100790, 100840, 100890, 100960, 
    101030, 101080, 101140, 101180, 101240, 101290, 101330, 101350, 101410, 
    101460, 101530, 101580, 101640, 101730, 101750, 101820, 101860, 101880, 
    101900, 101970, 102000, 102000, 102020, 102070, 102110, 102160, 102160, 
    102210, 102230, 102230, 102220, 102220, 102250, 102270, 102280, 102290, 
    102290, 102300, 102330, 102330, 102340, 102330, 102330, 102310, 102300, 
    102290, 102310, 102320, 102320, 102340, 102360, 102360, 102350, 102340, 
    102320, 102310, 102280, 102310, 102310, 102320, 102320, 102340, 102340, 
    102330, 102330, 102360, 102360, 102370, 102360, 102400, 102420, 102440, 
    102470, 102500, 102540, 102540, 102560, 102560, 102560, 102570, 102590, 
    102610, 102600, 102620, 102630, 102620, 102610, 102610, 102600, 102600, 
    102570, 102560, 102550, 102500, 102500, 102510, 102470, 102420, 102390, 
    102380, 102390, 102370, 102360, 102300, 102260, 102240, 102220, 102250, 
    102230, 102160, 102150, 102170, 102180, 102170, 102110, 102100, 102080, 
    102080, 102080, 102090, 102110, 102110, 102050, 102100, 102100, 102090, 
    102080, 102060, 102060, 102040, 102010, 102010, 102000, 102010, 101960, 
    101990, 102010, 101990, 101970, 101970, 101930, 101940, 101920, 101800, 
    101840, 101920, 101810, 101770, 101740, 101780, 101800, 101800, 101780, 
    101730, 101710, 101680, 101740, 101720, 101720, 101690, 101680, 101760, 
    101790, 101750, 101700, 101760, 101720, 101770, 101790, 101710, 101640, 
    101700, 101720, 101720, 101740, 101740, 101700, 101590, 101680, 101570, 
    101550, 101540, 101500, 101450, 101400, 101360, 101470, 101430, 101410, 
    101410, 101450, 101470, 101440, 101480, 101460, 101480, 101460, 101440, 
    101430, 101420, 101400, 101400, 101370, 101380, 101340, 101320, 101330, 
    101290, 101250, 101230, 101220, 101210, 101180, 101180, 101160, 101150, 
    101150, 101130, 101110, 101090, 101090, 101080, 101090, 101050, 101040, 
    101050, 101020, 101020, 101030, 101050, 101040, 101010, 101010, 101000, 
    101020, 101030, 100990, 100990, 101010, 101030, 100980, 100980, 100980, 
    100990, 101000, 100970, 100970, 101000, 100970, 100950, 100910, 100890, 
    100860, 100850, 100850, 100830, 100860, 100850, 100830, 100780, 100780, 
    100720, 100700, 100700, 100680, 100660, 100640, 100650, 100640, 100630, 
    100620, 100610, 100630, 100640, 100640, 100670, 100680, 100710, 100730, 
    100780, 100810, 100840, 100850, 100870, 100960, 101010, 101030, 101030, 
    101100, 101160, 101190, 101250, 101280, 101280, 101300, 101290, 101300, 
    101340, 101350, 101360, 101360, 101380, 101380, 101360, 101380, 101380, 
    101370, 101340, 101300, 101270, 101260, 101260, 101240, 101270, 101270, 
    101250, 101240, 101220, 101120, 101080, 101040, 101040, 100950, 100920, 
    100960, 100960, 100840, 100750, 100660, 100590, 100520, 100390, 100330, 
    100290, 100220, 100190, 100230, 100260, 100310, 100450, 100390, 100410, 
    100380, 100390, 100340, 100310, 100320, 100300, 100270, 100230, 100200, 
    100200, 100180, 100160, 100140, 100140, 100110, 100060, 100060, 100050, 
    100060, 100060, 100100, 100120, 100080, 100090, 100070, 100050, 100000, 
    99980, 99940, 99930, 99940, 100010, 100010, 100030, 100050, 100080, 
    100130, 100150, 100170, 100200, 100260, 100290, 100320, 100360, 100400, 
    100480, 100520, 100570, 100610, 100630, 100650, 100710, 100780, 100850, 
    100890, 100910, 100960, 101030, 101090, 101140, 101150, 101180, 101210, 
    101270, 101350, 101410, 101480, 101540, 101550, 101580, 101590, 101610, 
    101640, 101650, 101630, 101670, 101670, 101680, 101680, 101680, 101690, 
    101700, 101700, 101700, 101710, 101700, 101680, 101700, 101710, 101730, 
    101750, 101770, 101760, 101770, 101800, 101820, 101820, 101830, 101820, 
    101820, 101830, 101820, 101820, 101800, 101800, 101780, 101750, 101720, 
    101720, 101690, 101670, 101650, 101640, 101620, 101600, 101590, 101560, 
    101510, 101540, 101460, 101440, 101390, 101360, 101350, 101330, 101310, 
    101310, 101310, 101290, 101260, 101250, 101250, 101270, 101280, 101280, 
    101310, 101310, 101330, 101370, 101400, 101420, 101460, 101490, 101530, 
    101590, 101620, 101640, 101650, 101680, 101700, 101720, 101760, 101750, 
    101700, 101720, 101770, 101800, 101830, 101860, 101880, 101920, 101940, 
    101990, 102040, 102100, 102140, 102170, 102200, 102240, 102250, 102280, 
    102300, 102290, 102310, 102330, 102370, 102380, 102380, 102370, 102360, 
    102380, 102360, 102360, 102360, 102360, 102350, 102370, 102360, 102360, 
    102360, 102350, 102330, 102310, 102320, 102310, 102290, 102270, 102240, 
    102240, 102260, 102220, 102180, 102190, 102170, 102160, 102160, 102120, 
    102100, 102070, 102060, 102060, 102060, 102050, 102030, 101990, 101980, 
    101950, 101950, 101920, 101880, 101840, 101830, 101810, 101780, 101740, 
    101710, 101680, 101660, 101640, 101600, 101570, 101520, 101490, 101490, 
    101460, 101440, 101420, 101380, 101360, 101330, 101300, 101280, 101250, 
    101230, 101210, 101190, 101170, 101170, 101150, 101130, 101110, 101090, 
    101060, 101040, 101020, 101000, 100980, 100980, 101000, 101030, 101030, 
    101010, 100990, 100990, 100970, 100950, 100880, 100830, 100810, 100790, 
    100770, 100750, 100730, 100710, 100720, 100710, 100710, 100720, 100720, 
    100710, 100720, 100730, 100780, 100820, 100850, 100860, 100890, 100890, 
    100910, 100930, 100940, 100960, 100970, 100980, 100990, 100990, 101010, 
    101020, 101010, 100990, 100980, 100970, 100960, 100940, 100930, 100920, 
    100920, 100910, 100920, 100940, 100940, 100960, 100990, 101020, 101050, 
    101100, 101130, 101130, 101160, 101200, 101210, 101220, 101250, 101260, 
    101260, 101260, 101250, 101260, 101260, 101250, 101280, 101300, 101330, 
    101320, 101300, 101300, 101310, 101300, 101270, 101250, 101210, 101190, 
    101150, 101120, 101090, 101070, 101050, 101030, 101020, 101010, 101000, 
    100960, 100930, 100930, 100930, 100940, 100940, 100960, 100950, 100940, 
    100910, 100900, 100880, 100860, 100860, 100840, 100840, 100850, 100830, 
    100830, 100800, 100780, 100780, 100780, 100750, 100720, 100710, 100710, 
    100720, 100730, 100750, 100760, 100760, 100770, 100750, 100740, 100710, 
    100690, 100670, 100670, 100650, 100650, 100620, 100610, 100620, 100620, 
    100630, 100590, 100550, 100520, 100510, 100530, 100530, 100530, 100550, 
    100540, 100540, 100530, 100520, 100500, 100480, 100430, 100420, 100410, 
    100410, 100410, 100400, 100400, 100380, 100370, 100340, 100330, 100320, 
    100320, 100330, 100340, 100370, 100380, 100380, 100390, 100390, 100390, 
    100400, 100410, 100420, 100430, 100430, 100450, 100460, 100460, 100480, 
    100480, 100500, 100480, 100470, 100450, 100430, 100380, 100380, 100370, 
    100360, 100330, 100310, 100250, 100160, 100170, 100150, 100130, 100110, 
    100090, 100070, 100060, 100090, 100090, 100070, 100060, 100040, 100040, 
    100030, 100010, 100010, 100000, 100020, 100030, 100040, 100060, 100060, 
    100080, 100090, 100110, 100120, 100140, 100160, 100200, 100240, 100270, 
    100300, 100330, 100360, 100360, 100360, 100370, 100380, 100380, 100380, 
    100380, 100400, 100380, 100400, 100450, 100460, 100460, 100460, 100470, 
    100450, 100460, 100460, 100450, 100450, 100380, 100370, 100380, 100360, 
    100300, 100280, 100300, 100260, 100220, 100210, 100190, 100160, 100160, 
    100160, 100160, 100140, 100130, 100110, 100110, 100100, 100100, 100110, 
    100100, 100110, 100140, 100150, 100140, 100140, 100170, 100180, 100210, 
    100210, 100240, 100250, 100290, 100310, 100330, 100360, 100390, 100420, 
    100480, 100500, 100520, 100540, 100560, 100570, 100600, 100640, 100660, 
    100680, 100680, 100700, 100720, 100740, 100750, 100770, 100770, 100780, 
    100800, 100800, 100800, 100800, 100790, 100790, 100770, 100770, 100760, 
    100750, 100740, 100730, 100720, 100710, 100700, 100700, 100690, 100680, 
    100700, 100700, 100700, 100700, 100680, 100680, 100670, 100700, 100710, 
    100730, 100720, 100730, 100750, 100770, 100780, 100790, 100800, 100800, 
    100800, 100790, 100790, 100810, 100810, 100830, 100820, 100800, 100760, 
    100730, 100680, 100660, 100640, 100630, 100610, 100580, 100540, 100500, 
    100470, 100420, 100360, 100330, 100300, 100270, 100290, 100310, 100370, 
    100470, 100590, 100700, 100750, 100800, 100810, 100870, 100910, 100970, 
    101010, 101050, 101100, 101130, 101180, 101220, 101280, 101310, 101340, 
    101350, 101380, 101410, 101410, 101410, 101410, 101400, 101370, 101350, 
    101350, 101340, 101320, 101310, 101340, 101330, 101340, 101360, 101390, 
    101430, 101440, 101460, 101510, 101530, 101540, 101550, 101570, 101590, 
    101590, 101590, 101560, 101550, 101580, 101590, 101570, 101560, 101520, 
    101470, 101450, 101410, 101390, 101340, 101290, 101230, 101170, 101090, 
    101020, 100900, 100820, 100740, 100620, 100490, 100380, 100310, 100270, 
    100260, 100250, 100310, 100360, 100420, 100500, 100560, 100640, 100730, 
    100830, 100900, 100990, 101040, 101140, 101210, 101290, 101290, 101300, 
    101210, 101220, 101140, 101120, 101100, 100970, 100920, 100860, 100820, 
    100750, 100710, 100730, 100680, 100680, 100700, 100730, 100840, 100930, 
    100970, 101010, 101070, 101150, 101220, 101210, 101180, 101140, 101100, 
    101080, 101070, 101060, 101040, 101020, 101010, 100960, 100920, 100910, 
    100860, 100840, 100830, 100820, 100830, 100800, 100790, 100750, 100760, 
    100740, 100690, 100610, 100530, 100470, 100480, 100390, 100310, 100250, 
    100200, 100120, 100050, 99990, 99930, 99860, 99810, 99730, 99700, 99710, 
    99730, 99730, 99790, 99800, 99830, 99850, 99860, 99860, 99860, 99880, 
    99910, 99920, 99950, 99980, 99950, 100020, 100080, 100140, 100180, 
    100260, 100300, 100340, 100390, 100480, 100530, 100560, 100590, 100620, 
    100640, 100600, 100570, 100510, 100470, 100370, 100320, 100240, 100200, 
    100120, 100140, 100080, 100210, 100390, 100520, 100580, 100650, 100720, 
    100770, 100800, 100800, 100870, 100890, 100950, 101050, 101080, 101080, 
    101100, 101180, 101220, 101240, 101270, 101290, 101330, 101350, 101350, 
    101360, 101410, 101440, 101420, 101400, 101430, 101430, 101410, 101400, 
    101370, 101320, 101220, 101150, 101110, 101070, 101020, 100900, 100810, 
    100730, 100690, 100650, 100610, 100580, 100530, 100510, 100470, 100410, 
    100380, 100310, 100280, 100230, 100170, 100120, 100130, 100100, 100090, 
    100070, 100060, 100070, 100050, 100030, 100010, 99990, 99960, 99970, 
    99980, 99960, 99950, 99910, 99880, 99880, 99850, 99850, 99840, 99830, 
    99910, 100000, 100120, 100190, 100260, 100350, 100400, 100450, 100510, 
    100530, 100530, 100540, 100540, 100550, 100520, 100520, 100480, 100430, 
    100400, 100340, 100250, 100180, 100090, 100060, 99990, 99930, 99890, 
    99830, 99760, 99700, 99620, 99620, 99580, 99560, 99470, 99380, 99280, 
    99180, 99140, 99050, 98940, 98850, 98810, 98810, 98780, 98740, 98740, 
    98680, 98630, 98610, 98550, 98500, 98450, 98410, 98390, 98360, 98270, 
    98240, 98150, 98110, 98050, 97990, 97940, 97870, 97820, 97770, 97720, 
    97680, 97630, 97590, 97560, 97540, 97550, 97530, 97530, 97570, 97620, 
    97690, 97750, 97800, 97850, 97900, 97950, 98040, 98100, 98190, 98270, 
    98390, 98490, 98590, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    99440, 99440, 99460, 99470, 99470, 99480, _, 99490, 99460, 99460, 99450, 
    99420, 99400, 99400, 99400, 99380, 99370, 99370, 99350, 99320, 99280, 
    99240, 99210, 99180, 99190, 99170, 99150, 99160, 99160, 99170, 99200, 
    99210, 99220, 99200, 99190, 99180, 99180, 99200, 99190, 99180, 99150, 
    99100, 99050, 99000, 98890, 98890, 98850, 98840, 98860, 98870, 98880, 
    98900, 98910, 98900, 98880, 98820, 98740, 98690, 98640, 98570, 98550, 
    98560, 98600, 98640, 98710, 98820, 98940, 99080, 99180, 99270, 99380, 
    99520, 99660, 99780, 99870, 99960, 100050, 100120, 100180, 100220, 
    100270, 100310, 100380, 100420, 100490, 100560, 100620, 100680, 100740, 
    100800, 100860, 100910, 100970, 101000, 101060, 101090, 101110, 101140, 
    101170, 101190, 101200, 101190, 101180, 101170, 101190, 101180, 101180, 
    101160, 101160, 101180, 101140, 101120, 101100, 101090, 101080, 101070, 
    101070, 101070, 101020, 100990, 100990, 100970, 100960, 100980, 100980, 
    100980, 101000, 101040, 101070, 101100, 101140, 101170, 101200, 101230, 
    101250, 101290, 101320, 101350, 101370, 101380, 101420, 101450, 101470, 
    101500, 101500, 101510, 101490, 101490, 101480, 101470, 101460, 101450, 
    101430, 101420, 101410, 101370, 101350, 101320, 101290, 101280, 101230, 
    101210, 101190, 101150, 101130, 101110, 101080, 101040, 101000, 100980, 
    100950, 100940, 100890, 100870, 100820, 100790, 100760, 100730, 100700, 
    100670, 100640, 100620, 100600, 100570, 100550, 100550, 100570, 100600, 
    100640, 100670, 100700, 100760, 100800, 100850, 100880, 100920, 100980, 
    101030, 101110, 101170, 101230, 101250, 101300, 101340, 101410, 101440, 
    101450, 101500, 101550, 101600, 101640, 101660, 101720, 101730, 101760, 
    101770, 101770, 101790, 101790, 101810, 101800, 101850, 101860, 101860, 
    101870, 101900, 101900, 101920, 101930, 101930, 101920, 101950, 101950, 
    101920, 101990, 102000, 102030, 102050, 102050, 102040, 102030, 102020, 
    102040, 102070, 102040, 102050, 102100, 102090, 102110, 102160, 102110, 
    102110, 102120, 102090, 102070, 102070, 102070, 102050, 102050, 102050, 
    102020, 102010, 102020, 101970, 101950, 101960, 101960, 101890, 101860, 
    101880, 101890, 101880, 101830, 101820, 101800, 101780, 101760, 101730, 
    101730, 101720, 101730, 101700, 101710, 101740, 101730, 101730, 101700, 
    101710, 101710, 101690, 101670, 101670, 101680, 101690, 101670, 101660, 
    101670, 101650, 101610, 101590, 101510, 101490, 101440, 101480, 101510, 
    101510, 101510, 101500, 101500, 101490, 101470, 101460, 101510, 101520, 
    101530, 101480, 101530, 101540, 101530, 101530, 101530, 101580, 101520, 
    101520, 101620, 101630, 101550, 101590, 101570, 101560, 101580, 101540, 
    101530, 101480, 101460, 101360, 101300, 101230, 101190, 101140, 100990, 
    100930, 100880, 100760, 100600, 100530, 100450, 100330, 100210, 100090, 
    100030, 99930, 99800, 99680, 99620, 99600, 99530, 99400, 99450, 99390, 
    99320, 99250, 99280, 99230, 99190, 99240, 99260, 99270, 99330, 99370, 
    99460, 99560, 99670, 99760, 99860, 99960, 100070, 100170, 100300, 100430, 
    100550, 100590, 100710, 100820, 100890, 100990, 101070, 101150, 101240, 
    101310, 101420, 101480, 101530, 101610, 101680, 101750, 101810, 101830, 
    101870, 101940, 102000, 102000, 102050, 102050, 102050, 102060, 102060, 
    102090, 102060, 102040, 102010, 101970, 101960, 101940, 101890, 101840, 
    101800, 101760, 101710, 101670, 101650, 101580, 101520, 101490, 101430, 
    101360, 101320, 101280, 101270, 101240, 101240, 101210, 101190, 101160, 
    101130, 101100, 100980, 100980, 100980, 100910, 100860, 100880, 100800, 
    100750, 100730, 100730, 100680, 100700, 100680, 100680, 100690, 100630, 
    100610, 100550, 100450, 100310, 100230, 100110, 99850, 99720, 99590, 
    99600, 99350, 99230, 99170, 99040, 99060, 99140, 99200, 99330, 99450, 
    99630, 99790, 99950, 100180, 100310, 100350, 100470, 100460, 100500, 
    100570, 100600, 100660, 100660, 100720, 100780, 100870, 100950, 101030, 
    101090, 101140, 101230, 101270, 101350, 101370, 101500, 101500, 101580, 
    101600, 101650, 101660, 101670, 101660, 101660, 101680, 101690, 101690, 
    101730, 101750, 101770, 101780, 101780, 101800, 101750, 101740, 101700, 
    101650, 101610, 101520, 101460, 101350, 101170, 100930, 100730, 100670, 
    100630, 100600, 100570, 100590, 100630, 100690, 100730, 100810, 100870, 
    100910, 101020, 101100, 101180, 101180, 101120, 101100, 101170, 101110, 
    101070, 101020, 101020, 101020, 100980, 101010, 101090, 101150, 101240, 
    101320, 101390, 101440, 101530, 101610, 101700, 101780, 101850, 101870, 
    101890, 101890, 101880, 101930, 101930, 101950, 101950, 101920, 101910, 
    101900, 101860, 101840, 101830, 101800, 101780, 101780, 101800, 101810, 
    101830, 101860, 101880, 101920, 101910, 101970, 101980, 102040, 102060, 
    102090, 102110, 102100, 102110, 102090, 102080, 102050, 102030, 102000, 
    101940, 101850, 101800, 101780, 101750, 101710, 101700, 101710, 101680, 
    101690, 101690, 101700, 101680, 101710, 101710, 101710, 101730, 101740, 
    101760, 101780, 101790, 101790, 101820, 101820, 101800, 101800, 101810, 
    101820, 101840, 101850, 101830, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    100930, 100830, 100810, 100750, 100760, 100730, 100730, 100720, 100710, 
    100680, 100630, 100610, 100560, 100520, 100510, 100470, 100430, 100390, 
    100360, 100310, 100300, 100270, 100270, 100270, 100310, 100300, 100280, 
    100270, 100270, 100270, 100260, 100270, 100280, 100290, 100320, 100340, 
    100360, 100350, 100400, 100400, 100420, 100460, 100460, 100460, 100500, 
    100600, 100580, 100570, 100550, _, 100500, 100430, 100430, 100330, 
    100280, 100250, 100150, 100040, 100040, 99960, 99900, 99850, 99730, 
    99540, 99410, 99220, 99140, 99080, 98970, 98900, 98880, 98900, 98930, 
    98960, 98980, 98990, 99030, 99040, 99040, 99070, 99110, 99150, 99200, 
    99230, 99250, 99290, 99290, 99290, 99280, 99250, 99290, 99250, 99280, 
    99300, 99330, 99350, 99360, 99390, 99420, 99410, 99400, 99400, 99410, 
    99420, 99420, 99450, 99520, 99550, 99510, 99470, 99490, 99510, 99530, 
    99550, 99560, 99570, 99600, 99620, 99640, 99720, 99730, 99770, 99790, 
    99800, 99800, 99870, 99930, 99990, 100030, 100030, 100060, 100090, 
    100090, 100120, 100130, 100150, 100180, 100270, 100360, 100450, 100520, 
    100610, 100680, 100760, 100830, 100890, 100960, 101010, 101030, 101080, 
    101130, 101220, 101280, 101370, 101450, 101530, 101630, 101680, 101780, 
    101870, 101960, 102060, 102140, 102220, 102280, 102300, 102350, 102380, 
    102390, 102400, 102350, 102280, 102220, 102160, 102120, 102090, 102020, 
    101900, 101830, 101750, 101670, 101580, 101510, 101440, 101360, 101330, 
    101250, 101190, 101140, 101050, 100970, 100860, 100770, 100630, 100550, 
    100490, 100430, 100400, 100390, 100430, 100480, 100530, 100590, 100670, 
    100760, 100860, 100960, 101150, 101370, 101560, 101680, 101800, 101930, 
    102080, 102160, 102280, 102370, 102460, 102550, 102650, 102620, 102650, 
    102630, 102630, 102590, 102500, 102500, 102420, 102310, 102200, 102090, 
    101990, 101840, 101710, 101530, 101370, 101180, 101080, 100910, 100790, 
    100650, 100530, 100500, 100380, 100380, 100410, 100420, 100400, 100450, 
    100500, 100540, 100630, 100720, 100810, 100860, 100970, 101070, 101090, 
    101290, 101320, 101460, 101570, 101650, 101790, 101920, 102060, 102160, 
    102290, 102330, 102400, 102450, 102500, 102490, 102540, 102560, 102540, 
    102530, 102520, 102550, 102560, 102600, 102650, 102660, 102660, 102680, 
    102690, 102710, 102700, 102710, 102670, 102630, 102580, 102500, 102430, 
    102340, 102300, 102250, 102210, 102200, 102130, 102080, 102030, 101970, 
    101920, 101840, 101790, 101730, 101660, 101630, 101550, 101540, 101510, 
    101500, 101450, 101450, 101430, 101390, 101360, 101350, 101330, 101350, 
    101370, 101420, 101450, 101530, 101560, 101580, 101520, 101560, 101550, 
    101520, 101490, 101450, 101420, 101410, 101380, 101300, 101230, 101170, 
    101100, 101040, 100990, 100950, 100920, 100920, 100950, 100960, 100990, 
    101020, 101040, 101080, 101130, 101190, 101230, 101250, 101280, 101310, 
    101330, 101360, 101400, 101440, 101490, 101520, 101550, 101590, 101600, 
    101620, 101660, 101680, 101710, 101740, 101790, 101820, 101840, 101850, 
    101890, 101910, 101950, 101980, 102010, 102040, 102050, 102090, 102140, 
    102180, 102190, 102180, 102200, 102190, 102210, 102220, 102190, 102170, 
    102170, 102170, 102160, 102130, 102100, 102080, 102040, 102040, 101950, 
    101920, 101910, 101820, 101810, 101740, 101680, 101600, 101500, 101380, 
    101230, 101110, 100990, 100840, 100690, 100560, 100470, 100370, 100280, 
    100230, 100160, 100130, 100080, 100080, 100050, 100000, 99960, 99870, 
    99800, 99690, 99630, 99540, 99510, 99480, 99510, 99580, 99650, 99590, 
    99540, 99460, 99420, 99410, 99300, 99330, 99320, 99380, 99460, 99590, 
    99720, 99850, 99950, 100140, 100190, 100350, 100410, 100510, 100640, 
    100780, 100880, 100990, 101010, 101050, 101090, 101090, 101160, 101300, 
    101370, 101380, 101430, 101460, 101490, 101520, 101540, 101530, 101550, 
    101560, 101590, 101620, 101650, 101660, 101700, 101710, 101720, 101740, 
    101740, 101720, 101720, 101700, 101680, 101660, 101610, 101600, 101560, 
    101530, 101510, 101480, 101480, 101460, 101450, 101450, 101460, 101460, 
    101500, 101500, 101510, 101530, 101550, 101550, 101570, 101570, 101550, 
    101550, 101580, 101540, 101540, 101560, 101550, 101510, 101470, 101430, 
    101420, 101430, 101430, 101420, 101400, 101450, 101460, 101460, 101450, 
    101450, 101430, 101420, 101420, 101390, 101360, 101340, 101290, 101280, 
    101250, 101230, 101220, 101200, 101190, 101180, 101150, 101150, 101150, 
    101150, 101190, 101200, 101190, 101260, 101290, 101290, 101290, 101290, 
    101310, 101310, 101300, 101280, 101230, 101210, 101150, 101130, 101020, 
    100970, 100940, 100870, 100770, 100740, 100640, 100600, 100540, 100530, 
    100520, 100530, 100580, 100710, 100750, 100770, 100810, 100880, 101020, 
    101040, 101100, 101210, 101310, 101410, 101480, 101570, 101610, 101650, 
    101660, 101720, 101760, 101810, 101890, 101980, 102070, 102140, 102220, 
    102330, 102450, 102530, 102620, 102710, 102800, 102910, 102990, 103070, 
    103140, 103160, 103200, 103220, 103210, 103240, 103240, 103240, 103200, 
    103210, 103150, 103120, 103170, 103120, 103060, 103050, 102980, 102930, 
    102920, 102860, 102830, 102780, 102750, 102670, 102690, 102700, 102690, 
    102690, 102660, 102670, 102690, 102670, 102650, 102680, 102640, 102630, 
    102650, 102620, 102610, 102570, 102510, 102450, 102440, 102450, 102360, 
    102410, 102320, 102280, 102260, 102200, 102160, 102120, 102060, 102010, 
    101960, 101910, 101890, 101860, 101810, 101790, 101760, 101720, 101680, 
    101640, 101600, 101530, 101500, 101460, 101410, 101370, 101340, 101300, 
    101260, 101230, 101180, 101150, 101140, 101090, 101050, 101040, 101010, 
    100910, 100950, 101010, 100990, 101000, 101080, 101130, 101150, 101210, 
    101220, 101230, 101240, 101280, 101300, 101290, 101290, 101320, 101360, 
    101350, 101380, 101380, 101380, 101420, 101430, 101450, 101470, 101500, 
    101530, 101560, 101550, 101540, 101520, 101520, 101520, 101530, 101550, 
    101570, 101590, 101620, 101660, 101690, 101720, 101710, 101710, 101720, 
    101730, 101760, 101750, 101780, 101770, 101770, 101820, 101850, 101860, 
    101860, 101870, 101910, 101920, 101930, 101940, 101970, 102040, 102070, 
    102070, 102070, 102150, 102180, 102180, 102160, 102250, 102380, 102440, 
    102490, 102540, 102580, 102620, 102750, 102790, 102820, 102890, 102970, 
    103020, 103060, 103090, 103140, 103180, 103210, 103250, 103260, 103310, 
    103340, 103360, 103390, 103410, 103410, 103420, 103430, 103440, 103440, 
    103470, 103500, 103510, 103540, 103540, 103550, 103530, 103550, 103550, 
    103550, 103560, 103560, 103560, 103550, 103560, 103560, 103550, 103520, 
    103510, 103500, 103490, 103460, 103440, 103440, 103440, 103450, 103440, 
    103450, 103450, 103440, 103440, 103460, 103440, 103430, 103440, 103450, 
    103450, 103440, 103420, 103420, 103400, 103400, 103360, 103340, 103300, 
    103280, 103270, 103260, 103250, 103240, 103200, 103180, 103140, 103110, 
    103080, 103040, 103020, 103000, 102970, 102940, 102910, 102880, 102870, 
    102840, 102820, 102800, 102790, 102780, 102780, 102790, 102800, 102790, 
    102800, 102810, 102840, 102860, 102830, 102820, 102840, 102860, 102880, 
    102900, 102900, 102910, 102920, 102940, 102950, 102950, 102940, 102930, 
    102960, 102960, 102970, 102970, 102970, 102980, 102970, 103010, 103010, 
    103010, 103000, 102990, 102970, 102970, 102970, 102960, 102950, 102960, 
    102940, 102910, 102900, 102880, 102850, 102830, 102790, 102760, 102740, 
    102730, 102690, 102650, 102650, 102630, 102590, 102570, 102520, 102480, 
    102410, 102380, 102350, 102310, 102260, 102220, 102180, 102120, 102080, 
    102060, 102030, 102010, 102000, 102010, 102030, 102080, 102120, 102140, 
    102170, 102180, 102190, 102210, 102210, 102210, 102210, 102210, 102220, 
    102220, 102190, 102170, 102160, 102130, 102100, 102060, 102020, 101950, 
    101900, 101850, 101760, 101690, 101600, 101530, 101460, 101380, 101300, 
    101240, 101180, 101120, 101050, 100990, 100940, 100860, 100790, 100730, 
    100680, 100620, 100560, 100500, 100460, 100390, 100320, 100260, 100190, 
    100120, 100020, 99970, 99900, 99800, 99730, 99640, 99550, 99470, 99350, 
    99320, 99180, 99070, 99020, 98910, 98790, 98670, 98610, 98510, 98370, 
    98220, 98130, 98080, 98010, 98000, 98020, 98180, 98330, 98430, 98560, 
    98740, 98700, 98940, 98770, 98910, 99030, 99150, 99260, 99530, 99570, 
    99540, 99680, 99810, 99840, 99770, 99860, 99970, 100010, 100060, 100080, 
    100240, 100340, 100400, 100520, 100550, 100710, 100780, 100870, 100870, 
    100940, 101090, 101150, 101250, 101300, 101360, 101430, 101460, 101500, 
    101580, 101610, 101650, 101660, 101700, 101730, 101800, 101850, 101870, 
    101890, 101920, 101970, 101980, 102010, 102060, 102100, 102130, 102150, 
    102180, 102200, 102230, 102240, 102240, 102240, 102250, 102270, 102250, 
    102250, 102220, 102190, 102180, 102160, 102130, 102100, 102080, 102040, 
    102010, 101970, 101930, 101870, 101830, 101820, 101800, 101790, 101800, 
    101810, 101800, 101720, 101670, 101620, 101570, 101530, 101520, 101480, 
    101470, 101470, 101460, 101420, 101390, 101310, 101290, 101260, 101210, 
    101160, 101110, 101080, 101030, 100990, 100960, 100930, 100880, 100840, 
    100810, 100770, 100730, 100680, 100610, 100550, 100500, 100460, 100420, 
    100400, 100390, 100350, 100260, 100220, 100180, 100150, 100120, 100090, 
    100060, 100040, 100030, 100050, 100030, 100010, 99970, 99930, 99870, 
    99830, 99760, 99660, 99600, 99480, 99430, 99370, 99330, 99180, 99000, 
    98900, 98810, 98660, 98550, 98380, 98220, 98060, 97950, 97830, 97730, 
    97700, 97610, 97530, 97550, 97640, 97730, 97860, 97910, 98000, 98050, 
    98130, 98190, 98240, 98290, 98320, 98410, 98510, 98570, 98660, 98760, 
    98840, 98930, 99000, 99070, 99100, 99110, 99140, 99140, 99120, 99080, 
    98990, 98920, 98840, 98790, 98730, 98690, 98680, 98670, 98710, 98740, 
    98780, 98800, 98830, 98830, 98860, 98860, 98910, 98950, 98970, 99000, 
    99150, 99300, 99420, 99550, 99750, 99880, 100080, 100290, 100460, 100610, 
    100740, 100810, 100970, 101110, 101160, 101220, 101320, 101390, 101420, 
    101500, 101540, 101610, 101660, 101680, 101740, 101780, 101820, 101820, 
    101870, 101910, 101940, 101960, 101960, 101990, 101990, 101980, 101960, 
    101950, 101930, 101940, 101920, 101920, 101920, 101870, 101810, 101780, 
    101800, 101750, 101710, 101680, 101630, 101590, 101540, 101470, 101460, 
    101390, 101350, 101350, 101310, 101290, 101240, 101190, 101150, 101110, 
    101030, 100980, 100970, 100910, 100890, 100830, 100810, 100770, 100720, 
    100750, 100670, 100640, 100640, 100680, 100720, 100720, 100760, 100750, 
    100740, 100720, 100710, 100810, 100840, 100850, 100850, 100860, 100870, 
    100900, 100900, 100900, 100890, 100960, 100980, 101020, 101030, 101060, 
    101060, 101110, 101130, 101160, 101200, 101200, 101230, 101240, 101230, 
    101240, 101270, 101270, 101290, 101280, 101300, 101310, 101330, 101340, 
    101350, 101370, 101400, 101400, 101420, 101420, 101440, 101450, 101490, 
    101520, 101570, 101600, 101640, 101660, 101680, 101690, 101700, 101720, 
    101750, 101790, 101800, 101830, 101830, 101850, 101860, 101870, 101870, 
    101860, 101890, 101880, 101890, 101920, 101960, 101980, 101980, 101990, 
    101990, 101970, 102000, 102010, 101980, 101980, 101980, 101980, 101970, 
    101980, 101950, 101940, 101900, 101860, 101810, 101760, 101730, 101740, 
    101750, 101820, 101870, 101900, 101900, 101900, 101900, 101910, 101900, 
    101900, 101880, 101870, 101850, 101850, 101830, 101820, 101820, 101820, 
    101800, 101790, 101750, 101740, 101680, 101620, 101620, 101580, 101570, 
    101570, 101560, 101550, 101500, 101480, 101440, 101390, 101330, 101350, 
    101330, 101300, 101290, 101300, 101290, 101270, 101230, 101220, 101210, 
    101190, 101170, 101150, 101130, 101120, 101090, 101070, 101090, 101070, 
    101080, 101090, 101110, 101140, 101170, 101220, 101250, 101300, 101340, 
    101360, 101410, 101400, 101380, 101490, 101520, 101620, 101700, 101730, 
    101790, 101820, 101840, 101840, 101870, 101910, 101900, 101870, 101880, 
    101860, 101860, 101840, 101810, 101790, 101780, 101780, 101760, 101730, 
    101700, 101670, 101640, 101620, 101580, 101570, 101560, 101540, 101550, 
    101540, 101520, 101490, 101500, 101480, 101470, 101450, 101420, 101420, 
    101360, 101360, 101370, 101400, 101380, 101370, _, 101360, 101330, 
    101340, 101300, 101330, 101300, 101270, 101270, 101290, 101300, 101300, 
    101300, 101250, 101260, 101280, 101280, 101260, 101270, 101240, 101230, 
    101180, 101160, 101170, 101160, 101200, 101170, 101230, 101240, 101260, 
    101270, 101290, 101310, 101320, 101360, 101330, 101340, 101330, 101330, 
    101360, 101370, 101380, 101410, 101400, 101430, 101460, 101500, 101520, 
    101500, 101530, 101530, 101560, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 101620, 101620, 101580, 101540, 
    101490, 101470, 101390, 101340, 101330, 101310, 101350, 101290, 101240, 
    101200, 101160, 101130, 101080, 101040, 101000, 100970, 100950, 100910, 
    100880, 100850, 100810, 100790, 100790, 100760, 100730, 100700, 100660, 
    100620, 100600, 100580, 100560, 100550, 100560, 100560, 100580, 100600, 
    100630, 100640, 100660, 100670, 100680, 100670, 100660, 100740, 100670, 
    100660, 100680, 100680, 100670, 100590, 100530, 100490, 100410, 100290, 
    100220, 100110, 99930, 99840, 99690, 99520, 99370, 99360, 99400, 99550, 
    99660, 99760, 99860, 99970, 100030, 100120, 100190, 100220, 100220, 
    100270, 100280, 100360, 100390, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 100730, 100700, 100660, 100630, 100580, 100530, 
    100490, 100420, 100400, 100340, 100280, 100220, 100170, 100120, 100070, 
    100020, 99940, 99900, 99900, 99920, 99940, 99970, 99990, 100030, 100080, 
    100100, 100140, 100150, 100180, 100190, 100230, 100220, 100220, 100220, 
    100190, 100140, 100120, 100090, 100060, 99970, 99930, 99860, 99840, 
    99860, 99870, 99880, 99880, _, 99920, 99960, 100020, 100050, 100080, 
    100160, 100150, 100210, 100260, 100260, 100270, 100230, 100220, 100190, 
    100200, 100150, 100070, 100110, 100150, 100160, 100180, 100170, 100150, 
    100140, 100130, 100110, 100100, 100120, 100110, 100110, 100070, 100030, 
    100000, 99970, 99950, 99930, 99900, 99860, 99820, 99820, 99730, 99650, 
    99710, 99680, 99660, 99650, 99610, 99580, 99550, 99530, 99500, 99450, 
    99450, 99450, 99470, 99470, 99510, 99570, 99620, 99660, 99700, 99730, 
    99750, 99750, 99760, 99710, 99620, 99530, 99560, 99510, 99420, 99310, 
    99210, 99100, 98920, 98760, 98500, 98220, 97920, 97560, 97170, 96720, 
    96440, 96220, 96010, 95970, 95990, 96110, 96200, 96370, 96610, 96770, 
    97000, 97160, 97340, 97460, 97620, 97730, 97870, 97950, 98050, 98140, 
    98180, 98280, 98350, 98410, 98450, 98420, 98380, 98330, 98260, 98200, 
    98150, 98040, 97860, 97660, 97360, 97040, 96830, 96790, 96780, 96750, 
    96810, 96840, 96850, 96910, 96930, 96890, 96820, 96830, 96880, 96850, 
    96830, 96890, 96970, 97040, 97090, 97150, 97280, 97380, 97460, 97480, 
    97430, 97410, 97420, 97470, 97440, 97470, 97490, 97500, 97480, 97470, 
    97440, 97380, 97290, 97250, 97190, 97150, 97140, 97100, 97100, 97080, 
    97070, 97110, 97110, 97110, 97140, 97130, 97140, 97150, 97140, 97130, 
    97130, 97170, 97170, 97270, 97320, 97370, 97420, 97470, 97520, 97560, 
    97580, 97640, 97660, 97680, 97660, 97730, 97780, 97790, 97820, 97800, 
    97830, 97850, 97850, 97870, 97870, 97900, 97910, 97920, 97910, 97920, 
    97950, 97980, 97970, 98010, 98060, 98080, 98120, 98150, 98170, 98140, 
    98130, 98130, 98120, 98130, 98130, 98140, 98130, 98120, 98120, 98080, 
    98060, 98030, 98010, 98050, 98020, 97970, 97920, 97970, 97960, 97970, 
    98010, 98090, 98070, 98020, 98050, 98170, 98260, 98340, 98400, 98470, 
    98560, 98630, 98700, 98780, 98910, 98950, 99060, 99170, 99220, 99280, 
    99460, 99660, 99820, 99930, 100040, 100150, 100270, 100370, 100480, 
    100570, 100660, 100730, 100800, 100870, 100910, 100960, 100980, 101020, 
    101060, 101130, 101150, 101180, 101240, 101330, 101380, 101460, 101510, 
    101520, 101490, 101550, 101580, 101580, 101510, 101450, 101430, 101360, 
    101240, 101150, 101080, 100980, 100820, 100620, 100530, 100420, 100280, 
    100190, 100110, 100010, 100020, 99940, 99910, 99850, 99800, 99690, 99720, 
    99840, 99960, 100070, 100110, 100200, 100200, 100270, 100410, 100490, 
    100570, 100640, 100680, 100750, 100800, 100850, 100920, 100980, 101000, 
    101040, 101050, 101070, 101050, 101050, 101100, 101160, 101210, 101190, 
    101160, 101140, 101130, 101160, 101130, 101110, 101100, 101060, 101080, 
    101110, 101120, 101140, 101140, 101150, 101180, 101170, 101220, 101280, 
    101300, 101350, 101420, 101470, 101530, 101620, 101720, 101770, 101810, 
    101900, 101990, 102050, 102100, 102120, 102180, 102240, 102280, 102340, 
    102340, 102350, 102370, 102400, 102410, 102420, 102420, 102440, 102480, 
    102510, 102540, 102560, 102580, 102550, 102580, 102570, 102590, 102600, 
    102630, 102630, 102660, 102610, 102620, 102630, 102640, 102610, 102600, 
    102530, 102500, 102490, 102480, 102490, 102450, 102430, 102370, 102370, 
    102340, 102290, 102250, 102250, 102230, 102230, 102200, 102170, 102160, 
    102140, 102160, 102160, 102150, 102120, 102120, 102110, 102110, 102110, 
    102070, 102080, 102070, 102100, 102080, 102060, 102040, 102030, 102020, 
    102000, 101980, 101960, 101900, 101870, 101850, 101790, 101750, 101660, 
    101640, 101610, 101550, 101520, 101480, 101410, 101380, 101350, 101340, 
    101340, 101300, 101240, 101240, 101190, 101180, 101130, 101060, 100990, 
    100910, 100830, 100780, 100740, 100710, 100670, 100670, 100650, 100630, 
    100600, 100570, 100540, 100480, 100420, 100380, 100300, 100170, 99980, 
    99910, 99780, 99620, 99480, 99260, 99100, 98940, 98910, 98800, 98690, 
    98570, 98480, 98400, 98350, 98320, 98300, 98300, 98340, 98390, 98460, 
    98490, 98570, 98650, 98720, 98790, 98880, 98920, 98960, 98950, 98950, 
    98910, 98890, 98860, 98890, 98840, 98760, 98710, 98750, 98760, 98730, 
    98680, 98670, 98670, 98640, 98660, 98690, 98670, 98680, 98710, 98720, 
    98720, 98740, 98770, 98770, 98760, 98770, 98820, 98890, 98910, 98930, 
    98960, 98980, 99030, 99050, 99080, 99100, 99130, 99140, 99180, 99240, 
    99260, 99280, 99310, 99320, 99330, 99330, 99340, 99310, 99330, 99330, 
    99330, 99350, 99380, 99380, 99370, 99350, 99340, 99320, 99340, 99320, 
    99320, 99290, 99280, 99240, 99260, 99220, 99140, 99120, 99070, 99070, 
    99010, 98980, 98930, 98830, 98760, 98730, 98690, 98620, 98510, 98440, 
    98380, 98290, 98190, 98100, 98090, 98090, 98100, 98080, 98180, 98150, 
    98170, 98140, 98160, 98160, 98150, 98170, 98160, 98200, 98220, 98260, 
    98290, 98330, 98350, 98380, 98390, 98440, 98450, 98440, 98470, 98470, 
    98490, 98480, 98500, 98530, 98550, 98550, 98540, 98550, 98530, 98560, 
    98560, 98600, 98600, 98630, 98650, 98660, 98680, 98700, 98720, 98730, 
    98740, 98760, 98790, 98820, 98860, 98910, 98990, 99010, 99060, 99060, 
    99100, 99120, 99150, 99160, 99180, 99200, 99200, 99220, 99210, 99220, 
    99210, 99210, 99160, 99170, 99140, 99140, 99150, 99180, 99230, 99300, 
    99350, 99410, 99450, 99490, 99510, 99550, 99570, 99580, 99640, 99670, 
    99700, 99730, 99780, 99790, 99830, 99860, 99870, 99870, 99840, 99840, 
    99840, 99850, 99830, 99810, 99820, 99790, 99770, 99780, 99760, 99680, 
    99720, 99670, 99670, 99710, 99620, 99630, 99640, 99670, 99680, 99670, 
    99690, 99730, 99760, 99760, 99780, 99820, 99840, 99880, 99890, 99940, 
    99970, 100010, 100030, 100040, 100060, 100080, 100110, 100150, 100170, 
    100220, 100250, 100320, 100370, 100450, 100460, 100460, 100410, 100390, 
    100360, 100280, 100180, 100060, 99940, 99840, 99690, 99540, 99370, 99210, 
    99030, 98840, 98610, 98380, 98170, 98050, 97910, 97730, 97590, 97490, 
    97460, 97470, 97470, 97470, 97380, 97270, 97210, 97140, 97110, 97020, 
    96970, 96970, 96940, 96830, 96750, 96740, 96750, 96780, 96760, 96810, 
    97000, 97140, 97260, 97360, 97440, 97470, 97560, 97620, 97680, 97750, 
    97770, 97780, 97850, 97880, 97880, 97900, 97900, 97850, 97810, 97810, 
    97750, 97750, 97740, 97750, 97800, 97830, 97870, 97900, 97930, 97920, 
    97890, 97870, 97880, 97850, 97800, 97750, 97700, 97650, 97630, 97600, 
    97530, 97570, 97610, 97600, 97620, 97640, 97670, 97700, 97710, 97740, 
    97730, 97690, 97640, 97630, 97620, 97610, 97620, 97650, 97650, 97730, 
    97830, 97940, 98040, 98080, 98140, 98200, 98240, 98270, 98320, 98370, 
    98450, 98520, 98620, 98670, 98730, 98780, 98830, 98850, 98920, 98980, 
    99010, 99060, 99190, 99370, 99520, 99660, 99800, 99930, 100030, 100150, 
    100260, 100340, 100430, 100500, 100620, 100700, 100740, 100790, 100860, 
    100900, 100940, 100970, 101010, 101050, 101020, 101030, 101060, 101050, 
    101050, 101070, 101090, 101100, 101090, 101090, 101080, 101100, 101110, 
    101110, 101110, 101110, 101120, 101120, 101080, 101050, 101020, 100980, 
    100970, 100950, 100910, 100900, 100880, 100880, 100880, 100850, 100820, 
    100780, 100790, 100740, 100700, 100690, 100630, 100590, 100530, 100520, 
    100480, 100430, 100400, 100350, 100290, 100190, 100060, 99930, 99790, 
    99640, 99550, 99450, 99390, 99270, 99100, 98970, 98840, 98670, 98540, 
    98360, 98220, 98180, 98140, 98090, 98080, 98040, 98100, 98120, 98110, 
    98150, 98170, 98230, 98280, 98340, 98230, 98310, 98370, 98420, 98470, 
    98480, 98450, 98440, 98440, 98450, 98450, 98490, 98540, 98630, 98710, 
    98800, 98900, 98980, 99070, 99190, 99310, 99440, 99520, 99670, 99760, 
    99890, 100000, 100060, 100100, 100190, 100220, 100240, 100270, 100290, 
    100250, 100310, 100410, 100400, 100420, 100470, 100460, 100410, 100390, 
    100320, 100280, 100240, 100200, 100120, 100110, 100110, 100100, 100050, 
    100020, 99960, 99850, 99820, 99740, 99700, 99610, 99580, 99610, 99610, 
    99620, 99680, 99720, 99740, 99780, 99840, 99910, 99950, 100050, 100120, 
    100200, 100210, 100220, 100230, 100230, 100210, 100200, 100160, 100140, 
    100120, 100100, 100080, 100100, 100110, 100160, 100160, 100170, 100210, 
    100200, 100170, 100140, 100190, 100140, 100130, 100100, 100080, 100070, 
    100020, 99970, 99930, 99870, 99800, 99750, 99700, 99670, 99640, 99620, 
    99610, 99580, 99550, 99540, 99510, 99510, 99520, 99500, 99540, 99520, 
    99520, 99530, 99550, 99560, 99580, 99590, 99590, 99580, 99620, 99740, 
    99780, 99820, 99860, 99940, 100000, 100020, 100030, 100070, 100050, 
    100000, 100010, 100100, 100150, 100250, 100290, 100310, 100410, 100490, 
    100560, 100620, 100660, 100720, 100780, 100880, 100970, 101030, 101030, 
    101040, 101070, 101060, 101040, 101040, 101010, 101070, 101110, 101200, 
    101230, 101260, 101300, 101370, 101410, 101450, 101490, 101490, 101540, 
    101660, 101610, 101620, 101590, 101630, 101620, 101610, 101590, 101570, 
    101550, 101510, 101460, 101380, 101330, 101300, 101250, 101230, 101200, 
    101160, 101140, 101130, 101110, 101090, 101060, 101050, 101030, 101010, 
    100980, 100940, 100940, 100920, 100890, 100900, 100930, 100940, 100940, 
    100930, 100930, 100900, 100860, 100850, 100870, 100870, 100850, 100870, 
    100860, 100880, 100890, 100860, 100820, 100770, 100740, 100710, 100640, 
    100590, 100530, 100510, 100470, 100420, 100400, 100360, 100350, 100350, 
    100360, 100390, 100410, 100430, 100500, 100510, 100510, 100550, 100540, 
    100580, 100640, 100710, 100730, 100800, 100840, 100820, 100860, 100850, 
    100840, 100780, 100750, 100680, 100630, 100530, 100540, 100500, 100480, 
    100450, 100430, 100410, 100460, 100430, 100420, 100410, 100380, 100390, 
    100390, 100340, 100290, 100350, 100450, 100490, 100560, 100610, 100670, 
    100760, 100780, 100850, 100900, 100910, 100960, 100980, 101030, 101080, 
    101150, 101130, 101160, 101130, 101170, 101230, 101240, 101290, 101310, 
    101350, 101370, 101400, 101390, 101370, 101340, 101300, 101250, 101210, 
    101210, 101190, 101150, 101140, 101180, 101200, 101200, 101200, 101220, 
    101270, 101330, 101400, 101440, 101510, 101590, 101650, 101710, 101840, 
    101950, 102030, 102110, 102180, 102270, 102310, 102380, 102450, 102530, 
    102590, 102630, 102700, 102790, 102850, 102850, 102890, 102870, 102830, 
    102840, 102820, 102790, 102770, 102740, 102730, 102740, 102730, 102730, 
    102720, 102760, 102760, 102750, 102760, 102730, 102750, 102750, 102760, 
    102800, 102760, 102770, 102750, 102750, 102720, 102710, 102730, 102710, 
    102710, 102830, 102830, 102810, 102830, 102820, 102780, 102780, 102760, 
    102720, 102720, 102680, 102680, 102650, 102610, 102550, 102500, 102460, 
    102370, 102230, 102130, 102020, 101920, 101750, 101630, 101510, 101430, 
    101300, 101210, 101190, 101050, 100980, 100930, 100950, 100980, 101020, 
    101020, 100980, 100990, 100980, 100910, 100860, 100780, 100710, 100590, 
    100470, 100340, 100210, 100080, 99980, 99840, 99680, 99540, 99430, 99300, 
    99160, 99000, 98870, 98750, 98610, 98500, 98420, 98350, 98310, 98270, 
    98210, 98220, 98240, 98340, 98430, 98460, 98590, 98670, 98820, 98980, 
    99130, 99230, 99280, 99410, 99470, 99500, 99480, 99440, 99510, 99440, 
    99550, 99690, 99730, 99790, 99860, 99940, 100040, 100130, 100220, 100350, 
    100470, 100540, 100630, 100710, 100810, 100870, 100980, 101170, 101270, 
    101390, 101520, 101610, 101680, 101740, 101790, 101870, 101930, 101970, 
    102000, 102040, 102020, 101990, 101970, 101930, 101910, 101850, 101800, 
    101780, 101730, 101680, 101620, 101570, 101460, 101390, 101300, 101230, 
    101190, 101140, 101100, 101050, 101010, 100970, 100850, 100790, 100750, 
    100720, 100700, 100720, 100710, 100660, 100680, 100680, 100660, 100620, 
    100650, 100620, 100610, 100630, 100650, 100590, 100530, 100580, 100650, 
    100670, 100660, 100670, 100640, 100600, 100610, 100630, 100670, 100670, 
    100650, 100700, 100740, 100740, 100740, 100770, 100750, 100750, 100730, 
    100740, 100720, 100720, 100700, 100720, 100730, 100770, 100800, 100800, 
    100780, 100740, 100750, 100740, 100730, 100740, 100730, 100740, 100790, 
    100790, 100820, 100810, 100800, 100760, 100720, 100690, 100690, 100690, 
    100660, 100660, 100640, 100650, 100630, 100620, 100610, 100600, 100580, 
    100560, 100550, 100500, 100450, 100410, 100370, 100340, 100300, 100280, 
    100220, 100180, 100100, 100080, 100010, 99960, 99910, 99850, 99810, 
    99770, 99750, 99660, 99540, 99450, 99370, 99270, 99170, 99060, 98920, 
    98770, 98690, 98620, 98520, 98430, 98480, 98540, 98600, 98630, 98680, 
    98750, 98830, 98820, 98850, 98970, 99030, 99010, 98980, 99000, 99060, 
    99070, 99140, 99230, 99250, 99280, 99350, 99390, 99370, 99430, 99610, 
    99640, 99640, 99740, 99840, 99800, 99780, 99840, 99940, 100060, 100220, 
    100320, 100270, 100290, 100320, 100270, 100300, 100290, 100270, 100260, 
    100240, 100210, 100160, 100130, 100090, 100060, 100030, 99990, 99950, 
    99890, 99860, 99840, 99820, 99780, 99720, 99700, 99740, 99750, 99750, 
    99730, 99710, 99700, 99660, 99660, 99630, 99630, 99640, 99630, 99610, 
    99580, 99550, 99510, 99450, 99450, 99400, 99390, 99370, 99400, 99470, 
    99520, 99530, 99460, 99470, 99470, 99540, 99680, 99570, 99530, 99600, 
    99590, 99550, 99530, 99460, 99420, 99400, 99370, 99410, 99440, 99470, 
    99490, 99500, 99550, 99560, 99610, 99660, 99700, 99670, 99740, 99810, 
    99860, 99870, 99930, 99970, 99970, 99970, 100080, 100100, 100150, 100190, 
    100210, 100210, 100260, 100290, 100370, 100450, 100500, 100540, 100630, 
    100700, 100760, 100800, 100890, 100950, 100980, 101020, 101070, 101130, 
    101190, 101240, 101300, 101330, 101370, 101410, 101450, 101470, 101480, 
    101500, 101520, 101560, 101590, 101620, 101650, 101660, 101680, 101700, 
    101710, 101690, 101700, 101790, 101860, 101890, 101890, 101860, 101870, 
    101830, 101770, 101750, 101780, 101820, 101820, 101800, 101820, 101850, 
    101850, 101830, 101810, 101770, 101740, 101740, 101690, 101630, 101560, 
    101540, 101500, 101460, 101390, 101290, 101270, 101260, 101200, 101120, 
    101070, 101010, 100980, 100930, 100880, 100840, 100830, 100800, 100730, 
    100680, 100630, 100610, 100680, 100650, 100630, 100580, 100560, 100510, 
    100490, 100460, 100420, 100430, 100420, 100450, 100460, 100460, 100460, 
    100460, 100490, 100500, 100540, 100570, 100560, 100610, 100630, 100630, 
    100650, 100670, 100690, 100700, 100730, 100760, 100770, 100790, 100800, 
    100770, 100780, 100800, 100860, 100860, 100850, 100840, 100850, 100870, 
    100860, 100930, 100960, 100980, 101030, 101060, 101100, 101100, 101130, 
    101200, 101240, 101310, 101340, 101350, 101390, 101400, 101420, 101490, 
    101520, 101530, 101500, 101530, 101550, 101590, 101590, 101610, 101580, 
    101580, 101570, 101570, 101560, 101570, 101570, 101530, 101520, 101510, 
    101490, 101480, 101450, 101430, 101400, 101340, 101340, 101380, 101320, 
    101290, 101280, 101290, 101280, 101240, 101240, 101230, 101210, 101210, 
    101210, 101200, 101190, 101160, 101100, 101060, 101020, 101010, 100910, 
    100830, 100760, 100710, 100620, 100630, 100590, 100460, 100460, 100390, 
    100360, 100350, 100360, 100460, 100480, 100590, 100660, 100730, 100780, 
    100800, 100860, 100940, 101010, 101070, 100970, 100930, 101040, 101090, 
    101170, 101150, 101140, 101150, 101190, 101240, 101260, 101300, 101310, 
    101330, 101360, 101390, 101410, 101390, 101400, 101410, 101440, 101470, 
    101470, 101490, 101530, 101540, 101560, 101570, 101560, 101580, 101610, 
    101600, 101610, 101630, 101660, 101680, 101670, 101660, 101620, 101590, 
    101560, 101500, 101370, 101280, 101220, 101170, 101040, 100890, 100850, 
    100830, 100840, 100780, 100810, 100740, 100730, 100740, 100730, 100770, 
    100790, 100820, 100860, 100910, 100980, 101030, 101060, 101090, 101130, 
    101180, 101230, 101290, 101370, 101420, 101480, 101520, 101560, 101560, 
    101560, 101570, 101580, 101570, 101590, 101590, 101600, 101580, 101570, 
    101570, 101560, 101550, 101520, 101470, 101400, 101350, 101290, 101250, 
    101200, 101150, 101130, 101060, 100970, 100830, 100710, 100590, 100460, 
    100280, 100090, 99990, 99870, 99660, 99450, 99280, 99140, 98990, 98800, 
    98620, 98320, 97910, 97540, 97290, 97360, 97280, 97380, 97480, 97550, 
    97550, 97440, 97470, 97440, 97370, 97320, 97290, 97280, 97350, 97380, 
    97440, 97510, 97600, 97720, 97830, 98000, 98170, 98380, 98570, 98740, 
    98910, 99050, 99170, 99290, 99410, 99510, 99560, 99680, 99810, 99950, 
    100080, 100170, 100270, 100320, 100430, 100530, 100660, 100670, 100720, 
    100740, 100800, 100830, 100810, 100810, 100810, 100740, 100640, 100550, 
    100430, 100380, 100280, 100180, 99990, 99930, 99860, 99800, 99690, 99670, 
    99640, 99670, 99710, 99680, 99680, 99630, 99670, 99640, 99640, 99630, 
    99630, 99640, 99630, 99590, 99560, 99540, 99480, 99420, 99300, 99220, 
    99120, 99020, 98850, 98700, 98560, 98530, 98390, 98350, 98270, 98240, 
    98170, 98050, 97990, 97980, 97960, 97940, 97880, 97830, 97770, 97760, 
    97760, 97780, 97750, 97760, 97790, 97820, 97850, 97890, 97970, 97990, 
    98010, 98040, 98090, 98100, 98100, 98130, 98160, 98150, 98150, 98140, 
    98150, 98140, 98130, 98120, 98110, 98100, 98080, 98070, 98020, 98010, 
    98010, 97960, 97940, 97890, 97860, 97830, 97780, 97730, 97720, 97680, 
    97640, 97610, 97610, 97600, 97570, 97560, 97530, 97510, 97480, 97520, 
    97510, 97520, 97540, 97570, 97590, 97630, 97670, 97700, 97720, 97750, 
    97780, 97820, 97870, 97910, 97970, 98020, 98070, 98110, 98120, 98120, 
    98130, 98140, 98160, 98170, 98160, 98170, 98190, 98180, 98180, 98180, 
    98180, 98200, 98180, 98170, 98160, 98200, 98220, 98220, 98250, 98270, 
    98280, 98310, 98330, 98360, 98370, 98370, 98380, 98400, 98450, 98500, 
    98520, 98500, 98510, 98540, 98570, 98550, 98550, 98560, 98560, 98550, 
    98550, 98550, 98550, 98550, 98560, 98580, 98600, 98600, 98620, 98630, 
    98650, 98670, 98690, 98740, 98770, 98820, 98880, 98930, 98980, 99050, 
    99090, 99160, 99210, 99270, 99350, 99390, 99460, 99520, 99570, 99610, 
    99700, 99780, 99830, 99900, 99950, 100000, 100030, 100120, 100160, 
    100180, 100240, 100320, 100350, 100360, 100400, 100430, 100460, 100490, 
    100510, 100530, 100540, 100540, 100550, 100550, 100510, 100530, 100530, 
    100520, 100500, 100500, 100510, 100520, 100500, 100490, 100500, 100510, 
    100470, 100400, 100380, 100370, 100300, 100210, 100140, 100140, 100040, 
    100060, 99970, 99760, 99740, 99620, 99390, 99370, 99340, 99250, 99150, 
    99080, 99060, 99100, 99040, 98990, 98960, 98950, 98980, 99010, 99050, 
    99100, 99150, 99220, 99290, 99330, 99430, 99470, 99540, 99560, 99610, 
    99620, 99660, 99700, 99720, 99760, 99760, 99760, 99810, 99850, 99830, 
    99840, 99810, 99820, 99760, 99770, 99700, 99710, 99720, 99720, 99700, 
    99690, 99680, 99650, 99700, 99740, 99750, 99710, 99800, 99870, 99850, 
    99880, 99880, 99790, 99750, 99750, 99730, 99700, 99610, 99500, 99470, 
    99400, 99260, 99230, 99110, 99070, 99070, 99030, 98970, 98940, 98890, 
    98940, 98960, 99030, 98990, 99000, 99040, 99110, 99180, 99240, 99310, 
    99380, 99400, 99380, 99450, 99520, 99560, 99600, 99620, 99630, 99640, 
    99650, 99730, 99670, 99620, 99670, 99630, 99710, 99730, 99810, 99860, 
    99840, 99850, 99910, 99970, 100020, 100100, 100180, 100140, 100100, 
    100120, 100200, 100300, 100400, 100470, 100540, 100620, 100660, 100720, 
    100760, 100800, 100820, 100820, 100800, 100810, 100850, 100850, 100850, 
    100820, 100790, 100820, 100830, 100810, 100790, 100770, 100800, 100820, 
    100850, 100840, 100760, 100780, 100740, 100760, 100740, 100710, 100680, 
    100700, 100700, 100720, 100700, 100620, 100580, 100550, 100520, 100520, 
    100520, 100520, 100480, 100470, 100480, 100470, 100470, 100390, 100340, 
    100330, 100290, 100300, 100290, 100280, 100320, 100310, 100320, 100330, 
    100330, 100340, 100360, 100360, 100360, 100370, 100400, 100390, 100380, 
    100390, 100400, 100410, 100420, 100420, 100430, 100460, 100470, 100460, 
    100490, 100500, 100520, 100530, 100570, 100610, 100630, 100650, 100660, 
    100650, 100660, 100670, 100670, 100660, 100660, 100690, 100680, 100690, 
    100710, 100720, 100730, 100760, 100760, 100750, 100760, 100760, 100780, 
    100810, 100840, 100870, 100880, 100880, 100920, 100920, 100950, 100940, 
    100970, 100990, 100980, 100980, 101040, 101080, 101110, 101100, 101100, 
    101120, 101150, 101150, 101120, 101120, 101120, 101140, 101160, 101180, 
    101210, 101250, 101300, 101320, 101300, 101240, 101230, 101200, 101200, 
    101170, 101150, 101110, 101100, 101080, 101060, 100990, 100930, 100910, 
    100870, 100830, 100820, 100810, 100780, 100750, 100690, 100660, 100630, 
    100570, 100540, 100490, 100460, 100450, 100420, 100410, 100430, 100380, 
    100430, 100460, 100470, 100500, 100540, 100540, 100560, 100610, 100650, 
    100670, 100710, 100770, 100770, 100800, 100820, 100870, 100880, 100930, 
    100970, 100980, 100960, 100970, 101000, 101080, 101130, 101090, 101220, 
    101270, 101290, 101310, 101310, 101320, 101370, 101370, 101370, 101390, 
    101390, 101360, 101330, 101340, 101380, 101410, 101410, 101420, 101420, 
    101380, 101320, 101400, 101400, 101380, 101340, 101340, 101380, 101400, 
    101420, 101450, 101470, 101470, 101560, 101600, 101600, 101620, 101590, 
    101540, 101550, 101570, 101620, 101770, 101800, 101820, 101810, 101810, 
    101830, 101810, 101850, 101860, 101890, 101920, 101980, 101990, 101990, 
    102030, 102030, 102070, 102060, 102060, 102070, 102080, 102090, 102080, 
    102070, 102040, 102060, 102060, 102060, 102040, 102020, 101950, 101950, 
    101950, 101940, 101870, 101820, 101790, 101750, 101760, 101790, 101810, 
    101830, 101830, 101800, 101810, 101840, 101850, 101840, 101840, 101830, 
    101830, 101840, 101850, 101810, 101790, 101750, 101750, 101730, 101720, 
    101710, 101690, 101690, 101690, 101680, 101680, 101670, 101670, 101660, 
    101650, 101620, 101630, 101610, 101600, 101580, 101580, 101550, 101540, 
    101510, 101480, 101470, 101470, 101460, 101450, 101440, 101440, 101430, 
    101450, 101440, 101450, 101470, 101490, 101480, 101500, 101520, 101510, 
    101530, 101540, 101540, 101550, 101600, 101610, 101620, 101660, 101670, 
    101690, 101690, 101700, 101710, 101750, 101760, 101800, 101860, 101870, 
    101900, 101930, 101960, 101990, 102020, 102020, 102040, 102040, 102060, 
    102090, 102110, 102140, 102170, 102190, 102210, 102240, 102260, 102290, 
    102290, 102310, 102330, 102350, 102380, 102380, 102380, 102380, 102390, 
    102400, 102400, 102380, 102370, 102360, 102350, 102340, 102330, 102300, 
    102280, 102280, 102260, 102240, 102220, 102200, 102170, 102180, 102160, 
    102140, 102140, 102130, 102120, 102090, 102070, 102030, 101970, 101880, 
    101830, 101770, 101720, 101670, 101650, 101640, 101660, 101740, 101730, 
    101760, 101790, 101800, 101840, 101860, 101780, 101960, 101880, 102080, 
    102080, 102070, 102070, 102020, 101970, 102000, 102030, 102020, 102060, 
    102100, 102030, 102070, 102060, 102080, 102040, 102010, 102020, 101970, 
    101950, 101970, 101960, 101930, 101850, 101860, 101740, 101690, 101690, 
    101610, 101580, 101640, 101610, 101590, 101640, 101650, 101710, 101750, 
    101770, 101780, 101800, 101830, 101860, 101880, 101890, 101890, 101870, 
    101890, 101910, 101950, 101990, 102030, 102040, 102040, 102060, 102060, 
    102070, 102060, 102080, 102080, 102090, 102100, 102120, 102140, 102130, 
    102140, 102160, 102160, 102170, 102180, 102190, 102200, 102220, 102230, 
    102260, 102260, 102270, 102260, 102260, 102250, 102230, 102210, 102170, 
    102150, 102210, 102190, 102160, 102140, 102140, 102130, 102110, 102090, 
    102070, 102050, 102030, 102040, 102030, 102010, 102000, 101990, 101950, 
    101950, 101920, 101910, 101890, 101860, 101850, 101840, 101830, 101850, 
    101840, 101860, 101880, 101900, 101900, 101910, 101920, 101940, 101950, 
    101950, 101880, 101940, 101930, 101920, 101890, 101890, 101820, 101700, 
    101580, 101580, 101590, 101600, 101610, 101620, 101620, 101610, 101630, 
    101650, 101640, 101730, 101760, 101720, 101710, 101750, 101740, 101750, 
    101710, 101640, 101620, 101660, 101640, 101670, 101690, 101740, 101700, 
    101640, 101610, 101610, 101610, 101590, 101600, 101550, 101500, 101470, 
    101470, 101560, 101570, 101590, 101620, 101640, 101670, 101680, 101690, 
    101710, 101700, 101720, 101740, 101770, 101770, 101790, 101830, 101870, 
    101880, 101870, 101870, 101870, 101890, 101860, 101860, 101880, 101920, 
    101900, 101920, 101900, 101880, 101860, 101840, 101790, 101670, 101670, 
    101710, 101730, 101720, 101710, 101710, 101700, 101710, 101670, 101650, 
    101630, 101600, 101590, 101580, 101560, 101550, 101530, 101520, 101540, 
    101500, 101440, 101440, 101410, 101420, 101420, 101390, 101380, 101390, 
    101390, 101350, 101330, 101290, 101280, 101270, 101270, 101260, 101250, 
    101250, 101200, 101220, 101240, 101260, 101300, 101300, 101300, 101310, 
    101300, 101340, 101360, 101360, 101370, 101370, 101350, 101340, 101310, 
    101340, 101330, 101350, 101330, 101290, 101260, 101270, 101240, 101220, 
    101220, 101230, 101230, 101240, 101260, 101300, 101320, 101310, 101340, 
    101340, 101340, 101390, 101430, 101430, 101460, 101490, 101510, 101490, 
    101510, 101530, 101540, 101540, 101560, 101570, 101600, 101620, 101610, 
    101640, 101630, 101610, 101600, 101590, 101560, 101550, 101520, 101500, 
    101420, 101350, 101280, 101190, 101120, 101040, 100990, 100930, 100860, 
    100820, 100830, 100920, 100900, 100930, 100950, 100970, 101030, 101100, 
    101140, 101140, 101180, 101190, 101190, 101200, 101180, 101200, 101150, 
    101130, 101100, 101040, 101030, 100970, 100920, 100890, 100840, 100800, 
    100770, 100730, 100710, 100650, 100690, 100700, 100700, 100720, 100760, 
    100770, 100800, 100790, 100830, 100850, 100830, 100860, 100860, 100890, 
    100890, 100930, 100950, 101020, 101160, 101250, 101390, 101510, 101590, 
    101670, 101760, 101820, 101940, 102010, 102110, 102200, 102250, 102370, 
    102450, 102560, 102630, 102670, 102740, 102780, 102850, 102890, 102920, 
    102960, 103030, 103050, 103060, 103130, 103160, 103170, 103200, 103190, 
    103180, 103200, 103180, 103170, 103150, 103130, 103100, 103080, 103040, 
    103010, 102960, 102910, 102880, 102830, 102790, 102740, 102660, 102620, 
    102580, 102550, 102530, 102480, 102420, 102370, 102310, 102280, 102170, 
    102140, 102100, 102110, 102110, 102110, 102120, 102100, 102080, 102090, 
    102090, 102100, 102150, 102210, 102260, 102280, 102320, 102340, 102360, 
    102380, 102430, 102450, 102450, 102450, 102450, 102460, 102490, 102520, 
    102540, 102560, 102580, 102600, 102630, 102630, 102590, 102570, 102610, 
    102600, 102590, 102560, 102530, 102480, 102450, 102350, 102260, 102190, 
    102090, 101990, 101890, 101780, 101660, 101600, 101510, 101390, 101310, 
    101320, 101230, 101210, 101200, 101130, 101100, 101080, 101070, 101090, 
    101050, 101080, 101100, 101130, 101170, 101180, 101250, 101290, 101320, 
    101390, 101460, 101520, 101550, 101580, 101620, 101630, 101670, 101700, 
    101760, 101800, 101830, 101850, 101890, 101910, 101900, 101950, 102030, 
    102130, 102190, 102210, 102230, 102240, 102250, 102280, 102320, 102310, 
    102330, 102340, 102360, 102380, 102340, 102340, 102330, 102280, 102270, 
    102240, 102260, 102270, 102270, 102280, 102310, 102320, 102290, 102310, 
    102390, 102300, 102300, 102310, 102360, 102350, 102340, 102380, 102320, 
    102410, 102440, 102400, 102430, 102500, 102670, 102600, 102580, 102600, 
    102640, 102650, 102740, 102750, 102750, 102760, 102790, 102830, 102860, 
    102880, 102900, 102920, 102920, 102950, 102950, 102930, 102920, 102900, 
    102940, 102940, 102960, 102970, 102980, 102980, 103000, 103000, 103020, 
    103040, 103070, 103070, 103070, 103070, 103050, 103030, 103020, 103020, 
    103010, 102980, 102980, 102950, 102940, 102910, 102910, 102900, 102890, 
    102880, 102880, 102870, 102900, 102960, 102990, 103040, 103050, 103100, 
    103130, 103170, 103190, 103220, 103250, 103270, 103290, 103290, 103330, 
    103340, 103340, 103340, 103340, 103340, 103330, 103340, 103330, 103340, 
    103350, 103330, 103320, 103310, 103300, 103280, 103270, 103260, 103220, 
    103210, 103180, 103170, 103190, 103180, 103150, 103140, 103140, 103120, 
    103110, 103090, 103070, 103060, 103050, 103080, 103070, 103100, 103090, 
    103100, 103090, 103080, 103060, 103050, 103060, 103060, 103040, 103050, 
    103070, 103070, 103080, 103060, 103070, 103050, 103040, 103030, 103010, 
    103020, 103030, 103050, 103060, 103070, 103090, 103090, 103080, 103070, 
    103070, 103040, 103040, 103020, 103010, 103010, 103010, 102990, 102980, 
    102970, 102940, 102910, 102910, 102890, 102880, 102860, 102880, 102880, 
    102890, 102880, 102910, 102920, 102900, 102920, 102930, 102930, 102930, 
    102910, 102890, 102870, 102900, 102870, 102870, 102850, 102820, 102800, 
    102790, 102770, 102740, 102730, 102730, 102750, 102750, 102730, 102730, 
    102740, 102710, 102690, 102680, 102660, 102610, 102540, 102470, 102400, 
    102340, 102290, 102220, 102160, 102060, 101970, 101900, 101820, 101740, 
    101640, 101570, 101510, 101420, 101360, 101280, 101240, 101210, 101240, 
    101290, 101340, 101380, 101420, 101420, 101430, 101480, 101520, 101560, 
    101590, 101550, 101540, 101570, 101580, 101570, 101560, 101550, 101540, 
    101530, 101530, 101560, 101540, 101510, 101490, 101500, 101520, 101540, 
    101530, 101510, 101550, 101520, 101590, 101640, 101670, 101760, 101780, 
    101770, 101770, 101820, 101830, 101870, 101840, 101900, 102060, 102080, 
    102080, 102030, 102050, 102140, 102160, 102180, 102180, 102180, 102200, 
    102180, 102190, 102230, 102180, 102200, 102200, 102200, 102190, 102190, 
    102190, 102190, 102210, 102220, 102220, 102200, 102210, 102220, 102230, 
    102230, 102220, 102200, 102190, 102150, 102140, 102150, 102150, 102140, 
    102120, 102110, 102100, 102110, 102110, 102090, 102090, 102090, 102100, 
    102100, 102130, 102140, 102130, 102110, 102110, 102100, 102090, 102080, 
    102080, 102070, 102060, 102050, 102050, 102040, 102040, 102010, 102020, 
    102020, 102020, 102000, 101960, 101960, 101970, 101960, 101970, 101980, 
    101990, 101960, 101940, 101920, 101880, 101870, 101840, 101810, 101800, 
    101770, 101740, 101700, 101680, 101640, 101620, 101580, 101530, 101460, 
    101400, 101350, 101310, 101290, 101260, 101220, 101170, 101130, 101100, 
    101050, 101000, 100950, 100890, 100840, 100820, 100780, 100740, 100710, 
    100690, 100700, 100690, 100670, 100640, 100620, 100600, 100570, 100540, 
    100520, 100510, 100500, 100490, 100500, 100460, 100410, 100360, 100320, 
    100310, 100280, 100270, 100270, 100290, 100310, 100340, 100360, 100380, 
    100380, 100400, 100430, 100460, 100480, 100510, 100540, 100580, 100630, 
    100650, 100680, 100700, 100720, 100750, 100760, 100790, 100800, 100820, 
    100830, 100850, 100870, 100890, 100900, 100920, 100930, 100950, 100970, 
    100980, 100980, 100980, 101010, 101010, 101030, 101050, 101060, 101090, 
    101110, 101120, 101160, 101200, 101220, 101220, 101220, 101210, 101210, 
    101190, 101190, 101160, 101130, 101100, 101090, 101040, 101100, 101140, 
    101160, 101180, 101190, 101190, 101220, 101240, 101240, 101230, 101230, 
    101250, 101250, 101240, 101240, 101240, 101230, 101250, 101260, 101260, 
    101260, 101280, 101290, 101310, 101300, 101320, 101350, 101370, 101410, 
    101430, 101460, 101480, 101520, 101530, 101540, 101540, 101550, 101550, 
    101570, 101600, 101640, 101680, 101720, 101750, 101780, 101800, 101830, 
    101850, 101900, 101950, 101980, 102020, 102060, 102100, 102130, 102160, 
    102190, 102190, 102220, 102230, 102250, 102240, 102260, 102270, 102290, 
    102310, 102310, 102320, 102320, 102290, 102260, 102230, 102250, 102240, 
    102230, 102230, 102200, 102230, 102220, 102180, 102170, 102120, 102090, 
    102070, 102010, 101990, 101950, 101920, 101910, 101820, 101720, 101700, 
    101630, 101590, 101510, 101390, 101330, 101330, 101260, 101200, 101230, 
    101200, 101220, 101200, 101170, 101140, 101160, 101170, 101190, 101220, 
    101260, 101300, 101340, 101380, 101400, 101410, 101440, 101440, 101450, 
    101480, 101470, 101490, 101520, 101560, 101530, 101560, 101590, 101640, 
    101670, 101750, 101800, 101810, 101820, 101850, 101930, 101960, 102020, 
    101990, 101990, 102020, 102010, 102080, 102060, 102090, 102130, 102140, 
    102180, 102190, 102210, 102210, 102250, 102320, 102320, 102370, 102390, 
    102430, 102470, 102500, 102540, 102550, 102590, 102610, 102640, 102690, 
    102700, 102730, 102750, 102760, 102780, 102800, 102870, 102900, 102900, 
    102940, 102970, 102990, 103010, 103040, 103040, 103050, 103100, 103110, 
    103100, 103110, 103090, 103080, 103070, 103050, 103070, 103050, 103030, 
    103020, 103000, 102980, 102990, 102980, 102950, 102940, 102930, 102910, 
    102890, 102860, 102830, 102810, 102790, 102760, 102710, 102660, 102620, 
    102580, 102560, 102510, 102480, 102430, 102400, 102370, 102340, 102360, 
    102320, 102310, 102320, 102290, 102290, 102300, 102310, 102300, 102300, 
    102320, 102310, 102320, 102330, 102340, 102360, 102360, 102370, 102380, 
    102390, 102420, 102440, 102450, 102460, 102450, 102460, 102490, 102490, 
    102490, 102510, 102520, 102510, 102540, 102530, 102540, 102540, 102550, 
    102530, 102520, 102480, 102460, 102440, 102430, 102420, 102410, 102410, 
    102370, 102370, 102350, 102370, 102350, 102360, 102350, 102330, 102340, 
    102360, 102340, 102320, 102320, 102300, 102290, 102300, 102290, 102270, 
    102240, 102250, 102250, 102210, 102220, 102220, 102230, 102220, 102220, 
    102230, 102220, 102220, 102210, 102220, 102220, 102220, 102230, 102250, 
    102220, 102200, 102200, 102200, 102160, 102140, 102150, 102150, 102120, 
    102120, 102130, 102140, 102100, 102050, 102060, 102080, 102100, 102100, 
    102090, 102110, 102100, 102090, 102070, 102080, 102080, 102090, 102090, 
    102100, 102100, 102140, 102170, 102200, 102220, 102240, 102300, 102350, 
    102380, 102420, 102470, 102530, 102600, 102650, 102710, 102740, 102760, 
    102800, 102830, 102850, 102880, 102900, 102920, 102910, 102930, 102940, 
    102930, 102950, 102930, 102900, 102910, 102880, 102880, 102870, 102830, 
    102840, 102820, 102800, 102790, 102750, 102730, 102730, 102710, 102650, 
    102620, 102570, 102540, 102580, 102550, 102520, 102520, 102460, 102450, 
    102420, 102390, 102350, 102360, 102360, 102360, 102410, 102460, 102470, 
    102490, 102500, 102500, 102460, 102440, 102410, 102340, 102290, 102230, 
    102150, 102070, 101950, 101830, 101760, 101670, 101620, 101590, 101550, 
    101530, 101570, 101590, 101580, 101570, 101590, 101590, 101620, 101590, 
    101580, 101590, 101580, 101550, 101520, 101480, 101430, 101390, 101380, 
    101340, 101320, 101310, 101280, 101230, 101150, 101120, 101080, 101050, 
    101010, 101030, 101030, 101010, 101010, 101020, 101010, 100990, 100990, 
    100960, 100960, 100920, 100920, 100900, 100850, 100840, 100800, 100830, 
    100810, 100790, 100760, 100700, 100650, 100640, 100670, 100630, 100590, 
    100530, 100540, 100540, 100470, 100420, 100380, 100220, 100210, 100200, 
    100180, 100150, 100120, 100110, 100020, 99950, 99900, 99870, 99820, 
    99810, 99820, 99880, 99920, 99990, 100010, 100030, 100110, 100160, 
    100210, 100280, 100300, 100280, 100330, 100380, 100400, 100430, 100450, 
    100460, 100470, 100480, 100490, 100490, 100490, 100490, 100480, 100500, 
    100490, 100510, 100510, 100510, 100480, 100480, 100480, 100480, 100430, 
    100430, 100420, 100420, 100410, 100420, 100420, 100430, 100450, 100420, 
    100430, 100430, 100460, 100480, 100480, 100510, 100520, 100550, 100580, 
    100620, 100640, 100650, 100660, 100660, 100690, 100700, 100690, 100690, 
    100700, 100720, 100740, 100740, 100730, 100700, 100680, 100690, 100690, 
    100690, 100690, 100680, 100690, 100710, 100720, 100720, 100730, 100720, 
    100720, 100710, 100730, 100720, 100710, 100680, 100680, 100700, 100700, 
    100720, 100730, 100720, 100710, 100700, 100690, 100690, 100670, 100670, 
    100680, 100700, 100710, 100720, 100710, 100720, 100710, 100740, 100730, 
    100710, 100710, 100700, 100690, 100690, 100680, 100670, 100680, 100670, 
    100650, 100600, 100580, 100560, 100530, 100520, 100520, 100540, 100540, 
    100500, 100490, 100470, 100460, 100430, 100430, 100430, 100460, 100470, 
    100480, 100500, 100510, 100530, 100540, 100560, 100570, 100580, 100610, 
    100630, 100630, 100670, 100680, 100730, 100760, 100780, 100780, 100800, 
    100800, 100810, 100830, 100840, 100840, 100840, 100860, 100860, 100860, 
    100880, 100870, 100880, 100880, 100880, 100870, 100870, 100890, 100910, 
    100920, 100930, 100930, 100940, 100940, 100950, 100960, 100970, 100960, 
    100980, 100990, 100960, 100960, 100960, 100970, 100990, 100990, 100970, 
    100970, 100960, 100960, 100960, 100940, 100970, 100970, 100980, 100980, 
    100990, 101020, 101020, 101010, 101000, 101000, 101010, 101010, 101020, 
    101030, 101020, 101020, 101020, 101000, 101010, 101020, 101020, 101030, 
    101020, 100990, 101000, 101010, 101040, 101040, 101040, 101040, 101030, 
    101010, 101020, 101000, 101010, 101010, 101020, 101010, 101000, 101010, 
    101020, 101030, 101030, 101030, 101030, 101020, 101010, 101010, 101030, 
    101040, 101040, 101050, 101050, 101050, 101050, 101070, 101060, 101060, 
    101050, 101060, 101050, 101060, 101070, 101090, 101090, 101090, 101070, 
    101070, 101060, 101060, 101050, 101030, 101040, 101050, 101060, 101080, 
    101070, 101040, 101020, 100990, 100970, 100970, 100960, 100940, 100920, 
    100890, 100890, 100860, 100850, 100820, 100790, 100770, 100750, 100730, 
    100700, 100690, 100680, 100670, 100690, 100680, 100670, 100650, 100640, 
    100620, 100610, 100570, 100560, 100570, 100550, 100550, 100510, 100460, 
    100430, 100390, 100360, 100330, 100340, 100320, 100350, 100310, 100310, 
    100330, 100350, 100340, 100360, 100360, 100350, 100320, 100320, 100330, 
    100340, 100320, 100330, 100340, 100370, 100370, 100380, 100390, 100410, 
    100430, 100430, 100460, 100450, 100460, 100480, 100490, 100470, 100430, 
    100430, 100470, 100460, 100430, 100400, 100370, 100320, 100270, 100230, 
    100200, 100170, 100160, 100140, 100100, 100090, 100070, 100080, 100080, 
    100080, 100100, 100130, 100170, 100210, 100240, 100310, 100350, 100400, 
    100460, 100510, 100560, 100610, 100640, 100650, 100730, 100790, 100850, 
    100930, 100990, 101040, 101070, 101090, 101140, 101150, 101180, 101210, 
    101260, 101290, 101340, 101370, 101390, 101410, 101410, 101410, 101410, 
    101390, 101360, 101400, 101410, 101470, 101500, 101530, 101540, 101540, 
    101500, 101500, 101480, 101490, 101520, 101500, 101500, 101500, 101520, 
    101580, 101620, 101650, 101650, 101590, 101600, 101560, 101580, 101600, 
    101640, 101660, 101660, 101640, 101610, 101610, 101600, 101590, 101590, 
    101580, 101570, 101550, 101580, 101610, 101590, 101590, 101590, 101600, 
    101590, 101600, 101580, 101580, 101590, 101590, 101580, 101600, 101600, 
    101590, 101590, 101580, 101570, 101580, 101560, 101560, 101530, 101510, 
    101530, 101510, 101540, 101520, 101520, 101490, 101460, 101430, 101410, 
    101360, 101340, 101310, 101270, 101250, 101210, 101170, 101120, 101090, 
    101020, 100950, 100920, 100880, 100810, 100790, 100750, 100700, 100660, 
    100650, 100600, 100560, 100490, 100430, 100360, 100310, 100280, 100240, 
    100200, 100160, 100160, 100150, 100120, 100110, 100090, 100090, 100100, 
    100100, 100090, 100100, 100130, 100150, 100170, 100210, 100230, 100250, 
    100270, 100300, 100280, 100280, 100330, 100370, 100410, 100450, 100490, 
    100510, 100520, 100520, 100520, 100550, 100550, 100570, 100600, 100580, 
    100590, 100660, 100720, 100770, 100780, 100780, 100840, 100840, 100840, 
    100860, 100890, 100890, 100890, 100930, 100910, 100910, 100920, 100910, 
    100890, 100860, 100870, 100860, 100880, 100910, 100890, 100900, 100890, 
    100890, 100850, 100810, 100770, 100740, 100700, 100650, 100590, 100540, 
    100450, 100350, 100290, 100180, 100090, 100050, 99960, 99910, 99810, 
    99740, 99730, 99650, 99620, 99620, 99600, 99630, 99640, 99670, 99730, 
    99750, 99820, 99860, 99880, 99890, 99940, 99980, 100010, 100040, 100090, 
    100120, 100140, 100190, 100230, 100260, 100310, 100360, 100420, 100450, 
    100510, 100560, 100580, 100590, 100620, 100640, 100670, 100690, 100720, 
    100730, 100750, 100760, 100800, 100800, 100810, 100800, 100800, 100790, 
    100800, 100810, 100830, 100840, 100860, 100890, 100890, 100920, 100930, 
    100940, 100960, 100970, 100990, 101010, 101020, 101040, 101050, 101060, 
    101060, 101080, 101090, 101100, 101090, 101070, 101080, 101100, 101090, 
    101110, 101110, 101100, 101120, 101140, 101130, 101120, 101120, 101110, 
    101110, 101080, 101050, 101040, 101020, 101020, 101020, 101010, 100990, 
    100990, 100980, 100980, 100970, 100980, 100990, 100990, 101000, 100990, 
    101010, 101020, 101030, 101050, 101050, 101020, 101030, 101060, 101080, 
    101110, 101090, 101080, 101120, 101100, 101080, 101110, 101090, 101020, 
    101070, 101060, 101030, 100990, 100950, 100910, 100880, 100810, 100680, 
    100540, 100430, 100310, 100270, 100120, 99940, 99860, 99650, 99630, 
    99510, 99480, 99540, 99550, 99580, 99590, 99640, 99690, 99750, 99810, 
    99840, 99860, 99880, 99910, 99990, 100040, 100070, 100110, 100160, 
    100250, 100300, 100330, 100400, 100480, 100580, 100640, 100710, 100780, 
    100870, 100960, 101050, 101110, 101170, 101250, 101300, 101370, 101440, 
    101480, 101490, 101500, 101520, 101570, 101590, 101610, 101600, 101610, 
    101600, 101580, 101540, 101570, 101550, 101500, 101470, 101410, 101410, 
    101340, 101260, 101170, 101070, 101010, 100880, 100810, 100700, 100570, 
    100490, 100290, 100390, 100340, 100380, 100340, 100370, 100400, 100420, 
    100460, 100510, 100560, 100600, 100650, 100680, 100710, 100710, 100740, 
    100790, 100850, 100840, 100840, 100840, 100840, 100850, 100870, 100840, 
    100870, 100890, 100910, 100930, 100960, 101050, 101050, 101090, 101180, 
    101180, 101210, 101270, 101300, 101330, 101330, 101380, 101390, 101390, 
    101440, 101420, 101390, 101420, 101410, 101380, 101350, 101330, 101320, 
    101320, 101330, 101310, 101300, 101220, 101140, 101020, 101020, 100950, 
    100910, 100900, 100810, 100770, 100750, 100680, 100670, 100620, 100620, 
    100650, 100650, 100660, 100660, 100660, 100690, 100690, 100710, 100740, 
    100780, 100850, 100900, 100910, 100890, 100900, 100970, 101010, 101030, 
    101030, 101040, 101030, 100990, 100970, 100910, 100830, 100740, 100690, 
    100670, 100660, 100640, 100630, 100610, 100630, 100660, 100680, 100700, 
    100730, 100750, 100780, 100810, 100880, 100910, 100990, 101020, 101070, 
    101140, 101200, 101260, 101310, 101360, 101410, 101480, 101510, 101570, 
    101640, 101690, 101740, 101790, 101840, 101870, 101900, 101910, 101920, 
    101840, 101890, 101890, 101870, 101870, 101850, 101820, 101780, 101730, 
    101650, 101600, 101560, 101470, 101420, 101370, 101290, 101200, 101150, 
    101090, 101030, 101040, 101030, 101060, 101080, 101140, 101200, 101260, 
    101360, 101420, 101500, 101550, 101600, 101600, 101650, 101650, 101740, 
    101770, 101810, 101820, 101860, 101850, 101860, 101830, 101830, 101790, 
    101770, 101760, 101750, 101710, 101680, 101670, 101670, 101660, 101640, 
    101670, 101640, 101610, 101580, 101540, 101510, 101500, 101500, 101460, 
    101440, 101420, 101410, 101350, 101390, 101380, 101380, 101370, 101350, 
    101340, 101300, 101320, 101330, 101380, 101410, 101440, 101460, 101470, 
    101480, 101510, 101530, 101550, 101570, 101590, 101610, 101610, 101620, 
    101660, 101670, 101670, 101670, 101650, 101640, 101640, 101650, 101610, 
    101590, 101580, 101560, 101560, 101510, 101480, 101450, 101420, 101370, 
    101350, 101320, 101280, 101280, 101250, 101200, 101190, 101150, 101110, 
    101050, 101020, 100990, 100980, 100930, 100870, 100870, 100820, 100820, 
    100800, 100780, 100750, 100700, 100680, 100630, 100600, 100570, 100550, 
    100540, 100530, 100530, 100510, 100510, 100500, 100490, 100480, 100500, 
    100510, 100520, 100530, 100550, 100590, 100630, 100620, 100630, 100650, 
    100670, 100700, 100720, 100710, 100730, 100770, 100750, 100780, 100750, 
    100750, 100870, 100920, 100930, 100940, 100910, 100910, 100920, 101040, 
    101060, 101050, 101080, 101120, 101170, 101170, 101150, 101220, 101220, 
    101270, 101310, 101340, 101370, 101390, 101330, 101330, 101320, 101340, 
    101320, 101320, 101310, 101290, 101290, 101280, 101270, 101260, 101250, 
    101240, 101230, 101200, 101200, 101190, 101180, 101180, 101170, 101190, 
    101150, 101130, 101130, 101140, 101130, 101110, 101050, 101010, 100960, 
    100900, 100880, 100880, 100860, 100850, 100830, 100810, 100750, 100740, 
    100710, 100690, 100660, 100670, 100690, 100690, 100730, 100740, 100740, 
    100740, 100700, 100730, 100750, 100810, 100790, 100740, 100770, 100780, 
    100820, 100850, 100860, 100860, 100860, 100830, 100820, 100820, 100780, 
    100800, 100790, 100790, 100800, 100780, 100800, 100800, 100790, 100750, 
    100750, 100740, 100750, 100750, 100750, 100760, 100770, 100800, 100820, 
    100840, 100840, 100840, 100830, 100850, 100860, 100890, 100910, 100930, 
    100980, 101000, 101020, 101040, 101010, 101000, 101000, 101000, 101000, 
    100970, 100970, 100980, 100980, 100960, 100990, 100990, 100980, 100990, 
    100990, 100980, 100980, 100990, 101020, 101030, 101060, 101050, 101070, 
    101050, 101060, 101040, 101040, 101040, 101040, 101060, 101070, 101100, 
    101120, 101160, 101170, 101200, 101210, 101220, 101220, 101220, 101220, 
    101210, 101220, 101220, 101230, 101230, 101230, 101220, 101230, 101200, 
    101200, 101200, 101190, 101190, 101160, 101210, 101220, 101230, 101250, 
    101280, 101290, 101310, 101330, 101340, 101370, 101410, 101430, 101470, 
    101490, 101520, 101550, 101590, 101600, 101620, 101630, 101630, 101640, 
    101660, 101680, 101710, 101730, 101730, 101760, 101770, 101780, 101790, 
    101780, 101780, 101760, 101750, 101730, 101730, 101710, 101710, 101720, 
    101700, 101700, 101680, 101670, 101670, 101640, 101630, 101620, 101610, 
    101600, 101610, 101610, 101640, 101640, 101660, 101660, 101650, 101640, 
    101640, 101610, 101590, 101590, 101600, 101600, 101620, 101610, 101620, 
    101620, 101600, 101600, 101590, 101590, 101620, 101660, 101710, 101760, 
    101800, 101810, 101860, 101880, 101910, 101920, 101940, 101950, 101960, 
    101990, 102000, 102030, 102060, 102090, 102110, 102120, 102140, 102150, 
    102170, 102160, 102200, 102210, 102230, 102260, 102270, 102260, 102240, 
    102220, 102230, 102210, 102200, 102190, 102160, 102190, 102190, 102160, 
    102160, 102120, 102080, 102060, 102020, 101990, 101970, 101950, 101960, 
    101960, 101960, 101960, 101940, 101970, 101960, 101950, 101940, 101940, 
    101950, 101960, 101940, 101940, 101940, 101940, 101940, 101930, 101910, 
    101870, 101850, 101840, 101830, 101830, 101840, 101810, 101830, 101840, 
    101810, 101790, 101750, 101730, 101700, 101680, 101630, 101620, 101590, 
    101540, 101500, 101470, 101440, 101390, 101360, 101330, 101300, 101290, 
    101270, 101230, 101240, 101210, 101210, 101200, 101170, 101130, 101090, 
    101070, 101070, 101020, 100990, 100970, 100970, 100950, 100920, 100880, 
    100850, 100880, 100790, 100750, 100790, 100770, 100740, 100770, 100760, 
    100670, 100680, 100620, 100610, 100600, 100570, 100570, 100520, 100510, 
    100410, 100390, 100360, 100310, 100210, 100150, 100130, 100110, 100080, 
    99990, 99950, 99910, 99840, 99840, 99810, 99710, 99700, 99680, 99680, 
    99620, 99560, 99530, 99460, 99400, 99300, 99380, 99410, 99430, 99390, 
    99360, 99320, 99300, 99270, 99230, 99190, 99180, 99170, 99160, 99130, 
    99130, 99140, 99140, 99160, 99190, 99230, 99200, 99260, 99260, 99230, 
    99280, 99310, 99350, 99350, 99380, 99400, 99420, 99450, 99450, 99430, 
    99450, 99470, 99500, 99520, 99560, 99540, 99600, 99650, 99660, 99690, 
    99690, 99720, 99760, 99840, 99910, 99950, 99990, 100070, 100150, 100240, 
    100290, 100350, 100380, 100380, 100380, 100370, 100380, 100390, 100390, 
    100380, 100350, 100330, 100310, 100320, 100340, 100350, 100360, 100380, 
    100470, 100510, 100550, 100580, 100600, 100580, 100590, 100640, 100660, 
    100680, 100630, 100710, 100770, 100800, 100800, 100800, 100840, 100920, 
    100900, 100920, 100930, 100940, 100960, 100990, 101030, 101040, 101090, 
    101100, 101080, 101060, 101030, 101050, 101020, 100980, 100970, 100960, 
    100960, 100970, 100970, 100960, 100970, 100960, 100950, 100950, 100950, 
    100900, 100870, 100840, 100820, 100780, 100760, 100750, 100760, 100750, 
    100770, 100790, 100790, 100800, 100800, 100820, 100830, 100810, 100840, 
    100850, 100850, 100850, 100840, 100840, 100810, 100750, 100730, 100720, 
    100660, 100640, 100600, 100570, 100530, 100500, 100450, 100460, 100450, 
    100420, 100390, 100350, 100320, 100310, 100320, 100330, 100330, 100350, 
    100340, 100320, 100300, 100290, 100280, 100290, 100280, 100230, 100280, 
    100300, 100330, 100340, 100390, 100490, 100600, 100690, 100760, 100830, 
    100890, 100940, 101030, 101100, 101160, 101220, 101270, 101310, 101330, 
    101370, 101380, 101400, 101440, 101470, 101500, 101530, 101560, 101590, 
    101620, 101630, 101630, 101610, 101620, 101620, 101630, 101630, 101620, 
    101630, 101670, 101690, 101720, 101740, 101760, 101760, 101770, 101770, 
    101780, 101780, 101790, 101780, 101790, 101790, 101780, 101780, 101780, 
    101760, 101730, 101740, 101750, 101780, 101770, 101780, 101770, 101750, 
    101760, 101730, 101710, 101670, 101640, 101620, 101610, 101560, 101530, 
    101490, 101470, 101460, 101460, 101420, 101410, 101370, 101350, 101330, 
    101330, 101320, 101310, 101300, 101280, 101240, 101240, 101240, 101200, 
    101140, 101120, 101100, 101050, 101020, 100970, 100940, 100950, 100950, 
    100900, 100860, 100820, 100790, 100740, 100690, 100670, 100630, 100610, 
    100550, 100490, 100430, 100380, 100310, 100250, 100240, 100250, 100240, 
    100250, 100270, 100290, 100330, 100390, 100420, 100470, 100480, 100510, 
    100540, 100560, 100580, 100590, 100630, 100670, 100700, 100740, 100750, 
    100740, 100700, 100720, 100710, 100690, 100660, 100660, 100630, 100600, 
    100580, 100540, 100510, 100460, 100410, 100330, 100240, 100100, 100030, 
    99980, 99980, 99950, 99980, 99990, 100020, 100030, 100020, 100000, 99990, 
    99970, 99950, 99910, 99880, 99830, 99800, 99750, 99740, 99730, 99730, 
    99710, 99690, 99670, 99640, 99640, 99650, 99640, 99650, 99650, 99660, 
    99690, 99700, 99690, 99680, 99640, 99620, 99610, 99610, 99600, 99580, 
    99550, 99510, 99480, 99420, 99330, 99250, 99200, 99160, 99100, 99020, 
    98960, 98940, 98890, 98900, 98880, 98860, 98860, 98870, 98900, 98900, 
    98900, 98950, 98960, 98980, 99010, 99050, 99050, 99100, 99110, 99150, 
    99180, 99210, 99270, 99320, 99400, 99390, 99460, 99510, 99580, 99660, 
    99710, 99810, 99860, 99870, 99920, 99990, 100060, 100100, 100220, 100320, 
    100360, 100430, 100470, 100470, 100500, 100570, 100600, 100620, 100630, 
    100690, 100710, 100730, 100760, 100770, 100790, 100790, 100810, 100820, 
    100830, 100840, 100840, 100880, 100880, 100910, 100920, 100940, 100950, 
    100970, 100980, 101010, 101030, 101040, 101090, 101110, 101140, 101150, 
    101150, 101150, 101140, 101140, 101140, 101140, 101150, 101140, 101120, 
    101120, 101120, 101110, 101090, 101050, 101010, 100990, 100980, 100910, 
    100880, 100830, 100790, 100750, 100660, 100550, 100420, 100390, 100280, 
    100210, 100080, 99990, 99910, 99810, 99830, 99780, 99790, 99860, 99920, 
    99990, 100060, 100200, 100260, 100330, 100410, 100480, 100570, 100660, 
    100730, 100800, 100840, 100880, 100940, 100990, 101030, 101090, 101160, 
    101250, 101290, 101320, 101420, 101400, 101480, 101520, 101520, 101570, 
    101670, 101750, 101860, 101960, 102050, 102130, 102180, 102210, 102290, 
    102340, 102390, 102420, 102490, 102480, 102530, 102560, 102570, 102610, 
    102630, 102650, 102650, 102650, 102650, 102670, 102660, 102660, 102650, 
    102670, 102680, 102670, 102670, 102670, 102650, 102650, 102640, 102630, 
    102600, 102590, 102550, 102580, 102580, 102580, 102580, 102550, 102510, 
    102480, 102500, 102490, 102460, 102440, 102440, 102440, 102420, 102390, 
    102370, 102330, 102300, 102310, 102300, 102290, 102250, 102220, 102190, 
    102200, 102200, 102190, 102180, 102170, 102160, 102180, 102160, 102100, 
    102110, 102110, 102090, 102080, 102100, 102080, 102090, 102100, 102100, 
    102100, 102110, 102110, 102130, 102140, 102140, 102140, 102180, 102180, 
    102180, 102170, 102170, 102160, 102150, 102150, 102140, 102140, 102130, 
    102160, 102180, 102180, 102190, 102240, 102260, 102230, 102220, 102210, 
    102210, 102210, 102190, 102190, 102150, 102160, 102180, 102180, 102160, 
    102150, 102160, 102150, 102110, 102100, 102110, 102120, 102110, 102110, 
    102130, 102120, 102100, 102080, 102110, 102090, 102080, 102060, 102060, 
    102050, 102050, 102070, 102090, 102100, 102080, 102060, 102050, 102030, 
    102010, 102020, 102020, 102010, 102030, 102020, 102050, 102050, 102050, 
    102050, 102060, 101990, 101980, 101940, 101930, 101950, 101920, 101920, 
    101930, 101980, 101970, 101980, 101990, 101990, 101940, 101940, 101960, 
    101980, 102010, 102030, 102050, 102070, 102070, 102070, 102020, 102030, 
    102030, 102060, 102110, 102130, 102150, 102140, 102150, 102180, 102180, 
    102180, 102190, 102230, 102230, 102260, 102270, 102290, 102320, 102360, 
    102380, 102360, 102370, 102410, 102380, 102420, 102460, 102500, 102550, 
    102550, 102540, 102570, 102580, 102570, 102580, 102540, 102590, 102610, 
    102620, 102620, 102630, 102620, 102610, 102590, 102570, 102570, 102550, 
    102540, 102500, 102470, 102490, 102450, 102450, 102430, 102420, 102400, 
    102380, 102370, 102330, 102310, 102290, 102270, 102240, 102250, 102230, 
    102190, 102180, 102190, 102190, 102130, 102100, 102070, 102060, 102060, 
    101990, 101980, 101950, 101920, 101880, 101850, 101820, 101780, 101770, 
    101710, 101680, 101670, 101650, 101590, 101580, 101540, 101500, 101470, 
    101480, 101410, 101390, 101340, 101280, 101210, 101140, 101100, 101040, 
    100980, 100930, 100900, 100870, 100860, 100830, 100790, 100750, 100740, 
    100760, 100780, 100800, 100830, 100880, 100930, 100990, 101020, 101050, 
    101130, 101170, 101230, 101310, 101370, 101400, 101440, 101500, 101540, 
    101560, 101590, 101600, 101640, 101670, 101640, 101620, 101600, 101520, 
    101440, 101380, 101390, 101290, 101220, 101190, 101150, 101150, 101060, 
    100990, 100890, 100910, 100870, 100860, 100890, 100890, 100920, 101000, 
    100990, 101010, 101000, 101020, 101020, 101030, 101090, 101170, 101260, 
    101360, 101510, 101590, 101730, 101830, 101910, 102010, 102140, 102240, 
    102310, 102380, 102440, 102570, 102650, 102720, 102750, 102820, 102860, 
    102880, 102940, 102980, 102970, 103030, 103080, 103100, 103140, 103170, 
    103170, 103150, 103160, 103170, 103160, 103130, 103120, 103080, 103060, 
    103050, 103020, 102970, 102930, 102900, 102890, 102850, 102850, 102830, 
    102840, 102820, 102820, 102830, 102840, 102850, 102860, 102850, 102840, 
    102800, 102820, 102790, 102770, 102740, 102710, 102650, 102600, 102540, 
    102470, 102390, 102310, 102230, 102150, 102100, 102040, 101990, 101920, 
    101870, 101810, 101780, 101730, 101670, 101640, 101560, 101550, 101520, 
    101520, 101490, 101510, 101520, 101510, 101510, 101530, 101500, 101480, 
    101430, 101420, 101350, 101320, 101260, 101170, 101110, 101060, 100940, 
    100920, 100790, 100770, 100720, 100700, 100700, 100700, 100670, 100680, 
    100740, 100830, 100960, 101090, 101210, 101350, 101510, 101670, 101780, 
    101900, 102050, 102140, 102250, 102370, 102440, 102530, 102600, 102680, 
    102730, 102780, 102860, 102890, 102940, 102960, 102990, 102960, 102930, 
    102920, 102880, 102880, 102800, 102710, 102620, 102580, 102520, 102460, 
    102380, 102280, 102240, 102130, 102070, 101990, 101920, 101820, 101770, 
    101700, 101660, 101630, 101590, 101570, 101540, 101480, 101470, 101480, 
    101530, 101540, 101550, 101590, 101650, 101720, 101720, 101750, 101750, 
    101840, 101880, 101950, 101990, 102030, 102040, 102050, 102060, 102030, 
    102050, 102020, 102010, 101990, 101950, 101980, 101990, 102020, 102040, 
    102080, 102140, 102190, 102210, 102240, 102300, 102330, 102360, 102370, 
    102370, 102420, 102430, 102450, 102450, 102490, 102460, 102450, 102430, 
    102370, 102400, 102310, 102330, 102350, 102340, 102390, 102380, 102390, 
    102420, 102440, 102450, 102470, 102490, 102500, 102520, 102550, 102510, 
    102540, 102510, 102490, 102500, 102520, 102540, 102520, 102520, 102510, 
    102530, 102500, 102510, 102510, 102540, 102530, 102520, 102500, 102490, 
    102440, 102440, 102430, 102400, 102380, 102350, 102300, 102330, 102300, 
    102300, 102310, 102320, 102300, 102320, 102320, 102290, 102260, 102350, 
    102360, 102360, 102430, 102420, 102460, 102470, 102500, 102480, 102510, 
    102570, 102590, 102590, 102630, 102630, 102640, 102660, 102670, 102660, 
    102690, 102690, 102710, 102720, 102710, 102660, 102660, 102630, 102600, 
    102590, 102550, 102500, 102550, 102570, 102480, 102410, 102410, 102370, 
    102290, 102310, 102270, 102220, 102160, 102140, 102140, 102090, 102030, 
    102020, 102030, 102000, 101990, 102000, 101990, 101920, 101860, 101790, 
    101760, 101690, 101650, 101590, 101510, 101430, 101380, 101320, 101260, 
    101190, 101130, 101040, 100950, 100910, 100860, 100790, 100740, 100710, 
    100690, 100640, 100600, 100570, 100510, 100470, 100430, 100390, 100350, 
    100300, 100230, 100190, 100170, 100170, 100130, 100090, 100050, 100020, 
    100020, 100010, 100010, 99990, 99970, 99980, 99980, 99990, 100010, 
    100030, 100040, 100040, 100060, 100070, 100070, 100070, 100060, 100100, 
    100100, 100120, 100160, 100180, 100190, 100220, 100240, 100260, 100250, 
    100280, 100270, 100310, 100350, 100400, 100470, 100530, 100560, 100560, 
    100580, 100610, 100640, 100680, 100700, 100710, 100760, 100800, 100830, 
    100860, 100900, 100920, 100960, 100960, 100980, 101020, 101040, 101060, 
    101060, 101090, 101110, 101150, 101170, 101210, 101240, 101230, 101200, 
    101220, 101250, 101250, 101270, 101300, 101300, 101340, 101350, 101340, 
    101340, 101360, 101400, 101400, 101400, 101400, 101410, 101420, 101420, 
    101420, 101420, 101420, 101450, 101450, 101460, 101470, 101460, 101450, 
    101450, 101470, 101490, 101520, 101520, 101520, 101520, 101530, 101530, 
    101530, 101540, 101540, 101550, 101580, 101600, 101620, 101650, 101680, 
    101690, 101700, 101720, 101720, 101730, 101730, 101720, 101730, 101760, 
    101760, 101750, 101740, 101730, 101740, 101730, 101740, 101740, 101730, 
    101720, 101710, 101710, 101710, 101690, 101670, 101630, 101600, 101580, 
    101530, 101540, 101530, 101530, 101520, 101510, 101540, 101550, 101550, 
    101570, 101590, 101600, 101600, 101590, 101610, 101600, 101590, 101590, 
    101600, 101590, 101570, 101550, 101550, 101560, 101570, 101580, 101560, 
    101590, 101620, 101640, 101660, 101690, 101680, 101710, 101720, 101710, 
    101720, 101750, 101740, 101730, 101730, 101760, 101750, 101740, 101740, 
    101740, 101730, 101690, 101730, 101740, 101720, 101730, 101740, 101760, 
    101740, 101760, 101760, 101750, 101750, 101770, 101790, 101790, 101800, 
    101830, 101850, 101880, 101920, 101920, 101930, 101950, 101950, 101960, 
    102000, 102030, 102030, 102030, 102050, 102040, 102040, 102050, 102060, 
    102060, 102050, 102090, 102090, 102110, 102130, 102140, 102150, 102160, 
    102170, 102160, 102140, 102140, 102140, 102140, 102120, 102110, 102110, 
    102100, 102080, 102090, 102080, 102080, 102070, 102070, 102070, 102050, 
    102050, 102050, 102050, 102050, 102030, 102050, 102050, 102030, 102010, 
    102030, 102000, 101970, 101860, 101890, 101950, 102000, 102030, 102060, 
    102080, 102080, 102080, 102020, 102050, 102020, 102000, 101960, 101960, 
    101980, 102010, 102030, 102050, 102070, 102060, 102030, 102010, 102010, 
    102000, 101980, 101990, 102000, 101960, 101910, 101910, 101850, 101800, 
    101770, 101740, 101700, 101650, 101620, 101590, 101580, 101550, 101560, 
    101550, 101540, 101540, 101560, 101550, 101550, 101540, 101520, 101550, 
    101570, 101590, 101600, 101610, 101630, 101660, 101660, 101660, 101660, 
    101650, 101630, 101630, 101670, 101710, 101740, 101760, 101790, 101810, 
    101810, 101830, 101860, 101870, 101890, 101920, 101950, 101980, 101990, 
    102010, 102020, 102030, 102030, 102050, 102060, 102070, 102100, 102110, 
    102130, 102150, 102160, 102170, 102150, 102180, 102180, 102180, 102160, 
    102150, 102140, 102140, 102150, 102160, 102170, 102160, 102140, 102110, 
    102110, 102110, 102100, 102110, 102060, 102060, 102050, 102040, 102020, 
    102000, 101970, 101950, 101950, 101930, 101920, 101910, 101890, 101860, 
    101840, 101830, 101840, 101840, 101790, 101760, 101720, 101740, 101750, 
    101740, 101710, 101730, 101710, 101750, 101740, 101780, 101790, 101800, 
    101820, 101850, 101830, 101860, 101880, 101890, 101930, 101940, 101940, 
    101960, 101970, 101980, 101990, 101990, 101990, 102010, 101990, 102010, 
    102020, 102050, 102060, 102050, 102050, 102070, 102080, 102060, 102100, 
    102090, 102100, 102090, 102100, 102090, 102070, 102060, 102040, 102000, 
    101980, 101940, 101930, 101880, 101880, 101790, 101750, 101740, 101680, 
    101570, 101450, 101380, 101260, 101210, 101140, 101090, 101020, 100950, 
    100930, 100850, 100780, 100710, 100670, 100620, 100560, 100540, 100550, 
    100540, 100540, 100550, 100550, 100580, 100570, 100530, 100510, 100490, 
    100430, 100460, 100480, 100500, 100540, 100530, 100560, 100570, 100570, 
    100590, 100650, 100660, 100690, 100740, 100780, 100800, 100800, 100840, 
    100870, 100890, 100930, 100950, 100970, 100980, 100970, 100900, 100870, 
    100860, 100850, 100820, 100810, 100830, 100790, 100740, 100740, 100730, 
    100700, 100700, 100710, 100710, 100670, 100680, 100660, 100670, 100670, 
    100700, 100700, 100710, 100690, 100680, 100680, 100660, 100650, 100680, 
    100680, 100670, 100650, 100660, 100630, 100620, 100610, 100560, 100550, 
    100510, 100480, 100420, 100400, 100340, 100340, 100310, 100280, 100240, 
    100160, 100100, 100060, 100010, 99960, 99890, 99820, 99770, 99700, 99650, 
    99590, 99540, 99470, 99410, 99340, 99270, 99240, 99190, 99080, 99100, 
    99070, 99000, 98990, 98940, 98900, 98890, 98850, 98710, 98650, 98670, 
    98670, 98630, 98580, 98510, 98480, 98450, 98400, 98350, 98330, 98280, 
    98220, 98280, 98220, 98270, 98260, 98160, 98140, 98110, 98120, 98080, 
    98150, 98230, 98300, 98360, 98440, 98500, 98530, 98560, 98590, 98610, 
    98680, 98660, 98640, 98690, 98710, 98760, 98750, 98760, 98800, 98800, 
    98770, 98770, 98820, 98840, 98860, 98930, 98960, 98960, 99000, 99010, 
    99020, 99070, 99080, 99070, 99070, 99070, 99110, 99120, 99140, 99190, 
    99200, 99190, 99180, 99150, 99070, 99020, 98950, 98910, 98910, 98890, 
    98820, 98880, 98870, 98940, 98960, 98990, 98960, 98990, 98990, 99010, 
    99010, 99030, 99010, 99010, 99040, 99030, 99040, 99080, 99090, 99090, 
    99110, 99130, 99130, 99150, 99170, 99170, 99200, 99210, 99230, 99240, 
    99260, 99270, 99300, 99310, 99330, 99350, 99380, 99400, 99430, 99460, 
    99480, 99500, 99500, 99520, 99500, 99490, 99500, 99510, 99500, 99500, 
    99500, 99480, 99480, 99480, 99440, 99420, 99410, 99390, 99370, 99340, 
    99320, 99300, 99260, 99240, 99220, 99210, 99170, 99130, 99080, 99020, 
    98940, 98890, 98810, 98800, 98760, 98730, 98680, 98670, 98660, 98650, 
    98660, 98660, 98610, 98610, 98640, 98590, 98620, 98590, 98580, 98500, 
    98460, 98430, 98420, 98440, 98480, 98490, 98520, 98540, 98560, 98610, 
    98660, 98690, 98740, 98810, 98960, 98960, 99060, 99160, 99250, 99340, 
    99390, 99440, 99460, 99480, 99530, 99590, 99590, 99600, 99610, 99620, 
    99620, 99630, 99640, 99720, 99850, 99880, 99900, 99950, 99980, 100040, 
    100090, 100150, 100170, 100220, 100290, 100330, 100400, 100430, 100490, 
    100540, 100560, 100650, 100700, 100760, 100790, 100830, 100870, 100920, 
    100960, 101020, 101040, 101080, 101120, 101160, 101200, 101210, 101250, 
    101290, 101330, 101380, 101400, 101440, 101480, 101500, 101530, 101560, 
    101580, 101590, 101630, 101650, 101670, 101730, 101760, 101780, 101810, 
    101820, 101840, 101880, 101910, 101910, 101950, 101980, 102030, 102080, 
    102080, 102130, 102190, 102220, 102250, 102300, 102320, 102360, 102370, 
    102410, 102440, 102480, 102490, 102510, 102510, 102520, 102510, 102520, 
    102520, 102510, 102530, 102480, 102480, 102480, 102450, 102420, 102400, 
    102350, 102310, 102270, 102230, 102220, 102170, 102120, 102090, 102060, 
    102010, 101920, 101870, 101790, 101730, 101690, 101690, 101670, 101630, 
    101620, 101600, 101580, 101570, 101560, 101540, 101510, 101480, 101420, 
    101390, 101330, 101240, 101170, 101100, 101130, 101140, 101160, 101230, 
    101290, 101190, 101180, 101290, 101330, 101360, 101370, 101340, 101260, 
    101280, 101240, 101270, 101410, 101470, 101430, 101410, 101360, 101320, 
    101250, 101190, 101220, 101250, 101180, 101140, 101120, 101060, 100960, 
    100900, 100840, 100880, 100850, 100860, 100870, 100870, 100870, 100850, 
    100800, 100730, 100690, 100660, 100730, 100660, 100550, 100510, 100380, 
    100510, 100580, 100570, 100550, 100550, 100510, 100430, 100300, 100300, 
    100330, 100350, 100400, 100420, 100430, 100480, 100470, 100470, 100470, 
    100430, 100410, 100400, 100330, 100260, 100240, 100250, 100290, 100310, 
    100350, 100390, 100450, 100480, 100520, 100550, 100570, 100640, 100630, 
    100660, 100670, 100670, 100700, 100710, 100700, 100690, 100650, 100650, 
    100690, 100700, 100720, 100740, 100750, 100730, 100700, 100730, 100750, 
    100770, 100780, 100820, 100860, 100890, 100920, 100930, 100970, 101000, 
    101030, 101040, 101100, 101120, 101160, 101210, 101290, 101310, 101300, 
    101280, 101310, 101310, 101300, 101330, 101380, 101320, 101340, 101410, 
    101470, 101480, 101520, 101580, 101640, 101650, 101700, 101750, 101740, 
    101730, 101700, 101660, 101800, 101820, 101810, 101820, 101840, 101850, 
    101840, 101840, 101830, 101850, 101870, 101890, 101900, 101880, 101940, 
    101950, 101950, 101940, 101980, 101950, 102020, 101970, 101960, 102000, 
    102020, 102020, 102030, 102020, 102000, 101980, 101960, 101950, 101950, 
    101930, 101900, 101880, 101830, 101810, 101870, 101880, 101870, 101870, 
    101750, 101880, 101940, 102020, 102030, 102020, 102040, 102080, 102100, 
    102140, 102160, 102160, 102180, 102180, 102220, 102220, 102210, 102230, 
    102250, 102260, 102330, 102360, 102370, 102380, 102340, 102420, 102430, 
    102430, 102440, 102440, 102360, 102430, 102450, 102490, 102490, 102510, 
    102520, 102540, 102550, 102550, 102570, 102580, 102600, 102620, 102660, 
    102720, 102760, 102780, 102800, 102820, 102850, 102870, 102880, 102890, 
    102900, 102940, 102980, 102980, 103010, 103010, 103010, 103110, 103140, 
    103120, 103140, 103190, 103210, 103250, 103360, 103410, 103330, 103540, 
    103520, 103510, 103580, 103600, 103630, 103650, 103670, 103720, 103770, 
    103800, 103870, 103870, 103900, 103890, 103900, 103910, 103950, 103950, 
    103970, 103960, 103950, 103980, 104010, 104110, 104100, 104050, 104080, 
    104100, 104130, 104100, 104140, 104110, 104140, 104150, 104100, 104090, 
    104170, 104180, 104230, 104250, 104230, 104220, 104210, 104210, 104230, 
    104260, 104280, 104270, 104280, 104240, 104260, 104280, 104280, 104280, 
    104280, 104290, 104310, 104290, 104300, 104320, 104320, 104320, 104310, 
    104340, 104330, 104300, 104280, 104270, 104260, 104260, 104230, 104180, 
    104160, 104100, 104080, 104060, 104020, 104000, 103970, 103920, 103890, 
    103850, 103810, 103790, 103740, 103680, 103610, 103590, 103560, 103530, 
    103490, 103470, 103450, 103440, 103400, 103350, 103310, 103270, 103230, 
    103200, 103180, 103170, 103130, 103040, 102990, 102950, 102920, 102850, 
    102800, 102750, 102710, 102650, 102580, 102530, 102470, 102420, 102370, 
    102350, 102280, 102230, 102170, 102090, 102000, 101940, 101880, 101820, 
    101760, 101690, 101630, 101550, 101480, 101410, 101330, 101270, 101180, 
    101080, 101010, 100940, 100860, 100790, 100730, 100660, 100610, 100550, 
    100460, 100380, 100350, 100350, 100330, 100330, 100330, 100340, 100340, 
    100340, 100330, 100350, 100330, 100310, 100270, 100260, 100260, 100280, 
    100320, 100320, 100320, 100330, 100340, 100280, 100290, 100320, 100350, 
    100370, 100460, 100530, 100550, 100560, 100570, 100570, 100630, 100630, 
    100610, 100650, 100660, 100630, 100680, 100680, 100700, 100790, 101020, 
    101070, 101100, 101140, 101160, 101180, 101230, 101260, 101250, 101270, 
    101310, 101310, 101290, 101270, 101340, 101330, 101320, 101290, 101280, 
    101260, 101220, 101240, 101240, 101220, 101240, 101290, 101270, 101270, 
    101260, 101270, 101290, 101320, 101340, 101340, 101390, 101390, 101410, 
    101420, 101430, 101420, 101410, 101340, 101350, 101360, 101340, 101330, 
    101310, 101300, 101300, 101300, 101310, 101330, 101300, 101270, 101240, 
    101250, 101230, 101210, 101210, 101200, 101190, 101170, 101150, 101080, 
    101020, 100930, 100820, 100760, 100630, 100450, 100260, 100100, 99890, 
    99690, 99480, 99340, 99330, 99360, 99350, 99340, 99320, 99290, 99320, 
    99340, 99390, 99420, 99480, 99510, 99540, 99550, 99560, 99580, 99560, 
    99550, 99520, 99490, 99440, 99400, 99390, 99380, 99320, 99280, 99250, 
    99240, 99240, 99260, 99270, 99300, 99300, 99300, 99290, 99320, 99340, 
    99390, 99410, 99440, 99440, 99410, 99430, 99440, 99460, 99480, 99400, 
    99420, 99410, 99460, 99530, 99600, 99670, 99730, 99780, 99850, 99870, 
    99910, 99960, 99970, 100000, 99980, 99970, 99950, 100030, 100030, 100060, 
    100080, 100140, 100210, 100210, 100310, 100350, 100410, 100450, 100460, 
    100500, 100520, 100550, 100560, 100550, 100570, 100560, 100570, 100540, 
    100540, 100550, 100530, 100530, 100570, 100590, 100650, 100690, 100640, 
    100700, 100700, 100740, 100760, 100720, 100810, 100780, 100790, 100800, 
    100820, 100800, 100690, 100750, 100710, 100840, 100850, 100910, 101030, 
    101040, 101000, 101100, 101150, 101180, 101220, 101240, 101260, 101310, 
    101370, 101390, 101380, 101440, 101460, 101470, 101550, 101550, 101550, 
    101530, 101590, 101550, 101610, 101630, 101610, 101630, 101600, 101600, 
    101640, 101630, 101570, 101540, 101580, 101540, 101690, 101770, 101810, 
    101820, 101810, 101850, 101900, 101920, 101940, 101960, 101980, 102000, 
    102020, 102030, 102050, 102020, 102020, 102010, 102100, 102160, 102170, 
    102230, 102250, 102260, 102250, 102290, 102340, 102340, 102390, 102360, 
    102380, 102390, 102430, 102440, 102460, 102470, 102470, 102460, 102450, 
    102440, 102420, 102420, 102400, 102400, 102430, 102400, 102370, 102330, 
    102270, 102250, 102240, 102230, 102220, 102180, 102110, 102130, 102100, 
    102080, 102050, 102000, 101980, 101980, 101950, 101920, 101900, 101870, 
    101860, 101840, 101840, 101830, 101800, 101730, 101730, 101730, 101720, 
    101730, 101760, 101770, 101770, 101780, 101770, 101760, 101760, 101710, 
    101740, 101680, 101670, 101700, 101710, 101680, 101680, 101710, 101720, 
    101690, 101670, 101690, 101670, 101660, 101630, 101630, 101580, 101550, 
    101490, 101460, 101390, 101390, 101340, 101310, 101230, 101180, 101150, 
    101120, 101080, 101020, 100940, 100910, 100890, 100780, 100680, 100620, 
    100530, 100430, 100340, 100160, 100290, 99980, 99920, 99870, 99660, 
    99650, 99620, 99570, 99500, 99560, 99450, 99410, 99400, 99390, 99440, 
    99460, 99540, 99580, 99620, 99650, 99680, 99700, 99740, 99780, 99840, 
    99860, 99880, 99880, 99750, 99690, 99700, 99700, 99690, 99710, 99740, 
    99700, 99870, 100040, 100050, 100040, 100070, 100070, 100070, 100060, 
    100040, 100020, 99990, 99960, 99930, 99940, 99980, 99980, 99960, 99920, 
    99940, 99960, 100000, 100190, 100220, 100250, 100240, 100260, 100310, 
    100290, 100140, 100120, 100250, 100270, 100300, 100330, 100330, 100100, 
    100050, 100030, 100080, 100140, 100220, 100300, 100270, 100300, 100350, 
    100380, 100370, 100400, 100400, 100410, 100400, 100420, 100460, 100480, 
    100450, 100430, 100430, 100460, 100450, 100430, 100370, 100380, 100340, 
    100330, 100340, 100350, 100330, 100310, 100320, 100320, 100260, 100290, 
    100260, 100250, 100260, 100220, 100200, 100140, 100130, 100080, 100040, 
    99980, 99990, 100020, 100040, 100070, 100110, 100090, 100120, 100140, 
    100150, 100170, 100180, 100180, 100170, 100180, 100180, 100210, 100240, 
    100250, 100260, 100290, 100320, 100340, 100370, 100450, 100480, 100490, 
    100520, 100530, 100560, 100580, 100590, 100600, 100640, 100610, 100600, 
    100580, 100530, 100500, 100450, 100410, 100400, 100340, 100300, 100280, 
    100270, 100160, 100010, 99870, 99720, 99500, 99350, 99150, 98960, 98750, 
    98550, 98350, 98100, 97820, 97560, 97270, 96990, 96720, 96590, 96550, 
    96530, 96500, 96480, 96450, 96360, 96290, 96220, 96200, 96200, 96230, 
    96260, 96250, 96250, 96230, 96240, 96220, 96300, 96390, 96470, 96570, 
    96670, 96740, 96810, 96880, 96940, 97050, 97180, 97310, 97390, 97470, 
    97520, 97570, 97580, 97670, 97700, 97830, 97960, 98040, 98160, 98250, 
    98330, 98410, 98520, 98610, 98700, 98790, 98800, 98880, 98920, 98910, 
    98920, 98780, 98810, 98840, 98870, 98920, 98970, 98940, 98950, 99000, 
    99080, 99110, 99130, 99120, 99200, 99210, 99250, 99230, 99270, 99350, 
    99420, 99510, 99580, 99640, 99680, 99760, 99810, 99860, 99940, 99990, 
    100010, 100030, 100060, 100080, 100100, 100140, 100170, 100220, 100260, 
    100280, 100310, 100310, 100340, 100340, 100340, 100310, 100370, 100380, 
    100420, 100420, 100400, 100340, 100400, 100390, 100400, 100360, 100360, 
    100400, 100410, 100430, 100510, 100660, 100730, 100770, 100780, 100840, 
    100940, 101040, 101090, 101160, 101240, 101290, 101290, 101330, 101360, 
    101440, 101510, 101520, 101480, 101500, 101560, 101560, 101590, 101600, 
    101670, 101620, 101600, 101670, 101640, 101610, 101590, 101540, 101460, 
    101320, 101150, 100920, 100790, 100770, 100590, 100470, 100390, 100290, 
    100230, 100140, 100120, 100060, 100130, 100170, 100150, 100190, 100250, 
    100320, 100350, 100350, 100390, 100360, 100330, 100320, 100290, 100320, 
    100310, 100300, 100200, 100090, 100060, 100020, 99950, 99840, 99690, 
    99490, 99350, 99150, 98940, 98680, 98460, 98230, 98060, 98000, 97930, 
    97890, 97880, 97870, 97910, 97950, 98020, 98070, 98100, 98120, 98170, 
    98240, 98290, 98390, 98420, 98480, 98530, 98610, 98660, 98690, 98700, 
    98760, 98800, 98860, 98890, 98910, 98880, 98860, 98960, 98930, 98890, 
    98870, 98860, 98840, 98940, 99020, 99040, 99090, 99130, 99150, 99230, 
    99360, 99500, 99600, 99620, 99840, 99900, 100030, 100100, 100110, 100190, 
    100360, 100490, 100560, 100630, 100590, 100650, 100680, 100740, 100760, 
    100820, 100840, 100800, 100840, 100880, 100860, 100890, 100860, 100840, 
    100840, 100880, 100890, 100900, 100870, 100870, 100870, 100880, 100890, 
    100880, 100890, 100930, 100920, 100900, 100920, 100960, 100930, 100920, 
    100940, 100930, 100950, 100920, 100950, 100960, 100940, 100940, 100950, 
    100920, 100900, 100890, 100880, 100860, 100860, 100840, 100830, 100810, 
    100740, 100730, 100730, 100710, 100700, 100680, 100630, 100610, 100600, 
    100600, 100590, 100580, 100570, 100530, 100510, 100490, 100450, 100420, 
    100390, 100370, 100340, 100340, 100340, 100340, 100330, 100320, 100300, 
    100310, 100330, 100320, 100320, 100350, 100380, 100390, 100390, 100360, 
    100350, 100310, 100300, 100280, 100300, 100280, 100280, 100320, 100320, 
    100350, 100370, 100390, 100400, 100410, 100410, 100430, 100460, 100500, 
    100540, 100540, 100550, 100570, 100660, 100620, 100640, 100700, 100720, 
    100720, 100720, 100750, 100780, 100790, 100820, 100840, 100860, 100910, 
    100920, 100910, 100890, 100970, 100940, 100990, 101010, 101010, 101030, 
    101040, 101080, 101080, 101110, 101120, 101130, 101120, 101120, 101100, 
    101130, 101200, 101190, 101210, 101200, 101230, 101260, 101220, 101210, 
    101200, 101230, 101200, 101200, 101210, 101220, 101210, 101200, 101160, 
    101130, 101090, 101070, 100970, 100850, 100660, 100610, 100560, 100470, 
    100500, 100470, 100500, 100530, 100560, 100570, 100610, 100620, 100600, 
    100610, 100610, 100600, 100590, 100590, 100610, 100610, 100610, 100590, 
    100560, 100480, 100460, 100430, 100410, 100410, 100320, 100320, 100300, 
    100270, 100280, 100240, 100220, 100180, 100120, 100080, 100040, 100020, 
    100070, 100160, 100170, 100210, 100250, 100310, 100350, 100410, 100490, 
    100540, 100610, 100670, 100720, 100780, 100840, 100890, 100920, 100970, 
    101000, 101040, 101040, 101090, 101150, 101170, 101170, 101180, 101200, 
    101230, 101230, 101260, 101260, 101270, 101280, 101310, 101330, 101370, 
    101420, 101400, 101420, 101410, 101470, 101490, 101480, 101500, 101510, 
    101530, 101530, 101540, 101550, 101550, 101540, 101550, 101580, 101590, 
    101570, 101570, 101570, 101550, 101550, 101550, 101570, 101560, 101550, 
    101510, 101510, 101490, 101440, 101430, 101430, 101400, 101380, 101370, 
    101380, 101370, 101360, 101340, 101290, 101280, 101240, 101220, 101200, 
    101180, 101160, 101170, 101140, 101130, 101160, 101130, 101100, 101090, 
    101060, 101030, 101040, 101020, 100980, 100940, 100900, 100910, 100880, 
    100860, 100840, 100820, 100820, 100760, 100740, 100710, 100690, 100700, 
    100680, 100650, 100570, 100490, 100420, 100430, 100430, 100510, 100490, 
    100540, 100590, 100610, 100640, 100660, 100730, 100690, 100680, 100610, 
    100530, 100460, 100310, 100180, 100070, 99960, 99820, 99710, 99560, 
    99360, 99240, 99080, 98920, 98800, 98710, 98650, 98610, 98490, 98430, 
    98390, 98340, 98300, 98320, 98380, 98390, 98440, 98500, 98630, 98740, 
    98820, 98940, 99050, 99130, 99210, 99250, 99330, 99350, 99350, 99370, 
    99410, 99450, 99490, 99490, 99540, 99580, 99600, 99600, 99600, 99630, 
    99610, 99610, 99570, 99580, 99590, 99590, 99590, 99640, 99680, 99720, 
    99690, 99710, 99710, 99770, 99780, 99800, 99850, 99870, 99910, 99940, 
    99950, 99960, 99970, 99970, 99980, 100020, 100040, 100070, 100110, 
    100140, 100190, 100250, 100290, 100250, 100280, 100320, 100330, 100370, 
    100380, 100380, 100450, 100560, 100640, 100720, 100770, 100870, 100890, 
    100960, 101000, 101080, 101160, 101220, 101280, 101340, 101400, 101460, 
    101480, 101480, 101530, 101570, 101580, 101660, 101680, 101740, 101790, 
    101820, 101780, 101830, 101830, 101820, 101820, 101830, 101880, 101920, 
    101950, 101990, 102020, 102030, 102000, 101970, 101970, 101900, 101880, 
    101830, 101760, 101750, 101730, 101760, 101750, 101820, 101880, 101950, 
    102000, 102020, 102050, 102060, 102090, 102110, 102150, 102190, 102230, 
    102280, 102320, 102360, 102360, 102370, 102390, 102420, 102390, 102350, 
    102330, 102310, 102310, 102330, 102310, 102280, 102190, 102120, 102040, 
    101980, 101900, 101840, 101750, 101670, 101560, 101520, 101580, 101510, 
    101470, 101430, 101400, 101360, 101360, 101310, 101230, 101070, 100960, 
    100950, 100930, 100900, 100980, 101100, 101300, 101470, 101550, 101640, 
    101720, 101780, 101870, 101910, 101940, 101960, 101950, 101930, 101960, 
    101970, 102000, 102050, 102100, 102090, 102090, 102100, 102090, 102090, 
    102090, 102090, 102100, 102090, 102060, 102070, 102080, 102070, 102090, 
    102120, 102140, 102150, 102160, 102160, 102160, 102150, 102160, 102160, 
    102160, 102160, 102180, 102180, 102210, 102200, 102220, 102200, 102230, 
    102250, 102250, 102270, 102270, 102280, 102280, 102280, 102280, 102300, 
    102270, 102290, 102270, 102270, 102250, 102250, 102220, 102200, 102180, 
    102170, 102140, 102100, 102050, 102020, 101960, 101920, 101920, 101890, 
    101840, 101800, 101760, 101740, 101700, 101640, 101600, 101610, 101590, 
    101570, 101540, 101480, 101470, 101470, 101460, 101440, 101410, 101380, 
    101350, 101320, 101350, 101310, 101280, 101270, 101230, 101250, 101240, 
    101220, 101230, 101190, 101180, 101170, 101140, 101130, 101130, 101120, 
    101130, 101120, 101140, 101090, 101090, 101010, 100940, 100950, 100960, 
    100850, 100830, 100780, 100730, 100690, 100650, 100620, 100570, 100550, 
    100490, 100450, 100480, 100500, 100510, 100520, 100460, 100500, 100540, 
    100620, 100650, 100720, 100760, 100790, 100810, 100790, 100810, 100840, 
    100840, 100850, 100860, 100880, 100910, 100940, 100940, 100960, 101050, 
    101110, 101090, 101110, 101130, 101110, 101110, 101110, 101120, 101110, 
    101080, 101050, 101040, 101020, 100990, 100960, 100920, 100940, 100970, 
    101000, 100980, 101020, 101060, 101080, 101120, 101150, 101170, 101180, 
    101190, 101210, 101230, 101280, 101320, 101350, 101380, 101420, 101410, 
    101440, 101460, 101490, 101490, 101520, 101600, 101630, 101650, 101690, 
    101720, 101720, 101750, 101790, 101790, 101790, 101800, 101830, 101850, 
    101900, 101910, 101920, 101930, 101940, 101950, 101960, 101970, 101970, 
    101960, 101970, 101990, 102040, 102050, 102060, 102070, 102090, 102070, 
    102090, 102100, 102080, 102080, 102090, 102100, 102140, 102120, 102170, 
    102130, 102120, 102180, 102180, 102180, 102180, 102180, 102230, 102270, 
    102310, 102340, 102360, 102400, 102430, 102440, 102480, 102490, 102510, 
    102560, 102600, 102630, 102670, 102710, 102740, 102740, 102760, 102800, 
    102820, 102810, 102810, 102830, 102860, 102890, 102900, 102890, 102880, 
    102860, 102850, 102830, 102790, 102750, 102730, 102680, 102640, 102610, 
    102590, 102560, 102500, 102470, 102390, 102330, 102290, 102210, 102140, 
    102110, 102080, 102070, 102030, 101990, 101940, 101890, 101800, 101720, 
    101690, 101660, 101620, 101580, 101570, 101540, 101540, 101560, 101530, 
    101530, 101540, 101540, 101530, 101530, 101550, 101540, 101540, 101550, 
    101580, 101570, 101570, 101590, 101520, 101540, 101540, 101510, 101470, 
    101440, 101410, 101400, 101320, 101290, 101220, 101170, 101130, 101050, 
    100980, 100880, 100790, 100650, 100530, 100490, 100410, 100340, 100210, 
    100100, 100040, 99920, 99790, 99660, 99570, 99500, 99520, 99460, 99300, 
    99110, 98960, 98770, 98420, 98180, 97930, 97480, 97260, 97130, 97120, 
    97140, 97200, 97250, 97300, 97410, 97520, 97560, 97710, 97850, 98010, 
    98160, 98340, 98530, 98640, 98810, 98940, 99050, 99200, 99310, 99410, 
    99520, 99650, 99850, 100000, 100220, 100370, 100540, 100690, 100750, 
    100840, 100870, 100910, 100960, 100960, 100880, 100790, 100810, 100840, 
    100940, 101020, 101030, 101010, 101010, 101020, 100980, 100930, 100880, 
    100710, 100510, 100330, 100170, 100050, 99720, 99500, 99400, 99250, 
    99120, 98990, 98880, 98820, 98810, 98800, 98780, 98750, 98720, 98740, 
    98740, 98700, 98720, 98700, 98690, 98690, 98710, 98730, 98780, 98820, 
    98830, 98860, 98910, 98930, 98940, 98940, 99000, 99070, 99090, 99140, 
    99210, 99260, 99300, 99370, 99430, 99500, 99550, 99580, 99620, 99660, 
    99720, 99770, 99800, 99840, 99830, 99880, 99910, 99930, 99940, 100000, 
    100060, 100080, 100140, 100200, 100230, 100250, 100230, 100250, 100220, 
    100230, 100230, 100180, 100190, 100180, 100220, 100200, 100140, 100070, 
    100020, 99940, 99860, 99760, 99650, 99550, 99470, 99400, 99300, 99230, 
    99090, 99030, 98900, 98920, 99060, 99220, 99340, 99480, 99520, 99620, 
    99690, 99750, 99770, 99820, 99840, 99860, 99870, 99880, 99910, 99970, 
    100040, 100120, 100190, 100280, 100350, 100450, 100520, 100580, 100620, 
    100680, 100730, 100750, 100790, 100830, 100860, 100930, 100970, 101010, 
    101010, 101030, 101060, 101080, 101110, 101130, 101160, 101180, 101230, 
    101270, 101280, 101300, 101320, 101330, 101360, 101370, 101390, 101370, 
    101380, 101390, 101420, 101440, 101430, 101430, 101400, 101400, 101370, 
    101380, 101390, 101400, 101410, 101430, 101450, 101480, 101490, 101510, 
    101520, 101530, 101550, 101550, 101560, 101560, 101580, 101610, 101630, 
    101660, 101680, 101680, 101690, 101680, 101690, 101690, 101690, 101700, 
    101710, 101700, 101690, 101690, 101700, 101710, 101710, 101700, 101700, 
    101700, 101670, 101700, 101720, 101720, 101740, 101780, 101810, 101840, 
    101850, 101870, 101900, 101900, 101940, 101970, 101970, 102000, 102040, 
    102080, 102100, 102110, 102130, 102160, 102160, 102170, 102170, 102160, 
    102170, 102180, 102210, 102240, 102240, 102260, 102270, 102280, 102300, 
    102320, 102310, 102340, 102360, 102390, 102450, 102520, 102550, 102560, 
    102590, 102650, 102740, 102790, 102840, 102840, 102870, 102900, 102960, 
    103000, 103040, 103100, 103120, 103140, 103180, 103230, 103270, 103270, 
    103290, 103300, 103330, 103360, 103380, 103390, 103390, 103400, 103410, 
    103400, 103390, 103340, 103320, 103310, 103300, 103320, 103320, 103310, 
    103320, 103300, 103310, 103310, 103290, 103260, 103250, 103230, 103220, 
    103220, 103220, 103200, 103170, 103160, 103140, 103120, 103110, 103100, 
    103100, 103080, 103080, 103110, 103140, 103150, 103160, 103150, 103160, 
    103170, 103160, 103130, 103160, 103170, 103180, 103180, 103210, 103210, 
    103220, 103240, 103280, 103310, 103290, 103280, 103290, 103360, 103420, 
    103470, 103510, 103540, 103580, 103590, 103590, 103610, 103630, 103640, 
    103640, 103650, 103630, 103620, 103680, 103680, 103630, 103620, 103610, 
    103610, 103610, 103580, 103560, 103530, 103530, 103550, 103580, 103570, 
    103560, 103580, 103610, 103600, 103630, 103640, 103600, 103580, 103610, 
    103640, 103670, 103700, 103700, 103790, 103760, 103780, 103790, 103790, 
    103790, 103820, 103840, 103870, 103920, 103960, 103980, 104020, 104050, 
    104060, 104070, 104120, 104130, 104160, 104180, 104200, 104230, 104250, 
    104250, 104250, 104250, 104280, 104260, 104230, 104190, 104190, 104160, 
    104150, 104160, 104140, 104090, 104060, 104040, 104030, 104030, 103990, 
    103930, 103880, 103890, 103890, 103880, 103910, 103860, 103840, 103850, 
    103890, 103870, 103920, 103980, 103990, 104030, 104090, 104140, 104230, 
    104290, 104360, 104390, 104420, 104440, 104460, 104470, 104470, 104470, 
    104450, 104420, 104420, 104380, 104340, 104310, 104280, 104240, 104210, 
    104180, 104120, 104110, 104060, 104060, 104020, 103970, 103860, 103820, 
    103850, 103810, 103790, 103680, 103720, 103660, 103600, 103520, 103530, 
    103470, 103440, 103390, 103360, 103280, 103270, 103240, 103230, 103270, 
    103270, 103290, 103310, 103270, 103180, 103080, 103140, 103020, 102950, 
    102790, 102700, 102550, 102430, 102300, 102220, 102170, 102080, 102030, 
    101920, 101830, 101760, 101680, 101640, 101600, 101570, 101570, 101490, 
    101400, 101380, 101310, 101300, 101300, 101310, 101290, 101290, 101350, 
    101360, 101400, 101460, 101490, 101540, 101590, 101650, 101710, 101710, 
    101740, 101770, 101830, 101920, 102050, 102110, 102200, 102270, 102370, 
    102440, 102540, 102610, 102660, 102680, 102710, 102760, 102790, 102800, 
    102830, 102840, 102850, 102870, 102890, 102850, 102810, 102780, 102770, 
    102730, 102710, 102720, 102690, 102660, 102580, 102490, 102460, 102430, 
    102410, 102430, 102350, 102300, 102240, 102240, 102220, 102180, 102200, 
    102200, 102170, 102110, 102120, 102110, 102010, 102080, 102060, 102110, 
    102130, 102190, 102200, 102250, 102220, 102240, 102270, 102280, 102330, 
    102370, 102420, 102460, 102510, 102550, 102580, 102620, 102620, 102640, 
    102660, 102690, 102750, 102810, 102830, 102880, 102910, 102900, 102940, 
    102980, 103040, 103070, 103100, 103140, 103180, 103190, 103210, 103240, 
    103220, 103240, 103250, 103260, 103270, 103280, 103280, 103310, 103310, 
    103310, 103390, 103320, 103320, 103240, 103220, 103210, 103290, 103450, 
    103390, 103330, 103310, 103380, 103410, 103420, 103360, 103340, 103310, 
    103280, 103280, 103260, 103240, 103240, 103220, 103220, 103210, 103210, 
    103160, 103160, 103150, 103140, 103130, 103130, 103150, 103150, 103130, 
    103150, 103160, 103200, 103190, 103190, 103180, 103180, 103170, 103170, 
    103170, 103150, 103160, 103180, 103200, 103210, 103210, 103180, 103180, 
    103180, 103180, 103180, 103170, 103170, 103180, 103190, 103190, 103170, 
    103150, 103160, 103140, 103140, 103130, 103140, 103120, 103110, 103110, 
    103120, 103130, 103150, 103130, 103140, 103150, 103160, 103150, 103160, 
    103140, 103140, 103140, 103180, 103180, 103180, 103180, 103180, 103160, 
    103170, 103170, 103170, 103170, 103170, 103180, 103210, 103230, 103220, 
    103230, 103230, 103240, 103260, 103260, 103240, 103250, 103250, 103280, 
    103290, 103300, 103300, 103310, 103310, 103310, 103310, 103320, 103320, 
    103320, 103360, 103360, 103410, 103410, 103410, 103400, 103420, 103440, 
    103440, 103450, 103430, 103430, 103430, 103430, 103420, 103410, 103380, 
    103380, 103340, 103330, 103310, 103310, 103290, 103290, 103280, 103270, 
    103250, 103240, 103210, 103220, 103200, 103200, 103160, 103170, 103170, 
    103180, 103150, 103160, 103170, 103170, 103150, 103100, 103060, 103030, 
    103010, 102960, 102920, 102870, 102860, 102820, 102780, 102750, 102700, 
    102660, 102620, 102580, 102600, 102590, 102590, 102590, 102620, 102630, 
    102630, 102610, 102550, 102540, 102520, 102490, 102450, 102440, 102420, 
    102400, 102380, 102370, 102360, 102330, 102350, 102380, 102380, 102370, 
    102340, 102350, 102370, 102360, 102380, 102380, 102400, 102430, 102430, 
    102420, 102440, 102440, 102420, 102400, 102420, 102400, 102420, 102440, 
    102450, 102460, 102460, 102470, 102480, 102430, 102470, 102470, 102480, 
    102470, 102470, 102470, 102500, 102500, 102510, 102520, 102550, 102550, 
    102520, 102560, 102570, 102540, 102570, 102610, 102640, 102650, 102630, 
    102630, 102650, 102670, 102690, 102720, 102720, 102720, 102720, 102710, 
    102710, 102700, 102670, 102650, 102620, 102640, 102630, 102630, 102650, 
    102650, 102660, 102670, 102670, 102720, 102690, 102700, 102710, 102720, 
    102720, 102720, 102650, 102640, 102650, 102570, 102640, 102640, 102550, 
    102520, 102520, 102450, 102400, 102410, 102380, 102350, 102280, 102260, 
    102230, 102200, 102150, 102090, 102010, 102000, 101920, 101870, 101810, 
    101750, 101680, 101620, 101530, 101400, 101310, 101180, 101070, 101000, 
    100940, 100850, 100760, 100670, 100570, 100510, 100460, 100360, 100310, 
    100270, 100220, 100240, 100250, 100300, 100340, 100240, 100300, 100370, 
    100370, 100530, 100680, 100730, 100780, 100690, 100810, 100930, 101190, 
    101320, 101350, 101390, 101410, 101400, 101480, 101480, 101630, 101680, 
    101740, 101800, 101840, 101940, 102090, 102130, 102180, 102190, 102260, 
    102230, 102140, 102130, 102150, 102210, 102260, 102310, 102310, 102300, 
    102290, 102280, 102280, 102250, 102250, 102260, 102230, 102240, 102210, 
    102190, 102150, 102130, 102100, 102090, 102060, 102010, 101970, 101970, 
    101940, 101920, 101910, 101890, 101850, 101830, 101820, 101810, 101770, 
    101750, 101730, 101680, 101650, 101620, 101580, 101550, 101500, 101440, 
    101400, 101370, 101320, 101310, 101230, 101180, 101140, 101070, 101050, 
    101000, 100940, 100870, 100820, 100790, 100730, 100680, 100640, 100560, 
    100490, 100450, 100380, 100320, 100260, 100230, 100210, 100180, 100110, 
    100070, 99990, 99950, 99920, 99890, 99910, 100000, 100030, 99990, 99940, 
    99940, 99880, 99800, 99800, 99830, 99890, 99950, 99990, 100020, 100080, 
    100150, 100240, 100310, 100330, 100320, 100280, 100220, 100260, 100300, 
    100370, 100430, 100490, 100520, 100590, 100630, 100630, 100650, 100700, 
    100670, 100640, 100770, 100830, 100810, 100880, 100870, 100890, 100970, 
    100990, 101050, 101140, 101170, 101190, 101230, 101230, 101210, 101220, 
    101280, 101300, 101330, 101360, 101410, 101460, 101490, 101530, 101610, 
    101590, 101700, 101710, 101680, 101700, 101680, 101650, 101680, 101690, 
    101740, 101790, 101780, 101790, 101770, 101760, 101750, 101760, 101750, 
    101720, 101690, 101590, 101490, 101460, 101300, 101110, 100930, 100820, 
    100760, 100730, 100740, 100760, 100750, 100800, 100810, 100850, 100880, 
    _, 100860, 100840, 100830, 100830, 100800, 100750, 100720, 100660, 
    100640, 100670, 100720, 100740, 100740, 100760, 100780, 100840, 100850, 
    100870, 100890, 100880, 100880, 100880, 100880, 100860, 100860, 100820, 
    100810, 100810, 100800, 100780, 100760, 100760, 100730, 100720, 100710, 
    100690, 100640, 100610, 100590, 100570, 100550, 100530, 100510, 100510, 
    100480, 100460, 100490, 100490, 100490, 100490, 100510, 100550, 100580, 
    100620, 100610, 100640, 100660, 100680, 100690, 100700, 100710, 100720, 
    _, 100790, 100830, 100860, _, 100890, 100890, 100880, 100920, _, 100950, 
    100960, 100990, 101040, 101070, 101100, 101120, 101120, 101120, 101110, 
    101120, 101110, 101120, 101120, 101110, 101140, 101140, 101140, 101130, 
    101100, 101110, 101100, 101090, 101090, 101070, 101060, 101080, _, 
    101110, _, 101120, 101100, 101100, 101070, 101080, 101080, _, 101110, 
    101140, 101150, 101160, 101180, 101200, 101220, 101210, 101240, 101250, 
    101250, 101230, 101270, 101310, 101360, _, 101400, 101420, 101460, 
    101490, 101540, 101560, 101590, 101630, 101650, 101680, 101730, 101750, 
    101780, 101880, 101930, 101970, 102010, 102030, _, 102090, 102140, 
    102180, 102220, 102280, 102310, 102330, 102340, 102350, 102350, 102360, 
    _, 102410, 102430, 102460, 102510, 102540, 102590, 102610, 102660, 
    102690, 102720, 102730, 102780, 102820, _, _, 102930, 102950, _, 103040, 
    103060, 103070, 103070, 103100, 103120, 103140, 103150, 103150, 103190, 
    103200, 103190, 103190, 103200, 103190, 103190, 103190, 103170, 103170, 
    103150, 103160, 103150, 103150, 103160, 103160, 103130, 103110, _, 
    103100, 103090, 103100, 103070, 103080, 103060, 103080, 103070, 103030, 
    _, 102950, 102940, 102950, _, 102920, 102910, 102890, 102850, 102850, 
    102830, 102800, 102780, 102720, 102710, 102700, _, 102630, 102600, 
    102570, 102550, 102520, 102500, 102480, 102450, 102420, 102380, 102350, 
    102310, 102300, 102270, 102260, 102230, 102210, _, 102180, 102140, 
    102110, 102080, 102050, 102030, 102030, 102030, 102020, 102000, 101980, 
    101960, 101960, 101950, 101940, 101940, 101920, 101930, 101950, 101970, 
    101990, 101960, 101990, 102010, 102000, 102000, 101990, 101970, 101950, 
    101960, 101990, 101980, 102010, 101990, 102000, 101960, 101940, 101990, 
    101930, 101930, 101930, 101910, 101890, 101860, 101840, 101820, 101780, 
    101740, 101700, 101740, 101660, 101610, _, 101580, 101570, 101560, 
    101550, 101520, 101500, 101480, 101460, 101450, 101400, 101370, 101320, 
    101250, 101210, 101100, 101040, 100930, 100870, _, 100940, 100940, 
    100950, 100960, 100950, 100960, _, 100960, 100940, 100920, 100930, 
    100930, 100930, 100920, 100900, 100880, 100840, 100790, 100750, 100740, 
    100700, 100680, 100650, 100640, 100630, 100620, 100590, 100570, 100520, 
    100460, 100380, 100290, 100230, 100160, 100080, 100030, 99960, 99900, 
    99810, 99730, 99680, _, 99630, 99650, 99670, 99750, 99880, 99960, 100150, 
    100290, 100360, 100430, _, 100550, 100630, 100640, 100740, 100820, 
    100850, 100850, 100860, 100850, 100840, 100810, 100790, 100740, 100720, 
    100760, 100790, 100810, 100820, _, 100800, 100820, 100810, 100810, 
    100800, 100760, 100780, 100800, 100810, 100880, 100890, 100950, 100950, 
    101000, 101040, 101090, 101110, 101110, 101110, 101090, 101090, 101090, 
    101060, 101040, 100990, 100930, 100840, 100740, 100620, 100470, 100390, 
    100230, 100130, 100020, 99980, 99970, 99970, 99990, 100030, 100080, 
    100120, 100130, 100120, 100140, 100160, 100190, 100210, 100220, 100210, 
    100260, 100270, 100370, 100520, 100630, 100740, 100840, 100950, 100990, 
    101030, 101110, 101080, 101100, 101180, 101210, 101250, 101200, 101280, 
    101340, _, 101400, 101390, 101420, 101430, 101430, 101450, _, 101480, 
    101490, 101460, 101460, 101460, 101470, 101470, 101490, 101520, 101570, 
    101620, 101680, 101730, 101760, 101850, 101890, 101930, 101990, 102030, 
    102050, 102030, 102050, 102070, 102050, 102010, _, 101900, 101860, 
    101830, 101800, 101760, 101690, 101650, 101590, 101560, _, 101500, 
    101450, 101410, 101400, 101400, 101410, 101420, 101390, 101350, 101320, 
    101290, 101250, 101230, 101170, 101080, 101010, _, 100870, 100840, 
    100760, 100730, 100720, 100690, 100660, 100620, 100590, 100580, 100600, 
    100610, 100650, 100680, 100660, 100570, 100460, 100370, _, 100550, 
    100810, 100940, 101000, 101160, 101240, 101360, 101390, 101300, 101430, 
    101430, 101540, 101500, 101570, 101590, 101590, 101660, 101660, 101730, 
    101780, 101870, 101820, 101870, 101960, 102030, 102100, 102150, 102190, 
    102240, 102280, 102310, 102360, 102390, 102400, 102410, 102420, 102420, 
    102400, 102400, 102420, 102430, 102440, 102460, 102480, 102480, _, 
    102470, 102460, 102440, 102400, 102370, 102360, 102350, 102300, 102280, 
    102280, 102240, 102230, 102200, 102160, 102130, 102080, 102020, 101970, 
    101900, 101850, 101810, 101820, 101780, 101710, 101730, 101680, 101630, 
    101580, 101540, 101500, 101450, 101400, 101360, 101320, 101260, 101190, 
    101170, _, 101040, 101000, 100960, 100910, 100880, 100850, 100800, 
    100780, 100700, 100640, 100530, 100520, 100470, 100430, 100370, 100320, 
    100310, 100250, 100270, 100250, 100280, 100300, 100310, 100380, 100460, 
    100520, 100580, 100670, 100720, 100760, 100820, 100840, _, 100890, 
    100880, 100880, 100890, _, 100840, 100820, 100820, 100820, 100810, _, 
    100890, 100900, 100930, 100930, 100930, 100950, 100960, _, 100990, 
    101000, 101030, 101050, 101050, _, 101040, 101020, 101010, 101000, 
    100990, 100980, 101000, 101000, 100990, 100980, 100960, 100950, 100940, 
    _, 100910, 100900, 100900, 100900, 100890, 100890, 100880, 100870, 
    100870, 100860, 100850, 100830, 100810, 100810, 100810, 100810, 100800, 
    100800, 100780, 100770, 100770, 100770, _, 100750, 100750, 100750, 
    100750, 100790, 100780, 100780, 100810, 100820, _, 100840, 100850, 
    100870, 100870, 100880, 100900, 100920, 100940, 100960, 100980, 100980, 
    100990, 101030, 101040, 101030, 101040, 101050, 101070, 101100, 101140, 
    101160, 101180, 101210, 101240, _, 101280, 101260, 101300, 101340, 
    101360, 101390, 101410, 101410, 101410, 101420, 101440, 101450, 101450, 
    101460, 101460, 101470, 101500, 101510, 101530, 101550, 101560, 101570, 
    101590, 101590, 101580, 101580, 101590, 101590, 101580, 101600, 101600, 
    101590, 101580, 101570, 101560, 101550, 101520, 101510, _, 101480, 
    101460, 101450, 101440, 101420, 101400, 101350, 101330, 101290, 101270, 
    101230, 101190, 101140, 101100, 101070, 101030, 101010, 100970, 100940, 
    100910, 100900, 100900, 100890, 100880, 100870, 100880, 100890, 100920, 
    100930, 100940, 100960, 100970, _, 101000, 101020, 101020, 101040, 
    101030, 101030, 101050, 101070, 101080, 101070, 101090, 101120, 101130, 
    101150, 101150, 101170, 101180, 101200, 101230, 101260, 101290, 101330, 
    101340, 101370, 101380, 101420, 101430, 101420, 101440, 101450, 101480, 
    101470, 101480, 101510, 101510, 101560, 101610, 101640, 101640, 101620, 
    101670, 101720, _, 101790, 101830, 101880, 101930, 101950, 101980, 
    102020, 102040, 102080, 102070, 102090, 102140, 102170, 102190, 102190, 
    102210, 102180, 102200, 102210, 102180, 102180, 102180, 102190, 102170, 
    102160, 102200, 102200, 102190, _, 102230, 102200, 102190, 102180, 
    102180, 102180, 102220, 102210, 102230, 102220, 102190, 102200, 102180, 
    _, 102180, 102160, 102170, 102150, 102140, 102120, 102150, 102140, 
    102100, 102090, 102080, 102080, 102090, 102080, 102060, 102070, 102070, 
    102060, 102090, 102120, 102100, 102090, 102050, 102000, 101950, 101890, 
    101790, 101770, 101740, 101690, 101690, 101620, 101620, 101600, 101600, 
    101530, 101450, 101400, 101410, 101370, 101340, 101370, 101360, 101360, 
    101370, 101300, 101300, 101280, 101250, 101220, 101160, 101110, 101070, 
    101080, 101030, 100990, 100990, _, 100880, 100830, 100780, 100730, 
    100680, 100590, 100530, 100480, 100420, 100370, 100340, 100310, 100260, 
    100260, 100220, 100250, 100280, 100270, 100290, 100270, 100250, 100220, 
    100180, 100110, 100050, 99980, 99910, 99870, 99800, 99750, 99700, 99670, 
    99640, 99590, 99560, 99540, 99540, 99520, 99510, 99520, 99570, 99600, 
    99640, 99710, 99780, 99880, 99970, _, 100190, 100290, 100370, 100490, 
    100570, 100630, 100700, 100760, 100790, 100810, 100820, 100840, 100840, 
    100850, 100830, 100850, 100830, 100840, 100840, 100810, 100790, 100770, 
    100740, _, 100640, 100530, 100460, 100370, 100340, 100370, 100350, 
    100400, 100400, 100400, 100430, 100520, 100570, 100650, 100700, 100760, 
    100780, 100880, 100910, 100950, 100990, 100990, 100990, 100960, 100920, 
    100790, 100750, 100700, 100550, 100490, 100360, 100240, 100150, 100050, 
    99920, 99820, 99770, 99710, 99610, 99600, 99670, 99780, 99800, 99950, 
    100070, 100170, 100280, 100400, 100570, 100650, 100730, 100810, 100900, 
    100990, 101050, 101120, 101180, 101220, 101290, 101390, 101450, 101480, 
    101520, 101550, 101620, 101670, 101710, 101720, 101740, 101750, 101750, 
    101760, 101730, 101660, 101580, 101510, 101420, 101270, 101070, 100910, 
    100770, 100510, 100360, 100140, 99970, 99920, 99860, 99860, 99880, 99950, 
    100060, 100170, 100300, 100450, 100580, 100670, _, 100840, 100930, 
    101000, 101080, 101200, 101290, 101390, 101460, 101560, 101640, 101710, 
    101750, 101860, 101880, 101900, 101890, 101910, 101900, 101870, 101850, 
    101770, 101700, 101640, 101550, 101420, 101340, 101230, 101200, 101170, 
    101250, 101360, 101420, 101560, 101670, 101860, 102170, 102270, 102380, 
    102510, 102560, 102640, 102720, 102800, 102800, 102820, 102860, 102890, 
    102900, 102880, 102820, 102790, 102770, 102730, 102720, 102670, 102640, 
    102610, 102520, 102490, 102450, 102370, 102270, 102220, 102130, 102100, 
    102080, 102060, 102020, 101990, 101950, 101940, 101910, 101870, 101820, 
    101770, 101750, 101730, 101740, 101720, 101710, 101690, 101730, 101670, 
    101670, 101660, 101620, 101600, 101580, 101600, 101600, 101590, 101610, 
    101650, 101660, 101630, 101650, 101690, 101700, 101710, 101740, 101720, 
    101740, 101770, 101770, 101730, 101710, 101710, 101700, 101640, 101570, 
    101590, 101550, 101530, 101430, 101410, 101470, 101470, 101430, 101370, 
    101300, 101230, 101180, 101090, 101010, 101050, 101080, 101090, 101060, 
    101060, 101060, 101060, 101000, 101000, 100980, 100980, 100950, 100980, 
    100980, 100970, 100950, 100930, 100870, 100830, 100800, 100810, 100740, 
    100640, 100620, 100610, 100640, 100660, 100650, 100620, 100580, 100560, 
    100530, 100490, 100450, _, 100300, 100320, 100340, 100320, 100300, 
    100300, 100300, 100280, 100260, 100200, 100220, 100180, 100110, 100140, 
    100190, 100240, 100160, 100100, 100140, 100170, 100160, _, 100070, 
    100160, 100140, 100190, 100270, 100330, 100370, 100420, 100450, 100450, 
    100430, 100430, 100430, 100390, 100330, 100230, 100200, 100190, 100130, 
    100120, 100140, 100080, 100070, 100040, 100050, 100030, 100020, 100030, 
    100070, 100140, 100180, _, 100270, 100320, 100370, 100430, 100480, 
    100520, 100560, _, 100650, 100690, 100720, 100760, 100780, 100790, 
    100820, 100840, 100860, 100860, 100860, 100860, 100880, 100890, 100900, 
    100910, 100940, 100940, 100940, 100940, 100930, 100920, 100910, 100890, 
    100910, 100920, 100920, 100920, 100950, 100980, 101000, 101020, 101040, 
    101060, _, 101160, 101220, 101270, 101310, 101340, 101370, 101390, 
    101430, 101440, 101430, 101420, 101400, 101400, 101410, 101420, 101420, 
    101420, 101370, 101390, 101340, 101300, 101250, 101210, 101150, 101100, 
    101070, 101060, 101020, 100970, 100950, 100900, 100840, 100810, 100790, 
    100750, 100720, 100740, 100740, 100740, 100740, 100740, 100740, 100740, 
    100750, 100740, 100760, 100790, 100830, 100880, 100930, 100940, 100980, 
    101000, 101010, 101010, 100990, 100950, 100900, 100870, 100800, 100760, 
    100700, 100660, 100620, 100550, 100490, 100400, 100340, 100300, 100270, 
    100240, _, 100230, 100260, 100300, 100360, 100410, 100480, 100520, 
    100560, 100590, 100640, 100680, 100710, 100740, 100760, 100780, 100800, 
    100840, 100880, 100940, 101010, 101050, 101080, 101100, 101130, 101180, 
    101240, 101290, 101340, 101340, 101360, 101370, 101360, 101320, 101300, 
    101280, 101250, 101240, 101210, 101200, 101160, 101160, 101150, 101150, 
    101170, 101180, 101190, 101220, 101260, 101310, 101360, 101410, 101460, 
    101550, 101590, 101620, 101660, 101710, 101730, 101770, 101790, _, 
    101850, 101900, 101930, 101960, 101980, 101960, 101950, 101960, 101960, 
    101990, _, 102020, 102060, 102090, 102100, 102070, 102110, 102120, 
    102130, 102130, 102120, 102120, 102120, 102110, 102120, 102120, 102110, 
    102100, 102110, 102110, 102100, 102120, 102120, 102140, 102170, 102220, 
    102250, 102250, 102270, 102290, 102300, 102300, 102300, 102290, 102280, 
    102270, 102270, _, 102220, 102210, 102210, 102180, _, 102120, 102100, 
    102070, 102030, 102010, 101990, 101950, 101880, 101830, 101780, 101710, 
    101680, 101630, 101540, 101470, 101410, 101370, 101310, 101260, 101190, 
    101150, 101090, 101040, 101010, 100990, 100980, 100970, 100970, 100920, 
    _, 100940, 100940, 100940, 100950, 100950, 100920, 100910, 100860, 
    100830, 100800, 100810, 100810, 100810, 100810, 100770, 100740, 100710, 
    100670, 100650, 100630, 100580, 100550, 100520, 100510, 100490, 100480, 
    100460, 100470, 100460, 100470, 100460, 100450, 100450, 100400, 100370, 
    100330, 100270, 100260, 100230, 100220, 100200, _, 100180, 100170, 
    100150, 100120, 100130, 100150, 100190, 100210, 100240, 100230, _, 
    100230, 100200, 100220, 100150, 100210, 100290, 100350, 100420, _, 
    100510, 100570, 100650, 100640, 100750, 100850, 100920, 100970, 101080, 
    101130, 101180, 101210, 101290, 101330, 101390, 101430, 101480, 101510, 
    101500, 101520, 101530, 101550, 101550, 101560, 101550, 101530, 101510, 
    101490, 101480, 101470, 101460, 101380, 101370, 101330, 101340, 101350, 
    101330, 101260, 101280, 101210, 101240, 101260, 101120, 101180, 101140, 
    101040, 101070, 100950, 100900, 100910, 100790, 100700, 100690, 100620, 
    100600, 100600, 100570, 100520, 100590, 100570, 100540, 100520, _, _, 
    100480, 100470, 100430, 100390, 100380, 100360, 100320, 100240, 100150, 
    99980, 99900, 99850, 99810, 99690, 99580, 99550, 99330, 99220, 99120, 
    98930, 98770, _, 98540, 98370, 98260, 98130, 98070, 98050, 98060, 98110, 
    98110, 98080, 98170, 98290, 98380, 98450, 98500, 98570, 98630, 98670, 
    98570, 98740, 98870, 98940, 99010, 99100, 99240, 99420, 99420, 99600, 
    99700, 99830, 99950, 100090, 100200, 100330, 100400, 100500, 100600, 
    100700, 100780, 100810, 100900, 100960, 101020, 101060, 101120, 101180, 
    _, 101280, 101320, 101370, 101410, 101440, 101450, 101460, 101460, 
    101470, 101480, 101500, 101500, 101520, 101520, 101530, 101540, 101560, 
    101560, 101560, 101560, 101580, 101580, 101590, 101600, 101620, 101620, 
    101630, 101640, 101640, 101640, 101630, 101600, 101610, 101580, 101590, 
    101570, 101540, 101520, 101500, 101460, 101410, 101330, 101250, 101250, 
    101210, 101190, 101200, 101130, 101040, 100960, 100930, 100940, 100890, 
    100830, 100740, 100720, 100680, 100660, 100600, 100560, _, 100490, 
    100470, 100480, 100470, 100460, 100470, 100430, 100470, 100460, 100460, 
    _, 100400, 100360, 100330, _, 100230, 100170, 100090, 100000, 99950, 
    99910, 99850, 99830, 99760, 99760, 99720, 99700, 99610, 99600, 99660, 
    99660, 99650, 99650, 99630, 99620, 99610, 99610, 99580, 99600, 99580, 
    99590, 99620, _, 99640, 99670, 99710, 99760, 99800, 99850, 99920, 99940, 
    99990, 100050, 100120, 100170, 100210, 100270, 100330, 100360, 100420, 
    100490, 100540, 100610, 100670, 100710, 100750, 100780, 100790, 100820, 
    100820, 100840, 100880, 100950, 101000, 101030, 101070, 101130, 101180, 
    101200, 101250, 101330, 101350, _, 101440, 101430, 101450, 101480, 
    101460, 101440, 101440, 101420, _, 101340, 101330, 101340, 101340, 
    101340, 101290, 101270, 101250, 101190, 101100, 100980, 100910, 100790, 
    _, 100730, 100670, 100590, 100610, 100560, 100450, 100410, 100400, 
    100360, 100320, 100320, 100350, 100340, 100350, 100330, 100280, 100260, 
    100270, 100190, 100160, 100120, 100070, 100020, 100000, 99970, 99960, 
    99930, 99900, 99860, 99820, 99810, 99810, 99840, 99840, 99860, 99920, 
    99950, 100010, 100020, 100100, 100160, 100210, 100280, 100340, 100370, 
    100470, 100560, 100670, 100750, 100830, 100900, 101000, 101070, 101110, 
    101150, 101210, 101240, 101260, 101290, 101320, 101300, 101310, 101300, 
    101290, 101280, 101260, 101250, 101220, 101190, 101180, 101170, _, 
    101080, 101050, 101010, 100960, 100880, 100850, 100820, 100780, 100680, 
    100510, 100340, 100240, 100180, _, 99900, 99730, 99700, 99690, 99710, 
    99640, 99690, 99690, 99720, 99770, 99800, 99820, 99830, 99860, 99910, 
    99970, 100050, 100160, _, 100350, 100430, 100510, 100570, 100640, 100670, 
    100710, 100770, 100780, 100820, 100840, 100850, 100870, 100930, 100960, 
    100990, 101010, 101040, 101060, 101070, 101080, 101100, 101120, 101120, 
    101130, 101150, 101150, 101160, 101160, 101160, 101150, 101140, 101150, 
    101170, 101160, 101180, 101200, 101200, _, 101250, 101280, 101330, 
    101320, 101340, 101360, 101380, 101400, 101400, 101410, 101430, 101440, 
    101460, 101450, 101430, 101460, 101460, 101440, 101440, 101420, 101420, 
    101420, 101410, 101430, 101440, 101450, 101440, 101420, 101380, 101370, 
    101340, 101270, 101320, 101390, 101340, 101270, 101180, 101230, 101170, 
    100930, 101050, 101020, 100970, 100950, 100840, 100730, 100690, 100530, 
    _, 100460, 100320, 100280, 100170, 100110, 100030, 100030, 100010, 99950, 
    99940, 99890, 99880, 100050, 100020, 99990, 99940, 99950, 99880, 99890, 
    99840, 99830, 99820, _, 99780, 99760, 99730, 99730, 99720, 99680, 99640, 
    99610, 99580, 99540, 99560, 99520, 99490, _, 99450, 99420, 99400, 99390, 
    99370, 99380, 99350, 99330, 99350, 99340, 99350, 99320, 99340, 99320, 
    99290, 99280, 99250, 99210, 99170, 99140, 99130, 99120, 99100, 99070, 
    99050, 99030, 99000, 98980, 98960, 98950, 98970, 98990, 99010, 99040, 
    99110, 99160, 99200, 99240, 99260, 99300, 99330, 99340, 99380, 99410, 
    99460, 99490, 99530, 99540, 99590, 99610, 99620, 99660, 99670, 99670, 
    99690, 99670, 99700, _, 99740, _, 99790, 99810, 99800, 99790, 99810, 
    99820, 99830, 99820, 99810, 99840, 99830, 99830, _, 99810, 99810, 99770, 
    99750, 99750, 99790, 99820, 99860, 99880, 99910, 99930, 99950, 99980, 
    99980, 100000, 100020, 100030, 100030, 100060, 100060, 100100, 100110, 
    100150, 100190, 100090, 100060, 100100, 100180, 100260, 100300, 100300, 
    100380, 100400, 100420, 100500, 100550, 100520, 100560, 100590, 100610, 
    100620, 100610, 100590, 100570, 100530, 100480, 100460, 100460, 100420, 
    100400, 100350, 100310, 100300, 100290, 100320, 100310, 100280, 100280, 
    100280, 100250, 100260, 100270, 100240, 100260, 100270, 100260, 100250, 
    _, _, 100210, 100220, 100280, 100330, 100390, 100450, 100540, 100600, 
    100670, 100720, 100770, 100820, 100880, 100940, 100980, 101010, 101040, 
    101080, 101080, 101090, 101100, 101100, 101120, 101180, 101210, _, 
    101180, _, 101210, 101220, 101200, 101210, 101180, 101190, 101210, 
    101270, 101320, 101350, 101380, 101370, 101420, 101450, 101460, 101450, 
    101470, 101470, 101440, 101420, 101450, 101450, 101440, 101440, 101410, 
    101440, 101430, 101430, 101390, _, 101310, 101320, 101340, 101370, 
    101350, 101320, 101320, 101320, 101320, 101310, 101260, 101250, 101280, 
    101240, 101240, 101220, 101230, 101220, 101240, 101240, 101220, 101220, 
    101210, 101210, 101220, 101230, 101240, 101260, 101290, 101280, 101290, 
    101310, 101290, 101300, 101270, 101280, 101310, 101310, 101300, 101300, 
    101310, 101320, 101320, 101310, 101320, 101340, 101360, 101360, 101380, 
    101420, 101450, 101500, 101540, 101550, 101570, 101600, 101640, 101640, 
    101640, 101650, 101680, 101700, 101690, 101690, 101710, 101720, 101730, 
    101720, 101700, 101690, 101690, 101700, _, 101680, 101660, 101650, 
    101610, 101550, 101530, 101480, 101440, 101400, 101370, 101310, 101290, 
    101240, 101220, 101190, 101190, 101220, 101200, 101160, 101110, 101080, 
    101060, 101040, 101010, 100990, 100970, 100930, 100920, 100850, 100820, 
    100750, 100680, 100700, 100630, 100650, 100630, 100610, 100550, 100500, 
    100480, 100450, 100430, 100410, 100400, 100390, 100390, 100380, 100350, 
    100360, 100350, 100400, 100460, 100530, 100560, 100570, 100600, 100630, 
    100610, 100560, 100540, 100530, 100470, 100420, 100380, 100350, 100300, 
    100280, 100260, 100240, 100230, 100200, 100170, 100170, 100130, _, 
    100000, 100010, 99960, 99930, 99870, 99830, 99820, 99780, 99780, 99780, 
    99720, 99710, 99690, 99730, 99740, 99760, 99830, 99900, 99980, 100050, _, 
    100200, 100270, 100330, 100400, 100450, 100450, 100450, 100460, 100490, 
    100470, 100500, 100490, 100520, 100550, 100580, 100610, 100660, 100710, 
    100690, 100700, 100760, 100740, 100720, 100690, 100670, 100640, 100570, 
    100580, 100510, 100410, 100340, 100260, 100130, 100040, 99970, 99880, 
    99870, 99850, 99860, 99890, 99960, 100030, 100080, 100120, 100170, 
    100210, 100260, 100300, 100350, 100420, 100490, 100560, 100600, 100650, 
    100710, 100770, 100810, 100850, 100900, 100920, 100930, 100910, 100930, 
    100920, 100900, 100870, 100810, 100730, 100710, 100670, 100620, 100570, 
    100530, 100490, 100410, 100330, 100290, 100230, 100200, 100150, 100150, 
    100140, 100180, 100240, 100300, 100380, 100460, 100570, 100650, 100730, 
    100780, 100810, 100880, 100930, 100960, 101020, 101060, 101100, 101130, 
    101110, 101120, 101120, 101120, 101070, 101090, 101050, 101000, 100930, 
    100920, 100870, 100840, 100750, 100680, 100600, 100550, 100490, 100460, 
    100470, 100420, 100410, 100420, 100430, 100460, 100460, 100490, 100520, 
    100520, 100550, 100600, 100660, 100710, 100750, 100840, 100880, 100940, 
    101000, 101090, 101140, 101170, 101240, 101280, 101310, 101360, 101390, 
    101470, 101480, 101490, 101520, 101550, 101560, 101550, 101560, 101560, 
    101580, 101570, 101570, 101590, 101610, 101630, 101650, 101700, 101740, 
    101770, 101800, 101850, 101880, 101930, 101960, 101990, 102010, 102040, 
    102080, 102100, 102070, 102040, 102070, 102040, 102040, 101990, 101970, 
    101920, 101890, 101880, 101840, 101790, 101750, 101750, 101740, 101700, 
    101710, 101710, 101720, 101710, 101690, 101710, 101690, 101650, 101600, 
    101600, 101550, 101490, 101440, 101360, 101290, 101020, 101090, 100960, 
    100840, 100700, 100580, 100530, 100430, 100330, 100280, 100250, 100220, 
    100230, 100210, 100240, 100260, 100260, 100290, 100290, 100240, 100230, 
    _, 100200, 100220, 100250, 100260, 100280, 100300, 100320, 100310, 
    100330, 100350, 100410, 100370, 100420, 100470, 100510, 100560, 100580, 
    100600, 100640, 100680, 100690, 100720, 100780, 100810, _, 100900, 
    100970, 101010, 101050, 101120, 101160, 101180, 101210, 101220, 101200, 
    101230, 101240, 101220, 101190, 101160, 101130, 101130, 101100, 101050, 
    101010, 101010, 100980, 100910, 100870, 100810, 100780, 100790, 100760, 
    100760, 100750, 100720, 100710, 100660, 100600, 100610, 100580, 100590, 
    100580, 100550, 100530, 100550, 100520, 100510, _, 100540, 100560, 
    100520, 100520, 100510, 100510, 100510, 100460, 100450, 100410, 100400, 
    100370, 100350, 100340, 100320, 100300, 100290, 100280, 100270, 100260, 
    100270, 100260, 100250, 100240, 100240, 100230, 100230, _, 100270, 
    100280, 100310, 100340, 100380, 100410, 100470, 100500, 100520, 100590, 
    100690, 100740, 100800, 100910, 100980, 101010, 101050, 101090, 101130, 
    101140, 101110, 101100, 101070, 101040, 100990, 100940, 100930, 100910, 
    100860, 100800, 100770, 100700, 100640, 100630, 100590, 100580, 100620, 
    100590, 100550, 100590, 100630, 100660, 100690, 100710, 100710, 100750, 
    _, 100850, _, 100920, 100890, 100910, 100960, 100990, 100990, 100990, 
    101010, _, 101060, 101070, 101130, 101170, 101220, 101280, 101330, 
    101390, 101430, 101470, 101510, 101540, 101580, 101590, 101610, 101560, 
    101520, 101500, 101440, 101420, 101350, 101280, 101240, 101180, 101170, 
    101140, 101140, 101150, 101180, 101170, 101170, 101200, 101210, 101200, 
    101190, 101230, 101290, 101290, 101350, 101380, 101430, 101430, 101440, 
    101430, 101480, 101480, 101460, 101460, 101440, 101430, 101390, 101430, 
    101460, 101510, 101540, 101520, _, 101570, 101600, 101650, 101680, 
    101720, 101780, 101860, 101870, 101920, 101950, 101960, 101970, 102000, 
    102030, 102080, 102110, 102160, 102190, 102270, 102300, 102330, 102300, 
    102360, 102340, 102390, 102380, 102350, 102340, _, 102350, 102360, 
    102340, 102310, 102290, 102310, 102250, 102220, 102180, 102160, 102110, 
    102100, 102080, 102090, 102080, 102070, 102070, 102040, 102010, 102020, 
    102000, 101970, _, 101960, 101960, 101960, 101950, 101930, 101940, 
    101930, 101900, 101860, 101820, 101840, 101840, 101870, 101860, 101890, 
    101910, 101920, 101940, 101960, 102000, 101980, 101960, 101960, 102030, 
    102030, 102120, 102140, 102170, 102230, 102200, 102240, 102280, 102350, 
    102440, _, 102470, 102500, 102520, 102530, 102560, 102600, 102640, 
    102640, 102620, 102640, 102640, 102640, 102620, 102610, 102620, 102610, 
    102610, 102600, 102570, 102550, 102540, 102510, 102490, 102460, 102430, 
    102430, 102390, 102370, 102370, 102360, 102330, 102290, 102240, 102240, 
    102220, 102170, _, 102110, 102070, 102040, 102020, _, 101970, 101940, 
    101910, 101870, 101840, 101790, 101770, 101760, 101730, 101720, 101710, 
    101710, 101710, 101660, 101630, 101650, 101620, 101600, 101590, 101560, 
    101570, 101550, 101530, 101540, 101500, 101480, 101510, 101530, 101570, 
    _, 101610, 101650, 101660, 101670, 101670, 101680, 101660, 101610, 
    101580, 101480, 101400, 101320, 101340, 101300, 101310, 101230, 101080, 
    101020, 101000, 101010, 100960, 100960, 100900, 100840, 100810, 100740, 
    100720, 100660, 100570, 100500, 100410, _, 100490, 100390, 100330, 
    100320, 100280, 100280, 100280, 100170, 100080, 100010, 99950, 99850, 
    99750, 99720, 99660, 99650, 99600, 99570, 99580, 99520, 99570, 99560, _, 
    99570, 99530, 99530, 99520, 99500, 99470, 99510, 99510, 99520, 99630, 
    99660, 99720, 99760, 99810, 99830, 99870, _, 99890, 99890, 99870, 99860, 
    99900, 99920, 99960, 99990, 100020, 100060, 100130, 100150, 100140, 
    100150, 100180, 100220, 100250, 100280, 100270, 100280, 100290, 100310, 
    100330, 100320, 100330, 100350, 100390, 100420, 100470, 100480, 100500, 
    100510, 100530, 100550, 100570, 100580, 100580, 100590, 100610, 100630, 
    100650, 100680, 100700, 100730, 100720, 100740, 100750, 100750, 100760, 
    100780, 100800, 100860, 100900, 100920, 100940, 100950, 100980, 101010, 
    101020, 101050, 101050, 101060, 101070, 101140, 101150, 101130, 101140, 
    101130, 101120, 101110, 101120, 101130, 101100, 101080, 101060, 101090, 
    101080, 101070, 101090, 101030, 101020, 101010, 101010, 101010, 101050, 
    101010, 100970, 100910, 100890, 100840, 100820, 100820, 100760, 100720, 
    _, 100690, 100690, 100640, 100630, 100630, 100640, 100680, 100680, 
    100690, 100690, 100680, 100690, 100700, 100710, 100680, 100620, 100680, 
    100710, 100670, 100680, 100640, 100670, 100700, 100670, 100640, 100620, 
    100580, 100590, 100590, _, 100600, 100600, 100640, 100610, 100590, 
    100570, 100560, 100530, 100480, 100460, 100480, 100480, 100490, 100480, 
    100490, 100470, 100460, 100480, 100450, 100420, 100430, 100420, 100400, 
    100390, 100380, 100410, 100490, 100510, 100500, 100560, 100580, 100610, 
    100600, 100580, 100590, 100630, 100680, 100650, 100640, 100670, 100690, 
    _, 100740, 100730, 100770, 100770, 100800, 100810, 100840, 100870, 
    100910, 100930, 100910, 100920, 100920, _, 100940, 100940, 100960, 
    100970, 100990, 101000, 101010, 101030, 101060, 101060, 101070, 101090, 
    101120, 101130, 101150, 101160, 101180, 101190, 101190, 101190, 101210, 
    101200, 101170, 101180, 101180, 101200, 101210, 101210, 101180, 101180, 
    101190, 101190, 101180, 101160, 101130, 101110, 101100, 101100, 101060, 
    101060, 101020, 100990, 100950, 100930, 100880, 100850, 100820, 100760, 
    100720, 100620, 100590, 100520, 100390, 100190, 100030, 99890, 99800, _, 
    99430, 99310, 99220, 99040, 98870, 98760, 98750, 98850, 98870, 98950, 
    99010, 99040, 99050, 99070, 99070, 99050, 99080, 99080, 99070, 99090, 
    99070, 99040, 99010, 98970, 98960, 98910, 98910, 98890, 98880, 98870, 
    98850, 98840, 98850, 98870, 98880, 98890, 98900, 98900, 98890, 98870, 
    98830, 98720, 98720, 98730, 98730, 98750, 98770, 98810, 98750, 98800, 
    98830, 98850, 98770, 98790, 98760, 98820, 98880, 98820, 98860, 98940, 
    98960, 98940, 99000, 98960, 98930, 98980, 99000, 99030, _, _, 98980, _, 
    99010, 99000, 99040, 99120, _, 99140, _, 99180, 99160, 99210, 99250, 
    99250, 99280, 99280, 99280, 99300, 99320, 99400, 99440, 99440, 99450, 
    99490, 99530, 99580, 99630, 99680, 99730, 99770, 99800, 99830, 99900, 
    100000, 100040, 100090, 100140, 100180, _, 100280, 100320, 100380, 
    100430, 100480, 100500, 100550, 100590, 100640, 100670, 100700, 100710, 
    100760, 100800, 100810, 100830, 100860, 100880, 100900, 100930, 100970, 
    101000, 100970, _, 100960, 100960, 100980, 100930, 100930, 100920, 
    100970, 100960, 100940, 100900, _, 100910, 100910, 100890, 100870, _, 
    100880, 100890, 100890, 100880, _, 100850, 100850, 100830, 100790, 
    100810, 100840, 100860, 100870, 100900, 100900, 100950, 100970, 100960, 
    100960, 100940, 100900, 100900, 100880, 100910, _, 100950, 100930, 
    100920, 100870, 100810, 100810, 100770, 100750, 100670, 100620, 100550, 
    100460, 100400, 100330, 100230, 100120, 100060, 99970, 99890, 99830, 
    99780, 99730, 99700, 99650, 99650, 99630, 99650, 99670, 99700, 99720, 
    99760, 99820, 99880, 99940, 100020, 100080, 100140, 100210, 100300, 
    100350, _, 100460, 100500, 100570, 100610, 100670, 100700, 100720, _, 
    100780, 100810, 100830, 100850, 100870, 100860, 100890, 100890, 100880, 
    100880, 100880, 100870, 100860, 100870, 100880, 100860, 100850, 100860, 
    100910, 100920, 100930, 100960, 100980, 101020, 101040, 101080, 101110, 
    101140, 101150, 101190, 101200, 101250, 101280, 101310, 101330, 101360, 
    101400, 101430, 101460, 101470, 101470, 101450, 101430, 101410, 101380, 
    101360, 101320, 101300, 101310, 101300, 101280, 101280, 101260, 101250, 
    101250, 101260, 101260, _, 101230, 101210, 101180, 101160, 101100, 
    101030, 100960, 100840, 100770, 100710, 100610, _, 100400, 100300, 
    100210, 100120, 100010, 99860, _, 99550, 99370, 99250, 99140, 99110, 
    99080, 99040, 99130, 99120, 99090, 99110, 99090, 98980, 98840, 98800, 
    98810, 98750, 98750, 98780, 98800, 98850, 98850, 98970, 99070, 99210, 
    99360, 99500, 99690, 99820, 99830, 99970, 100180, 100380, 100520, 100590, 
    100670, 100740, 100830, 100910, 100980, 101050, 101120, 101190, 101260, 
    101300, 101320, 101320, 101320, 101310, 101320, 101300, 101270, 101230, 
    101170, 101120, 101090, 101030, 101020, 100990, 100960, 100940, 100880, 
    100870, 100820, 100800, 100750, 100670, 100630, 100550, 100480, 100360, 
    100280, 100240, 100190, 100150, 100090, 100050, 100010, 99980, 99940, 
    99910, 99900, _, 99840, 99840, 99830, 99820, 99800, 99800, 99830, 99750, 
    99630, 99580, 99450, 99350, 99230, 99150, 99110, 99040, 99050, 99050, 
    99130, 99220, 99330, 99470, 99600, 99750, 99870, 99980, 100070, 100180, 
    100320, 100450, 100560, 100680, 100780, 100850, 100940, 101050, 101130, 
    101210, 101290, 101370, 101410, 101460, 101500, 101500, 101500, 101510, 
    101520, 101550, 101560, 101580, 101640, 101680, 101710, 101740, 101730, 
    101750, 101730, 101710, 101640, 101590, 101550, 101480, 101400, 101330, 
    101280, 101240, 101170, 101090, 100980, _, 100860, _, 100720, 100670, 
    100640, 100640, 100670, 100710, 100750, 100800, 100860, 100910, 100990, 
    101090, 101190, 101250, 101290, 101340, 101380, 101420, 101490, 101510, 
    101530, 101580, 101590, 101620, 101630, 101640, 101680, 101750, 101760, 
    101740, 101760, 101730, 101680, 101670, 101640, 101610, 101550, 101510, 
    101480, 101430, 101420, 101420, 101420, 101420, 101450, 101470, 101450, 
    101460, 101470, 101490, 101510, 101510, 101500, 101530, 101560, 101530, 
    101520, 101510, 101480, 101460, 101390, 101340, 101350, 101280, 101250, 
    101190, 101180, 101170, 101130, 101120, 101110, 101130, 101140, 101150, 
    101140, 101160, 101190, 101210, 101240, 101240, 101270, 101310, 101340, 
    101370, 101370, 101430, 101450, 101480, 101490, 101510, 101530, 101530, 
    101540, 101590, 101600, 101630, 101660, 101640, 101650, 101640, 101680, 
    101720, 101730, 101750, 101770, 101780, 101810, 101810, 101820, 101830, 
    101860, 101870, 101900, 101900, 101920, 101910, 101930, 101930, 101940, 
    101920, 101920, 101940, 101940, 101940, 101910, 101920, 101940, 101890, 
    101850, 101880, 101900, 101840, 101780, 101770, 101720, 101690, 101670, 
    101650, 101610, 101560, 101530, 101500, 101490, 101480, 101430, 101390, 
    101370, 101380, 101340, 101330, 101300, 101310, 101340, 101350, 101320, 
    101290, 101250, 101220, 101200, 101170, 101110, 101080, 101030, 100970, 
    100900, 100870, 100810, 100740, 100670, 100580, 100500, 100420, 100380, 
    100340, 100310, 100270, 100230, 100200, 100160, 100120, 100090, 100040, 
    100010, 99980, 99970, 99980, 100010, 100030, 100030, 100000, 99980, 
    99980, 99950, 99930, 99950, 99970, 100020, 100080, 100160, 100230, 
    100290, 100350, 100410, 100510, 100550, 100600, 100650, 100710, 100780, 
    100840, 100900, 100940, 100970, 100980, 101010, 101050, 101080, 101100, 
    101120, 101110, 101140, 101140, 101190, 101210, 101190, 101210, 101200, 
    101170, 101190, 101210, 101210, 101190, 101220, 101230, 101260, 101300, 
    101320, 101360, 101410, 101450, 101510, 101560, 101580, 101600, 101620, 
    101680, 101700, 101730, 101800, 101830, 101830, 101840, 101860, 101880, 
    101900, 101920, 101930, 101940, 101920, 101930, 101920, 101910, 101890, 
    101890, 101890, 101890, 101890, 101890, 101880, 101870, 101840, 101820, 
    101810, 101770, 101750, 101730, 101690, 101670, 101650, 101610, 101590, 
    101570, 101540, 101510, 101480, 101460, 101450, 101440, 101430, 101410, 
    101400, 101400, 101400, 101400, 101400, 101410, 101420, 101430, 101450, 
    101440, 101450, 101460, 101470, 101460, 101450, 101480, 101500, 101510, 
    101510, 101510, 101510, 101510, 101550, 101540, 101550, 101540, 101540, 
    101540, 101560, 101570, 101580, 101560, 101560, 101580, 101580, 101570, 
    101550, 101550, 101550, 101540, 101530, 101490, 101470, 101460, 101440, 
    101430, 101420, 101410, 101400, 101360, 101340, 101320, 101310, 101280, 
    101290, 101260, 101260, 101210, 101220, 101190, 101150, 101120, 101030, 
    101020, 100980, 100930, 100910, 100850, 100840, 100820, 100810, 100770, 
    100760, 100740, 100710, 100700, 100690, 100680, 100670, 100660, 100650, 
    100670, 100670, 100640, 100620, 100610, 100550, 100500, 100490, 100500, 
    100500, 100510, 100480, 100410, 100370, 100370, 100340, 100410, 100430, 
    100430, 100500, 100550, 100560, 100530, 100530, 100570, 100500, 100450, 
    100390, 100390, 100370, 100390, 100370, 100320, 100280, 100320, 100270, 
    100240, 100140, 100070, 99960, 99910, 99810, 99600, 99440, 99370, 99290, 
    99320, 99280, 99000, 99030, 99030, 98920, 98770, 98610, 98550, 98330, 
    98210, 98230, 98210, 98280, 98290, 98250, 98250, 98220, 98150, 98160, 
    98160, 98190, 98160, 98150, 98090, 98040, 97980, 97990, 97930, 97930, 
    97960, 97920, 97950, 97970, 97950, 97920, 97920, 97900, 97880, 97860, 
    97830, 97830, 97850, 97860, 97880, 97890, 97900, 97890, 97880, 97900, 
    97890, 97870, 97870, 97860, 97860, 97870, 97890, 97920, 97950, 97950, 
    97970, 98030, 98080, 98120, 98150, 98170, 98220, 98230, 98290, 98330, 
    98390, 98410, 98440, 98460, 98480, 98500, 98520, 98540, 98550, 98560, 
    98590, 98620, 98620, 98650, 98650, 98670, 98680, 98680, 98690, 98700, 
    98700, 98730, 98770, 98820, 98880, 98910, 98930, 98940, 98970, 99000, 
    99030, 99050, 99070, 99100, 99110, 99140, 99170, 99160, 99170, 99180, 
    99200, 99210, 99230, 99250, 99270, 99280, 99300, 99340, 99390, 99430, 
    99460, 99470, 99470, 99470, 99480, 99460, 99460, 99480, 99490, 99520, 
    99560, 99600, 99610, 99640, 99650, 99680, 99700, 99720, 99740, 99800, 
    99830, 99870, 99910, 99940, 99960, 99990, 99990, 99990, 100000, 99980, 
    99990, 99990, 100000, 100000, 100010, 100000, 99980, 99950, 99950, 99940, 
    99940, 99970, 100000, 100050, 100090, 100120, 100160, 100210, 100280, 
    100300, 100320, 100330, 100360, 100340, 100310, 100310, 100290, 100200, 
    100180, 100180, 100090, 100050, 100020, 99940, 99860, 99800, 99790, 
    99690, 99730, 99710, 99660, 99750, 99690, 99630, 99570, 99620, 99660, 
    99670, 99650, 99680, 99680, 99640, 99630, 99540, 99550, 99550, 99540, 
    99560, 99680, 99690, 99740, 99750, 99770, 99790, 99890, 99910, 99930, 
    99950, 99950, 99950, 99950, 99980, 100010, 100030, 100050, 100090, 
    100100, 100090, 100050, 100070, 100050, 100050, 100000, 100040, 100070, 
    100100, 100070, 100070, 100140, 100210, 100210, 100260, 100250, 100280, 
    100260, 100240, 100190, 100130, 100120, 100080, 100070, 100060, 100070, 
    100100, 100120, 100100, 100120, 100080, 100110, 100100, 100100, 100110, 
    100110, 100120, 100110, 100100, 100070, 100060, 100020, 99970, 99920, 
    99870, 99830, 99790, 99750, 99690, 99620, 99530, 99430, 99340, 99240, 
    99160, 99110, 99050, 99010, 98960, 98920, 98870, 98820, 98770, 98710, 
    98680, 98640, 98600, 98540, 98530, 98520, 98510, 98510, 98490, 98510, 
    98510, 98500, 98500, 98480, 98490, 98520, 98560, 98600, 98640, 98650, 
    98700, 98700, 98740, 98770, 98750, 98680, 98680, 98670, 98690, 98700, 
    98740, 98720, 98700, 98700, 98670, 98650, 98640, 98610, 98600, 98580, 
    98580, 98590, 98590, 98590, 98620, 98620, 98630, 98640, 98650, 98670, 
    98690, 98680, 98700, 98680, 98690, 98680, 98650, 98610, 98600, 98540, 
    98500, 98480, 98450, 98430, 98440, 98460, 98470, 98470, 98480, 98500, 
    98520, 98510, 98520, 98540, 98540, 98560, 98590, 98610, 98650, 98660, 
    98650, 98650, 98650, 98650, 98640, 98630, 98640, 98660, 98670, 98680, 
    98700, 98720, 98720, 98720, 98710, 98700, 98690, 98680, 98680, 98690, 
    98680, 98680, 98690, 98680, 98700, 98720, 98740, 98750, 98760, 98780, 
    98820, 98850, 98870, 98910, 98960, 99030, 99100, 99140, 99230, 99260, 
    99300, 99340, 99360, 99410, 99460, 99510, 99570, 99680, 99760, 99830, 
    99890, 100010, 100070, 100160, 100250, 100310, 100410, 100520, 100600, 
    100690, 100770, 100860, 100950, 100990, 101060, 101130, 101210, 101270, 
    101340, 101400, 101480, 101530, 101550, 101600, 101610, 101610, 101610, 
    101610, 101600, 101620, 101620, 101620, 101600, 101630, 101630, 101630, 
    101630, 101660, 101700, 101710, 101730, 101750, 101790, 101830, 101860, 
    101860, 101860, 101850, 101840, 101820, 101760, 101750, 101690, 101620, 
    101610, 101560, 101500, 101480, 101430, 101400, 101390, 101300, 101220, 
    101170, 101100, 101020, 100910, 100850, 100770, 100650, 100620, 100550, 
    100450, 100340, 100300, 100300, 100240, 100130, 100080, 100030, 99950, 
    99890, 99820, 99780, 99680, 99730, 99730, 99670, 99590, 99560, 99590, 
    99570, 99600, 99620, 99640, 99630, 99560, 99410, 99470, 99530, 99470, 
    99410, 99380, 99360, 99380, 99390, 99340, 99370, 99380, 99410, 99420, 
    99460, 99490, 99510, 99550, 99610, 99620, 99620, 99650, 99710, 99710, 
    99720, 99750, 99770, 99780, 99830, 99850, 99890, 99920, 99950, 99990, 
    100010, 100030, 100050, 100090, 100110, 100170, 100190, 100200, 100240, 
    100270, 100270, 100310, 100350, 100360, 100380, 100400, 100410, 100460, 
    100470, 100470, 100490, 100530, 100530, 100520, 100510, 100500, 100490, 
    100450, 100420, 100390, 100330, 100300, 100270, 100260, 100230, 100200, 
    100170, 100150, 100100, 100060, 100030, 100000, 99990, 99970, 99950, 
    99950, 99970, 99970, 99950, 99940, 99940, 99920, 99920, 99920, 99930, 
    99930, 99950, 99980, 100010, 100030, 100040, 100070, 100090, 100130, 
    100160, 100190, 100220, 100250, 100320, 100380, 100450, 100530, 100570, 
    100630, 100680, 100730, 100800, 100850, 100880, 100920, 100950, 101010, 
    101060, 101110, 101130, 101140, 101170, 101160, 101150, 101140, 101160, 
    101190, 101190, 101170, 101150, 101140, 101100, 101060, 101020, 100990, 
    100940, 100900, 100850, 100760, 100710, 100670, 100620, 100540, 100500, 
    100410, 100350, 100290, 100280, 100240, 100210, 100170, 100130, 100100, 
    100030, 99940, 99880, 99810, 99760, 99730, 99700, 99670, 99620, 99550, 
    99500, 99430, 99400, 99360, 99350, 99330, 99300, 99300, 99330, 99350, 
    99380, 99410, 99450, 99480, 99510, 99500, 99530, 99540, 99550, 99600, 
    99660, 99690, 99730, 99750, 99800, 99870, 99920, 99960, 100000, 100040, 
    100080, 100150, 100230, 100300, 100370, 100450, 100500, 100560, 100610, 
    100660, 100700, 100770, 100800, 100830, 100890, 100940, 100990, 101030, 
    101080, 101120, 101140, 101150, 101180, 101220, 101260, 101260, 101310, 
    101350, 101410, 101470, 101510, 101550, 101560, 101580, 101590, 101620, 
    101600, 101610, 101650, 101680, 101700, 101740, 101750, 101770, 101780, 
    101780, 101810, 101840, 101860, 101870, 101870, 101880, 101940, 101960, 
    102000, 102040, 102080, 102100, 102140, 102160, 102180, 102250, 102250, 
    102300, 102340, 102360, 102430, 102480, 102500, 102520, 102550, 102570, 
    102620, 102660, 102700, 102730, 102770, 102780, 102800, 102840, 102840, 
    102860, 102870, 102860, 102860, 102840, 102810, 102750, 102690, 102640, 
    102550, 102510, 102490, 102470, 102440, 102390, 102390, 102380, 102350, 
    102350, 102340, 102340, 102300, 102270, 102210, 102100, 102020, 101980, 
    101940, 101910, 101860, 101810, 101780, 101750, 101680, 101630, 101590, 
    101510, 101490, 101440, 101470, 101470, 101480, 101450, 101410, 101400, 
    101410, 101400, 101380, 101350, 101360, 101330, 101300, 101280, 101240, 
    101190, 101160, 101100, 101110, 101060, 101000, 100950, 100910, 100860, 
    100830, 100760, 100670, 100600, 100540, 100430, 100380, 100310, 100310, 
    100320, 100330, 100320, 100330, 100310, 100320, 100310, 100310, 100300, 
    100310, 100330, 100350, 100330, 100380, 100410, 100520, 100630, 100710, 
    100770, 100830, 100960, 101130, 101290, 101480, 101540, 101690, 101800, 
    101840, 101980, 102060, 102090, 102120, 102150, 102180, 102180, 102170, 
    102140, 102090, 102000, 101960, 101870, 101790, 101710, 101630, 101570, 
    101500, 101440, 101380, 101320, 101240, 101180, 101120, 101070, 101020, 
    100970, 100950, 100940, 100920, 100880, 100850, 100850, 1008.4, 1008.6, 
    1008.8, 1009.4, 1010.2, 1010.9, 1011.2, 1011.6, 1013.1, 1013.9, 1014.2, 
    1014.8, 1015.1, 1015.5, 1015.8, 1016.4, 1016.8, 1017.1, 1017.2, 1017.6, 
    1018, 1018.2, 1018.5, 1018.8, 1018.7, 1018.6, 1018.3, 1017.9, 1017.3, 
    1018.2, 1018.7, 1019.2, 1019.9, 1020.4, 1020.2, 1020.5, 1020.7, 1021.2, 
    1021.7, 1021.7, 1021.6, 1021.8, 1021.9, 1022, 1022, 1022, 1021.9, 1021.9, 
    1021.8, 1021.5, 1021.3, 1021.1, 1021, 1021, 1020.9, 1021, 1020.8, 1020.7, 
    1020.3, 1020.3, 1020.2, 1019.7, 1019.5, 1019.2, 1018.9, 1018.8, 1018.7, 
    1018.7, 1018.5, 1018.2, 1018.2, 1017.7, 1017.3, 1017.1, 1016.8, 1016.4, 
    1016.3, 1016.1, 1015.6, 1015.3, 1015, 1014.7, 1014.6, 1014.3, 1013.9, 
    1013.3, 1012.6, 1012.3, 1011.8, 1010.7, 1010.2, 1009.7, 1009.2, 1008.6, 
    1008.5, 1007.9, 1007.8, 1007.3, 1007, 1006.9, 1006.3, 1006.2, 1005.9, 
    1005.9, 1006.2, 1007.5, 1007.4, 1007.6, 1007.9, 1008.3, 1008.3, 1008.6, 
    1008.9, 1009, 1009.3, 1009.9, 1010.5, 1011, 1011.5, 1012.2, 1012.6, 
    1012.9, 1013.3, 1013.8, 1014.3, 1014.9, 1015.3, 1015.9, 1016.5, 1017.3, 
    1017.8, 1018.6, 1018.9, 1019.3, 1019.6, 1019.9, 1020.2, 1020.5, 1021.3, 
    1022, 1022.5, 1023, 1023.6, 1024.2, 1024.7, 1025.2, 1025.5, 1026.3, 
    1026.8, 1027.3, 1027.6, 1028, 1028.6, 1029.4, 1029.9, 1030.2, 1030.5, 
    1030.7, 1030.9, 1031.1, 1031.2, 1031.4, 1031.7, 1031.9, 1032.2, 1032.4, 
    1032.5, 1032.6, 1032.9, 1032.8, 1032.7, 1032.7, 1032.7, 1032.6, 1032.4, 
    1032.4, 1032.7, 1032.7, 1032.4, 1032.3, 1032.1, 1032, 1031.7, 1031.1, 
    1030.9, 1030.4, 1029.8, 1029.7, 1029.3, 1029.1, 1028.8, 1028.4, 1027.9, 
    1027.8, 1027.4, 1026.9, 1026.2, 1025.7, 1025.5, 1025.1, 1025.1, 1024.5, 
    1024.2, 1023.6, 1022.7, 1022, 1021.5, 1021, 1020.2, 1019.7, 1019.2, 
    1018.8, 1018.3, 1017.9, 1017.4, 1016.7, 1016, 1015.3, 1014.7, 1014.4, 
    1013.4, 1012.9, 1012.2, 1011.6, 1011.7, 1010.8, 1010.5, 1010.1, 1009.3, 
    1008.8, 1008.1, 1007.3, 1007.1, 1006.1, 1005.6, 1004.9, 1004.6, 1004.2, 
    1003.8, 1003.4, 1002.6, 1002.5, 1002.7, 1002.6, 1002.2, 1002.1, 1002.3, 
    1002.6, 1003.1, 1003.4, 1003.6, 1002.8, 1002.7, 1003.2, 1003.3, 1002.6, 
    1002, 1001.8, 1001.2, 1001.6, 1001.4, 1001.5, 1001.8, 1001.6, 1001.3, 
    1000.6, 1000.4, 1000.1, 999.5, 999, 998.8, 998.4, 997.8, 996.7, 996.6, 
    995.7, 995.2, 994.2, 993.6, 991.6, 991.8, 992.5, 993.5, 993.7, 994.4, 
    996.1, 998, 999.4, 1000.3, 1001.5, 1003, 1003.8, 1005.1, 1006.1, 1007, 
    1007.8, 1008.2, 1008.9, 1009.4, 1009.9, 1010.1, 1010.6, 1011.1, 1011.6, 
    1012, 1012.5, 1013, 1013.7, 1014, 1014.5, 1015, 1015.2, 1015.3, 1015.3, 
    1015.6, 1015.8, 1015.7, 1015.8, 1015.1, 1015.1, 1015, 1014.8, 1013.9, 
    1013.3, 1012.7, 1011.6, 1010.7, 1010.1, 1009.6, 1009.1, 1008.6, 1007.7, 
    1007.3, 1006.9, 1006, 1005.4, 1004.8, 1004.1, 1003.9, 1004.3, 1003.7, 
    1004, 1004.2, 1004.8, 1005, 1005.6, 1005.9, 1006, 1006.2, 1006.5, 1006.6, 
    1006.8, 1007.3, 1007.5, 1007.9, 1008.1, 1008.9, 1009.2, 1009.6, 1010.1, 
    1010.5, 1010.8, 1011.5, 1012.1, 1012.9, 1013.5, 1014.2, 1015.1, 1015.8, 
    1016.3, 1016.1, 1016.7, 1016.9, 1017.5, 1017.6, 1018.1, 1018.5, 1018.7, 
    1018.7, 1019.1, 1019.4, 1019.6, 1019.9, 1020.2, 1020.2, 1020.4, 1021, 
    1021.5, 1021.9, 1022, 1022.1, 1022.5, 1023.3, 1023.5, 1024.7, 1025.5, 
    1025.5, 1025.4, 1026.4, 1026.3, 1026.2, 1025.1, 1025.1, 1025.4, 1024.4, 
    1024.3, 1023, 1021.9, 1020.4, 1019.3, 1018.2, 1016.8, 1015.4, 1013.7, 
    1012.2, 1010.7, 1010.1, 1008.4, 1007.6, 1006.7, 1005.7, 1005.4, 1004.8, 
    1004.8, 1004.2, 1004, 1002.9, 1002.1, 1000.8, 1000.2, 998.5, 996.9, 
    994.9, 993.6, 992.2, 990.6, 989.7, 989.1, 989.4, 989.3, 989.6, 990.7, 
    990.4, 990.3, 990.6, 990.4, 990.1, 989.7, 992.3, 996.5, 999.8, 1002.4, 
    1004.5, 1006.9, 1008.9, 1010.8, 1011.9, 1012.5, 1013.2, 1013.9, 1015, 
    1015.3, 1015.4, 1015.8, 1016.5, 1016.9, 1017.8, 1018.8, 1020, 1020.1, 
    1019.7, 1019.4, 1019.2, 1018.7, 1018.7, 1019.9, 1019.4, 1018.8, 1018.6, 
    1018, 1017.6, 1016.9, 1016.3, 1015.7, 1015.3, 1014.8, 1014.5, 1014.4, 
    1014, 1013.5, 1013.6, 1013.5, 1013.6, 1013.1, 1013.6, 1014.2, 1014.9, 
    1015.8, 1016.2, 1017, 1017.5, 1017.4, 1017.6, 1017.7, 1018, 1018.1, 1018, 
    1017.9, 1017.5, 1017.4, 1017.3, 1016.9, 1016.5, 1016.1, 1015.8, 1015.5, 
    1014.5, 1014, 1013.3, 1012.6, 1011.9, 1011, 1010, 1009.5, 1009, 1008, 
    1007.3, 1006.5, 1005.5, 1005.1, 1004.6, 1004.2, 1003.8, 1003.9, 1003.9, 
    1003.8, 1004.2, 1004.7, 1004.9, 1005.3, 1005.7, 1005.9, 1005.9, 1006.4, 
    1006.5, 1006.7, 1006.7, 1006.9, 1007.1, 1007.4, 1007.5, 1007.3, 1007.4, 
    1007.7, 1007.8, 1007.8, 1007.7, 1008, 1008.2, 1008.2, 1008.4, 1008.7, 
    1008.9, 1009.2, 1009.3, 1009.6, 1009.8, 1009.8, 1010.1, 1010, 1010.2, 
    1010.4, 1010.6, 1011, 1011.3, 1011.6, 1011.6, 1011.7, 1011.8, 1011.9, 
    1011.9, 1012, 1012.6, 1012.9, 1013.2, 1013.5, 1013.7, 1013.6, 1013.6, 
    1013.6, 1013.6, 1013.7, 1013.8, 1013.9, 1013.9, 1014.1, 1014.2, 1014.3, 
    1014.4, 1014.4, 1014.4, 1014.8, 1015.1, 1015.3, 1015.3, 1015.5, 1015.9, 
    1016.3, 1016.5, 1016.6, 1016.8, 1016.6, 1016.8, 1016.7, 1016.6, 1016.6, 
    1016.3, 1016.3, 1016.3, 1016.1, 1016.1, 1016.3, 1016.2, 1016, 1015.6, 
    1015.2, 1015, 1014.7, 1014.3, 1013.8, 1013.6, 1013.3, 1013, 1012.7, 
    1012.3, 1011.8, 1011.1, 1010.5, 1009.7, 1009.4, 1008.3, 1008, 1007.3, 
    1006.5, 1006.2, 1005.3, 1004.5, 1004.2, 1003.2, 1003, 1002.8, 1002.7, 
    1002.6, 1002.2, 1002.3, 1003.3, 1004, 1004.3, 1003.2, 1003.6, 1003.7, 
    1005.4, 1005.2, 1005.4, 1005.5, 1005.4, 1005.8, 1006.3, 1006.8, 1007.3, 
    1007.1, 1007.1, 1007.5, 1007.2, 1007, 1007.2, 1007.5, 1007.4, 1007.3, 
    1007, 1007.3, 1007.6, 1007.9, 1007.6, 1007.3, 1007, 1007.2, 1006.7, 
    1006.6, 1006.4, 1005.2, 1005.3, 1007.1, 1007.8, 1007.7, 1008, 1007.2, 
    1007.2, 1006.3, 1006.9, 1006.8, 1007.4, 1007.8, 1008, 1009.3, 1010.3, 
    1011.1, 1011.8, 1012.7, 1012, 1012.1, 1012.5, 1012, 1012, 1011.8, 1012.6, 
    1012.7, 1012.7, 1012.5, 1012.7, 1012.3, 1012.1, 1011.9, 1011.7, 1011.3, 
    1011.4, 1011.6, 1011.3, 1011.5, 1011.4, 1011.5, 1011.4, 1011, 1010.9, 
    1010.6, 1010.3, 1009.8, 1009.5, 1008.7, 1008.1, 1007.7, 1007.2, 1006.5, 
    1005.1, 1003.2, 1002.8, 1002.1, 1002.1, 1001.2, 1000.6, 999.2, 999.8, 
    999.5, 999.2, 999.1, 998.9, 998.7, 998.3, 997.7, 997, 996.2, 996.3, 
    996.6, 996.8, 996.7, 997.1, 997.7, 997.8, 997.9, 998, 998.3, 998.5, 
    998.4, 998.5, 998.6, 998.9, 998.9, 999.2, 999.3, 999.3, 999.5, 998.8, 
    998.5, 998.3, 997.5, 997.7, 997.2, 997, 996.9, 996.5, 996.9, 997.2, 
    997.3, 996.6, 996.1, 996.7, 996.6, 996.7, 996.6, 996.6, 996.5, 996.3, 
    996.5, 996.2, 996.3, 995.8, 996.3, 996.8, 996.9, 997.2, 997.2, 997.7, 
    997.8, 998.2, 998.2, 998.1, 997.8, 997.2, 996.7, 996.5, 996.2, 995.8, 
    995.7, 995.7, 995.6, 995.6, 995.4, 995.1, 994.7, 994.6, 994.5, 994.2, 
    993.9, 993.7, 993.7, 993.3, 993.2, 993.4, 993.9, 994.2, 994.8, 995.1, 
    995.4, 995.5, 995.6, 995.7, 995.9, 996.3, 996.7, 997, 997.2, 997.2, 
    997.2, 997.2, 997.1, 997, 996.8, 996.8, 996.5, 996, 995.9, 996, 995.6, 
    996.2, 996, 995.5, 995.4, 994.6, 993.7, 993.5, 993.7, 993.2, 992.8, 993, 
    992.8, 992.9, 992.8, 992.1, 991.8, 991.5, 991.6, 992.5, 991.5, 991.2, 
    991.2, 991.5, 991.2, 991.2, 991.5, 991.1, 990.9, 990.8, 990.6, 990.4, 
    990.3, 990.1, 990.1, 990, 990.2, 990.2, 990.1, 990.1, 990.2, 990.4, 
    990.5, 990.5, 990.6, 990.8, 991, 991.3, 991.4, 991.4, 991.4, 991.4, 
    991.6, 991.8, 992.1, 992.6, 992.9, 993.2, 993.8, 994.2, 994.5, 994.9, 
    995.1, 995.4, 995.9, 996.2, 996.6, 997, 997.1, 997.5, 997.8, 998.2, 
    998.8, 999.1, 999.3, 999.8, 1000.3, 1000.8, 1001.4, 1001.9, 1002.5, 
    1003.2, 1004.5, 1005.1, 1005.7, 1006.3, 1006.5, 1006.4, 1006.1, 1006, 
    1005.7, 1005.4, 1005.1, 1004.5, 1003.8, 1003.8, 1003.5, 1004.1, 1004.1, 
    1003.7, 1003.7, 1003.9, 1003.6, 1003, 1002.3, 1001.3, 1000.4, 999.2, 
    998.3, 997.1, 995.4, 994.3, 993.2, 992.3, 992.4, 993.4, 993.9, 994.9, 
    996.5, 997.4, 998, 999.3, 1000.5, 1001.2, 1001.3, 1001.4, 1001.4, 1001.9, 
    1002.5, 1003.2, 1003.8, 1004.5, 1005.2, 1005.3, 1005.3, 1005.4, 1005.1, 
    1004.7, 1003.9, 1003, 1001.7, 1000.9, 1000.2, 999.3, 998.4, 997.5, 996, 
    994.5, 993, 991.9, 990.5, 989.7, 988.8, 988.4, 988.4, 989.1, 989.7, 
    990.4, 990.9, 991.7, 992.2, 992.5, 992.7, 992.8, 992.8, 993, 993.4, 
    993.2, 993.2, 993.3, 993.6, 994.1, 994.9, 995.8, 996.8, 997.4, 998.4, 
    999.1, 999.9, 1000.5, 1001, 1001.6, 1001.6, 1001.5, 1001.3, 1001.1, 
    1000.9, 1000.6, 1000.6, 1000.6, 1000.3, 1000.2, 1000.1, 999.3, 998.4, 
    997.3, 996.2, 995.9, 994.9, 994.3, 993.6, 993.3, 992.8, 992.2, 992, 
    992.1, 992.2, 992.1, 992.2, 992.2, 992.4, 991.9, 991.6, 991.1, 990.9, 
    990, 989.7, 990.9, 991.9, 993, 993.7, 994.5, 995.4, 996.2, 996.7, 997.4, 
    996.8, 998, 998.4, 997.9, 998, 997.6, 996.6, 995.8, 995.5, 995.1, 994.7, 
    994.8, 994.8, 995, 995.4, 995.6, 996.6, 996.7, 998.1, 999.2, 1000, 
    1001.6, 1002.2, 1003.4, 1005.1, 1006.6, 1007.6, 1008.4, 1009.9, 1011.1, 
    1012.1, 1013.3, 1014.7, 1015.9, 1016.9, 1018, 1019.1, 1020.6, 1020.9, 
    1021.5, 1022.2, 1022.5, 1023, 1023.1, 1023.3, 1023.4, 1023.5, 1023.5, 
    1023.7, 1023.7, 1023.7, 1023.7, 1024, 1023.7, 1023.5, 1022.5, 1021.7, 
    1020.8, 1020.3, 1019.2, 1017.9, 1016.7, 1015.9, 1014.9, 1013.9, 1013, 
    1012.4, 1011.7, 1011.2, 1010.7, 1010.4, 1009.7, 1009.5, 1009.5, 1009.2, 
    1008.9, 1008.8, 1009, 1008.9, 1008.8, 1008.9, 1009.2, 1008.5, 1008.5, 
    1008.9, 1008.8, 1009.1, 1009.3, 1009.7, 1009.6, 1010.2, 1010.7, 1011, 
    1011.3, 1011.3, 1011.5, 1011.8, 1012.1, 1012.6, 1013.1, 1012.8, 1013.2, 
    1013.2, 1013.4, 1013, 1013, 1012.7, 1012.6, 1012.4, 1012.2, 1011.6, 1011, 
    1010.6, 1010.2, 1009.8, 1009.5, 1009.2, 1008.8, 1008.3, 1008, 1007.5, 
    1007.1, 1006.7, 1006.3, 1005.8, 1005.2, 1004.8, 1004.2, 1003.7, 1003.1, 
    1002.7, 1002.2, 1002, 1001.6, 1001, 1000.2, 999.6, 998.9, 998.2, 998.1, 
    997.7, 997.5, 997.2, 996.6, 996, 995.4, 994.3, 993.1, 991.1, 989.3, 
    986.7, 985.9, 983.9, 981.6, 981.5, 981.3, 980.5, 979.9, 979.2, 978.7, 
    978.6, 979.2, 979.6, 980, 981, 982, 983.9, 985.5, 986.8, 988.6, 990.2, 
    991.6, 992.1, 993.1, 994, 994.8, 995.7, 996.6, 997.6, 998.5, 998.7, 
    999.2, 999.9, 1000.1, 1000.7, 1001.3, 1001.3, 1001.4, 1001.3, 1000.9, 
    1000.6, 1000, 1000, 999.7, 999.9, 1000.2, 1000.3, 1000, 1000.6, 1000.1, 
    1000, 1000.2, 1000.1, 1000, 1000.2, 1000.6, 1000.5, 1001.2, 1001.3, 
    1001.3, 1001.4, 1001.5, 1001.6, 1001.9, 1002, 1002.3, 1002.5, 1002.8, 
    1002.9, 1002.9, 1003.1, 1003.2, 1003.2, 1003.1, 1003.1, 1002.7, 1002.7, 
    1002.1, 1002.2, 1002.1, 1002, 1001.5, 1001.4, 1001.3, 1000.9, 1000.6, 
    1000.3, 1000, 999.9, 999.7, 999.6, 999.3, 999.2, 998.6, 998.5, 998.6, 
    998.5, 998.1, 997.7, 997.8, 997.8, 997.5, 997.2, 997.4, 997.4, 997.4, 
    997.7, 997.8, 998.3, 998.8, 999.1, 998.8, 998.1, 998.4, 998.5, 999, 
    999.2, 999.4, 999.6, 999.7, 999.9, 1000.5, 1000.7, 1000.9, 1001.1, 
    1001.8, 1001.7, 1001.8, 1002, 1001.5, 1001.2, 1000.8, 1000.9, 1000.6, 
    1000.3, 1000, 999.4, 999.2, 998.7, 998.4, 997.9, 997.4, 996.7, 996, 
    995.3, 994.7, 994.2, 993.5, 992.9, 992.4, 992, 991.6, 991.1, 990.8, 
    990.4, 990.1, 990.1, 990.2, 990.5, 990.3, 990.5, 990.6, 991, 991.1, 
    991.6, 991.9, 992, 991.8, 991.1, 990.7, 990.4, 990.6, 990.7, 991, 991.1, 
    991.4, 991.6, 992.2, 992.6, 993.2, 994.8, 995.9, 996.3, 996.4, 996.9, 
    997.2, 997.3, 998.4, 999.3, 999.5, 1000, 1000.2, 1000.8, 1000.8, 1000.8, 
    1000.6, 1000.3, 1000.3, 1000.6, 1001.1, 1001.7, 1001.8, 1002.3, 1002.8, 
    1002.9, 1003, 1002.8, 1002.4, 1002.2, 1002, 1001.9, 1001.7, 1001.3, 
    1001.2, 1001, 1000.7, 1000.5, 1000, 999.8, 999.5, 999.4, 999.2, 999, 999, 
    999.1, 999, 998.8, 998.5, 998.5, 998.9, 999.1, 999.4, 999.4, 999.8, 
    1000.4, 1001, 1001.2, 1001.4, 1001.9, 1002.2, 1002.9, 1003.4, 1003.5, 
    1003.2, 1003.4, 1003.9, 1004.3, 1005.1, 1006.1, 1006.9, 1007.3, 1007.7, 
    1008, 1008.5, 1009, 1009.5, 1009.8, 1010.4, 1011, 1011.7, 1012.5, 1013, 
    1013.3, 1013.5, 1013.2, 1013.2, 1013.5, 1014.4, 1014.5, 1014.4, 1014, 
    1013.9, 1013.5, 1012.9, 1012.1, 1011.5, 1010.9, 1010.2, 1009.2, 1008.8, 
    1008.1, 1007.7, 1007.4, 1007, 1006.5, 1006.4, 1006.2, 1006, 1006.1, 
    1006.2, 1005.8, 1005.8, 1005.8, 1005.6, 1005.5, 1005.2, 1005, 1004.7, 
    1004.3, 1004.5, 1004.1, 1004.1, 1004, 1004.3, 1004.8, 1005.2, 1005.5, 
    1006.2, 1006.4, 1006.9, 1007.2, 1008, 1008.4, 1008.3, 1008.6, 1008.4, 
    1008.3, 1008.4, 1008.9, 1009.1, 1009.3, 1009.1, 1009, 1009.4, 1009.5, 
    1009.6, 1009.7, 1009.9, 1009.9, 1009.9, 1009.8, 1009.6, 1009.9, 1009.9, 
    1009.4, 1009.6, 1009.2, 1009, 1009.2, 1008.7, 1008.5, 1007.9, 1007.7, 
    1007.3, 1007.6, 1007.7, 1007.4, 1007.3, 1007.8, 1007.5, 1008, 1008.1, 
    1008.5, 1007.9, 1008.2, 1008.4, 1008.5, 1008.5, 1008.3, 1008.4, 1008.3, 
    1007.9, 1007.9, 1007.9, 1007, 1007.4, 1007.7, 1007.6, 1007.4, 1007.6, 
    1007.4, 1007.1, 1007.1, 1006.6, 1006.9, 1006.9, 1006.3, 1007.1, 1007.3, 
    1007.1, 1007.4, 1007.6, 1008, 1008.3, 1008.9, 1009, 1009.4, 1011, 1011.8, 
    1013.2, 1013.4, 1012.3, 1012.1, 1012.5, 1014.7, 1015.5, 1016.1, 1016.6, 
    1016.7, 1016.6, 1016.6, 1016.7, 1017.1, 1017.3, 1017.4, 1017.5, 1017.4, 
    1017.4, 1017.3, 1017.2, 1017.1, 1017, 1016.6, 1016.2, 1015.7, 1015, 
    1014.3, 1014, 1013.5, 1012.8, 1011.9, 1011, 1010.2, 1009.2, 1008.5, 
    1008.1, 1007.7, 1007.3, 1006.9, 1006.5, 1005.9, 1005.2, 1004.9, 1004.2, 
    1004.2, 1003.6, 1003.2, 1002.7, 1002.4, 1001.7, 1001, 1000.7, 1000.5, 
    1000.8, 1000, 999.1, 998.6, 1000.2, 1000, 999.2, 999.6, 999.6, 999.5, 
    998.5, 997, 996.9, 996.4, 995.4, 993.3, 994.1, 995.9, 997.3, 1000.7, 
    1002.1, 1002.9, 1003.4, 1002.8, 1002.7, 1002.4, 1002.3, 1001.7, 1002.4, 
    1002.1, 1002, 1001.6, 1002.5, 1002.9, 1001.9, 1001.7, 1004, 1005.1, 
    1005.2, 1004.8, 1005.1, 1004.2, 1003.9, 1003.6, 1003.5, 1003.7, 1004.8, 
    1004.6, 1003.9, 1004, 1004, 1003.9, 1003.4, 1003.1, 1002.8, 1002.4, 1002, 
    1001.7, 1001.5, 1000.8, 1000, 999.4, 998.9, 998.4, 997.8, 996.8, 996.9, 
    996.6, 996.6, 996.7, 996.4, 995.7, 995.7, 995.3, 993.7, 993.2, 993.9, 
    994.5, 994.3, 994.6, 995.2, 995.6, 995.5, 995.4, 995.3, 995.3, 995.5, 
    995.1, 995.3, 995.3, 995.4, 995.6, 995.7, 996, 996, 996.1, 996.2, 996.7, 
    997, 997.3, 997.7, 997.7, 998.1, 998.5, 998.9, 999.1, 999.2, 999.7, 
    999.9, 1000.3, 1000.6, 1000.9, 1001.1, 1001.3, 1001, 1001.5, 1002, 
    1001.7, 1001.9, 1002.1, 1002.4, 1002.5, 1002.5, 1002.4, 1002.2, 1001.9, 
    1001.9, 1002, 1002.3, 1002.6, 1002.5, 1002.6, 1002.4, 1002.5, 1002.6, 
    1002.8, 1002.8, 1002.6, 1002.6, 1002.6, 1002.6, 1002.7, 1002.7, 1002.7, 
    1003, 1002.4, 1002.6, 1002.9, 1002.9, 1002.9, 1002.2, 1001.7, 1001.5, 
    1002.2, 1002.4, 1003.5, 1003.5, 1003.4, 1003.1, 1002.2, 1004, 1004.1, 
    1003.7, 1004.1, 1004.5, 1004.6, 1004.8, 1004.7, 1004.6, 1004.2, 1004.3, 
    1004.3, 1004.5, 1004.5, 1004.3, 1004.5, 1004.8, 1005, 1004.9, 1004.7, 
    1004.7, 1004.6, 1004.6, 1005.1, 1004.8, 1004.8, 1004.8, 1004.6, 1004.3, 
    1004.2, 1004.1, 1004.2, 1003.8, 1003.7, 1003.6, 1003.5, 1003.3, 1002.9, 
    1002.6, 1002.5, 1002.4, 1002.4, 1002.3, 1002.7, 1002.2, 1002, _, 1001.3, 
    1001.2, 1001, 1001, 1000.4, 1000.5, 1000.8, 1000.6, 1000.1, 1000.7, 
    1000.3, 1000.5, 1000.6, 1000.6, 1000.7, 1000.6, 1001, 1001.3, 1001.8, 
    1001.7, 1002, 1002.1, 1002.4, 1002.6, 1002.9, 1003.4, _, 1003.8, _, 
    1004.5, 1005.1, 1005.4, 1006.3, 1006.7, 1007.2, 1007.4, 1007.3, 1007.9, 
    1008.2, 1008.2, 1008.8, 1009.3, 1009.8, 1010, _, 1010.7, 1010.9, 1011.4, 
    1011.7, 1012, 1012, 1012.4, 1012.9, 1013.2, 1013.6, 1013.8, 1014.3, 
    1014.7, 1015, 1015, 1015.3, 1015.5, 1016.2, 1016.6, 1017.2, 1017.5, 
    1017.6, 1017.7, 1017.6, 1017.7, 1018, 1018.3, 1018.7, 1019, 1019.1, 
    1019.2, 1019.4, 1019.3, 1020.1, 1020.5, 1020.8, 1021, 1021, 1021.3, 
    1021.5, 1021.6, 1022, 1022.3, 1022.5, 1023.2, 1023.6, 1023.6, 1024.1, 
    1024.6, 1024.7, 1024.8, 1025.2, 1025.3, 1025.7, 1025.8, 1026.1, 1026.4, 
    1026.7, 1027, 1026.9, 1027, 1026.9, 1027.1, 1027.1, 1027.2, 1027.3, 
    1027.4, 1027.5, 1027.7, 1027.6, 1027.4, 1027.2, 1027.1, 1027, 1026.9, 
    1026.6, 1026.5, 1026.3, 1026.3, 1026, 1025.7, 1025.6, 1025.4, 1025.3, 
    1025.2, 1025.1, 1024.9, 1024.8, 1024.7, 1024.5, 1024.6, 1024.7, 1024.7, 
    1024.4, 1024.4, 1024.3, 1024.3, 1024.2, 1024.1, 1024.1, 1023.9, 1023.9, 
    1024, 1024, 1024.1, 1024.1, 1023.9, 1023.4, 1023, 1023.2, 1023, 1022.5, 
    1022.8, 1022.4, 1022.3, 1022.3, 1022.3, 1022.2, 1022, 1021.8, 1021.5, 
    1021.2, 1021.3, 1021.2, 1021.3, 1021.4, 1021.2, 1021.3, 1021.3, 1021.6, 
    1021.4, 1021.7, 1021.8, 1022.1, 1021.9, 1021.7, 1021.4, 1021.5, 1021.4, 
    1020.7, 1020.4, 1020.6, 1020.5, 1020.1, 1019.8, 1019.4, 1019.1, 1018.9, 
    1019.1, 1018.8, 1018.5, 1018.1, 1017.8, 1017.7, 1017.3, 1017, 1016.7, 
    1016.5, 1016, 1015.8, 1015.4, 1014.9, 1014.6, 1014.5, 1014.9, 1014.8, 
    1014.8, 1014.8, 1014.8, 1015.1, 1015, 1015, 1015, 1015.2, 1015.4, 1015.6, 
    1016.1, 1016.4, 1016.6, 1016.8, 1016.8, 1017, 1017.1, 1017.3, 1017.3, 
    1017.2, 1017.3, 1017.5, 1017.7, 1018, 1017.9, 1018.1, 1018.1, 1018.3, 
    1018.7, 1019.1, 1019.3, 1019.6, 1019.8, 1020.3, 1020.5, 1020.7, 1021, 
    1021.1, 1020.9, 1020.9, 1021.1, 1021.1, 1021.3, _, 1021.5, 1021.8, 
    1022.2, 1022.4, 1022.3, _, 1022.2, 1022, 1021.9, 1021.6, 1021.3, 1020.9, 
    1020.7, 1020.3, 1020.4, 1020, 1019.7, 1019.5, 1019.3, 1019.4, 1019.1, 
    1019.1, 1018.8, 1018.8, 1018.8, 1018.9, 1019, 1019, 1019.1, 1019.3, 
    1018.9, 1018.5, 1018.3, 1018.3, 1018.1, 1018, 1017.7, 1017.7, 1017.6, 
    1017.6, 1017.8, 1017.3, 1017.2, 1017.1, 1017.1, 1017.3, 1017.4, 1017.6, 
    1018.1, 1018.8, 1019.6, 1020.4, 1021, 1021.7, 1022.3, 1022.7, 1023.3, 
    1023.8, 1024.2, 1024.9, 1025.5, 1025.9, 1026.5, 1026.9, 1027.4, 1027.6, 
    1027.8, 1028, 1028.3, 1028.5, 1028.8, 1029, 1029.5, 1029.7, 1030.1, 
    1030.4, 1030.8, 1031, 1031.1, 1031.2, 1031.3, 1031.5, 1031.5, 1032, 
    1032.2, 1032.3, 1032.5, 1032.8, 1032.9, 1032.8, 1032.8, 1032.8, 1032.9, 
    1033, 1033, 1032.9, 1033.1, 1033.4, 1033.5, 1033.8, 1034, 1033.9, 1033.6, 
    1033.5, 1033.4, 1033.2, 1033, 1032.8, 1032.7, 1032.5, 1032.1, 1031.8, 
    1031.5, 1031.2, 1030.6, 1029.9, 1029.6, 1029.3, 1029, 1028.3, 1028.3, 
    1028.4, 1028.5, 1028.4, 1028.4, 1028.2, 1028, 1027.9, 1027.8, 1027.5, 
    1027.6, 1027.5, 1027.5, 1027.4, 1027.8, 1027.5, 1027.4, 1027.3, 1027.1, 
    1026.9, 1026.4, 1026, 1025.8, 1025.3, 1025.2, 1024.6, 1025.1, 1024.9, 
    1025, 1025.2, 1024.8, 1024.7, 1024.2, 1024, 1023.8, 1023.6, 1023.2, 
    1023.1, 1023.2, 1023.1, 1023, 1022.7, 1022.7, 1022.5, 1022.7, 1022.6, 
    1022.6, 1022.7, 1022.7, 1023, 1023.2, 1023.5, 1023.7, 1023.8, 1023.9, 
    1023.9, 1024.1, 1024.2, 1024.1, 1024.1, 1024.4, 1024.4, 1024.3, 1024.1, 
    1024.2, 1024, 1023.9, 1023.8, 1023.5, 1023.3, 1023.1, 1022.9, 1022.8, 
    1022.8, 1022.7, 1022.3, 1022, 1021.4, 1021, 1020.5, 1020.2, 1019.9, 
    1019.5, 1019, 1018.6, 1018.7, 1018.2, 1017.8, 1017.3, 1016.9, 1016.4, 
    1016, 1015.7, 1015.5, 1015.2, 1014.9, 1014.6, 1014.4, 1014.3, 1014, 
    1013.7, 1013.9, 1013.5, 1013.1, 1012.9, 1012.5, 1012.4, 1012.1, 1011.9, 
    1011.8, 1011.4, 1011.2, 1010.8, 1010, 1009.9, 1009.7, 1009.5, 1009.4, 
    1009.2, 1009, 1009.1, 1009.1, 1009.1, 1009.1, 1008.5, 1008.2, 1008.2, 
    1007.5, 1007.3, 1007, 1006.9, 1007.6, 1007.8, 1007.3, 1007.2, 1006.7, 
    1006, 1006.2, 1005.9, 1005.4, 1005, 1004.1, 1003.3, 1003.1, 1002.7, 
    1002.4, 1002.7, 1002.6, 1002.2, 1002.2, 1001.9, 1002.1, 1002, 1002.5, 
    1002.4, 1002.1, 1001.8, 1001.5, 1001.4, 1001.7, 1001.9, 1002.3, 1002, 
    1001.2, 1001.1, 1000.7, 1000.4, 1000.2, 999.7, 999.1, 999.1, 999.5, 
    999.5, 1000, 1000.4, 1000.6, 1000.3, 1000.5, 1000.9, 1001.2, 1001.3, 
    1001.2, 1001.3, 1000.7, 1000.3, 1000.1, 1000.6, 1001.1, 1001.6, 1002, 
    1002.2, 1002.7, 1003.1, 1003.6, 1004.1, 1004.6, 1004.8, 1005, 1005.2, 
    1005.2, 1005.6, 1005.9, 1006.1, 1006.2, 1006.2, 1006.6, 1006.9, 1006.8, 
    1007, 1007.1, 1007.2, 1007.3, 1007.5, 1007.4, 1007.4, 1007.1, 1006.9, 
    1006.8, 1006.5, 1006.3, 1005.9, 1005.7, 1005.8, 1005.8, 1005.7, 1005.7, 
    1005.6, 1005.3, 1005.3, 1005, 1004.7, 1004.2, 1004, 1003.6, 1003.3, 
    1003.3, 1002.8, 1002.4, 1002.1, 1001.8, 1001.8, 1002, 1002, 1001.5, 
    1001.3, 1001.1, 1001, 1000.7, 1000.7, 1000.4, 999.9, 999.6, 999.3, 999.1, 
    998.9, 998.7, 998.8, 998.6, 998.2, 998.1, 997.8, 997.7, 997.4, 997.2, 
    997, 997.1, 996.9, 996.8, 996.5, 996.1, 995.6, 995.3, 995.4, 995.2, 
    995.3, 995, 995, 995.2, 995.3, 995.5, 995.9, 996.2, 996.5, 997.3, 997.3, 
    997.7, 997.9, 998.5, 998.7, 999.1, 999.9, 1000, 1000.4, 1000.6, 1000.8, 
    1001.3, 1000.9, 1000.8, 1000.3, 1000.1, 1000.1, 1000.2, 1001.6, 1002.5, 
    1003.3, 1003.3, 1003.3, 1003.7, 1004, 1003.6, 1003.6, 1003.5, 1003.2, 
    1003.4, 1003.8, 1003.8, 1003.9, 1003.9, 1003.9, 1003.8, 1003.6, 1003.4, 
    1003.3, 1003.1, 1003.2, 1003.7, 1004.2, 1004.6, 1004.5, 1004.9, 1005.2, 
    1005.3, 1005.4, 1005.3, 1005.5, 1005.7, 1006, 1006.3, 1006.9, 1007.4, 
    1007.8, 1008.2, 1008.8, 1008.8, 1008.5, 1008.9, 1009.2, 1009.5, 1009.6, 
    1009.7, 1009.8, 1010, 1010.4, 1009.5, 1009.2, 1009.1, 1009.6, 1009.2, 
    1008.7, 1009.3, 1009.7, 1009.4, 1009.8, 1009.6, 1009.3, 1008.8, 1008.6, 
    1008.3, 1008.1, 1007.7, 1007.8, 1007.3, 1006.6, 1006.2, 1005.4, 1004.2, 
    1004.3, 1004.1, 1003.9, 1002.9, 1002.3, 1001.9, 1001.5, 1000.7, 1000.2, 
    999.8, 999.6, 999.3, 999, 998.8, 998.6, 998.2, 997.6, 997.1, 996.4, 
    996.4, 996, 995.6, 995.4, 995.4, 995.5, 995.7, 995.9, 996.1, 996.2, 
    996.7, 997.1, 997.2, 997.7, 998.1, 998.8, 999.5, 999.7, 999.9, 1000.1, 
    1000.2, 1000.9, 1001, 1001.1, 1001.3, 1001.4, 1001.5, 1001.7, 1002, 
    1002.4, 1002.7, 1002.9, 1003, 1003.5, 1003.7, 1004, 1005, 1005.1, 1005.3, 
    1005.9, 1006.4, 1006.8, 1006.3, 1006.8, 1006.5, 1006.1, 1005.3, 1004, 
    1002.5, 1001.2, 999.6, 998.6, 997.5, 996.3, 995.1, 993.9, 993, 991.6, 
    991.1, 990.4, 990, 990.1, 989.7, 989.2, 988.8, 988, 986.7, 985.5, 984.9, 
    983.9, 983, 981.8, 981.7, 981.6, 981.3, 981.6, 981.8, 982.1, 982.1, 
    982.7, 983.2, 983.7, 984.7, 985.2, 986.4, 987, 988.3, 989.4, 990.3, 
    991.1, 992.4, 993.1, 994, 994.5, 996.1, 996.2, 996.9, 997.2, 997.9, 
    997.8, 998.4, 998.3, 998.4, 998.5, 997.7, 997.8, 997.8, 997.3, 996.6, 
    996.2, 996.1, 996.2, 996.4, 996.5, 996.4, 996.4, 997.1, 997.8, 998, 
    999.5, 1000.8, 1002.2, 1003.1, 1003.6, 1004.3, 1005.2, 1006.3, 1007.1, 
    1008.4, 1009.3, 1009.8, 1009.6, 1010.1, 1010.1, 1010.4, 1010.4, 1010.9, 
    1010.9, 1010.8, 1011.1, 1011.1, 1010.8, 1010.7, 1010.3, 1009.7, 1009.7, 
    1009.6, 1009.3, 1009.7, 1009.7, 1009.3, 1009.3, 1009.4, 1008.6, 1008.9, 
    1009, 1008.9, 1008.9, 1009.4, 1009.3, 1009.9, 1009.9, 1009.3, 1009.8, 
    1009.8, 1009.8, 1009.9, 1008.9, 1008.4, 1007.7, 1008.1, 1007.9, 1007.6, 
    1007.9, 1007.7, 1007.6, 1007.4, 1006.8, 1006.8, 1007.2, 1007, 1007, 
    1006.3, 1005.6, 1006.9, 1006.8, 1006.4, 1006.2, 1006.2, 1006.4, 1006.3, 
    1005.7, 1003.6, 1003, 1004.2, 1004.7, 1004.9, 1004, 1003.8, 1003.3, 
    1003.6, 1003.6, 1003, 1003.1, 1003.6, 1003.9, 1005.4, 1006.3, 1006.5, 
    1006.8, 1007.3, 1007.9, 1008.3, 1008.4, 1009.4, 1009.1, 1009.4, 1009.4, 
    1009.7, 1009.9, 1010.6, 1010.3, 1010.3, 1010.1, 1010.2, 1010.4, 1010.3, 
    1009.5, 1009.2, 1008.6, 1007.3, _, 1006.3, 1005.8, 1005.1, 1004.8, 
    1004.6, 1003.7, 1003.1, 1002.5, 1001.4, 1000.4, 1000.2, 999.4, 999.7, 
    998.6, 997.5, 997.3, 996.8, 996.7, 996.3, 995.8, 995.2, 995.3 ;

 wind_speed_10m = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 35, 30.9, 36, 26.2, 35, 30.9, 33.4, 3.6, 30.9, 3.6, 
    50.4, 26.2, 3.6, 3.6, 30.9, 17, 49.4, 30.9, 28.8, 33.4, 40.6, 35, 26.2, 
    35, 39.1, 40.6, 3.1, 5.3, 5.5, 5.9, 6.4, 6.4, 6.6, 5.9, 5.7, 6, 6.2, 6.8, 
    7.1, 7.2, 7.2, 7.4, 6.4, 6.5, 6.5, 6.9, 7.2, 7.2, 7.4, 7.3, 7.6, 7.7, 
    7.6, 7.4, 9.2, 11, 10, 9.8, 10.1, 7.4, 10.3, 9.2, 8.3, 9, 8.9, 9.6, 8.8, 
    7.5, 9.1, 7.4, 8, 7.2, 9.8, 8, 8.9, 8.6, 7.8, 8.2, 7.5, 7.3, 8.4, 5.7, 
    8.7, 7.8, 9.3, 8.2, 8.2, 8.4, 8.7, 9.2, 9.7, 8.9, 8.4, 9.2, 9, 8, 7.2, 
    8.7, 6.6, 8, 8, 6.9, 7.3, 7.4, 8.2, 7.9, 8.4, 10, 9.8, 8.9, 10.6, 9, 9, 
    8.8, 7, 7.3, 6.8, 7.2, 8.4, 8, 8.2, 7.6, 8.3, 7.9, 8, 9.3, 8.5, 8.7, 9, 
    9.5, 8.7, 5.8, 6.6, 6.9, 6.5, 7, 6.8, 7.3, 6.3, 7.5, 6.7, 5.8, 6.3, 6.3, 
    7, 6.5, 6, 6.9, 8, 6.8, 6.8, 6.4, 7.4, 7.3, 6.4, 6.3, 5.9, 5.3, 5.6, 5.6, 
    2.9, 4.1, 4.7, 5.1, 4.4, 2.2, 1, 1.2, 0.9, 0, 0.2, 1.8, 0.4, 0, 0, 0, 
    0.7, 0, 0, 0, 0.3, 0.1, 0.1, 0.9, 3.1, 1, 1.4, 1.8, 1.9, 0.9, 7.6, 2.9, 
    2.3, 9.9, 11.3, 11.1, 5.1, 6.4, 4, 3.6, 1.4, 1.5, 1.4, 6.5, 1.1, 2.2, 
    0.6, 1.2, 2, 3.1, 3.3, 2.3, 0.6, 2.2, 1.8, 2, 1, 1, 1.7, 2.1, 1.9, 1.6, 
    1.7, 2.1, 1.4, 0, 1, 0.6, 0.9, 0.3, 0.5, 0.1, 0, 0, 1, 0, 0.2, 0.8, 1.1, 
    2.9, 2.1, 0.3, 2.2, 0.6, 1.7, 0.1, 1, 2.2, 5.4, 5.4, 3.2, 0.8, 4.6, 5.3, 
    3.5, 4.7, 6.4, 4.6, 6.4, 5.9, 5.4, 4.7, 4.7, 3, 4, 2.4, 6.1, 4.8, 5.2, 
    6.2, 5.5, 5.3, 4.6, 3.1, 3, 1.7, 0.4, 0.1, 0, 2.9, 4.5, 3.5, 3.6, 2.9, 
    2.8, 2.9, 4.6, 4.3, 2.9, 3.7, 4, 3.2, 3.6, 2.6, 3.7, 3.7, 4.6, 4, 4.6, 
    3.8, 4.3, 3.5, 4.2, 3.1, 1.9, 1.8, 2.2, 2.5, 3.1, 2.1, 2.5, 3.2, 3.5, 
    3.1, 3.4, 3.4, 3.2, 4.1, 4.4, 5.5, 3.9, 4.4, 4.6, 4.3, 3.7, 4.1, 4.1, 3, 
    4.8, 5, 4.8, 2.8, 5.5, 5, 5.8, 5.3, 7.5, 5.3, 5.1, 4.5, 6.4, 6, 5.5, 5.3, 
    4.8, 4.6, 4.1, 2.9, 3, 2.2, 2.4, 2.4, 0.8, 0, 0.7, 0.9, 0.5, 0.5, 0.8, 
    0.7, 1.9, 1.4, 1.8, 0.7, 2.6, 3.1, 2.8, 4, 3.8, 4.3, 5.2, 6.2, 6.5, 5.6, 
    5.3, 5.5, 6, 5.3, 5.8, 5.9, 6.3, 6.8, 6.9, 7, 7.7, 7.8, 7.9, 6.7, 7.7, 
    7.6, 8.9, 8, 8.9, 7.1, 7.1, 7.6, 7.3, 6.9, 7.1, 7, 7.1, 7, 7.1, 6.5, 7.4, 
    5.9, 5.2, 3.2, 2.8, 2.6, 3.7, 2.8, 1.6, 1.1, 3.4, 3.3, 3.8, 3.1, 4.6, 
    4.8, 4.2, 4.6, 1.9, 3.1, 4.4, 5.7, 2.3, 4.1, 4.6, 3.4, 1.4, 0.8, 0.3, 
    1.9, 3.1, 4.8, 5.2, 6.3, 6.9, 4.6, 1.2, 3, 4.8, 4.8, 4.6, 6, 6.9, 5, 4.9, 
    5.2, 4.9, 2, 0.6, 0, 0, 3, 3.3, 5.4, 8.7, 8.6, 9.5, 11.4, 12.2, 13.4, 
    10.8, 10.7, 9, 8, 8.8, 9.2, 8.3, 8.3, 6.3, 7.8, 7.9, 9, 9.6, 8.4, 8.6, 
    9.6, 9.7, 9.7, 10.8, 11.5, 10.5, 12.3, 12.2, 9.1, 8.4, 8.5, 7.5, 6.9, 
    6.8, 6, 6.9, 5.4, 6.2, 4.9, 5.2, 4.1, 3.6, 3.2, 4.1, 4, 5.4, 5.4, 3.5, 
    2.1, 0.4, 5.6, 8.8, 7.1, 7.1, 7.2, 6.7, 6.6, 5.5, 5.7, 7.6, 1.4, 3.8, 
    3.6, 5.2, 3.3, 2.9, 3.3, 3.3, 1.7, 9.1, 9.3, 11.4, 8.9, 12.1, 11.8, 18.8, 
    19, 18.9, 18.9, 18.6, 18.4, 19.1, 17.5, 15.7, 13.4, 10.2, 8.1, 8.3, 6.6, 
    6.5, 8.1, 8.3, 8, 7, 6, 4.1, 5.7, 6.9, 4.4, 3.6, 4.6, 2.1, 1.2, 2, 3.4, 
    1, 0.8, 0.4, 3.5, 4.8, 6.9, 3.3, 5.5, 1.2, 0.9, 0.2, 0.7, 0, 0.6, 1.4, 1, 
    0.3, 1, 1.5, 0.4, 0.5, 1.1, 0.4, 1.6, 1.9, 1.3, 0.8, 1.2, 0, 0.1, 0, 2.1, 
    2.1, 4.5, 4.5, 6.8, 6.5, 6.7, 5.6, 8.5, 8.5, 6.9, 7.3, 8.3, 9.7, 12.4, 
    7.2, 4.8, 2.6, 9, 6.9, 5.8, 6.8, 6.1, 7, 7.3, 7.1, 5.4, 5.8, 3.6, 2.2, 
    1.2, 2.5, 4, 3.5, 3.1, 1.7, 1, 0, 0, 0, 0, 0.1, 0.8, 0.1, 0.4, 1.3, 1.9, 
    1.1, 2, 2.6, 1.7, 2, 0.9, 1.3, 0.5, 1.5, 2.8, 4, 3.1, 5.5, 6.2, 7.4, 8.2, 
    9.7, 9.4, 7.2, 8.5, 5.8, 3.6, 7.1, 5.1, 6.2, 9.6, 9.4, 7.3, 10, 8.7, 7.6, 
    7.2, 8.2, 8.4, 7.6, 7.2, 7.4, 5.4, 4.6, 3.4, 6.2, 6.1, 3.6, 6.2, 6.1, 
    8.1, 9.9, 10.1, 7.1, 9, 10.8, 12, 6.7, 18.9, 19.3, 13.6, 4.5, 15.3, 12, 
    11.1, 9.8, 10.3, 10.8, 9.2, 8.6, 10, 9.8, 11.1, 9.9, 8.4, 7.1, 7.3, 8.4, 
    8.9, 8.9, 9.5, 8.3, 8.7, 8.4, 9.1, 9.4, 10.8, 9.5, 8.4, 10.7, 10.8, 10.2, 
    10.1, 9.1, 9.8, 9.4, 9.1, 7.7, 7.3, 7.6, 5.7, 8.1, 7.4, 6.3, 1.9, 0.6, 
    2.2, 0.7, 1.2, 1.3, 2.9, 2.2, 0, 0.4, 1.1, 1.1, 1, 1.7, 1.2, 0.7, 1.4, 0, 
    0.1, 0, 0.4, 3.7, 2, 4.3, 6, 5.7, 6.2, 7.2, 6.2, 5.5, 5.9, 7, 7.2, 8.4, 
    9.2, 9.7, 10.3, 10.2, 9.8, 12.1, 11.7, 11.4, 12.4, 12.3, 11.5, 9.7, 10.3, 
    9.9, 9.6, 8.6, 6.9, 8.2, 7.4, 5.5, 3.6, 2, 1.3, 1.5, 1.7, 1.5, 4.4, 6.5, 
    7.5, 7, 8.1, 9.3, 10, 9.2, 8.4, 9.3, 8.3, 7, 7.7, 5.9, 4.2, 3.6, 3.6, 
    4.8, 4.5, 2.8, 0, 3.7, 10.3, 7.5, 6.2, 7.2, 7.9, 6.2, 6, 6.3, 6.1, 6.7, 
    7.2, 5.5, 0.9, 3.7, 0.3, 0.4, 2.1, 1.8, 2.5, 2.6, 3.2, 3.7, 3.7, 3, 4.8, 
    2.8, 3.6, 3.5, 4.5, 4.6, 5.7, 7.5, 7.9, 8, 8.3, 10.3, 9.7, 11.8, 11.7, 
    10.8, 9.5, 10.5, 7.4, 7.7, 9.8, 9.3, 8.5, 9, 8.5, 8.4, 7.2, 7.2, 6.7, 
    7.9, 7.4, 7.3, 5.1, 7.8, 7.8, 7.9, 7.9, 7.8, 7.2, 6.8, 6.6, 6.8, 6.5, 
    7.8, 7.1, 7.4, 7.9, 7.1, 8.2, 5.4, 7.1, 6.8, 7, 7.1, 6.9, 6, 6.4, 7.7, 
    7.5, 6.9, 7.4, 8.8, 8.8, 7.3, 8.8, 7.1, 7.2, 6.2, 5.8, 7, 6.7, 8, 6, 8, 
    8.6, 6.2, 7.8, 6.5, 6.6, 6.9, 7.1, 6.2, 6.2, 4.7, 5, 4.1, 3.2, 2.7, 3.1, 
    3, 1.4, 3.6, 4.1, 4.3, 4.9, 5.6, 5.1, 4.5, 4.7, 4.8, 6.8, 6.5, 7.8, 6.9, 
    7.4, 7.2, 6.3, 6.1, 7.8, 8, 6.8, 5.7, 7, 7.8, 7.9, 7.6, 7.7, 6.9, 6.5, 
    6.9, 8.1, 9.4, 9.4, 8.9, 10.7, 12.5, 12.9, 11.1, 10.8, 10.8, 9.9, 10.6, 
    10.5, 10.9, 11.2, 8.8, 9.1, 8, 7.5, 7.3, 8.4, 8.2, 6.8, 7.5, 6.5, 7.6, 
    9.1, 8.1, 10.3, 10.5, 11.7, 10.2, 9.8, 10.4, 10.7, 9.8, 10, 11.7, 11.8, 
    11.9, 11, 7.5, 7.7, 5.9, 6.1, 6, 5, 5.4, 5.7, 5.6, 6.1, 6.2, 6.5, 3.5, 
    7.1, 8.7, 8.6, 6.4, 6.7, 7.1, 8.6, 8.2, 7.7, 7.8, 7.5, 9.1, 8.4, 8.6, 
    8.6, 7.5, 7.8, 8.2, 5.2, 5.1, 10.3, 9.7, 11.1, 10.3, 11.4, 11.6, 8.5, 
    8.7, 10, 9.7, 9.2, 8.6, 7.9, 6.4, 6.9, 6, 1.6, 1.5, 0, 0, 0, 0, 0.5, 0.1, 
    2, 2.5, 7.3, 7, 7.8, 8.1, 8, 7.4, 6.6, 8.7, 7.5, 10.5, 10.6, 11.4, 11.2, 
    10.3, 8.2, 8.7, 9.2, 10.6, 11.2, 9.9, 9.5, 8.5, 8.8, 8.4, 7.5, 8.7, 6.8, 
    7.2, 5.4, 7.4, 8.2, 9.6, 7.8, 6.1, 5.8, 7.4, 8.3, 7.9, 7.2, 6.7, 6, 7, 
    7.1, 7.3, 4.5, 3.1, 4, 3.4, 1.9, 2, 2.4, 1.9, 2.8, 4.8, 6.4, 6.8, 7.6, 
    8.8, 11.6, 10.9, 13.4, 13.1, 13.5, 14.7, 15.4, 15.4, 15.5, 15.7, 15.4, 
    14.2, 12.4, 11.5, 13.2, 10.3, 11.8, 12, 10.8, 7.3, 12.1, 8, 10.5, 6, 4.4, 
    2.1, 3.1, 0.6, 1.3, 3.5, 4.1, 4.3, 3.2, 4.6, 4.9, 4, 1.2, 4, 2.5, 2.5, 
    4.4, 3.7, 3.3, 4.3, 2.4, 7.1, 6, 1.4, 1.1, 3.4, 5.5, 6.1, 5.5, 6.6, 6.2, 
    6, 9.7, 9.9, 8.9, 1.7, 2.6, 6.1, 4.6, 2.8, 1.2, 5.1, 5.8, 4.1, 4.5, 3.2, 
    3.5, 4.6, 5.6, 3, 3.4, 3.1, 3.5, 2.4, 1.9, 4.5, 2.6, 3, 2.5, 3.1, 4.4, 
    7.2, 5.4, 4.9, 6.9, 5.1, 4.5, 5.1, 6.3, 7.6, 9.4, 9.6, 10.8, 10.4, 8.3, 
    8.6, 9.3, 8, 8.2, 5.8, 5.2, 5.3, 6.7, 7, 6.9, 7.5, 5.4, 4.4, 7.1, 3.7, 
    6.7, 4.9, 7.1, 5.9, 5.5, 5.2, 6.2, 6, 6.4, 6.6, 6.6, 6.1, 6.5, 6.3, 7, 8, 
    7.8, 10.2, 11.1, 12.2, 10.7, 12.9, 10.3, 12.5, 13.6, 11.7, 13.1, 14.2, 
    12.6, 12.6, 12.1, 10.6, 10.7, 7.9, 8.6, 6.8, 5.2, 2.9, 0.6, 4.1, 7.3, 
    7.3, 5, 6.8, 9.9, 9.9, 11.2, 12.4, 9.6, 10.8, 10, 12.3, 10.4, 12.4, 11.5, 
    10.7, 11.1, 9.1, 8.8, 12.3, 12.1, 11, 13.8, 13.7, 14.6, 15.6, 13.3, 12.5, 
    12.9, 13.4, 13.1, 12.3, 14.4, 11.8, 13.6, 12.4, 12.3, 12.6, 12.1, 14, 
    14.9, 13.8, 12.4, 12.6, 11.4, 9.5, 8.4, 10, 10.3, 8.2, 9.3, 8.3, 8.6, 
    7.1, 10.1, 9.6, 8.5, 6.9, 6.7, 6.8, 6.9, 6.8, 6.7, 6.1, 5.4, 5.4, 6.5, 
    6.6, 5.6, 5.3, 7.5, 7.2, 6.4, 4.7, 6, 5.6, 4.8, 6, 6.1, 5, 5.3, 6.2, 6.8, 
    7.2, 6.7, 5.2, 4.1, 3.6, 2.7, 3.3, 3.3, 7.3, 9.1, 5.1, 6.5, 5.9, 8.4, 
    10.4, 7.7, 6.4, 7.4, 5.9, 7.5, 8.7, 6.4, 7.9, 5.8, 7.7, 8.2, 9.6, 9.6, 
    11.6, 12.6, 13.7, 13.6, 15.5, 12.8, 11.4, 9.5, 10.9, 11, 11.2, 12.4, 
    12.2, 11.4, 11.3, 11.1, 12, 12.9, 10.3, 10.2, 10.8, 11.8, 9.7, 10.5, 
    10.3, 10.6, 8.9, 7, 6.2, 5.4, 5.2, 4.3, 2.7, 3.2, 3.6, 2.2, 4.5, 6.5, 
    7.6, 10.7, 12.1, 13.5, 15.7, 17.5, 18.6, 18.2, 18.7, 21.3, 22.3, 21.8, 
    24.9, 23, 13.9, 5.8, 7.3, 4.2, 4, 6.1, 6.3, 4.1, 4.6, 4.8, 5, 2.7, 1.5, 
    1.5, 1.3, 2.3, 3.3, 5.1, 8.5, 9.1, 9.7, 9.9, 11.7, 14, 13.1, 13.1, 15.6, 
    15.8, 14.4, 14.8, 15.9, 15.5, 16.3, 17.9, 16.3, 13.4, 14.6, 13, 14.7, 
    16.6, 16.2, 16.2, 18.6, 18.6, 11.7, 16.5, 13.4, 13.3, 12.2, 14.5, 13.3, 
    _, 10.8, 10.8, 12.5, 14.9, 15.9, 14.4, 12.2, 10.9, 11.9, 13.1, 16.4, 
    14.4, 10.6, 13.8, 13.7, 14.6, 14.1, 12.7, 11, 12.7, 12.9, 14.9, 13.7, 
    14.4, 14.6, 12.9, 16, 15.2, 10.7, 11.1, 11.6, 11.9, 8.9, 9.8, 7.5, 8.5, 
    7.6, 7.4, 6.6, 4.9, 5.3, 5.2, 6.6, 5.9, 4.7, 4.4, 8.4, 8.7, 8.4, 6, 8.6, 
    7, 8.2, 1, 2.2, 3.3, 3.6, 6.8, 3.9, 3.8, 10.6, 9.6, 9.5, 11.2, 9.9, 9.5, 
    8.9, 9.4, 6.8, 7.5, 7.8, 5.3, 8.9, 4.6, 8, 8.3, 8.5, 11.1, 5.7, 7, 10.9, 
    11.3, 11.6, 11, 11, 11.7, 8.4, 10.3, 9.1, 9.1, 7.4, 6.9, 5.5, 6.5, 4.6, 
    4.8, 4, 5.5, 3.5, 3.6, 2.8, 5.5, 3.5, 2.9, 4.3, 5.2, 5.9, 8, 8.3, 8.8, 
    7.8, 5.5, 6.3, 5.1, 6.6, 3.9, 4.8, 4.6, 3, 3.5, 4.6, 5.9, 6.4, 7.7, 6.9, 
    6, 5.1, 3.5, 3.1, 5.4, 4.8, 3.5, 4.3, 3.4, 4.2, 4.2, 4.6, 4.3, 6.8, 7.1, 
    5.6, 6.6, 7.1, 5, 9.7, 8.7, 7, 9.3, 7.6, 10, 10.5, 12.8, 10.7, 12.5, 
    13.1, 14.5, 14.2, 13.7, 16, 17.4, 18.1, 17.3, 18.8, 20.7, 20.6, 21, 17.3, 
    21.4, 19.6, 16.9, 15.1, 13.1, 12.9, 10.8, 9, 7.8, 8.1, 7.5, 10, 7.6, 4.6, 
    2.3, 0.7, 2.7, 4.3, 7, 7, 10, 12, 12.6, 15.3, 13.9, 12.8, 14.7, 13.4, 15, 
    14, 13.6, 13.5, 11.1, 11.1, 10.5, 9.7, 10, 12.6, 9.8, 10.1, 8.9, 11.2, 
    7.9, 10, 8.7, 8.2, 7.3, 7.2, 4.1, 6.6, 6.1, 2.8, 1.2, 0.4, 3.6, 2.8, 3.8, 
    5.4, 7.6, 7, 8.6, 9.3, 9.3, 7.5, 6.2, 7.5, 7.3, 5, 4.9, 4.8, 5.6, 6.1, 
    7.5, 7.2, 7.5, 8.1, 7.8, 9.5, 10.6, 12.2, 14.2, 12.9, 14.2, 14, 15.8, 
    16.1, 16.3, 16.2, 16.4, 17, 17.4, 16.8, 14.7, 13.6, 13.2, 11.7, 11.7, 
    11.3, 12.2, 9.4, 7.9, 10.8, 12.2, 15.1, 11, 15.3, 11.8, 9.9, 9.8, 7.4, 
    6.5, 7.1, 9.1, 7.9, 5.7, 4.9, 3.5, 1.6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12.2, 13.3, 15.8, 11.9, 14.9, 16.8, 16, 17.4, 
    19.4, 18.1, 20.4, 19.9, 16.8, 18.7, 19.7, 22, 20.8, 23.9, 23.1, 22.9, 
    22.4, 23.7, 22, 22.8, 22.4, 20.6, 20.7, 22.1, 21.7, 20.1, 21.6, 19.6, 
    21.8, 18.3, 18.2, 16.5, 15.7, 16.6, 15.7, 15.9, 15.7, 18.1, 17.5, 17.8, 
    20.2, 19.8, 19, 19.2, 19.4, 20.3, 20, 18.2, 19.3, 19.9, 21.9, 22.3, 19.4, 
    25.1, 23, 22.7, 21.3, 20.5, 20.2, 18.3, 13.7, 18.8, 16.8, 17, 16.3, 13.8, 
    12.1, 12, 9.3, 10.2, 9.8, 8, 8.2, 7.3, 7.7, 5, 7.6, 4.3, 5.8, 6.6, 7.8, 
    7.8, 10.1, 9.5, 10.5, 9.2, 9.7, 6.4, 7.8, 6.3, 5.3, 6, 5.2, 5.1, 7.3, 
    5.9, 6.3, 7.3, 7.4, 4.6, 3.9, 2.9, 3, 2.6, 3.3, 3.5, 2.4, 2.8, 2.6, 1.5, 
    1.5, 1.1, 1.1, 1.5, 2.2, 3.5, 4.7, 3.9, 7.6, 6.1, 7.4, 9.1, 8.8, 8.1, 
    8.6, 9.4, 10.3, 9, 9.6, 6.4, 9, 9.4, 9.9, 11, 10.4, 11, 11.5, 13.6, 16.7, 
    14.9, 14.5, 15.9, 15.5, 14.1, 13.9, 13.3, 13.9, 12.6, 12.1, 12, 10.9, 
    9.2, 8.2, 7.9, 7.7, 6.9, 5.8, 6.7, 6.8, 6.5, 7.2, 7.4, 7.7, 8.7, 6.5, 
    5.7, 9.8, 9.5, 9.8, 10.1, 9.4, 9.1, 9.7, 7.4, 7.3, 10.4, 9.1, 10.2, 4, 
    3.8, 9.5, 7.7, 8.2, 4.9, 4.9, 5.9, 9.8, 8, 12.1, 10.3, 11.1, 11.8, 12.3, 
    12.6, 11.3, 12.7, 13.8, 15.2, 15.5, 14.7, 14.1, 13.3, 12.5, 8.9, 11.3, 
    8.6, 8.4, 8.1, 0.2, 0.5, 0, 0.1, 1.4, 2.3, 3.3, 4, 14.1, 18, 17.8, 18.6, 
    16, 16, 15.5, 14.6, 14.1, 17.6, 19.8, 15.7, 15, 16, 15.5, 14.9, 16, 14.9, 
    13.7, 14.5, 13.3, 11.6, 11, 9.2, 8.9, 11.4, 11.7, 11.1, 6.3, 8.7, 8.2, 
    5.9, 5.2, 5.6, 7.4, 6.9, 7.9, 6.9, 9.3, 8.2, 7.7, 6.6, 7.1, 6.6, 7.2, 
    5.9, 5.1, 3.8, 4.3, 7.1, 8.9, 11.3, 13, 14.4, 17.2, 16.3, 5, 4.1, 3.9, 
    3.2, 2.7, 2.6, 1.7, 1.1, 1.3, 1.1, 1, 2.9, 3.6, 4.2, 4.8, 5.2, 5.4, 4.9, 
    4.8, 4.5, 5.1, 6.4, 7, 8.1, 7.4, 7, 7, 6.7, 6.5, 6.4, 6.3, 6, 5.7, 5.3, 
    4.9, 4.9, 5, 5.4, 5.6, 5.7, 5.7, 5.5, 5.4, 5.2, 5.3, 5.4, 5.3, 4.9, 5.2, 
    5.3, 5.2, 5.2, 5.3, 5.7, 5.8, 6.1, 6.2, 6.1, 5.9, 6, 6.1, 6, 6.2, 6.3, 
    6.4, 6.6, 6.7, 6.7, 6.9, 7, 6.8, 6.5, 6.8, 6.8, 6.6, 6.6, 6.5, 7.6, 7.7, 
    7.6, 7.8, 7.6, 7.4, 7.9, 7.9, 7.7, 7.5, 7.4, 7.2, 7.3, 7.1, 7.1, 6.9, 
    6.7, 6.4, 5.5, 5, 4.8, 4.9, 4.8, 4.8, 5.1, 5.1, 5.3, 5.2, 4.8, 4.2, 4.4, 
    4.5, 4.5, 4.4, 4.4, 4.3, 4, 3.8, 3.3, 3.1, 3.1, 2.8, 1.8, 1.6, 1.5, 1.8, 
    2.2, 2.6, 2.9, 3.6, 4.4, 4.9, 5.6, 6.1, 6.3, 6.8, 7.2, 8, 8.6, 9.3, 9.5, 
    9.7, 9.7, 10.1, 10.2, 10.3, 9.6, 9.2, 9.3, 9.8, 10.1, 10.2, 10.1, 11.1, 
    11.9, 12.8, 13.7, 14.1, 14.2, 14.2, 14.1, 14.5, 14, 13.1, 12.6, 11, 9.5, 
    7.5, 6.6, 6.3, 6.7, 6.5, 6.8, 6.7, 6.4, 7.2, 6.3, 5.8, 6.8, 6.1, 6.1, 
    6.3, 6.8, 7.2, 7.4, 6.5, 6.1, 4.5, 3, 1.4, 2.6, 4.5, 6.4, 9.6, 9.9, 9.4, 
    6.9, 6.8, 7.3, 6.8, 6.6, 6.6, 7.3, 7.4, 7.2, 6.2, 6.2, 5.6, 2.6, 2.4, 
    5.6, 6.7, 7.1, 7.6, 8.7, 9, 9.4, 8.9, 9, 9.1, 9.7, 10.2, 9.8, 9.5, 9.3, 
    9.1, 9.4, 9, 9.3, 8.6, 8.1, 7.5, 7.1, 6.4, 5.4, 4.8, 4, 2.8, 2.7, 2.8, 
    3.4, 4.7, 4.8, 4.5, 4.4, 4.2, 4.5, 0.3, 1.7, 3.1, 4.6, 4.4, 4.4, 4.1, 
    3.9, 4.2, 4.4, 4.9, 5.3, 5.7, 6.7, 7.1, 7.2, 7.5, 8.2, 8.6, 8.8, 9.2, 
    9.7, 9.7, 10, 10.6, 10.8, 10.6, 10.8, 10.6, 10.4, 9, 9.1, 9.2, 8.8, 8.3, 
    8, 8.1, 8, 7.7, 7.7, 8, 8, 7.1, 7, 6.6, 6.8, 7, 7, 7.8, 7.7, 7.4, 7.4, 
    7.4, 7.1, 7.3, 7.3, 6.9, 6.9, 6.8, 6.8, 6.9, 7.1, 7.3, 7.4, 7.8, 8.2, 
    6.9, 6.7, 6.7, 6.8, 6.6, 6.1, 5.5, 5, 4.2, 4.1, 3.3, 3.3, 2.3, 2, 1.4, 
    0.9, 0.4, 0.3, 0.8, 0.5, 0.4, 1.2, 2.1, 3.1, 3.1, 4, 4.4, 5.3, 5.3, 5.4, 
    5.6, 6, 6.8, 7.8, 8.1, 8, 7.8, 8.1, 8.4, 8.1, 8.3, 9.2, 8.6, 9.6, 10.5, 
    11.1, 11.3, 11.4, 10.9, 11, 10.9, 10.8, 10.6, 10.3, 9.8, 9.3, 8.7, 7.9, 
    6.7, 5.5, 3.2, 1.2, 1.8, 3.7, 4.1, 4.4, 6.6, 6.4, 6, 5.4, 4.1, 2.7, 3.2, 
    3.7, 3.5, 3.7, 3.8, 3.8, 3.6, 3, 3.4, 5.3, 7.7, 8.4, 6.6, 6.4, 6.2, 6.2, 
    6.6, 6.6, 5.5, 5.4, 4.8, 4.4, 3.6, 3.1, 2.7, 3.6, 4.3, 5.1, 5.8, 6.1, 
    6.6, 6.3, 6.4, 6.4, 7, 7.5, 7.3, 6.6, 6.3, 7.7, 8.5, 7.7, 9.1, 9.2, 9.5, 
    9.6, 9.4, 8.7, 8.4, 8.1, 7.7, 7.4, 7.5, 7.5, 8.2, 8.1, 7.9, 7.8, 8.1, 
    7.6, 8.1, 7.6, 6.8, 6.9, 7.3, 7.2, 6.2, 6.2, 6.2, 6.6, 6.7, 7, 6.9, 6.9, 
    7.1, 7, 7.3, 7.3, 7.1, 7.1, 7.3, 7.4, 7.3, 6.9, 7.1, 7.3, 7.2, 7.4, 7.6, 
    7.5, 7.7, 7.8, 8, 8.1, 8.8, 8.9, 8.7, 8.8, 9, 8.8, 8.7, 9.2, 8.7, 8.6, 
    8.3, 8.8, 8.9, 8.3, 8.2, 8.1, 8, 8.1, 8.3, 8.4, 8.5, 8.4, 8.5, 8.5, 8.1, 
    7.7, 2.8, 2.4, 2.2, 2, 1.9, 3.2, 3.1, 3.1, 2.9, 3, 2.9, 2.5, 2.3, 2.9, 
    3.2, 3.2, 1, 3.6, 3, 2.8, 2.8, 1.3, 6, 1, 2.1, 6.9, 8.9, 8.7, 8.7, 6.9, 
    8.8, 8.5, 8, 7.4, 7.1, 7.4, 6.5, 5.7, 5.9, 6.2, 6, 5.5, 5, 3.9, 3.5, 2.9, 
    2.7, 2.5, 2.3, 2, 1.8, 2, 2.2, 2.4, 2.4, 2.2, 1.9, 1.7, 1.7, 1.6, 1.5, 
    1.4, 1.1, 1.7, 2.4, 2.1, 2, 1.6, 2.1, 2.8, 2.5, 2, 2, 2.1, 1.9, 2, 1.8, 
    1.7, 1.5, 1.8, 1.7, 1.1, 0.4, 0.4, 0.2, 0.4, 0.3, 0.5, 0.5, 0.3, 0.4, 
    0.6, 1.1, 1.3, 2.5, 2.7, 2.9, 3.6, 3.7, 4.5, 5.2, 4.8, 4.2, 3.5, 3.1, 
    2.7, 3, 1.8, 1.2, 0.8, 0.7, 0.6, 0.7, 0.4, 1.8, 2.1, 2.6, 2.9, 2.9, 2.3, 
    1.9, 2.6, 2.4, 2.5, 4.6, 4.6, 5.1, 4.9, 4.9, 5, 5, 5, 5.3, 5, 5, 4.8, 
    4.9, 5.4, 5.4, 5.3, 5.1, 5.3, 5.4, 5.2, 5.2, 4.8, 5.7, 5.5, 2.2, 1.6, 2, 
    4.2, 0.7, 0.8, 1.1, 1.4, 1.2, 1.4, 1.6, 1.4, 1.4, 1.6, 1.5, 1.5, 1.4, 
    1.2, 1.2, 1.4, 1.4, 1.5, 1.6, 1.3, 1.2, 1.3, 1.2, 1.4, 1.6, 2.2, 2.8, 
    3.1, 3.4, 3.4, 3.6, 3.8, 3.7, 3.8, 4, 4.1, 4.3, 4.3, 4.1, 4, 4.3, 4.2, 
    4.7, 4.3, 4.6, 4.9, 5.5, 6, 5.7, 6.6, 6.6, 6.1, 6.4, 6.6, 6.9, 7.2, 7.7, 
    8.2, 8.7, 9, 9.3, 9, 8.6, 8.5, 8.8, 9, 9.2, 10, 10.2, 10.8, 11.3, 11.6, 
    11.6, 11.7, 12, 12.2, 12.2, 12.7, 13.7, 14.3, 14.9, 15.6, 15.5, 15.3, 
    14.3, 14.2, 13.7, 13.2, 13.4, 13.7, 13.3, 13.5, 14, 13.8, 13.9, 13.5, 12, 
    11, 9.9, 10, 9.6, 9.5, 9, 8.6, 8.4, 8.4, 8.5, 8, 7.1, 6.6, 4.8, 3.2, 4.2, 
    5.1, 4.3, 4.2, 3.5, 3.7, 3.3, 3.2, 3.7, 3.7, 3.5, 3.3, 3.4, 3.7, 4.2, 
    4.2, 4.8, 4.7, 4.8, 5.5, 4.6, 4.7, 5.5, 5.5, 5.8, 5.8, 5.2, 5.1, 5.2, 
    5.6, 6.4, 7.5, 8.8, 9.1, 9.4, 9.2, 8.3, 7.7, 4, 5, 6.1, 5.9, 6.6, 7.3, 
    4.8, 6.5, 7.5, 8, 8.2, 8.7, 7.7, 7.9, 8, 8.5, 8.9, 9, 9.4, 9.7, 9.8, 
    10.4, 10.8, 11.2, 11, 11.4, 11.4, 11.9, 12.3, 12.4, 11.8, 12.1, 12.5, 
    12.6, 12.6, 12.7, 12.5, 12.2, 12.1, 12.2, 11.9, 11.5, 11.4, 11.2, 11.3, 
    11.2, 11.2, 11.1, 10.2, 10, 9.7, 9.8, 9.7, 9.5, 9.4, 9.1, 9.1, 8.9, 8.5, 
    8.6, 9.2, 9.5, 9.4, 9.3, 9.1, 9.1, 9.1, 8.9, 9, 9.4, 9.5, 9.1, 8.7, 8.5, 
    7.9, 7.9, 8.1, 7.8, 7.2, 6.8, 6.7, 6, 5.5, 5.1, 5.8, 5.9, 5.6, 4.9, 4.4, 
    3.9, 3.8, 4, 3.6, 3.2, 2.9, 3.3, 3.7, 1, 5.5, 6.6, 6.4, 6.6, 6.6, 6.6, 
    6.6, 6.2, 6.4, 6.6, 6.7, 7.8, 8.5, 8.1, 8.2, 8.4, 7.8, 7.2, 7, 7.6, 7.6, 
    7, 7.1, 6.8, 6.8, 5.8, 5.5, 5.2, 4.7, 5.1, 5.5, 6.1, 6.8, 6.9, 5, 4.7, 
    4.4, 4.9, 5.3, 6.1, 6.7, 6.7, 7.1, 7.5, 8.4, 9.5, 10.5, 10.9, 11.4, 12.6, 
    13, 12.9, 12.8, 12.8, 13.7, 12.5, 12.6, 12.3, 12.1, 11.9, 11.7, 11.6, 12, 
    11, 11, 12.2, 11.5, 11, 10.8, 11.3, 10.7, 10.2, 9.5, 9.2, 9.4, 10.9, 
    10.4, 10.2, 9.4, 9.6, 10, 9.5, 8.9, 9.3, 9.7, 9.8, 9.8, 9.1, 9.5, 11.1, 
    11, 10.8, 10.1, 9.1, 9.3, 9, 8.9, 8.8, 8.7, 7.7, 7.4, 7.2, 6.9, 6.8, 6.7, 
    6.9, 7.1, 6.6, 6.3, 5.7, 5.7, 5.8, 5.5, 5.4, 5.1, 5.4, 5.5, 4.7, 5, 5, 
    5.1, 5, 5, 4.4, 4, 4.3, 4.4, 4.5, 4.7, 4.5, 4.6, 4.8, 5, 4.9, 5.5, 5.2, 
    6.6, 5.9, 6, 5.4, 5.1, 5.4, 5.8, 6.1, 6.6, 6.3, 6.4, 5.7, 5.5, 5.3, 5, 
    4.8, 4.3, 4.9, 4.9, 4.8, 5, 4.8, 4.8, 4.4, 3.8, 4.2, 4.4, 4.3, 4.2, 4, 
    4.4, 4.4, 4.4, 4.4, 4.3, 4.4, 4.1, 4, 4.2, 4.2, 3.9, 4.2, 4.1, 4.2, 3.9, 
    3.7, 3.6, 3.3, 3.4, 3.3, 3.1, 3.3, 3.1, 3.1, 2.9, 3.3, 3, 3.2, 2.9, 2.2, 
    2.3, 2.1, 1.7, 1.4, 1.6, 1.3, 1.2, 1.3, 1.6, 1.5, 1.3, 1.7, 1.9, 2.1, 
    2.1, 2.3, 2.6, 2.4, 2.9, 3.4, 3.9, 3.6, 3.9, 4, 4, 3.9, 3.8, 3.5, 3.2, 
    2.7, 3, 3.4, 3.4, 3.4, 3.7, 4.2, 4, 4.5, 4.8, 4.9, 4.7, 5.7, 5.5, 5, 5.2, 
    5.1, 5, 5.4, 5.8, 0.2, 0.4, 0.8, 1.8, 2.5, 2.3, 2.5, 2.8, 3.8, 3.1, 3.6, 
    4.2, 4.9, 5.1, 4.7, 4.7, 4.9, 5.2, 6.6, 6.3, 6.3, 5.7, 5, 4.8, 5, 5.3, 6, 
    6.6, 7.6, 7.7, 8.2, 8.6, 9.8, 11, 12.4, 13.1, 13.9, 14.8, 15.3, 15.3, 
    14.9, 14.9, 14.6, 14.3, 13.8, 13.1, 13.7, 13.6, 14.8, 14.8, 15.1, 15.6, 
    15.8, 16.1, 16.7, 16.9, 16.6, 15.7, 13.7, 13, 11.9, 11.2, 10.1, 9.6, 8.4, 
    7.3, 5.6, 5.8, 5.4, 5, 4.5, 4.8, 3.9, 3.4, 3.1, 2.3, 1.9, 2.3, 1.5, 1.5, 
    2, 1.9, 3, 3.3, 3.3, 4, 5.2, 5.3, 5.7, 6.5, 6.7, 7.3, 7.4, 7.6, 7.2, 7, 
    5.9, 5.6, 5.6, 5, 3.9, 3.5, 2.7, 3.1, 4.2, 4.1, 3.2, 2.4, 1.9, 1.8, 1.5, 
    1.1, 0.5, 0.9, 1.6, 2.2, 2.7, 2.9, 3.1, 3.4, 2.7, 2.6, 2.7, 2.6, 2.4, 
    2.5, 2.7, 3.1, 2.5, 2.1, 1.5, 1.4, 4.6, 4.2, 3.7, 3.7, 3.6, 3.7, 3.8, 
    3.7, 3.8, 3.1, 2.7, 2.7, 3.7, 3.4, 3.1, 2.8, 3.1, 2.9, 3.7, 3.3, 1.9, 
    1.9, 2.6, 2.9, 3.4, 3.2, 2.9, 3.7, 3.7, 3.8, 3.2, 3.5, 3.9, 3.7, 3.9, 
    3.9, 3.6, 3.4, 3.1, 2.8, 2.7, 2.7, 3.4, 3.4, 3.3, 3.1, 2.6, 2, 1.8, 1.7, 
    1.7, 1.7, 1.8, 2, 1.8, 1.6, 1.2, 0.8, 0.6, 0.4, 2.3, 2.5, 2.8, 2.9, 3, 
    2.9, 3.2, 3.5, 3.5, 3.4, 3.4, 3.5, 4.1, 3.6, 3.3, 3.4, 2.8, 2.4, 2.2, 
    2.3, 2.7, 4.2, 4.7, 5, 5, 4.8, 5, 5.4, 5.2, 4.9, 4.9, 4.5, 4.1, 3.9, 3.5, 
    2.9, 2.5, 2.9, 2.9, 2.8, 2.7, 3.1, 2.9, 2.9, 2.5, 2, 1.8, 1.6, 1.6, 1.7, 
    1.8, 2.3, 2.7, 2.8, 3.2, 3.5, 4.1, 4.5, 5.1, 5.6, 5, 6, 6.2, 6.3, 6.5, 
    6.8, 6.4, 6.6, 6.4, 6.4, 6.4, 6.4, 6.4, 6.4, 6.5, 6.6, 6.5, 6.4, 6.1, 
    5.9, 5.4, 4.7, 4.5, 4.6, 5, 5.3, 5.5, 5.4, 5.5, 5.7, 5.2, 5.5, 5.7, 5.6, 
    5.7, 5.2, 4.8, 4.1, 3.2, 2.6, 1.9, 1.7, 0.7, 0.4, 1.2, 2.7, 3.6, 4.3, 
    3.6, 4.1, 4.3, 4.3, 4.7, 4.6, 5.3, 6, 6.9, 7.3, 7.5, 7.7, 8, 7.9, 8.5, 
    9.1, 9.5, 10.1, 9.5, 9.6, 8.5, 8.2, 8.6, 8.9, 9.1, 9.7, 9.7, 9.4, 9.4, 
    9.2, 8.8, 9.3, 9.5, 10.2, 9.8, 9.5, 9.1, 9.1, 9.5, 9.5, 9.5, 9.6, 9.1, 
    9.5, 9.8, 10.2, 10.8, 10.8, 10.7, 10.4, 11.2, 10.7, 9.9, 9.9, 8.3, 10.2, 
    10.4, 8.8, 7.5, 7.5, 8.1, 8.5, 8.3, 6.9, 6.3, 5.9, 7.1, 5.9, 4.6, 3.9, 
    4.5, 4.4, 5.9, 6.9, 7.5, 7.9, 8.2, 9.2, 7.7, 9.1, 10.3, 11.3, 11.6, 11.7, 
    11.4, 12.2, 12.8, 12.6, 12.1, 12.6, 12.5, 12.4, 11.7, 11.1, 11.9, 12.7, 
    13, 13, 12.8, 12.5, 12.3, 12.6, 12.7, 12.3, 12, 11.4, 11.2, 11.4, 11.8, 
    11.6, 11.7, 11.5, 11.2, 9.9, 8.8, 8.9, 9.5, 9.3, 10.7, 13.2, 13.3, 12.8, 
    12.3, 12.3, 12, 12, 12.4, 11.5, 11.3, 11, 11.5, 11.5, 11.9, 12, 12.4, 
    12.1, 11.9, 11.3, 11.5, 10.3, 9, 8.6, 8, 6.6, 4.4, 5.3, 6.1, 6.1, 6.8, 
    7.1, 8.1, 9.3, 10.4, 11.7, 12.6, 13.3, 13.4, 12.9, 12.8, 12.1, 11.4, 
    11.5, 11.2, 10.7, 10.5, 11.3, 11.5, 11, 10.7, 9.7, 8.6, 7.1, 5.9, 4.5, 
    2.2, 1.3, 1.8, 3.1, 4.2, 5.1, 5.3, 6.3, 7.8, 8.9, 9.7, 10.1, 11.9, 12.1, 
    10.9, 9.1, 8.1, 9.7, 11.3, 12.4, 12.1, 10.9, 10.3, 10.4, 10.6, 10.1, 9.2, 
    8.9, 10.5, 11.3, 11.5, 10, 9, 10.2, 15.1, 15, 15.8, 15.3, 15.4, 15.3, 
    15.2, 15, 13.7, 12.2, 10.3, 7.5, 6.5, 8.2, 9.9, 10.4, 10, 10.2, 11.2, 
    11.2, 12.4, 12.6, 12.4, 12.9, 13.6, 12.5, 12.3, 12, 11.5, 10.7, 10.2, 
    10.8, 9.7, 8.5, 7.2, 5.9, 4.6, 4.9, 4.1, 2.7, 1.6, 2, 3.2, 4.1, 5.6, 6.8, 
    7.8, 7.5, 6.2, 7.3, 6, 5.1, 4.4, 5.2, 6.6, 8.2, 8.2, 8.8, 9.6, 10.2, 
    10.6, 9.7, 9.5, 9.2, 8.6, 8.2, 8.1, 8.8, 9, 9.2, 9, 9.2, 9.4, 8.4, 8.8, 
    8.8, 8.6, 8.5, 8.1, 8.7, 8.5, 8.6, 8.9, 8.6, 8.6, 8.9, 8.6, 8.9, 9, 8.5, 
    8.9, 9.1, 8.8, 8.8, 8.9, 9.4, 9.7, 8.5, 7.9, 8, 8.9, 9.4, 9.7, 10.2, 9.8, 
    9.3, 9.8, 9.7, 9.4, 8.9, 8, 7.9, 8.8, 9.8, 8.7, 8.5, 9.4, 10, 10.2, 10, 
    10.4, 10, 10, 9.5, 9.5, 9.6, 9.7, 11.3, 10.7, 9, 9.3, 10.4, 11.2, 10, 
    9.3, 8.2, 8.4, 8.9, 11, 11.4, 11.5, 11.6, 11.3, 11.1, 9.8, 9.7, 9.7, 9.7, 
    9.6, 9.5, 9.1, 8.9, 8.7, 8.4, 8.4, 8.2, 7.5, 7, 6.6, 6, 5.5, 5.1, 4.8, 
    4.4, 4.4, 4.3, 4.2, 4.1, 4.3, 4, 3.8, 3.9, 4.1, 4.2, 4.2, 4.9, 5.3, 5.4, 
    5.6, 5.9, 6.2, 6.5, 6.7, 6.9, 6.9, 6.9, 7.3, 7.7, 7.8, 7.8, 7.5, 7.1, 
    7.4, 6.7, 6.2, 5.6, 5.3, 5, 5.4, 5.5, 5.3, 4.8, 3.8, 2.7, 3, 4, 4.5, 4.7, 
    4.9, 4.7, 3.8, 3.6, 3.9, 4.5, 4.3, 4.6, 4.2, 4, 3.6, 3.3, 3.2, 2.6, 4.3, 
    4, 3.9, 3.9, 4.1, 4, 5.1, 5.3, 5.4, 4.9, 4.5, 4.3, 4.6, 5.1, 5.7, 6.1, 
    6.3, 6.3, 6.4, 6.6, 6.1, 5.7, 5.2, 5.1, 5.9, 6.1, 6, 6, 5.7, 5.4, 5.8, 
    6.4, 7, 7.1, 7.4, 6.7, 4.6, 5.9, 7.1, 8.3, 9.6, 11.3, 12.3, 12.9, 13.3, 
    13.5, 13.5, 14.1, 12.8, 11.3, 10.4, 8.5, 6, 6.5, 6.8, 7.2, 8.6, 8.2, 7.9, 
    7.4, 8.4, 8.5, 8.1, 6.9, 5, 3.5, 3, 5.1, 10.6, 12.2, 11.3, 9.9, 9.1, 7.6, 
    5.4, 3.9, 3.8, 3.9, 2.4, 2.6, 4, 4.9, 4.8, 4.5, 5.3, 5.3, 5.6, 5.8, 5, 
    4.3, 3.9, 4.2, 4.5, 4.3, 4.6, 3.7, 2.9, 2.8, 3.3, 3.4, 3, 2.9, 3.9, 4.4, 
    4.7, 5.4, 6.1, 7.3, 7, 7.9, 8.6, 9.7, 9.8, 8.7, 8.1, 8.5, 8.8, 9.1, 9.1, 
    9, 8.7, 8.7, 9, 9, 9.4, 9.2, 8.8, 8.5, 8.8, 8.2, 8.6, 8.6, 8.3, 8.3, 8.2, 
    8, 7.6, 7.8, 7.4, 7, 7.1, 7.5, 7.6, 8, 6.7, 6.7, 6.8, 7.1, 7.5, 7.5, 5.9, 
    5.6, 5.4, 4.6, 4.6, 4.8, 4.7, 4.8, 5.4, 5.6, 6.3, 6, 6, 6.4, 7.1, 7.3, 
    8.4, 8.5, 8.3, 8.7, 8.6, 8.9, 9.4, 9.5, 8.3, 8.2, 8.6, 8.9, 8.7, 8.4, 
    8.6, 8.3, 7.6, 6.6, 5.5, 4.4, 4.2, 3.4, 2.8, 3.1, 2.9, 2.4, 3.8, 3.5, 3, 
    2.5, 1.3, 0.2, 1.9, 3.2, 3.9, 4.1, 5, 5, 4.4, 4.4, 4.6, 4.7, 4.7, 4.5, 
    3.8, 4.2, 6.3, 7.6, 7.8, 7.4, 6.9, 6, 4.9, 3.6, 4.1, 4.7, 6.1, 5.3, 4.7, 
    4.2, 3.9, 3.7, 4.2, 3.2, 2.3, 1.6, 1, 2.2, 3.9, 5.3, 6.9, 6.2, 5.7, 5.3, 
    5.4, 5.3, 4.6, 4.5, 4, 3.9, 3.3, 3.5, 4, 3.6, 3.3, 3.4, 3.9, 4.2, 4.3, 
    4.6, 4.5, 4.7, 4.2, 4, 3.5, 3.9, 4.2, 4.4, 2.6, 2.7, 2.9, 3.4, 3.6, 4.3, 
    4.3, 5, 5, 5.2, 5.4, 5.7, 6, 5.8, 5.7, 6, 6.3, 6.4, 6.9, 7.7, 8.2, 8.8, 
    9.2, 9, 7.6, 7.1, 6.8, 6.3, 6.6, 6.4, 5.6, 5.6, 5.7, 6.1, 6.5, 6.8, 8.1, 
    8.4, 8.6, 9, 8.7, 7.8, 11.6, 12.2, 12.2, 11.9, 12.1, 12.1, 11.7, 11.8, 
    12, 12.2, 12, 11.7, 10.8, 10.7, 10.7, 10.6, 10.4, 10.3, 10.2, 9.9, 9.7, 
    9.5, 8.8, 8.1, 8.3, 7.9, 7.4, 6.8, 6.1, 5.3, 4.5, 4.2, 3.7, 2.5, 1.5, 
    1.2, 2.8, 2.4, 2.2, 2.2, 1.8, 1.3, 3.4, 3.6, 3.7, 4.4, 4.7, 4.7, 4.4, 5, 
    5.7, 5.9, 6, 6.3, 7.5, 8.2, 8.8, 9.2, 9.2, 9.3, 9.3, 9.9, 10.2, 10.4, 
    10.8, 11.6, 11.4, 11.7, 11.9, 12.2, 12.7, 13.3, 12.8, 12.9, 13.1, 13.4, 
    13.6, 13.5, 13.2, 13.2, 13.3, 13.3, 13.4, 13.3, 14.5, 14.6, 14.8, 14.7, 
    14.6, 14.4, 13.3, 12.5, 11.6, 10.3, 9.1, 7.5, 4, 2.7, 3.4, 3.7, 3.4, 3, 
    4, 2.7, 2.1, 2.2, 2.2, 2.4, 10.5, 11.8, 11.7, 11.9, 11.8, 11.4, 10.8, 
    10.5, 10.7, 11, 11, 10.2, 9.4, 9.2, 9.5, 9.9, 10.3, 10.6, 10.4, 11, 11.5, 
    11.9, 12.1, 12.6, 13.7, 14.1, 14.3, 14.6, 14.9, 15.2, 15.3, 15.7, 15.5, 
    15.2, 14.5, 13.5, 12.2, 12, 11.5, 10.6, 11, 9.4, 10.4, 9.2, 7.9, 7.7, 
    6.5, 5, 5, 4.4, 4, 3.8, 4.8, 4.9, 4.3, 5.8, 6.7, 7.6, 7.8, 7.4, 6.8, 6.8, 
    6.4, 6.2, 6.9, 6.7, 6.6, 4.7, 6.4, 6.8, 7.4, 7.2, 8.8, 8.4, 7.6, 7.2, 
    7.4, 7.2, 5.7, 6, 6.5, 7.5, 8.3, 8.3, 8.7, 9.4, 8.4, 8.9, 8, 7, 7.2, 4.4, 
    6, 7, 7, 7, 7.4, 8.7, 5.4, 5.3, 7, 7.9, 7, 7.3, 7, 5.7, 7.8, 8.4, 6.1, 
    5.6, 6.5, 8.6, 5.7, 4.6, 3.3, 4.5, 4.6, 3.9, 5.4, 5.2, 4.1, 5.7, 4.4, 5, 
    3.6, 3.5, 2.6, 2.5, 3.6, 3.5, 2.1, 3.7, 2.5, 1.2, 6.3, 6, 7, 5.6, 9, 9, 
    10.5, 9.8, 10.8, 10.1, 8.7, 10.4, 9.6, 7.9, 8.7, 6.9, 7, 11, 10, 11.6, 
    12.4, 15.1, 15.2, 17.1, 16.6, 16.2, 14.3, 13.9, 14.7, 14.1, 14.9, 14.4, 
    14.6, 16, 16.9, 16.2, 16.5, 17.1, 16.5, 17.4, 18.7, 19.2, 19.7, 17.7, 
    19.5, 19.2, 13.3, 17.3, 15.9, 15.5, 13.3, 16, 15.3, 17.8, 17.5, 15.2, 
    16.8, 15.9, 14.6, 14.1, 14.2, 14.1, 13.5, 14, 13, 13.9, 14.1, 11.5, 13.1, 
    14.3, 14.1, 16, 15.4, 16.5, 17.9, 16.6, 18, 17.8, 18, 18.1, 18.2, 17.5, 
    16.1, 15.6, 18.3, 8.9, 15.7, 14.4, 13.3, 14.2, 13.4, 13.7, 10.3, 11.1, 
    7.8, 3.4, 4.6, 5.7, 4.1, 3.5, 2, 1.9, 2, 2.1, 2.2, 1.9, 2, 1.7, 8.2, 8.5, 
    5.6, 6.6, 6.9, 5.4, 6.4, 6.4, 6, 4.8, 5.4, 5.3, 5.1, 5.7, 5, 3.7, 4.2, 
    3.9, 1.5, 0.6, 1.9, 1.8, 1.9, 1.3, 0.9, 0.9, 1.2, 0.5, 0, 0.1, 1.7, 2.1, 
    2.8, 1, 7.2, 4.4, 9, 8.3, 6.9, 9, 9.6, 9.3, 9.3, 9.1, 9.6, 9.2, 9.2, 
    11.1, 10.5, 10.4, 10.9, 10.6, 11.9, 12.7, 12.7, 13.6, 12.3, 12.2, 10.8, 
    11.1, 10.4, 10.9, 10.8, 9.9, 9.2, 7.6, 9.5, 7.2, 8.9, 6.3, 5.6, 6.2, 5.1, 
    6.4, 8.2, 7.1, 6, 5, 4.3, 5.1, 4.9, 4.4, 2.5, 2.5, 2, 5.2, 3.3, 3.6, 3.9, 
    3.3, 6.2, 8.9, 10.2, 10.3, 7.7, 13.3, 15, 15.5, 17.1, 15.3, 16.2, 17.1, 
    16.2, 15.1, 17.5, 18.3, 15.3, 13.2, 10.8, 14.1, 13.1, 13.2, 11.3, 12.5, 
    10.2, 11.3, 9.6, 11.4, 9, 10.6, 9.5, 9.3, 9.6, 10.1, 9, 9, 10.5, 9.9, 
    8.9, 9.6, 9.3, 9.7, 9.2, 9.5, 10.7, 11, 11.3, 5.6, 6.3, 9.3, 12.1, 13.2, 
    12.5, 13.1, 9.7, 3, 5, 4.8, 7.1, 9.1, 8.8, 6.4, 2.3, 2.8, 3.8, 8, 3.4, 
    1.2, 7.1, 4.7, 6.9, 10.5, 6.7, 7.3, 7.3, 12.1, 9.4, 5.9, 4.3, 4.8, 5.7, 
    5.3, 5.4, 6.5, 10.2, 10.9, 13, 14, 14.4, 15.5, 17.8, 18.3, 18.5, 16.6, 
    15.3, 15.3, 16.4, 16.5, 16.9, 15.9, 16.3, 17.1, 15.9, 16.1, 15.5, 14.7, 
    12.9, 11.8, 15.1, 15.7, 16.1, 15.2, 15.7, 15.9, 15, 15.3, 14.4, 14.3, 
    13.9, 14.3, 12.3, 12.2, 14.2, 12.7, 14.7, 14.6, 14.2, 11.3, 14, 7.9, 8.2, 
    8.1, 9.2, 9.7, 10.6, 13, 13, 13.2, 9.6, 2.8, 3.6, 8, 9.6, 8.7, 7.8, 6.7, 
    6.8, 7.4, 8.1, 9.6, 10, 8.9, 9, 8.4, 9.4, 10, 10.8, 11.3, 11.3, 12.2, 
    12.4, 12.1, 11.9, 9.9, 10.1, 9.1, 9.9, 10.8, 11.1, 11.3, 8.9, 5.3, 8.5, 
    4.8, 4.4, 5.8, 3.6, 3.7, 2.5, 3.2, 3.5, 2, 2.4, 3.2, 3.5, 1.8, 3.5, 3.3, 
    3.6, 3.1, 3.2, 5.9, 4, 5, 8.8, 7.4, 9.2, 10.1, 9.4, 10.2, 10.3, 1.7, 8.5, 
    10.2, 9.6, 11.5, 11.3, 11, 8.8, 12.2, 10.9, 1.8, 1.8, 9.7, 10.4, 9.5, 
    4.6, 1.9, 7.3, 7.8, 8.4, 8.8, 10.1, 10.4, 9.3, 10.5, 5, 8.2, 9.4, 6.4, 
    9.7, 9.4, 9.1, 3, 8.7, 8.4, 7.7, 8.8, 8.4, 7.4, 7.7, 7.4, 6.9, 6.3, 5.8, 
    5.9, 7.5, 7.8, 7.5, 6.5, 4.9, 5, 5.1, 4.6, 3.9, 2.8, 5.9, 3.6, 5.4, 4.2, 
    6.2, 8.5, 7.9, 8.5, 7.7, 9.3, 10, 10.5, 10.8, 10.6, 10.8, 10.1, 10, 9.8, 
    9.5, 9.8, 10.2, 10.8, 11.6, 11.5, 12.1, 12, 11.7, 12, 11.7, 13.6, 13.5, 
    14.7, 13.7, 14.6, 14.6, 14.6, 14.8, 15.7, 16, 14.6, 15.5, 14.5, 14, 13, 
    11.9, 13.7, 12, 12, 12.9, 4.4, 11.8, 11.6, 11, 10.7, 11.6, 12.2, 13.2, 
    13.8, 13.3, 14, 11.9, 12.8, 13.3, 13, 13.4, 12.8, 9.7, 9.6, 8.1, 10, 6.4, 
    5.2, 6.9, 1.1, 2.9, 3.8, 5.2, 8.6, 12.8, 10.2, 8.4, 13.1, 11.9, 9.5, 
    11.1, 12.9, 11.1, 10.9, 12.7, 14.5, 13.3, 12.4, 12.5, 11.9, 13.3, 12.7, 
    15, 13.9, 16.8, 19.3, 14.1, 13.2, 17.4, 15, 15.7, 18.1, 16.9, 14.4, 19, 
    19, 16, 14.4, 14.1, 14.1, 14.6, 15.2, 15.2, 15.3, 14.2, 14.2, 14.3, 16.2, 
    16.2, 16, 15.4, 16.1, 19.7, 17.2, 19.2, 19.5, 18.1, 16.2, 16.3, 14.3, 
    15.8, 14.5, 14.7, 14.8, 14.3, 12.5, 14.6, 10.9, 12.2, 11.4, 7.2, 9.6, 
    8.7, 7, 4.5, 7.1, 2.8, 2.1, 2.1, 8.6, 10.9, 8.3, 9, 8.1, 9.1, 7.9, 7.8, 
    6.4, 7.7, 7.9, 7.5, 5.4, 5.3, 7, 6.7, 7.6, 8.1, 10.8, 8.2, 6.8, 6.4, 6.1, 
    5.9, 6.1, 6.6, 3.9, 2, 0.9, 1.9, 1.4, 1.2, 0.9, 1.9, 4.8, 6.4, 4, 3.1, 
    2.8, 0.7, 0, 0.5, 3.5, 1.6, 7.6, 10.1, 9.7, 9.4, 9.1, 8.7, 9.9, 9.3, 
    10.6, 11.3, 9.4, 10.6, 11, 12.6, 12.8, 8.6, 13, 13.7, 12.6, 15.7, 14.6, 
    15.1, 15.6, 14.3, 14.9, 16.3, 14.8, 11.6, 15.2, 13.4, 13.8, 12.6, 11.6, 
    9.8, 12.6, 10.8, 9.9, 11.3, 10, 8.6, 9.8, 9.1, 8.6, 7.5, 7, 5.4, 7.8, 
    5.5, 5.2, 8.2, 7.4, 8.2, 7.5, 5.4, 5.2, 5.6, 5, 5.1, 7.1, 7.3, 6.2, 1.9, 
    2.8, 0.7, 1.7, 3.1, 3.5, 2.9, 3.3, 3.4, 5.1, 4.8, 4.8, 5.1, 4.6, 5.3, 
    5.4, 1, 6.1, 7.3, 4.5, 7.2, 7, 10.4, 3.8, 1.3, 8.9, 10.1, 9.6, 8.8, 8.2, 
    7, 10, 9.7, 11.5, 10.3, 1.2, 1.9, 1.4, 1.2, 0.8, 1.7, 0.4, 0.9, 1.2, 5, 
    3, 2.9, 7.3, 10.1, 9.7, 3.9, 4.3, 5.4, 4.7, 6.9, 5.8, 7.4, 8.1, 8, 4.8, 
    6.7, 3.7, 7.4, 7, 1.7, 1.1, 7.8, 10.5, 11.9, 9.2, 10, 7.8, 6, 4.7, 4.2, 
    3.8, 5.8, 5.6, 7.4, 5.3, 3.1, 5.1, 3.9, 6.7, 9.6, 10.3, 8.3, 4.6, 7.6, 
    2.6, 6, 2.7, 7.7, 7.3, 8.6, 5, 6.7, 11.3, 9.8, 11.2, 10.4, 9.9, 9.3, 
    11.1, 8.9, 12.7, 10.9, 6.9, 7.7, 1.3, 5.1, 8.8, 7.7, 7.4, 7.4, 1.3, 2.7, 
    3.3, 6.3, 4.2, 6.9, 9.5, 9.3, 8.5, 7.4, 9.5, 9.1, 5.1, 6.1, 5.4, 4.2, 5, 
    5, 6.3, 5.6, 6.4, 5.1, 6.1, 6.5, 6.1, 4.7, 6.2, 6.5, 6.6, 7, 7.9, 8.4, 
    8.1, 6.6, 8.4, 7.9, 9.2, 7.7, 9.3, 7.8, 4.8, 10.2, 5.9, 1.2, 5, 7.4, 1.6, 
    7.3, 6.2, 4, 5.9, 4, 4.2, 6.3, 4.6, 5, 3.8, 4.8, 5.2, 5.9, 7.3, 6.4, 4.7, 
    3.6, 4.9, 4.8, 4.5, 3.2, 4.6, 4.6, 3.7, 4.2, 4.6, 5.9, 5.9, 3.5, 5.7, 
    6.4, 4.8, 3.6, 5.3, 4, 4.7, 3.4, 4, 4.2, 2.6, 2.9, 2.6, 1.7, 1.9, 3.4, 
    3.7, 4.3, 3.9, 6, 4.3, 4.2, 5.6, 5.5, 4.8, 4, 3.8, 5.4, 3.6, 4.4, 6.1, 
    6.1, 7.4, 8.3, 7.9, 8.3, 10.1, 6.7, 5.2, 7.3, 6.4, 4.8, 6.3, 5.6, 6.9, 
    5.3, 4.3, 7.3, 7.4, 8.3, 5.8, 5.7, 5.8, 6.5, 4.2, 2.6, 3.6, 3.1, 3.3, 
    6.6, 5.1, 5, 5.8, 4.2, 4, 3.8, 4.3, 3.8, 1.5, 1.4, 1.2, 2.2, 2.2, 3.8, 5, 
    4.1, 3.5, 4.3, 5, 5, 2.6, 4.1, 4, 2.8, 2.5, 1.3, 3.3, 2.3, 3.4, 5, 4, 
    1.8, 2.7, 5.4, 4.2, 0.1, 1.1, 1.8, 1.7, 1.7, 1.4, 3.1, 2.7, 6.8, 6.7, 
    7.3, 6.5, 9.3, 9.9, 8.5, 6.1, 7.4, 6, 4.3, 7.6, 8, 7.4, 7.6, 8.3, 10, 
    9.8, 10.8, 10.3, 8.2, 8, 9, 10.5, 10.3, 11.1, 11, 11, 9.3, 9.8, 8.5, 9.5, 
    8.2, 10.1, 11.5, 11.7, 12.2, 11.1, 12.1, 10.9, 9.2, 9.7, 9.1, 9.9, 10.1, 
    9.6, 10.5, 12, 11.3, 9.9, 10.9, 11.7, 13.4, 10.2, 12, 10.9, 12.3, 13.1, 
    8.3, 13.2, 12.6, 13.1, 13.1, 11.6, 13.1, 11.8, 11.1, 10.2, 11.6, 11.3, 
    10.4, 10.8, 10.1, 12.2, 13.6, 11.4, 11.4, 10.1, 10.4, 8.7, 8.6, 8.5, 8, 
    9, 7.9, 7.6, 5.2, 6.6, 4.6, 5.6, 5.8, 4.5, 4.4, 4.8, 4.5, 3.4, 3, 2.7, 
    3.1, 2.8, 2.4, 1.6, 3.6, 3.5, 1.7, 2.1, 4.8, 5.1, 2.4, 3.9, 4.2, 4.5, 
    5.3, 5.7, 4.6, 4.5, 5.6, 4.8, 5.9, 4, 4.9, 5.7, 5, 5, 3.3, 4.7, 4.1, 4.1, 
    4.6, 6.3, 6.7, 7.1, 7.6, 7.8, 6.9, 6.2, 6, 5.2, 5.1, 5.6, 6, 7, 7.6, 7.5, 
    7.5, 7.8, 6.7, 6, 5.6, 5.8, 5.5, 6.4, 7, 8, 8.4, 7.6, 7.8, 6.1, 6.8, 6, 
    5.4, 5.3, 4.3, 6.6, 4.9, 4.4, 4.4, 4.5, 5.3, 5, 2.6, 6.3, 7.8, 7.7, 6.8, 
    10.8, 7.8, 9.1, 8.8, 12.4, 11, 8.8, 9.3, 9.4, 10.5, 10.5, 10.5, 8.7, 12, 
    10.8, 14.1, 11.1, 12.3, 19.1, 13.4, 17.6, 13.3, 14.1, 13.9, 15.8, 21.4, 
    19.4, 21, 21.2, 20.1, 20.1, 19.8, 18.2, 18.7, 17.3, 16.8, 14.4, 11.5, 
    9.6, 8.3, 9.3, 10, 8.1, 7.9, 6.5, 8.3, 6.7, 6.2, 5.6, 3.7, 4, 6.2, 5.6, 
    4.6, 2.7, 3.9, 4, 2.4, 2.1, 2.5, 1.8, 0.5, 0.4, 2, 0.9, 0.4, 3.8, 4.1, 
    4.4, 4.5, 8.3, 10.5, 11.6, 11, 8.8, 10.5, 9.3, 9.7, 6.1, 9.7, 9.9, 11.9, 
    11.1, 11.1, 6.2, 12.5, 7, 11.3, 12.2, 14.3, 12.5, 12.5, 11.6, 11.9, 11.5, 
    12.3, 12.8, 11.4, 10.2, 11.3, 8.8, 10.1, 9.1, 7.2, 6.5, 7.9, 3.4, 1.7, 
    1.6, 2.9, 2.6, 2, 1.1, 4.8, 6.8, 6.8, 6.5, 5.8, 3.5, 3.9, 2.1, 0.8, 1.8, 
    3.7, 0.2, 3.1, 2.8, 4.5, 4.4, 8.9, 10.5, 12, 11.5, 12.6, 13.6, 13.9, 
    13.9, 13.5, 13.4, 13.5, 13.9, 15.1, 15.1, 14.7, 15.9, 15.9, 15.9, 14.3, 
    13.7, 14.2, 14, 14.3, 14.8, 16, 16.8, 16.7, 14.9, 14, 15, 15.5, 15.1, 
    15.6, 14.9, 12.2, 11.1, 10.7, 12.9, 11.7, 12, 12.1, 11.7, 12, 11.8, 11.4, 
    12.1, 12.9, 13, 14, 10, 11.4, 10.4, 10.2, 8.9, 6.7, 8.2, 9, 9.4, 8, 9.4, 
    8, 11.2, 10.8, 10.1, 9.5, 8.6, 4, 8.1, 8.7, 8.4, 6.9, 6.5, 5.5, 6.7, 6.8, 
    5.5, 5, 3.9, 1.2, 2.5, 2, 3.7, 0, 2.7, 2.6, 2.3, 3.7, 2.4, 4.2, 2.2, 1.9, 
    1.7, 2.5, 2.1, 4, 3.1, 0.4, 0.2, 0.1, 1.7, 1.5, 1.3, 2, 2.5, 0.7, 2.3, 
    0.3, 0.8, 2.6, 7.4, 6.8, 7.2, 7, 5.5, 7.3, 9.7, 8.9, 6.8, 7.3, 5.9, 5.7, 
    7.4, 8.6, 6.9, 7.7, 7.3, 9.1, 7.4, 7, 7.3, 6.7, 6.5, 5.7, 6.3, 5.9, 5.2, 
    5.5, 5.1, 4.4, 4.1, 3.6, 4.2, 4.7, 4.2, 4, 4, 4.1, 4, 3.3, 2.9, 2.8, 1.9, 
    1.7, 1.5, 1.3, 2.1, 3.5, 4, 4.3, 3.2, 2.2, 3.6, 4.7, 5.1, 6.5, 5.3, 5.1, 
    6.3, 5.6, 5.7, 6.9, 5.6, 5.6, 6.5, 6.1, 6.5, 6.4, 6.8, 6.5, 5.9, 7.3, 
    8.2, 7.8, 7.9, 6.9, 8.4, 7.3, 7.6, 8.1, 8.7, 8.8, 4.1, 7.2, 6.7, 7.3, 
    8.6, 8.5, 8.8, 9.5, 9.1, 8.6, 8.8, 9.8, 9.9, 9.3, 9.8, 9.7, 9.1, 9, 9.1, 
    9.6, 9.3, 8.6, 8.9, 7.9, 7.4, 6.7, 7.4, 5.4, 5.3, 5.5, 6.1, 5.3, 4.2, 
    5.8, 6.2, 6.5, 5.6, 5.9, 5.1, 5.2, 5.1, 5, 4.7, 5.4, 5.9, 6.2, 6.5, 6.5, 
    8.3, 10.3, 9.4, 9.4, 7.4, 6.1, 2.5, 8.7, 3.8, 5.7, 9.3, 6.1, 3.8, 1.9, 
    3.5, 4.5, 5.2, 5.1, 3.9, 3.9, 2.2, 4.2, 9.3, 9.7, 10.1, 9, 8.8, 7.4, 5.4, 
    6.7, 9, 8.4, 8.2, 7, 7.2, 8.5, 9.8, 8.9, 10.4, 7.6, 8.6, 9.4, 8.4, 10.6, 
    10.7, 8.8, 9.1, 7.2, 3.6, 6.6, 8.2, 8.5, 10.7, 12.4, 14.1, 6.4, 7.8, 4, 
    2.5, 3, 8, 7.9, 4.6, 2.3, 2.9, 3.3, 4.7, 1.8, 0.1, 1.3, 0.4, 1.9, 7.3, 
    4.8, 5.6, 0.4, 6.6, 1.1, 1.9, 8, 4.8, 6.7, 6.1, 8.6, 9.2, 7.8, 8, 7.6, 
    8.2, 6.8, 8.3, 6.6, 9.1, 7.9, 6, 5.4, 8, 10.4, 8.8, 8.4, 5.5, 2.2, 6.1, 
    4.6, 5.2, 5.4, 5.4, 3.2, 3.6, 5.6, 3.2, 4.7, 3, 3.2, 5, 3.3, 4.5, 5.2, 
    4.9, 5.3, 4.2, 4.3, 5.5, 3.4, 3.4, 2.7, 3, 1.9, 3.6, 0.8, 0.8, 0.8, 0.9, 
    1.8, 0.2, 1.1, 2, 2, 0.4, 2.4, 2.7, 1.7, 0.3, 0.5, 1.8, 1.7, 2.4, 2.1, 2, 
    1, 1.1, 2.1, 2.7, 1.4, 2.7, 3.8, 4.4, 3.5, 3.8, 4.3, 3.9, 4.1, 4.4, 4.4, 
    3.5, 4.2, 5.5, 3.7, 3.9, 2.9, 3.4, 4, 4.1, 4.3, 1.6, 2.9, 2.6, 3.5, 3.8, 
    3.8, 3.3, 1.9, 1.3, 1.8, 0.8, 0.9, 1.4, 0.2, 1.3, 0.7, 2.9, 4.5, 2.6, 
    1.7, 2.8, 2.6, 3.8, 1, 1.1, 1.7, 3, 4.2, 0.9, 9.8, 12.9, 15, 6.9, 5, 5.1, 
    6.1, 6.9, 5.6, 6.7, 4.8, 4, 3.6, 7, 2.6, 5.4, 6.3, 7.5, 4.7, 6.6, 10.9, 
    4.3, 4.3, 6.1, 7.7, 8.4, 7.9, 7.5, 7.2, 6.6, 6.3, 6.4, 7.4, 8.3, 6.5, 
    6.2, 3.9, 7, 3.3, 4.4, 6.3, 4.4, 6.6, 4.6, 5.4, 4.8, 6.3, 5.6, 5.1, 5.4, 
    4.9, 4.8, 5.8, 5, 6.2, 4.4, 4.5, 3.7, 3.6, 5.8, 4.3, 4.6, 4, 4.4, 3.4, 
    3.4, 3.9, 4.6, 4.5, 4.8, 4.1, 2.2, 3.1, 3.5, 3.3, 3, 3.3, 4.2, 3.8, 2.9, 
    3.1, 2.1, 2.2, 2.3, 4.8, 4, 3.8, 4.1, 3.5, 4.4, 2.6, 3.6, 2.8, 1.1, 0, 
    3.1, 2.8, 4.4, 5.9, 5.9, 6.2, 6, 6.3, 6.3, 5.7, 5.5, 3.9, 1.9, 2.7, 1.3, 
    1.7, 4.1, 4.2, 3.5, 5, 4.4, 4.4, 5.1, 5.4, 3.8, 3.2, 1.1, 0.9, 2.6, 2.5, 
    2.2, 3.2, 2.4, 6.5, 6.9, 8.5, 8.1, 7.1, 7.8, 8.3, 6.7, 6.8, 5.1, 2.5, 
    4.1, 3, 3.3, 3.3, 1.4, 1.5, 1.7, 0.4, 2.4, 0.2, 2.3, 3.6, _, 3, 4.1, 3.4, 
    4.8, 6.4, 7.8, 8.2, 8.1, 8.1, 8.2, 5.8, 9.4, 8.3, 10.1, 8.8, 8.9, 6.8, 
    9.8, 8.5, 9, 7.3, 6.9, 5.8, 5.5, 5.3, 5.8, 5.7, 4.8, 5.7, 6, 7.6, 7.6, 
    8.2, 7.6, 8.9, 11, 8.7, 10.4, 12.1, 9.6, 12.6, 11.4, 12.5, 11.2, 11.1, 
    12.8, 11, 10.7, _, 9.8, 10.7, 10.9, 9.8, 13.9, 11.5, 9.8, 8.5, 5.4, 6.9, 
    4.5, 6, 7.6, _, 12.5, 14.1, 14.5, 16, 16.6, 16.9, 17.1, 15.2, 13.1, 17.3, 
    15.7, 13.1, 14.1, 10.1, 11, 9.2, 9.6, 11.8, 14.4, 13.4, 11.1, 10.8, 13.2, 
    12.5, 12.9, 15.6, 14.3, 13.9, 13.8, 14.8, 15.4, 17.1, 15.2, 15.5, 14.3, 
    15.2, 14.5, 15.1, 15.6, 15.7, 13.7, 14.4, 15.2, 16.1, 17.2, 15.6, 17.3, 
    18.1, 18.9, 18.7, 18.1, 17.1, 14.8, 15, 11.4, _, 8, 10.9, 11.2, 10.5, 14, 
    12, 10.3, 10.7, 11.6, 11.5, 10.4, 11, 7.5, 8.6, 6.3, _, 6.2, 8.8, 6.6, 
    5.8, 6.1, 6.5, 7.1, 7.5, 7.5, 7.2, 8.1, 7.3, 7.5, 7.7, 11.1, 11.2, 11.4, 
    8.7, 8.3, 9.7, 9.7, 8.1, 7.8, 8, 8.1, 6.5, 6.2, 5.5, 5.4, 4.6, 4.8, 4.1, 
    5.5, 4.1, 3.9, 3.8, 2.7, 3, 3.6, 3.3, 3.7, 3.2, 2.8, 4.6, 3.9, 4.6, 4, 
    3.7, 3.6, 3.4, 3.4, 4, 3.4, 4.1, 4.2, 4.4, 4.4, 4.7, 6.4, 5.6, 5.4, 4.9, 
    4.8, 4.2, 6.7, 7.2, 7.4, 9, 7.8, 8, 8.2, 6.2, 5.3, 8.6, 5.7, 6.8, 6.3, 
    7.2, 6.8, 8.6, 7.7, 8.2, 7.6, 8.4, 11.1, 8.6, 6.2, 7.6, 7.7, 7.7, 5.7, 
    5.3, 5.7, 6.6, 8.9, 10.4, 7.8, 9.9, 10.5, 10.6, 12.3, 11.4, 9.8, 10.8, 
    8.9, 8, 9.7, 7.7, 8, 11.1, 11.9, 12.5, 13.3, 12.4, 12.5, 13.7, 14, 12.8, 
    12.1, 12.7, 11.3, 10.2, 7.3, 6.2, 7.2, 6.4, 5.9, 7.9, 7, 5.7, 9.6, 8.5, 
    5.1, 4.7, 5.4, 4.3, 8.6, 7.4, 7.6, 6.2, 6.5, 4.3, 3.7, 9, 6.9, 6.7, 6.9, 
    8.2, 5.2, 6.3, _, 6.8, 6.7, 5, 7.1, 5, 2.5, 2.5, 1.4, 2, 3.9, 2.2, 4.3, 
    5.3, 7.9, 9, 8.1, 6.7, 7.7, 5.4, 6, 5.4, 8.7, 10.5, 6.9, 8.7, 7.4, 9.3, 
    10.1, 9, 9.7, 5.9, 8.6, 9.1, 6.2, 6.2, 6, 7.7, 8.2, 8.3, 6.6, 9.8, 12, 
    8.9, 8.5, 4.3, 10.9, 4.2, 8.5, 7.2, 8.7, 8.1, 9.2, 8.5, 8.5, 8.5, 8.7, 
    6.6, 7.5, 5.1, 5.1, 4.7, 4.9, 7, 6.7, 6.3, 5.5, 7.1, 5.4, 5, 4.2, 5, 5.5, 
    5.2, 6.6, 6, 6, 5.4, 5.4, 4, 4.9, 2.9, 3.3, 4.4, 6.3, 5.4, 5.7, 5.7, 6, 
    4.9, 5.2, 6.5, 6.5, 6.8, 6.3, 5.9, 6.9, 6.7, 7.7, 7.1, 7.3, 7.3, 7.6, 
    7.6, 8.2, 6.2, 7.3, 6.8, 6.2, 6.1, 6, 6.9, 6.5, 7, 8.2, 6.2, 6.2, 6.4, 
    5.1, 4.5, 4.2, 3.4, 3, 1.8, 1.7, 3.6, 4, 4.4, 3.4, 3.4, 2.8, 2.3, 3.2, 
    4.1, 4.9, 4.6, 4.2, _, 2.9, 3.1, 3.6, 3.4, 2.9, 3.4, 3.6, 3.5, 4.4, 2.8, 
    1, 1.5, 3.2, 3.6, 2.7, 6.8, 4.6, 5.1, 1.4, 0.7, 1.2, 1.6, 1.2, 0.5, 1.1, 
    0.5, 1.1, 0.7, 1.4, 2.5, 7.6, 9.1, 11.3, 11.6, 12.5, 12.7, 13, 12.2, 
    10.6, 10.4, 9.9, 11.5, 11.8, 11, 9.8, 7.6, 6, 10.5, 10.8, 2.5, 11.3, 10, 
    9.1, 9.6, 9.3, 7.9, 5.8, 8.8, 10.8, 6.3, 7, 6.9, 1.2, 4.3, 1.6, 3.8, 5.6, 
    3.1, 1, 6.5, 7.2, 7.2, 8.9, 8.3, 7, 5.4, 7.1, 7.9, 8.8, 9.9, 9.7, 9.3, 
    7.7, 7.5, 10.7, 10, 10.6, 11.9, 12.7, _, 9.5, 10.5, 9.6, 9.1, 7.9, 8, 
    4.2, 4, 2.7, 1.5, 1.3, 1.7, 3.2, 3, 2.4, 2.7, 1.9, 1.2, 2.5, 1.1, 1.8, 
    2.9, 2.6, 2.7, 3.3, 3, 2.9, 2.7, 3.8, 5.5, 5.1, 5.2, 4.9, 5.3, 5.9, 6, 
    4.8, 4.1, 5.1, 5.2, 5, 3.8, 4.2, 2.7, 2.4, 1.4, 0, 3, 6.1, 4.6, 6.3, 7.1, 
    6.6, 7, 6.4, 5.5, 5.9, 4.9, 5.2, 3.9, 3.8, 3.6, 2.1, 1.9, 2.3, 1.3, 2.3, 
    2.1, 2.4, 2.8, 3.7, 5, 5.6, 7.4, 9, 10, 9.7, 10.4, 9.8, 8.9, 9.9, 8.2, 
    9.3, 8.9, 9.4, 9.2, 9.1, 10.1, 10.3, 11.4, 10.7, 12, 11.9, 12.4, 13.1, 
    12.5, 12.8, 11.4, 11.1, 11.4, 10.6, 10.4, 10.9, 10.5, 11.2, 10.1, 10, 
    9.2, 9.4, 9, 9.4, 10.2, 9.1, 8.7, 8, 8.1, 8.4, 8.7, 6.6, 4.5, 2.7, 1.4, 
    0.7, 0.8, 2.5, 3.3, 4, 4.3, 1.4, 2.8, 1.5, 0, 1, 5.5, 5, 4.8, 5.1, 3.7, 
    4.2, 4.6, 5.6, 4.9, 6.2, 5.9, 5.5, 5.7, 6.5, 6.5, 6.3, 5.5, 5.1, 3.8, 
    3.6, 3, 0.7, 3, 1.8, 3.3, 3.2, 4, 3.3, 3.2, 3.6, 3.8, 2.6, 2, 1.7, 2.1, 
    3.2, 4, 3.6, 5.4, 6, 5.8, 5.5, 5, 4.6, 4.5, 2.2, 1.9, 0.5, 0.5, 1.7, 2.1, 
    1.2, 1.3, 0.8, 1.6, 0.7, 1.5, 1.4, 1.4, 1.6, 1.6, 0.9, 0.8, 0.4, 2.3, 
    1.9, 1.2, 0.1, 2, 3.8, 3.4, 4.3, 6.5, 7, 5.2, 7.2, 7.6, 7.7, 9.4, 10.2, 
    11.4, 10.3, 8.7, 9.1, 8.5, 8.9, 8.2, 8.4, 6.4, 6.2, 4.1, 4.9, 4.5, 3.3, 
    3.5, 3.1, 2.5, 2.7, 3.3, 3.3, 1.6, 0.8, 0.6, 0.3, 0.4, 1.1, 3.5, 3.3, 
    3.7, 3.1, 2.5, 1.3, 0.7, 1, 0.6, 3.8, 3.1, 3.1, 1.8, 1.8, 1.5, 3.2, 3.3, 
    0.7, 2.1, 1.2, 2.1, 4.4, 7.3, 4.9, 3, 4.7, 4.5, 7.6, 5.1, 5.3, 5.9, 5.3, 
    4, 2.5, 2.2, 2.2, 4.8, 6.3, 4.9, 4, 2.8, 5.7, 5.9, 6.6, 5.7, 4.8, 4.2, 
    4.8, 4.4, 3.3, 2.8, 3.1, 3.5, 3.1, 4.5, 5.1, 5.4, 6.5, 6, 5.1, 4.4, 4.8, 
    4.9, 7, 8.2, 6.5, 6.5, 6.2, 5.5, 9.3, 7.9, 7.2, 6.3, 4.1, 3.8, 4, 4.4, 
    3.6, 1.3, 2.4, 3.5, 3.9, 4.2, 1.4, 3.1, 3.9, 0.9, 5.9, 5.7, 6, 7.4, 5.5, 
    4.9, 7.8, 9.6, 10.4, 9, 6.8, 5.9, 10, 11.3, 12, 12.2, 9.3, 8.7, 7.4, 5.2, 
    7.9, 7.7, 5.4, 4.9, 4.3, 3.9, 3.8, 3.8, 3.7, 4.3, 3.7, 5.4, 5.2, 4.9, 
    3.8, 3.6, 3.7, 3.9, 2.8, 3, 2.9, 2.1, 3.7, 3.2, 4.1, 3.4, 4.2, 4.1, 3.4, 
    3.5, 3, 2.3, 2.3, 2.9, 2.2, 1.9, 1.6, 2.6, 1.9, 3.2, 2.4, 2, 1.3, 2.5, 
    2.2, 1.2, 1.2, 1.5, 0.8, 1.2, 1.3, 0.4, 1.4, 1, 1.8, 1.7, 0.9, 0.4, 0.5, 
    0.6, 5.3, 0, 1.7, 1.4, 0.5, 1.2, 1.3, 1.9, 1.7, 2.5, 2, 1.7, 1.8, 1, 0.7, 
    0.3, 0.1, 0.8, 1.2, 1.4, 1, 2.1, 0.1, 0, 3.6, 1.7, 0.4, 1.5, 0.3, 1.6, 
    1.2, 1.5, 3.3, 4.7, 4, 3.7, 3.6, 3, 3.2, 4.5, 4.5, 4.4, 5, 5.3, 5.3, 6, 
    6, 7.7, 10.1, 9.5, 10.7, 9.7, 8.6, 8.5, 8.3, 8.9, 7.3, 8.4, 6.9, 8.3, 7, 
    7.7, 6.7, 6.4, 6.3, 6.5, 8, 6.4, 6.1, 7.3, 5.5, 6.9, 6.1, 4.5, 4, 2.1, 
    1.7, 0.9, 1.3, 2.7, 2.8, 4.8, 6.1, 6.8, 4.9, 7.2, 7.8, 9.1, 9.6, 10.7, 
    11.4, 11.9, 11.2, 9.8, 10.6, 12.2, 11.5, 12.1, 11.8, 11, 11.4, 11.3, 8.3, 
    7.9, 7, 5.7, 5.9, 6.5, 6, 4.8, 5.7, 6.1, 6.6, 6.3, 7.2, 5.7, 4.8, 4.3, 
    4.1, 4.1, 4.4, 4, 2.8, 3, 4, 1.9, 2.7, 3.9, 4.2, 4.1, 4.5, 5.5, 4.1, 4.3, 
    5.1, 8.4, 7.9, 10.1, 10.2, 11.3, 12.3, 12.8, 13.3, 9.2, 12, 9, 7.5, 8, 
    8.8, 10.2, 10, 9.8, 10.8, 10.8, 12.6, 13.8, 13.8, 11.6, 11.3, 11.7, 13.5, 
    13.1, 14, 13, 10.9, 8.9, 8.6, 8.8, 6.5, 7.2, 6.2, 7.2, 6.6, 8.1, 7.1, 
    7.1, 7.1, 6.6, 5.8, 4.7, 4.9, 4.6, 4.7, 3.9, 3.3, 3.4, 2.8, 3.8, 4, 4.1, 
    3.3, 4.1, 3.5, 3.9, 4.8, 6.5, 7.6, 8, 9.2, 9.8, 7.6, 6, 4.8, 5.5, 7.2, 7, 
    7.4, 8.7, 11.3, 9.6, 9.4, 9.8, 8, 7.2, 7.7, 8.6, 7.5, 6.8, 5.6, 7.4, 7.6, 
    6.8, 7.5, 7.2, 7.3, 6.6, 5.9, 5.1, 2.5, 1.2, 0.5, 0, 0, 3.9, 3.2, 0, 0, 
    2.7, 1.7, 2.1, 0.8, 3.9, 4.6, 4.6, 1.5, 1.9, 0.9, 0.9, 1.4, 2.5, 3.9, 
    4.5, 2.6, 4.4, 5.8, 5, 5.3, 6.8, 7, 5.2, 5.4, 3.8, 3, 3.5, 2.6, 3.5, 3, 
    4.1, 3.5, 2, 2.4, 3.3, 3.1, 1.5, 1.9, 2, 2.3, 2.2, 1.4, 1.4, 2.3, 2, 2, 
    2.4, 1.4, 1.7, 2.9, 3, 4.8, 5.7, 3.1, 2.3, 1.1, 3.8, 2.7, 1.6, 3.8, 5.6, 
    1.7, 4.4, 4.7, 4, 3.3, 2.1, 0.5, 6.9, 6.5, 6.3, 6.8, 6.8, 4.8, 8.1, 6.9, 
    6.7, 6.1, 8.7, 8.8, 9.5, 7.2, 5.2, 6.5, 5.8, 6.3, 7.7, 7.6, 5.5, 5.9, 
    5.2, 5.8, 5.6, 5.1, 6.1, 4.8, 4.1, 4.4, 5.4, 5.6, 4.9, 7.7, 5.5, 3.2, 
    3.3, 3, 3.3, 5.3, 5.8, 4.2, 4.8, 4.4, 4.1, 4.8, 5.4, 5.4, 5, 5.8, 6.4, 
    5.2, 4.4, 4.8, 4.7, 4.8, 4.1, 5.3, 5.1, 6.1, 7.8, 6.6, 7.9, 6.9, 6.8, 
    8.3, 8.2, 9.1, 9.2, 4.9, 4.5, 3.7, 4.6, 4.7, 3.7, 3, 3.2, 5.2, 5.1, 4.4, 
    4.8, 4.5, 3.1, 3.3, 4.2, 5.1, 5.9, 3.4, 4.6, 3.7, 3.9, 4.2, 4.2, 3.8, 
    3.7, 3.6, 3.4, 3.2, 4.4, 5.4, 3.2, 4.4, 2.3, 3.5, 2.1, 1.8, 2.5, 4.4, 
    4.3, 2.5, 2.2, 0.3, 3, 3.3, 4.8, 3.4, 2, 1.5, 1.5, 1.2, 1.1, 2.7, 4.3, 
    3.9, 1.7, 0.7, 0.8, 6.3, 4.3, 3, 12.2, 10.8, 11.5, 12.8, 3.3, 0.2, 7.6, 
    8.4, 7.9, 7.8, 11.5, 14.3, 9, 6.8, 8.6, 2.3, 1.3, 2.2, 2.7, 4.7, 2.5, 1, 
    1.3, 0.6, 0.7, 1.7, 1, 10.6, 9.7, 7.8, 1.9, 13.3, 14.7, 14.2, 11.9, 10.1, 
    9.7, 7, 7.9, 7.3, 10.7, 9.8, 2.7, 6.7, 12.1, 10.1, 13.7, 2.4, 12.2, 5.4, 
    13.9, 11.6, 11.2, 14.2, 13.7, 11.3, 11.6, 10.6, 11.5, 12.9, 10.7, 11, 
    10.5, 10.6, 11.3, 11.9, 10.8, 9.7, 9.6, 9.1, 6.5, 8.3, 8.5, 9.1, 9.2, 
    8.9, 9.2, 8.6, 9.7, 8.3, 10.6, 10.2, 10.1, 9.9, 9.2, 7.9, 7.3, 7.2, 7.5, 
    6.7, 5.6, 5.1, 7.4, 2.3, 1.9, 2.1, 2.2, 0.5, 12.7, 11.9, 12.9, 12.1, 
    11.7, 9.6, 9.7, 10.1, 10, 10.2, 8.4, 6.4, 6.6, 6.8, 5.8, 5.9, 6.1, 8.2, 
    9.5, 8.1, 9.4, 10.1, 10.7, 11.6, 9.6, 11.4, 13.5, 12.4, 12.4, 12.8, 11.4, 
    10, 10.8, 11.8, 11.7, 10.1, 10.6, 10.2, 9.4, 6.5, 3.1, 2.3, 2.8, 1.7, 
    0.4, 3.1, 0.7, 0.9, 0.8, 0.8, 0.2, 1.6, 0.4, 0.6, 1.1, 1.9, 5.9, 1.9, 
    4.9, 5.2, 2.3, 1.2, 1.6, 1.8, 1.5, 0.9, 4, 1.1, 0.9, 1.7, 1.1, 0.5, 0.5, 
    4, 5.3, 4.5, 5.7, 6.5, 6.7, 6.8, 5.9, 6.7, 6.4, 5.3, 4.7, 4.7, 5.2, 5.5, 
    2.7, 4.5, 5.2, 4.4, 3.7, 3.7, 3.7, 2.2, 0.5, 0.8, 1.3, 2.6, 2.5, 4.2, 
    5.4, 4.5, 6.1, 5, 5.2, 5.2, 5.1, 6.5, 8.4, 9.6, 10.3, 10, 9.1, 10.6, 
    11.9, 9.2, 8.7, 8.3, 4.9, 3.6, 3.8, 6.3, 2, 4.2, 8.7, 9.5, 9, 10.9, 9.1, 
    12.4, 9.2, 7.1, 7.6, 13.1, 11.6, 12.9, 12.8, 12.4, 12.1, 12, 14.8, 15.2, 
    13.2, 12.5, 14, 13.5, 14.2, 11.4, 10.4, 10.3, 9.2, 8.3, 5.7, 7.8, 7, 7.6, 
    7.6, 9.5, 10.7, 11.9, 9.8, 9.7, 8.4, 10.7, 7.4, 6, 6.3, 4.9, 7.4, 4.4, 
    4.5, 4.6, 5.3, 6, 5.9, 5, 2.8, 2.6, 2.9, 4.7, 1.6, 2.1, 2.8, 3.2, 4.5, 
    1.8, 1, 2.2, 2.3, 0.9, 0.6, 0, 0.9, 3.2, 4.5, 3.4, 4, 4.4, 4.6, 3.8, 4.1, 
    4.6, 3.2, 3.7, 5.2, 5.8, 7.8, 7.2, 8.6, 8.5, 8.6, 8.1, 6.1, 6.4, 5.7, 
    6.5, 8.4, 7.1, 6, 5.9, 6.4, 6, 6.7, 6.3, 5.9, 5.3, 5.9, 5.1, 5.4, 5.7, 
    5.2, 4.3, 4.1, 3.8, 3.5, 4.3, 4.5, 4.6, 5.2, 5.1, 3.8, 3.8, 6, 3.6, 5, 
    7.6, 3.9, 5.3, 1.6, 5.2, 3.6, 9.6, 9, 9.2, 8.7, 8, 9.5, 4.5, 1.4, 2, 0.5, 
    0.9, 3, 4.6, 3.8, 3.7, 4.1, 5.9, 5.3, 4, 4, 3, 4.5, 4.7, 4.5, 4.9, 5.6, 
    4.8, 4.6, 4.1, 4.6, 5.7, 4.6, 4.3, 6, 7.1, 7.3, 7.3, 6.3, 5.9, 5.6, 6.6, 
    6.4, 7, 7.8, 8.9, 7.8, 9.1, 7, 7.2, 9.4, 8.7, 8.5, 7.6, 7, 9.6, 10.4, 
    10.4, 10.2, 10.1, 9.4, 8.9, 6.5, 5.7, 6.6, 5.2, 5.2, 3.5, 4.9, 2.9, 3.3, 
    6.8, 0.6, 2, 2.2, 0.4, 0, 0, 0.7, 2.9, 3.1, 0.6, 0.7, 3.8, 7.4, 8.5, 7, 
    7.2, 7.1, 7.3, 7.6, 11.8, 11.9, 11.7, 11, 10.8, 9.9, 8.7, 11, 8.3, 7, 
    8.1, 5.5, 4.8, 0.2, 2.3, 1.9, 0.9, 1.7, 3, 1.4, 2.5, 3, 4.5, 5.3, 5, 7, 
    7.1, 2.6, 0.3, 1.7, 0.4, 2.8, 2.1, 1.6, 3.8, 4.1, 3.9, 5.1, 6, 7, 8, 8.3, 
    7.6, 8.4, 9.3, 7.3, 9, 10.9, 12.3, 11.3, 10.2, 10.1, 8, 10.2, 9.6, 8.5, 
    8.2, 7.3, 6.7, 7.1, 6.3, 7.3, 7.8, 7.3, 6.4, 6.5, 6.7, 4.6, 3.4, 3.2, 
    4.5, 1.1, 0.6, 0.2, 2, 2.5, 2.1, 2.4, 1.8, 2.2, 3.6, 5.1, 4.8, 5.7, 4.5, 
    5.5, 5.1, 6.1, 6.4, 8.6, 6.3, 7.6, 4.8, 9.2, 9.7, 8.7, 5.4, 6.9, 5.1, 
    5.1, 5.7, 4.9, 1.6, 2.3, 2.2, 2.8, 1.8, 2, 1.4, 3.1, 2.2, 0, 1.6, 2.4, 
    1.8, 1.9, 2, 2, 2.1, 2.9, 3.9, 3.5, 5.4, 3.9, 3.7, 3.8, 5.4, 6, 9.2, 11, 
    10.7, 11.7, 11.2, 10.6, 9.5, 10.3, 9.5, 9.1, 11.6, 11.5, 12.2, 11.4, 
    10.8, 12.9, 9.8, 10.2, 11.5, 8.1, 6.7, 5.1, 3.6, 6.2, 6.9, 5, 4, 5.4, 
    3.2, 3.4, 1.8, 0.6, 1.3, 1.7, 3.7, 4.7, 4.6, 6.9, 8.3, 8.7, 9.8, 9.9, 
    10.7, 10.5, 5.9, 6.8, 5.1, 4.8, 3.6, 5.8, 6, 6.8, 6, 6, 5.9, 6.1, 6.3, 
    3.9, 2.9, 7.2, 5.7, 5.5, 7, 7.1, 6.6, 6.5, 5.7, 8.1, 8.4, 6.2, 7.3, 7.6, 
    6.6, 6.4, 5.6, 7.3, 5.3, 5.4, 7, 8.6, 6.6, 8.3, 7.1, 8.9, 9.7, 9, 9.8, 
    10.8, 9.6, 9.4, 9.8, 12.3, 10.7, 12.4, 12.9, 8.9, 10.3, 10.5, 9.3, 7.5, 
    7.2, 6, 9.2, 5.4, 7.4, 6.5, 6.7, 7.2, 8, 8.7, 6.8, 5.1, 8.7, 6.7, 8.2, 
    10.6, 9, 7.4, 4.7, 4, 6.1, 4.3, 4.9, 2.6, 0.9, 2.1, 2.8, 4.2, 3.6, 3.8, 
    2.9, 2.9, 1.9, 0.2, 0.8, 0, 0.7, 1, 2.6, 2.5, 2.8, 3.3, 4, 5.1, 6.8, 7.9, 
    7.4, 6.8, 3.6, 2.5, 13.2, 13.7, 15.2, 14.8, 16.1, 15.5, 15.3, 17, 14.8, 
    11.6, 9.7, 10.5, 11.3, 10.5, 11.6, 9.2, 9.8, 10.5, 12.4, 11.9, 12.5, 
    13.5, 11.6, 10, 10.2, 11.2, 10.3, 13, 14.4, 15.1, 13.3, 11.1, 11, 13.6, 
    13.2, 14, 11.8, 12, 11.8, 12.4, 12.4, 10.5, 9.8, 10, 7, 6.2, 11.7, 9.3, 
    7.5, 5.9, 6.2, 6, 4.7, 6, 5.2, 5.4, 4, 6.4, 8.4, 7.5, 4.6, 4.1, 6.1, 5.7, 
    6.1, 6.6, 4.8, 3.2, 3.4, 3.7, 6.2, 5.3, 3.9, 3.5, 3.6, 5.6, 6.1, 3.2, 
    4.6, 6.2, 5.4, 6.4, 9.7, 10.5, 10.7, 9.5, 11.5, 10.1, 7.1, 7.6, 8.4, 9.7, 
    1.8, 0.4, 1.1, 1.4, 2.6, 2.9, 3.5, 4.3, 1.2, 2.9, 4.3, 3.4, 1.5, 2.5, 
    2.5, 1.6, 2, 1.8, 2.1, 1.6, 1.9, 1.2, 1.7, 1.6, 0.4, 0.7, 0.1, 0.4, 1.3, 
    0.8, 2, 2.1, 1.6, 1.8, 1.8, 0.7, 1.4, 1.4, 0.1, 2.3, 1.7, 2.7, 3.2, 2.3, 
    0.9, 2.8, 3.1, 2.3, 2.7, 2.8, 3.4, 2.5, 2, 1.5, 2.2, 2, 2.7, 2.2, 1, 2.9, 
    1.7, 3.6, 4.4, 5.3, 3.8, 4.1, 3.9, 2.8, 4.8, 5.7, 3.3, 4, 4.2, 4.5, 5.9, 
    4.7, 5.2, 4.9, 5.7, 6, 5.6, 8, 7.4, 6.7, 7.5, 7.9, 8.6, 8.4, 9.1, 9.5, 
    9.6, 8.3, 9.8, 9.6, 11, 10.4, 9.7, 11.4, 11.9, 10.1, 12, 11.8, 12.4, 
    12.2, 14.1, 14.3, 13.6, 14.3, 14.3, 12.9, 10.7, 9.6, 8.7, 8.3, 7.2, 8.4, 
    8.6, 7.6, 8.9, 8.8, 7, 6.6, 6.8, 6.4, 8.4, 7.6, 5.8, 8.5, 8.8, 9.2, 10.5, 
    8.4, 10.3, 10.4, 9.7, 11.6, 11.6, 13.3, 13.2, 13.4, 11.1, 11.7, 12.7, 
    12.1, 11.5, 11.4, 9.3, 8.9, 6.8, 6.4, 5.6, 4.7, 3.5, 5, 4.9, 6.3, 5.9, 
    5.9, 7.6, 6.7, 6.2, 7.8, 7.2, 9, 10.1, 6.9, 7.4, 4.5, 2.9, 2.7, 1.8, 1.3, 
    3.3, 0.1, 1, 4.5, 7.8, 7, 7.5, 9, 11.5, 12.4, 11.3, 14.1, 12.7, 11.3, 
    12.3, 12.3, 13.9, 12.1, 12.7, 12.4, 11.5, 10.7, 12.3, 9.4, 10, 7.8, 8.4, 
    7.8, 4.5, 4.8, 4.6, 5.4, 2.4, 2.7, 4.1, 4.6, 3.9, 5.7, 2.9, 2.3, 2.9, 
    0.9, 1.7, 3.2, 3.5, 3.3, 4.6, 5.1, 6.1, 7, 7.1, 8, 7.9, 7.6, 8.3, 10.2, 
    11.1, 13.5, 14.5, 14.3, 14, 13.3, 11.3, 10, 7.2, 5.6, 5.9, 5.1, 3.9, 2.9, 
    3, 2.7, 1.7, 0.6, 0.4, 0.4, 3, 3.8, 2.3, 0.6, 0.3, 0.2, 0, 3, 2.1, 2, 
    0.5, 1.7, 7.9, 9.1, 10, 9.1, 9.7, 8.3, 7.2, 5.1, 7.7, 7.2, 8.4, 7, 8.8, 
    9.6, 9.4, 11.5, 11, 11.5, 10.6, 10.8, 11.1, 10.3, 9, 9.5, 9.4, 8.4, 8.5, 
    8.9, 9.5, 10, 10.6, 9.7, 8.6, 8.1, 7.7, 7.6, 7.1, 6.6, 6.5, 7.5, 7.7, 
    7.5, 5.6, 5.6, 4.7, 2.8, 3.5, 2.3, 2, 1.6, 1.5, 2.7, 3, 4.5, 3.6, 4.4, 
    7.5, 7.4, 6.4, 6.3, 4.2, 3.4, 4.5, 2.1, 2.8, 2, 1.4, 1.3, 9.8, 8.7, 11.1, 
    10.8, 8.8, 11.1, 10.3, 8.6, 12.2, 13, 9.8, 10.1, 10.3, 10.4, 11.9, 8, 
    10.3, 9.9, 10.6, 12.7, 12.3, 15, 15.4, 14.9, 15.9, 16.1, 15.2, 2.1, 4.9, 
    9, 10.9, 11, 5.2, 3.1, 2.3, 2.4, 1.8, 7.1, 3.2, 2.2, 4, 4.2, 3.7, 1.5, 1, 
    5.5, 1.8, 2, 1.5, 1, 2.4, 0.8, 1.6, 0.9, 2.8, 5, 1.6, 2.8, 1.2, 1.8, 9.5, 
    2.7, 4.9, 11.7, 9.6, 1.7, 0.7, 0.5, 7.4, 7.2, 2.8, 1.2, 3.4, 0.9, 0.2, 
    0.8, 0, 4.3, 1.3, 2.1, 1.8, 3.8, 3.7, 4.7, 4.7, 4.5, 5.1, 4.9, 5.5, 7.8, 
    8.1, 7.5, 7.9, 7.2, 8.8, 8, 9, 9.1, 9.5, 9.5, 8.5, 6.9, 8.3, 8.5, 7.1, 
    6.5, 5.4, 4.4, 3.3, 2.1, 2.5, 1.8, 1.6, 4.1, 6.4, 6.9, 6.6, 8.7, 8.6, 
    9.8, 10.3, 11.6, 12, 12.1, 12.1, 11.5, 12.2, 11.1, 13.5, 13.5, 12.8, 
    11.8, 12.3, 10.4, 11.5, 12, 10.7, 11.6, 11.6, 10.7, 12.5, 12, 11.3, 11.8, 
    11.6, 12, 12.5, 12.8, 14.7, 14.6, 15.1, 13.2, 14.5, 11.5, 12.7, 13.6, 12, 
    13.1, 14, 12.6, 14.9, 11.6, 12.2, 12.6, 11.7, 11.9, 10.5, 9.7, 9.6, 11.1, 
    8.3, 11.2, 10.1, 12.5, 11.3, 8.7, 10.2, 10.1, 12.5, 6.8, 8.9, 11.7, 15.4, 
    12.4, 10.2, 12.8, 14.2, 14, 14.4, 15.9, 15.1, 12.8, 14.7, 14, 16, 14.5, 
    12.9, 16.4, 13.9, 13.2, 11.8, 13.7, 14, 13.7, 13.6, 12.5, 14.3, 13.4, 
    13.5, 12, 12.7, 15.1, 12.4, 14, 13.3, 14.2, 14.7, 16, 16.8, 18, 17.9, 
    17.1, 12.5, 19.9, 17.2, 16.1, 14.8, 15.7, 14.8, 15.7, 14.6, 13.4, 14.1, 
    15.2, 15.4, 14.7, 15.9, 14.2, 13.4, 15.6, 15.5, 16.7, 14.8, 13.8, 13.9, 
    12.8, 14.3, 14.1, 13.6, 13.6, 13, 12.8, 14.6, 14.8, 14.1, 13.8, 12.4, 
    12.1, 14.6, 15.1, 15.5, 15.4, 15.3, 19.2, 20, 19.7, 17.9, 14.3, 15.4, 
    11.9, 13.8, 14.3, 15.2, 14.6, 15.5, 14.8, 13.8, 15.7, 18.8, 17.3, 17.9, 
    15.2, 17.1, 17.6, 16.7, 15.6, 15.2, 16.1, 5.4, 4.4, 14.1, 13.4, 14.2, 
    14.9, 11.1, 15, 13.5, 11.1, 6.5, 6.5, 4.2, 1.9, 0.4, 0.2, 2.8, 1.8, 2.4, 
    3, 9.6, 6.7, 3.1, 3, 3.9, 4.6, 5.6, 4.7, 5.6, 5.9, 5.2, 4.9, 6.9, 8.9, 
    7.2, 6.9, 4.7, 5.3, 2.9, 5.4, 1.2, 3, 2.9, 5, 6.8, 4, 8, 6.3, 3.7, 2.5, 
    10.6, 12.9, 9.7, 8.4, 8.7, 3.8, 5.6, 8.6, 10.1, 11.6, 11.1, 9.2, 11.7, 
    10.9, 6.8, 8.3, 6.2, 7, 10.1, 10, 10.6, 9.7, 9.6, 7.2, 11, 9.3, 10.2, 8, 
    9.9, 10.6, 9.7, 8.4, 11.5, 9.9, 8.6, 8.2, 7.7, 7.3, 7.6, 7.7, 9.2, 9.7, 
    9.1, 8.7, 11.3, 9.1, 7.8, 7.2, 5.2, 7.1, 8.1, 7.2, 5.6, 5.3, 5.4, 5.7, 
    5.8, 6.6, 6.3, 3.3, 3.4, 2.7, 1.4, 1.8, 1.8, 2.2, 0.6, 1.3, 0.6, 0.5, 
    2.2, 3.1, 3.3, 2.6, 0.8, 0.1, 0.8, 1.2, 4.4, 4.8, 5.5, 6, 4, 4.2, 2.6, 
    5.4, 4.5, 5.4, 7.7, 5.9, 6.7, 7.6, 7.3, 7.9, 7, 6.6, 6.6, 9.4, 7.3, 4.1, 
    3.6, 4.8, 5.2, 11.1, 11.5, 10.1, 8.5, 8.5, 8.6, 8.1, 7.7, 6.6, 5.5, 5.5, 
    6.1, 6.1, 6.3, 4.6, 3.7, 4.9, 4.2, 5.5, 5.8, 5.6, 6.3, 7.9, 6.9, 6.6, 
    6.7, 7.1, 8.3, 8.4, 6.2, 6.7, 5.6, 5.1, 4.8, 3.8, 6.3, 4.4, 4, 2.9, 4.2, 
    4.2, 3.1, 2.8, 1.5, 3.2, 5.7, 6.7, 6.1, 5.3, 4.6, 1.2, 3.7, 3.6, 2.7, 
    2.4, 3.1, 2.5, 11, 10.8, 12.9, 12.1, 12.7, 10.3, 9.2, 9.4, 10.6, 8.7, 
    10.5, 9.5, 7.2, 7.1, 4.7, 2.7, 4.4, 2.6, 4.3, 4.4, 6.8, 6.1, 3.2, 3, 4, 
    4.5, 4.4, 3.1, 4, 6.3, 4.2, 5.1, 8.4, 8, 7.1, 7.5, 7.7, 6.6, 7.4, 6.3, 
    6.5, 7.1, 7.2, 5.7, 4.9, 5.1, 5.1, 5.8, 6.3, 6.5, 6, 6.4, 6.2, 5.4, 2.7, 
    2.2, 2.7, 3.7, 3.7, 6.2, 2.4, 4.8, 5.1, 5.7, 5.1, 7.5, 6.1, 6.5, 5.9, 
    6.3, 5.9, 5.6, 5.5, 3.7, 3.8, 4.7, 4, 3.1, 2.6, 1.8, 2.6, 3.2, 2.8, 3.6, 
    3.6, 3.1, 3.6, 3.1, 3.2, 3.2, 3.1, 2.4, 2.4, 3.6, 6.1, 4.7, 4.1, 4.5, 
    3.6, 3.7, 3.1, 3.8, 3.6, 3, 3, 2.8, 2.8, 4.7, 7.1, 3.9, 9, 9.6, 8.8, 
    11.6, 8.5, 9.8, 8.6, 11.1, 9.5, 9.8, 10.1, 7.5, 8.7, 3, 2, 9, 9.5, 9.9, 
    10, 9.8, 11, 11.1, 10.6, 10.5, 11.6, 11.5, 8.3, 6.7, 9.2, 8.8, 10.3, 7.1, 
    7.3, 10.2, 8.5, 11.4, 7.7, 7, 5.6, 4.5, 5.9, 4.5, 5.1, 4.4, 6, 7.1, 5.5, 
    6.6, 6.6, 7.4, 7.8, 2.6, 4.5, 0.8, 0.9, 2.6, 4.9, 5.8, 5.2, 2.2, 3.9, 3, 
    1.1, 1.6, 5.4, 5.6, 6.6, 7.8, 4.3, 6, 4.9, 5.6, 4.7, 5.7, 6, 7.1, 8, 8.8, 
    6.9, 7.2, 5.9, 8.4, 8.4, 7.6, 7.6, 6.6, 6.7, 5.2, 4.4, 4, 2.4, 3.8, 5.5, 
    8.3, 8.1, 12, 11.1, 11.2, 11.5, 12.3, 11, 12.1, 11.5, 11.6, 9.3, 8.1, 
    8.6, 6.7, 7.9, 4.2, 6.6, 6.7, 5.9, 5.9, 3.4, 2.5, 2.8, 2.3, 4.3, 2.1, 
    2.4, 1.3, 2.6, 1.4, 2.9, 2.6, 3.7, 5.6, 5.9, 5.6, 6, 5, 4.4, 4.9, 4.9, 
    5.7, 6.9, 5.9, 6.4, 6.7, 8, 5.7, 6.1, 5.6, 4.6, 3.8, 4.1, 5.3, 5, 3.9, 
    0.8, 2.3, 2.9, 5.4, 7.8, 8.4, 3.8, 3.8, 4.7, 5.8, 9.2, 7.8, 7.5, 8.3, 
    7.5, 8.4, 10.2, 9.1, 10.8, 11.1, 9.9, 10.6, 9.9, 9.3, 9.7, 10.1, 8.3, 
    8.9, 10.9, 9.8, 9, 9.7, 11, 11.4, 12.1, 10.9, 11.9, 10.9, 9.8, 9.2, 9.2, 
    10.5, 10.1, 9.6, 11.5, 8.4, 9, 10, 9.5, 8.2, 8.6, 8.9, 8.9, 8.5, 9.1, 
    9.2, 8.9, 9.7, 8.3, 8.9, 8.2, 7, 8.1, 7.5, 7, 6.7, 7.2, 9.3, 7.3, 5.9, 
    4.6, 1, 2, 4.2, 4.1, 4.6, 5.3, 4.9, 2.1, 3.3, 3, 4.4, 11.9, 11.7, 13.5, 
    14.8, 16.9, 17.2, 15.5, 15.3, 16.2, 13.5, 11.7, 11.2, 8.6, 9.1, 8.3, 8.7, 
    7.4, 4.8, 3.4, 3, 2, 2.1, 2.3, 3, 3.8, 2.8, 3.2, 5.5, 6.7, 6.8, 7.9, 6.2, 
    8.8, 8.1, 8.4, 7.4, 8.6, 6.9, 5, 6.4, 5.5, 6.2, 5.4, 6.2, 7.1, 5.9, 4.5, 
    6, 5.3, 3.8, 5, 7.6, 7.4, 7.9, 7.7, 7, 7.9, 4.6, 6.1, 6, 4.4, 3.7, 3.1, 
    1, 1.2, 2.1, 3.2, 4.9, 4.8, 5.8, 5.6, 5.6, 5, 4.4, 4.5, 6, 3.7, 3.4, 2.6, 
    3, 4.5, 3.5, 2.9, 4.3, 5.2, 5.8, 4.4, 6.8, 7.5, 6.4, 8.3, 8.2, 6.9, 6.3, 
    6.9, 7.7, 7.9, 6.2, 6.3, 7.2, 5.8, 5.6, 7.4, 7.6, 8.9, 8.1, 7.4, 5, 8, 
    8.3, 7.4, 7.1, 6.4, 8, 6.6, 8.6, 6.9, 7.2, 5.9, 5.9, 6.4, 6, 7.5, 7.7, 
    6.2, 7, 6.4, 5.9, 7.4, 8, 7.2, 9.7, 12.3, 12.6, 11.9, 9.1, 9.2, 11.3, 
    12.5, 11.7, 11.9, 10.8, 12.2, 11.5, 9.2, 8.8, 9.3, 10, 11.3, 11.7, 11.6, 
    13, 11.3, 11.1, 12.5, 9.2, 9, 8.2, 9.6, 10.9, 10.2, 10.5, 10.3, 10.2, 
    11.7, 9.9, 7.6, 7.7, 4, 6, 7, 5.4, 4.8, 6.1, 5.6, 8.5, 6.5, 6.2, 5.1, 
    5.4, 2.6, 0.9, 7.3, 2.6, 9.3, 9.8, 3.9, 3.2, 12.3, 6.7, 3.4, 7.2, 13.7, 
    13.4, 12, 13.1, 14.1, 13.4, 13.2, 12.5, 12.7, 12.2, 0.5, 2.1, 2.1, 4.2, 
    7.7, 10.3, 9.1, 8.6, 4, 3.9, 1.2, 1.8, 1.8, 2.2, 5.7, 7.6, 3.2, 6.9, 5.7, 
    2, 2.7, 2.9, 3.5, 4.1, 3.6, 4.6, 5.2, 4, 2.8, 5, 4.8, 3.4, 4.3, 4.8, 2.9, 
    4.2, 3.6, 2.4, 1.3, 2.1, 3.7, 2.4, 1.8, 1.6, 0.9, 2.5, 4.7, 4.3, 3.9, 
    4.6, 4.4, 6.2, 5.4, 4.5, 5.6, 7, 6, 6.3, 6.2, 5.8, 4.3, 5.4, 6.7, 5.9, 
    5.7, 6.2, 5.1, 5.2, 4.7, 4.1, 4.5, 6, 7.6, 6.2, 7.3, 7.3, 7.4, 12.9, 
    11.4, 9.8, 11.3, 12.8, 14.7, 17.5, 16.2, 18.8, 18.2, 17.5, 19.2, 17.4, 
    18.2, 17.9, 17.4, 18, 17.2, 20, 17.8, 15.3, 16.5, 13.6, 17.6, 15.9, 15.6, 
    14.1, 14.5, 14.8, 12.9, 13.4, 12.3, 12.8, 10.9, 11, 12, 13.8, 11.4, 7.1, 
    8.3, 5.7, 6.4, 5.8, 4.2, 4.1, 6.5, 5, 6, 5.1, 3.3, 2, 4.9, 4.9, 5.6, 7, 
    8.7, 8.4, 8.6, 11, 11.9, 13, 10, 6.5, 5.9, 6.6, 8, 10.7, 8.5, 10.6, 7.3, 
    10.6, 10.9, 9.2, 7.8, 7.9, 8.4, 9.2, 5.4, 6.1, 7.6, 5.6, 8.7, 9.3, 9.5, 
    9.3, 12.9, 11.5, 11.5, 13.8, 11.2, 7.7, 7.2, 4.5, 3, 2.5, 6.4, 7.8, 7.7, 
    8.1, 6.8, 7.6, 6.6, 7.4, 5.9, 7.5, 6.6, 4.5, 6.7, 7.7, 8.3, 7.2, 8.5, 
    8.2, 8.6, 9.5, 4.6, 9.4, 5.3, 7.5, 5.6, 3.2, 7.5, 7.1, 5.2, 5.1, 10.5, 
    4.5, 4.3, 7.3, 11.5, 11.7, 9.7, 9.2, 9.1, 10.3, 10.3, 8.5, 8.8, 7.6, 8.4, 
    9.6, 7.7, 9.3, 7.5, 6.6, 8, 7.5, 7, 6, 7.4, 7.9, 4.2, 5.4, 3.9, 7.4, 7.1, 
    6.9, 8.1, 7.3, 4.3, _, 1.1, 0.9, 3.3, 2.1, 2, 1.6, 2.5, 2.1, 2.3, 2.3, 
    4.1, 5.6, 5, 4.2, 5, 5.4, 4.8, 5.2, 6.3, 5.5, 4.8, 6.6, 8, 5.1, 3.3, 6.9, 
    6.7, 8, 7.7, 7.6, 8.1, 10.1, 8.9, 9.4, 11.6, 8.1, 6.8, 10.8, 17.5, 17, 
    18.9, 18.1, 14, 11.1, 9.3, 8.8, 8.7, 8.6, 8.9, 10.3, 9.9, 9.4, 9.7, 8.9, 
    8.9, 8.9, 9.4, 9.7, 10.5, 10.4, 10.1, 11.4, 12.4, 12.1, 11.7, 10.8, 11.4, 
    12, 9, 10.4, 10.4, 9.9, 10.1, 10.4, 9.5, 10.4, 10, 10.2, 10.3, 9.7, 9.8, 
    10.6, 10.2, 9.8, 11.2, 10.6, 9.3, 8.6, 9.3, 9.2, 8, 5.8, 5.1, 7, 6.4, 
    6.6, 7.2, 8.6, 8, 9.6, 9.7, 9.6, 9.3, 8.8, 9.2, 9.5, 8.9, 7.5, 6.9, 7.2, 
    7.2, 6.7, 6.8, 6.3, 5.3, 5.1, 4.2, 3.5, 4.2, 4.1, 5, 4.9, 5.4, 6.7, 5.9, 
    6.5, 5.3, 5.9, 7.1, 8, 8.5, 8.9, 7.3, 6.5, 7, 6.4, 5.1, 4.8, 5.4, 4.6, 
    5.4, 8.5, 7.5, 6.5, 10.4, 5.6, 5.7, 6.7, 6, 7.4, 8.3, 8.8, 9, 10, 10.8, 
    9.2, 9.7, 11.6, 13, 13.2, 12.1, 9.1, 10.8, 9.8, 10.8, 9.7, 12.6, 14.1, 
    9.5, 16, 17, 15, 16.9, 14, 15.2, 16.1, 13.4, 15.2, 13, 13.6, 14.3, 14.7, 
    15.3, 16.2, 14.8, 15, 15.1, 14.4, 15, 14.6, 13.6, 13.9, 13.8, 12.7, 13.8, 
    14.3, 12.4, 12.7, 12, 13.6, 14.1, 13.4, 16.2, 15.5, 15.8, 16.2, 19.4, 
    18.5, 19, 19.5, 20.2, 18.5, 19.8, 23.4, 22.5, 21.8, 22.5, 21.2, 22.2, 
    21.1, 21.7, 19.5, 20.8, 20.8, 19.4, 18.6, 20.2, 18.8, 18.1, 17.6, 18, 
    19.2, 17.1, 19.2, 19.6, 18.7, 18.9, 20.1, 19.5, 20.7, 20.4, 20.3, 21.2, 
    18.6, 21.6, 20.5, 19.2, 20.6, 21, 18.8, 18.6, 18.9, 19.3, 18.7, 17.4, 
    17.6, 15.6, 16.8, 14.5, 14.7, 13.4, 14, 11.9, 10.7, 9.6, 8.9, 9.5, 12.4, 
    11.8, 11.4, 12.6, 11.3, 12.7, 11.8, 14.3, 16.2, 14.6, 15.1, 14.5, 13.8, 
    14.4, 13.1, 12, 12.3, 12.3, 10.7, 9.3, 9, 6.5, 7.5, 6.7, 4.4, 5.5, 7.8, 
    6.8, 6.1, 5.6, 5, 3.8, 3.5, 3.3, 4.7, 4, 3.1, 5.5, 5.8, 5, 5.3, 6.7, 7.3, 
    8.3, 7.8, 6.5, 9.3, 9.5, 11.9, 10.9, 12.5, 8.3, 6.4, 7.4, 7.1, 12.9, 
    15.6, 11.4, 8.8, 9.3, 8.2, 8.2, 8.5, 9.9, 7.6, 6.1, 4.4, 6.2, 9.7, 11, 
    11.5, 12, 11.4, 11.8, 13.2, 11, 13, 13.2, 12.9, 14.5, 11.2, 13.1, 12.2, 
    12.3, 13.2, 12.5, 16.3, 12.2, 10.5, 8, 8.3, 8.5, 6.2, 6.5, 7.7, 4.7, 7.3, 
    8.4, 7.7, 8.6, 7.8, 8.9, 9.1, 11, 9.9, 9.8, 8.2, 5.9, 4.2, 5, 3.8, 3.7, 
    4, 3.1, 3.1, 6.6, 4.7, 5.2, 5.8, 6.1, 6, 5.7, 6.4, 8.1, 6.7, 6.7, 8.2, 
    7.5, 7, 7.2, 4.6, 5.5, 5.8, 5.2, 4.5, 6.1, 6, 10.1, 5.9, 4.1, 7.6, 7.3, 
    9, 9.3, 11.6, 10.5, 9.3, 6, 5.6, 6.9, 8.6, 12.5, 15.8, 16.8, 13.6, 16.1, 
    16.4, 14.7, 14.4, 12.4, 9.2, 9.5, 8.9, 10.2, 10.2, 7.9, 9.1, 8.3, 8.2, 
    7.1, 8.7, 10.7, 11.3, 9.5, 8.3, 8.6, 9, 8.2, 7.5, 8.3, 7.1, 7.7, 6.6, 
    4.7, 3.8, 2.8, 3.4, 3.5, 3.8, 6.6, 7.6, 7, 6.3, 5.3, 5.1, 5.1, 5.4, 5, 
    5.1, 3.4, 4.2, 5.9, 4.8, 5.4, 4.7, 4.3, 3.8, 3.6, 3.1, 2.5, 2, 2.3, 2.2, 
    6.3, 5.9, 7.3, 8.3, 9.1, 8.5, 8, 8, 9.1, 8.5, 7.8, 7.9, 9.3, 8.5, 8.6, 
    10.2, 10.6, 8.2, 9.1, 10.3, 6.8, 7.1, 6.1, 5, 7.7, 4.9, 6.3, 8.8, 6.1, 
    5.1, 5.1, 6.6, 8.5, 6.6, 7.7, 6.6, 6.5, 7.3, 9.5, 8.7, 9.3, 7.7, 9.1, 
    6.8, 5.5, 6.5, 5.2, 5.4, 4, 2.7, 1, 3.1, 2.1, 3.3, 5.5, 6.2, 10.2, 10.1, 
    5.3, 7.9, 6.5, 8.5, 8.6, 6.7, 6.8, 8.1, 8, 8.7, 8.2, 8.2, 8.2, 7.7, 7.1, 
    4.6, 3.3, 2.1, 5.7, 6, 6, 5.6, 7.5, 6.3, 6, 11.2, 8.5, 10.7, 10.8, 10.6, 
    10.8, 10.9, 10.9, 10.9, _, _, 11.7, 11.6, 13.4, 13.1, 12.8, 11.5, 11.3, 
    14.1, 13.7, 14.7, 11.3, 12.3, 12.6, 10.9, 9.1, 9.4, 8.6, 7.7, 8.7, 7.5, 
    7.9, 9.9, 10.6, 11.4, 5.3, 9.2, 9.2, 5, 5.7, 5.8, 5.3, 3.6, 5, 6.5, 6.8, 
    6.9, 7.6, 7.3, 8.2, 8.6, 8.1, 7.5, 7.6, 6.9, 8.5, 7, 8.9, 8.4, 8.3, 7.5, 
    7.5, 9.8, 9.4, 8.1, 10.1, 10.5, 10.2, 9.4, 6.9, 7.1, 7, 7.2, 8.2, 10.8, 
    11.6, 11.1, 10.1, 9.2, 8.3, 7, 7.7, 7.6, 7.6, 7.1, 7.5, 7.5, 9, 6.7, 8.4, 
    7.1, 7.5, 10.2, 9.4, 5.3, 10.1, 14.1, 8.4, 8.4, 9.3, 8.6, 9.2, 8.7, 6.7, 
    11.8, 9.3, 8.8, 7, 1.9, 6.6, 2.5, 3.8, 4, 4.7, 4.8, 5.5, 5.3, 4.4, 4.9, 
    3.9, 7.2, 6.2, 5.4, 8.5, 10.1, 8.1, 3.7, 6.1, 7.8, 10.1, 8.8, 8.9, 9.2, 
    10.1, 10, 9.3, 11, 9.2, 6.9, 6.8, 6.6, 7.6, 9.6, 8.8, 5.4, 1.5, 3.1, 2.3, 
    1.3, 1.1, 4, 2.8, 2.6, 3.1, 4.3, 4.8, 5.4, 4.5, 4, 4.7, 4.2, 4.6, 2.4, 
    4.4, 3.9, 5.6, 6.4, 5.8, 7, 8, 5.3, 3.5, 4.3, 4.6, 4.9, 3.7, 4, 4.8, 7.5, 
    3.3, 4.9, 6.7, 5.2, 6.2, 6.8, 5.9, 3.7, 4, 4.4, 6.2, 4.7, 4.8, 5.1, 5.7, 
    5.2, 5.3, 4.2, 5.3, 8.9, 4.7, 5.2, 4.7, 3, 6.5, 7.1, 7, 7.7, 7.4, 6.9, 
    7.5, 7.5, 6.3, 7.4, 5.9, 7.6, 7.5, 5.9, 6.7, 6.5, 8.5, 6.7, 8.9, 7.6, 
    7.5, 7.9, 7.9, 8.8, 7.8, 6.9, 6.9, 7, 5.5, 4.4, 5.8, 5.5, 5.6, 6.3, 5.3, 
    4.4, 4, 3.7, 3.5, 1, 1.8, 3, 4.1, 4.4, 6.4, 4.3, 3.8, 3.6, 2.4, 4.2, 3.7, 
    2.4, 2.1, 1.7, 2, 1.6, 3, 4.5, 5.9, 5.1, 2.8, 0.6, 2.2, 1.2, 4.9, 4.7, 
    8.2, 8.8, 10, 3.7, 5.4, 6.1, 8.2, 7.5, 7.9, 6.8, 5.8, 3.5, 4.3, 7.1, 7.5, 
    9, 7.9, 7.3, 8.6, 9.5, 8.7, 10.1, 10.7, 10.3, 10.3, 9.7, 8.7, 7.9, 8.3, 
    6.8, 8.5, 6.9, 8, 7.5, 8.3, 8.2, 7.2, 4.7, 5.4, 8.8, 9.4, 9.5, 8.4, 10.1, 
    9.9, 10.3, 9.4, 11.8, 13.2, 9.1, 12.9, 13.3, 12.7, 12.3, 12.8, 11.8, 11, 
    10.2, 9.9, 7.8, 8.6, 8.4, 9.3, 8.5, 7.3, 7.6, 8.4, 7.8, 8.1, 8, 6.6, 7.3, 
    1, 12.3, 11.2, 13, 13.1, 12.3, 14.1, 13.2, 10, 12.9, 13.9, 15, 16.5, 
    13.6, 16.1, 13.5, 6.2, 5.3, 11.4, 12.5, 13.2, 13.2, 13.5, 13.9, 12.5, 
    12.6, 10.8, 9.1, 0.6, 1, 2.1, 2.6, 3.5, 5.3, 4.6, 4.4, 3.7, 3.8, 4.4, 
    4.4, 3, 3.2, 3.7, 3.6, 3.9, 3.9, 5.8, 9.5, 10.6, 10.7, 10.4, 10.2, 12.1, 
    12.9, 14.9, 14.8, 15.6, 16.9, 16.2, 14.6, 13.2, 14.1, 12.4, 11.9, 11.9, 
    11, 10.9, 11, 11.4, 10.5, 12.1, 12, 10.6, 9.3, 10.6, 10.6, 9.2, 9, 9.4, 
    8.4, 6.9, 6.2, 4.9, 5.6, 8.4, 8.1, 8.7, 6.7, 8.3, 8.7, 7.1, 7.1, 8.2, 8, 
    8, 8.2, 9.2, 10.1, 10.4, 12.7, 11, 10.5, 10.6, 11, 10.4, 9, 8.3, 9.6, 
    8.6, 9.4, 9.2, 8.8, 8.7, 11.4, 9.3, 9.6, 10.2, 8.3, 9.2, 10.8, 11.8, 9.8, 
    9.6, 10.2, 11.7, 10.1, 10.4, 10.9, 10.4, 9.6, 9.5, 10, 7.9, 10.6, 10.2, 
    9.6, 8.3, 7.4, 9.5, 7.4, 7.8, 6.6, 8.1, 8.6, 7.6, 8.5, 6.6, 7.4, 6.8, 
    7.1, 7.1, 7.8, 5.7, 5.6, 6.3, 5.9, 7.5, 8.4, 6.7, 7, 7.2, 6.8, 7.1, 8.2, 
    8.7, 9.6, 10.3, 9.1, 9.6, 9.2, 8.4, 8.7, 9.9, 8.7, 8.9, 7, 8.9, 8.4, 7.1, 
    8.4, 5.1, 6.4, 6.7, 4, 5.1, 6.1, 6.9, 7.8, 7.4, 9.1, 10.2, 8.6, 8.2, 9.6, 
    9.8, 10, 10.9, 8.9, 10.3, 11.4, 10.4, 10.5, 11.3, 11.5, 10.3, 8.8, 9.1, 
    8.6, 5.8, 8.8, 4.3, 7.5, 9.1, 8.9, 8.9, 7.3, 7.5, 6.1, 7.2, 10.4, 12.6, 
    14.2, 16.1, 19.6, 18.8, 13.2, 14.5, 11.4, 13.1, 10, 10.3, 11.5, 8.2, 
    10.6, 9.7, 10.9, 9.6, 7.5, 11.2, 9.2, 9.6, 10.8, 9.2, 11.1, 11.3, 8.7, 
    8.4, 9.8, 9.5, 9.6, 6.6, 8.1, 7.1, 6.1, 5.6, 5.9, 4.9, 4, 4.9, 4.1, 4.7, 
    4.3, 2.8, 3.6, 2.8, 3.5, 4.5, 4.1, 6.7, 8.8, 9.2, 11.2, 12, 13.8, 11.1, 
    11.4, 13.7, 15.3, 15.6, 13.3, 12.3, 13.1, 8.1, 8.7, 16.7, 16.9, 15.3, 
    13.2, 15, 12.9, 11.5, 10.5, 12.2, 12.4, 11, 12.2, 10.6, 8.4, 10, 10.2, 
    9.9, 10, 8.4, 6.7, 5.2, 5.5, 6, 5.2, 5.3, 7.4, 5.9, 9.1, 7.3, 7.7, 5.8, 
    6, 4.8, 6.4, 5.4, 7.6, 9.2, 9.8, 11.4, 10.3, 10.1, 9.7, 14.2, 14.9, 17.7, 
    16.9, 18.8, 19.3, 20.7, 21.5, 23.7, 25.7, 27.8, 28.1, 26.2, 24.9, 14, 
    19.8, 8.4, 7.2, 8.5, 9.3, 9.7, 9.3, 8.2, 10.9, 11.5, 11.9, 8.9, 8.3, 9.4, 
    7.2, 9.9, 5.5, 5.1, 5.6, 7.8, 14.9, 20.6, 17.3, 17.7, 15, 15.5, 18.9, 
    18.7, 17.3, 18, 21.4, 20.1, 17.1, 14.1, 16.7, 12.2, 10.9, 11.2, 8.3, 9.9, 
    10.1, 8.5, 7.4, 6.1, 6.5, 5.9, 5, 5.2, 5.2, 4.7, 4.6, 4, 5.5, 6.2, 6.2, 
    5.8, 9.2, 7.1, 10.9, 11.1, 11.2, 12.9, 11.8, 10.4, 10.4, 11.3, 12.8, 
    11.9, 11.7, 10.6, 10.2, 10.4, 9.7, 11.5, 12.2, 9.4, 9.4, 9.4, 8.3, 8, 
    8.2, 5.6, 5, 6.2, 8.6, 6.1, 4, 4.3, 4.5, 3.9, 3.3, 4.6, 8.7, 3.5, 3.1, 
    4.9, 4.2, 4.6, 10.1, 9.2, 7.3, 8.8, 11, 8.1, 6.7, 7.4, 6.5, 8.3, 7.4, 
    7.3, 6.7, 4.3, 5, 7.1, 8.4, 8.5, 10.1, 10.1, 13.9, 12.6, 21.6, 14, 14.3, 
    19.6, 23.8, 23, 22.2, 17.5, 16.2, 14.5, 14, 13.2, 10.7, 11.3, 6.2, 5.7, 
    3.5, 2, 2, 2.8, 2.6, 2.9, 3.5, 3.4, 4.3, 3.2, 1, 0.8, 1.1, 2.7, 2.9, 1.6, 
    2.5, 2.5, 1.8, 2.7, 2.6, 3.9, 4.2, 3.4, 3.3, 3.1, 3.1, 3.7, 3.1, 3.5, 
    3.9, 4.9, 4.4, 7.2, 10.1, 10.6, 11, 16.6, 16.8, 14.9, 14.6, 15.2, 14.8, 
    15.4, 16.1, 16, 15.6, 15.2, 15.7, 17.7, 17.8, 17.9, 18.7, 19.5, 19.4, 
    17.1, 18, 19.7, 19.9, 19.8, 20.2, 19.6, 19.3, 20, 17.4, 18.2, 8.2, 7.2, 
    7.6, 8.3, 9.3, 8.8, 9, 6.4, 7.4, 7, 9.1, 9.8, 8.1, 8.3, 8.8, 9.7, 10.3, 
    10, 10.6, 10.9, 11.4, 13.2, 14.6, 13.4, 13.1, 14.2, 13.9, 14.2, 15.2, 
    15.2, 15.2, 15.2, 16.4, 16.6, 16.4, 18.5, 17.1, 15.7, 16.1, 16.1, 16.3, 
    18, 18, 18.3, 16.7, 15.8, 15.8, 15.6, 16.7, 18, 16.6, 17.7, 19.7, 19.6, 
    19.1, 18.6, 18.3, 18.5, 16.1, 18.2, 18.3, 17.2, 19.5, 18.4, 18.2, 19.5, 
    19.4, 19.5, 19.6, 20.5, 20.8, 20.4, 19.8, 20.6, 19.3, 19, 18.4, 18.6, 20, 
    19.1, 19.9, 18.1, 19.9, 19.6, 20, 20.5, 22.1, 20.8, 19.9, 19.7, 18.9, 
    19.5, 18.8, 17.8, 20.8, 20, 18.1, 17.3, 17.6, 19.2, 19.7, 18.2, 17.9, 
    19.4, 20.5, 16.9, 16.9, 16.7, 15, 16.3, 16.6, 17.2, 14.4, 16.5, 16.6, 
    15.5, 13.5, 10.4, 12.4, 11.8, 12.9, 12, 11.8, 9.8, 10.7, 11.7, 8, 7.4, 
    7.5, 12.8, 7.1, 7.6, 6.8, 8, 7.4, 7.4, 7, 6.7, 6.4, 11, 9.7, 10.8, 9.4, 
    13, 13.9, 10.5, 10, 9.4, 7.8, 7.1, 8.9, 8.6, 5.5, 5.4, 2.4, 4.1, 3.4, 
    7.9, 6.4, 7.1, 4.7, 5.6, 6.7, 8.2, 6.6, 7.7, 6.3, 7.9, 7.9, 7.8, 8.5, 
    9.5, 9.4, 10.6, 12, 12, 13.3, 12.3, 15, 15.8, 16.8, 17.4, 17.6, 18.9, 
    20.4, 20.5, 20.6, 20.3, 21.3, 20.7, 20.4, 20.7, 21.9, 21.1, 21.6, 21.4, 
    21.9, 20.7, 22.2, 19.2, 20.3, 20.6, 19.5, 19.4, 18.3, 16.4, 16.4, 15.4, 
    12.7, 8.7, 5.4, 1.2, 1.7, 1.5, 2.4, 4.2, 2.6, 4, 5.5, 4, 5.1, 5.9, 5.8, 
    7.4, 5, 2.1, 5.7, 4.1, 6.3, 7.3, 5.6, 6.9, 3.9, 2.4, 3.3, 10.4, 10.8, 
    10.5, 10.6, 11.2, 11.5, 11.2, 11.4, 10.2, 11.4, 10.6, 10.9, 9.8, 11.2, 
    9.6, 10.8, 12.6, 12.8, 8.5, 8.8, 7.9, 7.3, 6.6, 6.1, 4.8, 5.9, 7.2, 4.9, 
    2.5, 2.7, 1.8, 3, 5, 4, 4.3, 3.9, 4.3, 3.4, 2.6, 4.1, 6.1, 6.3, 6.2, 6, 
    5.1, 5.5, 6.3, 5.6, 6.8, 8.1, 8.3, 6.5, 7.8, 9.2, 8.7, 6.5, 5.1, 3.3, 
    2.2, 2.4, 7.9, 2.6, 13, 7.2, 13.7, 13, 12.2, 9.6, 7.4, 4.2, 11.3, 8.5, 
    10.2, 7.1, 7, 5, 11.2, 12.4, 12.7, 11.5, 11.4, 7.5, 7.6, 8.4, 10.1, 8.6, 
    12, 13.4, 15.3, 15.4, 14.6, 16.5, 15.7, 16.1, 20, 19.5, 18.9, 19, 20, 
    19.9, 21.2, 20.6, 16.4, 19.7, 19.7, 17.6, 18.1, 22, 18.2, 18.6, 16, 16.2, 
    15.5, 17.1, 18.3, 17.4, 17.1, 16.9, 15.1, 15.3, 17.4, 15.6, 15.2, 12.5, 
    13.6, 12, 8.8, 9.9, 7.8, 7.8, 8.7, 8.3, 6.8, 5.3, 5.6, 5.5, 5.7, 6.1, 
    5.9, 6.5, 6.6, 4.9, 7, 5.4, 4.8, 6.9, 4.9, 6, 4.1, 5.4, 5.7, 5.4, 3.9, 
    3.6, 5, 2.5, 4.4, 5.7, 5, 5.2, 5.6, 4.4, 4.2, 5.2, 4.6, 4, 4.3, 5.2, 4.1, 
    4.1, 4.6, 4.3, 4.3, 4.8, 4.9, 5.2, 6.5, 6.2, 7, 7.5, 7.5, 8.2, 7.9, 8.1, 
    8.1, 9.8, 9.5, 11.3, 9, 12.7, 11.4, 12.7, 11.7, 12.6, 13.7, 11.9, 14.2, 
    14.7, 14.2, 17.1, 18.8, 18.8, 17.6, 18.3, 18.2, 18.8, 17.6, 15.9, 17.5, 
    15.7, 15.6, 16.6, 18.3, 19.1, 21.2, 21, 22, 20.9, 22.9, 21, 18.3, 17, 
    17.4, 16.4, 14.1, 13.5, 14.8, 16.4, 15, 18.2, 14.8, 14.6, 13.1, 13.6, 9, 
    14.3, 13.8, 15.8, 18.2, 20.5, 19.9, 19.1, 9.8, 18.5, 17.3, 11.9, 13.4, 
    10.6, 10.5, 3.6, 2.8, 5.2, 4.7, 5, 6.5, 5.9, 6.3, 6.3, 6.1, 5.8, 4.5, 
    5.4, 7.5, 5.2, 5.3, 5.4, 4.8, 6.8, 5.7, 5.3, 5.8, 5.2, 3.7, 4.2, 4.7, 
    5.1, 6.1, 7.4, 7.2, 8.6, 9.1, 8.1, 8.4, 9.3, 11, 11.5, 12.1, 12.9, 14.8, 
    17, 18.5, 18.2, 20.1, 15.9, 22.5, 21.3, 19.3, 20.8, 22.1, 19.6, 16.4, 
    17.5, 16.7, 15.4, 14.9, 6.3, 10, 9.9, 12.7, 14.1, 10.8, 9.3, 10.7, 10.9, 
    11.1, 9.7, 10.8, 10, 6.5, 9.8, 10.2, 10.5, 11.1, 11.5, 14.1, 15.3, 15.1, 
    14.8, 15.2, 13.3, 14.9, 11.6, 10.8, 12.4, 10.8, 11.2, 10.3, 11.4, 10.7, 
    9.8, 10.9, 12.1, 14.4, 12.6, 13.2, 15.3, 16.3, 14.5, 15.1, 13.8, 15.8, 
    14.3, 15.7, 10.4, 13.7, 14.3, 17.2, 12.6, 10.4, 12.2, 11, 10.6, 9.5, 8.3, 
    11.1, 6.6, 4, 3.6, 8.6, 11, 6.1, 5.1, 8.4, 7.9, 8.3, 8.7, 8.3, 7.9, 5.1, 
    7, 7.8, 6.9, 7.1, 8.3, 9.8, 10.2, 6.1, 9.1, 9, 8.6, 8.8, 9.6, 2.8, 4.8, 
    4.7, 3.1, 0.8, 1.4, 1.3, 3.5, 2.1, 4.7, 5.6, 5.1, 5, 4.1, 3.9, 3.1, 3.5, 
    6.9, 4.2, 4.4, 4.1, 5.6, 5.1, 3.3, 4.3, 2.7, 1.5, 0.8, 1.1, 3.8, 6.1, 
    3.5, 2.3, 0.3, 0.5, 2.4, 7, 1.4, 0.4, 1.9, 5.4, 6.8, 6.3, 6, 6.3, 7.1, 
    6.7, 8, 8.7, 8.2, 6.5, 5.9, 5.9, 7.1, 6.8, 6.6, 6.9, 3.6, 3.2, 4.7, 4.1, 
    3.9, 5.9, 3.7, 1.6, 1.3, 4.6, 7.5, 3.6, 3.8, 2.9, 3.3, 2.9, 2.4, 5.2, 
    3.4, 2.5, 4.5, 3, 4.4, 7.6, 6.5, 5.2, 3.3, 3.1, 5, 5.1, 4.3, 4.4, 7, 6.1, 
    9.1, 7.8, 4.1, 4.5, 2.7, 3.6, 4.1, 4.5, 2.6, 3.6, 3.8, 4.1, 5.3, 6.1, 
    6.3, 6.5, 7.8, 4.8, 7.2, 7.5, 5.9, 8.6, 7.4, 5.2, 4.4, 6.7, 6.1, 4.7, 
    6.8, 3.2, 3.4, 3.3, 8.8, 8.2, 7.6, 4.4, 0.4, 0.5, 1.9, 3, 10.5, 11.8, 
    13.9, 14.4, 14.5, 1.7, 16.6, 12.3, 1, 2.3, 1.2, 1.8, 1.3, 1.7, 0.2, 10.9, 
    12.4, 13.3, 15.5, 12.8, 11.5, 0.4, 12.9, 11.7, 12.7, 12.7, 10.6, 10.4, 
    10.2, 10.7, 11.8, 12.4, 11.1, 11.4, 11.5, 9.4, 8, 10.5, 10.1, 10, 11.7, 
    10.7, 14.8, 14.4, 12.9, 9.6, 11.7, 11.2, 8.3, 8.9, 10.5, 9.6, 10.6, 11.2, 
    11.6, 12.1, 10.9, 10.4, 12, 12.8, 11.3, 13.6, 12.8, 14.1, 14.1, 15, 16, 
    16.2, 15.5, 16.1, 16.6, 14.7, 14.9, 16, 16, 15.9, 15.4, 8.5, 15.2, 3.3, 
    14, 15.9, 13.7, 15.6, 14.9, 14.3, 14.7, 17, 16.8, 17.7, 20.9, 17, 12.1, 
    12, 9.5, 7.7, 7, 7.4, 1.2, 7.7, 11.5, 9, 2.1, 2, 9.8, 10.1, 10.6, 10.5, 
    11.4, 10.3, 8.4, 8.8, 8.6, 9, 8.9, 8.6, 7.9, 8.8, 7.1, 8.2, 9.4, 8.5, 
    7.5, 9.1, 10.9, 11.2, 12.2, 11.9, 13.2, 12.1, 12.2, 11.1, 10.5, 10.7, 
    10.8, 9.9, 10.1, 12.4, 12.3, 13.7, 11.7, 10.1, 9.7, 8.4, 8.6, 11, 8.6, 
    7.3, 7.3, 8.9, 8.8, 8.5, 8.6, 9.3, 9, 9.5, 8, 9.3, 9.4, 8.9, 10.2, 9, 
    8.9, 8.7, 8.5, 7.3, 7.9, 7.3, 7.8, 7.2, 3.1, 6, 5.6, 3.7, 5.5, 6.2, 6, 6, 
    5.4, 6.1, 5.4, 6.2, 5.5, 4.9, 6.5, 3.9, 6.1, 6.1, 5.9, 6.1, 6, 6, 5.9, 
    4.4, 5.6, 6, 6.3, 5.8, 6, 7.2, 7.9, 7.7, 7, 7.8, 8.2, 5.5, 9.1, 8.3, 8.6, 
    8.1, 10, 9.2, 9.7, 9.5, 9.6, 7.9, 8.1, 7.5, 6.4, 7.6, 7.8, 7.6, 7.5, 7.9, 
    9.1, 9, 7.6, 7.2, 8.4, 7.8, 7.8, 7.4, 6.5, 7.5, 7.9, 5.2, 5.2, 8.2, 7, 
    4.9, 6.3, 5.4, 6.4, 5.6, 4.9, 5.1, 4.7, 6.5, 6, 4.1, 4.6, 5.5, 3.9, 3.5, 
    2.9, 2.7, 2.7, 1.5, 1.9, 1.4, 2.1, 1.7, 2.1, 4, 3.5, 2.9, 2.1, 0, 0.9, 
    1.5, 1.7, 2.9, 3.1, 4.2, 4.7, 3.8, 4.9, 4.6, 3.1, 8.8, 10.2, 11.9, 13.9, 
    12.9, 15.3, 16, 15.1, 12.4, 10.3, 9.4, 8.3, 11.1, 7.2, 5.8, 6.8, 5.2, 
    4.1, 5.7, 5.8, 3.9, 5, 5.5, 4.6, 8.5, 8.4, 7.6, 7.5, 6.2, 5.6, 5.8, 3.6, 
    2.4, 0.8, 1, 2.3, 2.6, 1.5, 6.3, 10, 8.1, 9, 5, 5.3, 1.8, 1.6, 3.5, 4.8, 
    4.2, 4.3, 7.7, 4.4, 4.5, 6, 6, 5.9, 5.9, 6.7, 2.8, 2.8, 3, 2.8, 2.6, 1.8, 
    2.1, 2.1, 3.4, 2.4, 1.4, 2.1, 1.3, 2.2, 2.2, 1.2, 1.9, 2.3, 1.8, 1.6, 
    2.1, 10.1, 11.3, 13.1, 12.8, 12.4, 11.4, 12.1, 11.4, 10, 10.2, 8.6, 8.7, 
    9.5, 9.9, 9.4, 2.8, 8.3, 7.5, 3.8, 3.1, 2.8, 4, 5.6, 13.6, 14.1, 14.5, 
    13.7, 13.7, 12.7, 13.7, 15.2, 12.5, 14.2, 13.4, 16.1, 16.3, 16.3, 13.7, 
    12.7, 14.4, 13.3, 15.4, 13.2, 12.1, 13.5, 10.3, 10.3, 8.7, 9.7, 8.7, 9.5, 
    9.8, 8.8, 8, 7.1, 6.5, 7.3, 6.1, 4.6, 2.2, 1.1, 6.5, 5, 7.9, 7.5, 6.7, 
    6.4, 7.4, 4.9, 8.1, 6.9, 5.7, 6.3, 2.4, 3.5, 4.6, 5.8, 6.9, 7.3, 7.3, 
    7.3, 7.3, 5.6, 5.4, 4.1, 2.5, 11.1, 11.9, 12.8, 16.5, 13.7, 12.2, 11, 
    10.7, 8.9, 12.3, 11.7, 11, 11.6, 12, 13.2, 14.1, 10.3, 7.3, 4.6, 5.9, 
    8.2, 0.8, 2.4, 4.2, 0.3, 6.1, 8.6, 9.8, 10.5, 10.7, 10.7, 12.7, 10.8, 
    10.9, 12, 10.4, 8.7, 7.9, 4.8, 13, 11.8, 13.4, 13.4, 11.1, 11.8, 9.4, 
    8.7, 6.9, 4.3, 3.5, 1.6, 1, 2.7, 4.3, 4.8, 5.9, 7.1, 4.7, 7.7, 8.2, 7.3, 
    8.8, 10.5, 10.7, 11.1, 11.1, 11.5, 12.8, 12, 10.9, 9.7, 8.3, 4.9, 11.2, 
    9.9, 10, 10.6, 11.1, 11.2, 9.7, 10.8, 10.8, 11, 8.8, 11, 12, 10.7, 12.3, 
    11.9, 10.3, 11.6, 12.1, 13.4, 12.9, 13.2, 10.6, 12.5, 12.1, 8.8, 10.3, 
    9.2, 9.9, 8, 9.1, 5.3, 7, 7.6, 9, 6.8, 5.5, 5.1, 5.8, 5.3, 4.7, 4.7, 4.3, 
    5.8, 5.3, 6.2, 7.5, 6, 7.4, 6.1, 4.8, 3.5, 4.1, 6, 5.7, 3.3, 6.7, 6.8, 
    10.2, 9, 7.8, 5.7, 8.4, 9, 9.1, 7.1, 6.2, 5.2, 5.3, 3.3, 4.4, 5.2, 8.3, 
    8.9, 8.9, 7.9, 6.9, 7.2, 6.6, 6.6, 4.8, 6.5, 8.9, 7.4, 10, 10.2, 9.5, 
    8.8, 10.4, 8, 6.3, 6.2, 8.3, 7.4, 6.9, 5.3, 5, 4.1, 3.1, 2.5, 3, 2.4, 
    1.8, 2.2, 1, 1.7, 2.4, 0.9, 2.3, 2.3, 2.2, 1.7, 1.7, 2.4, 5.8, 7.3, 7.6, 
    8.1, 9.9, 8.6, 8.5, 2.3, 8.9, 7.1, 3.4, 2.4, 1.5, 1.9, 1.3, 1.9, 2.2, 2, 
    1.9, 2.1, 2, 1.9, 0.8, 1.2, 1.5, 1.6, 2.5, 4.8, 4.8, 5.1, 3.5, 3.8, 5.7, 
    5.6, 6.1, 7.1, 6.7, 8.3, 8.3, 8.8, 9.2, 9.4, 9, 8.9, 5.6, 10.3, 8.1, 4.6, 
    3, 3, 4.9, 3.9, 4.5, 4.6, 1.5, 1.3, 1.9, 4, 0.6, 2.1, 1.1, 0.2, 0.5, 4.2, 
    0.7, 6.7, 2.6, 6, 6.8, 10.1, 2.4, 2.2, 5.9, 2.6, 3.1, 0.9, 0.2, 0.2, 1, 
    0.2, 2.7, 2.5, 1.2, 9.5, 8.6, 7.9, 8.7, 9.6, 9.3, 8.8, 8.1, 9, 8.8, 3.2, 
    8.7, 9.8, 10.1, 9.5, 9, 9.8, 9.8, 9.4, 8.7, 3, 8.5, 9.5, 8.9, 9, 8.6, 
    8.7, 8.7, 8.8, 8.3, 7.7, 7.7, 7.5, 8.1, 7.7, 7.2, 6.8, 7.2, 7.7, 7.2, 
    6.8, 6.7, 6.9, 7.7, 6.1, 3.8, 6, 5.2, 6.3, 4.4, 2.7, 1.5, 10.4, 10.2, 10, 
    10, 9.4, 12.4, 11.3, 10.8, 10.6, 11.7, 9, 9.9, 6, 7.8, 11.7, 11.5, 11.2, 
    8.4, 8.4, 6.6, 11.2, 12.2, 11.5, 11.7, 13.4, 7.1, 15.8, 13.9, 12.2, 8.9, 
    13.4, 11.7, 12.4, 13.8, 14.3, 11.5, 12.4, 14.5, 12, 12.8, 14.9, 10.8, 
    15.5, 12.2, 12.7, 12.7, 13.6, 10.9, 10.6, 12.9, 13.9, 14.7, 13.3, 12.9, 
    13.9, 13.4, 12.9, 11.9, 9.8, 11.4, 11.6, 13, 12.9, 11.9, 10.7, 11.4, 
    13.9, 14.6, 12.7, 13.1, 13.2, 13.4, 12.2, 11.3, 9.1, 8.7, 11.9, 7.9, 8.7, 
    11.4, 9.6, 8.1, 8.6, 10.6, 8.9, 8.4, 8, 3.7, 6.1, 7.3, 8.1, 8.6, 6.5, 
    6.5, 8.1, 0.9, 0.6, 1.7, 1.3, 0.2, 1.9, 1.4, 2.1, 2.4, 2.2, 2.5, 4, 7.4, 
    6.9, 4.8, 7.4, 6.8, 2.8, 5.6, 6.6, 7.1, 6.7, 8, 5.1, 8.8, 9.1, 4, 4.9, 
    4.7, 8.8, 10.7, 12, 14.2, 12, 17, 11.8, 14.2, 12.8, 15.2, 14, 9.7, 15, 
    14.6, 15.9, 15.7, 16.1, 15.4, 14.7, 11.2, 13.1, 14.1, 15.4, 13.9, 12.5, 
    12.3, 12.1, 12.3, 12.3, 10.6, 11.8, 11.9, 10.2, 9.5, 9.4, 8.9, 10.3, 
    11.2, 6, 6.5, 8.9, 5.4, 10.3, 1.8, 4.9, 2.3, 0.1, 1.7, 1.1, 3.3, 2.3, 
    1.5, 2.6, 3.5, 3.8, 8.6, 10.2, 2.1, 4.4, 3.3, 4.9, 4.3, 1.4, 11.3, 9.9, 
    10.7, 10.7, 13.7, 11.3, 9.3, 10.8, 15.4, 15, 10.3, 11.9, 7.7, 4.3, 7.4, 
    7, 9.1, 13.1, 10.9, 9.3, 10.4, 5.7, 9.3, 8.6, 9.3, 8.5, 10.5, 8.6, 7.1, 
    7.8, 6.1, 7.6, 6.3, 3.2, 8.1, 8.4, 7.7, 6.6, 6.2, 7, 4.9, 6.1, 3.8, 4.6, 
    7.4, 7.3, 8.1, 8.4, 8.8, 8, 9.5, 7.5, 5.7, 6.4, 7.9, 5.9, 6.3, 7, 7.7, 
    6.9, 8.1, 7.1, 6.4, 7, 6, 5.7, 6.3, 6.1, 6.5, 4.9, 6.8, 5.8, 4.8, 4.1, 
    4.6, 5.2, 3.4, 1.7, 1.4, 2.5, 1, 0.5, 0.1, 5.3, 5.7, 5.6, 5.1, 5, 5.8, 
    6.2, 6.2, 6.6, 6.3, 6.6, 3.8, 3.9, 7.4, 7.2, 7.2, 7.1, 7.2, 6.6, 6.1, 
    5.6, 6.5, 7.3, 6.6, 7.5, 7.7, 7.1, 6.6, 6.4, 7.2, 6.4, 6.7, 7.8, 9.4, 
    8.6, 8.7, 4.2, 9.7, 8.5, 5.6, 7.9, 6.6, 13.2, 15.7, 3.9, 4.5, 4.8, 16.4, 
    16.9, 6.6, 16.6, 15.2, 11.6, 9.9, 11.1, 8, 7.6, 8.4, 8.4, 7.9, 10, 10.3, 
    11, 9.3, 9.9, 8.6, 9.1, 9.6, 11, 11.3, 11.4, 11.3, 12, 11.6, 11.4, 13.2, 
    13.1, 12.2, 11.8, 10.7, 9.6, 9, 10.4, 11.6, 11.1, 10.2, 10.4, 10.5, 10.3, 
    9.5, 9.5, 6.9, 10.4, 10.1, 0.3, 2.2, 1.8, 8.4, 3.8, 10.9, 10.4, 9.3, 7.9, 
    8.8, 3.7, 10.4, 11, 12.8, 12.1, 6.2, 16.9, 12.3, 11.5, 14.3, 12.6, 7.8, 
    3.6, 6, 6.5, 4.5, 9.3, 9, 7.9, 9, 9.8, 9.1, 9.7, 8.5, 6.8, 5.4, 3, 1.7, 
    1.9, 0.8, 0.6, 2.1, 2.1, 2.2, 1, 1.1, 1, 1.9, 1.4, 1.9, 0.9, 1.4, 4.1, 
    1.5, 2.6, 2, 1.9, 0.3, 1.2, 1.2, 0.3, 0, 0, 0, 0, 0, 0, 0, 0, 5.8, 6.7, 
    5.9, 6.7, 6.7, 7.9, 7.5, 9.7, 10.8, 9.3, 9.7, 12, 14.9, 12.1, 13.7, 13, 
    8.8, 9, 6, 5.3, 5.1, 9.6, 10.3, 8.4, 6.5, 5.8, 10.7, 9.5, 10.2, 9.4, 9.4, 
    8.9, 7.9, 7.1, 8.7, 6.9, 7.6, 7.8, 7.5, 7.6, 9.2, 7.4, 8.4, 8.2, 10.7, 
    8.9, 8.2, 9.4, 11.8, 12.5, 8.9, 10.3, 10.4, 10.6, 10.4, 9.5, 8.4, 8.3, 
    8.5, 9.8, 10, 7.2, 7, 6.9, 5.7, 3.8, 4, 3.2, 4, 5.8, 5.2, 5.4, 6.6, 7.1, 
    9, 5.1, 6, 4.5, 6.5, 6, 4.9, 4.4, 3.6, 5.9, 4.7, 5.3, 2.3, 6.7, 3.8, 6.2, 
    6.3, 4.1, 4.8, 5.9, 6.8, 6.9, 8.2, 10.3, 5.9, 5.9, 9.8, 8, 14.1, 15.1, 
    14.9, 11.3, 7.8, 6.9, 6, 8.3, 5.3, 3.8, 0.6, 7.3, 4.5, 2.2, 12.9, 14.5, 
    5, 4.9, 3.7, 10.7, 11.6, 11.6, 11.5, 11, 9.2, 10.5, 13.1, 19.4, 20.5, 
    20.7, 19.2, 18.7, 19.4, 17.6, 17.1, 18.2, 18.2, 18.3, 18.2, 16.8, 16.7, 
    18.8, 18.7, 19, 16.9, 16.2, 16.3, 15.1, 16.6, 14, 13.2, 13.2, 13.8, 14.5, 
    15.9, 17.3, 18.5, 19.3, 18.7, 17.7, 18.3, 18, 18, 16.9, 16.2, 16.7, 15.4, 
    14.3, 13.6, 13.5, 13, 13.2, 12, 12.5, 12.5, 12.8, 14.5, 14.3, 14.4, 12.6, 
    12.4, 11.8, 9, 11.3, 10.9, 7.2, 5.7, 11.3, 11.2, 10.8, 5.1, 6.4, 5.9, 
    2.5, 2, 2.9, 6.4, 8.2, 8.2, 10.4, 10.2, 11.6, 12.7, 13.2, 13.7, 13.4, 
    13.2, 12.2, 11.7, 12, 12.2, 11.9, 11.2, 11.1, 9.6, 9.1, 9.2, 10.5, 6.4, 
    7.2, 7.5, 7, 9.1, 8.9, 9.6, 10.6, 13.4, 9.4, 0.7, 4.3, 2.2, 4.2, 1.9, 
    1.6, 0.6, 2, 4.3, 4.4, 6.7, 7.1, 11.9, 11, 11.5, 10, 13.8, 12.1, 10.2, 
    12.2, 11.8, 11.5, 13.6, 13.6, 16.2, 14.5, 14.5, 15.3, 15.5, 17, 15.8, 
    15.4, 12.2, 10.9, 9.7, 12.9, 13.8, 12.9, 12.2, 11.2, 11.6, 13.6, 15.2, 
    12.6, 12.7, 9.1, 8.5, 7.4, 9.1, 8.4, 8.3, 5.2, 8.6, 8, 6.2, 4.1, 7.6, 
    7.8, 7.3, 6.3, 9.5, 11, 10.1, 9.7, 11, 11.9, 14.8, 16.9, 3.1, 4.1, 2.5, 
    9.5, 7.1, 9, 0.6, 1, 4.1, 1.5, 1, 3.6, 2.6, 6, 5, 1.4, 4.2, 16.2, 10.1, 
    14.6, 13.8, 13.6, 10.2, 9.4, 13.9, 15.5, 14.3, 13.7, 7.5, 9, 8.9, 1.2, 
    8.8, 11.1, 8.9, 7.4, 6.4, 5.4, 6.6, 7.4, 6.7, 5.6, 8.2, 10, 7, 9.2, 8.6, 
    9.1, 7.1, 5.5, 7, 5.3, 15.9, 12.7, 10.9, 9.9, 9.7, 9.8, 12.4, 13.5, 14.7, 
    13.1, 10.6, 11.1, 10, 11.6, 14.5, 15.9, 13.7, 12, 10.6, 10, 11.4, 9.9, 
    10.7, 12.4, 11.6, 10.9, 13.3, 11.3, 11.2, 12.4, 11, 9.3, 9.3, 9.2, 12, 
    9.6, 9.8, 9.8, 8, 9.6, 7.5, 7, 7.9, 8.9, 9, 10.2, 9.6, 7.7, 3.8, 9.4, 9, 
    11.9, 13.6, 11.7, 8, 9.8, 9, 9.8, 10.3, 12.1, 12.9, 12.8, 15, 10.3, 10.4, 
    10.9, 9.6, 10.4, 10.6, 7.9, 8.1, 10, 11.8, 10.3, 8.2, 10.2, 8.7, 7.1, 10, 
    10.4, 7.9, 8.9, 8.8, 8.7, 7.2, 8.7, 8.6, 8.9, 9.8, 10.1, 8.5, 8.7, 9.8, 
    10.3, 9.9, 9.7, 9.1, 9.1, 10.6, 9.6, 9.7, 9.3, 9.4, 11.1, 10.2, 8.7, 
    11.1, 9.5, 8.8, 8.8, 9.7, 10.1, 11.1, 11.7, 10.9, 10.7, 10.2, 11.2, 11.6, 
    7, 9.7, 10.9, 11, 11.5, 11.2, 11.1, 11.3, 10.4, 11.2, 12.2, 13.1, 12.9, 
    12.9, 12.4, 12.4, 14.7, 12.2, 10.8, 13.7, 10.3, 10.5, 11.9, 12.8, 13.8, 
    12.9, 11.9, 14.1, 13.3, 10.1, 12.2, 12.3, 13.4, 11.3, 11.2, 11.3, 11.2, 
    13.5, 17.5, 7.7, 6.4, 8.1, 9.4, 7.2, 8.8, 9.4, 7.9, 8.4, 7.5, 7.2, 7.3, 
    7.7, 7, 5.6, 3.9, 6, 4.4, 3.5, 1.5, 0.4, 3, 3.8, 3.2, 4.4, 7.3, 6.8, 6.5, 
    6.2, 7.2, 7.6, 7, 6.7, 6.3, 6, 5.5, 5.1, 4.6, 4.3, 4.8, 4.3, 2.8, 1.8, 
    1.3, 0.6, 2.6, 2.4, 0.8, 0.9, 1.5, 1.8, 3.5, 2.6, 1.6, 0.3, 0.7, 0.7, 
    2.3, 4.3, 5.3, 6.5, 7.3, 7.2, 7.1, 5, 6.9, 6.7, 1.9, 0.5, 7.7, 2.9, 2.9, 
    4.7, 4.1, 6.8, 7, 6.6, 7.5, 8.7, 8.8, 9.2, 8.6, 9.7, 7.2, 7.3, 6, 5.4, 
    6.6, 5.9, 6.2, 4.4, 3.9, 4.8, 4.3, 1.7, 2.4, 2.1, 4.7, 4.1, 4.8, 7.1, 
    7.8, 8.8, 5.3, 6.9, 6.6, 7, 6, 4.7, 5.6, 4.7, 4.9, 5.3, 6.1, 5, 5.2, 3.7, 
    5.1, 5.8, 6.1, 5.2, 4.7, 6.1, 6.8, 6.5, 7.1, 6.8, 4.9, 5.4, 5.3, 7.1, 
    8.4, 8.2, 5.1, 5.7, 5.5, 6.4, 5.9, 4.8, 6.4, 6.3, 6.2, 7.3, 7.4, 9.2, 
    6.6, 6.1, 5.4, 9.5, 10.1, 7.7, 8.2, 7.1, 6.9, 7.1, 8.8, 9.5, 8.1, 10.1, 
    11, 12.4, 10.8, 8.2, 6.7, 6.7, 7.6, 8.5, 8.4, 9.6, 9.7, 9.3, 9.5, 8.5, 
    8.6, 8.5, 9, 7.5, 9, 8.2, 8.7, 4.6, 7.9, 4.4, 7.4, 6.9, 7.4, 6.6, 5.1, 
    6.1, 6.2, 6.8, 6.5, 5.9, 5.7, 6.5, 6.7, 5.4, 6.1, 5.9, 2.1, 1.7, 1, 0.7, 
    3.6, 2, 0.9, 0.4, 1.8, 3.4, 3.1, 4.3, 4.9, 5.9, 5.2, 5.1, 5, 4.2, 1.4, 0, 
    0, 1.1, 3.3, 3.3, 4.6, 4.5, 4.4, 5, 6.1, 4.3, 5.9, 3.8, 4.4, 2.8, 6.5, 5, 
    4.8, 5.9, 6, 5.8, 6.6, 6.4, 7.9, 9.1, 9.8, 10, 6.3, 11.3, 11.2, 12.3, 
    13.6, 14.4, 15.1, 15.2, 15.5, 17.4, 16.2, 17.9, 17.8, 20.2, 21.2, 20.1, 
    19.5, 18.3, 19, 19.4, 18.7, 21.4, 20.1, 19, 17.3, 18.7, 17, 17.8, 17.6, 
    17.6, 15.5, 16.2, 16.9, 16.9, 15.4, 15, 15.4, 16.5, 11.5, 11.4, 11.7, 12, 
    15.4, 14.9, 11.9, 11.9, 12.4, 10.8, 9.7, 9.6, 8.9, 9.5, 8.5, 10.5, 9.8, 
    8.8, 9.4, 10.5, 12.1, 11.1, 12.5, 7.8, 12.7, 10.7, 10.6, 11.3, 12.4, 
    12.6, 13.9, 14.9, 14.4, 14.6, 10.4, 14.1, 14.3, 13.7, 13.4, 12.6, 13.5, 
    12.6, 12.2, 12.7, 12.8, 12.8, 13.3, 12.8, 12.2, 12.9, 13.3, 12.4, 13.6, 
    13.1, 13.3, 12.8, 12.3, 12.3, 11.4, 12, 12.3, 11.3, 10.6, 11.7, 11.4, 
    10.3, 10.6, 9.2, 10.6, 10.2, 10.1, 9, 9, 9.8, 10, 9.1, 9.6, 9.8, 10.1, 
    10.4, 9.6, 9.5, 10.4, 9.4, 10.5, 10.3, 11.1, 10.8, 11.6, 11.7, 11.6, 
    11.2, 10.7, 9.9, 10.4, 12.6, 11.3, 11.9, 10.7, 10.7, 10.1, 7.9, 6.9, 7, 
    4.8, 2.9, 9.4, 9.8, 9.8, 9.8, 8.7, 9.1, 7.8, 6.7, 6.8, 7.7, 6.9, 4.7, 6, 
    7.9, 5.7, 10.5, 11.2, 10.6, 5.1, 3, 13.7, 11.9, 4.4, 1.7, 10.1, 14.4, 
    17.1, 17.6, 12.9, 10.6, 10, 10.4, 9.3, 10.2, 10.2, 10.1, 10.9, 13.3, 
    12.7, 13.7, 13.1, 14.6, 14.3, 12.6, 10.4, 7.7, 6.8, 6.7, 7, 7.5, 9.5, 9, 
    9.6, 10.2, 10.6, 5.8, 6.7, 8.1, 6.2, 7.9, 6.6, 6.4, 5.3, 5.3, 5.1, 3.4, 
    3.4, 3.9, 3.5, 2, 3.6, 5.1, 7.8, 7.1, 7.8, 8, 2.4, 8.8, 8.5, 6.9, 8.8, 8, 
    1.1, 6.7, 0.7, 5.5, 4.1, 3.3, 3.5, 4.5, 2.4, 0.6, 4.9, 7.1, 7.9, 7.9, 
    7.9, 9, 9.8, 9.2, 9.8, 9.2, 10.2, 9.4, 8.4, 9.6, 9.3, 8, 9.4, 8.5, 9.2, 
    9.6, 7.5, 9.2, 7.8, 8.1, 7.9, 7.3, 7.2, 7.9, 8.8, 8.3, 6.3, 6.4, 6.2, 
    6.3, 7.6, 7.8, 8.6, 8.7, 8.2, 7.9, 8.4, 8, 8.1, 7.7, 7.8, 7.4, 8.2, 6.9, 
    7.1, 7.3, 7.5, 7.3, 6.6, 6.2, 5.1, 7.3, 7.1, 6.4, 6.1, 6.1, 6.4, 6.6, 
    6.5, 6.4, 6.4, 6.1, 6.5, 6.4, 7.2, 6.9, 5.7, 5.4, 6.2, 5.8, 6.3, 5.3, 
    6.6, 6.2, 6.5, 2.8, 4.3, 2.2, 4.4, 3.6, 4, 3.6, 3.4, 5.4, 6.1, 6.3, 6.1, 
    7.3, 7.5, 4.9, 8.8, 6, 5.8, 5.6, 6.8, 7.6, 9, 5.7, 7.5, 6.9, 6.7, 7.9, 
    6.7, 6.8, 5.2, 4.4, 4.5, 3.7, 6.1, 5.7, 7.9, 7, 7.3, 6.3, 5.8, 5.5, 4.2, 
    4, 3.2, 2, 1.5, 1, 0.7, 1.2, 1.1, 4.1, 2, 1.6, 1.7, 4.7, 1.9, 1.9, 0.8, 
    0.6, 0.4, 0.5, 5.1, 3.9, 4.5, 5.5, 5.3, 6.1, 6.2, 5.8, 7.6, 8.8, 8.7, 
    8.2, 8.1, 8, 8, 8, 6.6, 6.4, 6.7, 6, 6.3, 7.2, 7.1, 5.8, 4.8, 4.1, 3.3, 
    1.5, 2.5, 1.4, 1.3, 0.7, 0.6, 2.9, 3.4, 3.7, 4.1, 5.3, 6.1, 5.1, 4.5, 
    4.4, 6.8, 5.7, 5.1, 5.5, 5.4, 6.6, 5.2, 5.5, 6, 3.8, 4.5, 4.3, 5.1, 3.9, 
    4.4, 6.2, 4.8, 6.7, 6.1, 6.3, 6.1, 5.9, 5.5, 4, 2.1, 4, 4.2, 5.5, 5.3, 6, 
    6.4, 9.3, 9, 8.6, 9.3, 8.8, 9.7, 8.4, 7.6, 6.7, 6.8, 5.3, 6.1, 9.2, 6.4, 
    6, 2, 3.6, 6.8, 3.6, 7.5, 5.6, 5.4, 6.5, 5.7, 4.4, 5.9, 5.1, 4.4, 4.7, 
    6.1, 6.3, 5.4, 7.2, 8.9, 7.3, 7.7, 5.4, 6.4, 6.9, 7, 6.7, 7.1, 7.3, 7.7, 
    7.8, 7.1, 7.1, 7.1, 7.4, 7.3, 6.5, 6.7, 6.9, 6.7, 6.9, 8.7, 8.3, 8, 8.5, 
    8.5, 7.3, 7.6, 7, 7.4, 8.1, 6.2, 6, 6.6, 5.3, 4.2, 4.6, 4.3, 3.2, 3.7, 
    3.2, 5.4, 3.8, 4.7, 3.4, 4, 3.5, 4.1, 3.3, 4.2, 3.7, 4, 5.1, 4.5, 5.6, 
    4.4, 4.5, 2, 3.4, 2.8, 2.4, 1.7, 0.8, 2.9, 0.8, 1.8, 1.3, 0, 2.4, 0.4, 
    3.1, 1.9, 3.5, 2.7, 2.7, 4.6, 5.5, 4.9, 4.6, 2.7, 0.5, 0.8, 1.3, 0.1, 
    2.8, 2.1, 3.2, 3.1, 2.6, 3.1, 1.5, 4, 3.6, 1.3, 2.8, 2.6, 1.1, 3.5, 0.4, 
    1.9, 3.4, 1.2, 0.8, 2.6, 2.8, 3.7, 2.1, 0.4, 1, 2, 1.4, 2.2, 2.4, 1.6, 
    1.6, 0.5, 1.6, 1, 2.9, 2.6, 2.1, 4.4, 2.9, 4.6, 3.2, 3.5, 4.5, 4.6, 3.7, 
    3.8, 3.8, 4, 8.5, 9.4, 10.3, 9.8, 10.3, 11.4, 11.5, 12.9, 11.1, 11.2, 
    11.2, 12.1, 12.3, 12.4, 12.5, 13.1, 13.2, 14, 15.5, 15.5, 14.1, 13.6, 
    13.7, 13.7, 14.6, 14.6, 14, 14.6, 15.1, 13.4, 14, 13.3, 13.5, 0, 1.3, 
    1.3, 1.5, 2.3, 4.3, 7.1, 7.1, 6.9, 7.9, 8.5, 11, 10.8, 12, 12.1, 13.9, 
    12.5, 12.8, 12.7, 12.7, 13.7, 11.2, 11.5, 9.7, 10.6, 10.2, 10.8, 8.6, 
    8.8, 7.6, 8.2, 5.8, 7.5, 6.4, 3.6, 1.6, 1.9, 1, 0.2, 0.8, 3.2, 3.6, 4.6, 
    6.5, 5.8, 6.2, 5.6, 6.4, 5.7, 5.3, 4.4, 3.7, 2.9, 2, 1.4, 1.6, 1.8, 2.3, 
    1.1, 0.7, 0.1, 6.4, 5.9, 6.3, 9.3, 10, 8.3, 7.4, 7.8, 7.9, 7.3, 6.9, 6, 
    4.9, 3.9, 2.9, 3.3, 3.3, 3.8, 4.6, 5.8, 5.5, 6.4, 5.4, 5.8, 4.2, 6.9, 
    5.2, 5.4, 6, 5.3, 6.4, 5, 6.6, 6.5, 5, 4.9, 5.9, 5.9, 4.6, 4, 4.4, 3, 
    2.6, 3.3, 0.8, 2.7, 1.1, 2.8, 2.4, 1.6, 3.2, 4.4, 4.8, 5.5, 6.7, 7.7, 
    7.7, 8.3, 8.1, 8.2, 8.4, 7.9, 8.3, 7.5, 7.1, 6.7, 6.4, 5.8, 5.9, 5.4, 
    4.1, 5, 5.3, 5.7, 7.8, 8.4, 8.9, 10, 9.9, 10.7, 8.8, 9.7, 9.2, 9.2, 10.3, 
    4.5, 5.6, 5.5, 8.2, 9.3, 10, 11.5, 10.8, 13.4, 14.9, 14.9, 11.3, 12.8, 
    13.1, 12.6, 10.6, 11.3, 10, 11.2, 11.8, 13, 10.3, 13.2, 11.3, 10, 12, 11, 
    11.4, 9.3, 10.2, 11.6, 13.2, 13.1, 10.5, 10.5, 11.2, 12, 11.7, 11.3, 
    10.6, 7.5, 9.2, 8.6, 10.5, 8.5, 7.7, 7, 9.5, 8.4, 8.1, 8.2, 13.1, 7.6, 
    7.5, 9.1, 6.9, 7.4, 6.1, 6.9, 6.2, 4.5, 5.5, 4.8, 4.9, 4.5, 4.3, 3.8, 
    3.9, 4.2, 3.9, 3.7, 4.8, 5.4, 4.7, 3.8, 4, 0.7, 2, 1.9, 2.9, 3.3, 5.3, 
    6.8, 6.8, 6.7, 6, 5.4, 6.8, 6.1, 5.9, 7.1, 6.8, 5.1, 5.7, 6.7, 5, 5.2, 
    5.7, 3.6, 3.2, 2.7, 1.6, 1.6, 3.9, 4.2, 4.2, 6.8, 6.9, 10.1, 8.5, 8.5, 
    8.2, 9.8, 9.6, 9, 7, 6.3, 7.8, 9, 8.6, 6.2, 1.3, 3.7, 1.4, 1.2, 1.9, 3.8, 
    7, 6.9, 4.7, 6.2, 6.3, 8, 7.8, 7.1, 6.5, 6.8, 7.2, 8.1, 7.6, 7, 7.3, 6.5, 
    6.4, 3.8, 4.9, 3.1, 2.3, 2.1, 2.2, 3.5, 3, 3.5, 4.2, 5.9, 3.9, 4.4, 4.6, 
    0.8, 0.9, 1.8, 1.8, 2.5, 3.5, 1.8, 2.7, 1.7, 3.1, 2.9, 3.6, 3, 2.5, 2.2, 
    1.3, 0.6, 0.5, 1.3, 4, 5.9, 7.6, 6.3, 5.6, 5, 4.2, 4.8, 4.9, 5.6, 5.2, 
    3.5, 3.8, 3.9, 2.2, 0.2, 3.2, 6.1, 5.7, 5, 4.9, 5, 4.4, 4.7, 4.7, 5.4, 
    5.9, 5.9, 6.6, 7.4, 8.3, 7.9, 6.1, 8.1, 7.9, 8.6, 9, 9.9, 9.9, 9.9, 11, 
    7.7, 10.3, 10.9, 11.4, 13, 13.2, 13.3, 14.4, 13.2, 14.1, 15.4, 18.3, 
    16.7, 13.5, 15, 15.8, 16.3, 15.8, 15.7, 14.9, 15.8, 11.1, 16.3, 15.1, 16, 
    15.5, 15.2, 14.3, 15.6, 15.6, 15.3, 16.5, 13.8, 14.8, 11.5, 8.2, 5.5, 2, 
    5.9, 5.2, 0.5, 3.2, 5, 7.4, 8.4, 8.1, 6, 7, 4.7, 2.9, 0.5, 2.6, 0.8, 3, 
    4.3, 5.9, 8, 9.7, 8.9, 10.3, 10.4, 10.3, 11.3, 8.1, 6, 4.5, 2.2, 3.3, 
    6.6, 6, 2.2, 1.6, 1.5, 6.8, 7.5, 6.8, 6.7, 4, 2.8, 3.3, 2.5, 1.9, 3.6, 
    0.2, 0.9, 2, 2.2, 0.6, 0.1, 1.4, 1.8, 1.2, 1.2, 4.6, 7.7, 3.8, 3, 3.1, 
    4.2, 5.2, 7.2, 6.7, 5.9, 8.4, 8.4, 8.6, 8.2, 5.3, 4.9, 6.9, 12.1, 14.3, 
    15, 14.9, 14.3, 13.4, 13.5, 12.7, 12.7, 10.5, 10.9, 11.1, 10.4, 9.1, 8.9, 
    10.2, 10.7, 9.7, 12.7, 12.2, 10.8, 10.1, 10.9, 8.7, 7.9, 6.3, 5.3, 2.7, 
    2, 2.9, 0.7, 1.5, 5.1, 4.2, 3.7, 2.7, 4, 6.1, 5.6, 4.1, 4.7, 4.4, 4.5, 
    2.9, 4.1, 3.3, 4.4, 5.8, 3.3, 1.9, 1.9, 3.2, 3.7, 6.5, 13.1, 13.9, 13.4, 
    11.6, 9.9, 8.6, 11.4, 12.2, 12.8, 12.7, 10.9, 8.6, 7.1, 8.1, 8.1, 8, 7.9, 
    7.9, 7, 9, 8.5, 9.9, 10.4, 9.9, 10.9, 11.2, 10.5, 12.2, 11.3, 11.3, 12, 
    15.6, 16.2, 15.8, 17.2, 10.9, 11.7, 13.8, 14.1, 14.8, 14.7, 10.8, 10.3, 
    10.2, 11, 11, 10.2, 11.9, 8.4, 6.6, 6, 6.8, 9.3, 4.8, 6.7, 8, 6.6, 8.1, 
    7.5, 9.7, 10, 8.3, 10.7, 9.4, 10.4, 11, 12.3, 10.8, 11.7, 12.4, 10.8, 
    10.1, 9.8, 7.6, 9, 9.6, 10.1, 6.8, 10.7, 10.8, 11.6, 10.7, 9.7, 9, 9.5, 
    9.2, 7.1, 10.4, 8.6, 7.7, 7.2, 7.1, 8.4, 7.9, 7.3, 8.1, 6.1, 5.7, 7.2, 
    5.2, 7.3, 9.3, 7.3, 4.8, 2, 5, 6.2, 9.4, 12, 12.1, 10.8, 11, 9.5, 8.9, 
    9.3, 11.1, 8.8, 7, 7.7, 9.7, 9.4, 9.4, 9.7, 10.2, 9.9, 9.7, 12, 10.6, 
    10.9, 11.4, 11.5, 11.7, 9.1, 8.8, 9.4, 7.3, 7.4, 8.2, 9.1, 7.8, 7.2, 9.3, 
    8.3, 6.1, 8.6, 7.8, 9, 9.4, 7, 8.8, 6.7, 8.4, 8.4, 8.5, 7.5, 8.2, 8.2, 9, 
    8, 6.7, 6, 7.5, 6.3, 9, 8.7, 8.5, 7.1, 6.5, 6.5, 6.2, 4.2, 3.4, 3.7, 4, 
    4.8, 5.4, 6.7, 7.2, 6.3, 6.8, 5.5, 3.1, 2.3, 2.2, 1, 2.2, 2.3, 2.7, 1.8, 
    1.5, 2.9, 3, 2.9, 2.5, 3.5, 3.8, 3.2, 2.4, 2.2, 0.4, 0.5, 0.3, 0.5, 4.2, 
    2.9, 2.8, 3.1, 2.6, 2.1, 1.7, 0.9, 0.6, 0.7, 1, 0.7, 0.7, 1.8, 2.6, 1.9, 
    0.9, 5.8, 7.9, 7.9, 4.6, 4.1, 4.1, 4.4, 1.2, 0.4, 3.4, 0.8, 0, 1.2, 3.4, 
    2.9, 2.4, 1.5, 0.4, 1.2, 0.7, 0.6, 0.6, 1.3, 1.3, 3.7, 4.5, 8.2, 8, 8.3, 
    8.1, 7.7, 8.3, 7.9, 6.9, 8.3, 8, 6.9, 5.5, 5.2, 6.2, 6.4, 7.7, 7.2, 6.4, 
    7.1, 6, 5.3, 5.3, 5.4, 5.9, 5.8, 5.7, 4.7, 4.9, 5.2, 6.2, 4.1, 4.3, 3.8, 
    4.5, 6.3, 5.8, 7, 9.4, 7.8, 9.1, 9.4, 8.5, 10, 6.6, 0.9, 0.6, 4.4, 1.4, 
    4.3, 1.7, 2.4, 2.2, 1.4, 0.7, 1.2, 1.2, 2.3, 0.9, 7.7, 4.9, 4.6, 5.2, 
    3.7, 4.9, 6.2, 5.5, 7.6, 8.5, 8.9, 9.8, 11.3, 10.8, 9.5, 13.2, 17.5, 
    17.7, 18.3, 17.5, 15.5, 16.1, 14.7, 12.6, 12.6, 8.7, 6.1, 4.9, 5.4, 5.2, 
    4.8, 4.4, 2.2, 0.9, 2, 4, 5.4, 2.7, 0.4, 1.8, 3.3, 5.3, 5.6, 7.9, 5.8, 
    7.4, 7.1, 9.3, 11.5, 12.5, 12.8, 11, 13.1, 14.4, 15.5, 12.8, 10.7, 9.6, 
    14.3, 14, 13.5, 13.1, 12.1, 8, 7.5, 8.8, 9.6, 6.7, 4.8, 4.8, 2.5, 2.7, 
    3.7, 2.6, 2.7, 1.6, 1.9, 3.5, 4.2, 7, 8.6, 8.6, 7.2, 6.4, 8.4, 7.8, 6.9, 
    7, 7.3, 6.7, 5.8, 4.2, 3.9, 3.7, 2.8, 2.9, 3.2, 4, 4, 3.5, 3.5, 3, 2.8, 
    2.8, 2.5, 2.6, 2.2, 2.9, 1.8, 3.3, 3.8, 3.3, 5.7, 6.9, 6.4, 4.9, 3.3, 
    5.4, 6.1, 6, 5, 5.2, 6.3, 6.1, 5.9, 7.2, 7.4, 6.9, 6.1, 5.5, 5.2, 4.5, 
    0.9, 0, 3.1, 1.4, 3, 7.7, 8.3, 6.3, 8.9, 10.1, 8.6, 6.6, 4, 3.6, 6.2, 
    5.4, 10.5, 2.1, 0.8, 0.8, 0.3, 1.7, 2.9, 3, 2.4, 2.2, 3, 7, 7.3, 7, 7, 
    6.3, 7.8, 8.4, 7.3, 8.3, 9.8, 12.5, 13, 3.5, 6.8, 6.3, 4.2, 1.9, 2.6, 
    3.3, 1.7, 1.1, 0.7, 2, 1, 3.2, 6.1, 6.5, 8.1, 8.1, 8, 9.6, 8.2, 7.9, 9.1, 
    10.3, 9.7, 10.5, 10.4, 12, 8.6, 12.4, 12.6, 13.7, 11.5, 9.9, 9.6, 9.8, 
    8.1, 4.5, 9.5, 5.4, 5.4, 3.3, 5.2, 5.1, 3.5, 1.5, 2.4, 3.6, 0.7, 2, 5.2, 
    4.2, 5.7, 5.9, 6.9, 7, 7.9, 9.4, 5.3, 5.6, 7.9, 8.2, 8.6, 8.6, 7.1, 5.9, 
    2.9, 0.6, 0.4, 2.4, 4.3, 6.2, 3.1, 1.4, 4.1, 4.3, 3.5, 3.6, 4.5, 3.9, 
    3.7, 3.9, 0.8, 1.2, 1.1, 0, 0.4, 0.6, 2.2, 1.7, 0.8, 4.8, 6, 10.4, 9, 
    5.6, 9.2, 10.9, 10.6, 2.5, 10.9, 9.2, 10, 9.5, 8, 0.8, 2.1, 2.7, 1.5, 
    1.5, 2, 3.6, 8.5, 9.3, 10.8, 6.8, 8.9, 6.5, 6, 6, 19, 22.4, 19.6, 20.2, 
    17.2, 15.6, 17.4, 15.5, 15.5, 14.2, 12.3, 14.1, 13, 10.4, 10.9, 11.7, 
    11.1, 10.1, 8.7, 10, 10.7, 10.8, 10.4, 10.8, 11.7, 10.4, 10.8, 9.7, 8.7, 
    9.9, 8.7, 9.9, 4.3, 7.8, 9.5, 8.5, 8.6, 7.2, 6.5, 6.5, 6.5, 7, 6.3, 7.4, 
    6.9, 10.9, 12.1, 12.4, 10.6, 10.3, 9.2, 9.8, 8.6, 10.7, 12.9, 11.3, 9.2, 
    7.7, 9, 6.4, 8.8, 7.3, 6.5, 9, 8.4, 8.6, 8.4, 9.6, 10.2, 10.7, 10.4, 
    10.2, 8.9, 10.5, 11, 12.4, 12.7, 12.3, 11.2, 9.9, 9.3, 9.6, 10.9, 8.7, 
    8.5, 8.8, 9.5, 10.8, 7.7, 8.9, 6.9, 7.4, 7.4, 7.5, 7.1, 6.7, 5.7, 4.8, 
    7.6, 6.5, 7.8, 8.2, 1.9, 1.3, 0.9, 2, 0.6, 0.9, 2, 1.6, 1.1, 2, 2.3, 2.4, 
    3.4, 2.4, 3.4, 3.1, 1.8, 2.4, 2.9, 2.7, 2.4, 2, 0.8, 0.5, 2.2, 1.3, 1.3, 
    0.9, 0, 4, 5.5, 5, 4, 6.7, 5.8, 5.8, 6.2, 8.7, 7.7, 9.2, 9.4, 11, 12.7, 
    12.8, 7.2, 9.9, 11.1, 11.3, 12.2, 13.2, 13.3, 9.8, 4.9, 0.7, 1.8, 4.2, 
    3.3, 4.9, 5.1, 3.6, 3.9, 5.6, 5.5, 6.9, 5.7, 4.3, 6.9, 8, 8.9, 7.1, 7.3, 
    4.7, 5.1, 5.6, 6.2, 5, 4.2, 5, 3.8, 3.4, 3.6, 2, 3.3, 3.8, 5, 4.9, 5, 
    4.4, 4.8, 5.3, 6, 6.4, 6.9, 6, 6.2, 7.4, 8.3, 7.4, 6.8, 6.8, 8.5, 8.6, 
    10.8, 9.4, 7.4, 9.2, 8.4, 9.3, 9.5, 9.3, 10.1, 9.9, 10.6, 9.3, 9.6, 10, 
    11.3, 10.5, 10.7, 11.4, 10.2, 11.9, 9.9, 10.8, 10.5, 9.2, 9.3, 7.9, 5.3, 
    7, 7.1, 6.5, 4.5, 4.1, 2.6, 8, 10.1, 5.9, 8.9, 12.3, 12.8, 13.9, 11.8, 
    11.7, 12.8, 10, 12.1, 11.3, 13.6, 10.1, 11.2, 9.4, 7.7, 5.7, 6.4, 7.1, 
    7.5, 5.6, 6.2, 8.2, 5.2, 7.3, 7.6, 3.4, 4.4, 4.4, 6.6, 4.8, 4.7, 3, 4.8, 
    5.8, 4.2, 2.8, 5.5, 4.2, 3.4, 4.9, 3.9, 4.8, 5.9, 5.9, 7.6, 5.6, 5.9, 
    5.4, 5.4, 5.4, 4.6, 4.8, 6.4, 5.6, 6, 6.1, 5.5, 4.2, 4.3, 4.2, 3.6, 2.6, 
    2.7, 1.7, 2.7, 2.8, 1.3, 2.1, 3.2, 3, 2.6, 2.7, 2.1, 1.6, 3.3, 2.1, 1.4, 
    3.6, 5.3, 6.1, 5.6, 3.6, 5.9, 2.9, 2.9, 1.7, 1.8, 2.8, 1.6, 0.5, 0.9, 
    2.1, 1.3, 2.6, 2.2, 1, 2.2, 2.1, 1.7, 0.9, 2.3, 0.6, 0.3, 2, 4.2, 3.2, 
    2.7, 0.2, 2.4, 2.5, 2.5, 2.7, 2.5, 0.9, 0.8, 0.8, 1.2, 4.9, 5.3, 1.7, 
    1.7, 2, 1.1, 2.2, 1.5, 7.3, 8.3, 9.2, 10.3, 9.2, 10.4, 13.2, 14.3, 4.5, 
    4.6, 15.9, 17.6, 15.1, 15, 12.3, 19.3, 17.3, 21.8, 23.7, 26.3, 24.9, 
    24.2, 22.5, 22.1, 23.9, 23.3, 22.5, 20.8, 18.7, 17.5, 18.3, 14.3, 13.3, 
    12.8, 10.3, 12.9, 15.2, 15.8, 16.9, 15.8, 16.3, 16.1, 15, 13.1, 11.3, 
    9.8, 8.8, 8.6, 9.6, 10.8, 11.6, 11.4, 8.8, 7.8, 9.2, 9.9, 9.3, 9, 9.9, 
    9.8, 9.5, 9.1, 9.3, 9.2, 10.6, 10.1, 10.6, 10.5, 9.1, 9.6, 10.7, 10.4, 
    8.8, 9.6, 7.9, 7.4, 5.3, 7.2, 6.6, 6.8, 6, 5.4, 5.8, 6.9, 3.7, 3.2, 1.7, 
    3.6, 2.7, 4.1, 6.5, 5.7, 5.8, 3.7, 3.6, 3.4, 3.7, 2.6, 2.5, 1.5, 1.4, 
    0.2, 0, 0, 1.8, 0.1, 1.7, 2.5, 0.6, 1.2, 2.6, 2.2, 1.1, 0.7, 0.8, 0.4, 
    0.2, 0.9, 1, 1.8, 1.6, 1.5, 1.3, 1.3, 2.7, 2.6, 3.7, 3.9, 4, 3.2, 3.3, 
    3.4, 3.8, 4.7, 4.8, 5, 4.5, 4.8, 3.8, 4, 4.3, 4.6, 4.3, 6, 3.8, 3.4, 2.3, 
    2.4, 2, 1.5, 1.4, 1, 2.2, 1.3, 2.7, 0.4, 0.9, 2.2, 2, 2.6, 2.8, 2.2, 2.6, 
    2.7, 2.1, 1.5, 1.3, 0.7, 2.6, 2.5, 3.2, 5.3, 6.2, 6.1, 7, 7.2, 6.4, 5.4, 
    5.1, 6.3, 5.9, 6.1, 6.2, 5.8, 5.8, 6.1, 7.2, 6, 6, 5.9, 6.2, 6.5, 6.6, 
    6.9, 5.8, 5.6, 4.9, 4.5, 3.8, 5.7, 5.8, 6.2, 4.9, 5.5, 4.8, 3.3, 6.7, 
    4.3, 3.9, 2.7, 3.9, 4.7, 4.6, 4.3, 3.9, 2.9, 3.4, 3.8, 3.9, 2.3, 4.3, 
    5.5, 6.8, 7.5, 7, 6.8, 6.6, 7, 7.7, 7.8, 6, 4.3, 5.2, 4.2, 3.6, 1.4, 1.9, 
    1.5, 3.8, 3.7, 4.6, 2.1, 0.8, 1, 2.5, 2.1, 5.9, 6, 6.3, 7.2, 7.5, 5.6, 
    6.5, 6.4, 6.8, 6.3, 4.9, 5, 5.8, 5.2, 4.4, 6.2, 7.2, 5.6, 6, 5.4, 4.6, 
    4.2, 4.8, 7.1, 5.5, 5.9, 6.3, 7.2, 7.4, 6.2, 5.8, 6.4, 6.5, 6.7, 6.1, 
    7.5, 8.8, 9.4, 8.6, 9.7, 9.1, 8.2, 8.3, 4.6, 2.2, 1.5, 2.8, 3.2, 4.4, 
    5.9, 6.4, 4.7, 6.8, 6.7, 7.1, 8.8, 9.4, 11.1, 9.7, 8.3, 9.3, 8.2, 10.6, 
    10.6, 10.4, 11.3, 13, 12.6, 9.2, 13.3, 14.5, 9.1, 11.1, 8.8, 9.3, 8.8, 
    9.9, 11.7, 9.6, 9.7, 10, 6.8, 6.9, 6.8, 6.1, 5.9, 4.3, 3.8, 3.1, 2.3, 
    0.8, 1.7, 3.4, 3.1, 2.1, 4, 3.6, 3.4, 3.4, 5, 5.9, 6.7, 6.8, 7.5, 6.8, 
    6.5, 6.1, 6, 6.8, 7.2, 6.7, 6.2, 5.8, 6.1, 5.5, 5.3, 4.8, 5.9, 4.5, 5.2, 
    4, 4.1, 4.2, 4.7, 5, 4.4, 3.2, 2.9, 3.1, 3.4, 3.6, 3.9, 2.6, 0.1, 2.2, 
    2.3, 1.7, 1.8, 2.7, 3.7, 4, 3.8, 2.7, 2.1, 2, 2.3, 2.7, 2.6, 2.6, 3.2, 
    1.1, 1.5, 0.9, 1.7, 0.9, 1.6, 0.3, 2.1, 0.9, 1.3, 1.9, 2.1, 3, 3.9, 3.4, 
    2, 3.4, 5, 6.2, 2.8, 1.7, 1.8, 0.2, 1.5, 0, 0.7, 1, 2.6, 2.1, 4.1, 4, 
    5.9, 6.3, 5.4, 6.8, 7.1, 7.1, 7.1, 6.9, 6.6, 7.1, 7.1, 7.4, 5.9, 6.2, 
    6.7, 6.6, 6.5, 6.2, 7.1, 7, 6.5, 5.8, 7.4, 7.4, 7.7, 8.1, 8.4, 7.8, 8.5, 
    9.1, 8, 8, 8.1, 7.6, 6.1, 0.5, 2, 2.2, 6, 6, 6.1, 8.3, 10.3, 11.2, 7, 
    8.5, 8.7, 9.1, 10.6, 9.3, 9.6, 8.7, 6.7, 6.2, 5.8, 6.8, 6.7, 3.8, 5.3, 5, 
    5.8, 5.6, 7, 4.1, 4.2, 4.6, 5.6, 5.9, 6.3, 5.8, 5.8, 7.1, 5.9, 6.6, 6.6, 
    6.4, 6.2, 7.5, 7.5, 7.3, 7.1, 7.6, 8.7, 6.7, 6.2, 2.5, 0.9, 2.3, 3.2, 
    5.1, 4.9, 4.8, 7.1, 6, 5.9, 5.1, 6.6, 4.9, 5.9, 6.5, 8, 8.7, 9.2, 8, 9.7, 
    9.6, 9.5, 9.4, 9, 8.4, 9.3, 9.8, 8.5, 8.7, 9.1, 8.5, 5.1, 8.2, 7.8, 10.3, 
    9.7, 11.5, 11.2, 9.8, 6.5, 6.5, 5.1, 5, 4.1, 4.8, 5.2, 5.9, 5.5, 4.7, 
    3.3, 1.6, 2.1, 4.5, 5, 4.6, 2, 3.7, 2.9, 1.9, 5.3, 5.6, 5.2, 5.6, 3.5, 
    5.1, 3.9, 4.5, 4.6, 6.9, 5.5, 2.7, 3.1, 4, 6.9, 7.6, 6.8, 6.6, 4.9, 4.7, 
    3.3, 2.4, 2, 0.8, 1.7, 0.8, 2, 4.2, 3.4, 4, 4.3, 5.9, 7.2, 7.5, 9.3, 
    11.3, 12.6, 11.9, 12.9, 12.7, 12.2, 12.3, 13.6, 12.1, 11.5, 11.1, 10.9, 
    9.8, 9, 7.2, 5.4, 4.2, 2.1, 0.9, 2.9, 7.9, 9.2, 10.1, 10.9, 11.1, 10, 
    9.7, 8.6, 8.6, 6.3, 6.2, 5.5, 4.6, 2.6, 2.8, 2, 1.2, 2.5, 3.9, 3.1, 4.2, 
    4, 4.8, 5.9, 6.1, 6, 7.3, 7.2, 8.8, 8.1, 8.8, 9.5, 8.8, 9.1, 9.2, 7.8, 
    8.8, 7.7, 9, 7, 7.9, 7.7, 8.2, 8.4, 7.4, 8, 6.7, 4.9, 7.4, 8.6, 9.2, 8.5, 
    7.8, 7.9, 8.8, 8.6, 8.3, 8, 7.7, 7, 7.7, 7.3, 7.2, 7.3, 6.3, 7.4, 7.3, 
    7.7, 6.4, 6.7, 7, 7.8, 8.2, 7.1, 8.2, 8.9, 8.4, 8.3, 9.2, 9.1, 8, 9, 9, 
    9.3, 9.2, 10.5, 10.6, 8.6, 9, 9.2, 9.7, 10.4, 9.7, 10.4, 10.4, 11.2, 
    12.8, 13.6, 15.7, 16, 16.2, 16.4, 16, 16.3, 16, 15.2, 14, 14.1, 14.7, 
    15.1, 15.6, 16, 14.6, 14.6, 14.4, 13.5, 15, 15.4, 16.7, 15.5, 13.8, 15.3, 
    14.1, 13.5, 13.8, 13.4, 12.4, 12.5, 8.7, 13.1, 14.7, 13.1, 12.6, 15.6, 
    16.5, 15.5, 16, 16.1, 14.6, 13.8, 13.4, 14.3, 13.5, 14.8, 14.2, 14.3, 
    16.6, 15.1, 13.2, 10.9, 10.6, 9.1, 8.7, 11, 10.2, 9.7, 10.2, 7, 10.3, 
    10.3, 9.7, 9.9, 8, 9.7, 8.6, 7.8, 6.7, 6.7, 7.6, 9.2, 8.2, 8.8, 10.1, 
    10.7, 8.8, 9.5, 9.4, 9.8, 5.7, 5.9, 4, 2.6, 3.6, 3.9, 5, 5.5, 4.8, 4.1, 
    4.6, 3.7, 3, 2.6, 5.3, 4.6, 3.8, 3.9, 7.2, 8.7, 9.1, 9.1, 8.9, 8, 7, 1.6, 
    0.7, 5.7, 2.7, 2.3, 4.6, 4.5, 4.9, 6.6, 4.7, 5.9, 6.2, 6.9, 5.4, 6.4, 
    6.1, 5.7, 3.7, 3.3, 2.8, 4.7, 3.8, 3.5, 2.4, 1.6, 0.8, 1.3, 2.4, 0.3, 
    1.6, 2.1, 2.4, 2.5, 1.7, 0.4, 1.2, 1.1, 2.7, 5.3, 4.5, 2.2, 2.2, 4.4, 
    3.8, 0.2, 0, 0.2, 0.7, 0.6, 0.7, 1.7, 2.7, 2.5, 2.7, 3.4, 4.3, 5.5, 5.3, 
    6.8, 8.1, 9.4, 9.1, 7.8, 7.9, 7.1, 8.8, 8.7, 9.7, 10.4, 13.3, 12.4, 12.9, 
    12.8, 12.9, 12.3, 13.9, 14.7, 13.5, 15.6, 15.3, 14.7, 14.3, 14, 14, 14.5, 
    14, 10.6, 12.7, 13.4, 13.5, 13.3, 13, 14.9, 13.9, 14.4, 13.8, 14.8, 12.7, 
    13, 12.4, 11.5, 12.4, 13, 13.9, 15, 13.9, 14.2, 12.5, 11.6, 11.6, 11.5, 
    11.9, 11.7, 12.1, 12, 12.5, 13.8, 15.3, 16.1, 16.3, 16.4, 17.2, 16.3, 
    15.6, 14.9, 14.9, 16.2, 15.6, 13.7, 12.5, 10.9, 10.4, 10.6, 10.2, 10.1, 
    11.5, 11.8, 11.9, 13.1, 12.8, 12.7, 14, 15.1, 15, 15, 12.5, 10.1, 10.4, 
    14.4, 18.9, 16.1, 16.6, 16.2, 18.5, 16.9, 14.9, 15.2, 19.1, 13.8, 17.2, 
    16.7, 15.5, 16, 14.1, 14.3, 13.1, 12.7, 11.1, 12.7, 13.4, 10.4, 11.8, 
    11.3, 13.4, 12.3, 9.9, 9.8, 7.5, 9.8, 9.7, 6.7, 6.5, 6.5, 6.4, 6.5, 5.7, 
    7.7, 8.2, 10, 11.3, 10, 9.4, 8.9, 9.8, 10.5, 9.3, 8.7, 8.4, 9.3, 9.9, 
    8.8, 9, 9.5, 10.1, 10.8, 10.9, 10, 6.8, 7.1, 7.6, 8.4, 8.4, 8.7, 8.5, 
    8.8, 9.2, 10.2, 10.3, 8.8, 8, 6.3, 4.4, 5.8, 5.4, 6.1, 8.1, 7.1, 8.5, 
    7.8, 9.5, 9.8, 8.6, 7.8, 7.5, 6, 5.6, 4.6, 4.4, 3.6, 5, 5.4, 5.2, 3.9, 
    3.9, 4.6, 3.5, 4, 4.4, 4.3, 3.9, 2.4, 2.7, 1.4, 1.5, 0.7, 0.3, 0.6, 0.7, 
    1.8, 2.4, 1.2, 1.2, 3, 1.6, 3.7, 3.3, 4.3, 3.2, 3.7, 2.8, 3.6, 3.9, 5.2, 
    3.1, 5.2, 3.8, 3.9, 4.7, 4.7, 5.3, 4.8, 5.1, 7.5, 6.9, 7.2, 7.5, 7.6, 
    6.8, 7.4, 7, 7.2, 8.2, 8.4, 9.1, 9.3, 10.2, 9.9, 8.4, 7.5, 5.8, 7.2, 7.6, 
    7.6, 8.2, 8.8, 8.5, 8.6, 8.9, 9.5, 5.7, 8.8, 7.7, 10.1, 7.4, 7.4, 6.4, 8, 
    8.7, 9.2, 8.7, 8.7, 8.7, 9.3, 7.7, 6.2, 5, 5.8, 5.8, 5.2, 4.5, 5.1, 4.6, 
    4.3, 4.5, 3.9, 4, 3.2, 3.3, 3.7, 3.2, 2.3, 2.2, 3, 3.5, 4.6, 3.9, 3.9, 
    2.8, 2.5, 1.3, 2, 1.7, 2.5, 2.1, 3.7, 3.7, 4.3, 3.7, 4.8, 5.9, 5.9, 7.1, 
    7.5, 8.3, 5.3, 2.3, 1.8, 2.7, 6.9, 7.6, 8, 8.6, 8.8, 7.7, 5.9, 4.1, 1.9, 
    1.3, 2.8, 3.6, 3.2, 3.3, 3.6, 4, 3.6, 3.6, 2.2, 1.5, 3, 2, 0.3, 2.1, 2.5, 
    2.7, 2.7, 3.2, 2.6, 2.9, 3.3, 2.4, 1.4, 1.1, 0.9, 0.1, 1.7, 1, 2.1, 4.4, 
    5.5, 7.3, 6.7, 6.3, 5.9, 5.5, 2.5, 3.9, 4.1, 5.4, 5.4, 6.8, 7.8, 8.8, 
    7.3, 9.1, 7.9, 7.2, 9, 9, 10.1, 10.1, 11.1, 12.8, 7.7, 6.9, 4.9, 5, 6.6, 
    6.1, 4.1, 3.5, 3.3, 3.4, 2.8, 2, 3.2, 5.2, 5.1, 3.5, 6.5, 5.2, 3.6, 6.1, 
    5.3, 7.9, 8.2, 8.2, 8.8, 7.2, 6.4, 6.2, 6.6, 6.4, 6.2, 8.1, 1.6, 15.4, 
    16.6, 16.5, 15.5, 12.6, 10.5, 8.5, 6.5, 7.7, 8.8, 9.6, 13.7, 13.5, 14.2, 
    13.8, 12.3, 12.7, 11.4, 11.2, 9.6, 10.4, 9.5, 7.2, 7.8, 7.1, 7.3, 6.9, 
    6.5, 7.6, 7.8, 7.7, 7.9, 7.3, 8.9, 7.5, 7.3, 8.1, 8.1, 8, 9.9, 8.8, 10, 
    9.6, 8.6, 8.6, 8.6, 8.6, 8.2, 12.3, 13.4, 10.9, 12.1, 11.7, 14.3, 13.8, 
    14.5, 16.1, 17.1, 16.5, 17.4, 16.8, 16.5, 15.2, 16, 16.8, 15.6, 14.8, 
    13.8, 14.5, 11.8, 10, 9.2, 7.8, 6.6, 7.2, 7, 8.3, 6.7, 7.8, 7.5, 7.4, 
    7.9, 9.3, 9.7, 10.9, 12, 10.2, 10, 8.2, 8.3, 7.4, 7.4, 8.1, 7.2, 7.1, 
    5.6, 5.3, 3.5, 3.2, 2.1, 1.6, 0.2, 0.1, 1.7, 4, 4.2, 3.7, 4, 4.1, 3.8, 
    3.1, 2.9, 2.7, 4.3, 3.1, 3.4, 2.7, 2.4, 3.5, 4.2, 4.9, 5.5, 2.3, 3, 1.7, 
    0.4, 1.2, 2.7, 3.1, 2.4, 3, 3.1, 4.5, 6.8, 6.9, 9.3, 9.7, 11.2, 11.9, 
    11.8, 12.7, 12.4, 13.1, 11.7, 10, 10.2, 10.3, 10.3, 10.4, 8.9, 9.6, 8.8, 
    9, 7.6, 8.1, 6.8, 7.9, 7.9, 8, 8.5, 9.6, 8.2, 8, 8.5, 8, 7.4, 5.3, 6, 
    4.9, 5.4, 6.6, 6.9, 5.6, 4.6, 4, 2.7, 1.6, 2.1, 0.1, 0, 1.3, 0.4, 0, 1.8, 
    2.9, 0.2, 0, 2.1, 1.4, 0.5, 2.1, 1.2, 3.7, 2, 1.1, 0.6, 5.4, 4.3, 3.3, 
    1.6, 1.6, 4.1, 3.1, 4.6, 2, 0.7, 0.8, 4.4, 5.2, 6.6, 6.7, 8.2, 8.3, 9.3, 
    8.4, 9.5, 8.2, 8.3, 8.7, 7.8, 8.1, 7.4, 8.9, 9, 12, 13.9, 12.1, 12.7, 
    13.3, 13.9, 13.3, 12.7, 12.8, 12.8, 13.2, 13.6, 13.4, 12.2, 9.9, 11.2, 
    10.8, 11.4, 10.5, 10.8, 11.3, 11.3, 11, 10.2, 10.1, 9.8, 9.3, 9.8, 8.8, 
    6.5, 8.2, 7.7, 8, 7.8, 7.6, 7, 8.5, 7.4, 7, 7.6, 8, 8.3, 7.9, 8.1, 6.7, 
    8, 6.7, 6.6, 5.9, 5.5, 5.8, 6.7, 7, 6.7, 6, 5.5, 6, 5.1, 6.1, 6, 5.9, 
    5.2, 5.2, 3.8, 4.1, 3, 3.4, 4, 0.3, 0.5, 0.3, 0, 0.3, 2.8, 4.8, 4.8, 5.5, 
    1.9, 0, 2.7, 5.3, 5, 4.3, 3.7, 3, 2.4, 0.3, 1, 2, 3.4, 3, 3, 3.7, 2, 2.6, 
    1.3, 1.2, 1.9, 4, 4.3, 2.9, 3.8, 4.4, 3, 5.8, 6.1, 6.4, 6.6, 6.5, 4.8, 
    3.9, 5.7, 5.4, 5.5, 6.7, 6.5, 5.7, 5.2, 5.1, 5.4, 5.3, 5.5, 6.1, 6.1, 
    7.3, 6, 5.7, 4.9, 4.9, 5.7, 5.8, 4.9, 4.8, 5.5, 5.4, 5, 5.6, 5.1, 5, 5.4, 
    4.3, 5, 5, 5.3, 5.9, 5.7, 5.8, 5, 4.9, 4.7, 4.6, 4.8, 4.8, 5.8, 4.7, 5.1, 
    5.2, 5.6, 5.9, 6.4, 6.1, 7.1, 4.5, 3.7, 3.8, 5.9, 5, 4.9, 5.1, 5.6, 4.6, 
    5, 4.5, 3.6, 4.1, 4.1, 4.7, 4.9, 5.3, 5.1, 5, 6, 6, 5.2, 4.8, 3.4, 3.9, 
    3.6, 4, 5.3, 5.3, 6.1, 5.4, 5.9, 6, 5.6, 4.2, 4.8, 4.4, 4.8, 5.3, 5.4, 
    5.1, 5.1, 5.3, 4.8, 4.8, 5.6, 4.7, 5.1, 6.2, 6.1, 5.3, 5.6, 6.1, 6.4, 
    7.2, 7.4, 5.6, 6.8, 5.7, 5, 4.5, 5.6, 5.8, 5.4, 5.4, 5.4, 4.5, 6.4, 6.1, 
    6, 5, 5.6, 7, 8.8, 8, 8.3, 8.5, 9.8, 12.2, 11.4, 12.9, 13, 11.4, 11.6, 
    11.9, 11.7, 12.6, 13.1, 14.6, 13.7, 13.7, 13, 14, 14.4, 14.4, 13.2, 13.5, 
    11.1, 10.6, 8.5, 7.3, 5, 3.8, 2.5, 0.8, 0, 8.1, 12.4, 12.3, 12.3, 9.1, 8, 
    8.4, 8.3, 0.1, 7.3, 4.9, 5.9, 6.9, 7.3, 6.9, 8.7, 6.7, 7.5, 8, 8.5, 10.3, 
    12.5, 12.6, 7.1, 4.7, 5.9, 17, 16.9, 16.9, 17, 15.2, 16, 14.5, 14.9, 
    13.3, 14.1, 14, 15.1, 15.9, 15.9, 15.9, 15.9, 17, 17.2, 15.8, 17.2, 16.6, 
    15.2, 15.2, 16.6, 16.8, 16.6, 18.8, 18.3, 17.3, 18.8, 17.9, 18, 18.4, 
    19.1, 18.7, 19.8, 19.7, 18, 18.4, 16.6, 15.9, 15.2, 15.5, 13.9, 14.6, 
    13.6, 16.4, 15.5, 14.2, 12.1, 11, 10.2, 10.6, 10.3, 9.2, 8.9, 8.4, 9.6, 
    7.8, 7.5, 5.2, 7.9, 3.6, 4.4, 5.5, 6.1, 4.3, 6.6, 7.1, 6.7, 7.6, 5.5, 
    8.5, 6.4, 6.4, 4.6, 3.8, 3.8, 2.7, 5.5, 2.5, 4.8, 3.9, 5.1, 4.1, 6, 4.1, 
    3.6, 5, 5, 4.5, 3, 3.6, 2.9, 3.8, 4.5, 4.4, 2.1, 2.7, 3, 1.2, 3, 4.5, 
    3.8, 4.7, 4.1, 1.5, 1.5, 1.4, 2, 1.4, 3.5, 2.2, 2.5, 1.5, 2.2, 1.1, 0.3, 
    1.8, 2.5, 2.5, 3.2, 2.4, 2.4, 4.1, 4.6, 4.1, 3.1, 2.6, 1.4, 2.5, 4, 4, 
    3.5, 4.8, 6.5, 4.8, 6.6, 7, 6.7, 6.6, 6.9, 7.2, 7, 5.8, 6.5, 5.7, 4.9, 
    6.1, 6.1, 6.4, 7.9, 5.8, 6.4, 5.1, 8.3, 6.8, 6.2, 7.6, 5, 6.2, 6.8, 6.5, 
    8.2, 7.2, 8.1, 6.9, 7.2, 10.8, 10.9, 13.8, 13, 11.2, 11.7, 9.7, 9.6, 9.2, 
    9.2, 11.5, 11.1, 11.5, 12.2, 13.4, 13.8, 11.2, 10.8, 10.6, 11.3, 9.7, 
    10.7, 11.5, 11.2, 13.6, 13.8, 13.4, 13, 13.1, 11.5, 8.5, 10, 9.4, 4.5, 
    3.5, 7.7, 4.1, 3.3, 3.3, 5.2, 6.7, 5.4, 3.4, 14.3, 15.7, 16.1, 16.9, 
    15.6, 11.1, 0.3, 1.9, 0.2, 6.9, 7.1, 8.7, 10.3, 10.6, 9.4, 10.8, 10.5, 
    10.8, 10.8, 10, 11.4, 10.1, 10.8, 8.2, 8.9, 8, 6.4, 9.2, 8, 6.1, 8, 4.7, 
    5.6, 6.9, 8.7, 8.8, 8.4, 6.9, 6, 7.1, 6.8, 7.3, 6.7, 6.3, 7.1, 5.4, 5.8, 
    3.5, 7.6, 2.9, 6.4, 5.3, 2.2, 8.6, 9.6, 8.6, 9, 10.2, 10.3, 7, 7.1, 5.2, 
    6, 5.2, 5.8, 5.1, 4.9, 4, 4.6, 4.4, 5.4, 7.7, 7, 8, 6.9, 8, 10.6, 9.6, 
    9.5, 8.5, 5.8, 9.6, 7.1, 8.4, 8.4, 7.5, 7.5, 4.9, 5.6, 4.5, 6.6, 5.7, 
    3.8, 6.4, 6.4, 4.7, 1.9, 2, 5.4, 5.2, 4.7, 3.8, 4.9, 2.1, 3.7, 6.5, 6, 6, 
    6.3, 5.4, 5.1, 4.4, 2.2, 5.1, 6.3, 5, 5.4, 5.4, 4, 3.1, 5.8, 6.4, 9.1, 
    8.1, 7, 7, 7.5, 6.2, 6, 5.8, 5.3, 4.7, 5.6, 5.2, 5.6, 5.7, 4.6, 5.2, 5.5, 
    4.8, 4.9, 5.1, 10.6, 8.3, 8, 8.5, 7.9, 4.9, 4.9, 5.3, 4.2, 4.2, 4.4, 4.3, 
    11.4, 10.7, 9.8, 10.6, 10.4, 7.9, 8.5, 6.5, 4.3, 4.1, 3.3, 5.9, 6.9, 5.7, 
    7.1, 6.1, 4.5, 5.9, 5.3, 4.6, 2.7, 3, 5.5, 4.4, 3.9, 4.7, 2.7, 4.7, 5.1, 
    5.7, 2.8, 2.6, 2.9, 5.4, 3.4, 4.6, 4.3, 5.2, 4.4, 6, 4.9, 3.6, 4.6, 2.7, 
    3.6, 4.4, 6.1, 4.4, 3, 3.6, 4.6, 4.4, 3.9, 2.5, 2.9, 3.6, 6, 6.3, 4.8, 
    3.1, 4.7, 3.7, 3.8, 4.2, 4, 2.8, 2.4, 0.9, 3.6, 2, 1.4, 2.1, 4.6, 7.2, 8, 
    7.7, 12.2, 13.7, 8.6, 9.9, 6.6, 6.1, 8, 6.7, 4.1, 10.7, 10.1, 10.3, 10.1, 
    10.7, 10.8, 10, 8.9, 8, 7.6, 6.5, 3.3, 2.1, 3.1, 7.1, 7, 8.9, 10, 10.2, 
    8.6, 6.9, 5.8, 6.5, 4.8, 7.4, 6.1, 8.1, 6.3, 6.1, 8.2, 8.5, 8.8, 8.6, 
    7.8, 6.8, 8.5, 8.2, 8.2, 7.9, 7.2, 8.3, 7.3, 6.6, 7.2, 7.9, 5, 5.6, 6.7, 
    7.5, 6.4, 5.3, 6, 6.5, 5.9, 9.4, 9.6, 8.6, 5.9, 6.4, 7.2, 8, 10.3, 10.8, 
    10.8, 10.8, 9.6, 10, 10.8, 10.1, 12.2, 12.4, 12.7, 11.6, 10.6, 11.7, 10, 
    9, 9.5, 9, 8, 10, 10.8, 11, 10.7, 9.8, 9.9, 10.9, 11, 12.4, 12.7, 10.5, 
    10.6, 10.5, 11.3, 10.6, 9.7, 10.3, 8.8, 10.1, 10.2, 11.4, 10.9, 10.4, 
    11.7, 10.5, 10.6, 10.6, 10.5, 9.7, 10.1, 10.3, 11.3, 12.6, 12.7, 12.8, 
    12.6, 13.5, 12.9, 12.5, 12.8, 11.7, 9.9, 9.8, 9.2, 9, 8.9, 8.8, 8.9, 9.4, 
    9.5, 9.3, 9.6, 8.7, 7.9, 7.4, 6.2, 6.4, 5.5, 5.7, 4.9, 4.9, 4.3, 3.8, 
    4.6, 4.5, 4.2, 4.2, 4.3, 4.6, 5.3, 3.9, 4.6, 3.7, 4.9, 4.6, 4.7, 4.9, 
    4.9, 5.3, 5.2, 4.7, 5.7, 5.7, 5.7, 5.9, 5, 6.1, 7.1, 7.6, 7.1, 8.3, 8.9, 
    8.3, 7.4, 8.5, 7.2, 7.2, 7.3, 7.6, 7.5, 7.1, 6.8, 5.1, 4.5, 5.4, 6.9, 
    5.2, 6.1, 4.9, 3.5, 3.8, 4.5, 4.3, 4.9, 4.5, 4.4, 4, 3.2, 4, 4.7, 4.6, 
    5.2, 4.7, 5.4, 4.5, 3.5, 2.9, 3.3, 2.6, 1.8, 1.8, 3.4, 4.5, 4.8, 4.3, 
    3.9, 5.5, 6.6, 7.3, 5.5, 6.4, 6.3, 8.1, 9.3, 8.5, 9.2, 9.5, 9.4, 9.5, 
    10.2, 10.5, 10.7, 10.9, 10, 10.2, 10.1, 9.3, 8.4, 8.2, 6.7, 5.9, 4.1, 
    3.7, 4.7, 4, 4.1, 5.4, 3.7, 4.3, 4.5, 4.3, 5.3, 5.5, 8.5, 8.6, 7.2, 7.3, 
    4.7, 5.6, 5.9, 7.4, 8.6, 9.8, 9.4, 9.8, 10.8, 11.6, 11.2, 11.4, 10.8, 
    8.9, 7.6, 7.7, 8.2, 8.7, 10.7, 9.6, 9.2, 9.9, 12, 10.7, 9.8, 9.3, 10.4, 
    15.1, 14.4, 16.8, 16.8, 16, 15.1, 16.1, 18.2, 20.6, 21.2, 20.9, 21.1, 22, 
    22.1, 22.4, 23, 19.9, 14.6, 8.8, 9, 8.6, 8.3, 7.3, 7, 2.7, 4, 3.3, 3.7, 
    6.2, 6.5, 7.9, 7.7, 10.5, 9.2, 10.4, 13.9, 12.9, 12.3, 10.6, 10.1, 7.7, 
    9.4, 12.1, 9.8, 10.9, 10.5, 8.3, 6.7, 2.8, 2.5, 1.9, 3.6, 18.2, 18.7, 
    18.3, 19.7, 21.3, 18.5, 20.9, 20.9, 18.9, 19.7, 23.6, 25.3, 25, 22.7, 
    23.4, 21.2, 20.5, 20.5, 20.1, 19.3, 19.1, 17.8, 17, 13.5, 13.6, 12.8, 
    12.9, 10, 4.5, 1.9, 0, 0.7, 1, 1.9, 3.4, 6.2, 5.8, 8.4, 7.7, 8, 9.5, 9, 
    9.1, 9.3, 8.4, 7.7, 7.8, 6.9, 7.4, 7, 6.4, 6.2, 5.7, 6.5, 5.8, 7.8, 8.4, 
    9.3, 6.8, 9, 8.6, 9.3, 9.9, 9.4, 7.8, 7.4, 5.6, 4, 4.5, 5.1, 6.7, 7, 4.2, 
    5.2, 5, 3.1, 2.1, 10.1, 10.1, 7, 9.1, 8.2, 10.5, 11.1, 10.8, 11.7, 12.3, 
    12.6, 12.5, 12.5, 12, 10.2, 12.3, 12.3, 10.4, 10.5, 7.8, 8.3, 7.9, 9, 
    8.3, 7.5, 6.5, 5.7, 4.3, 2.8, 3.1, 5, 6.6, 9.7, 7.5, 3.7, 2.7, 2.1, 5, 
    7.8, 9, 10.4, 7.6, 7.3, 8.6, 7.2, 5.4, 11.8, 11.4, 11.3, 10.6, 12.1, 
    14.3, 13.5, 12.4, 12, 11.1, 10.8, 10.2, 9.6, 10, 9.2, 9.2, 7.7, 8.6, 8.8, 
    9.5, 9.5, 10.8, 10.5, 10, 10.2, 10.5, 11.2, 15.5, 13.4, 14.4, 14.1, 13.7, 
    11.6, 9.5, 6.8, 4.5, 8.3, 9.4, 10.1, 11.2, 12.5, 13.2, 13.3, 13.1, 13.3, 
    12.2, 10.9, 10.3, 10.3, 11.2, 9.7, 10.5, 9.3, 9.1, 9.4, 8.8, 8.7, 10, 
    10.2, 10.3, 12.1, 13, 12, 12.4, 10.9, 11, 11.8, 12.5, 10.9, 11.8, 12, 
    11.3, 10.8, 11.7, 12.2, 11.4, 14.8, 14.8, 15.6, 16.1, 14.5, 13.8, 14.7, 
    15.5, 14.5, 13.7, 13.3, 13.3, 13.4, 12.8, 12.8, 12, 11, 11.9, 11.7, 11.8, 
    10.7, 11.6, 11, 10.9, 10.1, 10.1, 9.4, 10, 10.5, 9.3, 9.7, 10.2, 9.2, 
    7.1, 6.5, 6, 4.6, 3.9, 2.2, 3.8, 2.1, 6.5, 8.9, 6.6, 8.7, 10.3, 10.4, 
    9.6, 10.8, 14.1, 14.3, 14.7, 16.3, 17.8, 18.9, 20.8, 22.6, 23, 25.9, 
    24.3, 23.4, 23.2, 23.3, 21.7, 20.2, 18, 15.3, 13.7, 13, 11.5, 11.8, 11.1, 
    11.4, 11, 10.8, 11.4, 12.1, 8, 6.4, 6.7, 11.4, 12.8, 12.7, 13.2, 12.5, 
    12.5, 12.9, 13.1, 14, 14.7, 16.6, 13.3, 10.6, 2.3, 9.8, 10.7, 9.9, 10.4, 
    10.4, 11.1, 13.8, 14.8, 12, 5.6, 12.1, 10.7, 8.8, 8.9, 8.3, 8.6, 9.3, 
    7.4, 6.2, 5.7, 6.2, 6, 8, 7.2, 6.2, 9.7, 8.3, 7, 6.8, 6.5, 5.6, 3.8, 3.6, 
    3.2, 3.2, 3.9, 4.1, 5.1, 5.6, 4.7, 4.8, 1.2, 0.9, 2, 1.8, 1.2, 2, 1.6, 2, 
    1.7, 2.3, 5.8, 5.1, 4.8, 4.6, 4, 5, 3.7, 3.6, 4.8, 4.8, 5.9, 7.8, 8.3, 
    8.2, 8.2, 8.1, 7.5, 5.4, 3.5, 5.7, 5.7, 5.4, 6.2, 7.1, 6.3, 6.9, 7.7, 
    4.9, 4.1, 5.9, 5.4, 6.3, 7.3, 6, 6.1, 6.1, 6.3, 4.7, 6.2, 7.7, 4.9, 6.1, 
    5.6, 5.7, 4.9, 5.2, 5.2, 5.3, 3.1, 3.9, 4.8, 3.8, 3.6, 2.3, 3, 3.5, 3.6, 
    4.3, 4.6, 5.1, 6.3, 6.9, 7.4, 6.1, 7.4, 8.2, 9.1, 9.5, 11.1, 11.4, 12.2, 
    13.1, 13.1, 12.6, 11.7, 11.9, 11.5, 11.8, 12.3, 11.2, 11.5, 10.8, 12.1, 
    12.5, 12.7, 13, 13.7, 14.9, 14.8, 14.9, 13.9, 12.4, 11.8, 12, 10.7, 9.6, 
    13.7, 14.7, 15.6, 18.6, 19.5, 20.2, 21, 20.4, 19, 17.5, 15.1, 14.4, 14.9, 
    18.8, 18.3, 18.4, 17, 16.2, 15.7, 13.4, 14.9, 15.8, 16, 15.5, 13.6, 12.9, 
    10.3, 10.2, 10.1, 10.5, 11.2, 11.4, 12.1, 12, 11.8, 11.5, 11.1, 11.2, 
    11.5, 12.6, 12.4, 15.2, 16.4, 16.9, 16.6, 17.5, 17.2, 15.5, 16.2, 13.7, 
    15, 14.7, 15.2, 15.5, 16.1, 14.6, 15, 14.7, 15, 13.8, 14, 13.6, 12.6, 
    12.5, 12.4, 13.1, 12.5, 13.3, 12.1, 12.7, 12.5, 12.3, 11.1, 11, 11, 11.2, 
    8.5, 8.9, 8.6, 10, 9.3, 10.4, 10.1, 10.7, 10.4, 10.8, 10.5, 9.9, 9, 10, 
    9.5, 9.6, 10.6, 10.5, 8.4, 8.8, 7.6, 7.2, 3.4, 5.9, 7, 9.9, 9.5, 7.3, 
    7.7, 7.3, 7.4, 7.3, 6.5, 5.1, 7.5, 8.5, 8, 7.8, 8.5, 9.3, 9, 8.3, 8.8, 
    7.2, 7.6, 7.5, 7.7, 9, 7.8, 8.7, 8.6, 7.2, 7.7, 7.9, 6.3, 7.1, 9.4, 9.3, 
    8.9, 9.9, 9.8, 9.6, 9.4, 9.8, 9, 8.9, 10.1, 9.1, 8.5, 8.8, 9.4, 9.3, 9, 
    7.6, 7.8, 7.4, 7.2, 7.6, 7.1, 7.5, 8.2, 7.4, 6.9, 6.7, 8.5, 6.5, 4.3, 
    6.7, 4.1, 3.3, 4.6, 5.8, 6.7, 7.6, 8.5, 8.2, 7.7, 6.2, 6.9, 6.1, 7.2, 
    9.9, 9.4, 9.2, 10.3, 10.7, 10.3, 10.2, 12.7, 12.3, 11.3, 11.2, 10.7, 
    10.8, 11.7, 10.5, 9.5, 11.5, 9.5, 10.1, 9.3, 10.6, 9.2, 9, 9.7, 9.1, 9.9, 
    10.1, 10.2, 8.3, 9.4, 10.3, 9.8, 9.9, 11, 9.6, 7.7, 8, 8.4, 8.1, 9.3, 
    8.7, 7.5, 8.7, 10, 9.2, 10.6, 12.1, 14.2, 12.8, 11.6, 8.3, 4.1, 4, 9.1, 
    8.2, 8.4, 7.8, 6.6, 7.4, 10.5, 7.2, 9.2, 7.1, 7.1, 5.7, 6.3, 6.3, 4.9, 
    6.8, 6.7, 6.8, 6.1, 6.7, 7.5, 8, 8.2, 7.2, 7.2, 7.4, 7.9, 7.7, 5.9, 5.9, 
    5.3, 5.6, 5.5, 6.6, 6.2, 6.3, 8, 8.8, 9.2, 8.7, 9.6, 9.3, 9.5, 9.8, 9.3, 
    9.7, 9.5, 8.9, 8.7, 8.2, 9.1, 9.5, 9.9, 9, 8.7, 8.6, 9.8, 7.1, 7.2, 5.6, 
    7.2, 9.4, 9.4, 11.9, 9.4, 13.9, 13.8, 13.2, 13.7, 13.9, 13.3, 8.7, 10.3, 
    12.4, 12, 12, 11.4, 10, 10.6, 10.1, 10.1, 9.9, 11.6, 12, 12.1, 10.5, 
    10.3, 11.3, 10.2, 8.9, 10.8, 10.3, 11.5, 10.7, 12.3, 12.5, 12, 9.8, 11, 
    10.5, 10.1, 10.8, 9.8, 9.1, 10.3, 10, 9.7, 8.4, 8.1, 7.9, 7.5, 9.4, 7.1, 
    8.5, 9.1, 9.6, 9.3, 8.2, 9.4, 11, 10.7, 11, 10.7, 10.3, 8, 10.4, 11.6, 
    12.7, 14.8, 11.4, 12.9, 10.5, 11.4, 10.9, 12.2, 13.4, 13.5, 10.7, 11.9, 
    11.5, 12.2, 12, 10.5, 10.1, 10.8, 10, 10.7, 11, 10.1, 11, 10.3, 9.9, 
    10.3, 9.7, 8.4, 7, 5.9, 5.6, 5.3, 6.5, 5.4, 4.8, 4.2, 4.9, 5.6, 2.9, 3.9, 
    1.7, 4.5, 5.9, 4.4, 4.4, 3.5, 6.2, 5.7, 0.8, 3.8, 4.7, 3.5, 2.9, 0.9, 
    1.6, 2.4, 3.8, 5.3, 7.3, 5.4, 6.5, 5.6, 0.9, 1.3, 1.6, 1.4, 1.9, 6.2, 
    1.4, 1.5, 0.7, 1, 1.7, 2.7, 0.5, 0.5, 1.2, 3, 9.2, 4.8, 3.4, 10.5, 15.2, 
    16.8, 17.7, 18.8, 17.1, 19.7, 20.1, 18.4, 14.3, 13.4, 13.4, 11.6, 12, 
    12.5, 13, 15.7, 16.5, 17.8, 16.9, 16.1, 15.5, 14.5, 16.1, 16, 16.7, 16.5, 
    16.4, 16.3, 15.9, 14.7, 12, 8.2, 10.8, 8, 7.8, 7.5, 7.2, 6.9, 5.5, 5, 5, 
    5.1, 5.2, 5.7, 5.8, 5.3, 6.3, 8.7, 9.6, 8.5, 7.7, 7.5, 7.1, 6.3, 6.9, 
    3.1, 2.6, 0.9, 2.1, 3.2, 2.6, 4.9, 6.8, 6.3, 6.9, 8.7, 8.3, 8.7, 8.2, 
    9.2, 8.4, 9, 8.1, 6.1, 6.4, 4.9, 3.6, 4.5, 4.2, 3, 4.2, 5.3, 3.4, 4.3, 
    3.8, 2.7, 2.3, 0.6, 0.8, 3.7, 2.9, 4.6, 3.6, 3.7, 3.9, 5.6, 6.3, 6.7, 
    6.6, 8.6, 8.3, 9.1, 11.2, 11.5, 12.7, 12.7, 13.5, 14.2, 13.3, 13.5, 13.3, 
    13.9, 14.3, 12.5, 13.2, 13.9, 12.9, 11.7, 10.1, 11.2, 9.9, 11.9, 11.7, 
    13.4, 10.9, 8.5, 4.9, 7.2, 10.1, 10.1, 12.6, 16.5, 15.9, 15.9, 15.9, 17, 
    16.5, 17.1, 15.3, 17.5, 18.5, 17.6, 17.1, 17.4, 17.8, 17.7, 18.8, 18.3, 
    17.3, 17.1, 17.1, 17, 17.1, 17, 15, 14, 11.9, 11.3, 10.6, 10, 8.5, 6.9, 
    6.9, 5.2, 5.4, 7.1, 5.1, 3.3, 1.9, 2, 2.3, 3.2, 4, 5.8, 8.9, 10.5, 10.9, 
    9.2, 9.2, 12, 12.1, 11.9, 12.2, 12.4, 11.5, 10.6, 9.4, 9.5, 9.7, 10.1, 
    8.2, 9, 9, 9.4, 9.3, 8.8, 8.7, 7.9, 6.3, 6.5, 7.2, 7.6, 7.5, 8.3, 8.4, 
    8.4, 8.7, 8.6, 8.6, 9.4, 8.5, 8.8, 8, 8.3, 8.1, 6.7, 5.9, 5.7, 6, 5.8, 
    7.4, 7.2, 7.9, 8.1, 5.9, 7.5, 7.6, 7.3, 7.8, 6.4, 5.4, 4.4, 9.9, 8.9, 
    8.3, 6.2, 6.5, 7.3, 7.7, 7.5, 7.9, 7, 6.5, 7.5, 7.3, 6.7, 7.7, 7.2, 6.6, 
    7.3, 6.5, 5.9, 7, 6.6, 7.2, 8.4, 11.6, 8.6, 6.6, 6.5, 9.5, 8, 10.4, 15, 
    12, 1.4, 3.2, 6.4, 9.4, 11.8, 12.8, 15.1, 12.1, 12.4, 12.7, 11.4, 11.9, 
    10.3, 10.9, 11, 12.7, 11.2, 10.9, 11, 12, 11.4, 11.7, 13, 14, 14, 14.1, 
    12.6, 12.2, 12.8, 13.5, 13.8, 14, 13.2, 13.4, 14.8, 15.7, 14.3, 16.1, 16, 
    16.2, 15.1, 14, 13.8, 4.6, 0.9, 1, 9.8, 2, 6.6, 10.6, 12.1, 13.2, 15.9, 
    1.7, 4.6, 9.7, 11.3, 11.1, 11.5, 12.2, 12.1, 11.9, 12.6, 13.7, 16.7, 
    16.3, 15.1, 13.8, 13.9, 14.1, 14.9, 14.5, 13.5, 15.8, 15.7, 14.7, 14.4, 
    14.2, 14.2, 13.8, 14.5, 14.6, 14.3, 14.7, 15.7, 15.6, 16.6, 18, 17.8, 
    17.5, 16.7, 14.6, 14.4, 14.9, 13.4, 13.2, 14.6, 14.8, 14.3, 13, 12.8, 
    12.7, 11, 7.7, 3.1, 1, 0.9, 1.1, 1.2, 1.4, 1.5, 1, 3.5, 6.1, 6.4, 6.1, 
    6.8, 5.2, 5.1, 5.1, 5.2, 3.3, 5.4, 3.2, 3.2, 3.9, 2.9, 1.7, 2.2, 1.8, 
    2.1, 2.2, 2.3, 1.1, 13.3, 14.4, 14.8, 15.4, 16.5, 16, 15.7, 16.3, 17, 
    16.5, 15.7, 16.3, 15.8, 14, 14.5, 13, 14.5, 13.2, 13, 12, 12.4, 11.4, 
    10.9, 12.7, 12.4, 11.2, 11.5, 11.4, 10.5, 11, 11.2, 9.8, 9.1, 8.1, 10.7, 
    4, 8.3, 1.6, 4, 5.8, 13.2, 15, 14.5, 14, 14, 14, 14.6, 13.6, 13.4, 12.8, 
    13.4, 13.5, 12.6, 12.5, 12.4, 10.5, 10.9, 10.7, 11.3, 13.3, 13.9, 12.4, 
    12, 12.4, 11.8, 11.1, 11.7, 11.7, 10.8, 11.1, 10, 9.6, 9.5, 9.6, 10.2, 
    8.1, 8.1, 7.4, 7.3, 5.1, 3.8, 4, 3.7, 3.8, 2.6, 2.1, 1.5, 1.7, 0.2, 0.5, 
    1.3, 1.8, 4, 4.3, 2.5, 3.1, 2.3, 0.9, 1.4, 1.6, 4.7, 3.9, 3.9, 4.8, 5.8, 
    7, 7.5, 10.1, 12, 12.6, 13.6, 13.1, 11.8, 10.1, 9, 9.6, 9.6, 7.8, 7, 6.2, 
    7.7, 6.1, 4.5, 3.5, 3, 2.7, 2.9, 3.3, 1.9, 2.6, 2.9, 2.3, 1.9, 2.9, 3.1, 
    3.9, 2.9, 3.1, 3.1, 3.8, 5.7, 6.7, 5.6, 5.8, 6.2, 4.2, 4.2, 3.8, 6.4, 
    7.5, 6.1, 5, 5.2, 3.4, 2, 5.6, 1.8, 3.1, 2.1, 3.1, 2.1, 2.2, 3.9, 4.2, 
    2.9, 2.2, 4.1, 4.3, 4.2, 5.9, 5.2, 4.9, 5.5, 6.1, 6.8, 5.6, 5.6, 5, 4.9, 
    9.7, 9, 6.8, 7.8, 6.6, 4.9, 7.8, 6, 4.5, 4.8, 4.4, 5.9, 5.2, 6, 4.8, 4.2, 
    4, 4.8, 7.2, 7.1, 6.8, 6.2, 7.1, 5.3, 4.4, 3.9, 3.8, 3.8, 3.4, 3.9, 3.9, 
    5.6, 3, 3.8, 4.9, 6.2, 4.4, 9.4, 9.9, 8.1, 4, 7.3, 8.2, 6.6, 2.7, 2.9, 
    1.4, 6.5, 5.4, 5.5, 6.1, 3.7, 2.4, 3.6, 4.4, 4.3, 3.5, 4, 6.1, 4.2, 4.1, 
    7.1, 6.2, 4.8, 3.1, 3.7, 5.8, 5.9, 2.4, 1.8, 5.4, 4.8, 4.8, 4.8, 4.6, 
    8.4, 5.6, 5.7, 2.7, 11.6, 14.4, 14.2, 14.4, 15.2, 17.8, 18.4, 18.3, 18.3, 
    18.2, 0.9, 13.3, 13.6, 12.8, 12.8, 12.7, 12.3, 13.1, 12.1, 12.3, 12.5, 
    11.9, 10.3, 10.2, 10.4, 11, 11.1, 12.5, 12, 10.4, 10.9, 10.2, 11.2, 11.1, 
    11.5, 11, 11.2, 11.4, 10.5, 11.3, 10.6, 11.1, 10.9, 12.9, 11.6, 10.8, 
    10.5, 11.7, 11.2, 9, 9.4, 8.8, 9.7, 9.1, 8, 7.6, 8, 7.9, 8.1, 7.8, 7.2, 
    5.8, 5.5, 5.5, 5, 5.2, 5.4, 5.6, 6.1, 6.4, 7.2, 6.3, 6.2, 5.7, 4.5, 6, 
    6.3, 4.1, 4.8, 3.4, 3.5, 2.8, 2.2, 2, 2.4, 2.4, 2.3, 2.8, 2.8, 2.3, 2.3, 
    2.1, 1.7, 1.3, 1.3, 1.2, 0.2, 0.9, 0.7, 0, 0.4, 1.7, 0, 0.8, 1.3, 1.1, 1, 
    2.5, 3, 4.1, 4.8, 4.2, 5.2, 6.1, 6.3, 6.8, 5.4, 5.2, 5.1, 5.1, 4.9, 4.8, 
    2.4, 2.7, 1.6, 0.9, 1.3, 1.3, 2.3, 3.5, 3, 3, 2.3, 0.9, 0.8, 1.2, 3, 3.8, 
    3, 5.1, 3.2, 2.6, 1.9, 2.2, 0.9, 9.5, 10.1, 8.4, 6.8, 7.9, 8, 5.1, 4.9, 
    3.1, 0.5, 0.6, 2.1, 2.9, 1.9, 1.2, 0.1, 3.1, 3.1, 4.1, 5.7, 5.5, 6.2, 6, 
    7.2, 7, 7.7, 7.6, 7.5, 7.2, 5.1, 4, 5.3, 5.4, 5, 4, 3.5, 4.5, 3.5, 2.8, 
    2.6, 3.3, 4.7, 4.4, 4.1, 2.1, 2.4, 2.7, 2.4, 2.5, 3.5, 3.9, 4.2, 3.7, 
    3.7, 6, 5.7, 5.2, 4.7, 5, 5.8, 6.5, 6.2, 4.5, 4.4, 4.3, 4.8, 6.9, 7.3, 8, 
    7.2, 6.5, 7.1, 7, 6.3, 5.5, 5.3, 3.4, 3.6, 2.7, 2.8, 1.9, 3.9, 3.8, 4.2, 
    4.2, 3.8, 4.7, 4.4, 3.3, 3, 4.2, 3.2, 1.7, 3, 3.9, 3, 0.8, 3.4, 1.5, 0.7, 
    0.6, 1.3, 3.2, 3, 3.8, 4.1, 4.5, 4.6, 3.7, 2.5, 2.7, 1.5, 1.3, 10, 11.7, 
    11.7, 12.9, 11.8, 12.7, 14.1, 14.8, 13.8, 11.7, 12.9, 13.3, 14.3, 14.6, 
    14.5, 14.6, 14.7, 14.1, 13.4, 13, 13.4, 13.5, 15.2, 14.3, 12.5, 9.8, 8.8, 
    7.8, 5.8, 5.7, 5.9, 4.3, 4, 3.8, 2.6, 2.5, 1, 0.8, 1, 2.1, 2.9, 3.3, 3.5, 
    4.5, 4.5, 4.8, 4.7, 4.6, 4.8, 5.6, 6.3, 6.7, 7.1, 7.7, 7.6, 7.4, 7.3, 
    6.6, 6.8, 5.6, 4.7, 4, 3.7, 0.8, 0, 0, 1.4, 3.2, 2.2, 2.1, 3, 10.2, 10.6, 
    10.4, 8.8, 9.9, 10.6, 10.2, 11, 10.7, 9.2, 8.6, 8.5, 7.8, 7.4, 7.6, 8.2, 
    7.1, 7.8, 7.8, 7.5, 7.7, 7.9, 6.8, 7, 6.6, 5.9, 5.9, 7, 7.5, 6.9, 6.8, 
    5.9, 6.7, 5, 4.8, 3.9, 3.1, 1.2, 1.8, 1.3, 0, 0, 1.1, 0, 0, 1, 0, 0, 0, 
    0.3, 2.5, 5.7, 4.7, 4.2, 4.4, 5.2, 5.3, 5.6, 5.6, 5, 5.7, 4.8, 3.4, 3.3, 
    2.9, 2.2, 1.1, 1, 2.8, 3.8, 4.3, 4.4, 5.4, 5.8, 7.1, 9.2, 11.5, 11.7, 
    13.4, 13.7, 15, 13.8, 14.5, 14.4, 14.9, 14.2, 15.2, 15.9, 16, 15.9, 15.8, 
    14.9, 15.4, 15.4, 15.6, 16.3, 16.3, 16.8, 17.2, 17.1, 17.7, 18.1, 17.9, 
    17.8, 18.3, 19, 16.6, 15.7, 15.5, 16.6, 15.3, 14.6, 15, 14.1, 14.7, 13.9, 
    12.5, 13, 13.2, 10.8, 8.4, 9, 11.2, 8.6, 7.6, 10.8, 10.3, 11.2, 10.9, 
    8.7, 9.6, 8.1, 6.4, 6.3, 6, 7.2, 7.1, 6.2, 5.3, 5.2, 6.3, 4, 3.8, 4.7, 4, 
    4.6, 4.3, 4.7, 4.7, 4.3, 2.9, 1.7, 2.2, 1.1, 2.2, 1.8, 1.4, 0.7, 1, 1.4, 
    0.4, 0.4, 1.3, 0.9, 0.1, 1.5, 2.1, 3.3, 4.4, 5.4, 6.4, 6.6, 5.9, 6.8, 
    7.2, 6.2, 6.9, 7.1, 7.2, 8.1, 8.5, 8.6, 8.8, 9.5, 10.9, 10.4, 10.5, 10.7, 
    10.1, 11, 10.5, 10.9, 11.2, 11.6, 11.3, 12.4, 12.4, 12, 11.6, 10.3, 8.4, 
    6.3, 4.6, 0.7, 3, 2.4, 2.6, 4.3, 5.3, 5.6, 4.6, 3.5, 4.3, 4.1, 4.3, 3.4, 
    4.2, 4.1, 4.1, 5.5, 5, 4, 3.5, 3, 3.7, 3, 4.7, 6, 5.2, 5.5, 6, 7.1, 6.5, 
    7, 7.3, 7.3, 8, 8.7, 7.3, 6.9, 7, 7.1, 6.4, 6.9, 5.6, 5, 5, 5.9, 5.1, 5, 
    3.7, 5.7, 5, 5.1, 5.4, 5.7, 5.7, 5.8, 6.8, 5.8, 5.7, 4.7, 5.8, 6.1, 6.1, 
    7.1, 6.3, 7.9, 6.9, 5.9, 5.5, 5.4, 6, 6.3, 5.9, 7, 6, 6.7, 7.7, 7.2, 6.9, 
    6.8, 7.4, 7.6, 7.9, 8.2, 7.8, 8.1, 10, 8.3, 8.9, 9.2, 7.3, 8.5, 9, 9.4, 
    9.2, 10, 10.2, 10.7, 10.6, 11.1, 11.3, 11, 11.5, 12.4, 13.3, 13.7, 13.8, 
    14.4, 14.6, 14.2, 13.8, 12.7, 12.7, 12.5, 11.5, 11.4, 11.8, 10.8, 10.4, 
    10.3, 9.2, 9.1, 8.3, 7.4, 6.9, 6.7, 4.6, 4.3, 3.2, 2.6, 2.7, 2.1, 0.8, 
    0.2, 1.3, 1.1, 0.8, 1.6, 2.1, 2.5, 1.4, 1.5, 0.9, 2, 2.1, 2.7, 2.1, 1, 
    0.8, 0.2, 0.7, 3.5, 2.9, 4.2, 5.3, 4.8, 5.3, 6.4, 6.3, 6.8, 6.4, 6.6, 
    6.5, 7.2, 7.9, 8.9, 7.8, 8.4, 7.4, 7.3, 8.8, 9.2, 8.9, 8.4, 8.4, 7.2, 
    7.2, 7.6, 7.9, 7.8, 8.4, 8.7, 9.5, 8.1, 9.4, 9.4, 9.6, 9.4, 10.7, 10.8, 
    10.3, 11, 9, 8.6, 9.4, 9.4, 10.5, 11.4, 11, 10.6, 10, 10.5, 9.9, 9.6, 
    9.7, 8.8, 8.6, 8.8, 9.5, 10.9, 10.6, 11.5, 11.2, 11.5, 12.1, 11.7, 9.5, 
    9.8, 10.6, 9.9, 10.4, 10.4, 9.7, 9.2, 9.8, 9.9, 12.3, 15.4, 12.8, 11, 
    10.3, 11, 11.4, 11, 10.3, 10, 10.1, 10.2, 10.6, 11.6, 11.6, 11.9, 11.2, 
    11.5, 12.2, 13, 12, 12.5, 12.8, 13.1, 13.1, 13.3, 12.9, 12.8, 12.9, 12.1, 
    12.2, 11.1, 12.8, 12.3, 12.6, 12.9, 11.5, 10.2, 10.1, 14.3, 14.3, 14.5, 
    14.8, 15.2, 14.9, 13.4, 13, 12.4, 11.8, 11.7, 12.3, 12.2, 12.7, 12.3, 13, 
    13.3, 14, 14.5, 13.3, 13.3, 14, 13.9, 14.1, 14.2, 14.6, 14.8, 15.2, 15, 
    15.4, 15.2, 13, 14.2, 13.5, 11.5, 11.7, 12.9, 12.2, 11, 10.3, 10.3, 10.3, 
    10.9, 11.3, 11.8, 10.4, 11.1, 10.5, 11.7, 10.8, 10.9, 9.8, 9.3, 9.6, 
    10.9, 11.1, 11.5, 11.7, 12.3, 13.8, 13.4, 14.3, 12.9, 13.2, 13.6, 13.2, 
    12.2, 11.5, 11.4, 11.4, 11.7, 11.4, 11.3, 10.8, 10.9, 11.3, 12.4, 13.3, 
    15.2, 14.5, 16.4, 15.9, 15.9, 13.6, 14.4, 12.8, 13.3, 15.1, 14.6, 16.3, 
    18, 16.2, 17, 18.3, 14.6, 14.6, 14.3, 14.3, 14, 15, 15.2, 13.6, 12.2, 
    11.6, 12, 11.9, 10.6, 10, 9.8, 11.1, 9.9, 10.7, 12.6, 14.7, 14.5, 12.5, 
    10.1, 11.7, 11.2, 10.7, 10.8, 10.6, 10.4, 9.8, 11, 11.6, 13.9, 13.3, 
    11.7, 10.6, 10.2, 10.6, 11.6, 11.7, 12, 11.8, 12.8, 11.8, 12.5, 13.4, 
    14.1, 13.7, 12.5, 11, 9.8, 9.9, 9.7, 8.6, 9.3, 9.9, 9.7, 11.5, 11.3, 
    13.4, 13.7, 11.7, 12.6, 12.3, 10.6, 9.7, 8.1, 7.6, 8.8, 6.7, 9.1, 8.6, 8, 
    9.4, 10, 10.9, 11.1, 11.7, 11.7, 12.2, 12.2, 12.2, 12.6, 13.3, 13.3, 
    11.6, 11, 10.3, 10.5, 10.6, 9.7, 9.6, 9.5, 10.4, 9.9, 11.5, 11.1, 10.2, 
    8.5, 8.4, 8.4, 7.7, 8.4, 8.3, 8.8, 9.3, 8.4, 8.3, 8.3, 8.9, 7.8, 8.3, 
    8.3, 7.4, 5.6, 6.9, 7.8, 6.4, 7.1, 7.9, 7.6, 7.9, 10, 7.7, 7.1, 5.7, 5.8, 
    7.3, 7.6, 7.1, 7.1, 6.4, 7, 6.4, 7.7, 7.4, 4.1, 6, 6.5, 7.8, 8.1, 7.8, 
    8.2, 7.5, 7.2, 7.6, 8.1, 5.5, 4.1, 3.1, 2.4, 2.4, 3.1, 2.6, 1.9, 3, 2.9, 
    2.1, 3.1, 3.2, 2.8, 2.4, 2.9, 3.2, 4, 3.8, 4.9, 4.5, 3.1, 3.7, 2.5, 3.4, 
    1.3, 3.2, 3.1, 6.6, 6, 5.7, 3.8, 1.3, 4.9, 1.9, 3.6, 4.1, 5.2, 4.8, 3.9, 
    3.5, 1.7, 1.4, 4, 5, 5.7, 5.7, 4.2, 2.5, 2.2, 2.6, 4.7, 7.7, 8.3, 9.3, 
    8.5, 5.9, 6.3, 6.3, 5.3, 3.2, 2.5, 4.7, 6.9, 7.1, 7.3, 6.9, 5.3, 5.7, 
    4.6, 3.6, 4.6, 4.3, 5.6, 4.5, 6.5, 6.3, 7.2, 7.2, 8.5, 8.5, 8.8, 7.9, 
    8.1, 7.8, 9.7, 11, 9.4, 9.3, 9.4, 9.9, 9.2, 7.3, 7.8, 6.4, 8, 6.6, 7.4, 
    8.6, 7.5, 9.2, 11.3, 13.5, 14.7, 14.4, 15.6, 14, 14, 12.6, 10.6, 11.9, 
    8.4, 7.4, 9, 8.6, 11.4, 12.6, 13.1, 13.1, 9.6, 9.3, 10.2, 10.3, 12.3, 
    10.4, 11.6, 10.3, 12, 13.1, 11.5, 13.9, 12, 11.1, 12.1, 11.9, 11.9, 12, 
    12.5, 11.7, 12.5, 14.6, 14.3, 12.5, 8.9, 10.4, 11.5, 15.9, 16.5, 14.5, 
    13.4, 12.9, 12.5, 11.7, 12.5, 12.6, 4.7, 8.2, 7.2, 5.7, 5, 4, 2.4, 3, 
    2.6, 3.3, 2, 1.1, 1.4, 2.7, 3, 5, 6.7, 6.4, 5.9, 5.4, 4.2, 3.5, 4.6, 3.4, 
    5.5, 5.3, 6, 6.7, 7.6, 8.3, 8.2, 8.1, 11, 12, 13.3, 12.8, 12.8, 15.4, 
    15.3, 16.3, 13.3, 14.3, 13.2, 13.1, 16.7, 18.6, 17.8, 16.2, 16.8, 18.7, 
    18.1, 16.3, 15, 15, 16.7, 15.6, 15.4, 15.6, 17.9, 18.6, 15.9, 16.1, 15, 
    17, 17.4, 15.9, 16.2, 16.9, 17.1, 17.9, 15.1, 14, 11.6, 11, 10.3, 14.6, 
    13.5, 13, 11.7, 13.2, 10.3, 9.3, 10.1, 9.5, 9.2, 8.3, 5, 5.4, 3.4, 2.3, 
    0.8, 2.9, 2.3, 1.5, 0.9, 5.7, 8.6, 9.5, 9.2, 10.6, 11.6, 12.2, 13.5, 
    14.4, 14.5, 12.5, 10.4, 9.6, 8.2, 9, 9.2, 9.6, 11.9, 13.4, 14.3, 14.1, 
    15.2, 16.2, 17.1, 18.4, 17.7, 17.6, 18.6, 18, 17.3, 16.5, 15.1, 13.1, 
    8.7, 10.5, 12.1, 12.3, 13.3, 12, 12.6, 12, 12, 11.2, 12.5, 12.6, 12.5, 
    11, 10.1, 9.4, 9, 6.2, 3.5, 2.3, 1.8, 3.5, 5.4, 3.8, 7, 6.9, 5.4, 4.2, 
    5.9, 5, 5, 4.4, 6.2, 7.1, 7.6, 8.8, 10, 10.5, 10.3, 8.4, 7.3, 5.6, 2.7, 
    2, 4.1, 6.3, 6.2, 7.8, 6.6, 7.7, 5.8, 6.1, 6.6, 6.8, 9.3, 9.8, 10.3, 9.8, 
    11.3, 10.2, 11.1, 10.7, 13.7, 13.1, 13.7, 14.2, 13.2, 14.9, 15.5, 17, 
    16.9, 17.4, 16.1, 16.5, 16.6, 16.2, 16.3, 16.3, 14.2, 13.3, 14.5, 16.5, 
    17.4, 17.6, 17.9, 18.4, 17.4, 18, 17, 16.1, 14.4, 14.1, 13.6, 13.9, 14.4, 
    15.5, 15.1, 13.6, 13.3, 11.9, 11.5, 10.5, 11.1, 11.1, 11.5, 10.6, 9.8, 
    10.6, 11, 10.9, 11.8, 12.8, 13.7, 13.6, 14, 15.9, 15, 12.9, 13.4, 13.4, 
    11.8, 13.4, 13.8, 13.4, 12.3, 11, 10.6, 9.7, 6.8, 9, 9.3, 9, 7, 6.2, 8.1, 
    6.9, 5.4, 3.4, 4.7, 1.7, 5.6, 3.1, 4.5, 3, 1.2, 2.5, 4.2, 2.8, 4.7, 5.2, 
    5, 2.9, 2.2, 7.2, 8.6, 10.4, 11.8, 8.2, 4.5, 2.9, 6.8, 6, 9.3, 8.9, 7.7, 
    3.3, 10.2, 7.9, 7.5, 12.7, 12.1, 8.6, 10.6, 11.1, 10.5, 9.1, 11.5, 11.1, 
    10.5, 9.3, 8.7, 9.5, 9.1, 9.5, 8.6, 9.2, 8.9, 9, 8.5, 9.8, 9.6, 10.8, 
    9.1, 8.4, 11.7, 11.8, 12.7, 10.3, 10.1, 10.8, 11.2, 12.3, 12, 12.7, 12.5, 
    12.2, 11.9, 11.8, 12.2, 12, 11.3, 12.9, 12.8, 11, 13.4, 14.5, 12.9, 13, 
    13.4, 13.4, 13, 8.9, 8.6, 7.9, 10.5, 10.6, 9, 6.9, 5.5, 3.8, 3.8, 3.9, 
    4.4, 5, 4.1, 2.9, 2.1, 3, 2, 3.9, 4.3, 3, 3.3, 2.4, 3.1, 3.6, 2.4, 3, 
    3.4, 4.9, 5, 8, 8.9, 8.4, 8.7, 9.8, 9.6, 10, 9.6, 11.1, 10.9, 11.1, 11.3, 
    10.7, 11.5, 10.8, 11.9, 11.9, 11.6, 11, 11.5, 12.1, 12.9, 12.9, 12.3, 
    12.5, 14.1, 13.5, 12.5, 10.8, 10.7, 10.7, 9.5, 9.9, 9.6, 9.6, 9.7, 9.3, 
    10, 9.8, 10, 9.8, 9.4, 9.3, 9.8, 10.2, 10.2, 11.1, 10.9, 11.9, 12.6, 
    14.2, 14.8, 14, 14, 14.8, 14.9, 13.4, 12.5, 11.4, 13.2, 16, 16.8, 15.7, 
    19.5, 19.5, 20, 19, 17.8, 14.3, 17.6, 18.7, 19.4, 19.8, 18, 16.7, 16.6, 
    20.9, 20.9, 21.1, 20.1, 19.6, 16.1, 16.3, 14.8, 14.9, 13.5, 15.5, 14.7, 
    14.4, 15.8, 16.4, 16.1, 16.6, 17.1, 15.4, 16.4, 14.8, 13.4, 14.1, 14.5, 
    14.9, 14.2, 14.6, 11.8, 12, 13.9, 14.5, 14.2, 15, 14.7, 14, 14.8, 14.3, 
    13, 11.4, 8.8, 11.4, 11.7, 11.4, 10.6, 10.9, 8.9, 8.8, 8, 6.6, 7.3, 7.7, 
    8.5, 8.4, 7.7, 8.8, 9.1, 7.2, 5.8, 8, 9, 8.8, 9, 8.4, 8.3, 7.8, 6.6, 7.1, 
    6.2, 5.6, 6.3, 6.4, 6.2, 5.6, 5.7, 4.5, 4.1, 3.7, 5, 3, 3.5, 3, 3.7, 5.1, 
    4.5, 3.8, 4, 4.4, 3.4, 4.2, 1.9, 2, 1.2, 0.5, 5.7, 5.5, 3.7, 3, 5, 3, 
    2.4, 0.9, 1.7, 3.3, 4.8, 4.6, 3.6, 5.2, 5, 4.8, 6.6, 6.9, 5.8, 5.4, 6.7, 
    7.3, 7.4, 6.1, 5.4, 4.3, 2.8, 3.6, 1.8, 2, 3.5, 3.4, 2.9, 3.1, 2.8, 3.3, 
    4.8, 7.5, 9.1, 8.9, 9.5, 8.7, 8.6, 9, 9.3, 9, 8.8, 7.9, 7.2, 7.2, 6.7, 7, 
    4.8, 3.8, 3.8, 4.4, 4.3, 6.4, 5.6, 6.6, 6.6, 7.4, 7.8, 7.4, 6.6, 7.2, 
    6.8, 7.3, 6.5, 6.7, 6.6, 6.8, 6.3, 6.6, 7.4, 9.3, 9.2, 8.8, 8.5, 7.3, 
    8.2, 8.2, 8.2, 7.7, 9.4, 9, 8.7, 9.5, 7.2, 3.7, 2.2, 2.3, 4.3, 5.8, 3.8, 
    2.6, 7.7, 9.7, 8.7, 9.6, 10.2, 9.3, 9.7, 8.7, 9.5, 6.7, 8.5, 9.1, 10, 
    10.3, 13.5, 14, 13.1, 13.7, 13.6, 12.4, 11.1, 10.9, 9, 8.7, 7.3, 6.1, 
    4.9, 5.6, 6.7, 5.6, 6.4, 7.5, 8.9, 9.7, 5.6, 5.6, 6.4, 5.9, 5.3, 4.2, 
    2.3, 1.9, 0.5, 1.5, 0.4, 1.2, 3.6, 4.7, 5.3, 4.9, 6.4, 5.9, 7.4, 7.5, 
    8.3, 10.1, 11.1, 12, 14.8, 13.9, 13.6, 14.7, 14.4, 13.1, 13.1, 11.6, 10, 
    6.1, 0.8, 4.7, 5.1, 5, 9.8, 6.8, 5.5, 5.6, 8.2, 9.2, 9.5, 9.8, 8.6, 7.8, 
    8.5, 10.8, 9.2, 11.6, 15.4, 12.3, 14.4, 17, 16.3, 17.1, 18.7, 18.1, 17.6, 
    14.9, 16, 17, 18.2, 16.4, 19.2, 18.7, 18.3, 16.7, 17.4, 16.6, 17.5, 17.1, 
    17.9, 19.4, 21.2, 19.3, 17, 16.4, 16.4, 12.1, 12.3, 14, 14.6, 17.3, 14.1, 
    13.6, 14.6, 14.3, 16.1, 15.3, 14.6, 15.2, 16.1, 16.6, 17.1, 16, 15.7, 
    15.2, 14.2, 14.8, 13.2, 13.3, 14.4, 14.3, 15.7, 16.3, 15.3, 14.8, 15.2, 
    15.2, 15.4, 15.3, 15.3, 14.9, 13.3, 12.5, 13.2, 15.6, 15.5, 15.6, 15.8, 
    14.5, 14.2, 13, 12.2, 12.6, 13.9, 13.8, 12.2, 13, 12.5, 12.4, 11.2, 9.7, 
    11.2, 13, 11.2, 12, 11.7, 12.4, 12.5, 12.7, 11.5, 12.7, 12.6, 13.3, 13.6, 
    13.8, 13.9, 12.5, 11.9, 11.9, 11.2, 12.2, 12.5, 12.3, 13, 12.3, 11.2, 
    11.5, 11.1, 11, 9.3, 10.7, 9.4, 8.7, 10.2, 10, 9.5, 8.3, 6.2, 6.5, 5.9, 
    7.2, 8, 8.1, 8.7, 9.1, 10.2, 8.4, 6.7, 5.8, 3.8, 4, 6.3, 5.1, 6.2, 5.2, 
    9, 4.8, 6.1, 5.7, 5.9, 3.9, 3.6, 3.4, 4.2, 4.8, 3.6, 3.1, 3.4, 3.9, 3.6, 
    3.6, 5.2, 4.1, 3.4, 3.4, 3, 3.3, 3.3, 2.8, 3.3, 2.7, 4.7, 5.2, 4.8, 4.6, 
    4.4, 4.7, 3.8, 3.4, 2.3, 3.2, 2.3, 2.3, 7.3, 5.8, 5.8, 4.6, 4.8, 6, 5, 4, 
    7.8, 6.9, 10.3, 9.6, 11.5, 11.9, 12.4, 13.9, 13, 12.3, 11.9, 11.3, 11.7, 
    10.2, 10.4, 13, 12.7, 12.4, 12, 12.1, 12.4, 10.6, 9.8, 8.8, 9.4, 8.4, 9, 
    9, 9.2, 9.8, 8.7, 10.3, 8.7, 8.2, 9.6, 10.7, 10.3, 6.8, 7.4, 7.3, 7.4, 
    8.9, 7.3, 6.7, 9, 10.4, 9.8, 9.3, 8.9, 8.3, 9.2, 8.6, 7.6, 7.8, 8.6, 9.1, 
    8.6, 8.2, 7.9, 8.1, 7.6, 7.3, 5.1, 5.7, 5.6, 3.7, 3.8, 3.5, 1.9, 0.5, 
    1.5, 3.4, 4.2, 5.3, 5.5, 6.6, 6.8, 6.8, 6.7, 5.6, 5.1, 5, 6.9, 6.3, 5.9, 
    4.9, 4.6, 3.2, 2.7, 4.7, 3.1, 6.6, 5.3, 6.2, 5.7, 6.8, 3.8, 3.3, 0.2, 4, 
    5.5, 5.3, 10.6, 14.3, 14.2, 14.8, 16, 16.3, 14.6, 13.3, 14.4, 13.2, 9.5, 
    7.7, 4.1, 5.1, 2.7, 0.3, 0.2, 3.9, 2.5, 5.5, 2.2, 4, 2.6, 3.2, 17.1, 
    17.1, 16.7, 16.9, 15.5, 15.5, 12.2, 10, 12.8, 10.4, 12.7, 4.2, 7.7, 5.7, 
    8.1, 7.1, 5.7, 3.5, 5, 5.4, 2.8, 0.1, 0.9, 2.9, 4, 5, 3.1, 0.7, 0.1, 4.3, 
    5.7, 6.7, 5.6, 7.9, 8.6, 8.4, 8, 10, 11.3, 10.6, 11.1, 10.9, 10.2, 12.4, 
    11.3, 12.1, 9.9, 11, 13.6, 11.1, 8.1, 7.4, 7.1, 4.2, 7.8, 8, 7, 7.4, 6.3, 
    6.9, 7, 8.1, 8.5, 7, 4.8, 3.7, 3.8, 4.2, 5, 4.1, 5.3, 4.5, 4.1, 4.3, 3.8, 
    3.5, 3.7, 4, 3.5, 4.3, 4.3, 3.9, 4.1, 3.1, 3.1, 1.7, 2.4, 2.8, 2.2, 5.7, 
    6.4, 5.5, 7.9, 5.8, 7.9, 6, 8.8, 8.6, 7.2, 4, 5.9, 5.3, 3.5, 4.5, 5.5, 
    3.6, 3.7, 5, 7.1, 2.5, 2.2, 1.3, 2, 2.9, 5.6, 5.5, 6.8, 7.1, 5.8, 7.5, 
    3.3, 3.5, 3.2, 3.4, 2.6, 5, 3.2, 3.6, 3.5, 5.8, 6.5, 8, 7.5, 6.3, 6.1, 
    6.3, 7.4, 7.6, 9.8, 11.7, 13.1, 17.2, 13.9, 14.4, 14.9, 14.7, 15.9, 16.2, 
    14.9, 14.6, 14.6, 14, 13.8, 13.3, 12.3, 11.6, 11.6, 7.8, 4.6, 4.7, 4.8, 
    3.9, 6.3, 9.6, 12.7, 17.8, 16.7, 19.2, 17.8, 19.7, 19.5, 18.6, 16.3, 
    15.4, 18.4, 17.8, 17.6, 14.2, 14.1, 13.8, 13, 12.5, 13, 11.6, 9.2, 10.5, 
    9.8, 9.5, 9.6, 9.3, 7, 8.3, 9.4, 8.5, 9.8, 10.7, 8.4, 9.4, 8.4, 8.5, 9.6, 
    8.4, 9, 8.1, 9.1, 9.4, 10.4, 9.3, 12, 12.9, 13.3, 13.9, 13.3, 15.6, 14.3, 
    12.8, 13, 13.6, 11.6, 12.8, 13, 13.4, 12.5, 13, 14.4, 15.7, 14.6, 13.4, 
    14.4, 13.7, 13.7, 14.2, 12.7, 11.3, 10.8, 10.8, 9.9, 8.1, 9.1, 9.9, 8.4, 
    7.2, 6.3, 5.5, 3.4, 2.9, 1.8, 1.3, 1.5, 4.1, 3.6, 5.1, 4.2, 3.6, 4.5, 
    5.9, 6.2, 4.9, 5.4, 6, 6.2, 6.7, 6.1, 6.1, 6.2, 7.3, 6.9, 6.9, 7.9, 7.6, 
    8.6, 7.9, 9.3, 10.1, 11.1, 12.7, 11, 10.8, 12.2, 11.7, 10.7, 12.2, 12.5, 
    11.9, 11.1, 11.4, 11.5, 10.5, 10.5, 10.3, 10.5, 9.3, 9.3, 10.2, 8.4, 8.7, 
    9.1, 9, 8.4, 9.1, 7.4, 7.6, 7.9, 10.2, 7.6, 9.1, 9.3, 8.3, 7.5, 8.3, 7.5, 
    8.2, 7.7, 4.2, 3.9, 5.1, 6.9, 5.9, 8.3, 9.2, 9.8, 8.3, 9.3, 10.3, 10.6, 
    10.4, 11.7, 12.4, 11.7, 12.1, 10.5, 9.8, 12.7, 12.3, 11.2, 12.3, 11.4, 
    11.1, 10.4, 9.8, 11.4, 11.8, 11.6, 10.4, 10.7, 9.9, 8.9, 8.6, 8.6, 11, 
    11.5, 12.1, 10.5, 10.9, 11.3, 10.8, 9.8, 9.3, 10, 11.2, 10.7, 9.5, 9.6, 
    9.3, 12.4, 12.5, 14.6, 14.3, 14.3, 12.6, 13.9, 12.3, 11.1, 11.1, 12.5, 
    12.9, 12.8, 13.4, 13.2, 13, 12.8, 12.5, 12.5, 13, 12.9, 12.5, 11.3, 11.1, 
    11.2, 10.6, 10.8, 11.5, 9.8, 9.2, 10, 7.9, 5.7, 3.8, 5.6, 4.4, 4.4, 5.1, 
    4.2, 4.7, 2.8, 2.6, 4.5, 6.5, 7.3, 6.8, 6.6, 4.3, 3.6, 3.8, 4.2, 3.1, 4, 
    3.9, 4.3, 3.2, 3.7, 3.9, 5.7, 7.5, 8.8, 8.7, 9.4, 10.4, 11.2, 11.5, 11.1, 
    12.2, 15.6, 11.1, 14.5, 13.3, 14.8, 14.8, 12.7, 13.6, 8.6, 8.8, 8, 11.1, 
    10.5, 8.1, 7, 6, 6.7, 7.5, 7.1, 6.2, 7.6, 7.4, 6.9, 7.7, 6.8, 7.5, 6.6, 
    7.4, 7.2, 6.6, 7.6, 8.1, 7.6, 8.1, 8.9, 7.8, 7.3, 7.7, 7.3, 8.6, 7.8, 
    8.7, 9.2, 9.8, 10.8, 11, 10.6, 10, 9.3, 10.6, 9.6, 9, 8.8, 8.5, 8, 6.2, 
    6.9, 9.2, 9.3, 7.6, 8.2, 8, 8.7, 8, 9.6, 7, 5.6, 7.1, 5.5, 6.6, 6.7, 5.4, 
    6, 2.7, 2.4, 3.3, 4.6, 3.7, 5.9, 5.9, 7.3, 8.3, 6.2, 5.7, 6.3, 5.2, 5, 4, 
    5.7, 4.8, 5, 5.8, 4.8, 6.4, 6.8, 6.6, 6.3, 5.9, 6.4, 6.8, 7.1, 8.2, 8.5, 
    10, 9.9, 9, 8.8, 9.4, 9.7, 9.5, 8.7, 9.2, 10.3, 10.4, 10.6, 10.2, 9.3, 
    12, 10.2, 9.2, 10.8, 9.3, 9.1, 9.5, 9.4, 8.8, 8.8, 8.8, 9, 10.2, 9.1, 10, 
    10.2, 10.2, 9.6, 10.1, 10.3, 9.2, 8.8, 8.1, 7.6, 7.8, 7.7, 6, 5.1, 6, 
    3.5, 2.9, 1.5, 0.8, 1.2, 1.9, 1.9, 1.3, 1.2, 4.4, 3, 3.2, 4.3, 5, 3.9, 
    4.7, 4.9, 4.5, 4.1, 4.7, 5.5, 5.8, 6.6, 7, 7.2, 8, 8.6, 7.5, 6.3, 7.3, 
    4.9, 6.8, 4.6, 4.1, 4.8, 2.1, 1.5, 2.3, 3, 3.9, 4.2, 5, 4.2, 4.8, 3.4, 
    3.7, 1.8, 0.9, 1.3, 1.7, 0.5, 1.1, 1.9, 1.8, 2.8, 3.2, 2.1, 2.5, 4.5, 
    5.5, 6, 5.7, 5.8, 5.7, 4.8, 4, 3.8, 3.8, 3.9, 4, 4, 3.9, 4.8, 4.3, 4, 
    3.2, 3.8, 5, 14.1, 11, 9.7, 7.7, 12.4, 12, 13.1, 15.3, 14.6, 14.2, 12.1, 
    10.1, 10.3, 9.9, 8.5, 7.8, 6.6, 6.8, 7.3, 6.9, 1.9, 0.1, 1.5, 1, 0.7, 
    0.7, 0.7, 1.5, 1.7, 3.6, 3.4, 2.5, 1.8, 2.6, 1.7, 1.2, 1.4, 0.2, 1.1, 
    1.4, 2.5, 3.3, 3.1, 2.6, 2.1, 1.8, 4.6, 6, 6.1, 7.4, 6.3, 4.3, 3.4, 3.6, 
    2.7, 3.1, 6.7, 7.3, 7.9, 6.9, 6.2, 4.3, 4.3, 5.1, 3.7, 3.6, 2.6, 3, 3.2, 
    3.4, 2.5, 3, 3.5, 3.8, 2.6, 1.7, 1.6, 0.8, 0.8, 1.7, 2.1, 2.1, 2.3, 3, 
    3.7, 4.9, 6.6, 6.2, 7.8, 7.7, 7.8, 7.8, 10.5, 11.1, 12.7, 14.1, 13.5, 
    12.7, 11.9, 12.4, 12.9, 11.5, 11.6, 10, 8.7, 9.5, 9.6, 10.3, 3.5, 2.7, 
    2.2, 4, 5.5, 4.4, 4.6, 2.8, 4.3, 3.3, 4.2, 4, 3.1, 1.6, 1.7, 2.6, 1.9, 
    2.7, 2.7, 2.5, 1.4, 1, 1.4, 1.4, 2.5, 2.4, 3.5, 3.6, 3.6, 3.9, 3.6, 3.7, 
    2.9, 4.5, 2.9, 1.4, 5.3, 4.7, 6.1, 5.6, 7.2, 8.4, 7.3, 6.5, 6, 10, 10.3, 
    11.7, 10.5, 8.4, 6.6, 7.4, 7.1, 6.4, 7.6, 7.7, 6.8, 6.5, 7.4, 5.9, 6.1, 
    7, 7.9, 8.3, 9, 8, 9.4, 8.6, 8.3, 7.9, 6.7, 6.4, 3.8, 4, 2.4, 1, 2.5, 
    3.2, 3.3, 2.2, 0.5, 2, 0.4, 0.9, 1.7, 3.3, 3.6, 3.4, 2.5, 3.4, 4.3, 4.9, 
    4.4, 5.8, 4.1, 4.7, 4.7, 5.1, 5.3, 6.6, 7.5, 9, 9.8, 11.1, 10.4, 11.9, 
    10.9, 11.1, 8.2, 9.4, 12.7, 11.9, 12.5, 11, 9.3, 8.4, 5.7, 5.8, 8.2, 8.2, 
    8, 11.6, 9.7, 12.4, 14, 16.7, 17, 15.6, 16.1, 11.1, 10.6, 10.2, 8.3, 9.8, 
    10.5, 7.6, 9.2, 10.4, 10.5, 8.1, 8.2, 9.7, 10, 8.5, 8.5, 8.8, 8.9, 8.9, 
    7.1, 7.6, 8.7, 5.5, 6.3, 5.7, 4.8, 7.5, 8.1, 5.1, 5.9, 5.9, 7.1, 6.1, 
    4.2, 2.9, 0.4, 2, 0.5, 2.3, 4.7, 4.6, 2.7, 3.4, 3.5, 3.9, 3.4, 3.7, 1, 
    3.6, 1.7, 2.1, 3.7, 5.8, 4, 6, 6.5, 4.7, 5.6, 5.5, 6.6, 6.8, 7, 6.4, 6.8, 
    5.3, 5.5, 6.3, 6.5, 6.8, 5, 6.6, 5, 6.4, 6.7, 6.5, 4.9, 5.1, 5.5, 5.7, 
    6.6, 8.2, 9.1, 10.5, 10.3, 9, 10.4, 10, 7.1, 10.9, 11.4, 12.1, 10.5, 
    11.6, 11.7, 13, 11.7, 11, 9.8, 9.5, 7.8, 8.5, 10.4, 9.3, 8.8, 7, 6.1, 
    7.5, 8.2, 6.7, 8.7, 9, 9.7, 8.7, 7.6, 5.3, 6.6, 8.9, 7.7, 9, 10.6, 9.5, 
    8.1, 8.8, 9.1, 11.5, 11.5, 10.6, 9.2, 9.2, 8.9, 10, 9.4, 8, 8.2, 9.8, 
    9.3, 9.1, 8.1, 8.8, 9, 11.5, 11.7, 9.2, 4.8, 8.9, 8.7, 9.6, 7.7, 6.4, 
    6.6, 6.4, 5.9, 8.2, 9.1, 10.6, 11.2, 12.8, 10.8, 10.8, 11.7, 12.9, 12.6, 
    13.3, 11.9, 10.4, 10.7, 12.4, 14.1, 15.1, 14.5, 15.5, 15.6, 15.8, 15.3, 
    16.1, 17.4, 16.9, 16.7, 18.6, 17.8, 17, 16.4, 16.2, 16, 16.1, 16.1, 14.1, 
    14.7, 14.8, 13.2, 14, 13.6, 13.8, 12, 11.2, 11.7, 10.9, 11.8, 9, 9.2, 
    9.1, 8.8, 9.4, 9.2, 9, 8.5, 7.1, 5.5, 5.3, 3.9, 3.4, 4, 1.2, 1.3, 0.5, 
    1.9, 2.4, 2, 2, 4.1, 4.3, 4.7, 4.9, 6.1, 6.7, 6.8, 8, 8.9, 8.8, 8.8, 8.6, 
    7.6, 7.1, 5.7, 5.2, 3.5, 2.3, 2.6, 1.5, 0.6, 1.6, 1.7, 1.6, 2.9, 4.8, 
    5.4, 4.4, 3.8, 5.2, 6.2, 5.4, 5.6, 6.6, 3.6, 4, 4.1, 2.1, 3.9, 4, 4.1, 
    3.1, 0.9, 0.6, 1.1, 1.6, 0.1, 0, 1.4, 2.1, 2, 2.3, 2, 1.2, 1.2, 1.5, 1, 
    0.6, 0, 2.3, 1.2, 4.9, 4.1, 1.4, 2.7, 2.6, 3.5, 5.6, 4.5, 4.9, 3.3, 4.2, 
    4.7, 4.7, 5.2, 3.9, 2.6, 0.1, 2.5, 4.3, 3.8, 2.6, 4.8, 4.8, 3.9, 4.3, 
    3.1, 3.2, 1.9, 1.4, 1.1, 1.7, 3.3, 4.1, 4.7, 4.5, 4.3, 3.6, 4.1, 6.6, 
    5.6, 4.8, 5.1, 5.6, 4.3, 5.7, 6, 4.5, 4.9, 4, 5.3, 5.1, 5.2, 5.9, 5.2, 
    4.6, 4.3, 4.5, 4.6, 7, 6.6, 4.1, 4.4, 4.4, 3.4, 4.3, 3.2, 3.5, 3.7, 5.4, 
    4.9, 4.5, 7.1, 7.7, 7.1, 6.5, 6.4, 8.3, 8.4, 8.6, 6.6, 6.2, 6, 4.5, 4.7, 
    4.9, 3.8, 3.2, 2.8, 1.8, 0.5, 0.4, 2, 4.2, 4.5, 4.9, 4.7, 5.4, 5.3, 5.7, 
    5.8, 5.8, 4.9, 5, 4.4, 4.3, 4.2, 2.6, 1, 1.7, 1.6, 2, 5.8, 4.2, 6.2, 6.6, 
    8, 8, 7.3, 7.7, 6.6, 7, 6.6, 7.5, 6.7, 7.4, 5.7, 6.4, 5.6, 4.5, 5.9, 7.8, 
    7.4, 6, 5.8, 3.5, 3.9, 3.5, 1.8, 2.4, 2.4, 1.6, 0.1, 4.6, 5, 5, 5.7, 5.9, 
    6.1, 6, 6.5, 7.1, 6.3, 5.7, 3.7, 4.4, 4.9, 5.6, 6.1, 6.4, 7.6, 6, 7.2, 
    7.8, 8.5, 8.1, 8.1, 8, 7.2, 7.4, 8.8, 8.5, 9, 7.9, 7.6, 7.6, 8, 7.6, 7.3, 
    7.2, 6.7, 5.9, 3.8, 2.5, 1, 1.7, 3.5, 4, 5.5, 4.5, 5.2, 4.8, 4.3, 5.5, 
    5.3, 6.3, 5.7, 5.6, 5.5, 4.1, 5.1, 4, 3, 2.6, 2.7, 1, 0.1, 1.2, 1.1, 0.7, 
    3.2, 5.2, 6.4, 7.3, 7.8, 8.9, 9.7, 10.7, 11.5, 11.7, 10.6, 9.8, 8.3, 8.8, 
    8.1, 8.5, 10.1, 9.7, 8.7, 9.1, 8.5, 8.1, 8.1, 8.6, 8.9, 9, 9.2, 9.3, 8.8, 
    7.5, 6.1, 3.1, 7.2, 8.1, 7.9, 7.2, 5.3, 6.3, 6.7, 7.3, 7.3, 6.9, 6.5, 
    5.8, 5.9, 6.3, 6.7, 6.2, 7, 6, 7.1, 5.9, 6.1, 6.3, 5.1, 4.1, 3.5, 2.9, 
    2.2, 1.3, 0.2, 1.1, 1.2, 0.3, 1.8, 2.2, 1.8, 2.9, 4.2, 4.7, 5.2, 5.8, 
    6.3, 5.8, 5.9, 4.5, 5, 5, 3.9, 1.5, 3.1, 2.7, 5.7, 5.1, 6, 7.5, 8.9, 8.7, 
    7.2, 7.4, 6.7, 6.2, 7.1, 6.1, 6, 4.7, 4.7, 3.4, 2.9, 2.5, 2, 1.7, 2, 1.3, 
    0.5, 1.3, 2.9, 2.8, 1.7, 3.9, 3.7, 3.8, 2.4, 2.3, 1.2, 4.6, 7.9, 8.4, 
    7.7, 6.4, 6.1, 7.2, 7, 6.9, 6.5, 5.4, 5.8, 6.5, 5.6, 6.5, 5.4, 6, 4, 2.5, 
    1.9, 3.9, 5.3, 5.9, 7.4, 5.9, 6.3, 6.1, 7, 5.2, 3.2, 2.9, 1.1, 4.5, 3, 
    3.6, 4, 4.6, 5.8, 6.7, 6.1, 6.7, 6.1, 6.4, 4.5, 5.4, 4.4, 5.6, 6.7, 6.1, 
    6.5, 5.7, 5.9, 6.1, 5.8, 4.6, 3.8, 5, 4.8, 5, 5.4, 6.3, 3.9, 3.8, 2, 0.2, 
    1.4, 2.1, 6.8, 7.5, 9.6, 9.7, 6.6, 6.8, 7.9, 9.8, 12, 6.3, 8.7, 7.1, 6.6, 
    9.8, 13, 12, 11.8, 11.2, 11.6, 9, 7.2, 7.5, 8, 9.8, 10.2, 4.8, 2, 6.3, 
    4.6, 3, 6.8, 6.6, 6.4, 6.2, 7.8, 5.8, 6.7, 6.1, 7.1, 6.9, 6.8, 7.5, 7.1, 
    8, 8, 8.2, 8.3, 7.3, 8.3, 8, 8.4, 9.3, 8.9, 9.3, 9.3, 8.8, 8.5, 9.8, 8.9, 
    8.9, 9.5, 9.2, 9.2, 10.1, 11.1, 10, 3.2, 4.3, 6.2, 7, 4.9, 6.4, 6.5, 7, 
    7.2, 8, 10.4, 11.4, 12.9, 12.2, 13.7, 12.5, 12.1, 10.7, 11.4, 12, 11.3, 
    12.4, 12, 10.6, 10.4, 12.8, 14, 13.8, 13.6, 11.7, 12.1, 11.9, 11.8, 11.3, 
    11.1, 11.3, 11.2, 10.7, 10.1, 9.2, 8.5, 8.2, 7.8, 8, 7.8, 6.5, 5.3, 4.8, 
    7.3, 7.9, 9, 6.7, 5, 5, 4.4, 6, 6, 7.8, 5.2, 3.9, 6.1, 5.3, 4.9, 5.4, 6, 
    4.8, 6.1, 6.9, 7.8, 10, 9.7, 9.4, 9.4, 7.3, 5.6, 5.5, 4.9, 5.5, 7.7, 6, 
    5.5, 7.8, 6.6, 7.6, 7, 8.8, 8.9, 8.7, 8.5, 8.6, 7.5, 7.5, 7.6, 6.6, 6.1, 
    6.1, 7.3, 7.7, 6.8, 6, 5.7, 5.7, 5.1, 4.5, 4.1, 5.9, 6.9, 8.6, 10, 10.1, 
    9.2, 9, 9.2, 8.3, 7.7, 7.8, 8.5, 8.7, 8.6, 7.6, 7.5, 8.1, 6.7, 6.5, 6.5, 
    5.2, 5, 4.7, 5.8, 6.8, 4.3, 4.8, 6.4, 6, 5.9, 6.3, 7.4, 6.5, 5.6, 5.4, 5, 
    5.8, 6.6, 5.2, 5.6, 6.8, 6.7, 6.1, 6.3, 7.6, 7.9, 7.8, 7.1, 6.7, 5.4, 
    6.7, 6.8, 5.8, 6.1, 5, 4.2, 3.1, 2.2, 2.2, 1.4, 1.3, 0.4, 0, 0.1, 0.1, 
    0.4, 0.6, 0.4, 1, 1.4, 1.7, 1.7, 1.7, 2, 2.6, 3.1, 3.7, 3.7, 4.5, 3.4, 
    1.6, 1.6, 1.9, 0.3, 0, 0.9, 1, 0.1, 0.4, 0.3, 0.7, 1, 0.2, 0.3, 0, 1.1, 
    0.9, 2.2, 1.9, 0.9, 7.1, 9.2, 7.5, 6.5, 5.2, 6.4, 7.1, 4.8, 3.9, 2.6, 
    2.2, 1.9, 1.7, 1.4, 0.9, 2.7, 0.8, 1.6, 2.5, 1.6, 1.3, 1.9, 1.5, 2.9, 
    2.3, 2.9, 3.2, 2.2, 2.6, 2.8, 2.4, 3.1, 3.4, 2.9, 4.6, 3.2, 3.2, 2.5, 
    2.6, 2.6, 3.2, 3.5, 1.9, 2.1, 3.1, 3.2, 3.4, 3.8, 3.8, 3, 3, 2.4, 2.7, 
    1.9, 2.2, 1.6, 2, 2.6, 1.9, 1, 1.3, 2.1, 2.2, 2.2, 2.7, 2.4, 2.3, 1, 1.3, 
    1.8, 2.3, 3, 3.7, 3.2, 3.7, 3.8, 4.1, 4, 3.7, 4.1, 5, 5.3, 6.2, 6.6, 7.3, 
    8.3, 8.6, 8.7, 7.6, 8.2, 9, 9.6, 10.7, 9.3, 9.5, 11, 11.7, 13.1, 11.6, 9, 
    10.6, 10.8, 9.5, 8.7, 8.2, 10.1, 10.2, 10.2, 11.4, 11.6, 12.6, 12.9, 
    12.7, 13, 12.1, 12, 13, 14.1, 14.6, 14.5, 14.4, 14.4, 14.2, 14.1, 13.8, 
    13.5, 12.9, 13.1, 12.9, 12.1, 11.9, 11.7, 10.5, 10, 9.5, 9.1, 8.4, 7.2, 
    7.2, 8, 2.6, 2.4, 2.6, 2.6, 1.6, 0.9, 0.8, 0.7, 0.7, 0.1, 0.6, 0.8, 0.2, 
    0.2, 0.6, 1.5, 1.5, 3.3, 3.9, 5.1, 5, 4.9, 5.2, 5.4, 4.9, 4.8, 4.4, 5.9, 
    5.2, 4.9, 4.6, 4.2, 2.9, 2.7, 2.9, 3.9, 4, 5.1, 4.8, 3.6, 3.5, 2.1, 4.3, 
    4.5, 3.5, 3.5, 2.6, 2.9, 2.3, 2.5, 2.3, 2.1, 3.1, 2.1, 2.6, 2.2, 1.6, 
    0.9, 2.1, 1.5, 2.6, 3.9, 6.1, 6.8, 5.8, 6.8, 6.9, 7.3, 6.7, 5.5, 6.8, 
    6.8, 6.4, 7, 6.1, 6.5, 6.3, 6.2, 6.2, 5.1, 3.9, 4, 3.8, 3.4, 3.9, 2.7, 
    3.3, 3.2, 2.8, 1.8, 0.1, 1.1, 0.7, 0.7, 1.4, 1, 1.3, 0.7, 1.1, 1.6, 1.1, 
    2.2, 2.7, 2.4, 3.2, 3.6, 4, 3.8, 3.7, 4.1, 4.5, 4.6, 4.1, 4.4, 1.7, 1.1, 
    0.1, 1.4, 1, 3, 4.8, 6.5, 6.6, 6.9, 7.1, 5.7, 3.9, 3.5, 4.3, 5.2, 6, 7.8, 
    9, 8.2, 7.4, 5.9, 4.4, 5.5, 6.5, 5.7, 6.1, 6.8, 5.8, 5.4, 7, 5.8, 7.6, 
    6.5, 7.2, 7.8, 8.8, 8, 7.6, 8, 7.4, 5.9, 5, 5.7, 5.3, 4.9, 5.4, 4, 3, 
    0.3, 2.2, 2.4, 3.5, 4.4, 6.1, 4.9, 4.8, 5.7, 6.7, 6.6, 6.5, 6.9, 7.4, 
    7.2, 7.1, 6.7, 5.5, 4.2, 3.9, 2.1, 0.3, 0.9, 1, 1.1, 0.8, 1.4, 4, 3.8, 
    5.7, 5.9, 5.4, 3.1, 2.9, 1.2, 1.8, 2.4, 2.3, 3.4, 10.9, 8.1, 9.2, 11, 
    12.5, 11.2, 9.2, 7.2, 4.6, 1.1, 2.4, 5.9, 6.6, 8.1, 7.7, 6.6, 5.7, 4.3, 
    5.4, 7.3, 7.1, 7.4, 7, 6.5, 3.9, 1.6, 0.6, 0.7, 1.4, 1.2, 0.9, 0.9, 1, 
    1.2, 3.3, 2.2, 1.7, 1.3, 1.2, 2, 1.9, 1.8, 5.9, 7.8, 7.9, 7.2, 7.5, 8, 
    8.5, 7.2, 6.4, 5.5, 5.6, 6.8, 6.5, 6.8, 6.6, 7.2, 8.1, 9.1, 7.8, 7.3, 7, 
    6.4, 7.7, 8, 9, 10.3, 9.4, 10.4, 12.9, 11.3, 11.6, 11.1, 10.3, 9.3, 9.1, 
    8.6, 9.9, 10.6, 11.3, 11.1, 10.7, 12.8, 12.4, 11.1, 12.8, 11.8, 12.1, 
    11.5, 10.8, 10.1, 9.6, 9.7, 9.9, 10, 11.1, 12.3, 11.3, 9.7, 8.7, 8.4, 
    8.3, 9, 9.4, 8.1, 7.2, 7, 5.9, 4.5, 4.8, 4, 3.6, 4, 3.9, 2.7, 1.9, 2, 
    1.8, 1.8, 1.3, 0.6, 0.7, 0.7, 0.8, 1.4, 1.9, 2.6, 4.7, 4.7, 4.7, 5.2, 
    5.6, 6, 4.8, 4.1, 4.1, 4.5, 5.3, 4.7, 5.3, 5.8, 6.1, 6.1, 6.6, 7.1, 7.3, 
    8.7, 7.9, 8.5, 7.8, 8.2, 8.5, 7.7, 7.4, 8.3, 7.3, 8, 8.5, 7.9, 8.1, 7.4, 
    7.1, 7.2, 6.6, 5.5, 4.9, 4.8, 4.3, 2.9, 1.3, 1.4, 1, 2, 2.1, 3.7, 4.7, 
    5.4, 6.8, 6.5, 3.8, 4.5, 5.1, 5.7, 5.7, 5.5, 3.1, 3.1, 3.3, 3.2, 2.5, 
    1.5, 0.4, 0.2, 0.2, 1.4, 1.1, 1.5, 1.4, 2.5, 3.4, 4.4, 4.5, 4.8, 5.1, 
    5.6, 5.8, 5.1, 4.2, 3.3, 3.6, 2.9, 0.9, 0.6, 1.8, 4, 3.9, 3.6, 4.5, 4.2, 
    3.8, 3.4, 5.8, 7, 7.3, 5.8, 7.1, 4, 1.4, 5.1, 5.9, 5, 6.4, 6.3, 4.6, 3.7, 
    1.2, 1.2, 1.6, 0.8, 0.8, 2, 1.8, 2.6, 3, 1.4, 2.1, 2.9, 3.9, 5.1, 5.5, 
    5.9, 5.6, 5.9, 5.2, 5.2, 4.9, 1.1, 2.1, 3.9, 7.2, 6.3, 6.3, 6.1, 5.7, 7, 
    6.6, 7.2, 7.3, 7.4, 5.3, 4.4, 5.3, 5, 6.4, 7.8, 6.6, 5.5, 5.6, 6.9, 6, 
    5.4, 4.9, 5.7, 5.2, 3.6, 3.2, 3.1, 2.2, 0.6, 2.8, 4.2, 5.3, 6.1, 6.6, 
    6.3, 7.4, 8.6, 8.3, 8.2, 9.3, 9.8, 9.5, 9.7, 10.9, 10.2, 11.2, 11.1, 9.8, 
    9.6, 9.6, 8.6, 7.5, 5.9, 5.4, 3.9, 5.2, 4.1, 3.8, 4, 4.6, 1.4, 0.6, 4.5, 
    4.9, 1.4, 2, 0.2, 1.2, 4.6, 0.5, 2.4, 1.5, 1.2, 0.6, 3.6, 4.4, 4.6, 3.9, 
    0.3, 1, 3.3, 1.2, 2, 1.6, 6.2, 6.6, 5.7, 6.6, 6.6, 6, 5.7, 5.9, 5.7, 5.3, 
    4.4, 3.8, 4.6, 5.5, 6.4, 4.8, 6.3, 4.8, 6.3, 5.9, 6.3, 6.6, 4.9, 4.6, 
    3.8, 2.4, 2.5, 2.1, 2.6, 2.3, 2.2, 0.8, 2, 2.4, 3.8, 3.7, 3.6, 3.5, 4, 
    5.1, 5.2, 5.3, 5, 5, 5, 4.8, 4.8, 4.8, 4.2, 3.4, 2.6, 1.2, 0.9, 1.1, 3, 
    4.2, 3.7, 3.7, 3.5, 3.4, 4.5, 3.5, 4, 3, 3.5, 4.1, 4.7, 3.8, 5.2, 4, 4.4, 
    4.3, 3.9, 4.5, 4.4, 4.7, 4.3, 3.5, 3.8, 3.3, 3.5, 3.7, 3.1, 3.6, 4.8, 
    4.1, 3.8, 3.5, 3.4, 3, 2.8, 3.2, 2.8, 2.6, 3.8, 3.4, 4.1, 4.4, 4.3, 3.9, 
    4.6, 4, 4, 3.8, 4.8, 4.8, 4.8, 4.5, 4.1, 4.1, 3.4, 4, 3.6, 2.7, 2.4, 1.8, 
    1.7, 2, 5.5, 6.6, 6, 6.4, 6.5, 6.6, 5.6, 5.7, 5.1, 5, 6, 5.7, 7.1, 6.6, 
    7.1, 6.4, 7.2, 8.5, 8.3, 8.3, 8.9, 6.7, 7.6, 9, 7.2, 6.8, 5.3, 7, 6.5, 
    5.7, 5.7, 4, 4.7, 4.6, 6.2, 5.9, 5.5, 4.4, 5.7, 6.2, 6.9, 5.1, 4.4, 3.5, 
    1.8, 1.5, 2.3, 1.7, 2.1, 1, 1, 0.8, 0.2, 1.2, 0.4, 1.3, 2.1, 2.5, 3, 2.5, 
    3, 2.8, 2.7, 2.5, 2.3, 2.1, 1.9, 3.1, 4.6, 4.5, 2.5, 3, 3.1, 3.2, 3.8, 
    4.5, 4.3, 4.4, 5, 6.1, 6.9, 6.7, 5.9, 5.7, 6, 7.6, 7.5, 6.8, 7, 7.4, 6.9, 
    6.8, 6.7, 6.2, 6.3, 6.1, 6.2, 6.1, 5.8, 5.7, 5.6, 5.8, 6, 6.3, 6.5, 6.4, 
    6.9, 7.2, 7.6, 8.1, 8.3, 8.4, 8.6, 8.6, 8.6, 8.7, 8.8, 8.9, 8.4, 7.9, 
    7.6, 7.3, 7.2, 7.1, 6.8, 6.4, 6.3, 6.1, 6.4, 6.3, 5.8, 5.6, 2.7, 3.1, 
    6.1, 4.5, 3.9, 5.9, 5.7, 5.7, 6, 6.1, 5.7, 5.3, 5, 5, 5, 4.9, 4.8, 5.1, 
    5.2, 5.1, 5.1, 5, 6, 6.8, 3.1, 2.7, 4.5, 4.5, 4.6, 8.9, 10, 10.6, 6.5, 
    11.3, 4.9, 6.2, 5.5, 6.7, 8.2, 7.4, 8.9, 9.1, 9.2, 5.5, 8.1, 7.2, 6.4, 
    7.9, 7.6, 6.8, 5.2, 4.7, 4.8, 7.5, 6.4, 5.7, 5.9, 6.2, 3.9, 3.2, 3.1, 
    2.5, 3.6, 4.8, 5.5, 6.2, 4.1, 4.3, 7.5, 2.8, 4.2, 4.2, 7.4, 6.6, 7.9, 
    7.2, 7.2, 6.2, 6.5, 6, 5.1, 4.7, 5.4, 5.2, 4.5, 3.5, 3.5, 6.6, 6.8, 7.7, 
    8, 7.4, 9.2, 8.9, 8.8, 10, 11, 11.4, 11.4, 11.5, 9.3, 10.4, 12.4, 13, 
    12.7, 12.4, 10.8, 10.8, 10.7, 10.8, 10.8, 10.6, 10.3, 7.1, 4.4, 9.3, 2.4, 
    8.9, 1.9, 8.8, 8.7, 8.5, 8.4, 7.9, 7.5, 7, 6.6, 6.4, 6.3, 6, 5.7, 5.4, 
    5.3, 5.4, 1.9, 1.5, 4.7, 1.4, 1.5, 5.4, 4.3, 3.9, 3.7, 3.1, 2.8, 0.5, 
    1.7, 1.4, 1.9, 1, 1.1, 0.9, 0.7, 0.7, 1, 3.3, 3.1, 2.8, 2.9, 3.3, 3.2, 
    3.3, 3.4, 2.5, 2.6, 3.1, 3.7, 3.1, 2, 3, 2.5, 2.7, 3.3, 2.2, 1.4, 2.6, 
    1.6, 1.6, 1.3, 2.4, 2.5, 2.3, 2.1, 2, 2.8, 0.7, 1.2, 2.1, 2.7, 3.3, 2.8, 
    1.5, 2.7, 2.5, 6.8, 7.6, 7.5, 7.7, 6.4, 6.1, 8.2, 3.9, 4.1, 7.1, 7, 7.1, 
    7.3, 6.2, 5.1, 3.8, 3.5, 3.8, 4, 4.5, 4, 3.9, 4.7, 4.9, 4.3, 4.4, 3.2, 
    4.8, 5.1, 4.3, 4.5, 4.6, 5.1, 5.4, 5.2, 4.7, 5.2, 4.6, 3.6, 2.7, 3.2, 
    2.7, 3.1, 3.7, 5.5, 4.4, 4.5, 4.2, 5.1, 4.3, 4.8, 5.3, 5.9, 6.2, 6.5, 7, 
    7.5, 7.6, 6.6, 5.5, 5.7, 5.7, 8.2, 4.7, 4.3, 3.3, 7.1, 9.1, 5.6, 10, 8, 
    8.8, 6.4, 4.4, 7.4, 3.4, 4.7, 4.8, 6.4, 6.3, 5.8, 8.3, 7.9, 11.3, 9.5, 
    6.8, 7.6, 7.9, 8.3, 5, 5.1, 5.5, 5.7, 8.8, 9.6, 6.7, 6.4, 6.6, 7.4, 7, 
    5.6, 5.7, 6.6, 6.5, 8, 6.6, 6.1, 5.5, 4.2, 3.1, 4.4, 4.8, 5.9, 7.3, 7.7, 
    7.6, 7.9, 6.3, 7.3, 6.8, 6.2, 5.1, 5, 6.4, 5.6, 7, 7.2, 6.7, 6, 7.3, 7.5, 
    6.4, 5.7, 6, 7, 7, 6.1, 8, 7.3, 6.3, 7.4, 5.4, 5.4, 5.7, 9.4, 9.3, 12.5, 
    6.1, 5.6, 7.5, 8.5, 5.2, 4.6, 4.4, 4.2, 4.2, 4.1, 3.9, 3.9, 3.8, 5.8, 
    5.1, 5.4, 5.4, 3.9, 4.7, 4.6, 3.8, 4.1, 4.2, 6, 5.5, 5.6, 6.2, 5.8, 7, 
    5.6, 3.8, 4.4, 4.7, 4.8, 4.8, 4.8, 4.8, 8.2, 7.8, 5.2, 5.3, 8, 8.6, 8, 7, 
    5.2, 8.3, 8.4, 9, 8.6, 5.9, 10, 10.4, 9.4, 9.6, 5.5, 5.8, 11.3, 9, 8.6, 
    7, 7.3, 8.1, 8, 7.9, 7.3, 5.9, 6, 8.4, 8.8, 8.4, 6.3, 7, 7.4, 8.9, 9.2, 
    9.7, 9.5, 9.5, 9.8, 10.3, 10.7, 10.9, 11, 11.3, 11.7, 11.8, 11.4, 11.5, 
    10.9, 10.4, 10.2, 9.4, 9.1, 8.3, 7.8, 8.4, 6.6, 7.8, 7.8, 7.4, 7.1, 6.4, 
    5.9, 4.9, 5.5, 2.9, 2.8, 2.4, 2.3, 2.5, 4.5, 4.7, 2.2, 2.8, 2.5, 2.6, 
    3.2, 3.2, 5.5, 2.4, 5.8, 5.8, 5.8, 6, 6.2, 6.1, 6.1, 6.1, 2.4, 3.1, 2.4, 
    7, 3.1, 2.9, 3.6, 2.6, 7.1, 11.8, 7.1, 7.1, 8.3, 8.6, 9.2, 10, 9.6, 9.1, 
    9.4, 9.1, 4.8, 4.2, 4.3, 6.6, 5.3, 3.2, 2.6, 3.4, 3.3, 2.5, 3.7, 4.6, 
    4.3, 2.2, 1.5, 2.7, 2.7, 2.8, 2, 3.1, 3.5, 3.9, 3.2, 2.7, 2.9, 2, 0.9, 
    0.5, 0.2, 0.1, 0, 1.4, 0, 3, 2, 2.6, 2.2, 3.6, 6.2, 4.7, 4.9, 5.4, 3.3, 
    4.9, 3.7, 4, 3.9, 4.8, 5.3, 6.5, 7.4, 3.5, 3.5, 3.4, 3.8, 5, 9.1, 8.6, 
    10.2, 11.3, 12.9, 13.2, 13.2, 12.9, 13.1, 12.6, 11.4, 6.8, 6.9, 11.6, 
    6.7, 11.8, 11.3, 11.3, 10.6, 11.8, 12.1, 11.6, 7.3, 12, 11.4, 11.4, 11.8, 
    12.1, 12.3, 12.5, 10.9, 10, 9.1, 10.2, 9.7, 10.2, 10.5, 10.1, 10.5, 10.2, 
    8, 8.4, 7.7, 7.9, 8, 7.5, 7.1, 6.6, 6.2, 4.5, 3.1, 2.3, 1.4, 1.4, 0.8, 
    1.4, 2.8, 2.9, 3.1, 2.9, 3.4, 4.5, 2.6, 3.3, 2.7, 8, 3.1, 4.7, 7.5, 7.4, 
    7.8, 9.1, 10.3, 10.1, 9.8, 11, 11.9, 11.2, 12.1, 11.3, 10.2, 9.1, 9.7, 
    8.7, 6.9, 6.1, 4.7, 1.1, 1.9, 3.1, 4.1, 2.9, 4.1, 2.2, 0.9, 0.9, 1.1, 
    2.5, 2.6, 0.5, 4.2, 3, 3.7, 3.1, 6.9, 6.4, 6.3, 7.3, 6.4, 6.8, 6.4, 6.6, 
    7.7, 7, 8.1, 4.9, 4.6, 6.6, 7.3, 7.1, 7.6, 8.2, 8.8, 8.8, 8.8, 9, 9.6, 
    9.9, 11.1, 10.8, 9.2, 9.2, 9.6, 9.2, 10.3, 11.9, 12.1, 10.8, 10.4, 9.5, 
    9.1, 9.6, 9.8, 11.7, 8.9, 6, 7.9, 6.7, 4.6, 4.3, 4.7, 5, 3.8, 3.5, 0.6, 
    3.6, 2.1, 1.1, 2.5, 3.8, 3.9, 4, 4.1, 4.2, 5.1, 4, 3.5, 2.9, 4.4, 4.9, 
    0.7, 1, 1.5, 1, 0.5, 1.1, 2.1, 1.9, 1.5, 2, 1.8, 2.6, 2.3, 2.7, 3.1, 3.5, 
    3.9, 4.3, 4.8, 5.2, 5.6, 6, 6.4, 6.8, 6.1, 5.9, 5.7, 5.6, 4.8, 3.5, 1.9, 
    2.3, 2.5, 2.7, 3, 3.2, 3.4, 3.6, 3.9, 4.1, 4.3, 3.1, 1.7, 1.7, 1.5, 1.2, 
    0.4, 1.2, 0.9, 0.7, 0.4, 0.2, 1, 1.2, 2.1, 3.2, 3.4, 3.7, 3.3, 3.5, 3.9, 
    4.4, 4.3, 4.1, 4.6, 4.7, 5.1, 4.3, 4.5, 4.3, 4.3, 4.1, 5, 5.3, 5.6, 6.2, 
    6.1, 6.2, 6.1, 6.7, 7.5, 7.4, 7.8, 7.8, 8, 7.5, 6.2, 5.9, 6.3, 4.5, 2.5, 
    0.3, 2.2, 4.8, 6.6, 10.1, 13.1, 10.2, 11.3, 11.8, 12.4, 13, 13.3, 17.4, 
    18.1, 17.3, 17.6, 17.6, 15.1, 15.1, 14.2, 13, 13, 12.6, 11.8, 14.9, 13.9, 
    12.8, 13.7, 13.3, 11.6, 8.9, 9.1, 8.3, 9.4, 7.1, 8.1, 8.8, 9.6, 5.8, 3.1, 
    3.7, 5.6, 5.1, 3.5, 3.8, 2.8, 0.7, 2.7, 2.1, 2.9, 5.1, 2.5, 3.3, 5.1, 
    6.1, 6.8, 6.6, 5.8, 5, 6.1, 8.2, 5, 11.4, 12.2, 11.3, 10.2, 10, 10.9, 
    10.8, 11, 7.2, 7.4, 7.8, 8.1, 8.2, 8.1, 11.6, 11.7, 8.4, 7.8, 9, 7.6, 
    8.4, 5.9, 5.4, 6.2, 4.9, 5.7, 5.8, 6.6, 2.9, 1.3, 3.5, 5.5, 5.4, 5.2, 
    5.1, 5.1, 5.1, 4.8, 4.4, 1.4, 1.8, 0.9, 0.2, 0.8, 1.1, 0, 1.2, 3.4, 6.5, 
    5.5, 7, 4, 5.7, 5, 5.2, 5.5, 3.6, 4.2, 5.2, 5.8, 6.2, 5.4, 4.4, 3.4, 2.8, 
    3.1, 3, 3.2, 6.3, 4.2, 2.8, 3.8, 2.1, 1.4, 0.4, 1.1, 3.1, 2, 2.8, 4.2, 
    10.1, 11, 12.4, 12.1, 13.7, 13.5, 14.2, 14.5, 9.6, 9.5, 9.5, 11.7, 13, 
    12.2, 13.2, 13.3, 13.1, 13, 14.4, 14.9, 12, 13.3, 13.5, 14, 12.2, 10.7, 
    11.3, 9.9, 9.7, 8.4, 7.2, 4.5, 4.9, 3.2, 0.4, 1.6, 3.8, 5.9, 7.8, 9.7, 
    10, 11, 9.8, 11.4, 11.4, 11.4, 11.9, 10.2, 10.6, 10.9, 12.3, 11.4, 11.8, 
    8.9, 9.9, 6.9, 5.7, 6.6, 9.8, 8.1, 5.8, 5.2, 4.8, 3.9, 4.4, 4.8, 4.2, 
    3.7, 3.7, 3.6, 2.9, 2.6, 3.2, 2.6, 4.9, 6.3, 7, 9.2, 9.8, 11.2, 10.8, 
    9.5, 9.6, 9.5, 11.5, 10.8, 10.4, 10.9, 9.3, 9.6, 8.8, 8.1, 6.9, 8.4, 8.1, 
    6.6, 7.2, 7.5, 4, 2.9, 4.3, 6.6, 6.1, 5.8, 7.6, 8.5, 9.1, 8.2, 5.7, 4.9, 
    3.8, 7.2, 7.3, 4.9, 5.2, 4.1, 7.3, 6.5, 5.1, 6.2, 6.7, 7.5, 7.5, 6.9, 
    5.9, 7.5, 10, 10, 9.2, 7.7, 5.8, 3.4, 2.4, 9.9, 11.4, 12.6, 9.5, 13.3, 
    12.3, 10.5, 9.4, 8.9, 9.1, 8.7, 8.4, 5, 5.8, 7.2, 4.6, 4.2, 6.4, 5.6, 
    5.5, 4.8, 3.7, 3.6, 3.4, 3.1, 4.5, 5.8, 7.2, 7.7, 7.4, 5.2, 5.4, 4.6, 
    4.7, 4.8, 5.2, 5.8, 6.5, 7.1, 6.4, 8.6, 10.2, 10.7, 7, 6, 5.8, 3.4, 7.7, 
    11.9, 7.1, 9.3, 7.3, 7.4, 5.3, 7.1, 7.5, 6.8, 6.3, 6.6, 7, 7.5, 8, 8.2, 
    7.8, 7.3, 9.5, 7.1, 7.2, 10.1, 9.1, 8.4, 8.9, 6.5, 8.9, 8.7, 8.6, 8, 7.6, 
    7.5, 7.5, 6.8, 6.7, 3.2, 5.7, 5.5, 5.6, 5.5, 5.1, 4.6, 4.2, 3.9, 2.7, 
    4.2, 2.7, 1.4, 0.8, 0.8, 0.4, 0.4, 0.6, 1.3, 3.8, 3.2, 3.7, 5.4, 5.3, 
    6.1, 6.6, 7.4, 5.1, 7.2, 8.6, 8.8, 7.8, 8.3, 10.1, 9.3, 9.8, 9.2, 9.3, 
    9.6, 9, 8, 6.1, 6.6, 5.9, 6.2, 6, 8.5, 7.5, 6.9, 6, 7.1, 9.5, 7.7, 8.3, 
    10.2, 9.8, 6.6, 9, 7.7, 8, 7.6, 6.4, 6.1, 5.4, 5.8, 8, 8.2, 6.1, 6, 6.5, 
    6.4, 6.7, 9.6, 9.2, 7.6, 7.1, 9.1, 8.1, 5.9, 5.7, 6.5, 6.2, 7, 6, 7, 6.7, 
    7.3, 7.1, 7.8, 7.6, 8.2, 8.1, 9, 5.6, 5.1, 5.6, 11.7, 11.3, 10.7, 7.2, 
    7.4, 7.7, 7.6, 9.3, 11.6, 11.9, 12.6, 11.3, 10.3, 6.7, 12.5, 13, 12.7, 
    14.2, 13.8, 12, 10.7, 1.6, 7.9, 7.8, 7.9, 1.4, 4.8, 6.4, 7.5, 9.2, 6.5, 
    7.9, 8.5, 9.1, 11.5, 12.8, 8.9, 8.9, 8.8, 10.3, 8.8, 8.2, 9, 10.3, 9.9, 
    6.6, 8, 10, 9.9, 10.8, 10.7, 10.6, 12.9, 14.1, 10.7, 12.5, 11.6, 11.6, 
    10.7, 10.4, 10.7, 10.7, 10.8, 10.8, 10.7, 12.3, 10.8, 12.1, 10.3, 14, 
    9.7, 11.2, 9.6, 9.7, 10, 8.8, 7.1, 9.6, 9, 7.6, 5.7, 2.7, 3.1, 8.4, 7.6, 
    9.2, 9.1, 7.9, 5.2, 5.4, 4.4, 3.1, 6.6, 6.9, 5.8, 5.3, 6, 5.6, 5.3, 6.7, 
    6.8, 8.2, 6.6, 7.9, 7.5, 7, 7.8, 6.7, 3.9, 5.5, 3.2, 6.3, 4.3, 3.7, 8.3, 
    8.6, 5.9, 8.5, 8.1, 6.5, 8.1, 5.8, 7.6, 2.4, 8.6, 8.9, 9.2, 9.2, 9.3, 
    9.5, 10.8, 10.5, 5.7, 5.7, 5.8, 5.9, 5.3, 4.4, 3.3, 6.7, 3.4, 1.9, 2.4, 
    3.7, 3.8, 5.5, 4.4, 3.4, 3.6, 4.5, 5.2, 10.8, 12.5, 7.9, 15.2, 14.6, 9.5, 
    14.7, 15, 15.7, 15.9, 9.9, 15.3, 10.1, 12.9, 12.2, 8.3, 2.7, 3.3, 2.9, 
    1.5, 0.6, 0.3, 10.2, 10.4, 10.7, 9.3, 8.7, 9.4, 9.9, 10.6, 12.8, 12, 
    10.9, 11.9, 12.7, 11.6, 11.6, 11.5, 11.5, 10.5, 6.6, 5.7, 4.7, 5.4, 5.6, 
    4.5, 3.1, 2.8, 1.1, 1.9, 1.3, 12, 6.3, 16.9, 7, 16.9, 9.2, 17.4, 17.9, 
    17.4, 16.3, 10.7, 10.7, 11, 7.8, 14.1, 10, 7, 7.2, 5.6, 7.2, 6.5, 5, 5.1, 
    4.8, 4.9, 4.9, 5.4, 6.5, 6.5, 5.3, 4.4, 7.4, 7.3, 7.9, 8.4, 8.2, 8.4, 
    12.4, 15.7, 10.7, 9.3, 11.1, 2.7, 1.5, 5.9, 9.7, 8.6, 9.3, 12, 11.7, 
    10.5, 11, 11.1, 11.8, 10.5, 9.1, 8.6, 5.8, 13.6, 14.3, 12.2, 14.9, 15.4, 
    15.6, 15.9, 14.9, 16.7, 15.8, 16.6, 16.4, 19.1, 16.4, 16.7, 16.2, 17.4, 
    14.1, 13, 12.7, 14.2, 14.6, 16.5, 15.7, 13.7, 14, 13.3, 12.9, 14.8, 11.2, 
    10.8, 10.6, 10.8, 10.9, 11.2, 9.7, 8.8, 6.5, 5.1, 6, 5.3, 7.7, 6.2, 7.5, 
    6.3, 7, 7.5, 7.7, 8.5, 6.4, 2.4, 5.9, 6.1, 6, 5.2, 5.8, 5.1, 4.1, 3.9, 
    1.7, 1.6, 1.8, 1.9, 4.9, 5.3, 3.5, 6.6, 7.7, 7.3, 5.1, 5.6, 5.1, 4.8, 
    4.5, 5, 4.5, 4.6, 4.7, 5.5, 5.4, 5.4, 4.7, 4, 2.9, 2.5, 2.3, 5.6, 5.5, 
    2.7, 3.4, 5.3, 6.6, 7.1, 7.6, 7.8, 7.1, 4.3, 5.1, 8.2, 8, 7.4, 7.2, 8.7, 
    8, 8.5, 7.9, 9.1, 8.9, 9.2, 8.7, 10.7, 9.4, 9.7, 9.4, 8.5, 8.4, 10, 9.8, 
    6.8, 6.5, 7.7, 7.4, 7, 8.3, 8.2, 7.4, 7.7, 7.3, 9.8, 8.5, 6.8, 7, 7.3, 
    8.3, 8.1, 7, 5.5, 5.7, 5.7, 5.5, 7.8, 5.2, 4.7, 4.8, 7.9, 9.6, 6, 5.9, 
    8.5, 7.9, 7.4, 6, 9.5, 8.8, 9.2, 7.9, 7.9, 8.1, 3.9, 5.1, 4.3, 3.7, 4.9, 
    8.7, 8, 9.2, 11.1, 7.8, 7.7, 9, 10.7, 12.8, 11.4, 8.4, 10.5, 9.4, 8.6, 
    7.4, 7.6, 7.7, 7.5, 6.5, 7.9, 7.7, 8.2, 7.5, 8.8, 7.2, 6.3, 6.8, 6.8, 
    6.8, 8.4, 9.2, 10.9, 11.1, 11.8, 10.4, 11, 11.2, 9.5, 9.3, 9.8, 7.5, 8.9, 
    6.6, 7.7, 8.4, 8, 8.8, 10.6, 9.8, 10, 10.6, 10.3, 9.3, 8.9, 10.4, 9.4, 
    9.3, 7.1, 6.8, 6.6, 6.5, 6, 5.9, 5.6, 6.2, 3.6, 4.3, 4.1, 3, 3.4, 2.5, 
    2.3, 2.6, 2.1, 2.3, 0.8, 1.3, 1.1, 0.5, 0.8, 2.3, 2.5, 2.2, 1, 1.3, 1.8, 
    2.3, 0.2, 7.1, 11.8, 13.6, 6.8, 8.8, 17.7, 21.6, 23.9, 22.7, 20, 18.5, 
    17.5, 11.5, 10, 11.2, 4, 1.7, 0.2, 2.1, 4.2, 5.2, 4.9, 4.8, 5, 3.3, 3.2, 
    3, 3.8, 6.3, 7.1, 7, 7.1, 6.7, 6.7, 6.4, 5.9, 4.2, 4.3, 3.8, 2.1, 2.9, 
    2.5, 2.6, 2.6, 2.9, 6.5, 6.2, 6.1, 8.3, 8.5, 8.4, 7.4, 10.2, 7.8, 7, 9.1, 
    8.8, 8.8, 6.1, 6.5, 6.9, 5.1, 5, 4.9, 4.9, 4.7, 4.7, 6.6, 5.7, 7.3, 5.8, 
    5.8, 7.7, 7.9, 9.5, 3.4, 3.3, 6.7, 6.4, 5.3, 5.6, 5.5, 3.9, 2.2, 1.2, 
    3.4, 3.2, 4.6, 5.3, 4.9, 4.4, 4.2, 5.1, 4.7, 3.9, 2.8, 5.9, 7.2, 6.5, 
    5.7, 5.7, 5.5, 3.5, 3.6, 3.1, 3.9, 5.3, 5, 5.2, 4.5, 4.4, 4.8, 5.6, 5.7, 
    5.7, 8.4, 9.6, 10, 9.7, 9.4, 9.7, 10.7, 11.5, 7.8, 8.5, 8.7, 9.4, 9.6, 
    8.8, 10, 9.5, 9.3, 10.7, 10.7, 10.1, 11.1, 9.4, 9.7, 10.1, 10.1, 10, 9.9, 
    10.1, 9.5, 9.4, 12.8, 12.5, 12.6, 12.8, 13.2, 12.5, 12.4, 10.5, 8.5, 8, 
    7.4, 9.8, 9.5, 9.8, 9.1, 8.6, 8.3, 8.7, 8.1, 7.3, 7.9, 7.9, 8.8, 12.2, 
    12.5, 13.8, 13.5, 13.8, 13.4, 13.7, 14.3, 10.5, 10.9, 15, 13.4, 12.3, 
    12.6, 12.2, 9.9, 11.5, 12.9, 10.5, 10.7, 10.7, 10.7, 13.1, 11.5, 12.5, 
    12.2, 13.6, 13.9, 14.4, 12.3, 12.7, 13.1, 14.9, 14.1, 14, 14.4, 14.7, 
    13.4, 13.6, 13, 11.1, 10.7, 10.6, 12.9, 11.9, 11.2, 12.1, 12.4, 13, 14.2, 
    13.8, 10.3, 9.9, 13.9, 13.1, 13.3, 12.8, 12.7, 12.2, 12.9, 10.1, 10.5, 
    10.2, 10.6, 9.2, 10.7, 10.9, 14, 13.8, 13.5, 13.7, 13.8, 10.8, 10.9, 
    11.2, 11.7, 15.1, 16.5, 14.8, 14.4, 13.3, 13.8, 16.5, 15.4, 10.8, 10.5, 
    10.1, 10.7, 10.7, 12.3, 12.1, 11.1, 10.9, 10.1, 10, 11, 11.1, 10.9, 10.7, 
    10.4, 8.8, 7.8, 7.6, 7, 6.8, 5.7, 6.8, 7.1, 6.3, 5, 5.5, 5.5, 5.8, 5.8, 
    5.5, 5.5, 5.5, 5.5, 5.5, 5.8, 6.1, 6.2, 6.5, 4.8, 5.3, 5.2, 5.9, 5.4, 
    4.8, 4.7, 5.1, 4.7, 4.1, 4.7, 4, 4.7, 3.2, 4, 3.5, 4.9, 3.5, 4.1, 5.5, 
    6.6, 7.4, 7, 6.9, 4.2, 4.5, 4.9, 3.9, 4.2, 3.2, 3.5, 3.9, 3.7, 4.4, 3.5, 
    0.9, 1.5, 0.7, 1, 1.5, 2.4, 3, 3.1, 3.1, 2.8, 3.3, 3.4, 4.3, 4.2, 3.1, 
    4.1, 4.7, 5.8, 6.3, 6, 5.9, 5.1, 4.5, 4.6, 4, 5.4, 7.6, 6.9, 7.4, 8, 8.2, 
    7.8, 9.4, 9.4, 4.7, 6.8, 7.6, 7.7, 7.4, 11.4, 9, 7.4, 10.2, 6.2, 6.1, 
    6.1, 6.1, 6.4, 6.1, 5.3, 4, 6.1, 4.8, 6.2, 5.8, 6.3, 5.4, 6.2, 7.7, 5.1, 
    3.1, 5.6, 4.7, 5.9, 7.4, 8.3, 8.3, 6.7, 7.5, 9, 9.4, 8.6, 9, 9.1, 11.6, 
    9.6, 6.8, 7, 9, 9.5, 7.9, 9.2, 11.9, 12.1, 11.1, 12.4, 11.6, 12.8, 11.5, 
    10.9, 13.2, 14.4, 15.4, 15.2, 15.5, 14.8, 13.5, 13.6, 7.1, 8.2, 9.6, 7.6, 
    10.5, 10.1, 5.3, 8.9, 6.7, 6.6, 7.8, 6.1, 9.7, 6.5, 7.5, 4.3, 1.9, 2, 
    0.7, 0.9, 1, 3.6, 7.1, 6.7, 7.6, 7.5, 7.5, 7.8, 8.9, 9.8, 9.6, 9.1, 9, 
    8.4, 7.8, 8, 8.2, 6.3, 4.9, 4.1, 2.8, 1.8, 1.8, 1.5, 0.5, 3.3, 8.1, 8.1, 
    8.8, 10, 9.1, 9.1, 9.4, 8.5, 7.2, 8.6, 8, 9.1, 7.2, 6.6, 6.8, 7.2, 7.3, 
    6.2, 5.9, 8.1, 6.6, 5.5, 3.7, 4.3, 4.4, 4.6, 4.6, 4.8, 5.2, 5.6, 4.8, 
    3.7, 3.1, 2.9, 3.7, 2.6, 3.2, 3.4, 1.4, 2.9, 4.4, 5.6, 7, 8.8, 9.9, 7.7, 
    11.1, 12.8, 16.2, 18.1, 18.2, 19, 20.7, 22.2, 25.8, 27.3, 27.3, 23.8, 
    26.2, 26.6, 28.6, 30.5, 30.5, 30.5, 28.9, 30.3, 30.3, 28.6, 28.6, 26.5, 
    26.4, 27.8, 29.7, 27.7, 21.5, 18, 14.1, 14.3, 14, 14, 16, 15.9, 14.8, 
    16.2, 16.5, 12.9, 13.3, 13.8, 14.7, 17.2, 13.9, 15.1, 19.7, 14.2, 13.5, 
    10.5, 9.7, 11.4, 10.1, 9.8, 10.4, 11.4, 10.4, 10.7, 12.9, 10.9, 9.9, 9.5, 
    9.5, 8.3, 9.1, 8.5, 9.1, 8.8, 9.4, 9.7, 9.4, 8.4, 7.8, 8.3, 11, 9.3, 
    11.6, 11.2, 10.6, 8.4, 8.5, 8.5, 10.6, 12.1, 11.8, 10.4, 10.8, 11.8, 8.8, 
    10.4, 7.4, 7.5, 6.8, 7.4, 7.4, 7, 6.8, 6.5, 8.6, 7.6, 5.6, 6.7, 8.9, 9.1, 
    9.6, 7.5, 7.6, 9.3, 11, 10.5, 11.1, 12.8, 14.1, 10.2, 11.2, 11.5, 12.4, 
    12.1, 13.4, 13.5, 13.5, 12.8, 14.3, 15.8, 12.9, 10.4, 13, 14.3, 14.6, 
    13.4, 13.5, 9.7, 9.5, 10.1, 10.2, 14, 13.9, 11.9, 12.6, 10.3, 11.8, 12.8, 
    10.9, 6.5, 6.3, 7.8, 9.8, 12.5, 14.2, 8.8, 6.6, 5.5, 5.1, 6.3, 6.6, 6.1, 
    9, 8.6, 9.3, 10.7, 11.5, 11.7, 12.1, 10.8, 8.8, 5.2, 8.1, 9.8, 7.9, 8.8, 
    7, 8.8, 6.9, 2.7, 1.5, 3, 5.7, 5.3, 7.2, 6.4, 8.2, 9.4, 10.5, 10.2, 10.4, 
    9.1, 8.7, 8.3, 7.3, 3.2, 0.7, 11.8, 11.2, 13.3, 12.2, 12.6, 14.7, 13.4, 
    15, 16, 13.9, 15.9, 16.3, 17, 15.7, 16.9, 17.8, 16.5, 14.4, 13.2, 11.3, 
    10.4, 8.5, 6.7, 4.9, 12, 10.7, 10.1, 11, 10.9, 8.7, 10.4, 10.5, 8.6, 8.1, 
    4.5, 4, 3.8, 3.5, 4.1, 4.7, 4.8, 7.9, 8.4, 9.9, 9, 10.5, 10.2, 13, 14.5, 
    13.3, 14.1, 13.7, 15.6, 15, 14.9, 14.4, 15.2, 16.2, 15.3, 11.6, 8.9, 
    10.2, 11, 9.1, 8.4, 5.5, 5.2, 6.9, 5.2, 7, 5.2, 6.7, 6, 6.8, 4.3, 8.5, 
    12, 10.9, 8.3, 8.3, 7.5, 7.8, 7.9, 8.2, 10.9, 9.2, 7.2, 7.7, 8.7, 8, 8.3, 
    8.1, 9.9, 10.2, 11.1, 9.4, 10, 10.8, 10.7, 6.9, 11.1, 11.5, 8, 6.7, 9.4, 
    9.5, 7.2, 9.5, 10.8, 8.6, 8.3, 8.2, 7.2, 8.1, 7.7, 6.8, 6.8, 6.4, 7.3, 
    8.2, 8.9, 3.7, 5.2, 4.6, 2.5, 6.9, 7.2, 7.5, 6.8, 7.3, 7.7, 8.4, 9.5, 
    12.7, 11.8, 14.2, 14.4, 15.4, 15.6, 16.9, 16.1, 17.2, 16.6, 16.6, 17.6, 
    16.9, 17.5, 17.3, 17.4, 17.4, 16.2, 16.8, 17.6, 17.3, 16.7, 16.5, 15.8, 
    15.5, 15.6, 15.9, 16, 16.7, 15.2, 12, 9.7, 7.4, 6, 6, 4.7, 4.1, 2.3, 1.7, 
    0.5, 0, 1, 3.9, 5.4, 5.3, 6.6, 7.5, 6.8, 1.9, 1.7, 2.9, 3.5, 2, 2.2, 1.7, 
    0.8, 0.4, 2.4, 2.4, 3, 4.8, 3, 2.9, 2.9, 2.4, 1.3, 1.8, 3, 11.8, 14.7, 
    17.9, 14.9, 15.8, 13.2, 10.7, 11.5, 12.8, 13.3, 14, 14.4, 12.7, 15.6, 
    15.2, 15.4, 11.6, 12.2, 10.5, 11.3, 10.9, 10.9, 11.4, 9.8, 9.7, 8.7, 
    10.2, 10.2, 7.6, 7, 4.6, 5, 5.2, 3.3, 2.4, 1.9, 2.6, 7.1, 6.1, 5.5, 7.7, 
    7.5, 9.8, 11.7, 12.3, 12.3, 12.6, 11.6, 11.7, 11.8, 11.3, 10.6, 10.5, 
    10.5, 10.5, 10.6, 8.9, 8.1, 7.8, 7.9, 8.5, 10.3, 11.4, 12.6, 13.8, 13.1, 
    13.3, 14.5, 17.3, 16.4, 16.7, 16.2, 15.4, 14, 13.5, 12.1, 9.6, 9.5, 8.1, 
    7.4, 7.8, 7.9, 7.6, 8.2, 8.4, 7.6, 9.5, 9.9, 10.8, 10.5, 8.3, 9, 7.7, 
    7.3, 5.7, 7.7, 8.6, 7.9, 8, 8.6, 8.9, 9, 9.2, 8, 9.5, 10.5, 8.9, 9.2, 
    10.6, 11, 11.7, 13.6, 14, 16.4, 18.3, 17.1, 17.6, 18.1, 17.9, 17.5, 17.9, 
    19.3, 18.7, 19.7, 19.5, 18.2, 17.1, 14.6, 14, 15.6, 16.2, 10.5, 10.4, 
    8.4, 7.8, 5.4, 0.1, 2.8, 1.4, 4.4, 6.6, 7.3, 8.1, 9.5, 10.7, 11.9, 11.6, 
    10.6, 11.4, 10.9, 11.2, 11.2, 22, 10.9, 11.4, 11.3, 11.6, 11.6, 12.3, 
    11.7, 11.6, 11.4, 12.1, 12, 11.2, 10.4, 10.6, 11.5, 12.4, 12.2, 11.7, 
    11.1, 10.2, 10.4, 11.4, 10.5, 10.4, 10.3, 10.5, 11.9, 11.6, 12.4, 12.4, 
    13.1, 13.4, 14.1, 14.1, 14.5, 14.2, 14.1, 17.5, 15.6, 17, 17.5, 18.1, 
    18.9, 21.2, 19.4, 17.5, 14.7, 14.8, 14.5, 15, 15, 17.8, 19.5, 19.6, 18.5, 
    17, 17.3, 20.1, 22.4, 19.9, 17.8, 11.5, 18, 13.2, 14.6, 11.6, 13.7, 12.7, 
    15.2, 17.2, 21.7, 19.9, 14.3, 16.4, 14.9, 14.4, 13.1, 7.4, 9.1, 15.8, 
    13.4, 13.8, 13.7, 12.7, 12.8, 12.4, 12.4, 11.7, 11.8, 11.3, 7.7, 2.4, 
    7.7, 6.4, 10.3, 6.3, 7.1, 10.1, 6.9, 7.7, 7.6, 10.3, 9.8, 8.5, 7, 8.6, 8, 
    7.5, 6.6, 7.3, 6.9, 8.2, 10.9, 11.4, 10, 9.2, 8.2, 4.7, 6.7, 1.7, 2.2, 2, 
    1.7, 2.1, 0, 6.7, 5, 6.7, 6.4, 6.7, 6.5, 7, 7.3, 8.4, 14.1, 10, 9.9, 9.9, 
    11.9, 14, 17.4, 18.5, 17.1, 19, 20.1, 19.6, 22.4, 21, 27.5, 22.8, 21.6, 
    21.7, 21.6, 23.1, 23.4, 23.7, 24.3, 22.8, 23.8, 26, 22.9, 21.4, 20.5, 
    19.7, 19, 19.5, 19.7, 19.7, 21.9, 23.1, 24.5, 24.3, 26.6, 25.1, 17.2, 
    16.2, 17.8, 18.5, 18, 16.3, 18.7, 19, 17.8, 16.6, 15.8, 15.2, 15.1, 15.3, 
    14.1, 12.6, 14.4, 12.6, 6.6, 11.5, 8.9, 8.8, 9, 7, 10.5, 11.1, 12.6, 16, 
    12.9, 13.9, 12.7, 12.9, 13.3, 10.7, 10.6, 10.8, 10.2, 9.9, 9.5, 7.4, 5.6, 
    3.4, 3.5, 5.2, 8.7, 9.4, 8.2, 8.5, 7.8, 6.9, 5.6, 4, 5.1, 6.7, 6.4, 6, 
    6.7, 7.7, 6.4, 6.2, 6.4, 5.4, 6, 5.8, 5.9, 8, 8.6, 7.6, 7.3, 7.2, 6.4, 
    7.2, 8.4, 8.7, 7.6, 8.4, 7.7, 9.2, 9.2, 9.5, 9.5, 10.1, 10.4, 12, 11.8, 
    12.7, 11.1, 12.1, 13.1, 15, 16.4, 19.1, 19.8, 19.3, 19.3, 19.7, 19.5, 
    19.3, 20.9, 23.3, 24.4, 23.5, 22.9, 22.4, 20.9, 20.5, 19.1, 15.5, 14.1, 
    13.3, 13.2, 11.2, 10.8, 11.8, 10.6, 10.6, 8, 6.5, 5.9, 7.6, 6.6, 6.5, 
    6.6, 7.1, 5.1, 4.9, 4.8, 5.9, 7, 7.4, 7.8, 8.6, 8.9, 9.7, 10.6, 10.6, 
    9.7, 10.7, 11.2, 10.6, 11.1, 10.9, 9.9, 9.4, 10.8, 11.2, 12.2, 9.5, 9.2, 
    8.7, 8.9, 7.4, 6.7, 6.1, 3.7, 4.9, 4.9, 5.7, 5.8, 4.3, 3.7, 5.4, 5.3, 
    6.2, 7.5, 7.3, 6, 6.3, 6.6, 6.8, 5.4, 6.9, 6.7, 7.8, 10.1, 15.6, 15, 
    12.4, 11.9, 9.2, 10.6, 10.4, 10.8, 10.6, 11.3, 12.8, 11.6, 11, 11, 11.8, 
    11.8, 11.6, 13.4, 14.7, 15.5, 16.2, 15.6, 14.8, 13.8, 13.8, 13.6, 14, 
    15.7, 16.6, 16.9, 17.2, 16.2, 14.1, 12.7, 9.8, 7, 8.4, 8.3, 10.1, 8.3, 
    9.2, 10.3, 10.9, 9.2, 8.5, 8.1, 9.4, 8.6, 6.3, 5.6, 4.7, 3.2, 4.6, 5.6, 
    5.7, 7.5, 7, 7.2, 7.6, 6.3, 7.9, 8.4, 11.2, 12.9, 14.7, 13.6, 6.7, 6.1, 
    7, 6.5, 2, 3.5, 2, 2.7, 2.9, 5.8, 5, 3.6, 4.6, 2.8, 0.2, 3.2, 3, 2.3, 
    2.5, 1.7, 1, 2.6, 2.9, 0.8, 0.9, 2.6, 0.7, 4.4, 3.7, 2.3, 2.1, 2.4, 2.6, 
    1.8, 1.4, 0.1, 4.6, 3.5, 3.3, 0.1, 1.4, 6.6, 6.9, 9.4, 7.6, 7.2, 8, 9.2, 
    8.4, 8, 7.7, 4, 6.4, 4.3, 7.2, 6.2, 10.9, 9.5, 8, 8.5, 8.7, 9.6, 10.3, 
    12.5, 11.4, 10.7, 9.4, 10.3, 11.6, 11.9, 11.4, 10.1, 10.9, 11.2, 10.9, 
    12, 11.1, 10.7, 10.8, 9.4, 10.8, 10.2, 12.1, 11.5, 11.4, 11.8, 8, 7.9, 
    9.2, 9.5, 9.4, 9.6, 10.5, 11.2, 9.4, 8.2, 7.1, 7.3, 10.4, 6, 6.9, 6.8, 
    5.1, 4.5, 7.2, 9.5, 8.2, 7.3, 9.2, 8.8, 9.6, 12, 10.7, 11.2, 10.9, 8.1, 
    9.8, 13.3, 10.4, 9.6, 3.7, 6.3, 9.5, 8.8, 10.2, 10.3, 7.4, 8.2, 9, 10.5, 
    10.1, 12.6, 12.2, 7.9, 7.1, 8.2, 8.4, 9.7, 7.6, 6.9, 6.9, 5, 5, 8.7, 8.2, 
    6.3, 6.1, 5.4, 6.2, 6.6, 8.4, 4.6, 3.7, 7.1, 7.9, 8.6, 6, 6.4, 6.1, 3.9, 
    6, 7.5, 8.6, 5.9, 8.4, 8.4, 9.3, 7.8, 9.7, 8.7, 9.9, 11.2, 9.1, 8.1, 8.2, 
    10.5, 10.6, 10.6, 10.6, 8.5, 10.2, 7.3, 10, 10, 10.6, 11, 10, 8, 7.4, 
    9.8, 8, 9.3, 8.5, 7.8, 8, 8.3, 7.5, 8.1, 8.7, 8.4, 10.8, 7.3, 6.6, 11.4, 
    10.7, 10.5, 11.7, 12, 11.8, 10.9, 11.1, 8.9, 7.5, 7.1, 9, 8.9, 11.3, 
    11.8, 11.3, 11.5, 11.9, 12.1, 9.5, 9.4, 8.6, 8.1, 10.6, 11.3, 12.5, 12.1, 
    11.8, 10.2, 10.5, 9.8, 8.7, 8.1, 9.1, 10.1, 8.8, 7.5, 8.1, 8.9, 7.3, 9.2, 
    9.2, 11.1, 9.7, 8.2, 9.8, 6.3, 7.7, 6.6, 8.3, 7.9, 4.2, 6.3, 2.4, 3.6, 
    0.6, 3, 4.6, 5.3, 6.8, 7.6, 7.8, 7.7, 8.2, 9.9, 13.4, 13.5, 13.4, 14.3, 
    13.5, 15, 17.4, 18.3, 19.4, 17.5, 18.6, 17.9, 17.9, 17.4, 18.4, 21.4, 
    18.2, 18.2, 23.7, 25.9, 25.2, 24.9, 25, 24.2, 23.7, 24.5, 23.8, 25.2, 
    23.9, 22.3, 22.3, 21.5, 20, 20.4, 22, 24.8, 25.3, 25.5, 26.1, 24, 22.9, 
    22.1, 22.4, 20.5, 21.4, 20.3, 18.7, 17.9, 16.6, 14.5, 13.6, 12.8, 11.2, 
    11.5, 14.1, 16.9, 17, 14.5, 14.8, 15, 15.4, 13.5, 14.6, 19.2, 14.6, 17.9, 
    19.1, 18.7, 19.1, 17.6, 15.5, 15.9, 15.3, 15.2, 17.5, 17.8, 17.1, 16.7, 
    17.6, 17.8, 15.8, 15.2, 15.3, 15.1, 15, 14.1, 14.1, 15.7, 15.3, 14.4, 
    16.6, 18.3, 17.4, 17.6, 18.1, 17, 16.1, 16.8, 16.5, 16.2, 16.7, 16.5, 
    16.2, 17.3, 17.8, 18, 16.8, 16.2, 15.4, 16.2, 16.9, 17.2, 16.9, 17.8, 
    17.6, 17.7, 17.3, 18.3, 18, 18, 17.7, 17.5, 19.1, 20.9, 20.8, 20.8, 19.9, 
    18.9, 18.6, 18.3, 17.4, 17.3, 17.6, 17.1, 16.4, 15.4, 14.2, 13.3, 13.1, 
    12.5, 11.9, 12.1, 11.2, 10.1, 9.9, 10.1, 10.4, 9.8, 11.1, 9.5, 10.4, 10, 
    8.5, 8.9, 9.5, 11.2, 11.1, 10.9, 9.6, 9.7, 9.9, 10.2, 11.7, 11, 11.2, 
    10.9, 10, 11.8, 11, 10, 10.5, 9.5, 8.6, 9.2, 9.3, 8.1, 7.6, 7.5, 7.6, 
    6.8, 5.4, 4.2, 2.2, 2.3, 0.1, 2.5, 4.9, 5.3, 8.1, 3.6, 4.2, 7.1, 8.3, 
    7.3, 7.5, 6.6, 4.9, 3.8, 3.4, 3.4, 4, 4.3, 4.6, 3.9, 1.9, 3, 4.8, 4.9, 
    4.6, 6.1, 6.3, 7.5, 9.2, 9.7, 11.9, 13, 12.5, 12.4, 14.3, 14.6, 15.1, 
    14.7, 13.8, 15.9, 16, 14.6, 15.1, 14.3, 14, 13.3, 13, 13.9, 15.2, 14.2, 
    14.3, 15.1, 15.9, 15.8, 16.7, 16.5, 16.1, 18.6, 18.5, 18.4, 19.3, 18.8, 
    18.9, 17.9, 16.9, 15.4, 12.8, 7.5, 6.3, 4.3, 4.1, 4.1, 2, 1, 0.4, 1.8, 
    0.6, 2.4, 1.4, 1.2, 4.9, 5.6, 6.6, 7.6, 7.3, 8.6, 8.1, 8, 9.1, 8.1, 8, 9, 
    9.3, 9.8, 9.7, 10.5, 8.4, 9.2, 9.1, 9.1, 8.2, 7.9, 7.2, 6.8, 6.8, 6.4, 
    5.9, 5.4, 4.7, 4.7, 4.6, 4.2, 3.7, 3.4, 4.5, 3.1, 2.2, 1.7, 3.6, 7.4, 
    10.4, 13.9, 15.9, 15.6, 16.1, 17.2, 17.3, 17.9, 17, 16.9, 16.4, 14.1, 
    14.1, 14.9, 15.4, 12.4, 11.8, 12, 11.4, 14, 13.1, 11, 10.4, 8.8, 5.6, 
    6.6, 7.6, 7.8, 7, 6.5, 6, 5.5, 5.8, 4.8, 4.5, 4.9, 5.2, 4.5, 4.2, 3.9, 
    3.3, 2.4, 1.7, 1.6, 0.4, 0.2, 2, 1.3, 0.8, 0.2, 2.3, 4.1, 4.5, 3.5, 4.6, 
    5.6, 8.1, 7.5, 3.4, 2.8, 8.7, 4.4, 11.1, 11.3, 10.5, 12.9, 13.6, 12.7, 
    11.1, 10.3, 2.5, 9.5, 5.5, 6.1, 9.4, 9.9, 10.3, 9.9, 8.7, 8.9, 8.5, 1.4, 
    3.5, 2.4, 1.7, 7.1, 4.1, 1.9, 9.5, 10.5, 9.9, 7.3, 7.9, 6.1, 8.9, 8.1, 
    8.6, 9, 9.7, 9.2, 9.1, 0.8, 0.4, 0.7, 0.9, 0.4, 0.7, 0.3, 0.6, 0.9, 0.4, 
    1.6, 0.6, 1.5, 1.4, 1.9, 0.9, 1.3, 1.5, 0.2, 0, 0.9, 0.5, 0.6, 1, 2.1, 
    2.1, 0.1, 4.9, 2.1, 1.6, 4.4, 4.5, 5.2, 2.4, 3, 6.9, 4.5, 5.2, 5.5, 3.8, 
    3.5, 6, 6.9, 8.4, 7.9, 2.9, 1.8, 2.7, 7.9, 2.6, 7.2, 7.4, 7.4, 1.5, 2.1, 
    4.3, 3.9, 6.7, 4.4, 6.4, 8.6, 8.8, 8.6, 7.6, 5.8, 5.3, 4.8, 6.8, 7.9, 
    7.1, 5.2, 5.3, 5.3, 3, 2.7, 2.2, 2.9, 2.7, 0.9, 1, 1.6, 2.6, 4.3, 4.7, 
    5.4, 6.3, 6.8, 4.6, 4.2, 8.1, 6.3, 3.2, 4.1, 3.2, 3.4, 2.5, 3.6, 3.6, 
    3.6, 7.2, 6.1, 9.4, 9.2, 8.7, 8.1, 6.5, 6, 5.1, 2.5, 2.8, 2.1, 3.2, 6, 9, 
    10, 10.9, 11.7, 12.4, 12.6, 13, 12.8, 12.7, 13.6, 12.2, 12.2, 12.6, 13.7, 
    14.3, 11.5, 11.6, 10.2, 4.1, 6.3, 3.9, 0.7, 1.6, 4.1, 1.4, 3, 0.3, 4.3, 
    4.4, 8.6, 10.8, 10.5, 13.9, 12.6, 10.5, 2, 2.8, 4, 11.9, 1.7, 5.8, 8.9, 
    11.8, 11.3, 10.9, 11, 11.5, 12.3, 11.7, 12.3, 12.2, 13.2, 13, 12.7, 12.2, 
    12.4, 12.5, 11.7, 11.5, 12.5, 11.7, 11.6, 10.7, 11.6, 13.6, 13.3, 14.9, 
    12.1, 9, 5, 3.4, 4.9, 4.4, 5.6, 4, 3, 3.9, 2.6, 3.3, 3.7, 5.8, 6.6, 6.6, 
    3.5, 4.3, 5.8, 5.2, 7.7, 4.6, 6, 8.3, 7.2, 7.9, 9, 7.8, 4.7, 4.3, 5.2, 
    3.5, 2.4, 1.3, 2.7, 2.4, 0.9, 1.1, 3.6, 6.1, 1.9, 3.1, 0.7, 0.9, 1.9, 
    2.5, 3.6, 4.8, 5, 7.9, 8.8, 5.7, 7.1, 7.5, 7.4, 8.6, 8.6, 6.2, 4.6, 4.6, 
    0.9, 1.5, 2.9, 0.6, 0, 3.4, 3.2, 0.9, 4.1, 1.9, 0.9, 3.8, 3, 7.9, 3.3, 
    3.2, 3.5, 5, 4, 2, 1.8, 1.8, 2.1, 12.9, 5.9, 8.2, 13.8, 15.1, 13.2, 16.3, 
    16.2, 14.7, 14.7, 13.7, 11.1, 12.3, 13.8, 14, 13.9, 13.3, 12.3, 13.6, 
    13.1, 11.8, 12.2, 14.5, 14.7, 14, 2.2, 2.2, 2, 1.7, 3.8, 3.1, 1.6, 1.8, 
    1.4, 1.8, 3.3, 1.4, 1.8, 2.7, 3, 1.1, 0.8, 1, 1.9, 1.3, 8.8, 8.3, 7.9, 8, 
    9.1, 4.5, 7.3, 2.7, 3, 2.5, 1.2, 5.8, 2.9, 6, 5.9, 6, 1.9, 1, 4.2, 8.2, 
    7.3, 7.6, 6.6, 11.3, 9, 9.3, 9.5, 11, 10.8, 10.8, 11.1, 5.5, 0.7, 4.8, 
    4.8, 8.3, 5.6, 2.6, 3.6, 7.5, 0.3, 3, 6, 7.7, 6.1, 6.2, 4.6, 5.9, 5.4, 
    6.1, 4.6, 4.8, 4.5, 4.5, 4.3, 4.8, 5.9, 3.6, 4.4, 4.2, 3.1, 4.9, 5.1, 
    3.8, 3, 3.2, 3.3, 3.3, 3.7, 4.7, 4.8, 3.7, 4.6, 3.5, 3.5, 4.2, 4.3, 3.2, 
    3.9, 3.9, 3.9, 3.9, 4, 4.1, 4.3, 3.3, 2.5, 2.3, 2.3, 0.9, 0.4, 2.4, 0.7, 
    1.1, 1.6, 1.5, 2.4, 1.5, 1.4, 0.8, 1.2, 0.9, 0.7, 0.6, 1.2, 1.6, 1.9, 
    2.6, 2, 8.7, 9.5, 9.6, 10.2, 8.5, 11, 10.3, 10.9, 9.7, 9.8, 11.4, 9.8, 
    10.9, 10.4, 12, 11.8, 11.6, 10.9, 10.3, 11.9, 12.3, 11.5, 11.1, 6.6, 
    12.7, 13.3, 12.2, 16, 16.5, 16.1, 16.1, 14.8, 13.1, 15.2, 15.5, 16.3, 
    15.3, 14.8, 14.4, 14.5, 12.8, 14, 15.7, 15.3, 13.2, 13.1, 13.5, 13.7, 
    13.5, 13.9, 14, 14.6, 13.5, 13.5, 5.3, 5.7, 13.1, 14.2, 14.3, 13.6, 15, 
    16.1, 16.9, 16.4, 17.4, 17.5, 18.1, 16.5, 15.7, 14, 13.1, 10.7, 10.4, 
    11.1, 12.3, 11.7, 12.5, 13.4, 14, 14.6, 13.8, 13.4, 14.7, 13.2, 14.6, 
    15.8, 16, 16.7, 17.5, 17.8, 17.8, 18.5, 18.6, 18.4, 21.3, 20, 20.4, 20, 
    20.1, 19.6, 19.7, 19.9, 20, 21.4, 23.1, 22.3, 22.2, 21.6, 22.4, 19.8, 
    20.4, 20.7, 15, 12.8, 12.1, 9.1, 10.5, 8.4, 7.8, 6.9, 6, 9.3, 9.6, 10, 
    8.9, 11.2, 11.7, 13.5, 13.5, 13.9, 14.5, 13.7, 13.4, 14.1, 11.8, 14.9, 
    15.2, 13.8, 13.3, 17.5, 13.4, 17, 16.9, 17.5, 13.4, 17, 13, 15.9, 16, 
    15.2, 14.2, 15.1, 7, 15, 13.1, 6.5, 6.2, 6.2, 4.8, 9.7, 11, 8.8, 9.5, 
    0.8, 10.5, 12.2, 10.8, 11.6, 12.2, 12, 12.4, 10.9, 11.6, 12.8, 12.5, 
    11.9, 13.9, 13.7, 13.6, 14.8, 13.6, 15.1, 14.2, 14.3, 12.9, 12.9, 13.2, 
    13.3, 13.5, 14.6, 14.3, 12.7, 15.3, 16.3, 16.1, 15.7, 14.5, 14.8, 13.5, 
    12.6, 12.3, 9.8, 9.8, 10.3, 9.7, 9.3, 8.9, 8.5, 7.8, 7.9, 6.9, 5.6, 6.4, 
    6.4, 7.6, 7.3, 6.8, 6.6, 6.9, 7.1, 5.7, 6.4, 6.4, 5.9, 5, 5.2, 6.2, 6, 
    4.8, 3.4, 4.1, 2.6, 1.8, 2.2, 4.8, 4.7, 3.6, 2.7, 3.1, 2.1, 3.5, 3.7, 
    2.8, 2.9, 2.6, 2, 2.7, 2.4, 2.8, 2.4, 2.7, 3.8, 3.8, 0.2, 3.1, 3.1, 1.8, 
    1.6, 2.4, 5.2, 5.9, 3.8, 1.5, 6.7, 7.3, 8, 7.5, 7.5, 7.1, 7.1, 7, 7.3, 
    8.2, 7.3, 7.7, 9.3, 9.1, 9.1, 8.2, 1.9, 2.8, 2, 1.2, 0.1, 0.6, 1.7, 0.6, 
    1.3, 1, 2.2, 3.7, 5, 1.9, 1.8, 1.2, 2.3, 2.6, 0.8, 3.6, 7.9, 6.5, 6.2, 
    9.4, 9.4, 7.6, 8.5, 7.5, 9, 9.7, 9.2, 9, 8, 6.7, 5.7, 7.2, 6.1, 7.3, 7.3, 
    5.7, 4, 2.4, 1.1, 1.3, 3.6, 4.4, 2.8, 2.5, 3.3, 4.2, 3.7, 1.6, 1.4, 1.1, 
    5.2, 7.2, 8.5, 9.9, 8.3, 8.6, 7.7, 7.5, 9.1, 5.7, 4.5, 4.1, 4.2, 5.6, 
    7.3, 9.2, 10.8, 10.9, 14.8, 16.4, 19.8, 21.8, 23.7, 25.3, 25.8, 25.1, 
    27.2, 28.1, 28.7, 27.4, 27, 25, 22.5, 20.7, 19.2, 17.4, 12.1, 7.8, 7.1, 
    7.7, 8.6, 8.6, 9.2, 8.5, 8.2, 7, 6.7, 3.9, 4, 3.8, 6.6, 7, 4, 4.5, 4.5, 
    4, 1.4, 2.2, 1.5, 2.5, 5.4, 4.3, 6.2, 5.1, 5.3, 11.2, 11.7, 10.9, 1.7, 
    0.5, 1, 3.6, 4.2, 1.3, 7.4, 9.8, 9.3, 8.8, 10.6, 13.3, 14.5, 13.9, 11.7, 
    12.5, 12.5, 13.7, 14.5, 13.9, 15.1, 15.5, 16.5, 15.8, 13.5, 13.3, 13.4, 
    13.7, 12.5, 11, 11.8, 12.8, 12.3, 12.2, 11, 10.2, 9.8, 10.1, 11.2, 11.9, 
    10.7, 11.2, 11.3, 9.7, 9.4, 10.2, 11.6, 11.6, 11.3, 10.7, 9.7, 10.4, 
    10.8, 9, 7.6, 6.7, 6.4, 5.4, 7.7, 6.9, 7.4, 8.6, 8, 7.3, 7.3, 6.8, 5.7, 
    7.9, 5.1, 7.6, 6, 5.3, 4.8, 6, 5.3, 3.9, 2.6, 5.4, 2.8, 4.4, 1.8, 3.9, 
    9.5, 9.4, 9.1, 9.3, 6.3, 5.5, 4.1, 4.2, 4.2, 3.9, 3.8, 2.1, 1.3, 0.8, 3, 
    2.1, 4.3, 3.6, 0.8, 0.3, 0.4, 0.8, 1.5, 1.8, 2.3, 3.5, 5.5, 6.3, 6.6, 
    7.4, 5.4, 7.7, 11.6, 13, 12, 10.7, 11.6, 9.8, 7.9, 7.3, 5.1, 5.5, 6.2, 
    3.2, 3.1, 6.1, 2.1, 1.5, 4.4, 3.2, 3.4, 1.8, 2.2, 2.1, 2, 2.1, 1.7, 2.7, 
    2.2, 2.9, 3, 4.2, 3.7, 5.2, 6.9, 6.9, 7.1, 7.9, 7.5, 7.2, 6.7, 7.6, 7.3, 
    7.1, 8.4, 1.1, 2.7, 4.7, 8.8, 1.6, 1.3, 1.9, 1, 0.9, 0.8, 1.4, 1.2, 2.6, 
    0.4, 1.2, 7.8, 5, 16.9, 16.5, 16.1, 14.5, 14.1, 14.2, 14, 14.7, 14.8, 
    14.4, 14.1, 13.2, 10.7, 14.2, 13.6, 14.2, 12.6, 12.6, 13.4, 14.8, 15, 
    15.7, 16, 17.4, 15.2, 14.5, 12.3, 3.3, 1.9, 2.7, 2.2, 3.2, 5.8, 6.6, 7.7, 
    8.4, 6.8, 7.8, 8.4, 9.9, 12.1, 12, 13.1, 13.4, 13.2, 14, 13.8, 12, 10.5, 
    12, 12.3, 14.4, 13.1, 11.4, 11.3, 8, 9.7, 9.7, 8.1, 8.8, 9.6, 7.7, 6.3, 
    6.6, 7.4, 5.6, 5.5, 2.7, 5.6, 4, 3.8, 2.2, 0.9, 0.7, 0.7, 3.8, 4.2, 3.6, 
    0.9, 1.5, 1.8, 2.2, 0.3, 0.3, 0.5, 0.4, 1.9, 2, 1, 1.3, 0.4, 2.2, 0.7, 
    2.2, 0.9, 5.4, 7.3, 6.7, 4.9, 6.8, 10.4, 9.6, 2.7, 11.4, 10.1, 10, 15.6, 
    15.5, 15.8, 14.7, 13.5, 13, 13.7, 14.5, 15, 14.9, 14.7, 16.4, 16.6, 16.8, 
    17.4, 17.6, 18.1, 18, 18.3, 17.8, 17.3, 17.9, 18.6, 18.2, 18.1, 18.7, 
    18.6, 19.4, 21, 22.5, 23.2, 22.2, 26.3, 25.1, 24.4, 24.2, 24.1, 22.7, 
    24.9, 25.3, 24.3, 23.1, 21.8, 22.2, 22.4, 23.3, 23.2, 23.2, 21.3, 21.6, 
    20.7, 20.8, 18.5, 17.5, 16.2, 16.4, 15.7, 15.1, 14.1, 14.3, 14.2, 13.4, 
    12.5, 8.9, 8.6, 8.2, 8.4, 8.6, 9.2, 8.4, 7.5, 6.6, 6.2, 5.8, 5.5, 5.4, 
    6.2, 6.6, 6.6, 6.8, 8.5, 8.5, 8.5, 7.9, 7.4, 7, 6.6, 6, 8.3, 7.2, 7.4, 
    8.1, 7.6, 7.2, 7.1, 7.2, 6, 6.9, 6.5, 8, 7.4, 7.9, 8.2, 8.3, 6.6, 6.3, 
    5.9, 4.9, 4.7, 5.1, 4.8, 4.2, 4.3, 4.5, 4.3, 4.6, 4.6, 4.2, 4.8, 5.8, 
    6.6, 6.9, 7.1, 7.7, 7.7, 8.4, 8.6, 8.8, 8.7, 9.4, 9.3, 9.5, 10.2, 10.6, 
    10.3, 9.6, 10.3, 10, 8.5, 9.7, 8.4, 8.6, 9.5, 9.3, 9.5, 8.4, 8.5, 7.8, 
    7.9, 8.5, 9, 10.1, 8, 8.2, 9, 10, 10.8, 12.1, 13, 13.3, 13.9, 14.8, 15.5, 
    15.4, 15.8, 15.7, 14.4, 11.4, 9.7, 8.5, 8.1, 8, 7.1, 7.7, 7.3, 7.6, 8.9, 
    9, 9.9, 9.6, 9.9, 9.9, 10.7, 10.8, 10.4, 10.3, 10.7, 10.5, 10.5, 10.1, 
    9.4, 9, 7.8, 6.7, 5.7, 5.1, 5.3, 5.5, 5.9, 7.7, 5.7, 5.9, 5.9, 5.9, 5.5, 
    4.4, 3.4, 3.8, 4.2, 3.7, 2.8, 3.4, 3.7, 3.8, 4.4, 4.6, 4.6, 4.3, 4.5, 
    4.5, 4.9, 5.6, 6.9, 8.6, 9.8, 10.8, 9.5, 8.5, 10, 11.1, 11.3, 11.9, 12.5, 
    12.2, 11.8, 9.2, 9.3, 10.7, 11, 11.1, 11.8, 12, 11.5, 11, 11.3, 11.6, 
    11.1, 11.5, 12.2, 12.1, 11.6, 11.5, 11.4, 11.4, 10.8, 10.2, 9.2, 8.6, 
    7.9, 7.3, 6.6, 5.8, 5.2, 4.5, 3.7, 2.6, 1.5, 2.9, 4.2, 4.9, 5.7, 5, 5.8, 
    6.4, 7.1, 8.2, 9, 8.9, 8.8, 8.9, 8.4, 7.3, 6.6, 6.6, 5.6, 5, 4.1, 3.6, 
    3.2, 2.9, 3.2, 3.6, 4.1, 4.6, 4.8, 3.9, 4, 4.2, 4.5, 4.6, 4.2, 4, 2.9, 
    2.9, 2.7, 2.3, 2.1, 3.6, 3.8, 2.7, 5.1, 8.2, 7.3, 7.6, 8, 6.5, 6.8, 6, 
    4.2, 5.1, 5.9, 7.2, 7.4, 9.6, 10.6, 11.9, 14.6, 17.2, 17.2, 15, 12.7, 
    12.9, 11.8, 15.1, 14.3, 11.5, 9.8, 11, 13.5, 13.4, 12.8, 12.1, 11.8, 7, 
    7.8, 4.7, 4, 11.4, 8.4, 10.2, 11.4, 11.3, 13, 14.1, 15, 16.9, 22.8, 23.1, 
    23, 22.7, 22.5, 22.2, 21.7, 21.3, 20.7, 19.7, 18.9, 18.7, 17.2, 15.3, 
    13.9, 13.2, 12.8, 11.9, 10.9, 10.4, 9.3, 8.7, 8.9, 7.6, 7.3, 7.3, 8, 8.4, 
    8.5, 8.6, 8.4, 6.9, 7.5, 5.8, 7.1, 7.3, 6.9, 7.1, 6, 7.1, 5.6, 5.6, 4.8, 
    6.3, 6.5, 5.5, 5.2, 6.2, 5, 6, 5.7, 5.9, 7.1, 8.1, 10.2, 10.8, 7.5, 10.1, 
    9.2, 8.6, 8.5, 6.5, 8.8, 9.2, 9.4, 8.1, 6.8, 8.9, 9.5, 10.5, 10.1, 9, 
    8.2, 9.1, 8.8, 9.2, 10.7, 10.9, 10.1, 10.6, 12.7, 12.1, 12.6, 12.5, 11.6, 
    9.8, 10.7, 10.5, 13.2, 13.9, 13.1, 12.6, 13.5, 12.6, 12.4, 14.1, 13.8, 
    13.7, 11.8, 11.1, 11.5, 10.1, 9.8, 12.2, 13.3, 13.4, 12.3, 12.2, 12.2, 
    10.5, 10.6, 10.8, 9.4, 9.3, 8.6, 7.6, 7.6, 6.7, 8.6, 8.5, 8.4, 8, 8, 8.3, 
    7.7, 6, 6.1, 5.3, 5.3, 5.1, 5.8, 4.6, 5.5, 5.8, 5.1, 2.3, 4.4, 4.1, 5.3, 
    2.7, 7.5, 2.5, 2.9, 7.8, 7.2, 2.3, 0.4, 0.8, 2.6, 3.4, 3.9, 4.8, 3.2, 
    5.6, 4.8, 3.7, 5.6, 7.5, 4.3, 4.2, 4.5, 4.9, 8.1, 8.9, 6, 9.9, 6, 8.7, 
    11.7, 8.3, 12, 8.6, 11, 11.3, 10.8, 10, 12.1, 8.4, 9.8, 10.7, 10.8, 11.3, 
    10.2, 10.1, 9.5, 8.3, 10.6, 10.4, 9.5, 11.3, 10.1, 10, 12.9, 11.8, 11, 
    10.2, 7.7, 9.6, 10.6, 11.1, 9.7, 9, 9.8, 9.2, 9.2, 9.7, 9, 9.6, 8.5, 7.6, 
    6, 5.6, 5.2, 3.5, 0.5, 0.5, 3.4, 4, 5.3, 6, 7.4, 8.6, 8.6, 11.1, 9.9, 11, 
    10.5, 11.2, 10.2, 10.7, 11.6, 11.2, 9.8, 10.4, 9.9, 8.8, 6.3, 5.8, 4.8, 
    7.2, 4.2, 4.9, 5.8, 8.2, 7.5, 5.9, 4.4, 4.4, 5.1, 3.1, 5.1, 2.9, 1.1, 
    0.4, 1.9, 2.8, 2.5, 2.9, 3.9, 3.6, 3.7, 3.4, 4.5, 4.6, 5.7, 4.8, 7.7, 
    7.2, 7, 5.2, 6, 5.5, 7.2, 7.2, 7.5, 7.2, 5.8, 6.7, 6.4, 7.4, 7.5, 9.5, 
    8.7, 9.8, 10.5, 10, 9, 9.1, 10.7, 10, 12, 12.8, 13.3, 15.2, 16.5, 17.7, 
    17.8, 17.9, 18.1, 18.3, 18.1, 18, 13.9, 4, 6.8, 7.7, 7.9, 9.7, 4.2, 3.9, 
    2.2, 7.5, 6.6, 5.4, 4.8, 5.1, 5.3, 5.8, 5.5, 5, 5.4, 6, 6.4, 6.1, 6.1, 
    6.3, 6.7, 7.1, 7.9, 8.3, 9, 9.3, 8.9, 9, 9.6, 10.2, 10.5, 20.2, 22.7, 
    23.3, 20.5, 23.4, 22.2, 25.9, 26, 12, 24.6, 26.6, 26.5, 25.3, 27.9, 13.2, 
    13.2, 27.4, 26.4, 27.2, 26.1, 25.9, 24.5, 24.2, 24, 11.6, 21.4, 18.8, 
    17.3, 16.7, 10, 16, 13.5, 15.3, 13, 11.6, 11.6, 11, 12.2, 14.8, 13.6, 
    12.9, 14.5, 14.9, 15.4, 13.8, 17.3, 17.2, 16.9, 16.4, 18.1, 16.7, 17.7, 
    18, 15.9, 15.9, 16.5, 16.6, 18.4, 17.1, 16.9, 16, 15.3, 14.7, 15.1, 14.9, 
    14.3, 14.8, 14.7, 13.6, 12.7, 13.5, 13.7, 13.6, 14.3, 14, 13.9, 14.6, 
    15.4, 14.7, 14.6, 15.9, 14.9, 14.7, 14.2, 14, 13.3, 15.2, 14.2, 15, 13.8, 
    13.2, 11.5, 11.4, 11.5, 11.5, 12.2, _, 12.7, 13.3, 13.4, 12.4, 12.4, 
    11.7, 10.7, 12.9, 11.1, 10.2, 10, 9.3, 8.9, 9.7, 7.8, 7.5, 8.4, 8.5, 7.7, 
    7.5, 5.8, 2.5, 0.7, 0.5, 5.5, 4.3, 4.3, 4.9, 6.1, 6.9, 7, 7, 8, 7.8, 8.8, 
    8.8, 8.9, 9, 9.5, 7.8, 8.7, 11.2, 9.8, 10.7, 9.6, 9.2, 11.1, 12.2, 13, 
    12, 12.6, 11.9, 11.3, 11.6, 12.2, 14.2, 12.3, 12.7, 14.1, 14.3, 16.4, 
    14.2, 14.7, 16.6, 16.3, 16.2, 13.7, 13.7, 13.8, 12.5, 10.9, 11.6, 14.2, 
    12.3, 11.5, 10.6, 10.1, 10.8, 10.2, 10.5, 11.4, 9.6, 10.6, 11.4, 11.1, 
    11.1, 12.3, 11.8, 7, 9.3, 7.9, 8.3, 11.8, 10.1, 7.9, 6.8, 12.3, 12.2, 
    15.2, 14.1, 12.4, 13.1, 13.2, 14.1, 12.9, 12.5, 11.5, 9.7, 9.7, 8.8, 8.6, 
    7.5, 5, 2, 0.1, 1, 5.7, 7.8, 6.2, 6.6, 6.3, 6.1, 5.8, 5.1, 5.3, 4.5, 5.4, 
    4.4, 5, 5, 4.9, 3.6, 4.4, 3.7, 3.7, 4.4, 4.8, 4.6, 5, 3.6, 4.8, 7.6, 7.4, 
    5.1, 7.5, 8.6, 8.7, 7.3, 7.7, 9.2, 10.8, 11.2, 9.7, 8.5, 9, 9.6, 12.1, 
    13.1, 13.7, 11.6, 12.1, 11.7, 11.3, 10.5, 11.5, 12.9, 11.8, 11.1, 7.5, 
    8.5, 3.5, 5.1, 2.2, 0.6, 2.5, 2.5, 5.1, 2.6, 3.8, 3.9, 4.6, 4.4, 5.3, 
    6.6, 6.2, 6.9, 7.5, 6.3, 6.3, 6.8, 7.1, 5.8, 6.1, 7.1, 8.2, 7.5, 7.5, 
    7.9, 6.2, 6.2, 6.7, 7.6, 7.3, 7.5, 6.7, 6.4, 7.1, 6.4, 7.5, 6.5, 6.7, 
    6.3, 3.9, 4.1, 4, 2.9, 1.5, 1.9, 2.7, 1.6, 1, 0.9, 0.9, 0, 0.3, 0.9, 2.1, 
    2.1, 3.6, 3.4, 3.5, 4.2, 5.1, 6.2, 6.9, 7, 7.7, 7.9, 7.8, 8.8, 10, 11.3, 
    12.1, 12.7, 12.9, 14, 13.6, 14.5, 15.5, 15.3, 15.6, 15.1, 15.3, 15.8, 
    15.9, 15.7, 15.8, 14.4, 12.4, 11.3, 9.9, 9.4, 8.3, 6.9, 6.6, 6.6, 7.2, 
    6.9, 6, 6.7, 7.1, 6.6, 6.3, 7.4, 7, 6.6, 7.8, 6.1, 7.1, 7.4, 8.9, 10.1, 
    10.2, 10.5, 9.9, 9.3, 8.5, 13.5, 14.3, 14.9, 14.4, 14.4, 14.8, 14.7, 
    15.4, 15.3, 16.1, 16.5, 16.1, 15.5, 16.2, 16.1, 15.8, 16.5, 16.1, 14.6, 
    13.4, 9.7, 7.4, 9.6, 9, 10.9, 9.8, 8.9, 5.5, 3.3, 2.1, 2.3, 5.2, 3.2, 
    5.9, 4, 3.5, 1.2, 2, 6.2, 11.5, 11.2, 11.4, 12.1, 11.8, 12.2, 12, 11, 
    8.8, 7.8, 7.5, 7.1, 5.4, 4.5, 4.2, 3.4, 3.2, 3.8, 3.6, 5, 6.9, 10.4, 
    11.7, 13.4, 13, 12.1, 12.5, 13.5, 11.4, 10.8, 10.7, 11.3, 13.5, 13.1, 
    12.5, 11, 8.9, 7, 6.4, 8.8, 6.9, 4.4, 4, 3.3, 2, 1.7, 0.2, 4.6, 6.4, 6.7, 
    7, 5.5, 7, 6, 3.8, 2.3, 3.1, 2.3, 3.7, 1.9, 1, 5.5, 7.9, 7.1, 6.7, 3.9, 
    2.8, 1.5, 2.6, 5.1, 3, 4.6, 5, 2.9, 4.9, 4.2, 4.4, 5, 3.6, 5, 5.5, 6.7, 
    4.9, 3.3, 4.3, 3.6, 5.9, 5.8, 5.4, 4.8, 4.4, 4.5, 3.8, 2.9, 3.4, 3.4, 
    4.7, 5.3, 5.6, 5.5, 2.1, 0.6, 0.9, 1.2, 11.9, 11.3, 8.8, 10.9, 14.8, 
    16.7, 20.1, 20.4, 24.2, 25, 23.7, 23.2, 23.1, 21.7, 21.8, 18.3, 19.6, 
    10.4, 6.1, 2.6, 4, 3.1, 7, 13.4, 6.5, 11, 11.8, 14.6, 14.2, 14.6, 13.6, 
    15.8, 14.7, 13.6, 14.8, 13.4, 13.1, 15.7, 13.3, 11.9, 12.6, 18, 21.1, 14, 
    11, 12.3, 12.2, 14.3, 14.4, 14.4, 14.8, 15.1, 13.5, 14.3, 14.2, 12.5, 
    12.1, 11.9, 14, 12.8, 14.8, 10.7, 13.8, 14.5, 13.4, 13.1, 12.9, 11, 11.5, 
    10.4, 10.1, 12.7, 12.1, 7.8, 11.4, 10, 9.4, 9.4, 8.3, 12.5, 10.4, 8.3, 6, 
    8.7, 7.8, 9.2, 7.6, 9.9, 8.3, 7.7, 8.5, 13.6, 11.6, 12, 11, 9.5, 13.4, 
    10.6, 11.5, 11.2, 9.2, 9.5, 9, 8.6, 10.6, 9.6, 9.2, 8.4, 9.2, 8.4, 8.6, 
    6.4, 6.5, 6.3, 4.9, 4.1, 5.8, 5.1, 6.8, 6, 6.5, 6.1, 5.8, 4.7, 4.6, 5.1, 
    5.7, 4.1, 2.9, 5, 5.7, 4.3, 2.6, 3.8, 8.1, 6.8, 7.2, 5.8, 4.2, 5.4, 5.1, 
    5.2, 5.6, 6.4, 3.9, 2.8, 3.7, 0.4, 2.8, 2.3, 1.1, 1.6, 1.2, 1.7, 0, 3.9, 
    0.2, 0.7, 4.7, 3.4, 2.8, 4.5, 3.2, 4.1, 4.9, 1.8, 6.4, 7.3, 2.7, 1.6, 
    4.3, 4.7, 2, 2.2, 4.4, 4.8, 4.7, 4.7, 2.6, 1.8, 1.6, 1.6, 7.3, 6.7, 5, 
    4.6, 0.4, 1.4, 0.5, 0.9, 1.7, 1, 2, 3.4, 4.6, 4.3, 4.3, 4.6, 5.8, 6.1, 
    6.9, 6.5, 6.8, 6.5, 7.4, 6.2, 5.4, 6.3, 4.5, 4.3, 3.9, 3.6, 3, 4.7, 3.8, 
    3.2, 3.3, 5, 4.9, 4, 1.6, 0.8, 0.6, 2.4, 3.5, 5.8, 6.2, 6.8, 7.5, 9.8, 
    8.2, 9.3, 8.7, 8.5, 8.3, 7, 7.5, 7.7, 7.3, 6.9, 6.2, 4.8, 8.9, 8.2, 9.7, 
    9.4, 7.9, 7.2, 6.8, 3.5, 3.7, 6.1, 11.5, 13.6, 12.5, 14.4, 13, 11.7, 10, 
    10.8, 10.8, 10.4, 11.6, 10.5, 12.2, 12.5, 13.2, 12.5, 13.1, 12.5, 11.5, 
    11.2, 11.5, 11.1, 11.4, 12.1, 11.7, 11.9, 10.6, 9.6, 10.2, 10.7, 10.4, 
    10.6, 9.2, 9.5, 10.4, 10.7, 11.8, 12.1, 12.9, 14.1, 13.7, 10.7, 6.9, 7, 
    10.1, 10.7, 11.4, 8.7, 0.8, 5.3, 3.7, 3, 3.2, 6.1, 6.8, 7.1, 3.5, 4.4, 
    2.9, 1.5, 0.2, 1.1, 1.8, 2.9, 1.1, 3.5, 5, 4.8, 4.1, 5.2, 8, 8.1, 8.6, 
    8.9, 9.5, 9.8, 9.5, 9.9, 7.2, 13.7, 15.6, 12.3, 2.5, 1.3, 3.4, 3.8, 2.7, 
    3.5, 4.2, 2.8, 1.7, 2.6, 0.7, 3.6, 1.7, 3, 3, 4.1, 2.2, 2.9, 3.3, 5.6, 
    3.5, 4.4, 4.6, 4.2, 5.2, 5.6, 7.8, 8.8, 9.5, 8.6, 3.3, 3.8, 4, 6.2, 3.6, 
    3.1, 3.1, 6.9, 6.8, 7, 6.6, 6.9, 4.8, 5.8, 5.9, 6, 5.8, 5, 4.8, 5.4, 6, 
    5.2, 6.5, 5.4, 6.7, 5.5, 5.6, 5.3, 3.6, 3.7, 3.8, 4.8, 5.4, 4.9, 6.4, 
    7.9, 7.7, 5.2, 7.2, 8.2, 8.1, 8.5, 7.7, 7.6, 9.6, 6.5, 6.6, 8.2, 7.3, 
    6.5, 5.6, 5.1, 4.6, 4, 3.4, 3.7, 3.6, 2.8, 1.7, 2, 0.7, 0.3, 2.3, 1.2, 
    1.3, 2.9, 3.3, 4.2, 4.7, 4.2, 5, 5.4, 5.3, 5.9, 5.7, 6.5, 6.2, 6.1, 6, 
    6.3, 6.3, 6.8, 7.6, 7.6, 6.8, 6.7, 7.5, 7.3, 7.6, 6, 5.3, 5.5, 5.2, 5.4, 
    5.3, 4.8, 4.4, 4.5, 4.7, 4.9, 4.9, 5, 4.8, 4, 4.4, 4.6, 7.9, 7.7, 7.7, 
    8.4, 8.7, 8.7, 8.4, 8.8, 9, 7.5, 6.6, 3.7, 1.5, 0.8, 1.1, 2.4, 7.4, 8, 
    9.2, 10.3, 11.1, 11.3, 10.3, 9.9, 10.3, 7.8, 8.7, 7.1, 7.8, 7.1, 6.9, 
    6.8, 7.4, 6.7, 4.6, 3.7, 5, 2.3, 2.1, 2.6, 4, 4.8, 3.1, 1.2, 1.3, 1.8, 
    1.8, 1.1, 3.5, 3.3, 4.3, 5.8, 5.5, 6.5, 8.5, 9.5, 11.4, 13.2, 12.5, 12.3, 
    11.7, 9.9, 8.6, 8.7, 8.5, 7.5, 6.7, 6.7, 6.7, 6.9, 7.4, 8.2, 7.9, 8.3, 
    8.6, 7.5, 8.5, 9, 8.5, 7.6, 6.5, 6.5, 6, 5.9, 6, 5.2, 6.5, 6.8, 6.4, 6.4, 
    6.2, 5.8, 4.9, 5.9, 6, 5.6, 6.3, 6, 4.9, 4.1, 3.7, 6.5, 0.5, 5.1, 1.4, 
    1.9, 0.8, 6.1, 4.8, 1.9, 5, 3.6, 6.5, 8.4, 7.8, 7.5, 9.1, 8.6, 8.4, 9.2, 
    7.8, 4.6, 1.4, 1.8, 1, 1.7, 2.3, 5.8, 11.6, 10.4, 12.9, 11.3, 10.9, 11.7, 
    10.7, 11.5, 9, 7.4, 7.9, 3.6, 1.4, 0.6, 1.9, 0, 0.4, 0.9, 2.1, 7.6, 8.6, 
    11.3, 9.4, 7.7, 6.4, 8, 8.5, 10.3, 9.3, 9.7, 12.3, 12.5, 10.1, 10.4, 
    11.7, 11.2, 11, 10.9, 10.1, 10.1, 9.9, 9.5, 8.9, 9.1, 8.8, 8.2, 9.1, 8.3, 
    7.1, 8, 7.9, 6.6, 5.9, 5.3, 6.2, 5, 5.7, 4.4, 3.7, 5, 5.3, 2.9, 3.4, 3.1, 
    2.6, 1.6, 2.7, 3.4, 3.3, 3, 2.4, 3.6, 2.3, 2.9, 3.4, 4.5, 4.4, 4.6, 5.3, 
    4.7, 4.8, 4.4, 4.9, 4.6, 4.7, 4.1, 4.4, 5.4, 5.8, 5.3, 6.1, 6.1, 5, 3.1, 
    5.7, 4.4, 5.9, 6.5, 6.5, 6.2, 5, 1.9, 5.6, 4.8, 5.4, 3.8, 3.3, 6.4, 6.4, 
    5.2, 4.6, 5.7, 5.5, 4.2, 4.3, 5, 4.8, 3.4, 1.4, 1.4, 4, 3.7, 4.8, 5.7, 
    6.7, 6.1, 5.1, 5.1, 4, 2.6, 4.2, 2.6, 2.5, 2.3, 3.7, 3.4, 2.8, 1.5, 1.8, 
    2.6, 2.4, 0.9, 0.8, 0.5, 0.8, 4.5, 6.2, 5.1, 1.5, 1.5, 6.9, 3.9, 4.7, 5, 
    4.7, 5.7, 6.8, 6.7, 6.4, 6.6, 6.7, 4.7, 6.4, 5.9, 6.4, 6.7, 5.5, 3.8, 
    5.2, 5.1, 5.6, 5.9, 5.9, 5.7, 5.9, 6.9, 6.4, 4.1, 5.6, 2.6, 5.4, 5.5, 
    3.1, 0.9, 2.6, 7, 3, 1.9, 4, 4.2, 8.8, 8.7, 6.7, 10.2, 8.9, 9, 12.3, 10, 
    12.5, 12.6, 15, 12, 9.7, 11, 12.7, 13.2, 12.4, 13.4, 12.9, 12.7, 12.9, 
    9.3, 12.3, 8.7, 12.9, 13.1, 11.1, 10.8, 8.6, 10.7, 8.5, 11.8, 12, 13.3, 
    14.3, 11.8, 8.2, 10.9, 11.3, 10.1, 10.5, 9.9, 9.1, 8.4, 7.3, 5.2, 6.8, 6, 
    4.3, 5.3, 5.4, 4.6, 4, 4.4, 4.6, 5.4, 4.6, 3.9, 3.5, 5.9, 7.2, 4.7, 5.6, 
    5.1, 6.7, 8.6, 8.3, 10.8, 10.6, 10.5, 10.1, 11.4, 11, 10.7, 8.6, 7.3, 6, 
    8.3, 8.9, 8.6, 7.3, 10.3, 7.4, 5.3, 5.7, 7.3, 5.1, 8.7, 9.6, 12.7, 11.2, 
    12.5, 12.3, 12.3, 11.5, 11.2, 10.8, 12, 10.7, 12, 12.2, 11.8, 12.7, 11.2, 
    11.4, 11.5, 10.8, 9.6, 7.8, 7.5, 9, 9.7, 4.9, 8.1, 6.7, 7.8, 6.9, 4.7, 
    3.1, 6, 5.1, 6.9, 9.2, 7.8, 8.4, 7.1, 5.1, 8, 7, 6.5, 8, 8.3, 7.5, 7.7, 
    8.1, 10.6, 7, 8.5, 8.8, 6.8, 7.2, 7.2, 6.6, 5.6, 5.5, 5.2, 6.3, 6.5, 5.8, 
    10.1, 7.8, 7.8, 8.9, 8.2, 8.5, 8.8, 9.9, 10.3, 9.8, 8.5, 6.9, 6.8, 5.5, 
    4.1, 6, 6.2, 6.1, 6, 4.8, 4.2, 6.5, 6.2, 6.8, 5.4, 4.8, 3.6, 6, 6.2, 6.4, 
    4.6, 2.3, 5.1, 4.8, 3.4, 2.7, 3.7, 5.3, 6.2, 4.3, 4.9, 5.5, 5.5, 5.2, 
    4.7, 4.7, 4.3, 4, 3.8, 5, 4.2, 3.3, 1.8, 1.3, 1.2, 2.2, 1.2, 1.2, 0.5, 2, 
    2, 1.7, 2.9, 3.1, 4.3, 5.6, 6.6, 7.8, 8.5, 8.9, 9, 9.5, 9.3, 9.1, 8.3, 
    7.9, 7.8, 7, 7.5, 6.8, 6.9, 6.7, 5.8, 6, 5.4, 5.6, 5.8, 5.2, 5.6, 5.7, 
    6.4, 6.1, 6.2, 6.4, 5.8, 7.9, 8.3, 9.1, 9, 8.4, 7.9, 7.7, 7.8, 8.5, 10, 
    11.5, 10.6, 11.5, 11.6, 12, 11.4, 10.5, 9.3, 8.9, 6.7, 5.4, 7.3, 3.4, 11, 
    7, 4.4, 7.2, 3.7, 7.8, 9, 5.7, 4.9, 7.7, 8.8, 11.7, 15.3, 11.6, 13.4, 
    17.4, 17.2, 15.7, 15.5, 14.1, 18, 15.6, 17.3, 14.7, 14.8, 18, 16, 22.7, 
    20, 19.6, 17.3, 17, 17.2, 17.7, 15.9, 14.8, 11.7, 13.3, 15.2, 15.5, 11.6, 
    12.2, 13.5, 14.8, 14.5, 16.8, 14, 14.2, 16.6, 14.1, 16.8, 14.5, 12, 11.8, 
    11.6, 13.2, 14.4, 15.7, 12.6, 11.5, 9.3, 9.9, 8.8, 11, 12.3, 15.1, 12.4, 
    15.7, 16.9, 15.8, 15.9, 16, 15.4, 13.5, 12.8, 10.4, 8.1, 8.7, 4.9, 6.3, 
    1.1, 8.9, 1, 0.8, 4.1, 7.2, 8.5, 9.8, 6.5, 8.2, 10.2, 9.1, 8.7, 8.8, 8.6, 
    10.2, 9.9, 9.4, 6, 2.6, 2.1, 13.7, 11.2, 9.8, 11.5, 9.6, 8.4, 8.3, 12.8, 
    4.7, 2, 1.1, 2.1, 1.3, 0.7, 0.5, 2.1, 4.2, 6.7, 9.4, 7.8, 10.9, 12.6, 
    10.7, 8.3, 9.3, 11, 7.5, 9.9, 9.9, 8.8, 8.8, 8.6, 7.6, 7, 5.9, 6.9, 7.2, 
    6.6, 4.5, 5.6, 5.6, 5.8, 5.9, 6, 6.2, 5.6, 5.2, 6, 5.5, 4.6, 4.2, 2.8, 
    2.4, 1.8, 1.8, 1.7, 1.5, 1.5, 1.2, 1.2, 0.9, 0.7, 0.7, 7.5, 7.2, 6.4, 
    6.1, 4.5, 4.5, 4.9, 4.8, 4.9, 4.5, 4.9, 5.3, 4.6, 3.2, 3.6, 3.8, 3.9, 
    3.7, 4.5, 4.9, 5.5, 5.8, 5.3, 5.5, 6.3, 7.4, 6.5, 7.6, 7.9, 7.2, 7.5, 
    7.9, 7.1, 8.1, 8.1, 8, 8.7, 9.1, 9.1, 8, 7.8, 7.7, 7, 9, 7.5, 7.7, 8.1, 
    7.9, 8.4, 7.9, 6.5, 6.1, 8.3, 6.7, 7.2, 6.8, 6.7, 5.8, 6.2, 5.6, 4.6, 
    0.5, 2, 1.7, 1.9, 4.4, 1.7, 0.4, 1.6, 1.1, 1, 0.6, 1.5, 0, 0.2, 4.5, 5.5, 
    4.7, 2, 1.3, 1.6, 1.2, 1.7, 1.1, 1.8, 1.8, 1.5, 1.9, 2.3, 2, 2.2, 2.7, 
    4.1, 2.8, 3.3, 4, 2.7, 2.5, 2.1, 1.2, 2, 1.9, 1.2, 1.4, 1, 0.6, 1.4, 0.7, 
    0.6, 1.2, 1.4, 1.6, 1.1, 3.1, 1.7, 2.2, 2.6, 2.1, 2.7, 2.5, 2, 2.3, 1.6, 
    2.3, 1.5, 1.1, 1.4, 0.8, 0.4, 0.2, 1, 1.2, 1.9, 1.7, 1.5, 2.1, 1.9, 1, 
    1.2, 0.1, 0.7, 0.9, 1.7, 0.4, 0.7, 1.5, 1.7, 2.2, 1.7, 2.1, 3.1, 4.1, 
    1.9, 2.3, 2.2, 3.5, 1.9, 0.9, 1.9, 2.3, 2.1, 2.8, 2.5, 3.1, 3.1, 3.5, 
    3.8, 3.4, 3.3, 3.5, 3.7, 3.4, 3.5, 3.7, 3.5, 2.7, 1.9, 1.1, 3.7, 4, 1.2, 
    2.8, 0.6, 0.8, 1.1, 1.6, 2.2, 1.3, 1, 1.6, 0.4, 0.7, 1.9, 2.2, 2.7, 1.2, 
    0.4, 0.9, 1.5, 1.5, 1.8, 9.8, 9.5, 9.3, 9, 8.6, 2.7, 0.8, 2.8, 1.7, 0.4, 
    7.2, 2, 1.7, 1.8, 4, 3.7, 3.1, 3.9, 4.3, 4.6, 4.7, 5.8, 1.7, 5.8, 4.6, 
    5.1, 4.7, 5, 5.9, 6.1, 5.5, 4.2, 3.2, 3.8, 4.4, 4.6, 4.4, 4.1, 3.4, 1.9, 
    0.7, 0.5, 0.9, 0.7, 2, 3.2, 3.7, 1.2, 1.2, 0.8, 1.9, 1.1, 0.2, 2.1, 2.2, 
    3, 1.2, 1.5, 2.3, 1.5, 0.5, 1.1, 1.8, 4.6, 5.2, 4.7, 3.8, 3.3, 4.6, 4.8, 
    3.5, 3, 3.3, 4, 3, 4.9, 5.2, 7, 6.4, 6.8, 6.4, 6.5, 4.8, 4.5, 5.2, 6.1, 
    3.8, 5.3, 3.9, 8.3, 8.8, 7, 6.7, 7.6, 7.4, 6.8, 7.1, 8.5, 9.3, 7.7, 7.1, 
    8.8, 8.5, 8.8, 9.8, 9.7, 9.2, 9.8, 8.9, 10.1, 7.5, 7.2, 7.3, 8.2, 7.7, 
    6.8, 3.7, 4.7, 4, 3.7, 4, 5.1, 5.3, 4.2, 4.6, 2.6, 1.8, 1.6, 2.1, 2.2, 
    1.2, 1.4, 1.8, 1.9, 3.4, 3.9, 3, 0.9, 1.6, 0.5, 0.8, 1.6, 0.6, 1.7, 1.7, 
    0.2, 1.6, 2.2, 2.7, 1.9, 1.6, 1.6, 2.8, 2.1, 2.3, 0.5, 0.8, 1.7, 0.3, 
    0.4, 0.8, 1, 2.1, 3.9, 3.9, 5.1, 3.2, 3.2, 2.4, 1.7, 1.6, 0.7, 1.7, 3.1, 
    3.9, 4.5, 5.3, 5.6, 6, 6.3, 7, 6.3, 5.7, 6.1, 5.3, 5.8, 5.5, 4.7, 4.5, 5, 
    5.1, 5.1, 5.6, 6.3, 6.4, 7.3, 7.2, 7.8, 7.2, 8.3, 6.8, 7, 8.5, 7.7, 7, 
    7.4, 6.6, 7, 6.7, 5.5, 5.8, 4.9, 5.8, 5.4, 4.8, 4.9, 4.3, 4.5, 3.5, 4.4, 
    3.5, 3.7, 5.2, 5.2, 5.3, 5.4, 5.2, 7.7, 9.3, 8.2, 7.6, 6.1, 6.1, 6.6, 
    6.4, 3.3, 6.7, 5.3, 8.4, 7.8, 7.7, 6, 7.1, 6.6, 6.2, 6.5, 4.5, 6.3, 6, 
    5.5, 6.1, 6.4, 6.2, 7.2, 4.8, 4.2, 4.8, 6.5, 6.2, 7.9, 7.1, 8.6, 10.7, 
    9.9, 12, 9.6, 8.1, 7.1, 6.7, 9.5, 6.4, 5.4, 5.3, 8.2, 8.5, 8.8, 9.8, 
    10.1, 10.8, 7.1, 10.4, 10.1, 10.5, 10.8, 7.6, 3.6, 4.4, 6.7, 3.4, 8.1, 
    6.2, 2, 3.2, 3.2, 4, 2.8, 6.1, 0.8, 2.8, 5.7, 2.5, 3.7, 4.9, 0.5, 5.4, 
    6.7, 7.1, 6.7, 7.9, 6.5, 8.3, 8.1, 9.4, 7.7, 8.7, 9, 6.7, 6.4, 8.1, 6.1, 
    9.4, 8.5, 9.3, 9.9, 11.8, 6.7, 10.9, 7.2, 10.7, 7.1, 7.1, 8, 7.8, 6.7, 
    9.7, 7.2, 8.1, 7.1, 8.6, 9.8, 9.4, 6.4, 7.1, 10.2, 9.3, 6.4, 8.4, 8.4, 
    10.1, 5.6, 8.3, 7.9, 4.9, 8, 7.9, 9, 9.3, 8, 7, 9, 7.5, 9.7, 8.9, 4.3, 
    4.4, 4.9, 5, 7.5, 7.7, 5, 7.3, 8.5, 5.2, 9.2, 7.8, 9.3, 7.1, 6.4, 7.1, 
    8.3, 7.6, 6.9, 7.4, 4.9, 4.5, 9.5, 3.8, 6.5, 8.7, 7.1, 8.6, 5.5, 7.7, 
    9.1, 4.4, 7.9, 7.3, 5.4, 5.3, 6.8, 5.3, 7.6, 5.5, 5.2, 7, 8, 6.1, 5.3, 
    4.2, 5.5, 8.7, 9.7, 8, 8.1, 6.5, 8, 7, 5.5, 7.2, 4.7, 4.5, 5.3, 5.7, 5.1, 
    5.2, 6.2, 4.5, 3.2, 3, 4.8, 5.1, 4.9, 4.7, 4.8, 4.3, 3.7, 3.9, 4.6, 4.8, 
    4.8, 7.4, 7.1, 6.7, 7, 6.2, 9.3, 8.8, 7, 8.1, 8.9, 6.5, 5.7, 7.1, 9.8, 
    10.4, 9.4, 9, 10, 9.9, 10, 8.3, 7.7, 7.7, 6.9, 9, 10.5, 10.3, 7.8, 7.3, 
    8.9, 8.5, 9, 9.1, 9, 10.1, 7.4, 7.7, 8.1, 8.5, 7.7, 8.2, 6.8, 7, 5.2, 
    7.6, 7.9, 7.4, 8.6, 10.6, 9.8, 7.5, 10.5, 6.7, 7.4, 8.6, 6.3, 3.8, 4.5, 
    3.5, 8, 8.5, 8, 5.7, 8, 9.9, 8, 5.1, 5.7, 5, 4.5, 6.8, 12.6, 10.6, 10.4, 
    10.6, 10.3, 12.1, 10.9, 13.5, 11.5, 9.7, 9.5, 13.2, 12.9, 2.4, 6.9, 9.8, 
    10.4, 8.4, 8.2, 8.6, 7.2, 5.1, 5.5, 7.5, 7.4, 4.7, 8.2, 8.7, 7.7, 7.1, 
    8.4, 7.6, 4.7, 6, 5.4, 2.7, 1.3, 3, 2.4, 2.9, 1.7, 0.1, 6.3, 6, 2.4, 3.6, 
    3, 1.5, 6.3, 6.7, 6.8, 4.1, 2.1, 1.9, 1.6, 0.7, 2.8, 5, 3.6, 3, 3.7, 3.4, 
    6.2, 5.5, 6.9, 1, 4.2, 11.4, 11.8, 4, 4.8, 4.6, 2.7, 4.5, 6.9, 3.1, 4.4, 
    6.8, 5.3, 5.9, 4.3, 5.4, 5.9, 3.6, 2.1, 2.3, 0.7, 7, 7.1, 7.6, 7.2, 7.3, 
    7.5, 8.5, 5.9, 4.7, 4.1, 4.7, 3.8, 3.3, 3.9, 4.3, 6.1, 6.3, 5.8, 8, 7.7, 
    4.3, 6.1, 5.2, 4.3, 4.9, 5.2, 5.9, 6.6, 6.7, 7.7, 8.3, 7.5, 4.8, 10.3, 
    10.3, 12.5, 6.4, 6.2, 7.2, 8.7, 10.5, 12.8, 10.9, 14.5, 14.8, 13.5, 15.2, 
    15.5, 13.8, 16.1, 15.5, 15.8, 15.7, 14.2, 13.4, 13.5, 9.3, 10.1, 8.1, 
    7.1, 7.7, 7.6, 5.3, 4, 4.5, 2, 3.1, 3.1, 4.7, 4, 4.4, 6.2, 4.3, 9.1, 7.2, 
    7.3, 10, 7.8, 8.2, 11, 10.6, 8.4, 10.5, 11.5, 10.9, 6.9, 6.8, 12.4, 10.7, 
    11.5, 9.6, 8.1, 8.6, 9.1, 9.4, 4.6, 8.4, 8.4, 9.5, 8.7, 8.2, 6.5, 7.2, 
    7.6, 6.8, 8.1, 8.2, 8.6, 8.6, 8.3, 8.2, 7.1, 7.8, 8.9, 9, 8.5, 8.8, 8.9, 
    8.8, 9.2, 9.1, 9.4, 7.3, 7.8, 6.9, 7.6, 7.8, 4.6, 7.7, 8, 6.7, 6.4, 5.9, 
    5.7, 4.5, 5.1, 5.5, 5, 6.4, 4, 3.7, 5.9, 5.9, 4.2, 6.9, 6.5, 6.6, 5.9, 
    5.7, 5.5, 5.6, 5.4, 5.4, 5.9, 6.4, 3.7, 8, 7.9, 3.5, 4, 4.2, 6.5, 7.9, 
    8.1, 7.1, 4.9, 4.4, 5.7, 5.9, 4.8, 5.8, 5.5, 6, 6.2, 6, 4.2, 3.4, 2.8, 
    2.4, 3.6, 4.7, 4.7, 4.6, 5.6, 5.6, 5.6, 5.9, 5.1, 6.1, 5.7, 7.2, 6.4, 
    9.7, 14.1, 14.7, 13.9, 8.4, 13.7, 14.9, 14.7, 13.5, 13.7, 14.9, 14.6, 
    13.9, 13.7, 13.5, 12.1, 14.8, 7.6, 14.1, 13.1, 13.3, 11.7, 13.9, 12.9, 
    12.4, 14.4, 14.2, 13.8, 13.8, 12.7, 12.4, 13, 12.5, 12.4, 11.8, 9.7, 
    10.9, 11.2, 11.3, 10.5, 11.4, 12.2, 8.8, 10.9, 12.6, 5.6, 10.4, 5.1, 4.4, 
    10.8, 4.3, 13.1, 12.8, 6, 14, 5.1, 15.1, 13.2, 4.6, 9.6, 5.5, 9, 2.5, 
    2.5, 5.5, 5.6, 5.4, 5.5, 5, 4.8, 7.1, 9.9, 12.6, 4.9, 5.9, 9.1, 5.9, 6, 
    11.5, 12.1, 2.5, 5.5, 5.4, 0.4, 3.6, 1, 0.1, 1.8, 2, 0.7, 0.9, 0.7, 1.9, 
    1, 1.6, 0.7, 4.1, 4.8, 1.8, 5.2, 1.2, 0.8, 1, 5.3, 1.9, 0.9, 6, 5.8, 5.6, 
    0.8, 5.1, 5.1, 5.2, 5.2, 5.2, 5.6, 2.3, 2.5, 2.8, 3.2, 2.4, 2, 2.2, 5.5, 
    4.5, 2.4, 4.1, 1.5, 1.7, 6, 1.9, 1.9, 2.7, 5.6, 1.9, 3.8, 1.4, 0.9, 3.2, 
    6, 1.9, 4.5, 5.7, 5.7, 5.7, 6.5, 5.4, 6, 11.1, 10.5, 6.9, 7.5, 8.3, 9.4, 
    5.4, 8.6, 6, 6.1, 9, 8.6, 7.8, 5.2, 8.6, 7.5, 6, 4.3, 4.1, 5.1, 4.4, 5.1, 
    3.7, 4.6, 3.4, 3.6, 3.8, 3.8, 4, 2.9, 2.6, 2.4, 4.2, 3.2, 5.9, 5.4, 7, 
    6.8, 6.2, 7.2, 7.6, 8.1, 8.5, 7.7, 8.6, 7.5, 8.8, 8.8, 8, 8.1, 8.6, 8, 6, 
    8.5, 7.7, 8.1, 8.8, 9, 9.2, 9.6, 8.4, 8.3, 6.8, 7.2, 6.6, 6.5, 7, 6.7, 
    6.5, 4.8, 4.4, 3.5, 3.9, 3, 1.9, 1.5, 2.9, 2.5, 1.2, 0.4, 2.4, 2.4, 2.8, 
    3.7, 3.8, 1.3, 2.5, 2.2, 1.8, 2.9, 2.6, 2.1, 2.9, 3.4, 5.2, 0.6, 1, 0.4, 
    0.7, 0.3, 0.8, 0.7, 0.9, 1.1, 0.1, 1, 0.9, 1.9, 0.9, 0.8, 0.6, 0.8, 1.5, 
    1.7, 2, 1.8, 4.9, 7.1, 7.6, 7.8, 9.5, 9, 7.5, 8, 7.1, 7.8, 7.3, 7.4, 5.9, 
    5.8, 7.1, 6.8, 7, 7.5, 6.6, 8.2, 7.6, 7.8, 7.2, 6.7, 6.5, 6.6, 7.9, 6, 
    4.9, 6.2, 5.8, 4.6, 3.3, 2.7, 4.1, 3.9, 4, 4.3, 5.2, 6, 5.6, 5, 5.5, 5.9, 
    6, 5.7, 5.5, 4.5, 4.3, 3.2, 2.8, 2.9, 3.3, 3.6, 4.3, 4.6, 4.8, 4, 4.2, 4, 
    4.1, 3.7, 3.5, 3.5, 4.6, 5.3, 5.3, 6.5, 5.9, 4.7, 5.3, 4.7, 3.5, 4.4, 
    5.2, 6.2, 5.8, 6.1, 6.2, 6.8, 6.7, 7.5, 7.7, 7.9, 7.9, 8.3, 8.3, 8.4, 
    8.2, 7.7, 6.9, 6, 7.5, 5.4, 1.9, 0.3, 1.2, 0.1, 1.1, 0.1, 0.2, 0.1, 0.8, 
    0.2, 0.2, 1, 2.4, 2.4, 2.3, 2.5, 2.8, 3, 2.9, 3.1, 3.7, 3.4, 3.1, 4, 4.8, 
    4.2, 4.2, 4.4, 3.5, 4, 4.4, 3.6, 2.7, 2.3, 1.9, 1.6, 2.5, 2.9, 5, 7, 5.8, 
    9, 7.2, 7.5, 7.7, 6.3, 5.5, 5.2, 6.7, 6.6, 7.6, 8, 7.4, 5.1, 4.6, 3.4, 
    3.5, 1.6, 2.7, 2.4, 3.4, 2.4, 2.4, 3.6, 3.8, 4, 4.8, 5.5, 6, 5.3, 4.9, 
    5.1, 4.9, 3.4, 3.5, 3, 3, 3.1, 2.4, 2.4, 3.2, 3.2, 3.4, 3.6, 3, 2.7, 3.9, 
    3.3, 2.7, 2.6, 3.1, 2.9, 2.5, 2.1, 2.1, 1.8, 1.9, 0.4, 1.1, 1.7, 3.1, 
    3.1, 4.2, 4.6, 5.6, 6.2, 7.7, 6, 6.2, 6.2, 5.3, 5.8, 6.1, 7.2, 8.9, 8.4, 
    8.5, 8.9, 9.6, 10, 9.4, 7.4, 7.6, 6.1, 7, 6.2, 4.9, 2, 1.3, 0.2, 0.3, 
    1.4, 3.8, 3.9, 4.1, 5.4, 5.4, 4.3, 4.5, 5.8, 7.1, 7.7, 5, 5.1, 1.4, 2, 3, 
    3.9, 3.9, 3.9, 4.3, 4.4, 2.2, 3.2, 4.3, 2.8, 4, 4.3, 7.4, 4.6, 9.2, 5.7, 
    5.3, 6.7, 7.3, 7.6, 6.4, 5.8, 4.3, 2.9, 2.1, 2.1, 1, 1.3, 2.5, 2.7, 3.2, 
    4.1, 4.2, 4.8, 3.7, 3.5, 2.2, 2.8, 2.5, 2, 5.7, 5, 2.1, 3.6, 2.8, 2.7, 5, 
    4.2, 5.6, 5.9, 8.8, 8.9, 9, 9.6, 10.7, 9.2, 9.1, 9, 8.4, 8.5, 8.8, 9.4, 
    8.2, 10.5, 9.2, 9.5, 9.7, 9.9, 9.1, 10.7, 11.5, 10, 10, 9.1, 9.8, 10.2, 
    10.1, 9.3, 9.1, 8.9, 7.9, 7.7, 6.6, 6.9, 7.3, 6.2, 7.4, 8, 7.2, 6.2, 6, 
    5.9, 7.9, 7.1, 6.4, 6.8, 5.6, 3.9, 3.2, 2.4, 1.1, 0.2, 1.4, 0.8, 0.5, 
    1.5, 1.5, 5.4, 7.3, 7.3, 7.1, 8.4, 8.4, 7.8, 7.5, 7.3, 7.5, 8.2, 8.5, 
    8.4, 8.2, 8.5, 7.5, 6.1, 6, 4.5, 3.9, 5.8, 4.5, 2.4, 1.3, 0.7, 1.2, 0.9, 
    0.4, 0.2, 0.5, 0.6, 0.9, 0.6, 2.5, 2.8, 1.2, 3, 1.1, 0.9, 1, 2.5, 4.2, 
    2.5, 0.8, 1.4, 7.1, 6.3, 6.1, 7.4, 7.4, 7.2, 5.9, 6.1, 7, 7.8, 6, 7.6, 
    8.9, 10.3, 11.6, 11.5, 11.2, 12.2, 11.7, 10.9, 12.1, 11, 10.1, 10.6, 
    11.6, 13.1, 12.8, 13.2, 13.4, 12.6, 10.3, 10.4, 11.9, 12.2, 11.2, 11.3, 
    10.8, 12.8, 13.8, 10.6, 12.5, 13, 9.9, 10.3, 10, 9.7, 9.3, 9.8, 8.1, 7.7, 
    8, 8, 7.2, 6.9, 5.5, 5.5, 5.9, 6.9, 7.4, 8, 7.8, 7, 6.1, 5.8, 5.2, 5.3, 
    4.4, 3.7, 3.9, 4.9, 5.7, 5.3, 5.5, 5.4, 7.8, 8.4, 6.6, 6.8, 5.9, 4.9, 
    2.3, 3.8, 4, 4, 4.7, 5.4, 5.9, 6.2, 5.1, 5.1, 4.7, 4.4, 4.1, 3.6, 4.6, 
    4.9, 5.5, 4.7, 6.6, 6.6, 7.3, 7.1, 8.1, 6.8, 5.4, 7.4, 6, 7.3, 7.4, 7.5, 
    7.1, 6.6, 5.2, 2.8, 4.5, 6.4, 7.2, 8.3, 8.4, 8.6, 8.7, 7.4, 7.4, 7.2, 
    6.3, 7.5, 5.5, 2.8, 5.7, 6, 5.2, 4.4, 4.5, 3.3, 1.5, 2.9, 2, 4, 3.7, 4, 
    5.1, 3.7, 2.4, 2.7, 7.1, 5, 4.3, 3.3, 4, 4.8, 3.4, 4.3, 3.4, 3.1, 3.2, 
    4.3, 4, 4.6, 3.9, 3, 3.2, 2.8, 5.4, 2.1, 10.2, 10.8, 9.6, 9.7, 12, 12.9, 
    9.3, 10.9, 11.9, 11.6, 12.1, 12, 9.5, 12, 11, 9.8, 10.7, 11.6, 13.1, 
    11.3, 11.2, 13.4, 12.7, 13, 13.1, 13.5, 13.7, 13, 12.1, 12.3, 13, 13, 
    13.9, 14.6, 13, 15.4, 15.6, 14.8, 15.5, 14.2, 13.4, 13, 12.4, 11.8, 12.6, 
    12.4, 11.9, 14.9, 12, 14.3, 14.9, 15.9, 15.2, 14.3, 14.7, 15.8, 13.9, 
    14.9, 14.9, 12.3, 11.6, 12.2, 11, 11.4, 11.3, 12, 13.6, 10.1, 9.7, 9.6, 
    9, 8.2, 10.7, 10.8, 12.8, 13.6, 12.7, 12.4, 10.9, 13, 11.3, 12.8, 12, 
    11.4, 11.1, 11.5, 13.1, 13, 12.5, 13.7, 12.3, 12.2, 11.9, 12.9, 12.5, 
    12.6, 13.1, 10.8, 11.7, 11.8, 12.6, 10.9, 8.8, 7.6, 8.4, 7.4, 7.3, 7.8, 
    7.8, 6.5, 5.4, 5.1, 5.3, 5, 3.5, 3, 2.9, 3.3, 6.1, 5.9, 4.9, 5.4, 3.8, 
    2.5, 1.9, 0.2, 3.1, 5.2, 4.6, 4.5, 4.4, 2.7, 0.4, 1.1, 1.3, 2.7, 3.4, 
    3.6, 4.1, 3.9, 4.2, 5.3, 5.6, 4.9, 5.6, 7.7, 7.8, 7, 6, 8.4, 8.9, 9.6, 
    9.8, 6.9, 6, 6.7, 7.9, 8.5, 8.7, 9.3, 9.7, 9.5, 9.5, 11.4, 13.2, 14.2, 
    15.6, 12.8, 12.1, 15.9, 13.6, 15, 16.1, 16.2, 15.9, 15.1, 13.2, 10.5, 
    5.3, 7.1, 6.9, 6.3, 4.6, 3.1, 1.7, 1.1, 5, 4.4, 5.1, 6.3, 8.6, 8.6, 9.9, 
    9.6, 11.3, 12.8, 14.2, 14.9, 15.8, 14.3, 13.1, 14.8, 13.7, 11.8, 11.3, 
    10.7, 11.7, 11.9, 12.6, 10.9, 11.8, 13, 13.1, 12.3, 11.5, 11.4, 11.4, 
    11.7, 12.8, 11.1, 9.8, 9.2, 7.9, 7.8, 7.1, 7.2, 4.4, 2.6, 2.3, 3.7, 4.7, 
    5.2, 5.3, 6.7, 7.2, 6.6, 5, 6, 4.8, 5.2, 4.9, 7.6, 9.7, 9.8, 10.4, 12.7, 
    11.8, 11.4, 10.4, 8.7, 7.5, 6.1, 5.1, 5.2, 4.2, 1.6, 0.9, 2.9, 4.6, 6.1, 
    5.6, 5.4, 6, 6.4, 6.7, 6.8, 6.1, 6, 6.3, 5.7, 5, 4.7, 4.1, 3.4, 3.5, 3.1, 
    3.4, 1.9, 1.9, 6.6, 8.9, 5, 4.1, 4.1, 2.8, 2.4, 2.8, 3.9, 3.2, 3.1, 3.5, 
    4.8, 4.9, 8.3, 8.7, 8.4, 8.6, 9.6, 10.7, 8.8, 8.2, 5, 3.1, 0, 1.3, 2.4, 
    2.5, 3.3, 3.8, 3.9, 4.7, 3, 0.8, 1, 0.8, 1.4, 0.3, 0.6, 1.2, 1.2, 2.3, 
    4.5, 7.6, 8.8, 9.3, 10.1, 10.4, 10.2, 11.3, 10.9, 10, 10, 9.3, 9.1, 9.6, 
    9.1, 9.9, 9.9, 8, 7.7, 7.9, 7.4, 4.7, 2.6, 1, 6.4, 7.9, 10, 10.5, 11.7, 
    11.3, 11.1, 11.8, 10.9, 10, 9.3, 11.5, 9.5, 8.6, 7.3, 5.7, 5.4, 4.8, 2.2, 
    3.2, 3.4, 1.4, 5, 4.4, 4.3, 4.2, 4, 5.2, 5.3, 5.4, 5.8, 6.5, 7, 6, 5.9, 
    6.7, 7.5, 7.4, 7.6, 8.4, 8.1, 8.6, 9, 8.6, 8.4, 9.2, 8.4, 6, 7.3, 5.7, 
    4.2, 1.8, 1, 2.1, 1.7, 0.6, 2.3, 5.4, 6.5, 8.2, 12.1, 13.3, 10, 3.8, 1.2, 
    1, 1.2, 1, 0.5, 0.6, 2.7, 4.7, 2.7, 3.2, 3.7, 6.6, 8, 7.4, 5.1, 4.9, 4.4, 
    4.1, 4.3, 4.6, 2, 1.2, 0.5, 6.5, 6.2, 4, 7.5, 9, 8.7, 7.3, 8.7, 9.7, 9.3, 
    8.6, 8, 9.4, 8.5, 8.5, 7.5, 7.7, 7.2, 7.8, 7.4, 8.2, 9, 8.4, 8, 8.3, 7.5, 
    7.2, 7.3, 7.3, 7, 5, 5.7, 6.1, 6.3, 5.3, 5.6, 5.1, 4.2, 2.9, 1.4, 0.8, 
    0.6, 0.8, 1.7, 1, 2.2, 1.5, 2.9, 1.9, 1, 1.6, 2, 3.8, 6.7, 5.2, 4.4, 8.7, 
    9.5, 9, 6.9, 7.5, 6.6, 8.5, 7.9, 6.6, 7.5, 6.4, 7.2, 9.2, 7.8, 8.2, 7, 4, 
    2.3, 3.2, 1.6, 4.6, 5.5, 5.9, 6.7, 6.7, 8.7, 9.6, 8.1, 8.7, 10.5, 8.7, 
    8.2, 7.8, 7.6, 6.5, 6.8, 6.9, 7.4, 7.7, 9.4, 7.7, 7.8, 8.9, 7.3, 8.4, 
    6.7, 7.7, 6.6, 5.6, 5.1, 4.1, 3.5, 2.6, 2, 1.2, 3.1, 3.9, 5.3, 7, 7.8, 
    6.2, 4.2, 6.4, 9, 8.4, 3.6, 4.7, 5.2, 6.7, 4.8, 5.6, 5.9, 2.1, 1.2, 3.6, 
    2, 1.5, 1.1, 2, 2.5, 4.8, 5, 6.1, 6, 5.6, 4.3, 2.2, 2.5, 1.1, 4.5, 1.4, 
    0.1, 3.8, 1.9, 1.7, 0.3, 0, 0.9, 0.6, 2.6, 2.8, 4.8, 5.3, 3, 4.1, 5.4, 
    5.6, 5.1, 4.5, 4.4, 4.3, 4.9, 1.3, 1.7, 2.5, 3.7, 4.8, 5.4, 6.1, 4.2, 
    5.5, 5.6, 5.7, 6.1, 5.9, 6.4, 5.5, 4.9, 4.7, 5, 5.1, 5.1, 3.9, 5.1, 5, 
    5.2, 4.4, 5, 6.1, 5.1, 4.9, 5.2, 7.2, 6.4, 6.1, 5.7, 5.8, 6.8, 5.6, 3.3, 
    2.8, 2, 2.3, 1.6, 2.1, 2.4, 3.4, 4.5, 5.1, 6, 6.5, 6.8, 7.5, 7.6, 6.1, 
    4.4, 3.9, 4.1, 5.4, 4.7, 5.6, 7.7, 8.2, 9.8, 9.3, 9.5, 9, 7.4, 8.7, 8.2, 
    8.2, 8.9, 8.5, 8.7, 9.4, 9.2, 11, 11.6, 12.3, 10.4, 9.8, 6.1, 4.1, 5.1, 
    7.2, 10.8, 10.6, 9.8, 8, 8.9, 9.7, 9.8, 12.6, 11.3, 13.6, 14.2, 12.3, 
    13.8, 16.5, 16.5, 15, 13.2, 13.9, 13.8, 13.4, 13.1, 13.2, 13.7, 12.2, 
    10.8, 8, 5.4, 2.8, 1.3, 6.7, 12.6, 15.8, 18.8, 20.1, 21.1, 17.4, 17.7, 
    16, 15.9, 21.2, 15.9, 16.5, 16, 16.4, 17.3, 15.8, 15.7, 18.2, 17.8, 16.2, 
    16.7, 15.2, 15.2, 15.6, 14.4, 15, 12.4, 13.2, 16.4, 14.3, 12.5, 12.1, 
    11.6, 11.1, 10.9, 10.7, 10.6, 10.3, 10, 9.6, 9.1, 8.4, 8.9, 8.3, 7.8, 
    7.4, 6.8, 5.8, 4.9, 4.7, 4.8, 4.6, 4.8, 4.7, 3.9, 4.6, 4.6, 4.5, 4.2, 
    4.3, 4.5, 4.5, 4, 3.3, 3, 3.1, 3.7, 3, 2.8, 2.7, 2.9, 3.1, 3.4, 3.6, 3.4, 
    3.3, 3.2, 3.1, 2.8, 3.1, 3.3, 3.4, 3.1, 2.9, 2.9, 2.9, 3, 3.4, 3.8, 4.2, 
    4.8, 5.2, 6.3, 7.5, 8.1, 8.5, 8.1, 7.6, 7.3, 7.1, 6.9, 6.1, 7.5, 7.3, 
    6.6, 5.9, 5.5, 5, 4.9, 4.7, 4.6, 4.3, 4.1, 4.1, 4.9, 5.1, 4.9, 5.8, 6, 
    6.7, 6.6, 6.3, 5.9, 5.8, 6.2, 5.4, 5.3, 5, 4.3, 4.4, 5.5, 5.4, 4.6, 4.1, 
    5.1, 5.5, 5, 4.5, 5.2, 4.1, 2.6, 0.9, 0.2, 2.6, 6.6, 7.9, 7.7, 7.9, 6.8, 
    7.9, 8.8, 8, 7.6, 7.9, 8.1, 7.7, 7, 7.1, 6.7, 7.1, 6, 6.6, 6.5, 5.3, 5.6, 
    5.5, 5.5, 5.6, 6.1, 6.1, 6.3, 5.7, 6.4, 5.7, 6.1, 6, 5.5, 6, 6.7, 6.3, 
    6.6, 6.8, 7.2, 7.1, 6.9, 8.1, 8.3, 7, 7.7, 6.4, 7.3, 7.4, 6.6, 7, 5.2, 
    4.2, 3.4, 3.1, 4.4, 5.7, 4.1, 5, 5, 6.4, 5.1, 4.6, 5.8, 5.4, 5.2, 4.7, 
    5.2, 6.5, 6.4, 7.4, 6.6, 7.2, 7, 7.2, 8.8, 7.9, 12.1, 7.9, 8.7, 8.8, 9.1, 
    10.3, 7.6, 8.2, 7.6, 7.6, 6.8, 6.2, 6.5, 6.3, 4.9, 5.3, 4.6, 3, 2.1, 3.2, 
    4.7, 5.3, 6.9, 8.4, 4.5, 5.5, 6.4, 5.6, 6.2, 6.9, 9.1, 8.4, 7.2, 6.9, 
    7.1, 7, 7.8, 8, 8.5, 7.8, 6.7, 7.6, 8.1, 8.8, 8.4, 8.5, 9, 10.8, 10.9, 
    9.1, 8.9, 8.4, 8.3, 9.5, 8.9, 7.4, 8.1, 8.6, 8.6, 10.2, 10.5, 10.6, 7.7, 
    8.2, 10.5, 10.7, 7.8, 8.1, 7.3, 6.4, 5.8, 3.6, 6.7, 3.8, 4.7, 5.5, 5.4, 
    5.6, 6.5, 5.2, 5.1, 4.8, 5, 5.6, 5.6, 6.5, 5.1, 6.5, 7.7, 6.2, 6.1, 6.7, 
    6.9, 6.7, 6.1, 6.3, 5.7, 5.9, 6.4, 5.3, 5.2, 5.1, 4.1, 4.8, 6.2, 6.2, 
    5.8, 5.6, 5.9, 5.5, 5.1, 5.7, 5.6, 5.5, 7.1, 7.8, 7.8, 7.2, 8, 7.3, 8.7, 
    10.5, 10.5, 12, 11.2, 11.9, 13.2, 13.5, 13.2, 13.1, 14, 15, 14.5, 13.3, 
    15.5, 11.4, 14, 17.7, 18.1, 17.7, 17.4, 19, 19, 19.5, 20.9, 20.6, 21, 
    21.1, 22.2, 22.7, 25, 25.4, 23.8, 23.9, 22.5, 20.8, 20.1, 18.9, 17.8, 
    16.6, 15.4, 14.4, 14.4, 12, 12.9, 13.5, 14.3, 13.5, 12.8, 13, 12, 12.3, 
    11.5, 11.5, 12, 11.5, 7.1, 9.5, 7.9, 8.5, 8.4, 5.9, 6.2, 5.7, 7.5, 8.4, 
    5.1, 5.7, 5.6, 5.4, 4.9, 5.4, 4.5, 3.4, 1.9, 2.2, 1.7, 2, 2.3, 2.8, 2.9, 
    2, 1.8, 0.1, 1.3, 0.3, 0.9, 1.2, 1.4, 3.7, 3.6, 3.6, 2.4, 3.6, 4.1, 4.2, 
    4.9, 5.1, 6.8, 7.3, 7.1, 6, 6, 6.3, 6.5, 7.2, 7.7, 8.6, 5.1, 5.8, 2.8, 
    2.2, 0.9, 1.3, 1.8, 0.3, 1.7, 4.4, 4.5, 5, 5.7, 7.3, 10.6, 11, 12.1, 
    12.6, 13.2, 13.8, 13.2, 11.5, 12.1, 11.1, 11.9, 10.6, 9.7, 8.6, 10.9, 
    11.7, 10.9, 10.8, 10.7, 8.5, 9.1, 7.8, 6.2, 5.6, 7.9, 7.9, 6.8, 6.5, 5.4, 
    5.7, 3.2, 6.3, 7.9, 8.7, 8.4, 7.5, 7.8, 6.4, 2.7, 5.5, 6.1, 7.5, 7.1, 
    7.8, 7.8, 9.4, 9.6, 8.7, 7.6, 8.5, 8.8, 7.8, 7.3, 7.3, 4.5, 5.5, 7.7, 
    7.3, 6.2, 9.1, 7.3, 5.7, 5.8, 7.2, 10, 11.4, 10.7, 10, 10.2, 7.9, 7, 7.7, 
    7.9, 6.9, 8.3, 8.2, 7.3, 8.3, 8.5, 8.6, 8.4, 8.9, 8.9, 8.3, 6.1, 8.6, 
    7.9, 7.8, 7.4, 7.9, 8.5, 8.8, 8.1, 8.5, 8.7, 9.5, 8.2, 9.7, 9.3, 10.8, 
    10.7, 10.2, 10.5, 9.8, 15.8, 17.1, 19.5, 17.6, 18.4, 20.7, 20.6, 20.2, 
    14.4, 8.5, 9.6, 10.6, 13.5, 12.5, 11, 11.2, 10.4, 8, 5, 6.4, 5.9, 9.4, 
    14.4, 18.4, 17.9, 18.1, 12.7, 11.3, 11.8, 11.1, 10.6, 10.8, 10.1, 11.3, 
    11.6, 10.8, 12.7, 14.5, 13.4, 13.8, 13.9, 14, 13.9, 11.5, 13.4, 12.5, 
    15.6, 17.1, 15.2, 18.8, 18.4, 18.1, 15.8, 13.9, 14, 14.5, 13.1, 12, 11.3, 
    11.1, 12.6, 11.2, 10.8, 8.7, 10.1, 8.9, 8.8, 8.5, 8.5, 8.3, 8.2, 7.8, 
    7.4, 7, 6.4, 5.3, 5, 3.9, 4.9, 6.9, 5.4, 4.5, 2.9, 2.4, 4.1, 1.8, 1.7, 
    2.3, 6.6, 6.8, 8.7, 9.2, 7.7, 10.3, 9.7, 9.6, 10.2, 10.9, 10.1, 11.4, 
    9.7, 11.2, 12.8, 14.3, 14.3, 13.5, 13.1, 13.2, 13.1, 13.8, 14.9, 13.1, 
    13.4, 14.6, 13.9, 14.5, 14.3, 15.2, 15.5, 15.4, 15, 13.8, 13.3, 12.3, 
    10.9, 12, 9.9, 9.6, 8.8, 9, 9.2, 9.2, 8.2, 8.1, 7.7, 6.1, 5.5, 4.8, 5, 
    3.5, 3.9, 3.6, 4.2, 4, 5, 8.8, 10.2, 11, 10, 11.3, 10.1, 9.9, 11.1, 10.8, 
    11.9, 11.2, 11, 13.1, 13.9, 13.6, 10.8, 9.4, 10, 8.2, 7.3, 6.5, 6.6, 6.3, 
    6.4, 11.6, 9.3, 8.6, 8.2, 8.1, 7.9, 7.5, 7.6, 8.3, 8, 7.2, 7.1, 7.1, 6.4, 
    7.8, 8.8, 7.8, 7.4, 8, 9.2, 8.1, 8, 7.6, 8.9, 9.9, 9.1, 8.5, 9.3, 11.6, 
    11.5, 10, 8.1, 7.7, 6.9, 8.3, 8.2, 7.6, 7.5, 7.1, 8.3, 8.2, 4.9, 8.1, 
    7.5, 6.4, 4.7, 5, 6, 4.6, 2, 0.9, 2.4, 1.9, 0.9, 2, 10, 9.4, 8.1, 7.4, 4, 
    1.3, 1.1, 1, 4.7, 2, 3.4, 7.2, 9.5, 12.7, 13.8, 13.7, 13.4, 13.2, 13.8, 
    13.5, 9.5, 9.2, 10.3, 9.7, 8, 7.3, 7.6, 7.3, 6.1, 5.3, 6, 6.3, 7.2, 7.4, 
    6.3, 7.9, 7.6, 7.2, 7.6, 7.6, 7.1, 7.7, 8.5, 8.5, 10, 10.5, 11.3, 10.3, 
    11.7, 13.1, 13.4, 13.2, 13, 13.5, 11.8, 12.6, 12.6, 13.2, 14, 13.5, 13.7, 
    13.9, 12.8, 10.9, 14.9, 10.6, 10.5, 10.5, 9.3, 9.1, 9.7, 8.1, 7.3, 7.9, 
    5.8, 3.7, 2.3, 4.1, 5.3, 10, 12, 14, 13.3, 11.1, 9.4, 9.9, 12.1, 12.5, 
    14, 9.6, 12, 12.2, 12, 9.2, 8.7, 6.1, 10.9, 12, 13.6, 13.5, 13, 12.6, 
    10.3, 8.2, 4.9, 3, 3.2, 0.4, 7.9, 8.7, 10.2, 11.6, 9.6, 7.9, 7.6, 5.9, 
    5.4, 5.6, 5.4, 6, 6.2, 7.4, 6.6, 6.7, 6.9, 6.7, 8.4, 8.7, 8.2, 8.8, 11.3, 
    9.9, 11.4, 11.8, 9.9, 10.2, 8.3, 8.2, 8.5, 8.8, 9.6, 9, 10.2, 11.7, 12, 
    11.9, 12.3, 11.9, 12.7, 13, 14.5, 12.6, 13.3, 13.6, 13.1, 13.5, 13, 12.9, 
    11.1, 7.9, 7.8, 7.5, 8.8, 7.5, 8.4, 8.9, 7.7, 8.7, 10.2, 10.8, 11.5, 
    10.2, 10.9, 8.3, 7.9, 7.4, 4.9, 4.3, 5.8, 6.1, 6.6, 8.4, 7.6, 7.7, 7.7, 
    8.1, 8.3, 8.9, 9.5, 8.3, 9.4, 9.2, 10.5, 10, 10.7, 11.4, 12, 11.4, 12.1, 
    12.3, 13.5, 13.6, 12.8, 12.9, 12.5, 14.1, 13.6, 13.9, 16.4, 14.6, 14.5, 
    14.4, 14.2, 15.3, 15.2, 13.8, 13.4, 13.5, 14.1, 13.2, 12.7, 12.9, 14.3, 
    13.2, 14.2, 14.2, 15.2, 14, 14.1, 13.6, 14.3, 14.3, 14.5, 13.7, 13.5, 
    13.2, 11.9, 13.3, 12.9, 13.1, 12.3, 11.7, 12.3, 13.4, 11.5, 10.6, 10.8, 
    10.1, 9.3, 9.2, 9.7, 10.5, 12.1, 10.8, 10, 9.7, 9.5, 9.8, 9.6, 10.2, 8.8, 
    8.7, 8.7, 8.5, 8.4, 8.7, 8.1, 8.6, 8, 8.2, 8.1, 7.2, 8.2, 8.1, 7.1, 7.5, 
    9.1, 7.8, 8, 8.6, 8.8, 10.5, 11.6, 10.8, 11.6, 10.4, 11, 11.8, 10.4, 8.7, 
    8.7, 11.2, 11.3, 11.1, 9.8, 11.5, 11.6, 11, 10.5, 11, 11, 13.4, 12.8, 
    12.2, 12, 13.4, 14.2, 15.6, 18.2, 17.8, 18.7, 19.1, 19.5, 20, 18.3, 17.5, 
    15.4, 15.4, 14, 13.1, 13.6, 13.1, 13.8, 10.9, 10.9, 9.6, 11.5, 12.9, 
    12.9, 12.3, 9.1, 10.9, 10.4, 9.6, 9.2, 8.3, 7.8, 9.6, 8.4, 11.2, 9.4, 
    12.2, 11.9, 12.5, 12.1, 11.2, 11.4, 11.9, 11.8, 12.7, 12.1, 13.3, 14.5, 
    14.4, 10.7, 11.6, 11.2, 10.5, 9.2, 9.1, 9.3, 9.1, 9.6, 8.1, 7.6, 6.8, 
    3.4, 5.5, 4.7, 3.6, 4.3, 4.9, 4.3, 3.8, 3, 3.2, 2.1, 6.4, 13.2, 10.2, 10, 
    9.4, 10.7, 9.2, 9.7, 9.8, 10.2, 9.6, 10.3, 9.5, 8.4, 8.5, 8.3, 8.5, 7.9, 
    7.3, 5.9, 5.8, 5.9, 4.7, 5.2, 5.3, 4.3, 4.8, 5, 4, 5.8, 4.5, 5.3, 7, 5, 
    9.3, 9.7, 9.9, 11.6, 13.1, 14.8, 16.4, 16.8, 16.9, 17.1, 15.3, 12.6, 
    10.6, 3.3, 6, 2.4, 3.5, 3.5, 3.7, 5.2, 3.9, 5.2, 5.4, 15.8, 16.4, 17.8, 
    17.8, 18.1, 17.9, 16.7, 18, 16.2, 14.5, 13, 13.4, 12.8, 13.4, 12.5, 12.6, 
    11.6, 10.4, 10.5, 10.5, 9.9, 10.2, 9.6, 8.3, 7.6, 7.8, 7.4, 7.1, 8, 6.6, 
    3.5, 4.7, 3.9, 2.6, 1.4, 3.2, 2.9, 3.4, 4.2, 4.7, 9.4, 13.2, 11.6, 11.1, 
    8.9, 4.5, 6.7, 5.9, 7.7, 7.5, 7.2, 7.9, 9.5, 9.3, 11.9, 12.7, 9.7, 12, 
    13.3, 12.3, 11.6, 10.4, 11.6, 8.3, 7.2, 7.3, 7.3, 6.7, 5.9, 5.5, 5.4, 
    3.2, 10, 9.2, 9.4, 10.8, 11.9, 7.8, 8.7, 7.5, 5.5, 5.7, 6.5, 6.1, 7.5, 
    6.1, 7.3, 5, 13, 14.5, 15, 16.8, 14.2, 14.1, 13.9, 16.2, 17, 13.5, 11, 
    8.4, 5.6, 8.2, 3.4, 4.4, 4.7, 6.9, 6.8, 7.7, 6.6, 5.9, 3, 4.1, 2.2, 0.7, 
    7.8, 6.3, 3.2, 3.6, 6.2, 6, 5.1, 7.8, 8.8, 9, 10.5, 10.2, 7.9, 5.1, 5.8, 
    6.4, 6.6, 6.6, 7.1, 8.1, 8.5, 8.8, 9.6, 9.8, 8.5, 7.9, 9.5, 9, 7.2, 9.1, 
    10.8, 8.8, 9.4, 8.8, 8.1, 8.3, 8.8, 10.8, 11.2, 10, 9.9, 12.1, 12.1, 
    11.3, 11.6, 11.8, 13.5, 13.1, 10.1, 10.6, 12.3, 11.1, 10.6, 10.2, 9.5, 
    9.2, 9, 8.7, 8.9, 8.1, 6.3, 7.4, 6.8, 10.7, 9.3, 7.9, 7.5, 7.8, 7.7, 9.9, 
    10.2, 9.6, 10.2, 9.4, 8.7, 7.5, 7.4, 7.7, 7.4, 8.9, 8.8, 7.8, 8, 8.2, 
    6.1, 8, 9, 11.4, 9.5, 8.5, 9.9, 9, 7.1, 9.8, 10.6, 6.1, 5.9, 9.1, 9.4, 
    9.3, 6.5, 13.7, 15, 16.1, 15.3, 17.8, 19.1, 19.3, 19.9, 20.1, 19.9, 18.7, 
    18.7, 12.7, 19.3, 19.7, 18.2, 16.4, 16.3, 15.6, 14.6, 15.7, 15.2, 14.3, 
    12.9, 11.4, 10.7, 9.9, 9.7, 8.1, 7.6, 7, 8.4, 10.7, 12.9, 7.9, 10.3, 8.8, 
    8, 11.1, 9.5, 12.5, 12.4, 9.8, 10.2, 11.7, 11.8, 11.6, 12.8, 12.9, 13.1, 
    13.5, 12.6, 13, 10, 9.1, 11.2, 10.1, 11.5, 11.8, 11.7, 11.2, 11.3, 9.9, 
    9.9, 11.7, 11.2, 11.4, 10.9, 10.9, 11.8, 11.9, 11.5, 8.6, 12.1, 11.3, 
    10.9, 10.2, 11.4, 11.1, 10.5, 12.1, 12.3, 12, 12, 11.8, 12, 11.1, 13.3, 
    12.9, 12.9, 12.8, 11.8, 11.5, 11.5, 14.3, 14.5, 13.8, 14.5, 15.5, 15, 14, 
    12.2, 10.9, 10.7, 10.5, 13.4, 14.2, 13.8, 15.2, 16.4, 18, 19.6, 18.4, 
    15.9, 15.3, 16.4, 16.9, 16.7, 14.9, 13.4, 12.7, 14.5, 16.6, 16, 17, 18, 
    19.9, 20.7, 24, 24, 20.3, 17.9, 18.5, 18.2, 17.3, 15.4, 14.6, 13.5, 12, 
    11.2, 14.1, 16.2, 16.6, 16.6, 15.8, 18.7, 18.4, 17.4, 19.8, 16.3, 15.8, 
    18.3, 17.6, 17.5, 17.7, 17.4, 12.5, 8.5, 9.3, 8.4, 7.6, 11.2, 14.8, 14.1, 
    15.2, 14.5, 14.5, 14.5, 12.9, 11.8, 12.8, 8.5, 4.4, 1.2, 13.6, 15.3, 
    15.7, 10.7, 10.8, 7.1, 11.2, 12, 13.3, 11.9, 11.8, 11.8, 8.6, 4.6, 4.7, 
    7.7, 7.9, 8.4, 8.7, 9.3, 9.1, 9.2, 9.2, 9.7, 11.5, 11.5, 11.3, 10.5, 9.4, 
    9.2, 8.4, 7.9, 7.6, 6.9, 7, 6.3, 6.9, 5.6, 7.1, 5.9, 6.1, 4.8, 5.5, 4.6, 
    7.2, 6.4, 5.5, 6.8, 5.4, 7.8, 6.5, 5.6, 7.2, 6.6, 6.2, 5.6, 6.1, 6.7, 
    5.4, 3.6, 7.1, 6.7, 5.6, 7.5, 6.2, 6, 5.7, 6.5, 4.9, 5.7, 6.9, 6.8, 6.6, 
    8.2, 6.1, 7.3, 6.5, 6.6, 7, 5.7, 5.4, 5.4, 5.2, 3.4, 3.2, 3.8, 3.5, 3.6, 
    5.5, 5.5, 8.6, 10, 10.2, 10.6, 11.3, 11.5, 10.2, 9.6, 8.5, 9.7, 10.1, 
    10.5, 9.3, 8.8, 9.3, 8.1, 7.8, 11.3, 11.6, 11.5, 9.3, 3.3, 6.2, 5.5, 6.9, 
    7.6, 9.2, 10, 11.2, 10, 10.9, 10.1, 10.7, 10, 10, 10.1, 9.5, 9.6, 8.6, 
    9.8, 9.3, 9.8, 10.7, 10.5, 10, 9, 9.2, 9.3, 9.9, 10.5, 10.6, 10.4, 10.9, 
    10.3, 10.1, 10.6, 11.2, 10.8, 11.1, 11.6, 11.8, 11.8, 11.3, 11.6, 11.2, 
    10.4, 10, 10.7, 11.1, 8.7, 9.3, 8.4, 6.1, 9.5, 10.5, 11.4, 11.3, 9.8, 
    7.6, 6.8, 6.9, 8.1, 6.3, 5.7, 4.3, 5, 5.3, 5.9, 6.8, 7.1, 5.6, 3.2, 8.3, 
    7.1, 5.5, 5.7, 10.1, 7.2, 7.5, 11.7, 11.4, 12.1, 11.5, 11, 12.8, 13, 
    11.6, 12.9, 11.6, 13.7, 12.7, 9.8, 11.8, 13, 12.9, 12.6, 13.2, 13.1, 
    15.8, 15.4, 14, 16.7, 15.3, 16.5, 15.9, 15.9, 15.6, 15.4, 15.9, 15.8, 
    17.2, 17.7, 15.9, 16.9, 18.7, 14.9, 15.9, 14.5, 14.3, 13, 13.7, 13.2, 
    13.7, 15.6, 15, 16, 15.3, 12.5, 13.2, 11.9, 10.4, 11.1, 10.8, 10, 10.6, 
    7.2, 2.4, 4.3, 12.7, 3.1, 1.8, 2.2, 3.3, 4.3, 2, 7.2, 6, 7.7, 5.5, 6.3, 
    5.3, 2.2, 3.6, 3.9, 2.7, 4.8, 9.9, 7, 9.9, 15, 12.5, 13.4, 14.2, 17.6, 
    18.5, 17.4, 19.4, 19.2, 18.7, 18.4, 19, 18.5, 19, 20.5, 22, 21.1, 19.4, 
    19.3, 19.6, 20.8, 19.5, 18.7, 18.6, 20.4, 21.5, 21, 21, 21.8, 22.3, 21.7, 
    21.5, 21.7, 20, 19.5, 21, 21.6, 20.3, 22.3, 22.8, 23.5, 22.2, 23.6, 23, 
    23.6, 23.4, 23.3, 22.9, 23.3, 24.4, 23.1, 23.9, 20.3, 22.3, 21.2, 21.4, 
    22.1, 22.1, 23.6, 19.5, 17.3, 15, 13.9, 12.9, 13.1, 14.8, 14.7, 13.3, 
    12.7, 12.7, 14.8, 15.2, 15.2, 15.4, 15, 16.7, 17.5, 17.5, 14.5, 15, 13.5, 
    15, 15.5, 15.4, 18.7, 18.4, 20.4, 20.6, 18.2, 19, 15.7, 15.7, 16.1, 13.8, 
    16.1, 16.2, 17.4, 14.5, 16.7, 16.4, 16.3, 16.1, 15.8, 15.7, 15.6, 15.3, 
    15, 14.3, 14, 12.1, 13, 11.4, 13.7, 14.1, 13.1, 13, 11.5, 12.6, 13.3, 13, 
    11.8, 12.7, 12.3, 11.9, 11.5, 12.2, 11, 9.9, 10.6, 9, 7.9, 6.9, 6.8, 6.3, 
    4.9, 4.3, 3.4, 3.9, 4.8, 6.4, 7.9, 5.3, 11.9, 14.3, 17.3, 19.2, 14.1, 
    18.9, 9.3, 10.4, 10.8, 9.7, 9.7, 8.8, 8.8, 7.1, 7.4, 6.8, 5.1, 5.5, 3.7, 
    2, 11, 11.7, 14.7, 18, 21.3, 21, 21.4, 21.5, 20, 19.6, 18.7, 11.9, 16.3, 
    15, 12, 14.9, 11.5, 11.4, 13.6, 13.3, 12.2, 11.7, 10.7, 10.1, 10.1, 9.6, 
    9.3, 9.1, 9.2, 7.7, 11.7, 8.7, 10.9, 10.8, 10.7, 11.2, 11.6, 9.6, 13.4, 
    11.5, 13.4, 13.4, 15.2, 14.2, 14.3, 16.8, 17, 18.3, 17.8, 21.4, 20.9, 
    21.3, 21, 19.8, 22.5, 23.1, 23.5, 21.3, 21.2, 24, 20.8, 22.7, 22.7, 23.7, 
    20.6, 18.4, 16.9, 17.2, 16.5, 13.2, 14.3, 14.1, 13.6, 12.2, 12.1, 11.3, 
    10.4, 8.1, 6.6, 5.8, 4.9, 5, 3.8, 7.1, 5, 6.7, 7.8, 12.2, 11.7, 13.9, 
    14.6, 10.9, 12.2, 9, 8, 7.7, 3.7, 4.7, 5.1, 4.1, 7.3, 6.7, 6.6, 7.4, 6.2, 
    4.2, 4.3, 5.7, 6.4, 7.6, 7.9, 8.8, 10.9, 11.2, 12.5, 11.9, 12.5, 10.8, 
    10.4, 10.6, 10.4, 11.1, 12, 11.4, 11.4, 11, 11.5, 12.9, 13.3, 15.7, 11.6, 
    15.3, 13.5, 13.3, 13.6, 12.8, 13.2, 13.7, 11.6, 12.8, 12.5, 7.2, 7.1, 
    12.3, 7.6, 6, 7.1, 7, 7.2, 10.2, 9.2, 9.4, 8.8, 14.1, 9.1, 9.1, 8.3, 
    13.5, 14.6, 12.7, 12.5, 10.8, 9.4, 11.8, 3.2, 4.3, 12.1, 5.4, 12.7, 11.2, 
    2, 3.1, 6.8, 6.5, 7.1, 9.1, 8.2, 6.8, 7.7, 7.2, 9.4, 8.9, 11.3, 12.8, 
    10.8, 10.4, 13.8, 9.6, 14.8, 11, 14.2, 6.3, 4.6, 5.3, 7.7, 9.3, 13.1, 
    13.1, 9.2, 9.1, 15.8, 10.3, 15.9, 17.3, 15.5, 8.1, 11.6, 9.2, 8, 5.2, 
    5.2, 8.2, 3, 5.6, 5.3, 2, 4.1, 7, 8.1, 8.4, 7.3, 8.1, 10.9, 14.8, 11.8, 
    12.2, 11.7, 19.1, 20.2, 13.4, 13, 19.3, 19.1, 12.1, 18.5, 12.5, 18.1, 
    16.4, 9, 13.1, 6.9, 3.6, 5.2, 6.4, 5.2, 2.7, 1.7, 0.9, 0.4, 2, 2.5, 2.3, 
    2.4, 6.8, 7.8, 11.4, 7.1, 7.6, 7.6, 7.6, 6.4, 6.7, 7.9, 4.7, 4.5, 3.6, 
    3.9, 2.3, 2.4, 0.8, 1.8, 2.9, 5.6, 4.9, 6.1, 5.6, 7.2, 8.7, 8.2, 10.2, 
    8.6, 8, 4.8, 1.2, 1.3, 1.2, 0.3, 2.7, 3.1, 0.1, 1.2, 0.9, 4.9, 3.6, 4.5, 
    6.4, 5.8, 6.8, 9.4, 10.5, 10.2, 10.5, 9.7, 10.2, 10.9, 7.7, 5.4, 7.7, 11, 
    10, 8, 6.6, 7.3, 7, 8.2, 6.4, 7.1, 7.9, 5.6, 6.8, 7.2, 5.9, 6.8, 6.4, 
    4.5, 4.4, 3.8, 4.9, 5.5, 6.2, 7.7, 7.5, 7.5, 6, 6.3, 4.9, 5.6, 6.6, 6.6, 
    6.7, 6.3, 5.8, 6.9, 5.2, 6.9, 4.8, 4.8, 4.5, 5, 6.5, 7.6, 7, 6.8, 6.5, 
    6.4, 4.3, 5.2, 4.3, 4.1, 4.2, 4.9, 5.6, 6.3, 4.7, 6.7, 7.2, 7.4, 7.7, 8, 
    8.2, 8, 7.9, 7.3, 5.6, 5, 6, 6.8, 6.3, 5.5, 5.7, 4.2, 4.1, 4.6, 5.3, 5, 
    5.7, 4.3, 4.6, 4.8, 5.5, 4.5, 4.4, 3, 3.1, 4.1, 4.2, 4.3, 4.6, 4.6, 4.8, 
    3.7, 3.6, 2.8, 2.9, 3.1, 1.6, 3.2, 3.3, 2.9, 2.2, 2.9, 2.5, 3.4, 3.3, 
    3.4, 3.3, 3.6, 3.3, 3.5, 3.3, 3, 3.5, 3.3, 3.6, 2.7, 2.8, 2.4, 2.9, 2.5, 
    2.3, 2.1, 1.8, 1.4, 2.4, 2.6, 3, 2.4, 1.2, 3.6, 5.7, 7.9, 10.5, 9.6, 8.9, 
    7.9, 7.7, 4.4, 10.4, 10.8, 10, 10.9, 11.2, 10.1, 11.9, 12.1, 11.2, 12.5, 
    13.6, 13.6, 13.6, 12.4, 11, 11.1, 11.3, 10.1, 9.8, 9.6, 8.6, 9.6, 9, 6.8, 
    10.4, 10.5, 10.5, 10.7, 12.4, 10.8, 10.1, 9.6, 7.6, 9.2, 7.9, 5.8, 4.7, 
    11.2, 10.6, 8.8, 8.1, 2.9, 3.9, 4.7, 5.1, 4, 3.3, 3.5, 3.7, 4, 4.7, 6.4, 
    8, 8.9, 11.6, 14.7, 12.6, 9.6, 9.8, 9.3, 6, 6.6, 7.3, 7.9, 8.5, 7.9, 7.9, 
    5.1, 4.3, 4.6, 7.5, 9.4, 10.9, 12.4, 11.1, 12.2, 13.3, 12.8, 12.7, 12.6, 
    13.8, 12.6, 12.4, 11.3, 10.2, 9.8, 10.3, 11.1, 11, 10.8, 12, 10.7, 11.6, 
    11.1, 9.7, 10.2, 10.4, 10.3, 10.5, 10.3, 10.3, 11.4, 12.9, 12.5, 12.6, 
    12.3, 13.4, 12, 12.5, 14.3, 11.6, 9.9, 10.3, 11.6, 12.9, 11, 11.4, 10.8, 
    10.9, 8.3, 10.1, 10.4, 10.9, 12.8, 10.7, 10.6, 8.2, 11.5, 11.7, 11.1, 
    11.2, 10.9, 10.1, 10.6, 11.6, 11.1, 11.5, 11.2, 12.4, 13.4, 12.1, 12.7, 
    11.8, 10.9, 12.2, 11.7, 12, 11.7, 11.4, 11.7, 11.8, 11.2, 11.3, 10.6, 
    10.5, 10.7, 7.9, 7.7, 8, 8.1, 8.4, 8.8, 9.3, 9.4, 8.5, 8.7, 9.4, 8.1, 
    8.4, 8.1, 7.3, 7.8, 8.4, 8.4, 8, 8.2, 6.9, 6.8, 6.2, 5.7, 6.1, 6.3, 6.5, 
    6.3, 6.5, 5.8, 4.4, 5.6, 5.4, 4.4, 4.9, 4.5, 3.8, 0.9, 1.4, 1.1, 0.7, 
    0.3, 0.3, 1.8, 2.7, 3.3, 2.7, 1.6, 4.2, 4.6, 6.4, 7.1, 7.2, 7.9, 11.3, 
    10.1, 11.9, 7.7, 6.3, 5.6, 4.6, 5.2, 4.6, 4.2, 5.3, 4.2, 4, 4.3, 4.5, 
    4.4, 3.8, 4.7, 5.7, 6, 6.1, 5.8, 4.5, 1.7, 1.6, 2.3, 2.6, 4.3, 2.3, 1.2, 
    0.8, 2.2, 2.5, 4.4, 5.1, 6.2, 7.5, 10.6, 10.2, 11.3, 11.7, 10.9, 12.5, 
    9.6, 8.1, 6.6, 6.8, 6, 4.2, 3.5, 2.8, 2.5, 2.7, 2.5, 4.1, 3.9, 3.5, 2.5, 
    2.7, 3.6, 3.7, 3.9, 3.9, 3.4, 3, 3, 2.6, 3.8, 4.9, 7.4, 7.7, 7.7, 8.5, 
    9.8, 9.6, 9.6, 9.6, 10.9, 10.7, 12.1, 13, 12.6, 11.8, 11.8, 11.8, 10.3, 
    10.7, 13.5, 13.3, 12.6, 12.4, 13.7, 12.8, 13.4, 14.3, 12.6, 13.5, 14, 
    13.7, 13.8, 13.7, 12.8, 11.9, 12, 12.4, 12.5, 11.9, 11, 10.9, 10.1, 9.6, 
    9.6, 9.8, 10.3, 10.8, 9.6, 11.1, 11, 11.3, 10.2, 8.1, 7.5, 7.1, 7.3, 7.8, 
    7.3, 8.3, 9.2, 9.5, 9, 9.1, 9.2, 7.9, 7.5, 8.8, 10.1, 12.3, 14.6, 13.1, 
    10.3, 9.9, 9, 8.4, 9.6, 8.6, 9.2, 5.7, 6.4, 7.2, 8.9, 9.4, 9.4, 9.4, 8.7, 
    10.2, 10.2, 10.3, 10.2, 9.3, 8.9, 10.6, 11.7, 12.2, 14.1, 13.6, 13.2, 13, 
    13.1, 12.6, 15, 14.1, 12.9, 15.1, 15.8, 15.4, 19.2, 19.2, 17.3, 17.7, 21, 
    24.2, 25.5, 24.5, 22.2, 22.1, 20.4, 18.2, 16.8, 14.5, 12.7, 12.2, 12.1, 
    10, 7.7, 6.7, 5.9, 7.1, 10, 10.6, 13, 15.4, 13.8, 13.6, 14.4, 14.5, 15.3, 
    15, 16, 14.3, 14.8, 14.7, 16.3, 16.5, 10.6, 19, 19.5, 19.1, 20.6, 21.1, 
    21.4, 20.3, 18.6, 14.7, 13.5, 12.7, 10.8, 10, 10.3, 14.4, 12.7, 13.3, 
    12.9, 14, 13.7, 13.1, 11.2, 9.3, 16.3, 16.7, 14.9, 11.6, 10.4, 7.7, 9.9, 
    10.1, 11.1, 11.9, 14.1, 13.9, 16.2, 19.3, 17.3, 13.9, 11.8, 13.4, 16.5, 
    17.4, 18.3, 17.5, 14, 13.7, 9.7, 11.5, 11.9, 12.9, 11.7, 12.1, 11.8, 
    11.5, 12.3, 11.6, 13.8, 14.5, 12.7, 13.7, 13.3, 9.1, 5.7, 8.5, 9.3, 12.7, 
    10.4, 21.9, 24.7, 23.5, 21, 16, 13.1, 16.4, 14.2, 12.9, 13.3, 14.9, 17.9, 
    18.9, 19.7, 14.6, 19.8, 18.6, 19.3, 19, 19.6, 19.7, 17.9, 16.4, 11.2, 
    14.5, 11.5, 9.5, 9.4, 11.1, 12.8, 21.2, 20, 19, 20.2, 20.8, 23.6, 25.5, 
    26.9, 18.1, 7, 9.1, 9.1, 10.2, 11.4, 15.4, 12.5, 15, 5.9, 1.4, 11.4, 9.9, 
    10.3, 3.7, 4.6, 6.6, 4.6, 6.8, 7.8, 6.4, 8.7, 5.7, 6.3, 9.3, 9, 8.1, 6.7, 
    6.9, 7.8, 7.8, 8, 9.5, 9.8, 10.2, 6.2, 5.1, 6.6, 4.4, 6.2, 5.4, 4.4, 6, 
    8.3, 8.2, 5.8, 4.3, 2.7, 3.9, 3.1, 1.3, 4.3, 5.1, 5.4, 5, 4.2, 2.2, 0.9, 
    1.9, 5.4, 5.5, 3.2, 4.6, 4.4, 3.1, 2.7, 1.7, 2.5, 3.4, 2.2, 2.7, 6.2, 
    6.7, 5.3, 3.5, 4.4, 3.1, 1.5, 2, 3.8, 3.3, 4.1, 4.8, 3.9, 3.8, 3.4, 4.4, 
    3.8, 4.4, 1, 3.2, 3, 3.6, 3.2, 2.9, 2.5, 3.3, 3.7, 4.5, 4.8, 3.2, 2.9, 
    4.3, 6, 2.5, 4.2, 6.6, 8, 9.2, 8.3, 8.4, 9.6, 10.2, 13.1, 13.4, 13.8, 
    15.4, 16.3, 16.8, 19.6, 13, 16.4, 21.5, 19.6, 17.5, 15.5, 19.8, 18, 18.4, 
    14.5, 12.7, 13.6, 13.2, 14.2, 16, 16.5, 14, 12.4, 13.5, 14.7, 12.2, 15.8, 
    15.7, 13.9, 13.5, 13.4, 13.7, 13.4, 13.4, 10.9, 10.7, 11.8, 10.5, 12.9, 
    11.3, 10.9, 10.3, 10.2, 9.7, 10.5, 11.2, 14.8, 15.4, 14.3, 13.5, 12.2, 
    11.6, 11, 10.2, 8.6, 8.6, 7.8, 6.5, 5.2, 2.1, 4.5, 4.8, 3.9, 3.8, 2.8, 
    2.7, 3.4, 3.8, 6.4, 5.3, 4.8, 5.2, 3.5, 2.8, 5.6, 5.6, 5.2, 5.9, 5.7, 
    4.1, 2.3, 2.7, 4.2, 4.8, 4.1, 3.5, 2.7, 3.5, 2.1, 2.1, 0.6, 0.5, 0.9, 
    2.4, 3.2, 2.4, 4.2, 3.1, 4.5, 4.1, 3.3, 3.9, 3.6, 2.4, 5.5, 3.9, 3.6, 
    3.5, 4.8, 4.4, 5.7, 5.7, 4.9, 4.8, 4.6, 3.7, 5.1, 7, 7.5, 6.2, 8.4, 8.1, 
    7.4, 7.1, 7.1, 7.6, 6.6, 6.4, 5.1, 4.3, 3.4, 3.6, 4.2, 6.1, 6.4, 7.2, 
    8.1, 8.9, 8.3, 8.8, 8.4, 7.7, 7.2, 7.2, 7.4, 9, 8.5, 9.7, 9.4, 10.2, 9.6, 
    9.2, 11.8, 12.5, 13.8, 14.9, 15.2, 16.1, 16.8, 17.5, 17.1, 17.5, 17, 
    16.9, 17.5, 18.2, 17.8, 17.8, 18.3, 18.3, 18.2, 17.7, 17.2, 16.7, 16.4, 
    17.6, 16.5, 17.1, 17.2, 16.9, 16, 16.6, 15.1, 14.9, 14.2, 14.8, 15.1, 
    14.9, 14.1, 16, 15, 13.4, 11.9, 13.2, 12.1, 11.9, 11.6, 9.1, 8.6, 10.2, 
    10.9, 11.9, 9.9, 8.6, 10, 11.2, 8.6, 8.5, 9.8, 12.7, 12.1, 9.2, 7.5, 7.8, 
    7.1, 5.6, 5.6, 5.9, 5.3, 6.2, 7, 7.7, 6.4, 5.6, 6.5, 4.8, 3.1, 2.5, 2.5, 
    2.5, 3.3, 4.7, 3.6, 5, 6.2, 7.9, 8.7, 10.5, 10.3, 9.6, 9, 9.1, 10.2, 9.6, 
    10, 10.3, 8.4, 9.1, 9, 9.5, 10.3, 11.3, 12.3, 12.4, 11.3, 14.8, 16.1, 
    15.8, 16.9, 17.1, 16.6, 16.4, 15.5, 14.9, 12.3, 10.3, 9.8, 9.6, 10.1, 
    9.1, 6.9, 5.5, 5.5, 5.1, 5.4, 4.4, 3, 4.5, 4.4, 5.9, 6.2, 7, 7.3, 7.5, 
    7.4, 6.5, 6.7, 5.9, 5.6, 7.5, 7.9, 6.6, 5.9, 4.4, 5.2, 5, 6.1, 6.9, 6.5, 
    5.4, 4.4, 4.7, 3.3, 3.8, 2.2, 2.5, 3, 3.4, 2.2, 3.5, 3.3, 3.1, 0.4, 5.1, 
    7.6, 6.2, 5.9, 6.8, 8, 9, 10.5, 11.4, 9, 9.1, 10.3, 9.4, 8.7, 8.6, 8, 
    8.6, 8.7, 8.7, 9, 8.8, 9, 8.9, 9.6, 9.9, 9.1, 9.8, 9.7, 9.3, 10.1, 10.6, 
    9.8, 9.7, 8.6, 4.8, 9, 7.4, 7.8, 7.1, 7, 6.7, 5.1, 8.1, 9.9, 9.3, 6.5, 
    9.3, 9.2, 9.6, 11.1, 10.5, 9.2, 7.7, 7.5, 6.5, 6.2, 6.4, 5.7, 4.6, 3.9, 
    3.9, 3.9, 2.9, 3.4, 3.6, 3.6, 3.6, 4.4, 4.7, 4.7, 4.3, 4.8, 4.3, 5.3, 
    5.6, 6, 6.4, 7.3, 5.6, 5.8, 5.9, 4.8, 3.7, 3.8, 3.7, 4.1, 4, 5, 3.9, 3.6, 
    4.8, 5.3, 4.6, 5.4, 3.6, 4.3, 5, 7.2, 4.9, 3, 4.9, 5.4, 7, 5.2, 8, 8.2, 
    7.4, 7.7, 10, 8.6, 7, 6.1, 6.6, 6.7, 7.2, 7, 7.9, 5.8, 8.4, 8.1, 5, 8.1, 
    6.4, 7.1, 6.2, 6.6, 6.7, 3.2, 2.4, 0.9, 1.4, 0.8, 1.9, 1.3, 1.7, 1.5, 
    0.6, 2, 1.9, 1.3, 1.3, 1.9, 1.7, 1.4, 3.9, 4.9, 4, 5.8, 5.4, 6.2, 8.5, 9, 
    9.2, 8.5, 9.9, 7.6, 7.9, 8.8, 7.9, 8.9, 10.1, 9.5, 9.7, 9.1, 8.3, 4.4, 
    6.3, 2.6, 6, 5.5, 5.2, 3.8, 5, 4.5, 2.9, 2.6, 4.6, 5.7, 9.3, 10.3, 9.8, 
    8.4, 8.7, 8.6, 8.1, 8.3, 9.6, 8.9, 9.9, 9.5, 9.1, 7.6, 7.6, 8.9, 9.6, 
    9.9, 11.7, 12, 12.3, 11.4, 11.6, 11.6, 10.9, 10.8, 10.5, 8.4, 8.3, 8.2, 
    9.1, 9.3, 11.1, 12.4, 12.8, 13.4, 14.9, 16.9, 17.4, 16.8, 17.6, 16.3, 
    15.5, 13.6, 12.9, 8.8, 8.9, 10.8, 11.1, 12.2, 13.8, 16.1, 19.2, 20.9, 
    20.2, 19.3, 19.6, 18.4, 19.5, 19, 18.7, 18.1, 16.1, 15, 14.3, 13, 12.5, 
    12.3, 13.2, 14, 14, 14.3, 15.6, 15, 15.4, 16, 15.6, 16.4, 17, 16.5, 16.9, 
    15.6, 14.4, 14.7, 14.6, 14.5, 14.8, 14.4, 14.5, 14.7, 15.3, 15, 13.7, 
    12.9, 11.7, 13.2, 12.7, 12.7, 12.8, 12.5, 12.3, 12.2, 11.5, 12.4, 10.1, 
    10, 10.4, 10.5, 9.7, 8.3, 8, 5.7, 5.4, 4.7, 5.6, 6.4, 6.8, 5.9, 6.2, 7.3, 
    6.9, 5.7, 4.8, 4.4, 1.5, 2.3, 1.4, 3.5, 5.3, 4.8, 4.3, 1.5, 4.8, 3, 2.8, 
    1.3, 0.8, 0.1, 0.5, 0, 0.9, 4.1, 2.2, 2.2, 0.9, 2.6, 2.2, 1.2, 2.2, 3.3, 
    3.6, 4.2, 4.3, 3.1, 2.9, 2.3, 4, 4.7, 5.2, 4.1, 3.8, 3.4, 3.4, 2.7, 2.7, 
    5.5, 5.4, 5.4, 1.8, 4.6, 2.5, 3.1, 3.4, 5.8, 6.1, 5, 6.9, 6.5, 6.5, 4, 
    6.9, 6.3, 7.2, 7.1, 4.7, 4.4, 4.3, 4.2, 6.4, 6.6, 6.2, 6.9, 8.1, 8.7, 8, 
    6.6, 5.5, 6.2, 6.5, 4.6, 6.6, 5.9, 6.6, 7.1, 7.7, 7, 7.6, 8.7, 5.7, 7.9, 
    8.7, 11.6, 11.9, 10.7, 7.2, 6.8, 8.6, 8, 10.3, 9, 7.2, 5.6, 6.3, 5.8, 
    6.2, 8.5, 6.9, 5.9, 7.5, 7.8, 8.6, 8.6, 9.6, 9.3, 9.4, 9, 9.2, 8.8, 8.4, 
    7.2, 7.9, 8.9, 5.7, 4.6, 3.3, 3.5, 0.8, 1.3, 1.1, 1.5, 3.4, 4, 4.3, 5.7, 
    2.7, 1.6, 0.7, 1.4, 2.3, 1.9, 2.9, 3.5, 3.1, 3.7, 3.6, 3.8, 5.5, 5.6, 
    5.1, 6.2, 8, 9.8, 10.7, 11.3, 10.3, 9.7, 9.8, 10.5, 10.6, 10.4, 10.6, 
    11.3, 11.5, 11.4, 11.2, 12.2, 11.3, 10.5, 10.6, 10.1, 9.9, 9.7, 10.4, 
    6.8, 6.1, 6.9, 4.4, 4.1, 3.7, 3.5, 7.7, 3, 4.1, 3.6, 4, 3.4, 6.7, 6, 5.4, 
    4.3, 5.4, 6.1, 7.6, 5.4, 5.3, 5.5, 5.9, 6.7, 8.5, 10, 11.3, 12.7, 12.5, 
    12.5, 12.9, 11, 9.5, 6, 5.4, 6.3, 8.9, 7.2, 5.5, 2.7, 3.3, 1.4, 7.6, 
    14.8, 14.2, 15.3, 16.5, 16.2, 15.3, 13.7, 13.8, 13.4, 11.5, 9, 8.2, 5.8, 
    4.5, 1.7, 2.3, 6.3, 6.9, 9, 11, 11.5, 14.2, 14.3, 14.9, 13.2, 13.1, 11.2, 
    12.7, 13.4, 13.3, 12.2, 15.1, 14.4, 16.4, 13.3, 12.8, 14.2, 13.4, 13.4, 
    14.1, 14, 14.4, 14.5, 15, 16.6, 15.5, 14.7, 13, 10.8, 10.9, 10.4, 12.4, 
    10.7, 11.1, 11.9, 11.7, 11.3, 11.8, 12.9, 12.2, 13.4, 12.6, 11.6, 12.9, 
    14.1, 14, 13, 13.5, 12.9, 11.1, 12.1, 12.5, 12.1, 12.4, 13.4, 13.2, 13.6, 
    12.8, 14.2, 13.8, 14, 13.4, 12.4, 11.6, 11, 12.7, 13.8, 12.7, 12.8, 15.4, 
    15.2, 16.1, 17, 16.3, 16.9, 18.3, 16.4, 12.4, 13.4, 13.5, 12.2, 12.5, 
    10.1, 10.8, 11.6, 12.5, 12.5, 12.4, 11.7, 11.8, 13.4, 11.5, 12.2, 10.3, 
    10.5, 10.3, 11.8, 14, 13.6, 12.3, 12.2, 12.2, 11.4, 9.7, 9.3, 9, 7.3, 
    5.6, 5.2, 5.8, 5.8, 8.8, 11.5, 11, 10.5, 9.4, 7.1, 8.2, 6.4, 6.1, 6.2, 
    8.1, 9.1, 7.8, 9.5, 8.6, 4.5, 6, 10.2, 12, 13.5, 12.5, 13.2, 12.9, 12.2, 
    9.4, 11, 11.8, 14.3, 13.7, 12.1, 12.3, 10.9, 13.3, 15.3, 14.9, 13.3, 12, 
    14.2, 11.3, 14.3, 14.4, 14.7, 14, 13.3, 12.9, 12.1, 11.4, 11.9, 11.6, 
    10.5, 10.7, 9.8, 9.7, 9.2, 9.6, 8.8, 8.3, 8.6, 8.3, 8.2, 7.8, 7.7, 8.2, 
    7.1, 7.4, 6.9, 7.6, 6.2, 3.5, 2.9, 7.3, 4.5, 5.6, 4.9, 4.9, 3, 3.5, 4.9, 
    6.8, 0.7, 5.1, 6.6, 3.1, 5, 1.9, 6, 5.5, 4.4, 3.3, 2.4, 1.2, 1.3, 1.7, 
    1.7, 1.3, 2.2, 6.1, 5.9, 3.6, 1.4, 1.8, 3.2, 2.9, 3.5, 1.4, 1.4, 1.7, 
    2.1, 1.4, 3.5, 3.2, 2.9, 2.9, 3.3, 5.7, 1.6, 4.1, 3.8, 3.1, 2.5, 1.4, 
    2.5, 3.6, 2.9, 4.8, 5.3, 3.7, 4.3, 2.3, 1.3, 0.6, 1.4, 7.1, 7.6, 13.8, 
    13.5, 13.3, 11.1, 6, 10.7, 11.3, 11.2, 10.6, 11.2, 12.6, 12.9, 13.6, 
    14.4, 14.9, 13.4, 13.2, 13.2, 12.5, 11.9, 11.8, 10.6, 9.2, 8.9, 8, 6.4, 
    6.9, 6.2, 5.4, 4.2, 2.1, 0.8, 5.6, 8, 4.4, 8.1, 9.5, 9.7, 8.5, 9.6, 10.4, 
    9.7, 10.9, 9.6, 10.2, 9.4, 10.1, 9.6, 5.9, 10.5, 10.8, 11.2, 11.9, 11.5, 
    11.4, 12.7, 13.3, 12, 14.2, 14.1, 13.8, 15.6, 16.1, 18.9, 19.6, 19.2, 
    18.1, 19.9, 20.7, 22.4, 24.2, 24.5, 24.4, 21.8, 21, 19.4, 18.2, 17.9, 
    18.2, 18.4, 17.4, 14.8, 17.2, 16.8, 17.2, 16.9, 17.2, 21, 20.8, 18.7, 
    15.8, 16.1, 13.1, 12.7, 14.8, 14.7, 14.8, 12.9, 12.4, 11.6, 14, 13.6, 
    9.6, 13.7, 14.2, 13.2, 6.2, 5, 4.4, 5.3, 5.5, 6, 6.3, 6.8, 5, 5.4, 6.7, 
    7.5, 8.3, 6.7, 7.1, 6.9, 7.6, 7.7, 8.9, 7, 8, 7.1, 6.9, 8.1, 6.3, 9.4, 
    5.2, 6.4, 4.9, 7.1, 8.4, 8.8, 8.8, 9, 7.6, 9.1, 10.1, 9.9, 11.1, 10.5, 
    9.9, 9.8, 10.3, 10.3, 10.1, 10.6, 10.6, 7.5, 10.2, 11.1, 12.6, 11.9, 9.7, 
    7.6, 9.4, 11.4, 10.6, 12.1, 11.3, 11.5, 11.2, 11.2, 12.6, 11.2, 10.9, 
    11.4, 10.2, 9.6, 9.8, 10.2, 7.3, 5.7, 4, 6.3, 6.8, 7.1, 7.2, 7.1, 6.7, 
    6.2, 5.1, 4.4, 4.2, 3.2, 1.5, 1.1, 1, 1.4, 5.6, 2.3, 3, 3, 3.6, 3.4, 3.6, 
    3.3, 2.1, 4.1, 3.4, 3.7, 3.6, 3.9, 5, 3.6, 4.8, 5.2, 4.9, 3.9, 3.9, 4, 
    4.7, 4.5, 4, 4.1, 3.6, 4.3, 3.2, 3.2, 3, 4.9, 3, 2.6, 2.6, 2.6, 2.2, 1.7, 
    3.4, 2.2, 0.5, 1.4, 3.4, 2.6, 1.8, 3.2, 3.3, 2.9, 3.4, 3.7, 2.6, 3.7, 
    2.8, 3.7, 3, 3.9, 2.1, 1.3, 4.6, 4.7, 6.1, 4.3, 5.7, 6.5, 6.7, 6.7, 8.3, 
    8.8, 9.5, 11.1, 10.1, 11.6, 12, 3.5, 10.7, 9.6, 7.1, 8.2, 7, 6.8, 7.6, 
    5.7, 3.7, 5, 6.5, 5.1, 3.6, 2.8, 0.6, 1.4, 1.5, 2.9, 1.3, 1.8, 0.4, 1.4, 
    1.3, 1.3, 1.1, 2.2, 4, 3.5, 2.4, 3.1, 2.3, 0.5, 0.4, 0.7, 1.8, 2.2, 3.2, 
    4.6, 3.9, 5.9, 6.4, 3.5, 5, 5.1, 4.9, 5.9, 5.6, 5.4, 4.9, 4.2, 5.6, 6.1, 
    4.2, 5.1, 5, 2.1, 1.3, 2.6, 2.3, 3.8, 4, 4.4, 3.2, 2.6, 4.7, 4.4, 5.1, 
    4.6, 4.8, 6, 7.5, 4.7, 1.3, 1.9, 0.4, 1, 8.3, 8.5, 8.1, 6.6, 6.5, 5.7, 
    4.8, 5.6, 4.1, 5.3, 4.4, 3.9, 3.5, 4.6, 3.7, 4.5, 3, 6, 2.8, 5.1, 4.3, 
    2.8, 2.5, 3.3, 3.6, 3.1, 4, 2.7, 2.5, 3.5, 2.2, 0.1, 10.7, 12.1, 10.5, 
    8.9, 9.8, 8.7, 12.1, 10.9, 10.4, 9.2, 8.5, 7.7, 8, 6.9, 6.9, 8, 8.8, 8.8, 
    12.5, 11.5, 9.9, 10.3, 10.7, 10.2, 10.2, 9.7, 10.3, 11, 11.2, 12.5, 11.5, 
    14.5, 14.8, 17.1, 16.7, 16, 17.2, 17.8, 16.6, 17, 16.7, 15.4, 15.6, 14, 
    13.4, 13.9, 9.6, 12.2, 13.8, 12.8, 12.6, 13.5, 13.5, 14.7, 14.2, 14.6, 
    13, 13.9, 14.1, 13, 13, 12.3, 12.7, 12.2, 13.9, 12, 13, 13.8, 15.4, 17.7, 
    13.2, 12, 10.9, 11.8, 11.9, 10.6, 11.7, 11.4, 12, 13, 14.7, 14.1, 15.2, 
    14.4, 14, 13.4, 11, 12.2, 11, 11.4, 11.5, 10.6, 11.6, 11.9, 10.8, 12.2, 
    13.7, 15.2, 12.6, 11, 12.4, 12.5, 11.1, 12.3, 11, 10.8, 8.5, 9.7, 9.2, 
    10, 11.1, 12.1, 12.4, 9, 12.3, 11.2, 11, 11.9, 6.2, 4.6, 9.3, 8.7, 8.8, 
    9.6, 10.4, 8.4, 10.5, 10.6, 12.2, 11.4, 10.1, 11.3, 8.6, 7.6, 7.6, 9.6, 
    11.3, 12, 12.4, 12.4, 12.6, 9.5, 7.2, 7.8, 8.1, 10.7, 11.4, 13.8, 12.5, 
    6.8, 7.1, 7.7, 9.8, 7.1, 8.5, 7.5, 8.2, 10.2, 9.8, 11, 11, 8.5, 8.1, 8.4, 
    9, 7.3, 6.8, 6.7, 7.5, 5.4, 7.4, 7.8, 8.6, 6.9, 8.4, 8.7, 8.1, 6.7, 7, 
    4.4, 4.2, 7.3, 6.6, 6, 5.4, 6.1, 5, 5.2, 6.6, 5.6, 4, 2.8, 2.4, 4.1, 4.1, 
    5, 4.4, 4.4, 4.2, 3.1, 3.5, 5.9, 5.7, 7.3, 7.1, 7.2, 10.4, 11.2, 12.5, 
    11, 12.1, 11.2, 9.5, 6.7, 4.6, 10.1, 10.5, 10.2, 9.2, 9.6, 9.9, 9.3, 9.9, 
    11.1, 10.9, 8.7, 7.8, 6.5, 7, 6.5, 5.8, 5.8, 6.4, 6.5, 5.4, 5, 7.8, 7.6, 
    8, 8.4, 7.7, 5.9, 7.9, 8.8, 8.6, 8.2, 8, 8.2, 9.9, 11.7, 10, 10.7, 9.8, 
    14.8, 16, 10.2, 16.7, 14.1, 11.8, 11.3, 8.7, 8, 8.8, 9.8, 9.2, 9.4, 10.2, 
    10.8, 9, 8.8, 8.1, 7.8, 7.5, 7.8, 7.7, 7.9, 6.9, 7.2, 7.4, 7.7, 6.6, 6.8, 
    6, 6.1, 5.6, 4, 3.8, 3.2, 2.2, 2.2, 1.9, 1.4, 5.7, 2.9, 4.1, 2.3, 6, 8.3, 
    9, 10, 10.1, 11.6, 13.6, 14.2, 13.9, 15.3, 13.6, 13, 12.8, 14, 13, 13.4, 
    13.5, 7.8, 12.2, 10.9, 9, 9.4, 8.6, 10, 9.9, 9.1, 8.2, 5.5, 4.4, 3, 7.7, 
    3.2, 1.6, 2.9, 3.5, 5.8, 6.1, 7.4, 8.1, 8.7, 8.5, 10.5, 11.6, 10.2, 8.2, 
    8.8, 9.4, 10, 10.4, 9.8, 8.5, 7.8, 8.2, 7.7, 7.5, 8.4, 9.7, 8.8, 8.6, 
    9.2, 10.3, 11.6, 11.2, 11.8, 10.3, 9.4, 10.5, 11.1, 13.2, 14.5, 10.9, 
    10.7, 12.9, 13.9, 14.6, 15.1, 13.4, 12.7, 12.3, 12.3, 11.2, 11.8, 12.1, 
    11.5, 11.2, 11.8, 9.8, 9.2, 7.9, 7.3, 6.5, 6.5, 5.9, 5.1, 4.7, 4, 2.7, 
    1.5, 1.2, 1.3, 4.5, 4.5, 5.1, 4.6, 4.4, 3, 4.7, 4, 5.4, 6.1, 5.4, 6.2, 
    7.2, 8, 8.3, 8.7, 11.7, 11.7, 11.5, 9.4, 6.5, 10.1, 2.4, 11.2, 6.2, 5.1, 
    2.9, 3.6, 0.2, 1.4, 1.1, 3.2, 1.2, 2.4, 0.8, 0.5, 3.1, 0.9, 0.2, 1, 1.4, 
    0.9, 1.4, 0.6, 0.7, 0.8, 0.8, 0, 0.7, 0.1, 0.7, 0.8, 2.3, 5, 3.9, 2.4, 
    1.8, 0.7, 2.1, 6.2, 6.5, 6.9, 6.6, 4.9, 5.3, 4.7, 6.8, 6.5, 7.1, 7.3, 
    7.2, 6.7, 5.5, 6.4, 4.4, 4.1, 4.4, 3.1, 0.9, 0.5, 0.5, 1.9, 2.3, 2.2, 
    0.7, 3.4, 3.1, 3.6, 3.3, 4.5, 4.6, 4.6, 3.5, 1.8, 2.8, 2.6, 1, 1.1, 1.9, 
    2.5, 2.4, 1, 2.3, 3.7, 5.4, 6.5, 6.7, 7, 7.3, 7.6, 7, 7.7, 6.9, 6.3, 4.2, 
    2.1, 4.1, 4.2, 3.1, 2.4, 2.9, 1.5, 0.2, 1.8, 6.1, 8.3, 8.6, 8.3, 8.7, 
    8.9, 8.1, 9.4, 8.3, 7.9, 7.6, 10, 12.1, 10.2, 9.4, 9.3, 8.4, 8.9, 7.4, 
    6.9, 6.1, 5.9, 6.6, 7.2, 7, 7.1, 6.5, 5.7, 4.6, 5.1, 3.8, 4.9, 4.4, 4.5, 
    2.8, 3.1, 3.2, 3.8, 7, 3.4, 2.7, 3.3, 1.4, 3.5, 2.4, 2, 2.2, 2.7, 1.3, 
    2.8, 3.4, 3.6, 3.7, 3.7, 3.8, 4.2, 3.5, 3.5, 3.5, 4.1, 3.9, 4.5, 4.4, 
    7.7, 5.6, 6.1, 5.2, 5, 4.3, 4.3, 3.4, 3.1, 2.9, 2.1, 1.6, 1.8, 1.8, 2.6, 
    2.9, 3.9, 3.9, 5.1, 5.7, 6.5, 7.3, 6.8, 7.1, 7.1, 7, 6.2, 6.5, 6.3, 7.3, 
    6.8, 6.9, 5.4, 6.5, 6.8, 5.4, 6, 6, 5.7, 6.6, 6.1, 7.7, 4.1, 8.3, 7.4, 
    6.2, 7.2, 8.3, 8.4, 8.8, 8, 8.1, 8.4, 8.7, 8.4, 8.7, 8.4, 9.3, 9.8, 9.1, 
    10, 10.6, 10, 10.7, 10.2, 10, 10.3, 9.2, 9.5, 9.7, 9.8, 9.5, 8.6, 9, 8.5, 
    9.4, 8.5, 9, 8.6, 8.5, 9.6, 10.2, 11.6, 13.1, 15.1, 14, 13.3, 11.5, 10.3, 
    9.9, 9.1, 10.6, 11.1, 10.9, 11.1, 11.3, 12.3, 12.7, 12.6, 13.3, 12.3, 
    12.3, 10.2, 11.6, 14.6, 13.3, 13.5, 12, 12.9, 12.6, 9.3, 9.9, 11, 10.2, 
    7.9, 6.3, 8.1, 9.3, 8.9, 8.5, 7.1, 6.2, 6.4, 6.8, 6.6, 5.8, 8, 7, 6.1, 
    6.6, 6.4, 6.6, 6.9, 7.2, 7.5, 7.6, 7.9, 7.7, 7.8, 9.1, 8.8, 7, 7.4, 6.9, 
    6.9, 6.2, 6.1, 6.6, 6.4, 6.5, 6.8, 7.5, 6.2, 6.2, 5.8, 6, 6.4, 5.8, 6.3, 
    6.4, 6.5, 7.2, 7.1, 6.9, 6.9, 7.5, 7.4, 7.2, 7.3, 7.5, 9.2, 8, 7.8, 8.6, 
    8.3, 9.3, 8.4, 9.7, 9.5, 10.5, 10.2, 10.5, 10.2, 12, 10.7, 10.1, 10.7, 
    11, 11.8, 12.8, 13.9, 12.8, 12.2, 14.3, 15.7, 15, 15.3, 14.6, 14.5, 14.2, 
    14.9, 13.2, 13.3, 12.6, 12.1, 11.3, 10.3, 9.9, 10.5, 11.4, 11.6, 11.1, 
    11.8, 10.3, 10.3, 10.3, 9.4, 8.8, 8.9, 10.3, 10, 10, 10.2, 10.9, 11.6, 
    11.5, 10.9, 10.9, 10.3, 10.6, 9.8, 10, 9.7, 9.7, 9.2, 9.8, 10.1, 10.4, 
    9.3, 10, 9.5, 10, 10.4, 10.4, 11.3, 11.8, 12.3, 12.6, 12.4, 13.8, 13, 
    13.5, 14.1, 14.4, 13.8, 15, 16.1, 17.1, 18.2, 17.6, 17.4, 18.8, 19.8, 
    19.1, 18.3, 17, 14.9, 13.6, 12.1, 12.7, 11, 11, 9.8, 10, 10.1, 9.8, 10.6, 
    10.5, 11.3, 11.3, 10.4, 10.5, 9.7, 7.2, 6.9, 7.4, 7.5, 4.9, 3.3, 4.3, 
    3.7, 2.9, 7.2, 12.1, 13.5, 10, 14.3, 15, 15.7, 13, 13.3, 11, 2.8, 5.1, 
    5.1, 7.5, 4.8, 2.4, 4.2, 6, 5.8, 2.9, 1.3, 1.2, 2, 3.3, 1.1, 1.2, 0.4, 
    4.8, 3.3, 4.4, 4.5, 5.2, 2.7, 2.4, 3.1, 1.8, 3.3, 2, 2.5, 2.9, 2.8, 1.5, 
    2.3, 4.1, 4.2, 4.3, 4.5, 4, 4.8, 4.4, 6.1, 4.2, 4.8, 4.5, 5.5, 4.6, 4.3, 
    4.6, 4.6, 5.4, 5.7, 4.2, 5.3, 3.5, 3.4, 5.3, 3.3, 3.3, 4.1, 5.4, 5.5, 
    7.9, 8.3, 8.6, 6.4, 5.7, 6.3, 5.6, 5.2, 3.5, 3.4, 2.5, 2.5, 3.7, 2.8, 
    4.5, 3, 5.7, 6.1, 6.6, 5.7, 5.1, 5.6, 5.7, 3, 4.5, 2.9, 3.6, 5.4, 5, 4.5, 
    3.5, 2.4, 3.3, 6.3, 7, 5.8, 5.8, 7.7, 7.8, 12.3, 11.6, 12.1, 12.8, 13.4, 
    13.7, 14.1, 11.9, 10.5, 8.7, 7.3, 7.9, 6.4, 4.1, 2.4, 2, 1.6, 1.7, 4.9, 
    2.9, 4.2, 4.9, 5, 4.9, 4.4, 4.5, 5.3, 4.8, 5.1, 3.5, 2.7, 0.9, 3.3, 3.7, 
    3.3, 3.6, 4.6, 4.9, 4.9, 5, 5, 4.9, 4.9, 4.6, 5.6, 6, 6.5, 5.6, 6.4, 6.1, 
    5, 4.5, 4.9, 6.4, 7.8, 8.6, 9.1, 9.6, 9.4, 8.1, 8.6, 7.5, 7.5, 8, 6.7, 
    7.4, 6.9, 7.2, 7.8, 8.5, 6.1, 5.1, 5.3, 7.7, 10, 12.7, 11.7, 10.7, 11.1, 
    11.4, 5.1, 5.6, 3.5, 4.1, 4.6, 6.2, 12.1, 14, 17.8, 15.5, 15.6, 15, 14.3, 
    11.9, 13.7, 12.8, 11.7, 8, 11.2, 10.9, 12.2, 10.7, 1.3, 3.4, 3.3, 5.1, 
    8.3, 7.2, 9, 8.9, 6.1, 7.4, 8.9, 7.9, 6.8, 6.1, 6.9, 5.9, 4.4, 5.1, 6.1, 
    5.8, 5.7, 6.9, 6.7, 6, 5.2, 4.6, 4.9, 3.9, 3.2, 2.1, 2, 2.1, 1.2, 3.4, 
    3.2, 3.6, 3.9, 4.5, 5.1, 6.3, 6.9, 7.8, 7.7, 8.6, 8.9, 10.4, 11.2, 12, 
    12.3, 11.8, 11.3, 13.6, 13, 12.5, 13.8, 14.9, 16, 16.5, 16.6, 16.8, 14.4, 
    16.9, 15.6, 16.4, 15.9, 15.1, 13.2, 10.2, 9, 7.2, 7, 6.8, 7.7, 7.6, 6.5, 
    5.2, 4, 2.5, 1.6, 2.9, 2.5, 4.7, 7.4, 8.7, 9.3, 9, 7.7, 10.9, 7.4, 8.5, 
    10, 8.8, 5.3, 5.1, 5.4, 4, 3.4, 3.9, 4.2, 5.4, 3.9, 3.3, 2.4, 3.9, 3, 
    2.3, 1.4, 1.4, 0.9, 1, 0.8, 0.2, 0.2, 0.8, 1, 2.7, 3.7, 4.4, 4.1, 3.8, 
    4.1, 4.3, 4.8, 5.3, 5, 5.9, 5.2, 4.9, 4, 4, 3.6, 3.7, 4.2, 3.4, 3.9, 4.4, 
    4.4, 4.5, 4.6, 5.7, 5.9, 6.3, 6.3, 7, 7.8, 7.2, 6.2, 7.7, 7.6, 7.1, 6.6, 
    6.4, 6.3, 4.9, 5.4, 4.7, 4.5, 3.5, 4.2, 3, 1.4, 2.9, 1.7, 1.1, 8.1, 9.2, 
    12.4, 13.6, 15, 15.7, 12.8, 13.4, 11.3, 11.6, 10.5, 3, 4.4, 3.9, 4.1, 5, 
    6.4, 6.2, 6.5, 6.2, 7.2, 5.9, 6.5, 8, 7.2, 6.5, 5.2, 6.2, 6.6, 8.3, 8.7, 
    8.1, 9.1, 9.5, 10.1, 11.9, 11.3, 11.9, 10.7, 11.3, 11.7, 11, 11.9, 11.2, 
    10.9, 12.8, 14.5, 16.2, 14.4, 13.3, 13.5, 12.4, 13.1, 13.4, 12.7, 11.3, 
    11.4, 12.3, 10.6, 11.5, 11.2, 11.8, 11.5, 11.6, 12.9, 14.5, 14.9, 13.8, 
    14.4, 13.6, 13.4, 11.5, 11.7, 11.9, 12.9, 12.7, 12.3, 11.3, 12.9, 14.9, 
    17.2, 17.2, 13.6, 13.6, 13.7, 11.9, 11.1, 9.7, 10.3, 10.2, 12.4, 9.3, 9, 
    10.5, 7.9, 8.9, 10.2, 8.6, 8.4, 8.7, 9.5, 9.5, 8.4, 7.7, 9.7, 10.8, 7, 
    7.3, 7.9, 8.4, 8.6, 9.9, 9.3, 10.3, 8.7, 8.9, 9.6, 7.9, 9.3, 9.1, 10.7, 
    9.6, 6.4, 9.3, 9.5, 8.8, 7.3, 7.6, 6.9, 8.6, 7.6, 8.1, 7.6, 8.1, 9.1, 8, 
    6.8, 7.6, 8, 9.8, 7.9, 6.9, 6.7, 8, 8.1, 8.4, 7.5, 8.4, 7.3, 7.4, 7.4, 
    6.8, 8.4, 6.7, 8.3, 9, 8.9, 8, 7.7, 8.4, 10.2, 9.9, 9.1, 7.8, 8, 8.4, 
    8.3, 8.1, 8.2, 8.2, 8.6, 8.3, 8.5, 9.2, 10.1, 9.3, 9, 9.6, 7.8, 8.3, 8.9, 
    9.7, 9.8, 9.4, 8.9, 8.6, 8, 6.7, 7.1, 5.4, 6.4, 6.4, 6.3, 7.6, 6.3, 5.9, 
    6, 6, 7.3, 4.9, 6.8, 7.3, 7.9, 7.7, 8.2, 8.4, 11.9, 9.6, 9.6, 9.8, 9.2, 
    10.9, 11.2, 9.9, 9.9, 11.8, 11.3, 9.4, 8.6, 10.1, 9.8, 9.4, 8.5, 4.7, 
    9.3, 5.9, 9.8, 7.7, 7.8, 7.5, 5.8, 10.3, 5.8, 11.2, 9.1, 13.5, 10.9, 
    12.8, 10.6, 10.5, 8.9, 10.5, 10.6, 7.5, 8.6, 7.5, 7.7, 9.4, 9.7, 9.4, 
    8.9, 10.2, 9.4, 7.6, 7.8, 9.1, 8.4, 8.2, 8.5, 7.8, 7.9, 8, 7.7, 7.4, 8.1, 
    7.7, 6.1, 5.4, 6.3, 5.7, 4.2, 4.6, 3.5, 5.8, 2.4, 3, 3, 3.7, 4.9, 4.7, 
    4.3, 3.9, 3.7, 5.9, 3.5, 5.9, 2.3, 2.3, 6.3, 6, 2.4, 5.5, 1.3, 4.8, 0.7, 
    4.4, 1.1, 1, 4.2, 1.6, 2.9, 2.4, 2.5, 4.2, 3.3, 3.5, 4.8, 3.8, 4.8, 3.3, 
    2.9, 5.2, 2.9, 4.7, 4.1, 4.1, 4.9, 4.3, 4.5, 4.4, 6, 5.6, 5.7, 5.4, 5.7, 
    5.7, 4.1, 2.5, 4.4, 3.5, 4.9, 2.9, 1.9, 4.8, 0.7, 6.6, 7.3, 0.6, 2.2, 2, 
    2, 5, 8, 10.8, 15.7, 11.4, 13.7, 11.2, 12.9, 17, 12.7, 18.1, 19.2, 18.3, 
    18.1, 7.6, 7.1, 15.7, 6.2, 10.8, 5.5, 10.9, 10.7, 11.2, 5.8, 6.2, 13.1, 
    8.2, 13.3, 13.8, 9.8, 13.8, 14, 14.4, 14.7, 10.8, 15.9, 16.7, 15.6, 13.8, 
    12.3, 12.2, 11.8, 11.6, 11.6, 12.1, 10.7, 11.9, 9.8, 10.3, 10.5, 9.2, 9, 
    9, 9.1, 8.4, 7.1, 6.6, 6.3, 6.4, 6.8, 6.4, 6.6, 6, 6.3, 6.9, 6.6, 8.6, 
    7.9, 7.3, 8.4, 7.5, 9.2, 6.5, 5.6, 6.8, 7.9, 6.1, 7.8, 7.8, 8.1, 7.7, 
    5.6, 6.8, 4.7, 4.6, 8.6, 4.6, 2.3, 0.9, 1.2, 3.5, 3.4, 3.7, 4.1, 4.9, 
    5.9, 8.3, 7.8, 8, 8.3, 7.7, 9.9, 8.6, 8.4, 9.5, 9, 11.4, 9.3, 8.4, 8, 
    7.5, 11.2, 11.6, 8.7, 7.2, 4.7, 5.5, 6.7, 9.2, 7.2, 5.3, 6.5, 4.8, 5.7, 
    5.2, 5.3, 4.2, 5.7, 5.1, 4.9, 4.1, 1.5, 2.5, 3.6, 2.1, 3.1, 3.8, 2.8, 
    4.6, 4.1, 2.6, 3, 1.5, 2.2, 6.7, 7, 6.8, 3, 3.9, 2.1, 2, 3.6, 4.5, 6, 
    4.7, 5.6, 3.8, 5.9, 5.3, 6.4, 6.3, 3.9, 2, 5.2, 0.7, 0.9, 0.4, 1.2, 3.2, 
    3.5, 1.9, 4.5, 3.1, 4.5, 3.8, 4.3, 2.7, 2.9, 5.4, 2.8, 3, 2.5, 2.4, 2.5, 
    2.5, 5.5, 5.2, 5.4, 5.7, 6.5, 8.6, 7, 8.4, 7.7, 6.6, 6.8, 7.1, 7.7, 9.3, 
    8.6, 8.1, 7.9, 7.7, 8.3, 8.1, 5.3, 1.6, 2.9, 2.8, 3.1, 3.3, 3.7, 2.9, 
    0.6, 0.8, 2.1, 3.4, 4.7, 6.1, 6.9, 5.6, 4, 2, 3.4, 3.9, 3.7, 4.8, 3.6, 
    3.9, 1.5, 0.5, 1.3, 0.2, 0.7, 1.5, 1.9, 1, 2.2, 0.9, 1.3, 1.2, 0.9, 1.2, 
    0.9, 1.5, 1.7, 1.9, 1.4, 1.7, 1.6, 3.1, 3.5, 3.4, 2.7, 0.8, 2.6, 1.1, 1, 
    1.8, 2.3, 2.1, 0.1, 1.7, 3.4, 4.3, 4.7, 4.6, 5.6, 5.2, 5.6, 7.1, 7.3, 
    8.2, 8.3, 8.4, 8.9, 7.8, 8.8, 8.7, 8.6, 8.7, 8.7, 8.6, 9.5, 9.4, 8.9, 
    8.4, 8.1, 7.7, 8, 7.5, 6.5, 5.3, 4.9, 4.1, 2.8, 1.2, 1.3, 0.3, 2.5, 5.5, 
    6, 4.8, 4.9, 5.5, 5.3, 4.9, 4.4, 4.3, 2.7, 5.3, 4.6, 6.9, 8, 7, 7.4, 7.1, 
    5.3, 5.3, 3.5, 3.4, 4.3, 4.4, 5.2, 2.7, 2.5, 1.9, 1.5, 1.1, 1.1, 1.6, 0, 
    1.4, 1.7, 1.6, 1.8, 2.5, 3.6, 4.1, 4.6, 4.6, 7.8, 7.3, 7.2, 6.7, 6.5, 
    7.6, 6.2, 6.3, 4.7, 5, 5.3, 4.7, 3.9, 3.9, 2.8, 3.5, 3.2, 2.9, 3.3, 3.8, 
    3.7, 3.2, 3.1, 3.4, 4.6, 3.8, 3.3, 3, 2.5, 2.3, 2.5, 2.7, 2.5, 2.4, 1.8, 
    1.9, 1.4, 0.6, 0.6, 0.8, 1.9, 3, 2.3, 2.9, 3.1, 5.8, 4.2, 5.6, 6.4, 2.7, 
    6.7, 4.7, 3.9, 4.9, 4.3, 4.3, 3.9, 3, 2.7, 1.1, 1, 2.6, 3.3, 3.5, 2.7, 4, 
    4, 4.1, 4.4, 4.6, 4.4, 4.2, 4.8, 3.6, 4, 3.7, 3.4, 3.3, 4.4, 5.2, 4.2, 5, 
    5.9, 5.7, 4.8, 6.3, 5.9, 7.4, 9.2, 11.1, 12.2, 13.6, 9.6, 11, 11.2, 11.4, 
    10.8, 10.4, 6, 1.8, 5.6, 5.8, 4.7, 5.1, 5.1, 5, 5.2, 5, 5.4, 6.3, 2.5, 
    9.2, 10.7, 11.9, 10.2, 10.5, 11.2, 13.9, 13.6, 14.2, 7.6, 7.4, 6.3, 5.5, 
    6.7, 3.9, 2.8, 2.9, 3.8, 5.4, 4.6, 4.6, 5.2, 5.5, 6, 4.2, 3.7, 4.2, 3.5, 
    1.6, 1.1, 1.7, 2.6, 3, 3.4, 1.7, 2.8, 2.7, 1, 2.3, 3.3, 2.3, 2.6, 4.7, 
    5.6, 4.7, 4.9, 7.6, 5.8, 4.4, 4.4, 5.9, 4.4, 4.2, 5, 5.9, 4.2, 3, 2.7, 
    1.9, 1.8, 1.9, 1.3, 2.2, 2, 1.9, 0.8, 2.6, 1, 2.1, 0.9, 0.6, 0.6, 2, 1.8, 
    0.2, 3.4, 3.6, 1, 1.6, 1.1, 1.6, 1.6, 0.2, 1.4, 1.7, 4, 1.3, 2.8, 0.6, 
    1.4, 0.6, 1.1, 2.1, 0.5, 0.5, 2.1, 5.1, 3.9, 3.4, 2.3, 1.2, 1.6, 1.8, 
    1.7, 2.2, 1.4, 1.4, 0.6, 1.4, 1.9, 1.2, 1.3, 1.5, 1.3, 2.1, 1.2, 0.4, 
    1.6, 1.4, 2, 2, 1.4, 5.5, 3.3, 2.9, 5.3, 6, 3.8, 2.7, 6.3, 8.6, 7.3, 6.1, 
    7.4, 7.8, 7.5, 9, 9, 8.3, 6.8, 4.4, 6.5, 7.9, 3, 0.9, 0.4, 0.7, 1.3, 0.9, 
    6.2, 1.4, 1.4, 3.3, 2.2, 6.8, 2.8, 2.5, 1.6, 5.5, 5.4, 4.9, 7.5, 3, 3, 
    4.9, 1.7, 9.4, 2.2, 2.4, 4.1, 5.2, 3.1, 10, 3, 4.3, 14.4, 13.9, 10.6, 
    16.5, 17.1, 16.8, 15.6, 14.5, 14.1, 14.4, 15.2, 15.1, 16.7, 14.8, 16.5, 
    16.2, 15.8, 15.5, 13.6, 12.2, 13.6, 14.4, 12.1, 13.4, 2.8, 1.9, 8.1, 
    15.7, 10.7, 11.8, 12.1, 2.7, 1, 2, 13.1, 3.3, 12.8, 11.8, 12, 12.2, 14.1, 
    15.8, 15.6, 8.8, 9.3, 11.8, 12, 3.7, 1.2, 3.2, 3.3, 3.1, 1.5, 2.1, 2.5, 
    3.9, 3.4, 4.7, 1.6, 1.6, 1.7, 3.7, 2.5, 2.2, 1.5, 3, 2.6, 1.1, 1.3, 1.9, 
    2.7, 2.3, 1.2, 1.6, 1.6, 2.2, 1.6, 2.2, 1.5, 1.9, 2.6, 0.9, 2, 2.1, 4.1, 
    1.3, 1.9, 1.1, 2.6, 5, 7.3, 2.7, 2.4, 1.2, 1.8, 1.7, 1.1, 11.3, 11.1, 
    10.7, 10.6, 10, 9.9, 9.5, 8.4, 11.1, 10.6, 10.9, 10.3, 11.6, 11.4, 11.5, 
    11, 4.8, 1.8, 1, 1.5, 3.8, 2.7, 2.5, 1.6, 1.8, 0.3, 1.6, 1.5, 1.1, 1.9, 
    5.1, 5.4, 5.6, 6.8, 5.9, 5.7, 5, 6.5, 6.5, 7.2, 7.3, 7.1, 7.4, 7.7, 2, 
    5.2, 5.5, 4.9, 1.2, 0.1, 1.4, 1.2, 1.2, 1.2, 0.9, 1.3, 0.6, 0.2, 1.4, 
    0.8, 1, 1.3, 1.3, 1.1, 1.3, 1.6, 2.7, 1.5, 3.1, 1.4, 1.3, 1.1, 4.6, 4.3, 
    2.4, 2.3, 2.2, 0.9, 12.4, 12.5, 12.2, 13, 14.4, 15.1, 9.2, 4.4, 8, 16.3, 
    15.9, 18.4, 18.5, 20.7, 21, 20.3, 19.8, 19.8, 19, 14.3, 14.1, 3.2, 5.1, 
    6.4, 6.7, 6.1, 6.9, 9.3, 9.4, 9.1, 8.7, 9.9, 9.6, 9.1, 10, 10.4, 11.3, 
    9.3, 11.6, 12.4, 12.1, 11.8, 12.1, 12.3, 11.4, 10.9, 12.1, 8.1, 8, 7.4, 
    8.1, 7.9, 8.7, 8.8, 8.7, 2, 3.1, 2.4, 3.9, 2.7, 1.9, 2.3, 2.6, 2.4, 1.8, 
    2.6, 3.1, 3.4, 3.8, 3.2, 5.8, 5.8, 5.5, 7.4, 5.8, 6.9, 6.9, 7.7, 8.5, 
    10.2, 10.5, 9.7, 10, 10.3, 11.8, 11.8, 12.1, 12.6, 10.9, 9.7, 8.3, 6.4, 
    7.4, 7.3, 5.9, 7, 5.9, 5.4, 5.4, 3.8, 3.5, 3.5, 5.7, 1.6, 1.3, 3.5, 4.1, 
    3.4, 3.4, 6.1, 3.6, 3.5, 5.2, 6.1, 5.1, 5.6, 5.5, 5.4, 3.4, 2.1, 3.4, 
    3.4, 2.9, 2.5, 1.7, 3.8, 3.3, 3.9, 3.4, 3.2, 3, 3.4, 1.1, 0.3, 0.4, 1, 
    0.4, 0.8, 1.4, 2.2, 2.2, 3.4, 1.9, 1.8, 2, 1.1, 1.2, 1.3, 2, 1.1, 0.5, 
    1.6, 1.6, 3.2, 5.3, 5.4, 5.7, 5.9, 7.2, 6, 5.9, 6.8, 6.2, 5.5, 7.2, 7.8, 
    7.3, 6.2, 3.3, 4.4, 6.7, 7.9, 5, 4.4, 4.4, 3.2, 5.5, 7.2, 8.7, 6.5, 5.5, 
    5, 4.1, 3.7, 4.4, 5.6, 6.1, 6.1, 6, 5.9, 5.7, 6.9, 5.5, 7.2, 7.2, 7.6, 
    7.7, 7.8, 7, 6.8, 6.6, 5.2, 6, 6.1, 4.7, 4.6, 4.6, 4.2, 3.4, 2.6, 2.4, 
    1.6, 2.1, 1.1, 1.8, 2.5, 4.2, 4.1, 1.2, 1.6, 0.9, 0.8, 0.6, 2, 4.4, 5.5, 
    3.5, 3.6, 2.7, 3.2, 4, 3.3, 4.2, 4, 4.8, 4.7, 6, 5.3, 5.6, 3.7, 4.2, 3.4, 
    2.8, 2.5, 2.4, 1.6, 0.7, 1.2, 0.7, 1.7, 2.2, 1.4, 1.7, 1.2, 1, 0.4, 0.8, 
    1.2, 0.5, 1.3, 2.1, 1.1, 2.4, 2.6, 2.7, 3.5, 3.5, 4.3, 4.4, 4.3, 4.1, 
    4.3, 4.2, 3.9, 3.9, 3, 3.4, 3.2, 2.1, 0.8, 0.5, 1.4, 1, 2.9, 3.3, 4.6, 
    5.3, 4.1, 3, 2.9, 4.4, 4.1, 3, 2, 2.1, 1.4, 2, 2.9, 2.4, 1.8, 1.7, 1.5, 
    2.2, 2.2, 2, 2.9, 2.2, 3.9, 3.9, 4.3, 4.5, 4.7, 4.1, 4.2, 2.9, 2.6, 3, 
    3.8, 2.9, 2.7, 5.2, 4.8, 3.3, 3.8, 4.6, 4.1, 4.1, 3.4, 4, 2.9, 3.3, 3.8, 
    3.5, 2.8, 3, 2.1, 2.5, 3.9, 3.6, 4.1, 4.1, 4.1, 4.4, 2.8, 3.9, 4.5, 6.4, 
    6.1, 5.9, 6.9, 6.5, 5.7, 4.8, 2.9, 2.2, 1.3, 1.7, 2.4, 4.4, 6, 4.7, 4.8, 
    3.8, 1.1, 0.9, 0.8, 0.8, 5.4, 2.9, 0.6, 1.9, 7.1, 4.4, 6, 5.8, 4.8, 6.8, 
    4.4, 3, 4.1, 3.2, 2.4, 1.8, 2.2, 2.5, 5.8, 2.1, 2.9, 3.7, 4.1, 4, 4.5, 
    3.7, 1.5, 1.6, 2.2, 1.3, 1.3, 2, 2, 1.4, 1.9, 2, 2.7, 2.3, 2, 1.5, 2.1, 
    3, 2.9, 1.2, 2.6, 1.9, 2.4, 2.7, 3.8, 3.5, 5.9, 4.3, 2.7, 1.3, 1.2, 2.4, 
    2.8, 4.2, 4.4, 1.9, 2.4, 1.9, 2.2, 2.5, 1.4, 0.8, 1.6, 2.3, 2.5, 1.6, 
    0.4, 0.3, 0.8, 1.3, 1.8, 0.8, 1.6, 1.4, 2.4, 1.2, 2.7, 2.7, 2.8, 2.7, 
    3.3, 3, 2.4, 3.7, 3.4, 3.5, 3.9, 2.1, 2.2, 1.7, 1.9, 1.7, 0.7, 1.1, 1.4, 
    1.2, 2.3, 4.3, 4.2, 4.8, 5.2, 5.6, 6.4, 7.1, 8.3, 8.7, 9.5, 10.8, 8.2, 
    7.6, 7.6, 7.8, 8.6, 8.2, 7.3, 6.8, 7.6, 7.9, 7.3, 7.1, 6.8, 6.7, 6.5, 
    5.8, 5.4, 5.2, 4.8, 4.7, 4.6, 4.4, 4.2, 3.6, 3, 4.6, 2.4, 1.2, 2.1, 1.7, 
    1.8, 2.1, 1.8, 1.5, 2.1, 1.7, 0.6, 0.8, 0.3, 0.7, 1, 1.1, 2, 3.1, 3.7, 
    2.1, 3.5, 3.6, 3.3, 4.8, 4.8, 4.8, 5.5, 6.7, 7.8, 6.5, 5.6, 5.8, 7.7, 
    7.4, 5.3, 7.1, 7.2, 7.9, 7.7, 7.2, 7.4, 6.1, 7.8, 6.5, 7, 7, 9, 7.4, 7.3, 
    6.5, 7, 6.3, 6.1, 4.1, 4.7, 5.5, 4.7, 5, 4.3, 3, 5.8, 4.8, 2.7, 2.5, 2.9, 
    3.6, 3.3, 4.6, 5.8, 6.2, 6, 5.8, 6.5, 6.2, 6.3, 6.7, 5.8, 4.3, 6.2, 5.7, 
    5.6, 5, 4.4, 3.5, 2, 1.5, 1.8, 0.7, 1.8, 2.4, 3.6, 4, 5.1, 5.9, 6.6, 5.6, 
    4.6, 3.6, 3.4, 3.5, 2.9, 3, 2.7, 2.7, 0.8, 1.4, 2.1, 3.4, 3.2, 3.6, 3.6, 
    3.1, 2.1, 1.4, 1, 1.3, 2.3, 3.7, 1.3, 1.7, 4.5, 2.6, 3.4, 3.5, 3.6, 2.9, 
    1, 0.7, 2.3, 3, 3.3, 5, 5.7, 6.4, 6.2, 6, 5.2, 7, 8.3, 9.8, 8.9, 8, 9.6, 
    8.4, 7.8, 6.5, 6.4, 7.1, 6.1, 7.2, 10, 7, 7.4, 4.1, 8.7, 8, 7.8, 5.6, 
    4.3, 6, 3.2, 0.8, 1.1, 1.4, 5, 5.2, 4.2, 5.2, 4, 2.8, 3.9, 4, 6.1, 5, 
    5.8, 5.8, 4.6, 4.2, 4.1, 2.8, 1.1, 0.8, 1.6, 1.3, 0.9, 2.2, 1.8, 1.8, 2, 
    1.1, 1.4, 1.6, 3.8, 1.2, 2.1, 2.7, 2.4, 4.6, 4.1, 4.1, 4.2, 4.2, 5.1, 
    5.6, 6.6, 6.5, 6.2, 7.1, 7.8, 8.6, 8.2, 8.3, 9.6, 8.9, 9.8, 9.2, 9.1, 
    8.8, 9.1, 8.6, 6.5, 3.3, 0.8, 1.4, 3.7, 4.5, 4.4, 5.6, 6.9, 6.6, 4.6, 
    5.2, 4.6, 3.4, 4.2, 3.2, 1.2, 2.1, 4.7, 4.5, 7.8, 9.6, 8.9, 7.4, 9.3, 
    9.2, 8.6, 6.4, 7.3, 7.9, 4.7, 2.6, 2.2, 0.4, 2.7, 3.4, 3.4, 1.8, 2.2, 
    2.9, 2, 0.6, 1.1, 3, 4.7, 7.1, 9.3, 8.4, 6.5, 6.6, 6.4, 5.5, 5.1, 4.3, 
    4.7, 3.4, 3.2, 1.3, 1.6, 0.6, 3.8, 2.4, 3.8, 2.9, 2.2, 0.7, 3, 10.8, 
    11.2, 8, 8.2, 7.3, 8.3, 7.7, 8, 9.4, 7.4, 6.2, 5.9, 6.6, 7.1, 6.1, 3.5, 
    2.3, 0.5, 5.3, 4.9, 4.1, 3.9, 4.9, 6.3, 9.4, 7.6, 8.5, 8.6, 10.2, 9, 
    10.7, 8.8, 9.5, 8.1, 8.8, 9.5, 9, 9.3, 9.4, 8.7, 7.1, 6.4, 4.8, 5.6, 3.3, 
    2.5, 0.3, 3.1, 5, 7.9, 5.7, 5.3, 3.9, 6.4, 9.2, 11.1, 12.2, 10.5, 10.7, 
    12.5, 13.9, 13.4, 13.2, 15.2, 15.8, 14.9, 16, 15.1, 13.6, 14.8, 17.1, 
    16.6, 15.5, 16, 15.1, 15.7, 16.3, 15.6, 15, 15.8, 15.2, 13.8, 14.6, 15.5, 
    14.7, 14.8, 12.3, 10.3, 7.9, 6.3, 7.4, 9.4, 11.5, 9.7, 7.3, 9.1, 9.3, 
    7.6, 6.6, 4.8, 3, 3.2, 3.3, 3.5, 2.9, 2.1, 4, 4.3, 3.7, 5.5, 4.7, 4.6, 
    5.7, 4, 4.3, 3.4, 4.3, 4.7, 5.2, 6.8, 6.9, 8.7, 9.7, 8.5, 10.5, 9.2, 10, 
    9.8, 12.3, 12.6, 13.7, 13.1, 14.4, 13.1, 11.7, 9.5, 11.6, 10.8, 9.3, 9, 
    8.4, 10.1, 10.7, 11.9, 9.7, 10.6, 9.8, 10.5, 10, 11.3, 9.2, 10.3, 11.2, 
    7.6, 11.2, 9.9, 10.5, 12.3, 11.2, 11.5, 12.8, 11.9, 11.3, 11, 11.5, 13, 
    12.8, 11.2, 10.1, 10.9, 12.1, 13, 13.2, 13, 13, 13.3, 11, 13.4, 14.4, 
    14.7, 14.6, 13.4, 13.5, 11.6, 10.7, 9.1, 9.3, 10.6, 9.3, 8.2, 8.1, 8.8, 
    7, 7.1, 5.4, 4.8, 2.6, 3.5, 3.8, 4.1, 4, 5, 4.6, 4.3, 4.7, 4.1, 3.8, 3.8, 
    4, 3.5, 3.2, 3.7, 4.2, 4.2, 3.5, 3.9, 4.3, 4.5, 4.2, 3.6, 5.8, 8.3, 8, 
    9.1, 9, 9.1, 10.3, 10.3, 10.5, 11.9, 12.4, 10.9, 10.2, 9.4, 8.4, 8.3, 
    7.8, 7.4, 7.3, 6.8, 5.9, 5.7, 5.9, 4, 3.9, 2.3, 3.7, 5.5, 5.8, 3.2, 5.2, 
    5.6, 6.2, 6.5, 7.2, 7.5, 5.3, 8, 7.4, 7.5, 7.3, 7.5, 8.7, 7.7, 10.3, 3.2, 
    1, 0.7, 1.9, 3, 2.3, 3.7, 0.3, 1.1, 1.4, 4.8, 4.6, 5, 6.8, 6.5, 6, 5.9, 
    5.1, 4.4, 4.1, 4.4, 6.7, 4.1, 5.1, 6.4, 5.5, 5.3, 5.3, 5, 5.1, 5.3, 5.8, 
    3.5, 4.8, 7.3, 6.2, 7.8, 6.9, 7.2, 8.8, 9.5, 9.5, 8.8, 8.6, 6.8, 7.5, 
    7.6, 8.2, 8, 6.9, 7.3, 7.9, 6.9, 6.5, 7.4, 7.4, 4.8, 5.9, 3.5, 3.8, 3.7, 
    4.6, 3.2, 2.8, 2, 1.8, 0.1, 1.3, 0.9, 1.6, 1.4, 1.8, 4.1, 5.2, 6.4, 7.5, 
    6.6, 8.2, 3.7, 7.6, 8.3, 6.9, 6.3, 6.9, 7.7, 8.7, 5.5, 5.3, 6.9, 6.8, 
    6.5, 6.6, 4.2, 5.7, 3.2, 6, 8.1, 8.6, 9.3, 8.8, 8.6, 8.6, 9.1, 8.5, 7.4, 
    7.6, 8.1, 7.2, 6, 7.4, 7.1, 7.1, 6.1, 5.6, 5.1, 5.2, 4.6, 5.9, 4.4, 3.2, 
    1.4, 0.6, 1.4, 0, 2.6, 2.7, 5.3, 5.1, 5.9, 5.8, 7.1, 7.3, 7.3, 8.9, 8.7, 
    9, 8.6, 8.9, 8.8, 8.4, 8.3, 8.5, 7.9, 7.3, 7.4, 9, 8.3, 8.9, 8.2, 6.9, 
    6.2, 7, 7.8, 8.8, 9.6, 9.8, 8.8, 9.2, 8.8, 8.8, 10.1, 10.1, 8.9, 7.3, 
    6.5, 5.3, 3.2, 1.3, 2.1, 2.3, 1.6, 4.4, 3.4, 4.5, 6.4, 6.8, 6.4, 6.1, 7, 
    6.4, 6.8, 4.7, 5.7, 8.2, 5.3, 5.8, 5, 4.6, 4.9, 1.5, 2.6, 4.5, 4, 1.4, 
    1.4, 1.2, 1.9, 0.3, 1.3, 1.1, 2.2, 0.3, 1.2, 0.8, 1.5, 1.4, 1.6, 1.2, 
    0.8, 3, 8.3, 1.5, 6.6, 5.7, 3.8, 6.1, 6.8, 5.7, 6.4, 6.5, 5.2, 7.5, 9.5, 
    7.1, 7.8, 7.1, 6.4, 5.8, 6.6, 7.2, 8.3, 6.6, 9.4, 7.2, 4.8, 6.6, 8.1, 
    7.3, 8.7, 5.9, 7.8, 2.8, 4.7, 7, 6.1, 5.1, 5.2, 1, 2.5, 6.1, 6.1, 2.8, 
    4.5, 2.2, 2.4, 1.2, 1.2, 0.5, 1.4, 0.9, 1.1, 3.1, 2.5, 2.3, 3.9, 2.3, 
    6.8, 6.3, 5.6, 1.3, 3.8, 1.7, 0.3, 1.1, 0.6, 3, 0.4, 1.7, 6.1, 11, 9.7, 
    9.4, 9.4, 10.2, 9.1, 10.4, 9.5, 10.8, 7.8, 10.1, 9.1, 7, 10, 9.4, 8.6, 9, 
    9.3, 9, 8.7, 7.9, 5.9, 4.3, 3.8, 4, 2.9, 2.2, 1, 0.1, 4.6, 4.8, 5.7, 6.5, 
    7.6, 9.3, 9.8, 8.7, 9.1, 10.6, 10.9, 10.7, 11.2, 13.9, 12.6, 10.8, 12.2, 
    12.5, 15.1, 12.8, 10.3, 11.3, 11.3, 12.2, 9.2, 9.6, 11.3, 8.1, 9.2, 8.9, 
    8.8, 7.5, 9.5, 10.7, 7.2, 5.2, 3.2, 1.7, 1.2, 1, 2.9, 2.6, 4.6, 2.7, 2.1, 
    1, 3.5, 4.2, 6.3, 7.9, 9.9, 10.7, 10.5, 11.8, 11, 11.5, 12, 10.5, 9.7, 
    8.8, 9.1, 9.2, 8.3, 8.2, 7.2, 5.7, 6.6, 5.9, 3.1, 1.5, 2, 1.1, 0.5, 1.7, 
    2.6, 2.4, 3.6, 5.4, 5.8, 6.9, _, 8.7, 8.5, 9, 8.7, 9, 9, 8.9, 9.9, 10, 
    10.8, 11.6, 10.8, 11, 11.3, 12.1, 12.7, 12.2, 12.2, 11.7, 12.5, 10.8, 
    12.2, 12.2, 12.4, 13, 12.7, 17.2, 12.4, 11.9, 9.6, 9.6, 10, 10.4, 9, 9.7, 
    9.8, 10.4, 10.7, 9.9, 10.7, 10.7, 10.6, 10.6, 12.5, 13.1, 14.6, 17.2, 
    15.6, 15.1, 12.2, 13.5, 13.7, 12.8, 14.2, 13.1, 10.1, 11.3, 7.8, 6.1, 
    3.2, 4.7, 5.4, 4.9, 5.1, 7.9, 6.7, 6.6, 5.6, 6, 5.9, 4.6, 4.7, 4.7, 5.3, 
    6.6, 6.5, 7.5, 8.2, 8.8, 8.6, 8, 8.6, 7.2, 5.7, 6.1, 3.8, 4.4, 3.5, 2.1, 
    0.8, 1.1, 1.7, 2.9, 3.7, 4.8, 5, 4.9, 5.3, 5.6, 6.1, 6.7, 7.4, 7.8, 8.3, 
    9.2, 9.2, 9.8, 9.5, 9.2, 12.1, 13.3, 15.7, 9.5, 6.1, 5.4, 4.1, 3.6, 5.8, 
    6.4, 6, 2.1, 2, 8.1, 9.2, 7.4, 5.5, 3.8, 4.4, 4.4, 1, 0.2, 4.3, 6.1, 4.8, 
    5.4, 4.2, 2.8, 2.1, 1.1, 1.2, 4.9, 5.5, 7.1, 8.1, 10, 9.8, 7.4, 7.4, 6, 
    4.5, 3.7, 2.6, 0.4, 3.6, 3.5, 4.3, 5, 6.5, 5.2, 5, 4.3, 2.5, 2.8, 2.9, 
    2.5, 1.8, 1.6, 1.2, 2.7, 4.2, 4.2, 8.8, 6.6, 7.5, 0.9, 1, 1.1, 2.4, 8.3, 
    8.2, 9.2, 9.7, 9.9, 9.2, 9.2, 8.5, 9.8, 10.1, 9.3, 8.2, 7.3, 6.7, 2.9, 
    1.3, 2, 3.4, 3.5, 3, 2.8, 3.6, 1.9, 0.9, 0.1, 1.5, 2.3, 2.5, 0.9, 0.7, 
    2.1, 3.2, 2.1, 2.4, 2.6, 0.4, 0.8, 1.3, 3.9, 4.2, 4.1, 4.4, 5, 4.9, 4.6, 
    5.2, 6.2, 6.2, 6, 5.9, 6, 6.3, 6.3, 6, 5.7, 5.5, 5, 4.7, 5.3, 5.2, 7.7, 
    7.6, 8.1, 7.7, 8, 7.9, 8.1, 8.9, 9.4, 9.8, 10, 10.3, 11.3, 11.3, 11.1, 
    12.1, 12, 11.2, 9.5, 5.1, 6.2, 4.7, 3.9, 3.7, 5.3, 5.9, 5.8, 5.8, 7, 6.1, 
    5.8, 5.2, 6, 5.2, 5.6, 5.7, 5.4, 3.9, 4.4, 3.3, 3, 2.5, 1.8, 1.7, 1, 0.2, 
    5.2, 0.2, 1.7, 1.2, 2.6, 3, 1.3, 2.4, 5.2, 7.9, 7.9, 9.2, 10.8, 10.1, 
    7.2, 9.9, 8.3, 12.7, 8.4, 13.3, 14.7, 12.9, 16, 15.9, 15.7, 16.7, 17.6, 
    17.5, 16, 16, 16.4, 15.9, 18.6, 19.2, 22.5, 23.3, 20.8, 17.2, 16.1, 13.6, 
    12.9, 10, 9.9, 9.4, 9.5, 9.2, 8.9, 9.5, 9.3, 8.2, 8.5, 8.5, 8.4, 9.2, 
    8.8, 8.8, 9.3, 10.6, 10.9, 9.8, 11.4, 10.1, 8.6, 9.1, 10.6, 12.1, 12.1, 
    12.6, 12.3, 13.5, 13.9, 13.6, 13.6, 13.5, 13.7, 12.9, 11.4, 13.4, 15.2, 
    14.4, 12.5, 12.4, 12.6, 13, 13, 13.2, 13.9, 14.5, 13, 13.2, 13.2, 12.9, 
    13.2, 14, 10.6, 10.7, 10, 8.1, 10.2, 10.4, 10.9, 11.7, 10.9, 10.5, 9.8, 
    8.4, 5.3, 7.5, 9.3, 10.2, 10.4, 10.4, 11.3, 14.3, 12.3, 11.5, 12.4, 12.2, 
    12, 11.1, 11.2, 11, 10.2, 10, 10, 9.8, 9.8, 9.6, 9.5, 9.7, 8.9, 8.5, 7, 
    6.6, 3.2, 5.9, 6, 7.1, 7.6, 8.3, 10.1, 11, 11.9, 11.1, 10.4, 9.7, 9.9, 
    9.3, 9, 8.2, 8.9, 8.1, 8, 10.4, 9.3, 9.2, 9.6, 10.1, 10.3, 10.3, 10.1, 
    10, 11.7, 11.7, 10.3, 8.9, 9.2, 7.7, 4.2, 0.2, 2.6, 4.7, 7.3, 5.9, 6.2, 
    10.7, 12.3, 13.3, 12.8, 12.6, 12.3, 13.2, 12.1, 9.2, 8.6, 10, 8, 5.6, 
    4.5, 3.4, 2.3, 4.2, 4.8, 5.9, 7.8, 8.8, 8.9, 9.6, 10.4, 10.1, 9.9, 10.9, 
    10.7, 11.7, 10.8, 11.9, 9, 10.9, 8.4, 6.6, 6.9, 4.1, 10.1, 6.3, 2.2, 0.7, 
    0.5, 0.9, 6, 9.4, 9.1, 11.6, 15.4, 18.3, 17.6, 16.7, 17.7, 16, 17.4, 
    16.3, 15.2, 16.6, 16.2, 14.7, 14.1, 11.2, 9.9, 11.2, 9.8, 7.7, 6.3, 2.5, 
    4, 3, 6.7, 7.6, 5.2, 4.6, 7.4, 7.3, 6.5, 5.9, 5.1, 5.1, 3.4, 2.9, 2.1, 
    0.8, 3.6, 5.5, 7.6, 7.9, 9.7, 11.8, 12, 10.9, 10.3, 9.8, 9.9, 8.8, 8.1, 
    8.8, 8.3, 9, 7.9, 7.1, 7.2, 5.6, 5.6, 6, 4.9, 3, 2.9, 3.6, 2.8, 3.2, 2.3, 
    1.8, 1.4, 1.3, 4.6, 9.1, 7.6, 9, 6.2, 8.5, 11, 9.3, 8.2, 7.8, 7.4, 6.6, 
    5.4, 2.3, 1.3, 2.5, 4.2, 1, 3.9, 7.2, 8.3, 7.7, 7.9, 5.7, 4.4, 1.9, 0.9, 
    1.1, 1.8, 2.5, 5, 4.5, 4.1, 2.9, 3.2, 4.1, 4, 6.3, 5.8, 5.5, 6.1, 6, 6.6, 
    6.1, 6.1, 6.2, 5.5, 5.7, 5.5, 5.1, 5, 4.6, 4.6, 4.6, 3.9, 3.2, 2.7, 2.8, 
    2.6, 1.6, 0.7, 0.8, 2.3, 2.5, 2.4, 2, 1.6, 3.3, 4.7, 3.7, 3.5, 4.7, 4.8, 
    4.9, 4.4, 3.5, 2, 2.1, 2.6, 2.8, 3.3, 3, 2.9, 5.3, 5.2, 5.4, 6.3, 6.4, 
    7.7, 8.4, 9.1, 10, 10.8, 10.1, 10.4, 9.2, 7.6, 4.7, 3.8, 3.9, 2.6, 2.3, 
    2.1, 1.9, 5, 4.8, 4.4, 2.6, 0.8, 5.6, 2.9, 4.9, 2.1, 5.5, 5.8, 4, 3.2, 
    3.5, 3, 4.1, 8.3, 14.6, 16.2, 15.8, 16.5, 18.9, 17.4, 18.9, 18.6, 18.3, 
    19.3, 19.6, 18.3, 18.5, 19.2, 20.3, 19, 17.5, 16.9, 17.6, 17.7, 19, 18.8, 
    18.6, 16, 12.5, 10.2, 10.7, 9.1, 7.5, 5.6, 3.2, 3.8, 1.7, 1.2, 6.6, 5.7, 
    5.4, 6.2, 5.3, 5.8, 5.5, 4.8, 3.7, 3.1, 3.9, 4.2, 4.7, 5.5, 6.4, 6.8, 
    7.5, 8.2, 7.7, 5.6, 5.3, 5.3, 4.8, 5.1, 4.8, 3.7, 3.5, 1.1, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.7, 2.9, 4, 6, 6.4, 5.9, 6.4, 7.5, 7.7, 6.9, 5.3, 4.9, 4.1, 
    3.2, 2.9, 3.2, 1.4, 4, 3.6, 5.8, 6.3, 5, 6.3, 4.7, 5.6, 6.2, 6, 6.1, 6.5, 
    4.7, 3.4, 4.2, 3.9, 4.4, 2.2, 2.5, 2.6, 2.8, 2.1, 2.7, 2.2, 2.4, 2.1, 2, 
    2.7, 2.3, 2, 1.7, 5.6, 3.7, 4.9, 4.6, 7.3, 9.2, 11.1, 12.4, 12.9, 13.5, 
    4.1, 5.8, 6.5, 6.8, 6.6, 6.9, 8.6, 8.4, 4.6, 4.3, 4, 2.8, 1.9, 6.7, 6, 
    5.8, 2.1, 6.1, 6.5, 7, 5.5, 4.2, 6, 4.6, 5.2, 6.8, 7.9, 8, 10.5, 10.7, 
    11.1, 11.4, 11.4, 10.9, 11.1, 10.9, 10.1, 9.4, 8.2, 6.7, 5.7, 4.8, 4.2, 
    3, 1.6, 2.6, 3.9, 4.3, 5.3, 6.1, 6.1, 7.4, 9, 8, 8.4, 9.3, 9.6, 9.9, 
    10.5, 10.6, 10, 9.8, 9.3, 9, 9.3, 7.2, 5.1, 3.7, 2.8, 2.9, 0.9, 1, 0.7, 
    2.4, 1.5, 3.7, 3, 2.1, 2.9, 3.4, 4, 3.7, 4.6, 4.4, 3, 5.2, 3.2, 1.9, 1.3, 
    0.6, 2.1, 2.8, 3.4, 3.6, 4.4, 5.5, 5.7, 6.2, 3.9, 3.6, 3.1, 3.4, 3.7, 
    7.4, 7, 8.1, 9.1, 8.8, 8.4, 9.1, 10.2, 10.7, 11.2, 11.7, 12.5, 11.6, 
    12.3, 12.6, 13, 14.5, 13.2, 13.8, 17.3, 16.5, 14.9, 14.6, 14, 11.4, 10, 
    9.2, 5.3, 4.8, 6.4, 7, 5.6, 6.9, 6.9, 8.4, 8.4, 7.7, 7.9, 8.1, 8.4, 8.4, 
    8.1, 8.6, 9.2, 8.9, 9.3, 8.1, 8, 9.1, 10, 10.5, 10.7, 8.1, 10.5, 10.6, 
    10.6, 11.2, 10, 9.1, 6.4, 7.7, 7, 8.3, 8.6, 8.8, 9.4, 9.1, 9.3, 10, 12.6, 
    11.7, 9.6, 11.2, 12.5, 11.6, 9.4, 10.3, 9.1, 10.3, 9.7, 5.8, 8.3, 8, 9.3, 
    9.2, 10.4, 14.5, 17.2, 15.5, 13.6, 12.2, 12, 11.7, 13, 13, 8.8, 10.3, 
    10.7, 10, 6.2, 7.9, 6.7, 7.4, 8.1, 5.9, 4.9, 6.5, 8.3, 5.9, 2.6, 2, 1.5, 
    1.9, 2.4, 3, 1, 4.3, 5.4, 2.5, 0.5, 2.3, 4.1, 4.4, 4.3, 5, 4.5, 3.2, 1, 
    0, 2.5, 3.2, 2.5, 3.2, 4.2, 2.4, 2.7, 3.1, 2.4, 2.2, 2.6, 0.6, 1, 4.1, 
    2.2, 2, 4.7, 2.7, 4, 5.4, 4.8, 5.1, 4.1, 1.8, 0.8, 1.2, 1.1, 0.7, 5.2, 
    4.6, 4.2, 5.8, 4.2, 5.2, 4.5, 3.3, 5.1, 3.6, 3.1, 2.4, 2.7, 2.4, 2.1, 
    2.4, 2.7, 2.7, 3, 4.6, 4.9, 5, 6, 5, 5.5, 5.3, 5.5, 5.3, 5.3, 5.3, 5.7, 
    5.5, 6.1, 6.7, 6.9, 5.7, 4.7, 6.5, 7.8, 6.6, 7.8, 8.1, 7.5, 7.4, 7.7, 
    7.7, 6, 7.8, 4.8, 7.2, 7.5, 6.3, 7.2, 8.3, 8.1, 6.9, 8.1, 8.6, 7.3, 7, 
    7.8, 6.8, 5.9, 6, 6.6, 5.3, 4.8, 6.3, 5.6, 6.2, 6.8, 6.9, 7.3, 7.5, 7.2, 
    7.4, 6.4, 6.7, 6.5, 6, 6.5, 6.8, 6.7, 6.2, 6.9, 6.7, 6.8, 7.3, 9.2, 7.7, 
    6.4, 7.3, 7.4, 6.5, 6.4, 6.1, 7, 4.9, 3.9, 4.4, 1.4, 6.4, 8.5, 7.5, 8, 
    7.6, 6.7, 6.3, 5.9, 5.1, 5.1, 4.7, 4.3, 4.9, 3.4, 2.2, 2.8, 3.1, 4, 4.1, 
    2.2, 3.1, 5.3, 4.9, 6.6, 7.6, 8.6, 8.2, 8.8, 6.9, 10.2, 11.2, 9.7, 8.6, 
    7.9, 7.5, 7.4, 6.9, 7.5, 7.8, 7.8, 7.8, 7.7, 7.4, 8.1, 7.1, 6, 6.8, 11.1, 
    6.6, 6.9, 9.1, 8, 7.6, 9.8, 9.4, 10.6, 10.1, 10.1, 11.2, 11.5, 13.1, 
    14.3, 13, 12.4, 12.7, 11.8, 12.3, 12.4, 14.1, 13.1, 13.7, 12.1, 10.4, 
    9.9, 12.9, 7.9, 7.5, 13.1, 10.5, 11.1, 18.6, 14.3, 20.5, 21.2, 22, 19.5, 
    18.7, 15.5, 17.1, 18.7, 18.1, 16, 16.4, 17.4, 17.4, 17.1, 17, 17.3, 17.1, 
    14.9, 16, 16.6, 15.5, 16.8, 14.3, 14.5, 13.7, 14.7, 14.6, 10.8, 12.3, 
    9.6, 8.4, 8, 8.3, 8.1, 7.8, 7.8, 6.8, 6.4, 5.3, 5.2, 3.6, 1, 0.6, 0.5, 
    0.1, 3.7, 2.5, 5.3, 3.3, 1.4, 0.8, 0.8, 1, 0.4, 0.6, 0.8, 1, 2.6, 2.5, 3, 
    2.5, 3, 3, 2.7, 4.9, 6.8, 7.6, 7.9, 8, 8.1, 7.8, 7.1, 7.3, 7.7, 7.8, 6.7, 
    4.4, 4.8, 5, 5.8, 5.7, 5.8, 5.7, 8.1, 9.3, 11.1, 11.6, 10.8, 11, 11.4, 
    11.4, 11.5, 11, 11.7, 12.1, 11.4, 12.4, 11.7, 11, 11, 11.1, 11.1, 10.6, 
    11, 10, 10, 9.2, 9.3, 9.6, 9, 8.5, 8.6, 6.7, 7.6, 7.1, 6.9, 7, 6.7, 5.2, 
    7.6, 7.9, 7.5, 7.6, 7.6, 6.8, 8.4, 6.7, 6.1, 7, 6.5, 7.3, 6.9, 5.7, 6.8, 
    7.4, 10.2, 12.4, 12.8, 14.3, 13.3, 12.1, 12, 13, 16.1, 16.3, 15.4, 16.5, 
    16.7, 18.5, 19.9, 19.6, 19.1, 18, 16.3, 12.5, 13.2, 14.7, 15, 13.9, 12.9, 
    11.4, 14.1, 13.4, 14, 14.2, 13.9, 13.6, 13.4, 14.7, 12.7, 11.8, 10.6, 11, 
    9.9, 8.6, 9.2, 8.8, 9.2, 9, 9.4, 9.3, 9.9, 11.3, 12.2, 13.7, 15.2, 15.6, 
    15.4, 16.3, 16.9, 16.3, 16.3, 15.4, 15.2, 15.5, 15.6, 16.2, 16.8, 17.6, 
    18.4, 17.9, 18, 17.5, 16.2, 15.4, 12.9, 12.3, 13, 12.3, 12.6, 12.2, 9.2, 
    11.6, 8.5, 9.8, 11.1, 9.5, 9.4, 10.1, 10.6, 9.4, 9.7, 9.8, 10, 10.3, 9.3, 
    7.8, 8.3, 7.9, 7.4, 6.4, 8.8, 7.3, 7.1, 7.3, 7, 7.4, 6.2, 7.9, 5.9, 7.1, 
    7, 7, 5.9, 8.2, 7, 6.5, 7.6, 10.5, 10, 6.9, 6.7, 6.6, 7.4, 7, 7.7, 7.5, 
    7.3, 8.5, 9.6, 9.1, 7.4, 5.8, 4.2, 4.3, 6.4, 5.8, 2, 8.5, 8.6, 8.2, 9.3, 
    6.1, 9.4, 8.7, 8.9, 9.2, 2.4, 8.9, 10, 8.8, 7.7, 5.7, 7.7, 6.3, 6.1, 6.1, 
    8.6, 9.5, 7, 5.4, 6.4, 8.2, 7.7, 7.6, 6.9, 6.2, 7.4, 6.6, 5.3, 3.6, 3.3, 
    2.1, 1.5, 3.7, 4.4, 5, 6.4, 4.6, 4.1, 2.9, 2.9, 1.5, 2.2, 1.2, 2, 2.3, 
    3.1, 4.2, 3.3, 4, 3.8, 4.8, 4.4, 4, 3.1, 2.6, 2.2, 2.2, 1.9, 3.7, 4.3, 
    1.3, 2.9, 2.9, 3.9, 3.7, 3.7, 5.1, 4, 4.8, 5.6, 5.1, 5.4, 6.8, 6.8, 5.9, 
    7.1, 7.5, 8.6, 6.4, 9.5, 8.7, 6.8, 3.9, 2.5, 5.4, 4.1, 6.7, 7.7, 6.4, 
    6.5, 6, 5.1, 3.8, 3.4, 2, 1, 0.7, 1.2, 2.4, 2.6, 1.3, 7.5, 5.9, 5.4, 8.7, 
    4.9, 5.7, 5.2, 3.6, 6.6, 3.6, 1.8, 2.3, 2, 1.9, 1.8, 1.4, 1.9, 1.7, 0.8, 
    6.4, 7.2, 6.4, 5, 5.8, 6.3, 8.1, 7.9, 5.9, 7.4, 6.9, 6.6, 7.1, 6.9, 7.7, 
    7.4, 5.8, 7.5, 10.9, 11.2, 9.7, 9.1, 8.7, 8.6, 6.6, 7.9, 8.5, 8.6, 9.1, 
    7.5, 9.5, 6.7, 7.5, 7.6, 10.2, 11.1, 10.5, 7.8, 7.8, 5.5, 7, 9.4, 10, 
    10.7, 9.3, 12, 10.1, 10.7, 7.4, 12.5, 13.7, 12.1, 12.9, 11.8, 10.2, 9.7, 
    8.7, 9.2, 9.4, 10.7, 10.6, 7.4, 6.8, 6.8, 6.6, 6.9, 8.4, 5.7, 5.6, 6.3, 
    7.6, 6.9, 5.6, 5.7, 5.2, 4.7, 6.3, 6, 4.1, 4.9, 3.7, 3.7, 4, 4.1, 6, 7.6, 
    5.6, 7.4, 8.6, 6.5, 5.8, 3.6, 8.6, 9.2, 9, 9.7, 10.3, 10.2, 10.9, 9.9, 
    10.2, 7.8, 7, 9.3, 9.3, 11.5, 11.4, 11.2, 9.5, 9.6, 9.4, 11.8, 10.7, 10, 
    8.5, 9.2, 10.2, 10.6, 7.5, 10.1, 10.4, 9.4, 10.5, 10, 11.9, 10.2, 10.3, 
    10.3, 9.8, 6.3, 6.8, 9.5, 8.4, 11, 9, 10.3, 10.8, 10.4, 8.6, 9.9, 8.3, 
    10.5, 10.3, 9.5, 9, 8.9, 9.5, 8.1, 7.6, 9.4, 5.3, 4.7, 5.3, 6, 5.7, 4.9, 
    4.3, 3.6, 2.7, 2.2, 2.4, 1.6, 2.1, 3, 1.3, 0.6, 1, 2.2, 3.3, 4.4, 5.4, 
    4.9, 4, 3.9, 4.6, 5.1, 6.2, 5.5, 6.5, 7.2, 6.2, 6.4, 8.4, 9, 11, 7.8, 
    6.1, 5.8, 8.5, 7.9, 7.9, 8.2, 10, 8.6, 9.6, 8.2, 7.9, 7.4, 7.3, 7.9, 7.3, 
    6.7, 7.8, 6.8, 4.6, 6.4, 5.9, 6.7, 5.2, 8.1, 10.4, 9.8, 9, 9.2, 8.8, 8.9, 
    8.3, 8.4, 8.5, 7.7, 8.5, 10.4, 11.2, 9, 12.6, 12.5, 10.4, 10.2, 10, 12, 
    12, 11.9, 11.9, 12.3, 11.8, 13.6, 16.3, 14.7, 15.9, 17.1, 16.1, 16.7, 
    17.7, 17.6, 17.6, 18, 13.7, 10.4, 11.2, 11, 10.2, 7.7, 10.2, 10, 9.5, 
    12.3, 15.2, 11.7, 11.4, 11.8, 11.2, 10.7, 10.4, 9.5, 9.1, 9.5, 9.1, 8.6, 
    8.3, 8.4, 8.6, 8.2, 9.5, 9, 8.9, 9.2, 9, 9, 8.3, 7.9, 7.8, 7.5, 7.1, 6.7, 
    7.8, 7.8, 7.5, 7.4, 7.6, 7.5, 7.6, 8, 8.3, 8.6, 9.5, 10.1, 11.3, 11.6, 
    11.9, 12.1, 12.1, 12, 11.8, 11.8, 12.1, 12.4, 12.5, 11.6, 10.3, 9.8, 
    10.7, 12.5, 10.3, 2.4, 8.8, 12.9, 12.6, 10, 7.8, 5.7, 10.4, 8.6, 6.1, 
    3.8, 6.7, 10, 10.3, 10.4, 9.6, 10.5, 11.9, 12, 11.8, 12.2, 12.4, 12, 12, 
    12.4, 12.9, 13.8, 13.5, 13.6, 13.7, 13.6, 12, 11.6, 11.4, 11, 10.7, 10.6, 
    10.5, 10.3, 10.1, 10.2, 10.1, 10.3, 10.1, 9.8, 8.8, 7.7, 8.1, 8, 8.5, 9, 
    8, 8, 8.5, 8.8, 8.9, 9.1, 9.2, 9.1, 9, 9, 8.7, 8.5, 8.3, 7.8, 7.6, 7.7, 
    8, 9.2, 10.5, 11.2, 11.7, 12.2, 12.6, 12.6, 12.5, 12, 12, 12.2, 13, 12.8, 
    13, 12.7, 11.9, 11.3, 11.3, 11.6, 11.6, 11.5, 11, 10.2, 9.7, 9.4, 9, 8.7, 
    8.5, 8.3, 8.1, 7.6, 7.5, 7.7, 7.7, 7.8, 8.4, 7.8, 7.1, 6.6, 6.4, 6.2, _, 
    6, 5.5, 4.9, 4.3, 4.8, 4, 4, 3.9, 3.9, 3.8, 3.6, 3.7, 3.9, 4.2, 4.5, 4.7, 
    4.7, 3.9, 4, 4.3, 4.7, 4.9, 5.4, 5.7, 6, 6.5, 7.1, 7.1, 6.9, 8.7, 9, 9.3, 
    9.4, 9.3, 9.5, 10, 10.4, 9.9, 9.7, 10.2, 11.3, 11.7, 12, 12.4, 12.2, 
    11.9, 11.6, 11.4, 11.9, 10.1, 10.1, 8.6, 9.5, 10.6, 10.9, 10.5, 10.1, 
    10.4, 10.2, 10.3, 9.4, 8.2, 7.8, 6.5, 7.2, 6.9, 6.1, 3.7, 1.8, 2.7, 5.8, 
    9.8, 8.9, 10.3, 8.6, 8.3, 7.5, 6.5, 6.1, 3.6, 0.1, 2.2, 4.1, 2.9, 1.8, 
    2.7, 2, 6.2, 12.6, 12.3, 13.2, 12.9, 12.4, 11.9, 11.3, 7.8, 11.4, 10.8, 
    10, 10.3, 10, 3.4, 10.3, 9.7, 9, 9, 9.8, 10.2, 10.6, 9.8, 10.4, 9.9, 12, 
    9.8, 6.8, 8.6, 8, 7.6, 9.2, 9.3, 8.6, 5.8, 13.1, 11.4, 12, 12.2, 12.7, 
    13.8, 14.7, 14.4, 14.8, 10.5, 6.6, 7.6, 9.9, 7.7, 2, 1.8, 1.2, 1, 1, 0.9, 
    0.8, 0.8, 12.4, 0.6, 0.5, 0.6, 0.4, 0.4, 0.4, 0.4, 0.3, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9, 1, 1.1, 1.2, 1.3, 1.3, 1.3, 
    1.2, 1.1, 0.7, 0.7, 0.4, 0.6, 0.8, 0.8, 0.8, 0.7, 0.6, 0.4, 0.3, 0.4, 
    0.3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4, 15.4, 17.2, 20.6, 
    22.4, 22, 17.2, 14.4, 12.6, 13, 11.4, 11.8, 8.9, 10, 11, 13.7, 12.5, 
    11.4, 13.1, 15, 13.4, 10.1, 8.7, 9.2, 8.5, 8.7, 9.2, 7.4, 8, 10, 11, 
    12.9, 11.9, 11.7, 11.7, 9.7, 7.4, 8.8, 10.5, 9.3, 7.9, 11.4, 10.7, 10.7, 
    10.5, 9.7, 9.5, 9.4, 10.9, 12.3, 11.8, 12.9, 13.5, 13.2, 13.5, 12.5, 12, 
    12.9, 12.3, 11.4, 9.7, 9.7, 7.4, 8.5, 10.4, 11.1, 8.6, 7.4, 7.3, 8.3, 
    7.6, 6.7, 6.6, 9.1, 2.8, 1.8, 2.1, 1.5, 9.6, 7.6, 7.6, 7.2, 7.7, 5.6, 
    6.9, 6.7, 7, 7.3, 6.9, 6.2, 8, 8, 9.6, 9, 9.5, 8.7, 8.2, 6.1, 6.9, 9.8, 
    10, 11.6, 8.8, 8.3, 7.8, 6.4, 5.4, 6.7, 8.1, 8.6, 7.9, 12.1, 11.8, 13, 
    14.1, 16.9, 15.1, 14, 14.6, 14.9, 12.6, 14.8, 17.8, 17.7, 14, 11.7, 10, 
    10, 11.3, 10.4, 11.3, 14.5, 15.9, 15.9, 17.9, 16.7, 17.8, 20, 19, 17, 13, 
    8.7, 9.9, 9.1, 8.1, 6.6, 5.1, 7.1, 8.7, 7, 4.5, 5.3, 4.6, 4.3, 1.9, 1.6, 
    2.2, 2.2, 1.4, 3.8, 4, 9.9, 9.7, 8.7, 9.4, 6.2, 7.1, 8.3, 4.8, 4.5, 4.3, 
    6.1, 5.6, 4.5, 7.2, 8.2, 10.9, 9.9, 10.6, 11.4, 13.4, 14.5, 13.7, 14.9, 
    15.7, 15.3, 17.1, 16.7, 16.3, 18.2, 15.7, 18, 20.5, 20.1, 18.1, 15.8, 
    14.6, 14, 14, 16, 14, 10.8, 10.2, 11.4, 10.5, 11.1, 7.6, 9.4, 8.5, 8.2, 
    7.5, 8.4, 9.7, 7.4, 7.1, 7.6, 9.4, 12.3, 10.2, 7.4, 9.2, 7.8, 7.5, 11.5, 
    8.4, 8.3, 7.6, 9.1, 10.9, 9.2, 8, 9.1, 9.5, 10, 11, 9.3, 8.1, 9.8, 8.8, 
    8.7, 9.4, 8.7, 8.3, 9, 8.1, 6.1, 7.9, 8.5, 7.5, 6.6, 7.6, 9, 5.3, 5.4, 
    6.9, 5.2, 5.1, 2.6, 4.7, 6.8, 5.3, 6.3, 5.7, 4.9, 6.7, 6.9, 5.1, 5.1, 
    5.9, 5.1, 8.1, 7.3, 7.8, 7.9, 7, 6.3, 7.5, 6.2, 7.1, 7.3, 7, 7.9, 9, 8, 
    10.7, 11.6, 10.9, 9.9, 7.1, 8, 9, 10.8, 9.2, 10.1, 9.5, 9.2, 9.1, 7.1, 
    8.7, 9.4, 8.4, 8.8, 9.7, 9.3, 9.9, 8.7, 9.4, 9.1, 9, 9, 9.1, 9, 8.4, 8.2, 
    8.2, 8.1, 7.7, 7.4, 8.1, 8.7, 7.9, 8.2, 8.9, 9.4, 9.9, 10.1, 10.2, 11, 
    12, 12.1, 11.9, 11.5, 11.4, 12, 13.2, 12, 11.3, 9.1, 8.9, 7.9, 8, 6.7, 
    8.4, 4.9, 7.9, 7.2, 7.1, 6.9, 9.1, 6.8, 7.9, 5.8, 6, 5.5, 3.4, 3.5, 8.9, 
    8.6, 8.7, 10.4, 10.5, 11.5, 10.6, 8.4, 13.2, 9.4, 13.1, 14.4, 14.9, 14.9, 
    15.2, 13.8, 11.5, 9.6, 9, 7.9, 6.1, 8.4, 4.9, 3.3, 6.1, 8.3, 5.9, 8.1, 
    7.6, 9.6, 11.5, 13.2, 13.8, 13.2, 12, 9.3, 10.2, 9.4, 8.5, 9.3, 8.2, 8.1, 
    6.2, 5.4, 6.8, 6.9, 5.9, 6.3, 8.2, 8.5, 8.6, 8.4, 8.2, 8.5, 9.3, 10.8, 
    10.1, 10, 10.2, 8.3, 10.1, 9.4, 8.9, 9.2, 8.8, 8.4, 9.8, 7, 8.9, 9.6, 
    8.2, 8.5, 7, 6.2, 3.5, 8.2, 8.5, 8.6, 6.4, 4.7, 6.1, 7.4, 8.1, 5, 4.5, 
    4.8, 4.9, 4, 3.8, 6.2, 6.8, 6.4, 5.9, 4.7, 4.9, 4.4, 8.3, 6.3, 7.5, 7.6, 
    7, 8.2, 9.3, 9.2, 9, 11.2, 9.7, 10.7, 10.6, 13.1, 13.1, 12.8, 16.2, 16.7, 
    17.4, 15.9, 16.9, 19.8, 19.7, 17.3, 16, 17.3, 22.6, 22.9, 21.2, 21.2, 21, 
    17.2, 17.1, 15.8, 16.7, 14.5, 14.6, 14.6, 13.8, 13.3, 12, 11.3, 10.2, 
    9.4, 8.5, 6.3, 7.2, 3.7, 7.6, 5.9, 4.9, 3.8, 2.1, 1.3, 2.8, 2.1, 3.6, 
    3.5, 4.8, 5.2, 4.8, 4.8, 5.3, 5.8, 5.1, 4.7, 5.3, 5.3, 5.8, 5.4, 5.4, 
    8.2, 6.4, 7.8, 6.4, 6.7, 7.4, 8.7, 6.9, 7.7, 8.4, 5.1, 8.1, 7.9, 7.7, 
    6.4, 6.2, 6.3, 5.9, 5.5, 5, 4.2, 1.2, 1.9, 0.6, 3.2, 3.6, 5.1, 6.3, 5.1, 
    10.3, 6.9, 8.8, 9.3, 9.3, 7.1, 6.6, 5, 5.6, 5.8, 4.1, 4.8, 3.8, 3.4, 3.1, 
    2.7, 4.5, 3.5, 3.9, 3.7, 5.8, 7.5, 8.9, 10.3, 10.5, 9.5, 11.7, 12.3, 
    14.2, 14.7, 13.8, 13.2, 17.5, 14.6, 15.7, 13.7, 8.8, 15.8, 14.7, 15.8, 
    12.9, 12.5, 12, 11, 9.7, 9.4, 10.1, 7.7, 8.8, 7.2, 5.2, 6, 5.8, 7.4, 6.2, 
    6, 6.1, 5.6, 6.4, 5.8, 4.9, 6.4, 7.9, 11.6, 9.7, 8.9, 6.8, 5.9, 2.7, 4.9, 
    4.9, 4.9, 7.9, 11, 13.5, 15.2, 14.8, 15.1, 16.6, 15.6, 15.2, 16.1, 17.2, 
    18.2, 19.1, 19.3, 17.9, 15.3, 14.1, 12.1, 10, 6.4, 5.2, 8.4, 4.2, 8, 10, 
    12.2, 10.5, 12.2, 13.3, 13.1, 12.5, 11.3, 11.4, 13.4, 9.4, 14.1, 10.6, 
    10.6, 10.1, 13.2, 15.7, 14.2, 13.2, 13.4, 15.5, 14.7, 15.7, 14.2, 14.2, 
    14.2, 17.1, 16.3, 15.9, 16.5, 16.8, 16.6, 15.9, 15.1, 13.5, 13.2, 13.3, 
    12, 13.1, 11.8, 13.9, 14.1, 13.5, 13, 9.4, 7.5, 10.2, 8, 7.6, 8.2, 7.2, 
    2.6, 6.8, 5.6, 9.3, 10.2, 7.8, 7.4, 11.7, 12.4, 11.1, 10.1, 9.1, 7.4, 
    8.3, 6, 7.1, 8.9, 8.8, 10.7, 10.5, 10.8, 11.6, 10.8, 13.1, 12.8, 13.3, 
    14.9, 14.4, 14.6, 13.9, 10.1, 11.1, 10.6, 8.4, 8.7, 8, 8.1, 7.8, 8.7, 
    8.5, 10.6, 11.4, 11.7, 13.6, 11.7, 7.5, 9.9, 8, 9.1, 8.3, 8.6, 9.7, 10.3, 
    9.5, 8.9, 9.6, 8.8, 9, 6.7, 8.6, 10.1, 10.3, 9.5, 9.1, 7.1, 5.5, 2.4, 
    4.8, 12.7, 11.5, 9.9, 8.4, 10.1, 8.3, 5.9, 5.2, 9.1, 9.8, 8.2, 7.9, 6.5, 
    6, 5.5, 5.5, 5.6, 4.8, 4.9, 4.9, 5.1, 6.2, 6.4, 6.5, 8.2, 7.7, 7.4, 9.1, 
    9.2, 8.5, 9.1, 10.6, 10.6, 10.6, 11.2, 10.4, 9.6, 11.1, 9.6, 10.6, 10.6, 
    11.4, 10.3, 9.8, 10.2, 11, 12, 12.1, 11.8, 11.7, 12.6, 12.8, 12.2, 12.5, 
    12.8, 12, 12.3, 12.9, 12.3, 11.3, 11, 11.6, 12.1, 13.4, 13.8, 18, 14.9, 
    16.4, 15.4, 15, 17.1, 16.6, 15.3, 13.6, 17.6, 15.7, 13.9, 13.4, 11, 11.6, 
    10.1, 11.8, 11.4, 10.6, 11.2, 12, 11.9, 11.6, 12.6, 12.9, 12.2, 12.9, 
    13.4, 13.9, 14.5, 14.4, 14.6, 14, 14, 14.7, 13.9, 15.1, 16.2, 16, 16.8, 
    17.3, 16.8, 15.5, 17.1, 17.1, 15.2, 15.8, 15.9, 14.9, 14.6, 14.5, 15.2, 
    16.5, 16.2, 16, 16.8, 17.6, 17, 16, 14.5, 15.4, 14.4, 14.1, 14.3, 13.6, 
    14.6, 15.1, 15.7, 16, 14.5, 13.9, 13.7, 11.8, 10.9, 11.1, 13.3, 12.4, 
    11.6, 12.6, 12.8, 10.6, 8.5, 7.5, 7.9, 11.7, 8.1, 9.5, 10.7, 10.7, 12.2, 
    13.1, 12.8, 13.1, 12.6, 14.4, 13.2, 13, 14.2, 13.4, 14.6, 13.2, 13.5, 
    11.4, 12.2, 10.8, 11, 10.1, 10, 9.7, 11.2, 9.3, 9.8, 10.5, 11.2, 11, 9.6, 
    9.9, 10.3, 9.7, 10, 11.9, 11.6, 11.6, 11.9, 11.3, 11.3, 8.7, 10, 11.1, 
    10.8, 11.3, 12.4, 12.2, 12.3, 12.8, 13.1, 13.4, 9.3, 5.5, 9.5, 7.9, 7, 
    4.3, 3.2, 16.4, 14.2, 16, 19.2, 20.8, 14.7, 11.2, 7.4, 8.6, 17.2, 12.6, 
    14.5, 15.5, 14.6, 18.4, 18.9, 18.1, 17.6, 16.9, 16.7, 17.4, 18.3, 17.9, 
    19, 19.6, 21, 21, 20.4, 20.2, 19.3, 18.3, 17, 17.4, 17.4, 16.7, 15.9, 
    15.9, 16.7, 14.4, 11, 12, 10.9, 10, 7.1, 7.3, 4.5, 1.8, 1.1, 1.8, 3, 4.7, 
    6.2, 6.9, 6.1, 7.4, 7.9, 9, 10.1, 9.1, 8.7, 8.6, 8.8, 9, 9, 9, 9.6, 9.6, 
    11, 11.1, 12.7, 13.6, 13.7, 14, 13.1, 13.4, 12.7, 12.8, 12.6, 13.1, 13.6, 
    12.4, 12.1, 12.5, 12.7, 12.9, 12.4, 12.5, 12.3, 12.5, 12.8, 12.7, 12.2, 
    13.3, 14.2, 14.1, 14.1, 14.3, 14.9, 13.9, 13.8, 14.3, 13.4, 12, 8.5, 6, 
    5.1, 3.3, 2.4, 1.5, 1.5, 7.4, 8.8, 12.5, 11.6, 10.9, 7.5, 7, 7.3, 4.3, 
    3.4, 5.6, 5.4, 5.4, 5.7, 7.8, 7.1, 6.7, 7.3, 7.4, 6.2, 5.6, 5.3, 5, 4.9, 
    5.3, 4.7, 2.8, 3.1, 3.4, 4.9, 6.4, 5.5, 1.4, 3.9, 5.3, 6.2, 5.5, 3.2, 
    3.4, 3.3, 0.7, 1.3, 1, 1, 4.4, 1.5, 3.1, 3.6, 3.3, 4, 8.4, 5.7, 4.4, 3.2, 
    3.7, 3.2, 3.2, 2.9, 3.3, 4.2, 5.1, 4.7, 5.7, 5.9, 4.3, 2.7, 2.8, 3.6, 
    3.2, 7, 2.7, 4.4, 2.7, 6.5, 5.6, 0.5, 5.6, 4, 3.4, 3.3, 5.2, 7.1, 9.5, 
    10.4, 9.3, 10.8, 9.4, 9.3, 9.3, 11, 11.5, 10.3, 9.2, 8.4, 5.5, 3.4, 1.3, 
    0.5, 3.3, 4.3, 4.8, 4, 4.4, 4.3, 5.8, 5.4, 5, 3.1, 2.8, 3.4, 1.3, 0.8, 
    1.2, 1.6, 1.9, 2, 1.8, 3.9, 3.3, 2.1, 1.9, 0.6, 0.9, 3.7, 5.8, 4.4, 8.1, 
    11.7, 7.5, 6.2, 6, 6, 5.1, 4.3, 1.9, 2.6, 2.2, 2.1, 1.7, 0.7, 1.7, 3.4, 
    3.8, 3.5, 4.6, 6.5, 9.3, 8.8, 8.7, 8.5, 8.7, 9, 9.7, 6.7, 8.7, 7.7, 5.1, 
    4.9, 10.7, 9.3, 9.8, 7, 2.1, 4.1, 2.2, 3.4, 3.2, 7.2, 4.3, 2.6, 4.2, 3.7, 
    4.2, 2.3, 6.3, 9.5, 4.2, 6.7, 6.8, 6.7, 3.6, 3.2, 3.8, 2.4, 2.5, 2, 2.8, 
    3.3, 3.1, 2, 2.6, 4.6, 10.6, 9.9, 14, 13.7, 11.3, 12.6, 9.2, 12.7, 14.9, 
    16, 13.9, 14, 11.7, 12.1, 11.1, 9.1, 11, 15.9, 14.7, 16, 14.5, 12.9, 
    11.4, 12.5, 15.5, 16.1, 15.1, 16.1, 16.6, 16.7, 16.6, 17.1, 17, 19.4, 
    19.2, 20.6, 19.5, 19.1, 18.8, 18.7, 18.1, 18.9, 18.6, 17.7, 15.6, 15.4, 
    17.8, 17.5, 15.7, 14.7, 12.7, 12.6, 12.5, 11.2, 7.9, 8.5, 9.7, 8.2, 6.8, 
    6.6, 5.4, 7.2, 7.8, 8.9, 9.4, 10.7, 10.5, 10.8, 10.1, 11.3, 11.4, 11.5, 
    11.7, 11.9, 12.5, 13, 12.7, 13.5, 13, 13.5, 12.7, 12.7, 13.5, 14.6, 13.9, 
    14.3, 14.6, 14.2, 13.7, 15, 17.3, 15.8, 15.1, 14.9, 15.4, 15.7, 16, 16.9, 
    17.8, 16.3, 15.2, 15.5, 15.8, 14.2, 13.4, 13.9, 13.8, 12.9, 12.7, 12.2, 
    13.3, 11.7, 12.8, 12.6, 13, 12.8, 10.4, 9.1, 8, 9.2, 10, 11.2, 10.7, 
    10.5, 11.2, 10.3, 9.5, 10.1, 7.4, 7.4, 8.3, 7, 6.4, 7.8, 8.1, 7.5, 8.1, 
    8.1, 8.4, 8, 7.4, 7.5, 7, 6.8, 6, 4.4, 5.7, 2.9, 3.8, 3.9, 5.4, 5, 4.9, 
    4.7, 3.6, 3.1, 4, 6.7, 8.7, 8.3, 6.6, 7.6, 7.5, 8.7, 11.3, 10.4, 9.4, 
    12.1, 14.3, 15.8, 17.3, 17.6, 19.5, 21, 23.5, 22.7, 25.2, 25.6, 26.9, 27, 
    25.5, 23.7, 20.5, 20.3, 19.5, 19.5, 18.2, 19, 20.4, 18.7, 16.3, 16.6, 
    18.4, 17.7, 16.6, 18.2, 17.4, 16.3, 19.2, 18.9, 18.6, 19.4, 21.1, 21.8, 
    19, 19, 20.3, 19.5, 18.9, 19, 21.4, 19.9, 18.1, 16.2, 9.5, 3.5, 11.6, 
    11.6, 8.4, 11.9, 9.5, 9.8, 9.1, 6.7, 6.8, 7.4, 9, 10, 9.5, 8, 9, 9, 9.1, 
    10.3, 7.8, 7.7, 4, 9.3, 10, 7.2, 10.6, 9.8, 8.9, 8.5, 8.4, 8.5, 9.6, 9.6, 
    9.2, 9.3, 10.4, 10.3, 9.6, 11.1, 10.4, 11.6, 12.7, 13.7, 17.5, 18, 20.4, 
    19.9, 19.3, 18.1, 16.3, 19.1, 20, 19.6, 16.4, 4.3, 14.5, 17.4, 12.3, 
    11.1, 14, 12.1, 12.6, 15.9, 15.9, 15.6, 13.4, 10.4, 12, 12.6, 12, 10.4, 
    10.7, 9.8, 9.8, 8.1, 10.1, 8.8, 4.8, 7.8, 7.5, 8.9, 8.3, 10.8, 12.4, 9.2, 
    9, 9, 8.3, 10.3, 10.9, 10.6, 12.1, 13.5, 13.5, 13.2, 15.3, 13.6, 12.3, 
    12.1, 12.8, 12.1, 12.3, 9.9, 10.3, 10.9, 12.6, 9.7, 9.6, 9.7, 10, 11.1, 
    11.5, 9.1, 8.5, 8.4, 7.8, 4.7, 3.7, 3.1, 3.4, 3.3, 10.8, 11.3, 11.6, 
    12.3, 12.9, 14.5, 11.1, 10, 9.2, 8.7, 7.9, 5.3, 3.6, 9.8, 11.1, 10.5, 
    9.3, 8.2, 6.9, 6.8, 5.5, 5.3, 6.3, 5.7, 6.9, 8.5, 7, 6, 6.3, 6.5, 6.2, 
    5.5, 5.7, 7.2, 9.6, 6.5, 4.7, 5.9, 7.9, 9.9, 9.7, 7.6, 9, 7, 7.9, 6.9, 
    3.6, 9.4, 10, 10.5, 9.1, 2.3, 6.7, 7, 9.1, 8.4, 9.2, 9, 10.8, 11.9, 10.4, 
    11.3, 10, 8.5, 8, 8.1, 8.7, 8.3, 7.4, 6.7, 5.1, 3.5, 3, 4.3, 3.6, 4.6, 
    2.6, 2.6, 3.2, 1.8, 2.9, 1.9, 2.9, 2.7, 3.4, 4.1, 4.9, 1.9, 3.8, 4.5, 
    7.1, 7.4, 8, 9.9, 9.5, 9.2, 8.8, 6.9, 7.2, 7.7, 10.4, 10.9, 10, 10.1, 
    8.4, 8.9, 10.7, 6.5, 8.6, 7.1, 5, 3.8, 1.7, 7.1, 7.5, 6.7, 4.8, 4.6, 3.2, 
    4, 4, 3.2, 2.7, 3, 4.6, 3.5, 3.5, 3.7, 4, 4, 4, 5.2, 5, 5, 7.7, 7.3, 5.9, 
    6, 7.5, 7.6, 7.6, 7.6, 8.8, 8.7, 8.5, 9.1, 9.9, 9.8, 9.9, 9.7, 9.8, 10.9, 
    11.5, 11.8, 10.9, 11.7, 11.9, 12.2, 11.6, 12.5, 10.7, 10.1, 9.5, 8.5, 
    7.9, 6.3, 4.9, 10.8, 12.3, 14.4, 11.1, 12.9, 13, 14.6, 15.2, 16.1, 16.6, 
    15.3, 15.8, 21.1, 22, 21, 19.1, 17.6, 17.5, 18.1, 16.4, 17.3, 15.7, 13.8, 
    13, 13.1, 13.2, 12.9, 11.6, 11.5, 11.3, 10.8, 9.9, 8.9, 8.8, 8.9, 8.7, 
    8.2, 8.1, 8.3, 7.9, 7.1, 7.3, 7, 6.4, 5.8, 4.8, 4.5, 3.7, 3, 3, 3.3, 3.8, 
    3.1, 6, 9.1, 8.9, 7.9, 9.1, 10.4, 13.1, 11.8, 11.9, 10, 9.9, 7, 7.5, 6.3, 
    5.8, 3.9, 2.1, 2.6, 1, 1.5, 4, 1.8, 4.9, 3.9, 3.9, 6.4, 7.2, 5.7, 6.9, 
    6.5, 5.8, 6.6, 7.3, 6.8, 6.5, 6.4, 5.8, 4.8, 4.4, 3.6, 2.7, 2.5, 3.3, 
    3.8, 4.3, 4.7, 4.9, 5.5, 6.2, 6.7, 6.8, 6.8, 3.6, 5.1, 6, 5.3, 5, 5.1, 
    8.3, 9.2, 10.5, 11.4, 12.9, 14.3, 14.8, 14.5, 15.7, 18.6, 18.8, 18.5, 16, 
    15.2, 14.2, 13.8, 9.2, 11.9, 10.4, 2.9, 29.1, 30.6, 29, 28.6, 27.5, 28.4, 
    27.7, 28, 28.3, 26.5, 27, 25.7, 23.2, 12.8, 12.1, 11.8, 1.2, 13.5, 13.1, 
    12.4, 12.4, 12.4, 8.9, 8, 7.8, 8.7, 8.9, 8.8, 8.9, 6.9, 12.4, 12.9, 11.3, 
    11.5, 10.3, 12.4, 13, 13.9, 13, 12.7, 10.2, 12.3, 10.9, 10.2, 7.6, 6.2, 
    5.7, 5.5, 2.4, 2.7, 5, 7.1, 7.8, 8.7, 9.3, 9.3, 8.8, 9.7, 8.9, 9.1, 7.4, 
    9.5, 9, 9.9, 8.7, 10.4, 8.6, 9.9, 8.7, 11.5, 7.7, 8.3, 7.2, 6.1, 6, 7.8, 
    5.8, 4.6, 5.6, 8.4, 9.2, 13.6, 15.2, 16.2, 18.5, 19.8, 20.7, 19.7, 19.9, 
    19.2, 16.8, 15.7, 15, 15.6, 15.3, 13.4, 11.2, 11.2, 11, 11.8, 12.5, 11.6, 
    10.9, 10.5, 10, 8.5, 7.8, 7.2, 5.9, 3.6, 5, 6.2, 7.8, 8.9, 8.7, 9, 9.5, 
    9.6, 9.6, 11, 11.8, 12.2, 11.3, 11.9, 13.1, 14, 14.6, 13.9, 13.6, 14.1, 
    15.1, 15, 14.7, 16.1, 15.7, 16.8, 17.5, 17.1, 16.6, 17.2, 16.7, 17, 17.4, 
    17, 16.3, 16.4, 15.9, 16, 15.6, 16, 16.7, 15.4, 16.5, 16.5, 15.5, 15.9, 
    16.1, 16.6, 15.5, 15.8, 14.7, 14.9, 15.2, 15.3, 14.6, 14.1, 13.5, 12.9, 
    12.4, 11.7, 11.6, 11.9, 11.2, 11.1, 11.2, 11.6, 11.5, 11, 10.7, 10.5, 
    11.4, 11.3, 11.4, 11.3, 11.3, 11.3, 11.1, 10.7, 11.1, 11.1, 10.1, 9.7, 
    9.3, 10.2, 8.8, 8, 7.8, 7.7, 7.9, 8.2, 6.8, 6, 5.9, 7, 6.7, 6, 5, 5.1, 
    5.7, 6.6, 6.7, 7.3, 7.7, 7.8, 8.6, 8.5, 8.3, 8.3, 7.9, 7.2, 7.5, 8.6, 
    8.3, 8.6, 8.3, 8.4, 8.9, 8.2, 8.8, 8.6, 9, 8.4, 8.5, 9.1, 8.6, 9.4, 9.5, 
    9.9, 9.5, 8.9, 10.2, 10.2, 9, 9.7, 10.2, 9.7, 8.8, 8.9, 8.4, 7.5, 8, 9.5, 
    8.8, 8.1, 7.5, 7.7, 6.8, 6.9, 5.8, 6.1, 6.4, 5.6, 5.7, 7, 6.5, 5.8, 9.1, 
    8, 3.3, 5.5, 3.6, 3.9, 0.6, 0.2, 2.6, 1.8, 0.2, 0.9, 2.8, 5.7, 4.1, 4.4, 
    4.3, 13.9, 14.3, 15.1, 15, 14.5, 15.6, 19.7, 18.6, 19.6, 23.3, 22.2, 
    21.5, 21.4, 20.6, 19.8, 17.3, 13, 11.1, 10, 8.4, 6.5, 3.2, 5.2, 4.4, 5.9, 
    9.8, 10.1, 10.9, 12.9, 10.9, 11.5, 9.7, 9.9, 8.4, 8.5, 10.1, 9.8, 7.6, 
    5.7, 6.4, 7.8, 6.1, 7.5, 9, 8.4, 7.3, 8.4, 9.2, 8.8, 9.8, 10.4, 10.8, 
    11.1, 13.5, 13.7, 14.7, 15.8, 14.2, 13.8, 14.4, 15.1, 13.2, 11, 11.6, 
    12.2, 11.4, 12.5, 11.9, 12.1, 9.9, 8.5, 8.4, 7.4, 7.4, 7.5, 8.5, 5.8, 
    10.1, 10.4, 8.1, 5.1, 5.5, 7.8, 8, 7.9, 8, 6.5, 10.7, 14.6, 15.3, 15, 
    15.4, 14.9, 14, 12.3, 14.3, 17.1, 16.5, 14.7, 15.5, 14.8, 14.6, 15.3, 
    15.8, 16.3, 14.2, 14.5, 18.4, 16.6, 19, 16.9, 17.3, 15.5, 15.5, 16.6, 
    17.8, 16.1, 16.6, 15.8, 13.9, 13.6, 15.3, 18.7, 19.3, 19.1, 17.5, 15.2, 
    15.8, 12.8, 12.1, 11.1, 12.5, 11.8, 11.9, 12.4, 13.1, 14.3, 13.1, 12.4, 
    13.1, 14.4, 14.3, 15.2, 15, 12.7, 11, 13.6, 15, 13.1, 12.8, 12.8, 14, 
    14.6, 14, 14.1, 13.9, 13.7, 13.6, 14.7, 13.4, 10.8, 9.5, 8, 7.6, 7.7, 
    8.8, 9.9, 10.2, 11.5, 9, 11.3, 11.5, 8.7, 7.1, 5.7, 6.6, 7.2, 6.1, 6.5, 
    5.5, 5.5, 8, 7.9, 7.6, 7.2, 6.6, 6.8, 8.8, 9, 9.2, 9.3, 9.1, 8.3, 6.4, 
    5.6, 4.7, 5.4, 7.3, 7.4, 7.8, 7.6, 7.9, 7.4, 8, 7.3, 8.7, 6.3, 7.2, 6.9, 
    6.7, 6.3, 5.2, 7, 6.8, 7, 7, 7.5, 6.3, 6.6, 7.9, 7.8, 7.3, 7.2, 5.7, 7.7, 
    8.9, 7.6, 5.8, 8.5, 9, 9.6, 9.7, 9.6, 9.4, 9.6, 10.5, 9.6, 10.1, 10.1, 
    11.7, 10.6, 10.6, 10.1, 10.4, 7.4, 6.3, 4.1, 5, 9.4, 9.9, 6.1, 7.1, 8.1, 
    9.6, 8.5, 8.5, 10, 9.8, 8.9, 7.4, 5.6, 4.7, 5.3, 6.3, 5.5, 5.4, 2.6, 3.3, 
    0.4, 1, 1.9, 0.2, 0.2, 0.5, 0.5, 1, 1.8, 2.1, 4.1, 5.5, 3.4, 4.2, 6, 6.4, 
    5.9, 7, 6.7, 6, 5.9, 5.8, 7.7, 10.5, 9.2, 11.4, 9.1, 10, 11.8, 10.3, 
    10.4, 10.9, 12.3, 12.5, 11.9, 12.9, 12.8, 11.7, 13.2, 11.2, 8.7, 6.8, 9, 
    7.7, 6.9, 6.9, 10.3, 11.5, 11.7, 8.7, 7.5, 11.9, 4, 2, 1.1, 2.3, 3.1, 
    5.9, 2.2, 1.8, 3.8, 3.1, 3.6, 7.2, 12.7, 9.3, 10.4, 8.7, 6.8, 5.6, 9, 
    10.9, 12.6, 2.7, 1.7, 3.1, 7.6, 5.1, 4.3, 1.6, 4.7, 4.1, 5.7, 8.5, 6.8, 
    6.4, 8.4, 8.3, 11.8, 15.4, 14.9, 15.1, 13.9, 1, 0.8, 3.1, 8.4, 10.4, 
    10.6, 11, 8.5, 8.9, 8.9, 9, 4.4, 5.3, 4.4, 3.1, 8.4, 7.3, 9.5, 9, 9.2, 
    8.7, 9.1, 10, 10.7, 10.8, 9.7, 8.8, 8.6, 8.6, 8.8, 11.7, 11, 10.7, 10.5, 
    11.1, 13.2, 12.2, 14.2, 12.1, 11.1, 10.2, 9, 8.8, 10.2, 10.1, 9.5, 8.9, 
    10.5, 9.4, 10.2, 10, 10.1, 8.8, 8.8, 9.3, 8.6, 8.3, 8.3, 8.5, 8.1, 8.9, 
    8.9, 9.5, 9.6, 9.3, 9.2, 8.5, 8.3, 9.2, 9.5, 8.8, 9.1, 8.4, 8.6, 8.3, 
    8.5, 8.1, 8.7, 9.4, 9.1, 10.1, 8.1, 9.7, 8.3, 9.9, 9, 8.2, 9.5, 9.2, 9, 
    9.1, 9.6, 9.3, 8.7, 7.8, 9.1, 9.3, 10.1, 9.6, 7.2, 8.1, 8.3, 2.5, 1.4, 
    2.1, 5.6, 4.4, 4.2, 0.6, 6, 3.7, 3, 1.1, 0.8, 1.1, 3.6, 3.1, 1.1, 1.8, 
    6.8, 8.6, 8.5, 9.1, 9.4, 6.8, 5.1, 1.1, 0, 0, 3.3, 0, 0, 2.4, 2.6, 1.6, 
    0, 1.1, 4.1, 5.1, 5.9, 5.1, 3.3, 3.2, 3, 2.7, 1.1, 0, 0.4, 0.4, 2.2, 2.8, 
    2.3, 1.1, 0.2, 0, 0, 0, 4.5, 4.2, 3.7, 3.3, 3, 3.9, 1.4, 1, 0.7, 1.5, 
    1.6, 0.4, 2.8, 5.5, 6, 9.7, 11.5, 9.8, 9.7, 9.7, 9, 8.8, 10.7, 11.1, 
    14.3, 10.7, 13.8, 9.5, 10.9, 10.9, 12.5, 13.5, 14.6, 13, 10.9, 12.4, 
    12.8, 8.5, 12.2, 10.7, 9.3, 9.5, 9.8, 11, 11.9, 14.1, 15.5, 13.2, 13.1, 
    14.7, 17.6, 15.1, 17.2, 17.6, 16.8, 18.7, 18, 16.5, 16.3, 16, 15.2, 14.1, 
    11.5, 10.2, 10.3, 9.8, 9.5, 9.5, 8.3, 8, 9.4, 10.3, 11.5, 11.3, 12, 11.2, 
    10.7, 9.9, 10.2, 10.2, 10.1, 10.2, 10.5, 10.8, 10, 9.3, 9.6, 9, 9.4, 7.7, 
    7.7, 8, 7.4, 6.9, 7, 8.5, 9.2, 7.4, 9.9, 8.7, 8.1, 7.3, 4.6, 5, 4.4, 4.9, 
    6.1, 7.7, 9.9, 9.4, 2.8, 3, 1.7, 2, 3, 2.5, 1.6, 3.1, 4.1, 3.7, 4.1, 3.2, 
    3.2, 4.5, 4.2, 3.7, 2.9, 2.2, 3.8, 3.2, 1.5, 2.9, 2.1, 3.5, 4.3, 4.2, 
    4.9, 4.2, 2.3, 1.9, 2.4, 3.5, 4.7, 4.8, 4.6, 3.5, 12, 10.7, 10.1, 11.4, 
    13.2, 10.8, 13.8, 15.6, 19.9, 18.8, 17.7, 17.8, 17.7, 17.4, 17.8, 17.7, 
    17.2, 16.2, 15.8, 13.3, 13.2, 14.2, 13.8, 12.9, 14.2, 13.8, 15.4, 17.3, 
    17.3, 15, 14.4, 12.1, 10.8, 7.6, 7.1, 10.2, 11.4, 10.3, 11, 11, 11, 11.5, 
    12.1, 12.2, 11.7, 1.4, 5.7, 3, 3.4, 5.2, 6.2, 6.2, 6.6, 6.2, 5.9, 6.5, 
    8.3, 7.8, 11.3, 12.3, 9.5, 8.5, 7.8, 7.9, 8.6, 5.5, 6, 8.7, 9.6, 7.3, 
    5.3, 6.3, 5.5, 7.8, 7.9, 8.4, 7, 9.2, 14.2, 13.8, 11.9, 10, 8.9, 8.8, 
    8.6, 9.4, 6.7, 8.9, 9.4, 7.9, 7.9, 8.4, 7.4, 7.7, 8.3, 9.6, 11.4, 9.1, 
    9.8, 11.6, 12.3, 11.1, 8.5, 11.2, 10.9, 10.3, 9.1, 8.9, 10.1, 11.4, 10.6, 
    9.9, 11.1, 10, 10.3, 10.9, 9.1, 11, 10.4, 10.4, 10.2, 9.1, 10.6, 9.9, 
    9.6, 9.6, 7.7, 8.1, 7.1, 6.5, 6.9, 8.5, 8, 10.4, 7.6, 8.5, 6.2, 6, 5.4, 
    9.9, 7.8, 7.1, 7.9, 7.9, 8, 8.4, 8, 8.9, 7.9, 6.9, 8.1, 6.9, 8.5, 8.8, 
    6.6, 6.9, 7.2, 5.9, 5.8, 5.2, 6.2, 5.3, 4.6, 4.5, 4.1, 3.5, 3, 2.5, 4.7, 
    4.7, 4.6, 3.7, 3.9, 3.6, 4.5, 3.2, 3.1, 2.3, 2.7, 2.5, 5.4, 5.6, 6.7, 6, 
    5.8, 4.5, 4.2, 4.9, 5.8, 10.2, 7.9, 11.9, 11.2, 11.4, 11.6, 10.9, 8.9, 
    8.8, 8.5, 6.4, 5, 4.5, 3.2, 3.9, 1.2, 1.9, 1, 3.8, 5.5, 5.8, 7.8, 8, 8.7, 
    9.1, 10.1, 10.7, 10.9, 10.9, 11, 9.4, 7.6, 8, 6.2, 3.5, 2.6, 0, 0.8, 1.1, 
    1.2, 0, 0.9, 0.5, 2.1, 4.1, 7.6, 7.3, 9.6, 10.6, 9.7, 8.6, 6.1, 7, 7.1, 
    6.9, 7.4, 9.2, 9.1, 8.9, 9.3, 10.5, 8.4, 8.5, 7.2, 7, 8.3, 7.6, 8.1, 7.2, 
    7.4, 7.6, 7.6, 6.9, 6.5, 5.5, 4.5, 3.5, 2.7, 1.7, 1.9, 3.3, 2.4, 3.7, 
    2.7, 3.9, 4.4, 6, 6.3, 7.5, 8.6, 9.4, 9.5, 10.3, 11.7, 11.5, 11, 11.1, 
    10.7, 12.1, 12.7, 11.8, 11.1, 10.6, 11.6, 12.1, 10.8, 11.3, 10.7, 10, 
    9.7, 8.1, 6.3, 5.6, 4.1, 1.9, 8.4, 9.8, 11.6, 9.9, 7.8, 8.3, 7.7, 7, 8.1, 
    8.4, 8.7, 7.4, 8.6, 8.6, 8.8, 10.3, 11.2, 9.9, 11, 9, 9.8, 9.5, 9, 8.6, 
    8.4, 9.6, 10.6, 5.2, 4.2, 3.6, 2, 2.1, 0.7, 1, 4.6, 6, 7.4, 8.3, 8.2, 
    8.3, 8.9, 8.1, 7.7, 6.9, 8.9, 9, 8.1, 8.2, 8.9, 5.5, 5.5, 5, 1.1, 0.6, 
    1.3, 1.5, 1.8, 6.2, 9.7, 8.3, 11.6, 10, 8.9, 9.7, 10.9, 9.4, 8.5, 10, 
    10.7, 9.6, 10.5, 13.8, 12.8, 12.3, 10.9, 12.1, 12.8, 10.1, 11.8, 15.1, 
    15.4, 14.2, 13, 11.3, 13.4, 14, 14.8, 13.3, 13.8, 12.7, 11.7, 10, 10.8, 
    11, 8.7, 11.2, 10.3, 10.5, 12.2, 12.2, 12.2, 11.6, 10.9, 10.3, 8.8, 8.9, 
    10.1, 13.5, 13.8, 13.1, 14.6, 15.5, 15.1, 13.4, 16.7, 17.4, 16.3, 17.8, 
    17.8, 13.8, 18.7, 18.1, 17, 13.5, 17, 16.4, 16.5, 16.3, 16.3, 15.8, 15.7, 
    15.7, 16, 14.9, 12.9, 11.8, 13.2, 12.9, 11.6, 11.1, 11.5, 10.2, 11.7, 
    11.3, 11.1, 11.9, 12.1, 11.1, 10.9, 10, 10.5, 9.6, 8, 9, 9.7, 9.5, 8.2, 
    8.2, 6.8, 6.5, 6.9, 7.6, 7.5, 7.8, 7.4, 6.3, 7.5, 7.6, 8.2, 6.8, 6.4, 
    7.4, 8.2, 8.8, 10.5, 9, 8.3, 7.2, 7.3, 7.6, 8, 7.2, 8, 7.4, 7.2, 6.4, 
    6.5, 6.3, 6.9, 6.5, 6.1, 6.4, 6.4, 6.2, 7.3, 6.9, 6.2, 6.9, 6.4, 6, 6.7, 
    6.9, 6.7, 6.8, 7.7, 7.3, 6.1, 7.1, 6.5, 7.1, 5.1, 2.7, 2.1, 1.1, 1, 0.8, 
    1.7, 0, 1.3, 0.5, 1.7, 1.6, 1.8, 2.2, 1.3, 2.2, 2.2, 2, 2.4, 2.3, 2.3, 
    3.4, 3, 3.9, 3.7, 2.5, 3.6, 1.9, 1.1, 0.1, 2, 0, 0.8, 1.5, 1.9, 3.8, 1.7, 
    2.4, 1.2, 1.1, 2.3, 2.7, 3.3, 3.7, 3.9, 4.7, 3.7, 4.7, 3.9, 4, 5.2, 4.3, 
    4.7, 4.8, 3.7, 4, 2.8, 4.2, 4, 3.4, 4.3, 3.6, 4.4, 3.3, 3.1, 3.2, 2.6, 
    2.8, 3, 3.2, 3.8, 4.4, 5.7, 4.8, 6, 5.1, 5.3, 4.5, 5, 5.3, 4.2, 4.7, 4.4, 
    2.9, 3.4, 2.3, 3.5, 3, 3.4, 3.8, 3, 3.8, 4.4, 4.1, 5, 6.1, 6.3, 7.5, 7.1, 
    7.5, 7.5, 7.5, 7.9, 8.2, 6.9, 6.7, 7.3, 5.5, 6.1, 6.5, 4.9, 4.1, 3.6, 
    4.4, 8.4, 10.4, 10.8, 11.7, 13.1, 13.6, 14, 13.4, 12.9, 13.3, 13.9, 13.5, 
    12.5, 10.8, 10.5, 10.6, 11.1, 10.5, 10.9, 11.5, 13, 11.6, 13.1, 14.9, 
    15.7, 15, 15.2, 16, 16.3, 16.8, 15.4, 15.5, 13.8, 13.6, 13, 9.1, 8.7, 
    9.7, 11.8, 9.9, 11.1, 11.6, 14.5, 13, 9.4, 9.3, 10.6, 13.3, 12.3, 9.1, 
    7.1, 7.1, 6.8, 7, 6.7, 7.9, 9.4, 6.4, 8.9, 5.8, 6.5, 5.2, 5, 6, 5.6, 6.1, 
    5.8, 5.4, 5.9, 6, 5.9, 6.4, 4.9, 5.4, 5.4, 3.8, 4.8, 3.9, 4.5, 4.3, 3.2, 
    2.8, 2.7, 3.9, 3.8, 4, 3.3, 4.2, 3.4, 3.9, 3.6, 3.1, 2.7, 2.9, 3.2, 2.9, 
    3.1, 3, 2.4, 4.1, 2.7, 2.8, 4.7, 2.9, 4, 3.1, 3.1, 2.1, 1.2, 1.5, 0.4, 
    0.2, 1.9, 1.7, 1.8, 3, 3.1, 3.4, 3.5, 4.7, 4.2, 4.6, 5, 5.2, 5.1, 4.7, 
    4.5, 5.4, 4.9, 5.5, 4.3, 5.9, 5.2, 5.8, 6.1, 5.3, 7.1, 7.4, 8.3, 8.3, 
    8.1, 8.9, 8.3, 6.9, 6.4, 5.7, 5.7, 5.4, 5.1, 5.2, 4.4, 3.8, 3.6, 3, 0.8, 
    7.6, 7.8, 8.8, 8.8, 6.7, 9.8, 8.6, 9.5, 9.6, 10.5, 10.5, 10.9, 9.1, 8.3, 
    7.9, 7, 4.9, 3.7, 2.9, 5.9, 3.6, 4.8, 5.6, 7.7, 6.4, 5, 3.6, 2.7, 2.3, 
    2.6, 2.8, 5.3, 6.3, 6.7, 7, 7.1, 7.4, 7.1, 7.5, 6.9, 6.2, 5.1, 5.1, 2.9, 
    3.5, 3.8, 3.3, 3.9, 4.9, 4.8, 6.3, 4.5, 3.3, 4.7, 6.1, 5.8, 4.8, 6.1, 
    6.7, 5, 3.3, 3.6, 4.4, 6.6, 8.3, 7.2, 6.5, 5.5, 7, 6.3, 8.2, 8, 6.7, 8.5, 
    10, 11.8, 10.8, 12.6, 10.3, 8.9, 9.8, 10.6, 10.2, 9.8, 8.8, 8.1, 8.2, 
    8.3, 7.8, 7.8, 6.9, 8.7, 8.2, 8, 7.7, 7.4, 6, 7, 6.4, 4.9, 4, 3, 5.6, 6, 
    4.9, 4.7, 5.4, 3.5, 3.1, 4.8, 3, 3.1, 3.1, 2.7, 2.6, 3.1, 3.8, 3.6, 1.6, 
    1.6, 0.7, 0.6, 0, 0, 0.2, 2.5, 1.7, 0.8, 1.1, 0.7, 0.9, 1.1, 1.3, 1.3, 
    1.3, 1.5, 1.7, 1.8, 2.1, 2.5, 3, 4.7, 4, 3.8, 3.8, 4.4, 4.6, 5.1, 5.4, 
    6.9, 4.1, 4.2, 4.5, 4.5, 5.1, 5.2, 5.7, 6.3, 5.5, 6.8, 6.6, 7.7, 8.8, 
    8.5, 8, 7.5, 5.2, 4, 4, 3.7, 6.2, 8.1, 8.6, 11.9, 15.3, 14.2, 13.5, 15.3, 
    13.9, 16.1, 12.8, 13.4, 11.2, 11.7, 9.8, 9, 8.7, 9.3, 8.8, 8, 9, 6.7, 
    7.1, 7.5, 8.3, 9.6, 9.3, 6.9, 12.1, 13.6, 12.9, 11, 15.4, 16.1, 15.8, 
    15.2, 14.5, 14, 12.5, 13.8, 13.6, 11.9, 9.7, 9.8, 5.8, 8.4, 10.1, 6.8, 
    11, 2.9, 2.5, 4, 8, 7.9, 2.8, 6.1, 4.9, 5.3, 5, 4.2, 4.3, 4.6, 4.9, 5.2, 
    6, 6, 4.9, 4.3, 4.4, 6.5, 4.9, 5.5, 5.8, 5.5, 6.5, 6.6, 3.6, 4.1, 3.5, 
    3.5, 2.3, 1.8, 2.5, 3.6, 0.6, 2.9, 3.3, 2.5, 2.5, 2.7, 2.6, 2, 1.8, 2.1, 
    1.6, 2.5, 1.5, 1, 0.3, 2, 1.8, 1.7, 1.8, 1.6, 0.6, 0.6, 1.9, 2, 1.9, 2, 
    2, 2.5, 1.6, 2.3, 3.2, 2.9, 3.8, 4.9, 5, 4.4, 4.6, 5.8, 6.1, 7.3, 6.5, 
    5.8, 5.6, 5.6, 4.7, 5.3, 4.8, 2.7, 2.3, 3.1, 3, 2.6, 2.5, 2.6, 3.4, 3.5, 
    3.5, 3.5, 3.1, 2.4, 1.7, 1.4, 1.5, 2, 3, 4.2, 5.6, 7.1, 7.6, 6.9, 5.5, 
    5.5, 5.8, 4.5, 3.1, 4.4, 4.4, 4, 3.7, 3.7, 3.8, 3.3, 3.5, 3.7, 3, 2.9, 
    3.1, 2.3, 1.7, 1.4, 1, 0.8, 1.7, 1.6, 0.7, 0.6, 2.4, 0.5, 1.7, 0.8, 1.8, 
    1.1, 2.2, 0.7, 0.1, 0, 0.9, 1.2, 4.7, 4.9, 5.1, 4.7, 5.3, 5.4, 6.6, 6.2, 
    7.4, 8.1, 7.6, 8.9, 8.5, 9.7, 6.5, 6.8, 6.5, 7, 8.3, 8.7, 8.3, 8, 7.7, 
    7.7, 6.9, 5.8, 3.7, 2.6, 6.4, 7, 4.9, 3.2, 2.9, 2.3, 2.7, 1.8, 1.1, 0.1, 
    3.2, 3.3, 3.7, 4, 4.1, 3.9, 2.8, 3.1, 2.6, 1.9, 3.8, 4.9, 4, 4.7, 3.5, 
    3.7, 5.7, 5, 4.3, 2.3, 2.8, 2.8, 2.6, 2.3, 1.8, 2.6, 1.5, 1.2, 0.6, 1.7, 
    2.7, 2.9, 3.3, 4.3, 5.3, 4.8, 4.3, 4.6, 5, 5.3, 5.6, 6.1, 6.1, 6.9, 6.6, 
    7.2, 7.8, 7.6, 8.4, 9.7, 8.6, 8, 5.7, 7.1, 7.7, 5, 6.1, 6.8, 6.8, 7.9, 
    8.3, 9.7, 8, 8.3, 7.9, 6.6, 6.4, 6.5, 4.7, 4.5, 3.8, 3.5, 2.4, 3.3, 1.5, 
    1, 1.4, 1.3, 0.7, 0.9, 5.4, 6.4, 8, 10.2, 11.6, 11.9, 9.5, 8.7, 9.4, 8.4, 
    8, 8.3, 6.7, 6.5, 6.8, 5.9, 5.3, 5.1, 5.2, 6.3, 6.4, 6, 6.7, 6.8, 6.4, 
    5.2, 5.2, 5.5, 7, 8.1, 8, 8, 7.9, 7.4, 8, 8.2, 7.3, 6.7, 5.6, 7.7, 8.2, 
    8.6, 7.9, 8.5, 7.7, 8.7, 9.9, 10, 10.8, 8.9, 8, 7.3, 8.6, 9.7, 11.4, 9.6, 
    7.1, 7.9, 7.8, 10.2, 7.9, 6.6, 7.6, 9, 8.9, 13.6, 11.6, 11.7, 10.6, 11, 
    11.1, 8.4, 10.5, 12, 12.9, 12.1, 12.4, 12, 10.6, 8.8, 7.5, 6.2, 6.7, 6.3, 
    4.8, 2.4, 1.5, 5.3, 4.9, 8.6, 6.8, 4.5, 5.4, 4.5, 3.9, 4.4, 4.4, 5.7, 
    5.8, 6.3, 6.8, 5.9, 5.5, 4.5, 5.8, 5.4, 5.4, 6.1, 5.8, 6, 5.1, 4.9, 4.9, 
    4.4, 4, 3.9, 3.3, 3.3, 3, 2.5, 2.3, 2, 1.9, 2.1, 1.2, 2.2, 0.5, 1.1, 1.2, 
    2.5, 2.5, 1.9, 2.4, 2.5, 3.4, 3.7, 4.3, 4.9, 4.5, 5.2, 5.7, 6.6, 6.8, 
    6.5, 6.4, 7.4, 8.8, 8.6, 7.7, 8.2, 8.2, 8.2, 8.2, 6.4, 8.8, 7.3, 9, 7.9, 
    9.6, 9.7, 8.3, 8.5, 7.6, 8.4, 9.4, 8.7, 8.1, 7.5, 7.8, 8.2, 6.9, 6.1, 
    6.9, 6.7, 7.8, 7, 8.2, 6.3, 6.2, 6.3, 6.2, 6.2, 6.7, 5.3, 5.4, 4.9, 6.2, 
    6.1, 6, 5.5, 5, 5.2, 5.1, 5.4, 3.8, 3.5, 2.9, 3.4, 3.5, 3, 2.2, 1.9, 1.5, 
    1.1, 0.8, 1.4, 1.3, 3.1, 5, 6.1, 6, 5.5, 5.3, 6, 5, 6, 6.1, 7.3, 5.9, 
    5.8, 5, 4.2, 4.2, 3.3, 6.1, 4.3, 3.5, 3.5, 3.7, 3.6, 6.2, 3.4, 4, 3.9, 
    5.7, 4.5, 3.1, 4.5, 4.9, 4.4, 4, 4, 5.9, 4.7, 6, 6.8, 5.2, 4.5, 5.8, 6.3, 
    6.5, 7.9, 7.1, 9.1, 7.9, 8.4, 8.4, 6.9, 5.7, 5.9, 6.9, 6, 6.2, 5.6, 5, 
    5.9, 5.2, 5.8, 5.7, 7.5, 6.4, 3.7, 3.9, 4, 4, 6.2, 6, 4.9, 6.4, 6.9, 6, 
    4.8, 4.2, 4, 3.8, 3.9, 3.6, 3, 4.6, 4, 2.9, 2.9, 2.6, 3.2, 3.6, 3.6, 3.7, 
    2.3, 2.9, 2, 3.7, 3.6, 3.1, 3, 2.9, 4.1, 4.4, 3.5, 3.6, 5, 4.3, 4.9, 3.2, 
    3.6, 3.4, 4.2, 3.9, 6.4, 5.8, 3.8, 4.6, 4.2, 4.5, 3.8, 3.8, 3, 3.4, 3.8, 
    3.5, 3.6, 2.6, 2.5, 2.3, 2.6, 2.5, 2.4, 2.7, 2.9, 2.7, 3.4, 4.1, 3.3, 
    3.2, 3.2, 2.5, 1.5, 1.5, 0.7, 0.9, 0, 0, 1.2, 2.1, 1.6, 1.9, 2, 2.2, 2.5, 
    2.8, 2.5, 1.7, 1.2, 1.8, 3.1, 2.8, 4, 4.5, 4.6, 4.9, 4.2, 4, 3.4, 3.3, 
    3.9, 4.2, 4.4, 3.7, 5.3, 4.7, 5.5, 5.3, 6.2, 8, 8.8, 9.4, 8.7, 8.1, 7.8, 
    8.4, 7.6, 9, 8.7, 8.5, 7.8, 8, 7.6, 7.5, 7.8, 8.6, 8.5, 8.2, 7.6, 7.4, 
    7.1, 7.1, 6.9, 6.8, 6.6, 6.2, 6.1, 6.4, 6.9, 7.3, 7.8, 7.8, 8.2, 9, 8.6, 
    9.9, 9.3, 8.4, 7.8, 9.2, 9.5, 11.1, 11.3, 12.1, 12, 11.9, 11.2, 11.2, 
    11.1, 10.6, 9.5, 9.5, 8.1, 6.9, 6.3, 5.9, 5.2, 3.9, 4, 2.3, 0.3, 2.6, 
    4.1, 5.6, 5.3, 8.1, 8.1, 8.1, 8.1, 8.7, 7.8, 7.7, 7.7, 6.9, 6.5, 5.9, 
    7.3, 6.9, 7.3, 8, 8.8, 8.1, 8.2, 8.9, 8.1, 7.2, 5.9, 6, 6, 5.9, 3.1, 5, 
    5.2, 5.6, 7, 5.7, 5.7, 5.5, 5.5, 7, 7.3, 8, 7.9, 6.9, 6.8, 7.2, 7.7, 7, 
    6.8, 4, 4.4, 3.7, 4.1, 6.9, 7.7, 6.6, 5.7, 5.2, 4.5, 3.7, 4, 4.3, 3.6, 
    3.1, 3.2, 2.9, 2, 2.1, 3.6, 1.6, 2.5, 2.2, 1.9, 2.6, 2, 2.1, 2.5, 2.6, 2, 
    2.4, 1.5, 1.7, 0.7, 2.2, 1.5, 1, 0.7, 0.7, 2.2, 1.7, 1.6, 2.4, 3.1, 4.7, 
    4.4, 5.4, 4.6, 4.6, 4.7, 5.2, 4.7, 4.7, 4.2, 4.3, 4.5, 4.9, 5.6, 6.2, 
    6.5, 6.6, 6.9, 7.9, 7.1, 8.7, 5.5, 7.8, 6.1, 7.8, 10.4, 9.9, 8.2, 7.6, 
    7.4, 6.6, 6.5, 5.9, 5.5, 4.7, 3.5, 2.4, 1.1, 1.9, 1.4, 1.6, 1.7, 1.3, 
    3.5, 3.4, 3.2, 2.8, 2.7, 3.1, 3.2, 2.3, 2.6, 2.3, 3.8, 3.4, 3.4, 5.5, 
    5.3, 5.2, 2.2, 1.6, 0.1, 1.2, 0, 0.5, 0.6, 1.1, 2.2, 4, 4, 4.6, 5.8, 5.5, 
    3.7, 1.5, 0.6, 0.4, 0.9, 4.7, 3, 1.2, 1.1, 3.2, 3.2, 3.5, 1.8, 5.5, 6, 
    1.6, 1.1, 0.9, 4.4, 2.6, 1.3, 3, 1.1, 1.7, 1.8, 1.6, 1.6, 0.8, 1.2, 0.4, 
    0.7, 0.6, 3.5, 6.9, 3, 8.7, 8.6, 8.5, 8.5, 9.4, 7.6, 8.6, 7.7, 9.6, 9.5, 
    6.3, 8.1, 7.7, 8.2, 9.3, 9.9, 9.8, 9, 8.7, 8.9, 7.7, 7, 7.2, 8, 8.6, 7.8, 
    7.5, 7.4, 7.2, 6.8, 5.5, 5.3, 4.4, 5, 4.9, 4.2, 5, 4.4, 5, 3.9, 2.4, 3.1, 
    4.2, 4.3, 3, 2.8, 1.4, 3.9, 2.8, 1.8, 1.3, 1.2, 1, 1, 1.4, 1.5, 0.4, 1.3, 
    1, 0.5, 0.9, 1, 0.7, 0.9, 0.7, 0.7, 1.2, 2.2, 1.2, 0.5, 1.1, 2.1, 1.5, 2, 
    2.6, 1.3, 1.5, 2.3, 3, 2.8, 3.3, 3.5, 4.2, 4.2, 5.4, 6, 6, 5.6, 6.1, 7.4, 
    7.4, 7.8, 7.4, 6.1, 6.1, 7.9, 9.2, 8.5, 7.8, 6, 7.1, 7.6, 6.7, 6.7, 5.8, 
    4.9, 4.2, 4.1, 4.5, 3.3, 3.3, 3, 3, 3, 3.2, 3.2, 2.6, 2.7, 3.1, 2.8, 2.7, 
    3.6, 2.1, 0.6, 1.7, 2.1, 0.7, 3.7, 0.8, 1.9, 2.1, 2, 2.6, 3.1, 1.7, 3, 
    13.2, 16.6, 17.7, 18.6, 17, 17.3, 18.9, 18.9, 20.3, 16.8, 17, 13, 8.4, 
    3.9, 1, 3.8, 4.4, 2.9, 0.7, 1.1, 2.4, 3.6, 5.6, 6.2, 2.9, 1.2, 2.2, 4.6, 
    1.7, 3, 3.2, 2, 2.1, 2.7, 1.6, 1.1, 1.1, 1.8, 2, 1.8, 2.3, 0.3, 2.2, 4.3, 
    6.2, 5.2, 5.8, 3.3, 6.3, 9.7, 9.7, 7.9, 8.6, 6.4, 6.9, 6.1, 6.6, 8.2, 
    7.8, 8.8, 6.8, 6.2, 5.8, 8.7, 9, 10, 8.1, 9.8, 10.8, 12.2, 14.6, 14.1, 
    14.4, 15.7, 13.6, 16.6, 14.6, 11.8, 7.9, 7.1, 8.1, 7, 6.2, 6.2, 5.8, 5.8, 
    5.8, 5.3, 5.8, 8.3, 7.4, 7.8, 8.8, 8.8, 9.6, 9.9, 11.1, 10.8, 12.3, 10.9, 
    11.6, 9.7, 10.4, 9.9, 8.5, 9.8, 8.7, 9.4, 8.6, 7.9, 7.8, 7.8, 6.6, 5.5, 
    4.5, 4.8, 6.1, 6.6, 8.6, 8.9, 7.2, 5.9, 3.7, 2.4, 2.5, 2.2, 5.2, 3.8, 
    2.4, 2.4, 2.2, 1.3, 1.2, 1.4, 11.4, 5.4, 11.3, 5.4, 2.1, 3.2, 1.4, 3.8, 
    6, 10.3, 10, 8.5, 1.7, 2.3, 2.7, 1.6, 3, 1.5, 2, 4, 4.7, 4.4, 5.1, 4.7, 
    4.7, 6.2, 6.1, 5.3, 3.6, 3.1, 1.4, 3.5, 4.4, 5.8, 7.5, 8.4, 10, 12.2, 
    12.5, 12.1, 11.1, 9.5, 8.8, 8.3, 6.1, 4.8, 4, 3.4, 3.4, 3.3, 3.2, 2.5, 
    1.7, 2.2, 1.4, 4.4, 5.5, 6.4, 6.3, 6.1, 6.6, 6.4, 5.5, 5.2, 4.5, 3.8, 
    2.9, 2.1, 1.6, 1, 0.4, 0.8, 1.9, 4.4, 5.4, 8.4, 9.1, 9.8, 10.7, 11.5, 
    11.8, 11.9, 12, 12.1, 10.1, 11.1, 10.8, 10.6, 9.8, 9.9, 9.3, 9.3, 9.4, 
    8.3, 8.2, 4.6, 2.3, 3.1, 1.9, 2.6, 4.5, 6.3, 5.3, 3.6, 8, 5.5, 2.6, 7, 
    1.2, 6.4, 2.2, 4.5, 1.3, 0.9, 0.6, 1.4, 2.1, 2.5, 4.4, 3.5, 5, 5.1, 5, 
    5.4, 4, 2.4, 2.2, 2.6, 2.8, 2.8, 1.8, 1.6, 1.3, 1.1, 0.9, 2.2, 3, 1.8, 1, 
    0.9, 1.6, 0.7, 0.3, 0.2, 0.6, 1.2, 1.7, 1.6, 4.1, 4.2, 3.3, 3.5, 1.4, 
    2.8, 2.5, 1.2, 1.5, 0.6, 0.5, 0.3, 0.3, 0, 0.4, 0.2, 0, 0, 0, 0, 0, 0, 
    0.5, 1, 0.9, 2, 3.7, 5.3, 5.7, 3, 6.3, 6.5, 6.4, 7.6, 8.7, 7.4, 8.7, 7.9, 
    8.9, 9.3, 9.4, 7.9, 8.3, 6.9, 8.3, 7.7, 7, 6.9, 6.7, 7.2, 3.9, 5.2, 7.7, 
    6.5, 7.2, 7, 7.4, 6.5, 4.4, 3.6, 5.5, 3.3, 3.1, 2.9, 3.6, 3.4, 2.7, 3.1, 
    1.5, 0.5, 0.5, 0.1, 0.1, 1, 2.2, 2.6, 2.2, 2.7, 3.1, 3.4, 2.8, 2.2, 2.3, 
    4, 4.3, 3.4, 4.8, 4.3, 6.8, 8.1, 4.5, 3.5, 2.5, 2.5, 1.9, 1.8, 1.9, 1.5, 
    1.6, 2, 1.7, 1.6, 1.4, 1.1, 1.2, 1, 1, 0.8, 0.7, 0.7, 0.8, 0.6, 0.9, 1.2, 
    1.1, 0.9, 0.9, 0.8, 0.7, 0.5, 0.7, 0.8, 0.6, 0.9, 0.9, 0.8, 0.7, 0.8, 
    0.9, 0.8, 0.9, 0.8, 0.7, 0.8, 0.8, 0.9, 0.8, 0.7, 0.5, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    3.5, 1.4, 0, 0, 0.2, 0.1, 0.8, 1.2, 0.2, 0.4, 0.6, 0, 1.6, 1.7, 0.7, 0.3, 
    0.9, 1.7, 0.8, 0.3, 0.2, 0.7, 0.7, 1.4, 2.8, 2.8, 4, 2.5, 2.4, 3.6, 3.2, 
    4.5, 5.5, 5.5, 5.6, 5.2, 4.9, 3.4, 2.2, 2.1, 2.7, 3.3, 2.5, 1.9, 0, 0, 0, 
    0.2, 1.5, 0, 0.2, 1.2, 0.3, 0.6, 2.7, 2.9, 3.1, 1.6, 2, 0.1, 0, 0.1, 1.5, 
    1.1, 1.3, 0.5, 0.7, 2.6, 3.2, 2.9, 2.3, 1.6, 2.7, 2.8, 2.7, 3.3, 2.3, 
    2.6, 3, 3.2, 2.5, 2.2, 1.7, 1.1, 1.2, 1, 1.3, 0.1, 0.9, 0.8, 0, 0.3, 0, 
    0, 0, 0.2, 0.1, 0.3, 0.7, 0.6, 0.1, 0.1, 0.2, 0.8, 1.4, 1.8, 4, 4.1, 2.7, 
    3.4, 3, 3.4, 3.3, 2.5, 2.5, 2.4, 3.1, 2.5, 1.6, 1, 0.4, 0.1, 0.5, 0.1, 
    0.3, 0.3, 1, 2.2, 3.2, 2.3, 2.7, 1.7, 2, 2, 2.9, 2.6, 1.8, 1.6, 3, 2.5, 
    1.9, 2.9, 3.1, 2.5, 1.9, 2.3, 3, 3.2, 3.6, 2.5, 3.2, 2.9, 3.3, 3.5, 3.4, 
    3.6, 4.6, 4.7, 4.6, 4.5, 4.2, 4.1, 3.8, 3.6, 4.3, 4.2, 4.8, 5, 5.2, 5, 
    2.1, 0.9, 0, 0.2, 0.3, 0.9, 1.2, 1.5, 0.8, 1, 0.8, 0.4, 1.2, 1.6, 1, 0.5, 
    0.1, 0, 0, 0.1, 0.4, 0.9, 1.9, 1.7, 2.7, 2.4, 2.2, 3.9, 5, 5.4, 4.3, 3.9, 
    3, 2.8, 1.9, 5.7, 4.2, 5.5, 5.2, 5.8, 6.2, 5, 5.2, 5.3, 5.1, 6.6, 7.4, 
    7.2, 7.6, 8.1, 9.3, 7.9, 7.6, 7.6, 7.7, 7, 7, 6.8, 7.2, 7.7, 8.2, 8.1, 
    7.6, 7.7, 8.1, 8.9, 8.1, 9.8, 9.6, 8.9, 7.8, 8.1, 7.2, 5.8, 6.1, 6.9, 
    7.5, 7.4, 8.4, 7.3, 8.8, 8.2, 7.4, 7.9, 7.9, 8.5, 7.8, 7.5, 6.5, 6.8, 
    7.5, 7.9, 7.3, 7.9, 7, 7, 6.6, 6.9, 9.4, 9.6, 9.6, 10.1, 9.1, 8.2, 9, 
    8.9, 7.5, 8, 8, 10.4, 10.3, 8.4, 13.1, 11.9, 11.1, 9.8, 10.2, 9.8, 6.8, 
    10.5, 9.9, 11.6, 12.2, 12, 11.3, 10.7, 10.6, 10.5, 11, 12.1, 13, 13, 
    13.3, 15.3, 15.4, 14.1, 13.3, 14.3, 14.4, 14.2, 15.4, 12.9, 14, 16, 15, 
    14.6, 13.7, 13, 14.4, 13.5, 14.4, 14.4, 15.9, 12.1, 2.3, 0.5, 3.2, 1, 0, 
    0, 0, 1, 4, 3.7, 3.9, 7.2, 7.8, 7.7, 8.6, 9, 8.7, 9.8, 8.4, 9.1, 6.5, 
    7.3, 7.2, 7.6, 5.9, 4.3, 5.3, 5.7, 5.1, 4.9, 5.6, 4.6, 4.9, 4.4, 4.4, 
    3.7, 2.3, 2.6, 3.7, 2.4, 1.2, 1.2, 1, 1.5, 1.1, 0.5, 0.9, 2.4, 3.5, 4.1, 
    6, 8.5, 8.1, 6.8, 5, 5.9, 6, 6, 6.4, 5.8, 6.7, 7.3, 6.6, 7.4, 6.1, 8.5, 
    6.6, 7, 8.7, 10.1, 11.3, 10.6, 10.2, 8.7, 9, 9.9, 11.4, 11.7, 10.3, 9.1, 
    9, 10.2, 7.6, 5.6, 4.8, 6.2, 7.1, 8.4, 6.7, 7.7, 7.9, 6.7, 8.5, 9.2, 8.3, 
    5.8, 7.4, 4.4, 6.2, 5.9, 6.6, 7.9, 7.7, 8.3, 8.5, 8.2, 8.2, 8.2, 6.1, 
    4.4, 4.7, 4.8, 5.5, 5, 4.8, 3.2, 3.1, 0.6, 1.1, 0, 0.8, 1.4, 3.5, 5.1, 
    5.9, 6.3, 5.4, 5.8, 5.9, 6.3, 6.2, 6.2, 6, 4, 4.4, 3.8, 3.1, 3.1, 3.7, 
    3.9, 4.2, 3.8, 2.6, 3, 3.2, 1.1, 0.5, 3.6, 4.9, 6, 4.1, 3.7, 4.3, 5.1, 
    6.3, 8.2, 6.5, 4, 2.4, 3, 1.7, 3.7, 4.1, 4.9, 4.8, 4, 4, 6.7, 9.1, 7.5, 
    8, 9.2, 10, 9.4, 6.5, 5.6, 4.5, 4.8, 4.5, 3.9, 4.7, 4.6, 4.5, 4.8, 3.5, 
    4.1, 4.9, 4.8, 3.6, 4.2, 4.6, 2.7, 1.4, 2.6, 1.5, 2.7, 0.7, 0.9, 0.1, 
    0.1, 0.1, 0.3, 2, 2.3, 2.9, 2.1, 1.9, 0.3, 0, 0, 2.5, 0.6, 0.1, 0.1, 0, 
    0.9, 0.9, 0.3, 0.5, 1.6, 2, 3.2, 3.3, 3.3, 3.4, 4.7, 4.7, 5.6, 4.2, 3.5, 
    2.3, 2.9, 2.3, 3.5, 4.2, 6.5, 5.8, 5.7, 6.6, 6.1, 6.5, 7.2, 7.2, 7.7, 
    8.4, 8, 7.8, 7.2, 7.9, 7.1, 7, 6.6, 7.3, 7.9, 8.2, 8.5, 9.2, 9, 8.3, 8.1, 
    9.1, 9.6, 9.4, 10.1, 10.2, 10.7, 11.1, 9.9, 9.6, 10.3, 11.3, 11.4, 10.3, 
    11.2, 10.2, 8.6, 8.1, 7, 7.2, 6.6, 5.8, 4.5, 5, 2.8, 2.5, 1.5, 0.1, 0.6, 
    3.2, 3.4, 3.7, 3.3, 3.6, 1.8, 0.8, 2.5, 1.2, 0, 0, 2.5, 2, 2.7, 2.5, 1, 
    1.7, 3.9, 6.5, 6, 6, 5.3, 6.3, 5.4, 6.2, 6.4, 6.8, 7, 6.7, 7.4, 6.6, 8.2, 
    10.3, 13, 13.9, 11.1, 8.7, 8, 6.4, 5.2, 4.4, 5.1, 5.1, 4.9, 5.4, 4.6, 
    5.9, 6.3, 4.1, 5.3, 6, 6.4, 4, 2.7, 2.1, 3.4, 3.8, 5.4, 7.1, 7.7, 7.2, 
    7.2, 7.1, 6.9, 7.5, 7.4, 6.3, 6.1, 5.6, 6.6, 6.7, 6.2, 5.9, 4.2, 5.1, 
    5.5, 6.8, 6, 7, 8.4, 10.8, 11, 10.9, 10.8, 10.6, 11, 10, 8.6, 7.4, 5.5, 
    4.5, 1.9, 0, 0.2, 3.1, 4.8, 5.5, 5, 3.4, 2.1, 2.1, 2.2, 2.2, 2.3, 2.4, 
    2.4, 2.6, 2.5, 2.8, 2.7, 3.1, 3, 3.7, 3.7, 3.8, 4, 3.7, 3.7, 14.2, 14.6, 
    14, 12, 13.9, 12.5, 9.3, 6.5, 6.8, 7.3, 9.1, 7.4, 4.9, 4, 3.8, 5, 3.6, 
    2.4, 1.1, 2.1, 0.7, 0, 0.3, 0.9, 2, 2.6, 2.4, 4.1, 3.4, 5.4, 6.3, 6.3, 
    7.5, 8, 7.4, 7.4, 7.5, 6.5, 7, 7.3, 7.2, 7.6, 8.3, 8.3, 8.1, 8.1, 10.9, 
    10.1, 11.1, 9.6, 9, 9, 8.3, 7.8, 8.6, 8.9, 9.7, 10.7, 11.5, 11.1, 13.3, 
    12.9, 13.9, 13.4, 14.9, 15.7, 15.8, 15.4, 13.7, 13.6, 12.5, 14.3, 14, 
    12.8, 14.2, 9.2, 8.8, 8, 3.4, 2.7, 0.3, 0, 2.9, 3.4, 2.3, 1.9, 1.9, 2.1, 
    3.1, 0.2, 0.2, 5.1, 4.8, 3.6, 3.4, 5.4, 9, 9.8, 10.5, 8.4, 12, 11.9, 
    13.7, 14.2, 14.2, 14.5, 14.9, 13.4, 12.2, 11.6, 10.9, 11, 10, 10.3, 9, 
    8.3, 7.5, 6.6, 5.6, 3.3, 3.7, 2.2, 2.8, 0.8, 1.3, 4.6, 5.1, 4.7, 5.7, 
    5.1, 6.5, 6.9, 7.4, 7.8, 7.7, 8.5, 8.8, 9.3, 9.9, 9.4, 9, 9, 10.4, 11.1, 
    10.1, 11.9, 11.7, 10.5, 9.2, 5.9, 6.8, 6.2, 5.4, 4.3, 9.7, 9.2, 8.8, 6.3, 
    6.8, 6.8, 11, 10.6, 10.5, 8.7, 9.3, 11.7, 13, 14.2, 14.3, 14.5, 14.5, 
    15.1, 15.8, 15.5, 15.1, 15.1, 13.9, 13, 13.5, 15.6, 14, 13.4, 12.8, 13.9, 
    13.7, 13.9, 12.2, 10, 9, 8.3, 8.4, 7.6, 7, 7.2, 7.2, 5.9, 5.7, 7, 6.9, 
    6.7, 6.8, 5.8, 7.2, 6.1, 7, 8.2, 7.5, 7.1, 7.5, 7.9, 5.7, 5.2, 7, 8, 7.2, 
    7.2, 6.8, 8.2, 8.9, 10.5, 9.5, 9.5, 9.4, 8.5, 8.6, 8.3, 8.6, 8, 8.9, 8.8, 
    8.7, 8.9, 8.7, 7.8, 8.8, 8.8, 9.6, 8.5, 10.1, 9.4, 8.9, 9.4, 10.1, 9.8, 
    9, 9.6, 10, 9.5, 10.8, 10.8, 10.9, 11.1, 11.6, 11.4, 11.9, 11.1, 11.7, 
    11.1, 12, 11.9, 10.5, 10.4, 11.2, 12.8, 12.5, 11.8, 11.5, 11.2, 11.2, 
    11.7, 9.6, 9.3, 9.6, 9.1, 8.7, 10.8, 11.5, 9.9, 9.5, 9.9, 9.9, 9.4, 8.7, 
    9.9, 9.8, 12.8, 11.7, 11.1, 9.4, 8.6, 8.4, 6.7, 7.8, 9.4, 8.6, 9.2, 7.4, 
    8, 8, 7.1, 7, 8.4, 8.7, 9.1, 9.9, 9.1, 9.6, 10, 8.8, 10.3, 9.3, 7.9, 9.2, 
    7.8, 7.9, 8, 8, 9.1, 9, 7.9, 9.4, 3.9, 1.8, 0.7, 2.1, 3.6, 3.6, 2.4, 2.1, 
    1.7, 0, 0.1, 0.2, 1.2, 2.9, 0.6, 0.2, 1.3, 0.3, 0, 0, 0.2, 0.1, 0, 0, 0, 
    0, 0, 0.1, 0, 0.2, 0, 0, 0, 4.6, 0.7, 0.1, 0.1, 3.7, 7.3, 6.8, 7.2, 6, 
    6.9, 6.5, 6, 5.5, 5.6, 6.4, 6.4, 5.7, 6.5, 6.3, 6.5, 6.7, 6.9, 6.7, 7.7, 
    7.5, 7, 7.2, 7.4, 9.2, 10.3, 9.1, 9, 9, 9.3, 8.2, 8.5, 7.5, 6.7, 6.5, 
    7.3, 6.5, 6.2, 5.6, 5.2, 4.9, 3.6, 3.1, 2, 0.5, 1.1, 0.6, 0.3, 0, 0, 0, 
    0.2, 0.2, 0, 0.6, 3.6, 4.1, 5.9, 5.6, 6.5, 6.9, 5.9, 8.9, 10.6, 12.4, 
    12.7, 12.5, 11.9, 12.6, 11.8, 11.9, 9.7, 10.2, 9.6, 9.6, 8.6, 7.6, 6.8, 
    3.7, 3.7, 1.4, 0.9, 3.4, 1.3, 1.3, 0.4, 2.1, 2.7, 3.7, 5.2, 8.2, 12, 
    13.7, 15.5, 13.6, 13.1, 13.8, 13.9, 12.5, 12.3, 12, 12.6, 13.1, 10.9, 
    10.1, 8.7, 10, 8.4, 8.3, 7.2, 8, 7.8, 8.4, 7.8, 8, 7.7, 8.1, 7.3, 7, 7.4, 
    5.5, 4.4, 4.1, 3.6, 3, 2.9, 3.3, 3.3, 2.4, 2.3, 3.1, 2.6, 2.7, 2.3, 2.7, 
    2.6, 3.2, 3.5, 4.3, 6, 6.2, 6.2, 6.5, 6.3, 5.5, 4.8, 2.3, 1.2, 0.5, 0.4, 
    0.1, 1.2, 3.9, 5.4, 4.9, 5.6, 5.3, 5, 5.1, 4, 4.2, 5.1, 4.1, 4.3, 4.1, 
    4.2, 4.2, 4.1, 3.9, 4.8, 3.2, 2.6, 2, 1.5, _, _, _, _, _, _, _, 0.9, 2.8, 
    3.4, 4, 3.6, 3.8, 5.4, 5.6, 4.6, 4.7, 6.6, 5.6, 4, 2, 1.3, 1, 0, 0, 2.1, 
    3.4, 4.7, 5.2, 4.4, 4.2, 5.1, 5.8, 5.3, 6, 6.5, 4.9, 5.9, 6.5, 6, 6.7, 
    4.5, 4.1, 2, 2.7, 1, 2.2, 2.6, 1, 1, 4, 4.8, 4.4, 4.5, 4.6, 5.5, 7.1, 
    8.9, 8.9, 7.5, 7.5, 7.4, 8.1, 6.5, 6.5, 6.6, 6.4, 6.2, 7, 6.3, 5, 6.4, 
    4.9, 3.5, 3, 5.7, 4.7, 2.4, 1, 0.8, 0.6, 0.8, 0.3, 0, 1.2, 2.5, 2.3, 0.1, 
    2.7, 0, 4.1, 2.5, 3.8, 0.7, 0.3, 2.7, 4, 3.8, 3.7, 3, 2.5, 3, 0.6, 0, 
    2.8, 4.5, 5.5, 4.6, 4.4, 6.4, 3.5, 3.2, 3.4, 3, 2.8, 1.2, 2.2, 2.9, 3.3, 
    4.7, 4.6, 2.6, 2.5, 3.4, 5, 3.5, 4.1, 2.4, 2.3, 2.4, 0.2, 0, 0, 2, 0.9, 
    0.1, 0.6, 1.2, 1.3, 2.5, 3.5, 2.3, 2, 2, 0.1, 1.3, 0.9, 2.7, 2.4, 2.3, 
    0.7, 2.6, 2.6, 2.7, 2.4, 2.6, 2.4, 4, 3.5, 3.3, 3.6, 4.1, 2.4, 4.6, 4.6, 
    4.6, 5.7, 2.1, 1.9, 2, 0.8, 1.2, 1.7, 1.9, 2.5, 1.2, 4, 3.4, 3.3, 0.5, 2, 
    0.5, 1, 1.1, 0, 0, 0, 0, 2, 2.6, 3.6, 3.6, 2, 4.1, 4.6, 4.7, 3.6, 2.3, 
    3.4, 3.4, 4.4, 5.6, 5.6, 7.1, 7.5, 8.2, 7.4, 9.3, 8.6, 9, 9.2, 10.5, 9.7, 
    9, 8.7, 9.5, 9.3, 9.7, 10.4, 9.5, 8.6, 9, 10.4, 10.7, 9.1, 10.2, 8.9, 
    8.3, 6.2, 8, 9, 9.3, 9.1, 10, 10, 9.9, 10.4, 10.9, 11, 10.8, 10.7, 10.8, 
    10.6, 10.7, 10.9, 10.3, 10.1, 10.1, 10.2, 10.1, 9.2, 9.1, 9.2, 8.7, 9.3, 
    8.8, 7.8, 7.2, 5.9, 4.8, 6.5, 6.3, 6, 5, 4.4, 4, 4, 0, 1.1, 0.1, 0.1, 2, 
    0, 0, 3, 3.4, 3.4, 3.6, 4.7, 4.8, 5.5, 4.9, 5.4, 5.1, 5.8, 6, 9.1, 7.8, 
    8.1, 7.7, 8.1, 7.7, 6.5, 5.7, 6, 8.5, 8.1, 7.9, 7.9, 7.7, 5.5, 4.9, 5.8, 
    7.3, 7.7, 7.5, 5, 6.4, 6.4, 8.4, 6.3, 5.6, 4.1, 5.1, 4.4, 4.1, 3.3, 5, 
    6.4, 4, 2.7, 4.7, 6.2, 7.2, 6.7, 7.5, 7, 6.2, 4.2, 5.5, 7.6, 7.1, 5.4, 7, 
    7.1, 6.8, 6, 4.5, 3.5, 5, 7.4, 5.7, 5.3, 4.9, 4.8, 4.8, 4.3, 4.8, 4.8, 
    5.6, 6.7, 6.7, 6.1, 5.7, 5.7, 5.3, 5.3, 5.7, 6.5, 5.4, 5, 3, 1.4, 1.5, 
    2.6, 2.3, 3.4, 4.4, 6.3, 5.1, 5.6, 3.5, 4.8, 3.7, 4, 3.7, 3.2, 2, 1.7, 
    0.7, 1.9, 0.2, 0, 0.4, 1.2, 0.5, 0, 0, 0.2, 1.7, 1.7, 2.7, 1.4, 3.6, 3.8, 
    4.9, 5.1, 7.1, 8, 7.5, 10.7, 10.8, 10.1, 9.3, 6.4, 3.5, 3.2, 2.5, 0.9, 0, 
    2.2, 2.9, 2.6, 1, 0, 1.2, 1.3, 2.1, 2.7, 3.6, 4.3, 4.5, 3.9, 3, 3.1, 1.3, 
    1.2, 1.1, 1.2, 2.3, 1.4, 0.2, 0, 0, 0.3, 3.3, 0.2, 0.4, 0, 0, 0.5, 1.5, 
    2, 5.5, 5.2, 5.6, 5.8, 5.7, 5.8, 5.1, 4.7, 4.1, 2.7, 3, 3.3, 3.9, 3.1, 3, 
    2.8, 2.6, 2.5, 1.5, 1.9, 2.1, 2.5, 2.6, 2.6, 2.6, 2.8, 2.5, 4, 3.7, 3.6, 
    3.4, 4.2, 3.1, 4.1, 3.9, 4.4, 4.1, 5.5, 5.9, 6.2, 6.2, 7.1, 8.7, 7.7, 
    8.2, 9.2, 9.4, 9.8, 10.2, 9, 7.8, 10.2, 11.6, 11.9, 11.6, 11.7, 10.9, 
    10.2, 9, 7.8, 9.2, 9.5, 9.7, 8.7, 7.6, 9.5, 12.8, 12.7, 11.4, 10, 11, 
    11.1, 12.5, 12.9, 12.8, 14.2, 13.9, 12.2, 13.4, 14, 16.2, 15.7, 13.7, 
    12.7, 12.1, 11.5, 10.8, 11, 10.6, 12.6, 12.2, 12.5, 13.4, 14.1, 14.5, 
    13.2, 12.5, 11.7, 12, 12.4, 12.2, 12.9, 13.9, 13.5, 13.9, 14, 13.8, 12.9, 
    12.8, 14.2, 12.3, 13.8, 14.5, 14.6, 14.6, 15, 15.8, 15.9, 15.9, 15.1, 
    14.6, 13.6, 12.8, 12.3, 12.5, 11.5, 12, 10.7, 10.9, 12.1, 12, 11.7, 11.5, 
    11.9, 11.2, 10.7, 10.2, 9.4, 10, 9.4, 10.1, 11.9, 12.7, 12.5, 13.8, 13.5, 
    13, 12.2, 12.5, 12.6, 11.4, 10.7, 10.3, 9.9, 9.9, 9.6, 8.2, 8.4, 8.7, 
    9.3, 8.3, 8.4, 8, 7.1, 6.8, 5.9, 6.4, 5.2, 6.2, 7.2, 7.3, 8.4, 7.5, 8.2, 
    6.7, 8.1, 8.6, 9.7, 9.1, 7, 7.5, 5.9, 6.8, 3.6, 8.5, 6.4, 4.1, 4.2, 3.5, 
    3.8, 1.7, 3.2, 2.6, 1.4, 2.1, 2.7, 1.4, 3.1, 2.7, 4.4, 1.3, 1.9, 3.2, 
    2.3, 1.9, 2.9, 0.4, 0.4, 2.6, 4.4, 3.5, 3.5, 3.2, 3.2, 0.7, 3.7, 3.5, 
    4.9, 3.4, 5.4, 4.5, 1.4, 3.5, 4.9, 3.1, 2.4, 4.3, 0.6, 0.4, 4.8, 2.2, 1, 
    1.1, 1.4, 1.3, 2.9, 0, 2.8, 3.9, 3.6, 4.4, 4.1, 4.8, 5.5, 5, 5.6, 5.9, 
    6.3, 6.9, 6.7, 7.3, 6.3, 7.1, 7.5, 7.3, 7.4, 7.9, 8, 8.5, 9.5, 7.8, 7, 
    6.7, 6.1, 5.7, 5.3, 6.2, 7.3, 7.8, 8.7, 7.7, 6.7, 4.5, 3.4, 1.9, 1.9, 
    2.2, 4.4, 5.8, 5.2, 3.9, 2.5, 2.5, 2.5, 0.1, 1.4, 2.7, 3.3, 3.3, 4.8, 5, 
    5.9, 6, 7.7, 7.8, 11.1, 11.6, 12, 12.1, 11.9, 11.8, 12.9, 14, 13, 12.6, 
    12.3, 12, 10.5, 11.3, 11.4, 11.2, 11.4, 10.1, 10, 8.9, 9.1, 8, 8, 9.6, 9, 
    6.8, 7.2, 7.3, 6.9, 4.6, 5, 4.8, 4, 4.1, 4.3, 5.1, 3.7, 3.4, 5, 4, 4.8, 
    4.8, 5.4, 4.4, 4.8, 4.1, 4.1, 4.5, 2.5, 1.3, 4.1, 2.3, 2.2, 0.9, 1.6, 2, 
    2.4, 2, 4, 4.1, 6.6, 7.1, 7, 7, 6.7, 7.9, 4.4, 7, 7.5, 7, 7.3, 7.6, 7.5, 
    8.9, 8.6, 8.8, 9.7, 10, 10.5, 11, 11.3, 11.3, 12.4, 11.6, 11.9, 12.7, 
    10.9, 10.7, 14.4, 11.8, 9.6, 10.6, 11.7, 11.5, 11.3, 10.1, 10.4, 15, 
    16.5, 15.5, 13.9, 14, 15.9, 16.7, 15.6, 16.1, 17.5, 18.6, 18.4, 20.2, 23, 
    20.7, 20.8, 20.9, 21.5, 23.6, 23.1, 22.9, 21.7, 22.1, 22.5, 21.1, 21.1, 
    21.8, 21.3, 20.8, 21.8, 21.8, 21.2, 21, 20.7, 20.5, 20.3, 17.2, 17.7, 
    15.3, 15.4, 14, 10.7, 10.4, 14.1, 15.3, 15.2, 15.7, 15.3, 13.8, 14.7, 15, 
    14.8, 14.9, 14.4, 14.2, 13.3, 13.2, 14, 14.4, 14.1, 14.4, 14.4, 13, 12, 
    13, 13.8, 11.6, 12.9, 12.4, 13.5, 13.8, 13.7, 12.4, 13.1, 7.5, 6.2, 5.1, 
    5.3, 1.3, 7.6, 7.1, 7, 4.9, 6.7, 4, 6.9, 6.6, 6, 4.9, 5.6, 4, 2.5, 3, 
    3.2, 2.7, 2.2, 3.2, 2.1, 0.8, 4.5, 7.2, 7.9, 8.3, 7.8, 8.4, 6.6, 5, 1.6, 
    3, 3.5, 5.2, 3.4, 1.7, 1.8, 1.3, 1.2, 2, 1.5, 1.4, 1.8, 1.4, 0.3, 0.5, 
    0.3, 1, 0.3, 0.3, 0.3, 0.9, 1.3, 0.8, 0.4, 0.6, 0.7, 0.8, 0.6, 0.6, 0.7, 
    1.8, 0.8, 0.9, 0, 5.3, 5.5, 9.1, 11.1, 8.7, 8.2, 7.1, 8.2, 8.8, 8, 8.5, 
    8.7, 8.1, 8.3, 10.2, 6.7, 12.5, 11.7, 12.7, 11.4, 14.8, 15.5, 17, 18.7, 
    17.5, 17.5, 17.6, 16.9, 16.4, 16.6, 16.9, 15.9, 16.5, 16.4, 15.2, 12.1, 
    14.4, 14.5, 10.9, 8.8, 8.1, 6.6, 7.8, 8.9, 9.3, 5.5, 6.7, 9.3, 9.8, 10.7, 
    12, 15, 15.1, 15.4, 12.5, 2, 5, 2.6, 4.8, 4.4, 4.5, 1.4, 0.2, 1.3, 4.4, 
    0, 6.4, 5, 5.6, 4.5, 4.2, 6.1, 4.3, 0.5, 0, 4.5, 3.5, 4.3, 4.6, 3, 2.6, 
    3.2, 3, 3.6, 2.2, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0.8, 0.1, 1, 1.3, 0.3, 
    1, 2.4, 1.7, 1.6, 2.2, 0, 0, 0.6, 2, 3.3, 6.9, 5, 6.8, 5, 5.7, 7.9, 8, 
    6.1, 5.2, 6.7, 5.8, 5.3, 5.8, 6.5, 6, 4.7, 2.7, 0.8, 0.7, 0.7, 0.5, 2.3, 
    4.1, 4, 3.9, 3.2, 4.4, 6.3, 5.8, 6.6, 5.9, 6.1, 8.3, 9.1, 9.2, 8.3, 7.1, 
    9.2, 7.5, 5.7, 5.1, 6.8, 9.7, 9.6, 9.6, 9.9, 9.7, 9.4, 9.4, 9.7, 9.5, 
    9.6, 9.6, 9.6, 10.3, 9.8, 8.9, 10, 9.7, 6, 9.1, 10.7, 12, 12.1, 11, 10.5, 
    11.2, 12.1, 13.3, 17.4, 19.2, 16.7, 15, 13.2, 14, 16.2, 19.8, 19.2, 21, 
    18, 13.2, 9.8, 11, 9.5, 9.9, 9.2, 12.4, 15.1, 12.8, 11, 12.1, 12.4, 10.1, 
    11.5, 14.3, 14.1, 17.1, 15.4, 13.4, 13.1, 11.3, 11.3, 10.5, 10.8, 13.1, 
    14.9, 14.9, 14.9, 12.3, 13.4, 18.2, 18.4, 21.4, 18.2, 14.7, 14.5, 14.3, 
    13.6, 13.4, 14.5, 18.3, 17.2, 14.2, 13.1, 10.8, 11, 11.9, 10.6, 11.5, 
    11.9, 11.5, 11.3, 11, 10, 10, 11.3, 10.2, 9.1, 8.6, 8.3, 7.2, 7.6, 6.6, 
    7.7, 8.4, 8.3, 8.3, 6.7, 9, 9.6, 10.3, 10.5, 9.3, 7.9, 8.2, 7.4, 8.7, 
    7.7, 5.4, 4.9, 4, 6.1, 7.4, 6.4, 9.3, 8.7, 8.1, 8.5, 8.8, 7.8, 6.4, 6.6, 
    6.4, 7.6, 6.9, 7, 8.7, 11.2, 10.5, 11.5, 12.3, 13, 11.5, 10.9, 11.8, 
    13.4, 12.2, 12.2, 12.3, 10.8, 7, 10.6, 9, 8.2, 6.1, 9, 7.2, 7, 5.9, 8.8, 
    7, 7.4, 7.5, 10.8, 11.8, 12.6, 4.8, 2.2, 3.5, 5.8, 5, 0.9, 6.7, 5.5, 7.5, 
    5.7, 2.7, 4.3, 4, 7.2, 5.7, 6.4, 8.2, 9.1, 9, 10.1, 6.6, 12.3, 10.6, 9.1, 
    8.7, 7.6, 6.4, 7.3, 5.9, 6.8, 6.9, 6.5, 5.4, 7, 7.1, 8.8, 9.5, 11.1, 9.2, 
    10.8, 12.4, 13.5, 16.9, 12.8, 9.6, 7.5, 7.8, 9, 9, 8.9, 8.5, 7.8, 7.4, 
    8.5, 7.7, 8.6, 6.9, 7.3, 10.1, 8.2, 7.6, 7.7, 7.5, 7.3, 7.3, 8.5, 10.1, 
    7.9, 6.3, 7.2, 5.2, 7.2, 10.5, 7.6, 7.9, 7.3, 7.8, 7.5, 8.7, 8.7, 9.4, 
    10.5, 11, 11.6, 11.7, 10.9, 10, 9.6, 8.3, 8.7, 8.6, 6.6, 8.3, 8.4, 6.2, 
    9, 9, 10, 7.8, 12.2, 13.5, 15, 16.4, 14, 13.3, 13.3, 13.9, 10.3, 9.9, 
    10.2, 8.6, 8.9, 8.1, 8.1, 9.4, 9, 8.7, 7.8, 10.1, 10.5, 10.5, 10.7, 9.4, 
    10.4, 9.3, 9.1, 8.3, 10.4, 11.8, 11.6, 10.5, 10.2, 10, 10.7, 13.3, 14.1, 
    12.4, 8.4, 6.3, 8.7, 8.5, 4.8, 6.4, 10, 10.5, 11.3, 11.3, 10.5, 13, 12.8, 
    9.6, 8.3, 4.4, 1.2, 3.8, 3.8, 6.4, 7.2, 8.2, 7.7, 8.3, 7.9, 7.1, 9.8, 
    9.6, 7.8, 8.6, 7.7, 7.7, 7.7, 9.6, 11.5, 11.1, 10.4, 9, 8.2, 8.5, 5.4, 
    4.3, 3.3, 3.3, 4, 2.7, 3.3, 2.9, 3.9, 3.7, 2.2, 3.9, 1.3, 1.9, 2, 4, 2.7, 
    2.3, 3.8, 3.9, 1.8, 3, 2.2, 2.5, 2.2, 3.7, 2.5, 2.4, 2.6, 2.8, 3.3, 3.4, 
    2.9, 3.4, 2, 1.9, 2.1, 1.6, 1.3, 2.3, 1.7, 2.1, 2.8, 3.2, 2.1, 2.8, 3, 
    1.3, 2.1, 2.3, 1.4, 3.5, 2.1, 4, 2.6, 4.5, 3.3, 2.6, 1.8, 3.2, 3.1, 2.9, 
    3.4, 3.6, 4.3, 4.5, 2.8, 2.2, 2, 2, 2.2, 0.5, 4.7, 2.5, 1.8, 1.9, 3, 3.6, 
    4, 4.1, 4.2, 5.1, 4.8, 3.8, 3.9, 4, 4, 7.5, 7.7, 6.1, 5.8, 6.4, 3.6, 7.3, 
    6.9, 8, 6.6, 8.8, 6.9, 8.3, 7.8, 6.4, 4.7, 3.5, 7.2, 10.9, 9.4, 12.1, 
    14.1, 13, 10.4, 9.4, 10, 8.8, 8.9, 7.2, 7.9, 8.5, 7, 5.9, 8.8, 11.3, 
    13.5, 15.9, 15.3, 9.5, 10.1, 11.3, 11.3, 11.1, 11.1, 8.3, 9.2, 10.8, 
    11.7, 10, 8.6, 10.3, 11.2, 7.3, 8.7, 7.9, 6.7, 5.8, 6.9, 7.9, 1.9, 3.1, 
    2.6, 2.4, 1.4, 1.5, 3.2, 7.6, 5.7, 6.7, 8.4, 8, 6.1, 3.8, 2.8, 1.3, 2.5, 
    0.8, 1.2, 0.2, 7.2, 6.9, 6.3, 8.5, 10.4, 11.8, 12.5, 11.5, 12, 11.4, 11, 
    11.7, 11.4, 12.2, 11.3, 11.6, 11.5, 11, 9.5, 9.3, 9.1, 8.3, 9.5, 9.8, 
    10.2, 12.5, 13.4, 14.8, 17.8, 21.2, 21.8, 24.1, 23.7, 24.7, 23.7, 19, 
    9.1, 8, 8, 6.9, 8.5, 11.9, 11.9, 13.5, 13.9, 14, 13.9, 14.4, 15.1, 15.3, 
    14.8, 13.6, 13.1, 13.5, 13.9, 15.4, 16.2, 16, 15.4, 15.5, 16.4, 16.9, 
    17.1, 17.6, 17.6, 17.9, 17.5, 17.2, 16.7, 18, 16.9, 16.2, 16.1, 15, 14.3, 
    14.2, 14.7, 14.2, 14.4, 15.1, 15.8, 17.8, 17.7, 18.7, 18.5, 15.9, 14.4, 
    12.6, 11.4, 11.9, 10, 9.5, 8.5, 9.5, 11.2, 11.4, 13.5, 14.3, 15.3, 14.5, 
    15.4, 15.6, 15.3, 15.1, 13.7, 13.9, 11.4, 10.8, 10.1, 9.9, 9.8, 8.6, 7.3, 
    6.9, 6.1, 7.4, 6.6, 8.1, 6.2, 7.6, 8.3, 7.7, 8.6, 8.6, 8.7, 10.8, 9.9, 
    10, 12.7, 10.5, 10.2, 8.7, 9.2, 12.7, 7.1, 10.1, 10.5, 11.5, 11.9, 13.4, 
    17.1, 15.7, 17.6, 16.2, 15.6, 15.4, 11.7, 10.8, 14.7, 11.9, 11.1, 11.4, 
    11.3, 12.2, 13.1, 12.7, 12.4, 12.3, 13.8, 12.7, 14.2, 13.5, 10, 12.4, 
    13.1, 13.9, 12.1, 12.8, 9.9, 9.1, 10, 7.6, 8.4, 8.4, 8, 7.8, 11.7, 14.6, 
    14, 15.1, 11.9, 9.2, 9.6, 9.1, 10.3, 13, 12.6, 12.9, 13.5, 13.5, 12, 13, 
    12.1, 11.8, 11.8, 11.9, 13.1, 14.2, 11.5, 8.4, 10.7, 9, 9, 8.7, 10.3, 
    10.2, 10.2, 11.7, 9.4, 12, 11, 11.1, 10.4, 10.4, 8.9, 8, 7.9, 7, 5.3, 
    6.7, 7.6, 5.9, 7.8, 8.4, 7.9, 7.9, 8.7, 7.9, 9.6, 9.3, 9, 7.7, 7.9, 7.5, 
    9.1, 9.2, 10.3, 9, 9.6, 10.6, 10.3, 7.7, 6, 5.9, 6.3, 7.4, 7.8, 9.1, 9.1, 
    9.2, 10, 11.1, 10.5, 10.2, 10.2, 9.8, 9.6, 10.1, 9.3, 9.8, 10.6, 11.9, 
    11.9, 12.9, 10, 12.5, 13.7, 12.5, 10.5, 11.2, 11, 11.2, 11.4, 12, 12.5, 
    10.6, 11.2, 10.6, 10.6, 10.8, 11.6, 11.1, 11.2, 11.4, 13.5, 11.8, 12.1, 
    12, 11.6, 10.2, 10.1, 9.6, 8.8, 10.8, 11.6, 10.6, 10, 11.6, 13.4, 12, 
    13.4, 13.5, 14.6, 16.5, 7.8, 17.1, 14, 9.6, 20.3, 18.2, 17.3, 16.5, 17.4, 
    12, 13.9, 14.9, 14.6, 13.8, 11.1, 10, 9, 7.8, 8.2, 7.4, 8.2, 8.7, 8.4, 
    9.1, 7.3, 8.5, 9.8, 8.7, 15.7, 18.8, 18.4, 18.3, 19.2, 19, 18.3, 20.6, 
    16.5, 4.9, 2.4, 5, 4, 4.7, 6.1, 7.4, 10.2, 12.5, 12.8, 13.9, 14.8, 16.2, 
    13.4, 14.2, 15.1, 15.9, 15.7, 14.2, 14.7, 3, 2.2, 1.6, 3.8, 3.4, 3.4, 
    3.8, 13.4, 13.6, 3.7, 5.3, 3.3, 4.7, 2.8, 17.3, 19.1, 20.2, 20.3, 18.8, 
    17.4, 14.8, 15.8, 15.2, 15.5, 13.9, 14, 13.8, 14.2, 13.9, 14.4, 14.1, 
    14.1, 13.1, 12.7, 13.2, 12, 9.9, 9.9, 11.4, 12.4, 11.6, 12.6, 13, 12.4, 
    12, 11.7, 12, 11.9, 12.2, 12.6, 11, 11.1, 10.8, 11.3, 12.2, 12.5, 14.5, 
    14.5, 15.4, 16, 17.1, 15.7, 14.7, 13.7, 12.3, 11.6, 11.2, 10.1, 9.1, 8.2, 
    8, 9.2, 9.4, 11, 10.3, 10.3, 10, 9, 9.9, 9.8, 8.9, 8.3, 7.9, 7.1, 2.4, 3, 
    3.5, 3.9, 5.7, 4.9, 3.5, 3.5, 3.6, 4, 5.2, 6.5, 6.7, 7, 7.9, 8.3, 7.4, 
    8.1, 7.5, 8.2, 8.3, 10.3, 11.4, 14.1, 15, 14.5, 16.1, 15.5, 16.6, 18, 19, 
    19.9, 20.2, 21.4, 22.3, 22.9, 24.5, 26.3, 26.8, 24.8, 18.3, 14.1, 14, 
    13.4, 13.7, 14.9, 16, 17, 16.4, 14, 12.4, 11.8, 11.5, 11.2, 12.3, 12.5, 
    14.1, 13.1, 9.1, 7.8, 8, 8.5, 9.4, 9.4, 10.5, 13, 11, 9.5, 6.3, 7.2, 7.9, 
    8.3, 9.7, 11.6, 11.4, 13.5, 11.9, 8.7, 8.7, 8.5, 8.2, 7.6, 7.2, 7.3, 8.5, 
    7.3, 6.9, 9.3, 8.8, 8.9, 10.5, 9.1, 16.1, 14.7, 12.8, 12.2, 12.5, 11.2, 
    13.1, 12.4, 11.3, 8.9, 11, 10.1, 13.4, 10.6, 11.4, 11, 12.3, 10.6, 12.5, 
    13.3, 12.3, 11.4, 11.5, 12, 10.8, 9.9, 9.5, 7.2, 5.1, 0.5, 0.5, 0.9, 1.7, 
    0, 5.6, 4.3, 3.9, 2.1, 2.1, 2.4, 3.7, 0.8, 1.1, 6.4, 9.1, 7.9, 8.3, 7.6, 
    8.8, 10.2, 14.4, 10.5, 11.9, 11.7, 14.6, 16, 14, 16, 14.4, 13.9, 10.2, 
    10.2, 5.8, 10, 8.3, 6.4, 2.7, 5.4, 0.9, 1.9, 5.4, 10.1, 9.8, 11.4, 9.6, 
    9.7, 10.2, 9.7, 9.7, 8.9, 9, 9.6, 11.1, 10.4, 13.9, 15.1, 9.6, 14.4, 
    12.9, 10.4, 10.6, 13.2, 13.3, 15.8, 18.5, 21.3, 16.4, 17.1, 14.3, 14.1, 
    15, 12.7, 11.9, 13.3, 12.4, 11.3, 12.9, 14.3, 14.8, 14.2, 14, 13.8, 14, 
    11.6, 12.7, 13.2, 13.2, 12.9, 11.8, 12.4, 10.7, 12.6, 15.4, 14.4, 10.4, 
    8.3, 5.9, 3.7, 2.2, 2.2, 6.8, 11, 12.5, 13.3, 13.8, 11.9, 7.3, 5.9, 4.3, 
    5.3, 0.7, 0.3, 2.1, 5.5, 4.9, 5.3, 5.7, 4.6, 4, 4.2, 6.9, 7.8, 8.1, 6.9, 
    6.8, 5, 10.8, 12.2, 10.6, 10.9, 7.8, 9.2, 9.6, 11.6, 14.5, 14.2, 14.3, 
    16.4, 18.2, 19.8, 21.4, 21.7, 19.7, 20.2, 21.4, 21.3, 22.4, 22.5, 22.2, 
    19.6, 18.8, 19.3, 16.5, 16.5, 14.6, 14.3, 16, 14.8, 12.4, 11, 10.4, 9.8, 
    12.6, 9.9, 9.8, 8.9, 8.4, 9, 8.1, 9.2, 8.8, 8.4, 9.1, 7.7, 8.7, 8.8, 9.6, 
    8.5, 7.9, 7.9, 7.9, 7.4, 8.3, 7.8, 7.4, 8.7, 8.1, 6.6, 6.5, 6.3, 4, 5.7, 
    7.3, 7.3, 9.2, 9.4, 9.1, 9.6, 4.2, 1, 1, 2.6, 4.6, 0.3, 0.5, 0, 0.5, 1.9, 
    0.6, 1.1, 1.1, 0.3, 7.3, 8.5, 6.8, 6.9, 5.4, 1.6, 0.5, 0.1, 0.7, 0.2, 
    0.8, 0.9, 1.4, 1.2, 1.1, 1.4, 1, 0.3, 0.4, 1, 6.7, 7, 8.4, 9, 10.1, 10.7, 
    11.2, 10.9, 11.4, 12.3, 13.2, 11.9, 11.1, 13, 12.6, 12.5, 15, 15.5, 15.6, 
    14.7, 13.8, 14.7, 14.5, 14.5, 15, 15.4, 14.8, 15.6, 15.2, 14.6, 14.2, 
    13.9, 13.7, 12.8, 12, 12.7, 12.7, 11.8, 10, 10.8, 10.6, 8.8, 6.6, 7.1, 
    8.4, 6.6, 6.7, 7.7, 6.6, 8.3, 8.3, 6.4, 7.2, 7.2, 8.4, 7.3, 9.1, 7.8, 
    7.1, 6.7, 7.1, 7.5, 6.2, 6.9, 5.1, 3.9, 5.7, 5.4, 5.1, 5, 4.4, 4.7, 4.3, 
    4.9, 4.8, 5.8, 5.4, 6.8, 6.7, 4.7, 6.5, 5.9, 3.6, 2.2, 2.1, 1.4, 0, 0, 0, 
    0.8, 2.7, 2.6, 13, 16.6, 17.9, 17.1, 20, 18.3, 17.1, 16.6, 15.1, 13.2, 
    11.3, 9.1, 7.8, 10, 10, 10.2, 10.1, 9.9, 9.7, 6.8, 6.6, 5.2, 3.6, 2.8, 
    9.3, 8.6, 8.9, 10, 9.2, 10.3, 9.9, 7.8, 7.9, 6.8, 7.3, 7.8, 8, 11.6, 
    13.2, 14.4, 15, 13.4, 11.4, 11.7, 12.2, 10.6, 9.1, 10.3, 10.1, 9, 8.3, 6, 
    5.7, 6.8, 5.8, 6.7, 6.8, 5.2, 5.1, 5.3, 5.4, 4.9, 4.6, 3.9, 2.8, 0.7, 
    1.8, 3, 3, 3.8, 3.3, 4.4, 3.8, 4.5, 4.6, 5.5, 5.6, 4.7, 5, 4.2, 4.6, 4.1, 
    3, 3.5, 5.4, 3.8, 5.2, 6.1, 7.2, 8.4, 8, 8.8, 8.1, 9, 9.4, 8.9, 10.1, 9, 
    6.7, 6.8, 7.3, 6.9, 5, 5.4, 5.8, 5.4, 5.3, 5.7, 5, 7.1, 4.6, 6.5, 4.8, 
    3.8, 4.6, 3.3, 2.3, 3.1, 2.3, 1.6, 0.6, 1.2, 0.6, 1.1, 0.6, 0, 1, 0.3, 
    4.6, 3.2, 5, 6.2, 5.4, 4.3, 1.6, 0.5, 1.1, 0.2, 1.3, 1.3, 1.9, 0.4, 0.2, 
    0.1, 0.9, 1.3, 0, 0.6, 0, 0, 5.4, 8.1, 12.5, 13, 13.6, 12.5, 10.2, 8.7, 
    3.8, 2.3, 0.5, 0.3, 4.6, 4.3, 4.2, 0.7, 1.1, 7.9, 8, 9, 12.4, 11.1, 10.7, 
    10.4, 9.1, 8.6, 9, 9.1, 7.5, 7.7, 7.8, 6.2, 3.6, 2.7, 4.2, 5.3, 3.7, 6.5, 
    7.9, 6.4, 1.8, 3, 1.3, 3.8, 2.8, 3.7, 3.5, 4.6, 4.1, 6.7, 7.5, 9.7, 4.3, 
    2.4, 3.3, 5.6, 0.6, 6.1, 6.2, 4.7, 3.8, 3.6, 2.7, 2.4, 2.5, 0.8, 1.9, 
    3.9, 6.7, 10, 10, 11.8, 12.4, 11.6, 9.7, 9.1, 10.5, 9.1, 9.2, 9.5, 12.1, 
    11.9, 10.6, 10.2, 9.7, 9.7, 8.6, 10.3, 10.1, 9.1, 8.8, 7.6, 8.1, 8.1, 
    8.4, 11.2, 9.7, 6.9, 7.2, 11.5, 11.4, 11.2, 11.8, 13.5, 15.4, 15.6, 15.6, 
    15.5, 15.5, 15.5, 15.6, 15, 14.4, 14.7, 15.5, 14, 12.9, 14.2, 14.2, 14.5, 
    14.3, 14.7, 14.2, 15.9, 16.1, 15.5, 16.7, 16, 15.7, 15.3, 16.2, 16.6, 
    17.9, 17.6, 17.8, 17.3, 17.7, 17.7, 15.5, 13.4, 12, 10.5, 11, 11.4, 13.9, 
    15.5, 14.3, 15, 14.7, 14.4, 16.1, 13.3, 13.9, 12.8, 13.3, 11.8, 11.6, 
    9.8, 8.5, 7.3, 8.2, 8.9, 9.6, 10, 9.9, 11.4, 12, 12.7, 11.7, 11.9, 11.5, 
    11.2, 11.8, 9.3, 8.9, 8.5, 10, 10.2, 11.2, 9.6, 9.6, 8.8, 10.3, 10, 10.1, 
    10.5, 11.2, 11.9, 12.4, 12.6, 15, 15.9, 10.4, 9.8, 9.4, 9.1, 9.8, 9.2, 
    8.7, 8.5, 9.7, 12.5, 13.9, 14.1, 12.9, 12.7, 8.8, 7.8, 9.4, 5.7, 6.2, 
    5.6, 5.9, 6, 6.8, 4.9, 5.7, 5.7, 6.2, 8.8, 8.8, 7.5, 7.1, 5.7, 5.3, 4.2, 
    5.3, 6.4, 7.7, 7.6, 9.7, 9.7, 10.3, 9.7, 10.4, 9.5, 9.4, 9.7, 10.9, 11.4, 
    10.9, 10.5, 9.2, 9.1, 9.2, 9.3, 9.5, 10.1, 10.4, 10.8, 11.5, 12.1, 10.5, 
    11.2, 11.2, 11.2, 10.3, 10.3, 10.6, 9.6, 8.9, 8.2, 8.1, 8.8, 10.5, 9.9, 
    10.4, 10.5, 9.3, 8.8, 9.2, 8.5, 9.2, 8.9, 9, 8.9, 9.3, 9.6, 10.6, 10.1, 
    11, 12, 10.7, 9.6, 9.8, 10.7, 10.5, 10.3, 11.1, 10.6, 10.4, 7.6, 8.2, 
    9.3, 9.1, 9.5, 9, 7.4, 6.1, 7.8, 7.8, 7.3, 7.7, 7.7, 1.3, 6.7, 7.8, 8.1, 
    9.5, 9.1, 8.7, 10.5, 11.4, 12.7, 12.2, 12.6, 12.7, 13.2, 12.4, 11.6, 9.8, 
    8, 2.2, 3.3, 3.6, 8.5, 11.2, 12, 10.8, 13.2, 9.3, 11.8, 10.1, 9.6, 9, 
    8.2, 9.1, 9, 10.5, 11.7, 11.3, 10.8, 10.5, 10.1, 14.1, 13.9, 13.3, 11.2, 
    11.4, 9.9, 9.6, 8.6, 9.4, 9.3, 9.6, 7.5, 6.6, 6.1, 4.4, 2.8, 1.8, 3.5, 
    2.9, 6.3, 9.4, 7.5, 7.8, 9.6, 3.6, 0.3, 2, 3.7, 3.1, 4.3, 3.1, 4.4, 2.4, 
    3.6, 2.4, 1.8, 1.2, 1, 0.9, 0.9, 5.5, 3.9, 5.2, 4.3, 3.1, 1.8, 1.3, 1.6, 
    0.7, 0.6, 1.2, 1.2, 1.2, 1.8, 4.1, 1.4, 4.4, 1.5, 2.5, 1.7, 3, 2.9, 1.1, 
    0.6, 3.1, 3.4, 0.1, 1, 1, 0.7, 0.4, 1.2, 1.3, 2, 2.7, 1, 2, 1.3, 0.1, 
    0.4, 0.5, 1.4, 1.8, 2.6, 1.1, 0.6, 1.4, 0.4, 1.6, 0, 1.5, 2.7, 5.3, 4, 
    3.7, 5, 2.6, 1.9, 2, 1.1, 0, 0.4, 5.1, 5.3, 4.3, 3.1, 1.4, 3.7, 4.1, 0.3, 
    0.2, 0.5, 3.8, 3.2, 1.1, 0.7, 0.7, 1.4, 0, 0.9, 1.5, 0.8, 0.1, 1.1, 1.1, 
    0.4, 1.6, 1.2, 0.9, 1.1, 2.6, 2.1, 0.7, 2.9, 1.7, 1.7, 1.5, 2.7, 1.3, 
    1.3, 1, 1, 1.3, 1.2, 0.6, 1.5, 3.5, 3.6, 3.1, 2.9, 3.6, 3.8, 4.5, 4.2, 
    4.1, 3.5, 4.3, 5.2, 5.5, 6.2, 6.7, 7.4, 7.2, 8.3, 8.9, 9.4, 9.6, 9.6, 
    9.6, 9.3, 8.4, 8.3, 7.9, 7.8, 6.9, 5.9, 6.3, 6.5, 7.9, 8, 8.9, 8.7, 10.1, 
    11.3, 11.1, 11, 10.9, 11, 11.5, 10.9, 12.6, 11.9, 11.8, 11.1, 10.4, 11.2, 
    10.5, 11.3, 11.4, 11.3, 12.3, 12.4, 13.3, 12.7, 12.4, 12.6, 11.7, 11.3, 
    11.1, 14.1, 14.1, 13.7, 14.2, 14, 15.3, 12.7, 11.5, 9.3, 11, 12.8, 15.7, 
    18.7, 16.6, 18.7, 19.4, 20.4, 23, 20.8, 18.9, 15.4, 14.3, 13.2, 12.6, 
    13.6, 14.2, 12.4, 13, 12, 10.8, 7.1, 7.3, 11, 10.5, 9.6, 7.9, 9, 7.6, 
    5.4, 7.5, 7.5, 6.8, 8.1, 10.3, 10, 8.9, 10.8, 8.6, 6.5, 4.6, 2.8, 2.4, 
    0.1, 3.3, 5.7, 6.2, 9.3, 8.6, 6.4, 1.8, 3.2, 2.9, 4.5, 2.2, 1.4, 3.7, 
    4.1, 4.9, 5.6, 10.3, 11.6, 14.1, 9.8, 13.6, 18.4, 13.6, 11.3, 11.8, 13, 
    13.4, 11.6, 8, 7.9, 7.3, 6.8, 6.9, 5.3, 5, 4.6, 4.6, 3.8, 3.5, 3.5, 2.1, 
    3, 1.2, _, _, _, _, _, _, 3.6, _, _, _, _, _, _, 6.5, _, _, _, _, _, _, 
    _, _, _, 4.6, _, _, _, _, _, _, 6.5, _, _, _, 5.4, _, _, _, _, _, _, _, 
    _, _, 11.1, 10.7, 10.2, 11.3, 12, 12.3, 12.8, 13.8, 14.8, 15, 15.2, 14.5, 
    14.4, 14.6, 15.2, 16.2, 15.4, 16.9, 16.6, 14.4, 12.6, 10.1, 9.8, 10.9, 
    10.7, 9.9, 9.5, 10.3, 9.1, 8.2, 7.6, 7.6, 7.5, 6, 5, 4.7, 1.9, 0, 2.8, 
    4.2, 3.3, 5.3, 4.6, 5.7, 6.1, 4.8, 3.7, 3.2, 1.1, 0.7, 0.5, 2, 1.9, 2, 
    3.5, 3.3, 2.4, 2.6, 2.9, 3.6, 4.3, 4, 3.9, 3.8, 3.5, 4.4, 3.9, 3.3, 4, 
    3.3, 3.9, 4.6, 5.1, 5.1, 4.8, 4.2, 3.9, 5, 5.9, 6.6, 3.6, 4, 5.1, 4.5, 
    3.8, 6.1, 5.9, 3.1, 4.6, 4.8, 3.7, 3.1, 3.8, 3, 3.9, 3.7, 6.1, 5.9, 5.3, 
    5.5, 4.6, 3.9, 4.9, 4, 6.3, 5, 4.4, 3.8, 3.6, 4.2, 5, 4.9, 0.4, 1.1, 1.8, 
    0.3, 1.6, 6.8, 3.3, 2, 2.5, 0.9, 0.4, 2, 0.9, 1.3, 1.9, 1, 4.5, 1.7, 1.3, 
    2.9, 1.4, 0.8, 0.4, 1, 1.3, 3.2, 2.6, 4.6, 4.3, 4.3, 3.8, 4.1, 4.3, 4.6, 
    4.9, 5.1, 7.4, 5.8, 6.2, 7.2, 7.9, 8, 8.8, 10.9, 12, 12.9, 12.4, 13.4, 
    14, 14.8, 13.9, 13.1, 11.8, 11.5, 12.5, 13.7, 14.5, 14.3, 14.3, 14.1, 
    12.8, 12.8, 12.9, 12.2, 10.6, 9, 8.9, 7.1, 5.4, 3.2, 2.5, 1.9, 1.8, 1.5, 
    1, 2.1, 3.4, 3.1, 2.4, 1.9, 2, 1.4, 1.1, 0.8, 0.7, 0.2, 1.2, 1.8, 1.6, 
    2.2, 2.3, 1.9, 1.5, 1.8, 2, 1.9, 2, 1.6, 1.5, 2.1, 2.2, 2.1, 2, 1.5, 1.5, 
    2.2, 1.9, 1.8, 2.1, 1.7, 2.3, 2.6, 2.7, 2.8, 3.5, 3.7, 8.7, 7.7, 10.8, 
    11.3, 12, 12.7, 12.9, 12.3, 12.2, 13, 13.5, 14.8, 13.8, 13, 11.9, 11.2, 
    11.4, 10.6, 9.7, 9.9, 10.1, 9, 9.3, 9.1, 8.4, 9.7, 10.3, 9.4, 9, 9.4, 
    9.7, 10.1, 10.5, 10.2, 9.9, 10.2, 10.8, 11, 11.7, 11.6, 11.3, 11.6, 11.8, 
    11.3, 11.4, 10.9, 10.7, 12.2, 12.8, 12.3, 11.8, 12.9, 11.2, 11.7, 9.3, 
    8.8, 9.1, 9.7, 10.7, 11.5, 10.7, 11.5, 11.6, 11.1, 11.6, 11.9, 11.6, 
    11.3, 11.5, 11.5, 11, 10.4, 9.3, 8.9, 9.2, 8.7, 8.7, 8.6, 9.3, 8.9, 9.3, 
    9.6, 10.1, 11, 11.7, 12.1, 11.9, 12.4, 12.5, 13.3, 13, 13.3, 13.6, 12.9, 
    13.3, 13.9, 14.5, 13.9, 13.9, 14, 12.5, 13.9, 14, 13.8, 12.4, 13.2, 12.6, 
    11.2, 11.1, 10.7, 9, 9, 6.9, 7, 5.2, 5.5, 5.2, 5, 5.8, 6.1, 6.2, 7.7, 
    8.8, 9.9, 9.4, 9.2, 9.5, 10, 10, 10.3, 9.8, 9.4, 10.5, 9.6, 10.7, 10.3, 
    11.1, 11.5, 12.5, 12.2, 9.8, 10.1, 9.6, 10.3, 11.3, 11, 10.3, 11.3, 9.6, 
    9.4, 7.8, 7.6, 6.6, 7.9, 6.1, 6.1, 5.4, 5.1, 4.1, 5.5, 2.1, 2.5, 0.5, 
    1.9, 4.2, 5.3, 4.9, 5.3, 4.1, 6.4, 6.9, 7, 8, 9, 9.4, 6.1, 6.4, 6.1, 6.4, 
    6, 2.3, 6.3, 9, 7.5, 7.9, 7.6, 8.4, 5.7, 9.5, 8.6, 8.7, 8.7, 10, 9.9, 
    11.2, 11.3, 11.8, 11.9, 13.3, 14, 14.1, 14, 14.6, 15.5, 16.4, 16.6, 16.4, 
    16.4, 16.5, 16.2, 15.7, 14.5, 13.8, 13.9, 13.2, 12.4, 12.7, 13.5, 13.3, 
    13.9, 14.4, 12.8, 12.8, 12.7, 12, 12.4, 13, 13.3, 14.8, 13, 15, 14.3, 
    15.6, 16.9, 17.7, 17, 17.9, 18.8, 18.8, 18.2, 18.4, 19.4, 19.5, 18.9, 
    19.4, 19.5, 20.3, 19.1, 18.3, 19.2, 19.3, 18.5, 20, 20.3, 18.1, 18.3, 
    17.3, 15, 12.9, 13, 11.8, 12.6, 11.8, 9.1, 8.5, 9.3, 7.7, 6.9, 7.1, 7.2, 
    5.7, 9.4, 7.5, 8, 9, 7.8, 9, 6.9, 6.7, 9.4, 8.1, 4.3, 9.5, 8.8, 7.5, 7.1, 
    6.6, 5.1, 4.1, 4.2, 4.2, 3.4, 3.4, 6.4, 3.7, 0.8, 0.1, 0.1, 5.1, 7.2, 
    8.6, 9, 11.1, 9.5, 11.7, 11.8, 14.6, 15.8, 16.5, 13, 1.7, 7.9, 11.3, 
    13.1, 11.7, 9, 8.8, 9.8, 6.1, 7.1, 7, 6.9, 8.4, 7.8, 8, 8.3, 9.2, 9, 8.4, 
    10.3, 8, 9.5, 8.5, 8.4, 8.5, 7.5, 6.5, 7.2, 6.2, 6.3, 0.1, 3.8, 0.2, 2.5, 
    2.1, 4.6, 5.1, 5.8, 5.5, 7.1, 8, 7.9, 6.4, 6.1, 5.9, 4.1, 5.2, 4.3, 5.2, 
    5, 4.8, 4.5, 3.2, 2.5, 5.1, 4.3, 4.8, 4.3, 5.6, 4.5, 5.2, 4.5, 4.3, 3.5, 
    1.6, 2.5, 3.3, 4.4, 3.8, 3.6, 3.7, 4.4, 4.5, 3.8, 3.9, 5.4, 3.9, 5.1, 
    5.3, 5.1, 5.7, 5.1, 5.1, 5.1, 5.3, 4.9, 5, 5.5, 5.5, 5.1, 4.6, 5.3, 4.9, 
    5.1, 5.7, 5.6, 6.6, 6.4, 6.8, 6.7, 5.4, 4.6, 6.4, 5.5, 6.4, 5.7, 6.5, 
    7.1, 7.3, 8.3, 7.3, 7.2, 7.2, 7.2, 7.6, 8.9, 8, 7.6, 6.6, 5.8, 6.7, 6.5, 
    6, 4.9, 5.4, 6.2, 5.6, 6.1, 5.6, 5.5, 5.8, 5.1, 3.8, 2, 1.6, 1.5, 1.3, 
    0.1, 0.3, 1.4, 0.3, 1.4, 7.6, 7, 7.3, 7.4, 7.9, 5.9, 5.3, 0.7, 0.9, 1.5, 
    4.3, 2.7, 1.7, 2.5, 1.6, 1.8, 1.9, 1.8, 1.6, 0, 1.1, 3.5, 7, 9, 7.9, 7.4, 
    6, 6.5, 2.4, 2.9, 3.5, 3.2, 7, 5.6, 5.2, 3.6, 2.5, 1.9, 2.4, 0.3, 5.2, 
    6.4, 5.2, 6.5, 8.6, 7.1, 5.2, 3.6, 5.2, 5.8, 5.4, 5.6, 5.9, 6.7, 7.2, 
    5.4, 4.8, 3.8, 1.1, 2.4, 3.5, 4.6, 3.2, 3.5, 1.7, 4.4, 4.7, 4.1, 4.5, 
    3.8, 3.7, 5.6, 3.3, 3.8, 3.9, 4.4, 3.2, 5.6, 3, 5.2, 5.2, 5.2, 5.9, 7.3, 
    7.8, 7.9, 9.4, 10.6, 10, 9.7, 9.3, 9, 8.1, 10.1, 8.6, 8.5, 7.9, 6.6, 6.8, 
    7.3, 7, 6.5, 5.4, 6.2, 6.4, 5.9, 5.2, 4.4, 2.4, 2.7, 1.8, 1.5, 1.7, 2.2, 
    2.6, 1.6, 0.3, 2, 0.2, 1.2, 0.4, 0.2, 9.9, 10.5, 9.4, 12.6, 10.6, 11.9, 
    14, 13.9, 13.4, 15.2, 15.8, 14.6, 14, 15.1, 17, 17.2, 17.1, 16.4, 16.5, 
    17.4, 17.7, 17.9, 18.6, 18.2, 18.3, 18.5, 17.8, 17.5, 17.6, 19.2, 20.2, 
    20.5, 20.1, 18.5, 16.5, 16, 17.6, 17.6, 18, 18.9, 20.3, 21.2, 22.8, 22.9, 
    23.6, 23.3, 23.2, 23.2, 22.5, 24.8, 23.8, 23.3, 24.2, 22.9, 19.8, 19.1, 
    19.1, 22.5, 21.5, 20.1, 13.4, 11.2, 15.7, 15.7, 17.4, 18.9, 18.3, 19.4, 
    17.3, 16.8, 16.9, 17.5, 16.1, 14.8, 9.3, 7.6, 6.9, 7.2, 1.4, 9.5, 13.6, 
    14.5, 14, 12.7, 10, 4.5, 4.4, 7.7, 7.5, 8.3, 7.9, 8.8, 8.4, 7.4, 8.1, 
    5.7, 7.9, 7.5, 7, 7.6, 5.9, 2.3, 6.9, 7.8, 6.9, 6.1, 4.4, 4.2, 4.5, 3.2, 
    3.7, 2.7, 2.2, 1.4, 3.8, 3.6, 4.4, 4.1, 3.4, 3.2, 3.4, 2.9, 2, 4.2, 5.4, 
    4.5, 5, 5.1, 7.6, 6.7, 6.9, 6, 5.8, 4.5, 3.6, 2.1, 5, 5.9, 5.8, 6.3, 4.2, 
    4.4, 2.8, 7.6, 7.6, 10.3, 11, 10.7, 10.6, 9.6, 10.1, 10.1, 11.9, 12.2, 
    10.8, 11.3, 13, 8.7, 5.9, 6.3, 7.9, 6.3, 4.9, 11.7, 11.6, 11.8, 9.9, 9.7, 
    11.7, 10.8, 11.2, 12.4, 10.6, 8.4, 8.6, 7.7, 6.7, 8.9, 10.8, 10.1, 10.8, 
    9.1, 8.7, 9.6, 10.8, 8, 8.9, 11.7, 10.8, 12.8, 14.1, 12.3, 12.7, 12.6, 
    12, 15.1, 14.7, 13.3, 13.7, 13.8, 12.8, 12.7, 12.9, 13.1, 13.4, 15.1, 15, 
    15.1, 14.3, 14.5, 14.3, 13.5, 13, 14.1, 14.2, 12.1, 14.7, 11.8, 10.6, 
    11.8, 10, 12.8, 14.3, 13.3, 12.9, 11.2, 8.8, 9.4, 9.4, 7.9, 8.9, 9, 8.3, 
    9.8, 8.2, 8.4, 8.7, 12.9, 9.5, 13.6, 16.2, 17.7, 17.8, 16.5, 14.6, 13.8, 
    14.4, 13, 12.8, 12.2, 11.3, 8.5, 8.5, 8.8, 8.2, 7.5, 5.4, 4.2, 4.1, 3.6, 
    5.8, 8.9, 9.1, 7.1, 6.6, 7.9, 7.7, 8.1, 4.3, 3.8, 3.7, 2.7, 2.9, 2.9, 
    2.2, 1.7, 0.2, 1, 1.7, 0.8, 0.2, 0.3, 2.8, 3.1, 2.2, 2.9, 4, 2.1, 2.2, 1, 
    0.4, 0.9, 0.2, 1, 0.9, 1.2, 1.8, 5.8, 6.3, 5.9, 4.4, 4.1, 3.4, 5.7, 5.5, 
    4.6, 2.5, 2.2, 1.1, 2.4, 2.1, 0.8, 1.3, 0.5, 0, 0, 2.7, 2.1, 3, 3, 4.3, 
    3.9, 6.3, 4.8, 4, 3.4, 1.5, 4, 4.2, 3.8, 3.9, 4.8, 4.1, 4, 2.8, 3.6, 2.3, 
    1.1, 3.4, 3.1, 2.4, 1.2, 1.4, 2.4, 0.9, 1, 1.3, 1.6, 1.2, 0.6, 1.4, 0, 0, 
    0.8, 1, 2, 0.9, 1.5, 1.9, 1.7, 0.7, 1, 1.8, 1.6, 6.1, 3.7, 2.4, 1.6, 0.3, 
    4.1, 0, 0.6, 4.6, 7.2, 7.1, 6.9, 6.4, 6.4, 6.4, 6.4, 6, 4.1, 1.4, 0.4, 
    3.7, 2.2, 3.4, 8.3, 9.1, 9.9, 11, 0.3, 0.1, 2.1, 1.9, 8.1, 7, 6, 5.1, 
    0.5, 3.4, 3.2, 3.4, 1.9, 3, 1.7, 1.2, 1.4, 1.5, 3.8, 5.7, 5.3, 5.9, 5.9, 
    4.7, 4.3, 3.6, 3.6, 3.4, 5, 1.9, 2.6, 2, 1.8, 1.1, 2, 1.2, 1, 0.7, 1.2, 
    0.3, 1.2, 0.9, 1.8, 2.1, 1.4, 1.4, 1.2, 1.6, 1.8, 1.3, 0.6, 1.6, 2.4, 
    0.6, 2.4, 6.1, 4.7, 5.4, 5.9, 5.4, 5.8, 7.5, 7.4, 6.5, 6.5, 5.9, 0.6, 
    0.6, 0.1, 1.2, 1.3, 2, 7.4, 7.2, 7.1, 6.2, 5.8, 2, 2, 1, 1.2, 1.6, 1.6, 
    1.1, 0.5, 1.2, 2.7, 1.7, 0.2, 0.6, 0, 0, 0.3, 0.2, 1.2, 0.9, 0.8, 2.2, 
    0.9, 1.4, 1.7, 1.2, 0.5, 1.6, 0.9, 1.5, 0.4, 0, 0, 0, 1, 0.4, 0, 0.8, 
    1.3, 1.1, 0.3, 0, 0.1, 1.3, 0.4, 1.2, 1, 0.6, 0.2, 0, 1, 0, 0.3, 6.8, 
    4.8, 2.8, 4.1, 4, 4, 9.5, 9.3, 8.5, 6.1, 8.4, 4.7, 5.9, 1.8, 2.7, 1.9, 
    1.1, 9.2, 8.8, 7.9, 6.8, 6.9, 7.5, 7.1, 6.3, 6.9, 9.1, 9.8, 6.5, 7.4, 
    8.1, 7.5, 7.3, 7.6, 6.4, 5.4, 5.3, 4.4, 3.8, 3.3, 2.6, 2.1, 0.7, 0.6, 
    0.2, 0, 1.6, 2.3, 1, 6, 6, 5.5, 4.6, 6.8, 5.8, 4.5, 5, 4.5, 2.9, 3.3, 
    4.3, 4.1, 2.8, 2.3, 1.8, 2.2, 0.3, 0.1, 0.6, 3.5, 5.1, 2.6, 3.1, 4.1, 4, 
    4.4, 3, 4.1, 4.9, 5.9, 7.8, 8.2, 10.1, 10.8, 10.8, 10, 8.1, 6.6, 5.8, 
    5.9, 7.6, 7.1, 5.5, 5.2, 3.5, 8.7, 8.4, 10.8, 11.9, 14.5, 13.6, 14.9, 
    14.8, 13.5, 13.2, 11.9, 11.1, 7.3, 5.6, 3.4, 1.4, 0.1, 0.9, 4, 3.5, 4.1, 
    4.8, 5, 4.1, 0, 0, 0.5, 1, 1.2, 0.5, 1.8, 2.8, 3.7, 7, 6.7, 6.7, 7.7, 7, 
    7.3, 5.2, 6, 5.6, 4.7, 5.2, 4.1, 2.9, 4.2, 5.4, 6.4, 6.5, 6, 6.2, 7.5, 
    8.6, 9.5, 10.1, 10.7, 11, 9.2, 11.2, 10.5, 9.3, 6.5, 3.5, 0.6, 2.2, 4.3, 
    9.2, 6, 9, 9.2, 9.7, 11.6, 8.9, 10.3, 10.1, 10.8, 10.2, 9.2, 12.5, 12.4, 
    10.9, 10.3, 10.5, 7.9, 8.5, 10.5, 11.1, 11.6, 11.2, 11.4, 10.6, 8.6, 
    11.2, 10.3, 8.1, 7.3, 7.9, 9, 8, 8.5, 8.2, 8.3, 6, 2, 2.3, 0.3, 1, 0, 
    0.2, 1.8, 2.6, 6.1, 8.4, 7.5, 8.2, 8.4, 7.9, 0.8, 0.2, 0, 1, 2.3, 3.1, 
    2.4, 3.5, 3.9, 4.5, 6.3, 6.5, 7.7, 8, 8.1, 8.2, 8.8, 9.5, 9.4, 10.1, 
    10.6, 9.5, 9.6, 9.3, 8.9, 8.4, 8.8, 8.8, 7.4, 8.3, 7.6, 7.6, 6.7, 6.2, 
    5.8, 5.6, 6.4, 7.8, 7.8, 9.2, 8, 8.6, 7.3, 3.8, 0.8, 2.5, 10.3, 10.4, 
    10.7, 12.2, 12.9, 12.1, 11.9, 12, 13, 12.8, 11.8, 14, 17.7, 16.1, 12.4, 
    14.5, 10.6, 9.8, 12.1, 12, 15.9, 11.9, 14, 12.3, 15, 13.9, 11.9, 12.2, 
    10.1, 11.7, 10.7, 11, 11.7, 14.5, 14.2, 12.3, 10.6, 9.6, 6.5, 7.7, 8, 
    8.5, 8.9, 7.4, 5.3, 7.8, 6.7, 7.3, 7, 8.6, 9.8, 9.2, 9.2, 10.2, 9.2, 7.6, 
    8.5, 8.6, 9.2, 8.8, 8.4, 10.6, 10.6, 9.6, 9, 10, 9.9, 8.8, 7.6, 7.2, 5, 
    7.5, 4.5, 4.4, 6.7, 8.7, 9.2, 9.3, 9.6, 7.1, 8.1, 9.8, 4.9, 4.3, 4.4, 
    5.4, 5.7, 3.8, 6.3, 5.8, 5.7, 6.4, 5.8, 4, 0.3, 1.6, 4, 4, 3.7, 3.1, 4.6, 
    4.7, 6.1, 5.7, 7.4, 9.5, 11.3, 10.9, 11.9, 11.7, 12, 13.3, 13, 13.3, 
    12.2, 12.3, 12.1, 11.8, 12.3, 11.6, 8.5, 8.4, 7.1, 1.7, 1.9, 3.8, 3, 3.6, 
    3.6, 4.9, 3.3, 2.9, 1.3, 0, 0, 2.2, 2.8, 2.8, 4.1, 5.1, 5.3, 7, 6.6, 6.8, 
    6.9, 6, 6, 4, 3.9, 2.3, 1.3, 2.4, 1.8, 1.8, 2.9, 3.6, 3.7, 4, 4.6, 5.5, 
    5, 4, 4.8, 4.6, 3.9, 3.4, 3.2, 3.2, 3, 1.8, 1.2, 1.4, 0, 2.5, 2.8, 5.5, 
    4.7, 4.5, 3.1, 2.5, 3.4, 4.2, 4.7, 5, 4.6, 3.7, 4.8, 5.3, 6.8, 6, 6, 6.5, 
    6.3, 5.5, 5.6, 4.2, 4.2, 5.5, 3.9, 2.7, 2.5, 3.5, 2.5, 1.3, 0.7, 0.4, 
    0.7, 1.8, 1.2, 1.9, 4.3, 5.4, 6, 2.3, 2.8, 2.2, 1.3, 0, 0.5, 2.2, 1.3, 
    1.2, 1.9, 2, 2.7, 2.8, 4, 5.3, 2.9, 4.2, 3.7, 3.4, 3.5, 5.8, 6.3, 5.5, 
    3.8, 5.1, 5.2, 0.9, 0.3, 0.3, 0, 1, 0.3, 0.8, 0.7, 0.5, 0.1, 0, 0, 0, 0, 
    0, 0.7, 1.2, 0.7, 0.1, 0.6, 1, 1, 1.7, 2.2, 2.2, 2.5, 4.5, 4.4, 4.8, 4.6, 
    4.5, 5.1, 5.3, 5.3, 5.4, 4.9, 4.6, 3.9, 4.2, 3.5, 3.3, 4, 4.3, 4.5, 3.4, 
    3.6, 3, 2.8, 2.1, 0.8, 1.1, 0.2, 0, 0, 0, 0, 0, 0, 0, 0.9, 3.4, 2.9, 2.7, 
    3.1, 2.7, 2.1, 1.8, 0.8, 2.7, 3.7, 5.1, 4.6, 6.6, 5.4, 5.8, 6.2, 5.9, 
    5.5, 7.6, 7.4, 6.9, 7.8, 8.6, 7.8, 6.8, 7.1, 8.3, 7.3, 7.4, 8.2, 8.9, 
    7.7, 7.4, 6.9, 7, 4.7, 5.6, 6.6, 8.4, 9.4, 8.2, 7.5, 7.5, 7.8, 7.3, 6.5, 
    7, 7.5, 6, 5.2, 5.1, 6.5, 5.6, 3.4, 1.4, 0.3, 0.2, 5.2, 5.8, 4.7, 5.8, 
    6.6, 7, 7.2, 7.1, 6.8, 7, 6.2, 5.7, 6, 6, 5.7, 5.6, 5.2, 4.8, 4.3, 3.9, 
    3.8, 4, 3.7, 3.5, 4.4, 4.5, 4.2, 4.5, 4.9, 4.6, 3.6, 4.3, 7, 8.7, 8.6, 
    7.5, 8.5, 8.5, 7.3, 8.8, 7.5, 6.6, 8.7, 8.2, 7.9, 7.7, 7.3, 7.1, 7.4, 
    7.9, 7.4, 9, 8.8, 9.2, 11.6, 12.1, 11.7, 13, 13.2, 13.9, 13.3, 12.7, 
    10.5, 10.1, 11.6, 11.7, 10.2, 10.7, 10.9, 9.7, 9.6, 8.8, 7.2, 10, 9.6, 
    9.6, 8.7, 8.8, 9.6, 10.4, 11, 10.4, 10.5, 10.3, 10.7, 11, 12.1, 11.2, 
    12.1, 11.5, 10.6, 11.7, 12.3, 12.8, 12.9, 13.5, 12.5, 12.1, 11.9, 10.7, 
    10.5, 8.7, 7.2, 6.8, 7.6, 8.2, 8.9, 9.1, 11.2, 12.4, 12.8, 13.5, 14.2, 
    14.5, 14.4, 14.3, 14.7, 14.8, 14.6, 14.8, 14.6, 14.4, 13.2, 12, 11.1, 
    10.2, 7.2, 4.6, 1.8, 2.3, 5.4, 6.2, 6.9, 6.5, 5.6, 3.1, 1.6, 0.4, 0.2, 
    0.8, 2, 2.7, 3.3, 3.8, 5.3, 5.2, 5.7, 7.6, 7.7, 8, 8.3, 8.6, 8.6, 9.9, 
    9.8, 10.4, 9.5, 9.3, 10.9, 12.1, 13.3, 13.1, 11.4, 7.3, 8.9, 4.7, 5.2, 
    4.2, 3.1, 1.6, 2.2, 2.6, 2.1, 0.5, 4.2, 1.4, 4.4, 3.7, 1.6, 0.2, 0.1, 
    1.4, 4.2, 7.5, 9.8, 8.8, 11.3, 12.7, 13.7, 13.5, 14.5, 16.1, 16.9, 17.8, 
    16.5, 16.5, 20.1, 20.4, 19.5, 19.3, 19.4, 18.1, 16.8, 16.4, 15.2, 14.9, 
    11.2, 10, 9.4, 8, 6.1, 4.5, 2.7, 1.8, 0.4, 3.4, 4, 3.9, 5.7, 4.6, 4.7, 
    4.3, 2.8, 2.3, 2.6, 3.3, 2.4, 0.2, 0.1, 1.5, 1.5, 3.1, 6.3, 5.9, 5.2, 
    7.9, 12.4, 12.7, 8.4, 10.3, 11.9, 12.5, 12.7, 9.9, 9.9, 10, 11, 11.9, 
    12.2, 11.8, 11.3, 11.9, 11.5, 11.6, 12, 12.1, 11.1, 11.6, 12.1, 9.9, 10, 
    9, 9.3, 8.3, 7.1, 6.8, 8.5, 5.3, 3.1, 2.1, 2.3, 2.2, 5.1, 6.9, 8.7, 9.3, 
    11.7, 11.5, 11.6, 14.2, 13.2, 13.7, 13.1, 13, 11.8, 10.3, 12.8, 12.7, 
    12.4, 11.6, 4.7, 2.8, 3.4, 5.3, 4.7, 4.5, 4.8, 1.2, 3.1, 2.6, 2.1, 0.3, 
    0.9, 1.8, 3.2, 3.6, 4.9, 5.1, 5.8, 6.7, 6.5, 6.1, 5.5, 6.6, 6.7, 4.5, 
    5.3, 6.5, 6.3, 5.6, 4.7, 4.7, 3.7, 3.5, 2.6, 3.4, 3.3, 1.9, 1.7, 0.6, 
    0.8, 0.3, 0.4, 1.5, 1.5, 2.9, 2.7, 2.4, 3.4, 4.1, 5.9, 6.1, 7.6, 7.3, 
    9.1, 11.4, 11.1, 11.1, 11.6, 12.5, 13.4, 13.6, 13.6, 13.3, 12.9, 13.6, 
    14.8, 11.4, 10.6, 11.3, 16.2, 15.7, 15.1, 16.4, 18.9, 17.7, 17.9, 18.5, 
    21.8, 22, 18.9, 18.6, 18.9, 19.6, 19.6, 20.3, 20.4, 21.3, 22, 19.2, 17, 
    15.5, 14.8, 14.2, 13.1, 12.4, 13.2, 12.5, 12.5, 12.1, 12.4, 11.3, 11.1, 
    12.3, 12.7, 12.9, 14.2, 13.6, 14, 12.5, 11.5, 14.7, 12.6, 12.7, 11.8, 
    10.1, 10.8, 9.9, 10.8, 10.9, 10.8, 11.8, 11.3, 11.5, 15.3, 15, 14.2, 
    14.1, 14.5, 13.4, 12.9, 13.7, 13.5, 13.5, 12.1, 12.2, 13.7, 11.3, 9.8, 
    7.7, 11.3, 13.4, 12.8, 11.3, 11.6, 11.8, 15.1, 11.3, 12.6, 11.7, 10.5, 
    9.6, 9.8, 2.3, 4.4, 3.7, 6.3, 2.4, 2.6, 1.3, 2, 10.9, 11, 9.4, 10.5, 8, 
    1.8, 3.5, 3.4, 2.7, 0.8, 2.7, 3.7, 6.3, 5.6, 5.4, 5.8, 5.5, 4.9, 6.2, 
    4.4, 3.6, 3.1, 2.3, 2.2, 1, 0.4, 1.4, 1.6, 1.2, 1, 0, 0, 0, 1.1, 1.8, 
    3.4, 4.4, 5.1, 4.1, 3.8, 3.6, 2.5, 2.4, 2.5, 3.3, 4.1, 4.4, 3.8, 3.6, 
    3.8, 3.3, 2.3, 1.6, 0.9, 1.6, 1.8, 4.2, 4.7, 5, 5.5, 5.8, 3.7, 3.6, 1.3, 
    1.1, 1.5, 3.3, 3.4, 1.6, 2.1, 3.1, 3.3, 4, 4, 3.1, 2.7, 2.1, 1.9, 1.8, 
    2.6, 3.7, 5.5, 7, 8.9, 9.9, 10.8, 10, 10.8, 11.2, 10.5, 10.4, 11.7, 11.6, 
    11, 10.1, 9.5, 7.3, 6.5, 7.3, 5.6, 5.6, 5.2, 5.1, 4.9, 5.5, 3.9, 2.6, 2, 
    8.6, 8, 9.3, 9.5, 9.1, 8.7, 6.6, 5.9, 5, 4.4, 4.1, 4.8, 4.2, 4.4, 3.6, 
    3.4, 2.7, 2.6, 4.7, 6.2, 5.8, 6.9, 7.2, 7.5, 8.7, 10, 10, 9.1, 8.6, 8.2, 
    8.1, 7.7, 7, 6.5, 6.1, 6.9, 5.2, 6.8, 6.8, 7.2, 8.2, 6.4, 8.6, 9.5, 8, 
    9.7, 9.1, 7.2, 5.6, 6.6, 6.2, 4.2, 2.7, 1.5, 1.3, 1.3, 2.5, 3.2, 3, 4.3, 
    5.8, 6.9, 7.4, 9.4, 9.1, 8.8, 8.4, 8.4, 9.1, 9.5, 9.3, 8.6, 7.2, 8.3, 
    8.7, 9.6, 8, 8.3, 8.8, 8.5, 8.7, 8.2, 8.9, 9.6, 7.9, 7.9, 6.3, 5.9, 5, 
    4.9, 4.4, 4.7, 3.2, 4.3, 3.9, 3.3, 3.3, 2.2, 2.7, 1.9, 1.5, 1.6, 0.1, 
    1.7, 1.3, 0.1, 1.2, 0.4, 1.3, 0.1, 0.9, 0.2, 1, 0, 0, 0.8, 1.9, 0.9, 1.1, 
    0.3, 2.5, 0.5, 0.6, 0.2, 0.3, 1.4, 2.1, 2.6, 2.1, 3.3, 1.8, 2.5, 2.5, 3, 
    2.6, 2.2, 1.6, 2.5, 2.5, 3.6, 4.7, 4.7, 3.9, 6.2, 6.1, 7.8, 8.8, 8.5, 
    9.7, 9.8, 10.3, 10.9, 11.2, 11.1, 11, 10.8, 11.6, 11, 11, 12.3, 11.7, 
    11.2, 10.7, 10.6, 10.6, 10.4, 11.7, 11.5, 11.2, 10.3, 10.3, 10.2, 10.5, 
    11.8, 11.2, 11.6, 10.5, 10.3, 8.2, 8.5, 8, 7.8, 9.3, 10.4, 10.5, 10.6, 
    9.9, 10.3, 11.1, 11, 9.3, 8.5, 11, 10.4, 11.1, 11.4, 12.1, 10.4, 9.2, 
    7.5, 5.2, 2.3, 2.5, 2.6, 13.2, 12.4, 12, 10.6, 10.3, 7.7, 7.6, 9.7, 8.2, 
    7.5, 7.9, 7.7, 7.5, 7.4, 7.7, 9.6, 9.8, 13, 15.1, 11.9, 13.6, 12.5, 11.7, 
    8.5, 8.8, 9.8, 10.4, 11.2, 11.3, 14, 10.5, 9.4, 9.3, 8.5, 5.3, 5.4, 3.6, 
    6.7, 5.5, 5.5, 6.2, 4.4, 5, 5, 4.8, 4, 4.1, 4.8, 2.8, 5.9, 7.1, 5.9, 7.1, 
    7.9, 10.2, 8.8, 8.5, 10.6, 11, 12.3, 12.3, 9.3, 10.9, 12.6, 9.9, 12.6, 
    9.9, 6, 13.3, 9.1, 10.9, 15.6, 12.2, 14.4, 13.5, 13.1, 16, 16.4, 16.6, 
    16.7, 16.7, 15.1, 13.9, 14.9, 12.1, 11.6, 10.1, 10.9, 9.4, 9.2, 5.9, 9.6, 
    9.2, 8.1, 7.4, 8.6, 7.9, 8.3, 11.7, 15.4, 18.8, 16.8, 15.8, 14.8, 19.4, 
    13.9, 16.7, 16.9, 15.9, 16.6, 21, 20.5, 19.4, 20.1, 20.8, 22.3, 21.8, 
    20.9, 19.1, 15.4, 16.7, 18.3, 16.9, 15.1, 12, 12.2, 11.7, 11.2, 11.2, 
    11.7, 15.2, 13.7, 10.7, 10.8, 12.2, 12.5, 12.5, 10.8, 12.8, 12, 13.2, 
    12.1, 11.7, 11.5, 13.6, 10.7, 11, 9.3, 8.7, 7.3, 7.1, 6.8, 5.7, 6.5, 6.7, 
    6.8, 9.4, 9.5, 7.5, 7, 7.1, 7.8, 5.9, 5.3, 5.8, 5.3, 5.8, 6.3, 5.5, 5.9, 
    6.4, 4.9, 5, 5.7, 6, 5.4, 5.4, 4.6, 5.9, 5, 5.3, 5.1, 6.5, 7.2, 7.2, 5.7, 
    6.2, 6.1, 4.7, 3.7, 4.7, 4.4, 7.8, 6.9, 8.5, 7.4, 6.9, 9, 9.3, 10.8, 
    11.9, 12.4, 12.9, 12, 12, 9.7, 9.8, 13.2, 13.6, 13.6, 11.7, 11.4, 11.9, 
    12.5, 10.5, 9.5, 7.1, 6.5, 5.8, 5.4, 4.7, 3.1, 0.6, 1.9, 1, 0.4, 6.7, 
    3.8, 0.4, 2.7, 3, 5.9, 7.1, 6.2, 6.5, 7.6, 6.5, 7, 8.3, 5.2, 3.7, 3, 3.6, 
    5.1, 3.3, 3.9, 0.4, 11.3, 10.4, 1.7, 0.4, 0, 0.3, 2.1, 0.1, 3.2, 1.3, 
    6.3, 2.1, 4.5, 6.4, 5.1, 5.1, 5.3, 4, 3.4, 2.4, 2.5, 5.1, 6.4, 8, 8, 9.4, 
    8.9, 8.4, 9, 9.4, 9.7, 9.8, 9.2, 8.7, 8.6, 9.2, 10.4, 9.4, 9.2, 8.8, 9.2, 
    10.3, 10.6, 10.3, 9.1, 7.5, 6, 7.7, 7.1, 6.9, 6.6, 7.8, 7, 6.4, 5.8, 6, 
    5.1, 8.2, 8.1, 7.3, 8.9, 10.4, 12.1, 11.5, 12, 14.4, 13.6, 14.5, 15, 
    13.9, 13.8, 14.5, 14.1, 14.4, 15.1, 17.3, 17.9, 19.6, 19.5, 19.3, 19.2, 
    19.3, 18.7, 18.8, 20.2, 20.7, 19.4, 18.4, 17.2, 16.2, 13.7, 13.6, 12.2, 
    12.3, 12.3, 11.7, 11.3, 11.9, 13.2, 13.3, 12.4, 14.3, 14.2, 13.2, 13.7, 
    14.5, 14.6, 13.6, 13.9, 13.3, 11.7, 10.2, 9.1, 7.1, 5.9, 3.6, 1.9, 0.1, 
    2.1, 0.1, 0.2, 1.1, 0, 6.7, 2.9, 1.7, 4.9, 2.7, 4.8, 3.4, 2.1, 0.3, 0, 
    1.1, 2.4, 3.2, 5, 4.8, 4.1, 4.7, 4.7, 4.6, 6.5, 7, 7.5, 6.5, 7.6, 9.5, 
    10, 9.5, 10, 11.6, 11.9, 12.8, 12.9, 13.9, 14.7, 13.9, 13.3, 13.5, 16.5, 
    18.9, 19.9, 17.7, 19, 20.8, 21.4, 19.2, 17.4, 14.6, 15.4, 11.5, 12.9, 
    12.3, 12.4, 11.8, 11.8, 12.5, 12, 11.7, 10.8, 8.5, 6.6, 3.8, 2, 1.7, 0.7, 
    0.6, 1.4, 1.5, 3, 1.2, 1.5, 1.2, 0.3, 0.9, 1, 0, 0, 0.9, 0.6, 0.6, 1.8, 
    2.5, 1.1, 0.1, 1.1, 0.5, 0, 0, 0, 0, 0, 0, 0.6, 1.3, 0, 0.9, 1.2, 0.3, 
    0.7, 2.1, 0.4, 0.3, 0.1, 1, 0.6, 0.7, 0.3, 0, 0.2, 3.2, 2.9, 4.2, 4.1, 
    3.4, 2.5, 3, 0.9, 2.7, 2.1, 2.6, 1.4, 1.7, 2, 2.2, 1.6, 1.2, 3, 2.4, 1, 
    1.8, 2, 1.6, 1.7, 0.4, 4.1, 3.7, 3.9, 4.1, 3.6, 4.6, 14.4, 1.8, 1.5, 2, 
    2.7, 3.1, 5.6, 1.1, 13.6, 13.6, 13.9, 15.8, 15.8, 17.6, 18, 19.2, 18, 
    16.4, 17.2, 16.4, 16.6, 17.1, 1.2, 3.3, 1.4, 7.2, 1.3, 8.9, 2.1, 1.6, 
    1.6, 1.8, 1.7, 1.1, 1.3, 0.7, 3.3, 1.7, 0.3, 0.4, 0.2, 1.2, 0, 1.4, 0.5, 
    1.9, 1.7, 0.9, 0, 0.1, 0.1, 0.7, 0.4, 1.5, 2, 0.1, 0.5, 0.1, 1.2, 1, 0.7, 
    0.9, 0.5, 0.9, 1.3, 2.2, 0.8, 1.7, 1.1, 0.1, 2.1, 0.5, 1, 2.3, 4.3, 5.8, 
    7.4, 7.6, 7.4, 6.4, 7.4, 6, 5.7, 5.1, 5.2, 5.9, 5.2, 6.4, 7.3, 7.5, 6.4, 
    4.9, 5, 4.4, 7.1, 5.5, 5.5, 6.4, 3.2, 2.8, 4.9, 4.6, 5.9, 5.7, 6.4, 6.2, 
    6.1, 6.1, 5.6, 6.7, 8.6, 7, 5.9, 6.4, 6.7, 8.8, 7.3, 8.5, 7.4, 7.4, 6.8, 
    7, 7.3, 9.2, 10.9, 9.7, 9, 8.2, 7.2, 7.1, 7.4, 7.2, 7.9, 8.9, 9.6, 9.3, 
    8.5, 7.6, 7.3, 7.3, 7.2, 7.2, 6.4, 5.6, 12.2, 13.6, 13.4, 12.1, 10.2, 
    9.3, 10.3, 9.5, 10.4, 10.3, 9, 7.5, 9.9, 9.3, 7.4, 7.4, 7.3, 8.3, 8.2, 
    8.8, 9.4, 11.9, 11.8, 10.3, 7.1, 7.7, 9.3, 11, 10.9, 9.7, 7.4, 6.7, 7.8, 
    7.5, 6.9, 7.5, 7.2, 7.3, 7.4, 6.2, 6.1, 5.5, 4.3, 5.8, 5.8, 5.6, 6.2, 
    5.1, 5.9, 6.2, 6, 4.3, 4.6, 4.8, 6.5, 7.8, 7.5, 6.9, 5.8, 5.3, 6.7, 7.1, 
    7.5, 7.9, 8.9, 10.2, 11.1, 11, 9.9, 8.5, 8.6, 8.9, 8.5, 8.4, 8.6, 10.3, 
    10.5, 11.5, 11, 10.6, 10.4, 9.5, 10.1, 8.7, 9.8, 7.9, 7.2, 8.6, 7.6, 7, 
    6, 7.4, 6.7, 6.3, 5.8, 6.3, 6.9, 6.4, 3.3, 1.6, 1.9, 3.4, 4.5, 6.5, 5.5, 
    4.7, 4, 4.8, 3.7, 3, 2.5, 2.4, 2.1, 3.7, 4.7, 3.6, 4, 3.6, 2.5, 1.7, 2.1, 
    2.1, 2.1, 1.6, 0.6, 0.4, 0.3, 1.2, 2, 1.7, 2, 2.6, 2, 0.8, 0, 0.1, 0.3, 
    0.2, 1.5, 2, 1.9, 1.9, 2.7, 3.3, 2.5, 2.3, 2.7, 2.9, 2.7, 3.2, 3.5, 0.3, 
    0.8, 0.6, 0.7, 0.4, 2.2, 3.5, 4.2, 4, 4.8, 5.8, 6.6, 7.2, 6.5, 8, 8.4, 
    9.1, 7.9, 7.5, 7.8, 6.9, 8, 8.2, 7.4, 8, 9.7, 10.3, 10.6, 11.5, 11.9, 
    12.7, 13.9, 13.2, 13.3, 13.4, 14.2, 13.6, 13, 12.6, 10.5, 9.7, 8.9, 8.3, 
    9.4, 10.6, 11.4, 12.1, 11.8, 11.7, 11.9, 12.2, 11.8, 10.7, 11.4, 11.6, 
    13.1, 12.6, 11.1, 10.2, 8.6, 8.8, 8.6, 9.4, 9.2, 7.7, 9.1, 7.8, 7.1, 7, 
    6, 5.5, 5.6, 6.5, 5.8, 5.5, 3.1, 0.5, 2.6, 1.6, 2.4, 3.2, 2.3, 1.9, 6, 
    6.1, 5.2, 6.1, 6.5, 7.6, 7.3, 7.1, 6.1, 3, 3, 2.4, 3.8, 5.1, 5, 6.6, 7.3, 
    9.1, 7.2, 7, 5.1, 6, 5.8, 6, 2.2, 2.9, 3.4, 4.3, 4.8, 3.2, 2, 1, 0.3, 
    0.7, 2.3, 4, 4.7, 4.2, 3.7, 2.7, 1.5, 2.2, 2.4, 1.9, 3.4, 4, 2.3, 0.4, 
    1.7, 4.9, 6.3, 1.2, 0.6, 0.3, 1.9, 1.1, 5.2, 6.7, 5.3, 4.2, 8.5, 6.7, 
    7.6, 7.9, 8.6, 7.2, 5.8, 6.6, 7.9, 8.8, 8.2, 8.8, 6.4, 6.5, 6.2, 3.9, 
    1.6, 0.2, 4.4, 2.6, 2.2, 2.9, 2.1, 2.2, 2.6, 1, 0.8, 0.7, 5.5, 2.2, 0.4, 
    3, 3.4, 3.8, 3.9, 3.9, 4, 2.9, 0.8, 3.1, 4.3, 5.9, 6.4, 6.7, 7, 7.9, 6.4, 
    6.4, 6.4, 6.5, 7.2, 6.5, 7.2, 9, 7.5, 6.9, 5.8, 4.6, 2.2, 0.4, 2.7, 3.9, 
    5, 3.1, 3.8, 3.8, 2.4, 5.2, 4.6, 4.3, 3, 0.1, 0.6, 0.3, 1.2, 3, 4.8, 7.8, 
    8.5, 8.9, 8.6, 9.7, 8.5, 7.9, 10, 12.3, 13, 12.6, 11.7, 12.6, 12.2, 12.7, 
    11.8, 10.9, 8.1, 6.7, 5.3, 4.8, 3.3, 2.6, 0.5, 0.3, 1.4, 2.4, 4.9, 4.5, 
    6.9, 8.7, 9, 9.6, 9.8, 9.4, 8.2, 7.8, 7.1, 5.9, 5.9, 5.9, 4.9, 5.8, 4.1, 
    4.3, 2.9, 2.4, 2.4, 1.2, 1.4, 0.7, 1.4, 2.3, 3, 3.8, 3.2, 3.5, 2.7, 1.4, 
    1.8, 0.5, 0.7, 2.6, 2.3, 2.5, 1.1, 0.9, 1.1, 1.8, 0.8, 0.7, 1.7, 1.7, 
    2.4, 3.5, 4.9, 5.3, 5.6, 4.8, 4.6, 4.9, 6.1, 7.8, 7.5, 7.1, 8.3, 7.5, 
    7.2, 5.8, 5.3, 5.7, 4, 3.6, 3.8, 5.3, 4.3, 3.4, 3.5, 5, 5.2, 5.4, 6.3, 
    6.5, 6.3, 7.8, 9.7, 10.9, 11, 10.7, 11.7, 11.5, 8.9, 8.9, 8.5, 7.5, 7.1, 
    5.7, 5.4, 6.8, 7, 7.5, 6.4, 4.1, 3.6, 4.5, 4.9, 4.6, 4.4, 4.2, 2.8, 1.9, 
    2.2, 3.6, 2.9, 4, 2.3, 2, 1.3, 5.5, 3.4, 1.5, 2.6, 0.1, 1, 2.1, 0.6, 0.4, 
    2.9, 1.6, 0.8, 1.1, 0.7, 0, 0.2, 0.4, 0.9, 1, 1.3, 0.2, 1, 0.4, 2.6, 1.3, 
    0.7, 1.8, 1.5, 1.7, 8.7, 7.8, 8.3, 7.9, 9.3, 7.7, 9.2, 9.1, 8.1, 10.8, 
    11.9, 9.7, 7.8, 5, 4.1, 3.2, 1.7, 6.1, 7, 6.5, 6.4, 0.9, 0.2, 6.1, 9.2, 
    7.2, 8.8, 6.8, 1.8, 1.1, 2.6, 2.4, 2, 0.7, 0.8, 0.1, 3.9, 0.1, 0.2, 2.1, 
    1.6, 1.7, 0, 1.8, 1.7, 1, 0, 0.9, 3.2, 1.4, 5, 5.6, 5.1, 5.3, 5.4, 5.1, 
    5.1, 5.1, 4, 3.5, 2.8, 2, 2.1, 1.8, 0.9, 2.3, 2.6, 3.8, 5.7, 4, 2, 2.1, 
    3.3, 2.8, 1.2, 1.1, 2.3, 2.5, 4.9, 5.9, 8.5, 9.9, 9.5, 9.8, 9.9, 10.5, 
    11.9, 10.2, 9.7, 8.8, 8.5, 7.7, 7.6, 5.6, 5.7, 7.5, 6, 4.3, 2.4, 1.6, 
    1.1, 0.7, 0.6, 1, 1.2, 2.1, 3.6, 6, 5.2, 4.1, 1.4, 1.9, 2.9, 3.3, 2.2, 
    2.2, 3, 2.5, 2.8, 3.1, 3.3, 0.3, 2.2, 2.7, 3.2, 1.5, 0.4, 2.1, 1.9, 2.3, 
    4.1, 5.4, 5.4, 4.6, 5.6, 6.3, 7.4, 6.4, 7.6, 4.1, 3.3, 1.4, 2.1, 1.5, 
    2.9, 3.4, 2.7, 5.1, 3.7, 3.1, 0.6, 3.1, 6.3, 5.6, 4.4, 4.3, 4.5, 4.7, 
    3.7, 3.6, 3.5, 2.1, 0.9, 0.2, 0.2, 0.4, 0.5, 1, 1, 0.8, 1.3, 2, 5.3, 
    10.1, 7.6, 8, 7.8, 9.6, 6.5, 8.8, 8.6, 8.5, 6.5, 6.8, 6.7, 7.6, 7.7, 5.7, 
    6.4, 4.2, 2.4, 1.3, 1.7, 3.3, 1.4, 0.2, 3.1, 3.9, 4.2, 4.8, 5, 5.4, 5, 
    5.9, 6.4, 6.6, 6.1, 5.9, 6.3, 6.2, 5.7, 5.6, 5.7, 5.1, 5.8, 6, 5.3, 4.9, 
    5.9, 5.8, 5.2, 5, 4.5, 4.1, 3.3, 3.5, 3.4, 3.3, 4.6, 3.7, 3.3, 4.3, 4.1, 
    4.1, 5.7, 1.1, 1.6, 1.9, 0.2, 1.5, 0.5, 1.3, 2.4, 1.9, 1.7, 9.9, 11.7, 
    9.6, 10.6, 4.5, 10.9, 11.8, 11.4, 11.9, 13.1, 11.8, 10.1, 7.7, 10, 10.5, 
    10.3, 9.6, 12.3, 11.6, 11.1, 10.3, 10.1, 11.4, 10, 10.4, 9.5, 9.1, 9.9, 
    10.5, 9.3, 8.8, 9.4, 8.9, 8.8, 8.4, 8, 8.2, 7.6, 7.6, 7.8, 7.6, 8.3, 8, 
    8.7, 7.6, 8.1, 8.4, 8.2, 7.5, 6.9, 6.9, 7, 8.3, 6.9, 6.5, 6.5, 6.7, 6, 6, 
    5.6, 5.8, 6.5, 5, 4.4, 3.4, 4.5, 3.1, 2.6, 2.2, 2.6, 2.5, 1.1, 1, 1.5, 
    2.6, 2.6, 0.8, 1.2, 1.1, 0.3, 4.8, 8.3, 9.4, 10.5, 7.6, 7.8, 7.9, 1.9, 
    2.7, 2.4, 3.1, 2.5, 1.6, 4.7, 4.9, 8.9, 9.7, 8.8, 6.8, 9.9, 4.4, 2.9, 
    12.1, 12.4, 11.9, 11.4, 11.2, 9.2, 8.5, 9.2, 6.2, 7.4, 5.1, 8.3, 8.3, 
    12.6, 12.9, 11.2, 5.7, 11.6, 11.2, 12.4, 10.2, 10.5, 7.1, 10.9, 12.3, 
    11.4, 10.9, 11.5, 11, 11.6, 11.2, 8.5, 10.3, 8.8, 7.3, 9.3, 5.9, 4.6, 
    4.6, 5.6, 8, 9, 7.8, 5.6, 7.5, 1.8, 5.5, 8.6, 5.9, 2.8, 1.4, 3, 1.9, 0.7, 
    1.2, 1.2, 2, 6.8, 8.3, 10, 11.8, 11.8, 9.4, 8.3, 8.2, 6.7, 8.6, 6.3, 7.9, 
    7.2, 6.5, 5.3, 5.3, 5.1, 4.5, 4.3, 4.9, 5.2, 3.7, 2.7, 3.5, 2.9, 2.2, 
    1.4, 1, 0.8, 1.4, 0.7, 1.2, 2.2, 2, 2, 1.7, 1.7, 2.1, 1.4, 2.2, 2.6, 2.3, 
    2.5, 4.3, 3.5, 2.5, 5.1, 5.8, 6.2, 5.2, 5.1, 5.1, 4.2, 6.3, 7.4, 6.6, 
    5.8, 6.5, 6.4, 6.8, 6.4, 7.7, 6.4, 5.8, 6, 6.7, 8.8, 8.5, 9.7, 9.6, 9.6, 
    9.7, 9.5, 8.5, 7.5, 8.1, 8.8, 9.4, 10.5, 8.6, 8.2, 8.2, 6.7, 5.6, 0.8, 
    2.8, 6.3, 6.8, 9.4, 10.5, 8.7, 11.2, 11.1, 9.5, 9.5, 8.6, 8.5, 8.7, 8, 
    7.3, 5.3, 6.8, 7, 7.6, 8.7, 9, 6.3, 5.2, 10.6, 12, 10.3, 6.2, 6.1, 8.6, 
    10.5, 9.4, 7.9, 10.2, 10.4, 10.3, 12.1, 10.6, 12.1, 10.5, 10.7, 10, 8.1, 
    9.2, 10.1, 10.6, 9.8, 10.6, 11, 12.3, 10.1, 9.3, 8.5, 7.9, 8.6, 8.5, 7.9, 
    6.6, 7.4, 7, 6.2, 6.3, 8.1, 9.5, 9.5, 8.6, 4.8, 4.2, 5.2, 4, 4, 4.4, 5.2, 
    6.9, 7.4, 6.1, 5, 5.8, 6.1, 5.2, 5.2, 4.6, 4.6, 4.3, 2.8, 2.8, 2.9, 3.8, 
    3.1, 1.9, 0.7, 1.2, 4.7, 1, 0.4, 2.6, 3, 3.6, 0.1, 0.9, 0.9, 1.6, 5.7, 
    1.4, 0.2, 0.1, 1.5, 4.2, 2.9, 0.8, 1.1, 2.4, 1.5, 0.8, 1.2, 0.6, 1.2, 
    0.2, 2.8, 2.3, 0.5, 1.1, 1.5, 2.3, 3.5, 3.1, 3.5, 2.9, 1.9, 1, 3.6, 4.7, 
    4.1, 4.1, 4.3, 5.4, 5.6, 6.3, 7.7, 7.8, 7.2, 8.7, 8.3, 7.7, 8.5, 10.7, 
    10.7, 10, 11.7, 17.9, 20.1, 19.6, 20.7, 21, 22.2, 21.5, 19.4, 20.5, 22.4, 
    22, 20.4, 15.9, 14, 10, 9.3, 8.8, 11.4, 10.5, 11.9, 14.4, 12.5, 11.9, 12, 
    11, 8.8, 10, 10, 10.8, 10.5, 11, 9.9, 10.4, 9.7, 10, 10.4, 11, 11.1, 9.9, 
    10.7, 9.4, 9.7, 10.1, 9.8, 9.5, 10.5, 13.8, 15.5, 13.6, 13.5, 13.9, 13.3, 
    12.9, 15, 15.7, 12.5, 12.5, 15.5, 15.8, 16.8, 15.7, 14, 15.4, 15.2, 13.5, 
    11.3, 11.8, 4.7, 7.1, 12.3, 12.3, 10.6, 10.6, 10.8, 11, 11, 11, 11.6, 
    12.1, 11.8, 7.4, 10.7, 10.5, 10.3, 9.4, 11.8, 11, 9.6, 9.6, 9, 10, 10.5, 
    9.6, 9, 6.3, 5.9, 7.7, 9.6, 8.9, 8.3, 7.6, 6.2, 5, 5.3, 6.1, 5.8, 7.5, 
    6.4, 3.9, 4.9, 3.6, 2.5, 2.2, 2, 2, 2.4, 2.4, 1.7, 1.8, 2.5, 0.3, 2.8, 1, 
    0.6, 0, 0, 0.1, 1, 0.5, 2, 2.2, 4.2, 4.8, 4.1, 4.6, 3.9, 3.8, 3.6, 5.9, 
    6.9, 4.7, 5.5, 8.7, 11.1, 5.6, 6.4, 5.6, 7.8, 6.8, 4.8, 7.3, 7.5, 7.4, 
    7.5, 7.9, 7.5, 9, 9.3, 10, 11, 11, 10.6, 13, 12.7, 9.4, 10.2, 10.7, 11, 
    10.7, 9.7, 8.1, 9.3, 9.2, 9.4, 10.3, 9.4, 11.3, 9.3, 8.2, 8.2, 7, 6.3, 
    7.4, 9.3, 9.2, 8.4, 8.1, 8.5, 7.2, 7.9, 7.6, 7.7, 6.7, 7, 9.5, 6.8, 6.8, 
    7.7, 8.1, 7.3, 7.7, 7.4, 8.8, 8, 7.7, 7.3, 7.4, 6.3, 8.2, 7.9, 8.2, 7.9, 
    6.3, 5.7, 5.6, 7.6, 6.9, 5.3, 4.5, 2.2, 0.9, 0.6, 1.8, 2.7, 3.1, 3.6, 
    1.9, 1.8, 1.8, 0.9, 0, 0.8, 0.6, 2.3, 1.6, 0.1, 0.1, 0, 0.1, 1.8, 0.3, 0, 
    0.7, 5.4, 7, 6.9, 3.2, 0.5, 0.4, 2.1, 2, 1.5, 2, 2.1, 1.9, 1.6, 0.8, 0.7, 
    0, 0.4, 0.5, 0.6, 0.5, 1.8, 1.7, 0.7, 1.2, 2.3, 4.3, 4.8, 5.4, 6, 7.4, 
    7.8, 7.4, 7.5, 7, 5.9, 5.8, 4.8, 5.1, 7.2, 5.7, 5, 4.1, 5.1, 5.4, 7.1, 
    6.9, 7.3, 7.7, 8.3, 8.9, 9.3, 9.4, 9.4, 10.6, 10.6, 10.7, 11.2, 11.3, 
    10.3, 11.1, 11.4, 11.5, 14.9, 15.6, 14.7, 14.8, 11, 8.6, 9.5, 6.5, 7.7, 
    6.1, 3.4, 4.6, 8, 12.1, 9.8, 7.8, 6.8, 7, 6.3, 7.8, 8.6, 6.7, 10.5, 11.2, 
    9.8, 12, 13.6, 13.6, 14.2, 16.3, 16.1, 13.2, 13.9, 10.8, 12.5, 8.4, 11.5, 
    9.1, 6.8, 6, 5.9, 3.8, 2.7, 2.6, 1, 1, 2.1, 3.3, 4.2, 5.8, 6.4, 7.2, 9.4, 
    11.2, 12.5, 11.9, 10.4, 7.8, 7.7, 7.5, 7.3, 7, 7.9, 6.6, 7, 7.3, 6.4, 
    9.1, 8.7, 8.3, 8.8, 9.3, 6.6, 6.2, 5.4, 6.9, 5.5, 3.2, 3.7, 3.9, 4.1, 
    2.1, 3.1, 3.7, 5, 5.2, 5.1, 4.9, 2, 1, 1, 2.5, 1.2, 0.6, 1.9, 0.7, 7.3, 
    7.1, 5.5, 8.5, 7.6, 7.8, 7.3, 9.7, 9.5, 8, 6.4, 7.6, 9.2, 8.1, 9.1, 6, 
    3.2, 3.7, 1, 1.4, 4.5, 5.8, 6, 4.8, 0.1, 1, 0.7, 0.2, 2.5, 2.9, 4.4, 4.4, 
    4.5, 4.1, 1.3, 0.5, 5.8, 0.3, 4.6, 4.7, 3.5, 2, 1.1, 2.4, 4.7, 4.6, 4.7, 
    5.2, 5.2, 6.6, 6.8, 6.3, 5.3, 4.8, 4.5, 6.8, 4.2, 4.2, 2.4, 0.8, 0.5, 0, 
    1.5, 3.3, 2.9, 2.8, 4.8, 4.6, 5.3, 10.9, 10.6, 7.4, 6.5, 5.9, 4.7, 5.8, 
    7.3, 7.4, 6.6, 8, 8.1, 8.5, 5.7, 8.9, 9.7, 7.4, 5.3, 3.4, 3, 3.1, 2.9, 
    3.7, 2.8, 2.6, 3.1, 4.2, 3.2, 1.5, 2, 2.6, 0.5, 0.1, 1.6, 0.2, 0, 0, 1.1, 
    3, 2.9, 2.9, 2.1, 0, 0.8, 2.4, 2.9, 2.9, 3.6, 5, 5.6, 6.1, 6.1, 6.4, 7.1, 
    5.1, 6, 5.3, 5, 6, 4.9, 3.2, 1.7, 0.2, 0.8, 0, 0.5, 0.2, 1, 1, 1.5, 1.5, 
    1.6, 3.5, 3.9, 5.1, 4.4, 2.8, 4.1, 5.9, 4.9, 5.8, 7, 6.1, 5.1, 4.9, 4.5, 
    5.1, 4.6, 5, 4.4, 3.4, 2.5, 2.8, 3, 2.4, 2.5, 1.9, 1.2, 0, 0.9, 0.6, 1, 
    0.9, 0, 1, 4.1, 1.6, 6.1, 6.9, 8.9, 7.6, 6.4, 6.3, 7.1, 7.3, 7.2, 6.8, 
    7.1, 9.4, 6.4, 4.4, 6, 6.6, 6.3, 6.1, 5.5, 5, 5.3, 5.8, 7, 7, 6.5, 4.4, 
    3.2, 4.5, 6, 5.4, 5, 4.9, 6.6, 7.6, 8.1, 5.8, 3.5, 3.9, 3.9, 4.3, 3.6, 
    2.1, 1.6, 2.3, 2.2, 4.7, 5.6, 6.5, 4.9, 5, 5.9, 6.3, 7.3, 7.7, 8.7, 9.4, 
    10, 10.5, 10.4, 10.7, 9.8, 10.8, 11.1, 10.9, 9.5, 9.5, 9.6, 9.1, 9.4, 
    9.1, 8.4, 7.4, 7.8, 8.1, 7.7, 8.9, 9.7, 8.6, 8.6, 10.3, 10.5, 9.9, 9.6, 
    9, 9.5, 9.5, 8.1, 8, 6.5, 5.1, 3.7, 4, 2.3, 0.4, 0, 1.4, 1, 2.7, 4, 3.4, 
    2.8, 4.7, 6.7, 7.3, 8.9, 7.2, 5.8, 6.4, 7, 8.6, 10.8, 8.5, 7.3, 9, 9.7, 
    8.9, 9.5, 9.8, 9.5, 9.2, 9.1, 8.5, 8.4, 7.9, 6.6, 7.8, 10, 8.2, 8.4, 8.1, 
    7.9, 6.2, 6.4, 7.2, 7.3, 6, 5.5, 5.2, 4.2, 3.5, 2.5, 2.3, 5.2, 3.9, 4, 4, 
    4.5, 5, 5.3, 5.4, 3.4, 4.2, 3.3, 1.7, 2.9, 5.5, 3.5, 2.8, 1.8, 2, 3.3, 
    3.4, 4.7, 4.1, 5.2, 2.6, 2.9, 2.3, 3, 2, 1.7, 3.4, 2.5, 3.2, 3.3, 2.6, 
    2.3, 1, 4.9, 3, 3.1, 4.1, 4.8, 3.9, 3.1, 0.9, 1.3, 3.2, 2.3, 2.1, 4.1, 
    4.7, 5.1, 3.9, 4.9, 2.9, 2.1, 2.7, 1.2, 2.4, 1.8, 2.8, 1.5, 1.5, 1.6, 2, 
    3.4, 2.9, 3.2, 3.3, 1.5, 1.2, 2.1, 2.6, 3.9, 4.2, 4.2, 4.3, 3.6, 5.3, 
    4.5, 2.5, 4, 2.9, 4.7, 4.2, 6.7, 5.7, 4.9, 5.5, 5.3, 3.3, 3.8, 2, 4, 6.8, 
    6.3, 8.9, 9.2, 7, 9.4, 7.9, 7.8, 7, 7.1, 6.6, 6.7, 7.1, 7.8, 6.6, 7.8, 
    6.1, 8, 7.7, 7.9, 6.4, 6.8, 6.3, 6.1, 8.4, 10.8, 10.3, 9.7, 9.8, 9.9, 
    10.3, 12.6, 14.4, 14.7, 14.8, 12, 13.7, 13.3, 12.4, 10.7, 11.3, 11.1, 
    9.7, 7.4, 10.2, 14.3, 15.8, 15, 14.3, 13.8, 13.9, 14.3, 14.2, 9, 11.5, 
    13.4, 13.9, 13.3, 15.2, 14.2, 15, 19.2, 21.6, 20.1, 22.8, 19.8, 19.2, 23, 
    21.1, 19, 18.6, 18.6, 19.8, 19.6, 22.9, 22.3, 19.8, 18.9, 15.2, 13.2, 13, 
    12.7, 12.5, 14.5, 14.5, 14.3, 12.2, 12.5, 11.7, 13.2, 13.9, 13.9, 13.2, 
    13.2, 10.2, 9.7, 10.4, 9.8, 10.4, 10.2, 10.2, 10.3, 11.5, 12.1, 12.7, 
    12.8, 13.1, 12.1, 11.3, 9, 7.7, 8.4, 8.5, 8.2, 6.5, 5.6, 5.4, 5.4, 5.4, 
    2.6, 0.9, 1.4, 1.6, 5.7, 9.8, 10.5, 9.6, 8.1, 6.6, 7.1, 6.6, 6.2, 5.8, 5, 
    4.9, 4, 4.5, 4.3, 4.3, 5.2, 5.8, 5.8, 6.3, 7.1, 6.8, 7.1, 6.9, 7, 7.2, 
    7.1, 6.6, 6.5, 6.6, 6.4, 5.7, 5.9, 6.4, 5.3, 4.8, 5.6, 5.1, 4.4, 3.4, 
    3.8, 3.4, 4, 4.3, 5.6, 5.2, 5.5, 5, 4.4, 4, 3.9, 4.5, 4.8, 6.3, 6.5, 7, 
    7.2, 6, 7.3, 6.1, 5.1, 3.9, 4, 3.8, 3.1, 8.5, 4.4, 5.9, 7.4, 8.2, 9.3, 
    8.8, 6.1, 9.2, 7, 8.7, 9.2, 7.2, 6.1, 6.1, 3.7, 3.5, 3.3, 3.8, 3.8, 4.1, 
    3.8, 3.6, 3.1, 4.4, 4.9, 4.5, 3.9, 4.3, 3.1, 5.1, 4.9, 5.6, 5.5, 6.8, 
    5.8, 7.2, 6, 6.6, 7, 6.2, 6.8, 6.7, 6.3, 8.9, 9.9, 10.5, 10.2, 11.2, 
    11.5, 13.3, 13.3, 13.7, 14.8, 17.1, 16.3, 17, 17.7, 17, 17.4, 16.7, 18.3, 
    18.9, 17.4, 18.4, 16.7, 16.2, 14.7, 11.8, 11.6, 12.5, 11, 10.9, 7.9, 8, 
    9.5, 7.8, 8.8, 10.4, 9.9, 14.8, 11.8, 14.1, 15.1, 15.7, 12, 11.8, 9.8, 
    9.7, 10, 9.5, 6.1, 7, 8.4, 8.3, 9.1, 8.5, 8.5, 9.2, 9.2, 9, 8.3, 9.5, 
    9.3, 10.4, 11.9, 11.7, 12.3, 12.8, 15.1, 14.3, 13.3, 14.7, 15.7, 16.9, 
    14.1, 13.1, 11.7, 9.8, 11.1, 8.2, 8.1, 8.9, 10.7, 12.6, 12.2, 12.7, 13, 
    13.1, 11.5, 8.6, 7.8, 7.5, 5.8, 7.1, 6.8, 6.6, 6.8, 5.2, 6, 5.8, 4.7, 
    3.3, 3.9, 3.1, 5.1, 5.2, 7.2, 7.7, 6.8, 7.3, 5.9, 4, 1.8, 2.7, 8.7, 8.1, 
    7.4, 7, 3.9, 4, 6.2, 6.9, 6.9, 6.2, 6.6, 6.4, 5.4, 6.4, 6.3, 7, 5.9, 6.4, 
    8.3, 7.8, 7.7, 8.4, 7.8, 7.6, 7.8, 8, 9.4, 8.3, 9.5, 9, 9.7, 9.2, 9.9, 
    6.2, 9.4, 7.4, 3.1, 5.5, 9.7, 10.3, 10.9, 10.6, 10.1, 8.5, 9.2, 9.2, 9.7, 
    10.4, 11.4, 11.8, 11.8, 9.7, 9, 9, 8.7, 10.1, 9.7, 7.6, 8.6, 11.5, 12.1, 
    13.2, 14, 14.1, 14.6, 13.6, 14.2, 13.4, 13, 12, 12.4, 11.6, 11.2, 11.5, 
    11.4, 10.6, 9.8, 8.9, 8.7, 8.5, 8.3, 8.9, 9.7, 9.3, 10.2, 8, 7.6, 7.5, 
    5.8, 4.1, 1.5, 0.7, 1.8, 2.7, 3.2, 3.5, 2.9, 5.6, 5.6, 6.1, 5.8, 5.3, 
    4.8, 3.9, 2.8, 3.6, 2.4, 2.5, 1.5, 2, 2.5, 4, 2.7, 2.3, 3.7, 3.7, 5, 5, 
    3.4, 2.1, 2.5, 3.7, 4.5, 4.8, 5.1, 6.9, 11.9, 13.4, 13.6, 13.8, 14, 14.4, 
    15.4, 14.8, 16, 16.2, 17.3, 16.1, 18, 17.6, 17.6, 17.6, 17.8, 18, 17.7, 
    17.5, 16.6, 15.3, 15, 14.2, 14, 13.5, 13.9, 13.4, 12.8, 11.8, 10.6, 10.2, 
    9.9, 8.3, 8.5, 7.5, 6.1, 2.4, 1.2, 0.8, 1.1, 3.7, 3.5, 3.8, 4, 5.3, 4.9, 
    5.2, 5.8, 6.2, 6.2, 3.9, 4.9, 5.8, 4.8, 0.5, 2.8, 4.8, 7.7, 5.9, 6.1, 
    3.9, 1.5, 0.9, 4.5, 7, 9, 10.2, 9.6, 9.4, 10.9, 10.8, 10.4, 10.2, 10.7, 
    10.8, 9.7, 8.7, 10.1, 12.2, 11, 10.6, 11.7, 12.3, 12.5, 14, 13.8, 13.8, 
    13.1, 15.4, 16.9, 16.6, 15.4, 14.6, 16.2, 16.7, 17.3, 17.8, 18, 20, 20, 
    20.2, 18.6, 17.1, 16.9, 18.1, 18.1, 16.7, 16.7, 15.7, 14.6, 13.3, 14.3, 
    16.1, 19.1, 16.2, 12.2, 14.6, 15.8, 15.5, 13.6, 10.8, 7.4, 9, 6.9, 8.3, 
    9.2, 10.1, 9.7, 8.9, 10.1, 10.4, 10.5, 12.1, 11.8, 12.4, 10, 11.2, 9.7, 
    9, 10.2, 10.1, 10.5, 9.6, 9.2, 8.4, 7.4, 5.3, 6.8, 6.9, 7.6, 6.8, 6.4, 
    3.7, 3.7, 5.7, 7.3, 7, 7, 7.9, 7.3, 8.6, 8.8, 8, 8.2, 6.8, 6.7, 6.5, 6, 
    6.8, 6.6, 6.2, 5.6, 5.9, 5.5, 5.6, 6.5, 6.1, 7, 6.9, 7.1, 6.8, 7.6, 7.9, 
    7.6, 8, 8, 8.2, 8.2, 6.7, 7.3, 7.2, 8.9, 8.9, 5.1, 4.9, 4, 3.6, 3.2, 2.7, 
    2.3, 1.7, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 1.6, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 11.7, 9.8, 11.4, 12.2, 12.2, 
    14.4, 15.2, 16.2, 15.9, 17.6, 16.1, 16.1, 15.5, 15.4, 14.9, 16, 16.8, 
    16.8, 16.6, 16, 16.2, 17, 16.3, 16.2, 16, 15.6, 15.9, 15.7, 15.7, 14, 
    15.3, 14.6, 14.2, 14.2, 13.7, 12.1, 12, 12.1, 13, 13, 11.2, 11.7, 12.2, 
    11.7, 11.9, 11.9, 9.4, 7.9, 6.3, 6.7, 6.4, 7, 6.8, 6.8, 7, 6, 5.4, 5.4, 
    6.3, 5.1, 6.9, 5.2, 5.7, 5.5, 5.8, 7.5, 8.5, 7.1, 8.2, 7.9, 8.7, 8.4, 
    6.9, 3.3, 4.1, 2.7, 2.7, 1.7, 3.2, 5.1, 5.7, 8.6, 9.2, 7.6, 7.1, 6.3, 
    4.7, 5.4, 7.7, 7.3, 8.4, 7.6, 6.9, 7.5, 8.7, 9.9, 10.3, 7.9, 8.1, 7.8, 
    8.1, 8.7, 8.5, 8.7, 8, 9.3, 8.4, 10.5, 11.3, 11.2, 11, 9.3, 7.7, 8, 9.3, 
    5.7, 7.8, 9.2, 8.1, 9.4, 9, 6.9, 6.5, 5.7, 7.2, 7.5, 8.7, 9.8, 10.6, 
    10.6, 11.2, 12.6, 13.3, 13.4, 13.6, 14.3, 14.5, 12.5, 12.9, 12.3, 11.2, 
    10.7, 11.9, 11.3, 9.7, 10.2, 10.3, 9.6, 10, 11.3, 11.8, 12.9, 13.3, 13.4, 
    13.3, 13.4, 13.9, 13.4, 12.4, 12.9, 14.2, 14, 14.8, 15.3, 15.3, 13.4, 
    11.9, 9.9, 9.6, 9.1, 8.3, 6.1, 5.7, 3, 1.9, 1.4, 1.5, 2.6, 5, 6.4, 7.1, 
    8.2, 8.5, 7.9, 8.3, 7.4, 9.4, 9.1, 9.5, 9.6, 11.4, 12.8, 13.4, 14.8, 
    15.1, 15.2, 14.9, 12, 8.9, 8.6, 7.9, 7, 7.5, 6.8, 6.5, 5.7, 4.5, 2.6, 2, 
    1.8, 0, 0, 7.1, 11.5, 12.9, 12.2, 12.9, 13.1, 12.2, 12.7, 13.6, 14, 14.5, 
    12.4, 12.1, 12, 9.6, 7, 6.6, 5.5, 3.6, 1.1, 1.3, 1.1, 2.5, 4.7, 6.2, 6.7, 
    7.7, 8.5, 8.1, 8.1, 8.9, 9.3, 9.3, 9.8, 9, 8.6, 8.3, 7.9, 6.6, 5.7, 5.5, 
    4.2, 3.9, 3.2, 3.7, 3.3, 1.9, 3.2, 3.6, 4.6, 12, 12.4, 11.5, 11.2, 11.9, 
    9.1, 9.1, 8.9, 5.9, 6.6, 7, 6, 5.5, 5.9, 4.8, 3.3, 4.6, 4.2, 4.4, 4.5, 
    3.6, 3.7, 2.8, 1.8, 3.7, 5.5, 10.1, 10.7, 9.2, 9.4, 8.6, 10.7, 10.5, 9.5, 
    9.5, 8, 8, 6.8, 6.7, 5.3, 6.1, 5.8, 5.4, 5.2, 3.2, 4.2, 3.8, 4.5, 1.9, 
    2.7, 4.1, 3.3, 2.4, 1.6, 2.8, 2.3, 0.9, 0.8, 2.1, 2.7, 4.4, 3.4, 4.4, 
    4.8, 4.4, 4.2, 4.3, 4.9, 5.8, 5.4, 5.9, 3.8, 6.6, 5.6, 4.1, 4.7, 5.5, 
    5.9, 7.9, 6.8, 6, 5.1, 7.3, 7.4, 6.1, 6.4, 10.4, 10.1, 11.5, 11.9, 10.8, 
    11.4, 11.1, 11, 10.9, 11.5, 10.8, 12.3, 11.6, 12.9, 11.7, 8.8, 6.1, 8.5, 
    10, 8.6, 6.9, 8.5, 6.6, 4.7, 3, 5.4, 3.6, 5.3, 5.5, 7.2, 7.2, 5.7, 7.3, 
    7.7, 7.7, 7.7, 7, 7.6, 6.3, 6.5, 5.3, 6.8, 3.1, 4.9, 4.8, 4, 3.3, 4, 4.8, 
    5.2, 4.4, 7.1, 6.4, 4.5, 6.4, 4.6, 6.4, 6.4, 5.6, 5.9, 5.3, 5.6, 7.9, 
    7.7, 6.4, 7.8, 8.1, 9.5, 9.8, 10.1, 9.7, 9.4, 10.7, 10.5, 10, 10.5, 10.2, 
    10.6, 10.1, 10.2, 9.3, 10, 10.1, 9, 8.6, 9.4, 9, 8.7, 8.4, 9.6, 9.3, 10, 
    10.1, 10.1, 10, 11, 10.6, 11, 11.6, 11.1, 11.6, 11, 11.3, 10.6, 10.1, 
    9.9, 9.6, 10.3, 11.4, 13.1, 13.8, 13.8, 14.4, 12, 13.3, 13.5, 12.6, 11, 
    10.5, 11.3, 10.9, 9.6, 9.1, 10.1, 8.9, 8.2, 9.7, 8.2, 8.7, 6.8, 5, 4.8, 
    4.1, 4.4, 4.2, 2.9, 3.2, 2.9, 2.5, 2, 4.5, 6.3, 5.7, 7, 7.9, 8.2, 8.5, 
    8.8, 9.6, 8.8, 8.5, 9.4, 8.8, 8.8, 9.4, 10, 10.9, 10.6, 10, 9.1, 7.9, 7, 
    9.7, 10.7, 7.9, 7.2, 8.6, 8.6, 7.3, 5.5, 2, 10.7, 9.9, 10.9, 11.6, 10.6, 
    10.2, 10, 10.3, 11, 10.4, 11.1, 10.4, 10.8, 12.4, 11.5, 12.2, 12.1, 12.3, 
    10.3, 11.6, 14.7, 14.5, 13.3, 16.5, 17.9, 16.5, 13.7, 12.6, 15.2, 14.6, 
    12.7, 12.1, 11.8, 9.8, 9.4, 8.1, 11.1, 10.5, 10.6, 9.8, 10.5, 10.6, 9.5, 
    10.3, 10.6, 10.1, 8.8, 6.1, 5.5, 4.2, 3.2, 3, 3.2, 2, 2.6, 2.7, 0.3, 0.2, 
    0.9, 4.2, 5.6, 6.3, 8.2, 7.9, 10.3, 11.9, 13.6, 12, 11.7, 12.2, 12.4, 
    13.6, 12.6, 11.7, 12.4, 12.3, 12.4, 9.2, 8.4, 6.7, 4.1, 8.8, 10.5, 11.8, 
    11.5, 11.3, 10.8, 10.2, 11.7, 11.6, 11.3, 11.6, 11.1, 12, 10.7, 11.3, 
    9.3, 9.3, 9.4, 10.5, 9.8, 10.4, 10.5, 8.8, 8.9, 8.7, 8.6, 8.1, 6.7, 6.9, 
    7.5, 6.4, 4.7, 4.4, 4.5, 2.1, 2.1, 3.5, 3.9, 4.1, 4.7, 5.6, 6.4, 8.1, 
    9.1, 9.9, 4.9, 5.7, 5.3, 6.1, 5.7, 8.6, 6.6, 6.5, 9.3, 7.7, 7.7, 0.7, 
    6.6, 11, 11.5, 10.5, 10.5, 10.3, 9, 9.7, 8.4, 8.7, 8.3, 6.5, 6.1, 7.7, 
    5.7, 5.9, 8.6, 10.1, 8.2, 8.2, 8.1, 6.3, 2.4, 2.4, 1.3, 0.3, 3.5, 4.9, 5, 
    2.4, 4.1, 1.3, 2.8, 3.4, 9.1, 9, 7.8, 10.7, 12.3, 12.9, 7.6, 7, 6.3, 1.1, 
    1.3, 3.5, 11.6, 11, 9.8, 3.3, 17, 17.2, 16.2, 13.2, 16, 15.9, 15.5, 16.7, 
    15.8, 16, 17.6, 18.4, 17.9, 18.6, 18.6, 19.5, 19.1, 20.3, 20.4, 18.9, 17, 
    16.5, 17.7, 18.2, 18.4, 17.7, 16, 12.5, 13.8, 12.9, 12.1, 11.6, 11.3, 
    13.4, 14, 14.3, 15.2, 15.6, 16.4, 16.5, 17.7, 18.2, 18.4, 19.3, 18.6, 
    18.9, 18.7, 18, 17, 14, 14.2, 11.9, 12.2, 11.1, 11.7, 12.1, 11.3, 9.8, 
    11, 8.8, 9.2, 7.5, 4.6, 4.1, 4.8, 4.3, 4.8, 4.2, 4.8, 5.9, 5.1, 5.8, 6.4, 
    7.2, 7.1, 6.4, 4.3, 4.2, 5, 5.6, 7.9, 7.4, 6, 4.1, 3.3, 4, 3.4, 4.3, 3.9, 
    4.7, 4, 4, 2.8, 2.1, 5.1, 4.6, 6.1, 8, 8, 7.2, 6, 6, 5.5, 6.5, 6.2, 6.1, 
    6.5, 6.2, 8.3, 8.3, 6.9, 9.8, 9.7, 9.7, 8.8, 8.6, 9.3, 8.3, 8.4, 8.1, 
    7.8, 8.1, 6.9, 6.5, 5.4, 5.6, 5, 4.4, 4.6, 5.6, 5.7, 4, 10, 9.9, 7.5, 
    7.5, 7.4, 6.3, 6, 5.4, 6.8, 7.5, 7.1, 6.8, 7.2, 6.2, 5.9, 7, 6.7, 6.3, 
    8.1, 7.3, 6.7, 6.2, 4.9, 3.4, 4.8, 6, 4.7, 0.6, 1.7, 1, 0.8, 2.7, 2.8, 3, 
    2.5, 1.2, 1.6, 2.6, 2.9, 2.9, 2.7, 2.4, 1.5, 2, 1.4, 1.6, 3, 2.8, 5, 5.9, 
    6.4, 7.3, 7.5, 8.5, 9.1, 10, 11.3, 12.1, 12.4, 11, 12.3, 11, 10.4, 13.8, 
    15.6, 16.9, 17.4, 16.8, 18, 17.5, 17.2, 16.8, 16.4, 18.1, 18.5, 16.8, 
    15.4, 14.9, 18.1, 17.3, 17.9, 11.6, 12.2, 12.3, 13.2, 14.4, 14.2, 13.9, 
    12.9, 12.8, 13.6, 13.9, 12.6, 13, 12.2, 10.8, 8.1, 10.1, 8.7, 8.7, 9.9, 
    10.1, 10.1, 9.8, 10.9, 11.9, 11.9, 12.2, 12.6, 13.9, 17.8, 19.7, 14.2, 
    11.2, 13.4, 13.9, 14.9, 16, 18.9, 18.6, 19.8, 17.8, 17.6, 18.2, 15.5, 
    13.2, 11.6, 8.3, 6, 12.3, 10.9, 7.9, 12.6, 13, 14.7, 11.3, 11.1, 12.5, 
    14, 12.2, 12.3, 12.5, 14.1, 14.5, 15.9, 14.9, 13.2, 13.6, 13.5, 13.7, 13, 
    11.7, 11.6, 12.3, 11, 8.8, 10.7, 11.7, 10.9, 11.6, 8.8, 9.7, 10.8, 14.3, 
    16.9, 18.1, 17, 15.4, 16.3, 15.2, 17.2, 13.6, 13.1, 13, 11.2, 10.3, 6.1, 
    6.2, 5.4, 7.7, 13.4, 10.6, 10.2, 8.2, 9.9, 10.3, 8.9, 8.6, 9, 9.8, 9.2, 
    8, 7.7, 9.2, 8.4, 9.4, 8.5, 7.5, 7.6, 8.7, 4.7, 7.8, 8.5, 9.5, 10.5, 
    10.7, 11.7, 11.7, 11.1, 11.9, 11.2, 11.3, 9.4, 12.8, 13.4, 12.4, 12.5, 
    11.9, 10.5, 7.9, 12.2, 13.5, 13.7, 13.6, 12.7, 14.8, 12.4, 11.4, 10.6, 
    10.4, 9.6, 8.6, 7.9, 8.4, 9, 9, 9.2, 10.8, 12, 10.5, 9.7, 11.3, 9.5, 9.7, 
    10.4, 10.3, 11.5, 11.3, 11.5, 11, 10.8, 11.6, 11.6, 11.6, 10.5, 10.6, 
    10.9, 9.2, 6.8, 6.9, 8.7, 6.3, 7.2, 6, 6, 6.3, 6.2, 5.1, 4.8, 5.1, 5, 4, 
    5.3, 4.6, 5.2, 6.7, 6.9, 7.5, 9.4, 11.8, 10.7, 10.2, 11.4, 9, 7.4, 9.5, 
    8.6, 11, 12.7, 12.8, 11.6, 13.4, 14.7, 13.3, 12.1, 11.2, 10.5, 13.1, 
    13.3, 13.9, 12.6, 7.4, 10.5, 11.6, 11.8, 10, 10.3, 9.6, 5.3, 4.8, 4.4, 5, 
    2.8, 3, 3.1, 5.1, 4.7, 4.8, 4.4, 6.7, 6.8, 5.3, 4.8, 5.5, 3.3, 3.6, 1.6, 
    2.9, 3.6, 2.7, 0.5, 4.7, 7.4, 8.5, 11.1, 12, 11.6, 10.1, 8.6, 9.3, 9.5, 
    9.5, 10.1, 10.2, 11.6, 12.2, 11.7, 11.5, 11.3, 11.5, 10.9, 11.9, 12.6, 
    12.8, 13.3, 14.1, 13.8, 13.5, 11.5, 12.9, 13.6, 12.5, 14.7, 15.1, 13.3, 
    13.3, 13.3, 11.9, 10.6, 6.8, 7.4, 7.7, 10.7, 10.1, 8.9, 9, 9.1, 7.6, 8.3, 
    7.1, 8.7, 9.6, 11.5, 11.2, 11.6, 5.9, 3.7, 5.9, 7.9, 7.1, 7.5, 8.1, 7.9, 
    8.3, 9.9, 12, 13.4, 16.5, 16.6, 15.9, 14.8, 14.6, 13.5, 16.1, 15.5, 12.9, 
    11.2, 13.2, 15, 12.8, 13.6, 12.3, 10.6, 9.8, 9.6, 8.6, 7.8, 8, 4.8, 4.2, 
    3.4, 4.3, 4.9, 6.3, 7.6, 6, 6, 6.6, 6.2, 6.8, 7.8, 8.3, 8, 8.1, 9.7, 10, 
    9.1, 8.4, 9.3, 9.1, 9.5, 9.2, 10.4, 10.7, 10.8, 10, 8.6, 9.9, 9.2, 9, 
    9.7, 9.5, 9.4, 8.5, 8.5, 8.5, 8.3, 7, 6.5, 5, 3.9, 5.1, 5.8, 6.7, 6.1, 
    6.1, 6.5, 7.5, 7.8, 6.4, 6.6, 5.3, 3.2, 1.3, 1.4, 3.4, 6.9, 7.2, 10.2, 
    9.2, 8.7, 8.5, 8.8, 8.1, 7.2, 9.5, 9.2, 9.1, 7.4, 7.2, 3, 0.9, 0.6, 3.5, 
    3.3, 3, 3.6, 5, 5.3, 13.1, 14.2, 13.8, 14.6, 14.3, 14.3, 14.4, 14.4, 
    12.8, 16.4, 14.7, 14.7, 16, 15.3, 15.2, 17.5, 16.4, 16.6, 17.5, 17.8, 19, 
    19.8, 18.1, 18.7, 19.9, 19.5, 19.6, 20.3, 18.3, 19.2, 16.9, 18.7, 17.6, 
    17.4, 17, 16.1, 15.9, 15.4, 15.9, 14.8, 14.7, 12.7, 12.3, 10.3, 10.6, 
    10.3, 9.4, 8.1, 7.5, 6.3, 5.5, 5, 4.7, 3.9, 5.6, 5, 5, 3.7, 3.6, 0.4, 
    1.9, 0.4, 1.5, 2, 6.2, 8.3, 9.1, 10.5, 10.1, 12.3, 12.5, 11.7, 10.5, 8.9, 
    7.7, 5.2, 4.8, 6.6, 6.1, 6.2, 6.8, 7.5, 6.3, 5.2, 5.6, 5.1, 8.9, 6.9, 
    7.6, 11.2, 11.5, 13.9, 15.1, 13, 14.1, 15.4, 14.8, 14.6, 15.5, 14.8, 14, 
    14.2, 13.6, 14.1, 12.6, 13.7, 12.9, 10.7, 9.2, 9.2, 4.9, 2.9, 1.9, 2.5, 
    1, 2, 2.5, 4.1, 6.7, 8.2, 10.1, 10.9, 10.4, 9.7, 9.5, 7.5, 7.1, 7.1, 6.7, 
    6.3, 6.2, 5.7, 6, 5.7, 5.2, 4.4, 4.6, 4.6, 4.4, 2.8, 5.2, 5.5, 4.2, 4.2, 
    4, 3.7, 2.4, 1.2, 7.6, 7.4, 7.4, 5.6, 3.5, 2.1, 4.8, 8.5, 11.9, 15.3, 
    14.4, 17.9, 15, 16, 17.4, 12.1, 5.4, 4.1, 3, 4.8, 4.6, 9.7, 17.3, 19.5, 
    21.1, 25, 23.7, 22.9, 21.9, 20.4, 18.8, 18.5, 16.8, 16.6, 16.7, 16.4, 
    15.4, 15, 13.6, 12.9, 11.3, 11.3, 11.3, 10.9, 11.4, 12, 10.2, 9.7, 8.5, 
    7.1, 4.1, 0.6, 8.5, 7.3, 10.5, 8.7, 9.8, 9.9, 8.9, 5.1, 6.4, 7.8, 7.8, 
    8.9, 9.6, 10.6, 11.4, 11.6, 10.8, 10.1, 10.3, 10.1, 10.3, 9.6, 8.7, 8.8, 
    9, 9.3, 9.5, 9.7, 9.6, 9.7, 9.4, 9.5, 8.9, 8.5, 7.9, 6.4, 8.5, 7.8, 8.1, 
    8, 9.2, 9.3, 10.4, 10.3, 10.4, 10.8, 11, 11.5, 11.2, 11.7, 12.6, 12.6, 
    15.3, 14.3, 15.1, 14.2, 16.5, 18.8, 19, 18.8, 17.5, 20.3, 18.6, 20.4, 
    19.7, 19.5, 18.8, 17.1, 16.7, 14.9, 15.1, 17, 15.9, 15.2, 15.1, 14.8, 
    15.1, 14.4, 14.3, 15, 13.5, 13.8, 14.8, 15, 13.9, 11.8, 10.8, 12.5, 9.9, 
    11.4, 11.4, 12.7, 11.1, 10.7, 9.3, 9.4, 7.7, 8.1, 6.1, 7.4, 4.5, 4.6, 6, 
    5.6, 5.5, 6, 1.5, 6.5, 6, 1.6, 3.1, 5.1, 4.7, 8, 8.8, 9.8, 10.3, 10.2, 
    10.2, 10.7, 11, 10.2, 9.2, 9.2, 9.8, 9, 7.8, 7.6, 9, 8.6, 10.8, 12.1, 
    12.9, 14, 15.1, 17.3, 18.3, 18.5, 18.8, 16.4, 16.6, 17.4, 18.3, 17.7, 
    17.4, 18.3, 16.5, 14.8, 15.3, 14.2, 13.5, 12.3, 11.7, 10.1, 11.9, 11.4, 
    10.2, 10.1, 10.3, 12.2, 13.2, 12.2, 11.6, 11, 11, 8.5, 8.2, 9.3, 7, 8.5, 
    8.3, 7.9, 9.3, 11.4, 10.5, 10.8, 11.2, 10.3, 8.3, 6.8, 8.9, 8.9, 9, 8.5, 
    9, 8.3, 9.5, 10.8, 11.8, 12, 11.6, 13.8, 13.7, 12.7, 12.8, 14.5, 14, 
    14.7, 13.6, 12.2, 13.5, 14.6, 14.4, 14.5, 14.6, 15, 16.2, 13.2, 13.9, 
    13.6, 14, 14.7, 14.1, 14.3, 13.8, 13, 13.6, 12.6, 11.9, 11, 9.5, 9.1, 
    8.9, 9.8, 9.3, 8.7, 3.7, 4.1, 3, 2.6, 1.6, 1.9, 2, 6.3, 7.7, 5.9, 8.9, 
    10.4, 9.4, 10.7, 9.9, 9.7, 9.7, 10.5, 9.5, 9.9, 10.3, 9, 8.5, 8.7, 7.9, 
    6, 5.6, 6, 5.8, 6.4, 5.5, 3.9, 4.1, 4.7, 9, 7.8, 8.6, 7.3, 7.3, 7.1, 8.2, 
    8.5, 8.7, 7.3, 7, 6.7, 8.3, 7.9, 8, 8.6, 7.9, 5.9, 5.4, 6.8, 8.6, 9.2, 
    10.1, 9.6, 9.4, 9.6, 8.1, 8.1, 8.9, 8.3, 7.5, 6, 5.2, 5.6, 1.9, 2.6, 6.2, 
    4.9, 3.9, 3, 3.5, 5, 6, 6.3, 4.9, 5.6, 8, 3.6, 3.1, 2.5, 6, 2.4, 1.2, 
    2.7, 5.5, 1.3, 2.4, 4.2, 2.6, 4.1, 4.5, 1.4, 6.3, 11.8, 10.2, 7.9, 7.9, 
    8.8, 7.4, 6.9, 8.2, 6.8, 11.5, 9.1, 10.6, 14.3, 11.7, 11.7, 14.2, 14.6, 
    15.8, 15.4, 16.1, 14.9, 15.4, 16, 12, 9.3, 0.9, 7.1, 14.4, 16.3, 16, 8.1, 
    0.3, 2, 3.6, 2.1, 1.8, 2.3, 3.2, 5, 2.6, 2.1, 2.6, 3.8, 3.1, 3.3, 3.5, 
    3.1, 4, 3.6, 4.3, 5.7, 7, 8.5, 9.5, 8.6, 9.2, 10.3, 11.6, 12.5, 14, 14.9, 
    15.3, 14.6, 14.4, 14.6, 15.2, 14.7, 15.1, 14.4, 14.6, 14.4, 15.4, 16.3, 
    17.7, 17.2, 19.3, 20.7, 21.5, 22.4, 21.6, 22.3, 23.1, 24.5, 21.2, 19, 
    19.5, 18.7, 19.5, 19.3, 21.9, 23.5, 23.6, 24.5, 25.7, 28, 26.6, 23.2, 
    20.9, 14.6, 8.9, 9.1, 8.8, 12.6, 11.9, 13.1, 13.1, 16.1, 15.4, 15.1, 17, 
    17.9, 16.5, 15.3, 18, 18.8, 10.6, 5.2, 4.5, 8.5, 4.4, 10.4, 11.9, 14.2, 
    14.7, 11.1, 5.1, 5, 10, 7.5, 1.5, 1.1, 2.9, 3, 4.1, 8.6, 8.8, 7, 3.2, 
    7.3, 9.4, 10.6, 11.2, 10.9, 11.7, 13.7, 12.2, 10.5, 5.1, 4.1, 5.2, 7.8, 
    1.4, 3.8, 14.2, 15.6, 12.5, 7.9, 9.5, 9.2, 4.5, 1.9, 0.6, 3.1, 2.6, 1.1, 
    0.1, 7.8, 7.9, 6.3, 4.5, 8.2, 8.7, 7.2, 4.1, 4.9, 6.8, 6, 5.8, 5.5, 5.1, 
    6.6, 5.7, 7.3, 7.2, 5.9, 8.2, 8, 3.3, 4.1, 5.6, 5.3, 3.5, 0.6, 7.4, 6.5, 
    3.2, 8.6, 8.9, 9.3, 7.8, 7, 6.7, 5.3, 5.2, 6, 5.9, 5.8, 7.2, 7.3, 8.6, 
    6.6, 8.4, 7.6, 6.9, 6.2, 7.1, 6.8, 7.4, 7.2, 7.3, 7.3, 7.2, 8, 7.1, 9.9, 
    9.9, 7, 5.4, 3.8, 10.5, 12.6, 15.4, 15.5, 13.5, 6.4, 1.5, 0.6, 6.5, 13.5, 
    0.5, 2.7, 8.9, 7.7, 7.5, 8.2, 8.1, 7.3, 7.9, 9.1, 8.6, 7.5, 6.9, 6.4, 
    6.3, 6.8, 6.3, 4.5, 3.8, 4.1, 5.1, 7.3, 6.2, 1.2, 6.3, 6.2, 5.6, 7.5, 
    7.5, 6.5, 6.3, 4.3, 5.4, 5.6, 8.5, 7.5, 6.6, 8.2, 9.6, 9.7, 9.8, 9.1, 
    8.6, 5.8, 3.2, 1.3, 6.1, 9.2, 9.2, 9.5, 8.2, 10.4, 9.6, 8.7, 7.7, 8.2, 
    6.5, 8.2, 6.5, 8.1, 8.5, 8.3, 9.7, 8.9, 8.5, 6.8, 9.7, 9.6, 9.2, 8.9, 
    8.6, 10.1, 7.5, 6, 7, 6.1, 8.4, 8.5, 9.9, 7.9, 9, 6.8, 7.7, 10, 9, 9.1, 
    10.2, 10.5, 9.1, 8.5, 9.9, 8.1, 10.2, 10, 9.4, 8.9, 8.1, 9.6, 9.9, 10.5, 
    11.2, 11.2, 12.2, 11.6, 9.7, 8.6, 11.4, 10.5, 11.4, 9.2, 9.4, 6.1, 7.1, 
    8, 8.7, 9.5, 9.9, 8.2, 6.5, 8.2, 6.8, 7.4, 8, 9.2, 11.7, 8.1, 5.1, 4.1, 
    5, 7.9, 5.9, 6.8, 7.3, 5.9, 7.3, 7.3, 4.6, 3.6, 5.9, 3.8, 1.6, 3.6, 2.6, 
    2, 1.7, 1.4, 1.8, 1.2, 0.5, 1.9, 2.7, 1.9, 1.8, 1.5, 0.6, 1.5, 1.2, 1.3, 
    1.1, 2.1, 1.5, 2.7, 3.4, 4.2, 4.8, 4.9, 4.9, 4.2, 3.3, 2.2, 0.6, 0.9, 
    0.3, 1.3, 1.4, 0.3, 1, 1.1, 1.8, 2.1, 1.5, 1.7, 1.2, 2.9, 2.4, 1.1, 1.5, 
    2.1, 3.5, 3, 3.5, 2.6, 2.4, 1, 2, 1.7, 3.3, 2.7, 4, 3.9, 7.5, 5, 5.1, 
    5.1, 4.3, 4.2, 5.5, 5.5, 6.2, 5.1, 5.6, 5.6, 4.4, 4.6, 4, 3.8, 2.9, 2.8, 
    2.7, 2.2, 2.9, 2.4, 0.5, 0.2, 0.3, 0.3, 0.6, 2, 7.4, 8, 9.4, 13.2, 13.4, 
    10.8, 9.3, 9.3, 10.3, 9.4, 10, 9, 6.5, 5.9, 5.6, 7.1, 6.5, 6.2, 6.2, 6.8, 
    7.1, 7.3, 8.6, 8.3, 8.3, 9.6, 9.3, 9.5, 8.8, 9.3, 8.1, 9.2, 8.8, 7.6, 7, 
    8.2, 8.5, 8.4, 7.8, 8.3, 7.6, 7.1, 7, 8.1, 8.4, 8.8, 8.6, 7.7, 8.1, 8.9, 
    9.4, 8.2, 7.9, 8, 7.5, 8.2, 8.3, 7.7, 8.6, 7.8, 8.1, 8.2, 8.4, 8.9, 8.8, 
    8.6, 8, 7.8, 9.4, 10.4, 9.8, 9.2, 8.6, 6, 8.4, 8.2, 8.6, 8.7, 9.8, 6.9, 
    10.4, 9.7, 10.5, 11, 11.7, 13.1, 11.7, 13.4, 12.5, 13.7, 13.6, 13.3, 13, 
    12.1, 12.3, 12.3, 11.9, 11.7, 11.2, 11, 12.4, 12.1, 12.5, 12.1, 12.2, 
    13.6, 11.9, 12.3, 11.7, 13, 13.1, 14.2, 13.9, 14.6, 13.6, 15, 15, 15, 15, 
    15, 15.3, 15.6, 14.8, 13.3, 14.2, 13.7, 12.8, 11.5, 10.7, 10.5, 10.4, 
    9.2, 9.5, 8.4, 7.9, 7.2, 7.4, 7.4, 6.2, 6.7, 7, 6.4, 6.4, 6.2, 6.4, 6.2, 
    5.2, 4.9, 4.6, 4.8, 5.5, 5.5, 5.7, 6.8, 6.6, 5.3, 6.5, 6.1, 5.4, 6.2, 
    5.3, 5.6, 5.6, 6.4, 6.3, 6.9, 7.4, 7.5, 6.6, 5.6, 5.9, 5.8, 5.8, 5.5, 
    5.9, 5.8, 6.9, 6.9, 6.6, 6.5, 8.6, 8.5, 8.8, 9.1, 9.7, 10.3, 10.9, 10.7, 
    11.9, 13, 13.5, 12.4, 12.9, 13.9, 14, 15.1, 14.4, 14.6, 13.9, 13.9, 13.8, 
    13.4, 12.9, 13.7, 13.5, 12.5, 11.7, 11.1, 11.6, 12.8, 12.8, 12.1, 10.6, 
    11.2, 12, 12, 11.7, 10.8, 10.7, 11.6, 11.5, 10.9, 10.9, 11, 11.2, 11.5, 
    12.1, 11.6, 11.6, 11.8, 12.3, 12.5, 13.1, 12.9, 11.9, 12, 12.6, 11.4, 
    9.8, 9, 8.5, 8.7, 7.3, 6.2, 5.6, 5.6, 5, 5, 4.7, 3.5, 3.4, 3.5, 3.8, 3.6, 
    3.5, 3.7, 3.7, 4.2, 4.1, 4.9, 5.3, 5.7, 5.3, 3.6, 5.4, 5.9, 5.5, 5.4, 
    6.4, 6.8, 6.2, 6.8, 6.9, 6.6, 5.9, 5.7, 6.3, 6.5, 6.6, 4.6, 6.3, 5.5, 
    7.4, 7, 6, 7, 6.9, 5.5, 6, 6, 6, 4.6, 6.2, 5.9, 9.4, 7.3, 6.6, 7.2, 5.9, 
    6.8, 5.4, 6.8, 6.6, 5.8, 7.1, 7.8, 8.2, 10.2, 10.6, 11.1, 10.4, 10.9, 
    11.8, 12.1, 11, 11.4, 12.1, 11.1, 11.5, 11.9, 10.6, 11, 13.4, 13.8, 14, 
    10.3, 10.3, 11.2, 10.8, 12.2, 14, 13.3, 11.8, 10.1, 13.6, 15.1, 16.5, 
    17.2, 17.9, 17.9, 17.2, 16.8, 17.1, 16.9, 16.3, 15.2, 14.4, 13, 12.2, 
    13.4, 13.5, 14.3, 14.2, 13.3, 10.7, 6.6, 7.5, 9.4, 9.4, 10, 11, 11.1, 
    12.1, 13.7, 14, 13.7, 12.9, 9.5, 6.7, 4.5, 8.2, 7.2, 1.1, 3.3, 1.9, 2, 
    1.4, 6.2, 9.5, 9.7, 8.9, 9.4, 10, 10.5, 10.1, 10.6, 9.9, 9.2, 9.8, 10.3, 
    9.6, 9.4, 10, 10.5, 10.5, 10.2, 9.7, 9.4, 9.6, 9.4, 7.5, 6.6, 6, 6, 5, 
    4.6, 5.1, 5.6, 5, 4.5, 2.9, 2, 0.9, 2.2, 3.7, 7.8, 6.8, 5.3, 5.5, 5.1, 
    4.8, 1.3, 0.1, 0.6, 1, 0, 2.6, 0.8, 3.4, 2.4, 4.8, 5.6, 6, 7, 7, 5.2, 
    6.4, 6.4, 6.3, 7.2, 6.9, 6.7, 6.8, 8.4, 9.1, 8.3, 8.1, 8.7, 7.9, 8, 6.4, 
    6.7, 7.4, 7.6, 7.8, 7.8, 4.2, 4.7, 3.9, 4.6, 4.1, 2.8, 4.9, 5.6, 7.7, 
    6.7, 6.1, 4.4, 1.8, 5, 4.4, 6.7, 7.2, 6.9, 7, 8, 9, 7.9, 8.6, 7, 8.4, 
    6.1, 5.5, 4.5, 2.9, 3.9, 5.2, 4.4, 3.9, 2.2, 2.4, 1.2, 3.5, 5.3, 4.4, 
    1.2, 10.5, 9, 7.6, 9.2, 9.1, 9, 7.4, 8.6, 7.8, 8.2, 7.4, 5.4, 4.8, 5.8, 
    5, 6, 5.7, 6.5, 5, 4.5, 4.6, 5.5, 6.9, 8.2, 9.3, 10.4, 10, 11.4, 9.3, 
    10.2, 10.2, 10.4, 11.2, 10.5, 13.8, 13.9, 14, 14.5, 13.8, 14.6, 13.4, 
    12.3, 15.5, 15.4, 14.6, 13.5, 14, 13.9, 13.9, 13.3, 12.2, 14.5, 14.5, 
    12.5, 10.1, 11.1, 11.3, 10, 8.4, 8.4, 7.4, 8.2, 7.3, 8, 9, 9.3, 8.6, 6.9, 
    6.3, 7.9, 8.8, 9.6, 11.4, 15.5, 13.7, 10.7, 8.6, 8.6, 9.6, 9.3, 8.8, 8.8, 
    7.2, 6.8, 7.7, 8.7, 9.5, 8.4, 7.2, 6.6, 10.7, 11.2, 12.5, 11.6, 11.7, 
    11.5, 12.2, 13.6, 12.6, 9, 8.6, 9.8, 10.9, 10.6, 10.6, 11.2, 9.2, 8, 8, 
    8, 9.9, 13, 12.2, 11.6, 11, 9.5, 9.6, 10, 8.9, 9.1, 10.4, 11.9, 10.4, 
    8.8, 9.8, 9.8, 7.8, 6.6, 4.2, 2.8, 6.1, 5.8, 6.3, 4.4, 0.2, 1.9, 6.6, 
    5.4, 5.4, 6.3, 8.2, 9.4, 9.9, 10.4, 9.5, 9.1, 8.7, 8, 6.8, 4.4, 8.4, 6.5, 
    5.1, 4.9, 7, 5.6, 7.2, 5, 5.3, 6.1, 4.6, 3.8, 1.8, 1.4, 7, 5.4, 3.5, 2.9, 
    0, 1.1, 1, 0.5, 0.9, 0, 0.3, 0.9, 4.3, 2.9, 5.1, 1.7, 4.6, 7.2, 7.1, 6.3, 
    6.5, 5.7, 7.8, 4.6, 8.2, 2, 1.7, 2.3, 3.8, 4.6, 0.6, 2.2, 0.2, 0.9, 2.5, 
    1, 1.7, 0.6, 0.4, 0.1, 1, 4.2, 6.1, 9.4, 10.5, 12.6, 13.1, 16.6, 15.3, 
    14.7, 14.9, 14.3, 14.6, 17.2, 17, 16.5, 14.7, 12.4, 11.9, 11.6, 13.1, 
    13.7, 13.5, 13.5, 13, 11.9, 10.6, 10.2, 10, 9.2, 10.4, 9.7, 10.2, 9.8, 
    9.9, 10.1, 12.4, 13.1, 12.4, 11.5, 12.9, 15.3, 14.8, 15.5, 13.6, 13.6, 
    13.5, 12.4, 12, 11.4, 10.2, 11, 9.9, 8.4, 7.9, 6.8, 8.3, 8.9, 8.8, 9.5, 
    10.4, 10.7, 8.5, 8.4, 8.8, 7.7, 8.8, 9, 6.7, 6.8, 7, 7.6, 15.4, 8.9, 7.6, 
    7.9, 12.1, 11, 10.8, 11.2, 13.4, 17.4, 19.3, 17, 15.9, 14.3, 16.7, 16, 
    15.9, 14.9, 16.5, 17.3, 16.8, 13.6, 13.5, 11.8, 11.6, 12.8, 13, 12, 11.9, 
    12.7, 13.4, 11, 12.4, 12.1, 12, 10.7, 12.6, 9, 9.9, 9.5, 12.2, 10.1, 9.7, 
    5.1, 6.4, 7.8, 6.3, 9.9, 11.5, 10.3, 9.9, 12.7, 11.6, 10.9, 13.1, 13.4, 
    14.3, 13.7, 15.8, 14.5, 14.1, 12.6, 12.8, 15, 12.6, 13.5, 13.2, 13.3, 
    13.4, 13.7, 13.7 ;

 wind_from_direction_10m = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 90, 110, 100, 140, 140, 110, 170, 130, 110, 
    130, 90, 140, 130, 130, 110, 170, 140, 110, 50, 170, 0, 140, 140, 90, 10, 
    0, 80, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 112, 121, 114, 110, 118, _, 115, 119, 123, 111, 116, 127, 
    132, 135, 135, 138, 134, 136, 123, 132, 128, 135, 134, 130, 127, 120, 
    102, 108, 116, 114, 115, 112, 111, 117, 120, 119, 121, 119, 120, 122, 
    127, 133, 132, 127, 138, 125, 130, 132, 129, 128, 113, 116, 114, 110, 
    106, 107, 109, 112, 118, 113, 118, 122, 127, 124, 120, 122, 132, 135, 
    141, 138, 132, 133, 133, 113, 109, 106, 109, 113, 111, 114, 110, 112, 
    116, 118, 121, 126, 124, 126, 117, 117, 116, 114, 117, 114, 118, 120, 
    122, 129, 120, 134, 139, 131, 127, 103, 101, 108, 120, 102, 94, 86, 86, 
    296, 327, 326, 318, 0, 356, 122, 291, 355, 358, 0, 319, 0, 0, 343, 329, 
    300, 356, 323, 259, 249, 152, 250, 292, 189, 50, 40, 22, 54, 54, 60, 66, 
    37, 46, 235, 218, 357, 272, _, 224, 259, 320, 318, 51, 77, 44, 24, 351, 
    329, 346, 319, 283, 118, 180, 315, 241, 265, 266, 240, 193, 204, 180, 
    201, 191, 268, 275, 301, 0, 0, 347, 0, 32, 321, 341, 317, 318, 331, 318, 
    203, 196, 298, 268, 309, 317, 314, 322, 98, 321, 320, 329, 318, 324, 333, 
    313, 314, 319, 311, 300, 310, 310, _, 318, 317, 313, 320, 320, 308, 317, 
    320, 322, _, 332, 308, 0, 135, 137, 137, 136, 136, 120, 125, 111, 116, 
    113, 125, 127, 133, 115, 102, 96, 98, 94, 114, 108, 114, 104, 96, 77, 98, 
    81, 139, 98, 95, 128, 88, 130, 115, 98, 125, 140, 151, 149, 152, 151, 
    132, 108, 107, 99, 103, 123, 128, 115, 123, 88, 78, 90, 76, 66, 66, 63, 
    57, 61, 67, 80, 68, 58, 57, 69, 64, 59, 65, 61, 58, 56, 54, 63, 67, 18, 
    0, 18, 97, 83, 97, 308, 310, 30, 25, 352, 238, 150, 141, 152, 144, 127, 
    122, 110, 99, 103, 104, 120, 117, 116, 117, 130, 124, 124, 114, 114, 111, 
    114, 112, 109, 119, 122, 123, 123, 118, 111, 120, 121, 119, 123, 124, 
    132, 136, 126, 124, 132, 127, 127, 133, 181, 96, 111, 110, 110, 116, 130, 
    251, 323, 313, 338, 309, 292, 311, 296, 308, 320, 267, 270, 271, 263, 
    258, 262, 266, 254, 190, 110, 113, 117, 131, 111, 93, 80, 74, 46, 347, 
    329, 326, 323, 322, 326, 324, 329, 322, 324, 131, 314, 0, 0, 146, 317, 
    83, 61, 71, 72, 80, 83, 69, 71, 69, 81, 86, 80, 83, 92, 87, 99, 102, 106, 
    108, 114, 109, 110, 113, 102, 101, 95, 99, 100, 92, 90, 89, 94, 111, 119, 
    118, 124, 119, 112, 121, 116, 118, 117, 119, 130, 132, 128, 133, 123, 
    125, 167, 118, 272, 320, 342, 341, 335, 345, 346, 354, 353, 4, 17, 39, 
    135, 110, 108, 131, 113, 117, 146, 306, 58, 52, 57, 63, 50, 59, 62, 61, 
    59, 59, 61, 61, 71, 72, 75, 89, 97, 101, 117, 110, 113, 105, 123, 119, 
    128, 123, 120, 119, 131, 119, 113, 109, 108, 117, 328, 320, 219, 330, 
    344, 327, 330, 303, 351, _, 156, 94, 127, 133, 0, 44, 187, 26, 345, 98, 
    306, 3, 260, 331, 3, 110, 117, 131, 132, 109, 0, 7, 0, 334, 130, 69, 86, 
    94, 74, 73, 76, 84, 78, 95, 108, 94, 90, 73, 79, 102, 139, 111, 109, 118, 
    105, 104, 98, 125, 117, 120, 114, 104, 114, 96, 294, 323, 299, 315, 309, 
    288, 0, 0, 0, 0, 356, 63, 331, 95, 78, 92, 124, 109, 111, 96, 81, 44, 
    108, 39, 342, 332, 338, 339, 317, 341, 324, 323, 324, 328, 336, 330, 346, 
    349, 346, 339, 340, 343, 343, 347, 348, 352, 358, 355, 359, 355, 356, 
    356, 354, 353, 9, 355, 341, 354, 318, 30, 342, 25, 49, 38, 12, 298, 306, 
    290, 335, 47, 48, 40, 325, 48, 54, 57, 57, 59, 59, 78, 86, 99, 103, 108, 
    109, 101, 97, 99, 96, 80, 84, 84, 83, 95, 87, 72, 80, 78, 88, 97, 80, 91, 
    96, 82, 89, 79, 72, 70, 80, 77, 73, 82, 64, 67, 63, 320, 355, 324, 325, 
    332, 246, 303, 325, 358, 143, 290, 297, 296, 109, 130, 305, 314, 0, 359, 
    0, 330, _, 335, 319, 313, 320, 306, 314, 314, 324, 316, 312, 314, 313, 
    316, 319, 318, 317, 320, 321, 320, 319, 314, 315, 314, 319, 318, 318, 
    312, 321, 325, 329, 334, 328, 330, 321, 250, 358, 184, 153, 140, 140, 
    138, 131, 121, 115, 115, 116, 115, 114, 114, 115, 107, 111, 108, 108, 
    108, 114, 117, 107, 21, 306, 21, 359, 347, 339, 354, 329, 321, 329, 322, 
    319, 326, 330, 354, 357, 94, 229, 108, 122, 123, 123, 115, 116, 118, 115, 
    _, 123, 114, 123, 118, 123, 124, 113, 95, 96, 120, 107, 103, 94, 102, 
    125, 129, 119, 122, 117, 105, 106, 111, 110, 112, 110, 128, 138, 128, 
    111, 120, 125, _, 122, 124, 121, 115, 120, 118, 116, 119, 117, 119, 116, 
    117, 109, 109, 117, 110, _, 114, 105, 111, 113, 120, 124, 109, 115, 108, 
    106, 98, 99, 98, 111, 126, 123, 118, 133, 128, 116, 115, 101, _, 104, 91, 
    110, 114, 134, 127, 113, 114, 121, 114, 118, 113, 162, 139, 123, 132, 
    131, 146, 131, 129, 131, 138, 135, 123, 97, 118, _, 122, 121, 114, 114, 
    116, 116, 118, 124, 116, 113, 117, 119, 110, 98, 117, 116, 115, 119, 119, 
    122, 126, 113, 115, 117, 113, 113, 109, 107, 112, 122, 114, 113, 114, 
    111, 111, 116, 113, 122, _, _, 115, 112, 105, 109, 111, 119, 113, 110, 
    110, 108, 115, 107, 109, 106, 103, 109, 95, 97, 86, 89, 90, 99, 98, 97, 
    99, 116, 128, 109, 106, 102, 87, 100, 79, _, 73, 68, 75, 84, 83, 81, 63, 
    71, 71, 66, 60, 64, 70, 69, 69, 67, 65, 79, _, _, 71, 82, 81, 71, 70, 76, 
    51, 54, 69, 65, 66, 68, 37, 52, 50, 51, 336, 276, 0, 0, 0, 0, 246, 357, 
    302, 322, 313, 324, 327, 327, 324, 329, _, 309, 300, 312, 316, 308, 317, 
    306, 309, 295, 304, 295, 308, 313, 322, 324, 321, 314, 309, 300, 290, 
    283, 290, 274, 270, 276, 261, 244, 241, 253, 261, 236, 237, 236, 238, 
    216, 209, 205, 201, 180, 161, 156, 95, 104, 126, 100, 117, 91, 71, 69, 
    68, 68, 63, 65, 59, 54, 52, 53, 53, 53, 55, 55, 52, 53, 52, 51, 52, 53, 
    54, 54, 51, 51, 47, 52, 49, 31, 303, 19, 352, 240, 319, 28, 49, 38, 36, 
    31, 21, 5, 54, 17, 24, 21, 36, 33, 17, _, 360, 27, 27, 326, 319, 314, 21, 
    21, 37, 42, 37, 47, 58, 56, 54, 127, 339, 36, 68, 84, 41, 33, 39, 38, 65, 
    42, 15, 17, 42, 26, 47, 34, 32, 35, 26, 40, 357, 34, 29, 22, 21, 36, 37, 
    33, 36, 28, 10, 24, 7, 7, 5, 1, 352, 347, 340, 335, 351, 359, 6, _, 342, 
    2, 5, 351, 26, 20, 8, 1, 18, 4, 359, 354, 360, 357, 360, 347, 342, 339, 
    350, 349, 345, 345, 335, 339, 340, 330, 337, 332, 334, 331, 333, 329, 
    334, 329, 324, 326, 327, 322, 325, 326, 326, 334, 344, 359, 354, 3, 5, 0, 
    8, 251, 307, 297, 311, 311, 309, 313, 295, 283, 279, 284, 289, 284, 299, 
    296, 300, 300, 304, _, 300, 300, 301, 311, 294, 292, 292, 296, 300, 286, 
    282, 286, 278, 275, 278, 278, 285, 278, 278, 271, 278, 281, 285, 277, 
    288, 291, 291, 289, 286, 289, 293, 300, 285, 296, 305, 303, 306, 307, 
    302, 306, 310, 318, 314, 313, 320, 323, 322, 327, 318, 332, 325, 326, 
    317, 323, 323, 333, 333, 330, 328, 319, 307, 306, 309, 311, 301, 312, 
    309, 311, _, 347, 356, 5, 14, 56, 38, 20, 10, 0, 15, 14, 10, 20, 25, 8, 
    18, 12, 8, 9, 4, 354, 347, 337, 333, 326, 319, 320, 313, 312, 318, 312, 
    311, 303, 300, 304, 301, 302, 300, 306, 299, 295, 306, 296, 297, 307, 
    305, 305, 297, 304, 309, 315, 315, 324, 330, 320, 326, 307, 343, 40, 48, 
    95, 93, 114, 98, 88, 92, 94, 85, 81, 85, 81, 78, 80, 79, 83, 80, 93, 127, 
    _, 124, 135, 111, 98, 108, 97, 126, 137, 108, 92, 1, 1, 315, 329, 332, 
    334, 341, 325, 336, 335, 329, 334, 333, 323, 323, 320, 318, 314, 309, 
    309, 309, 312, 318, 317, 315, 314, 312, 316, 308, 309, 314, _, 315, 320, 
    314, 316, 313, 316, _, 320, 333, 325, 328, 326, 323, 321, 327, 318, 322, 
    321, 329, 327, 325, 325, 321, 317, 318, 327, 328, 326, 325, 326, 325, 
    325, 332, 327, 332, 334, 333, 334, 340, 339, 345, 346, 342, 344, 338, 
    346, 345, 341, 344, 357, 352, 16, 20, 26, 46, 50, 70, 56, 51, 60, 29, 64, 
    46, 55, 67, 59, 355, 53, 48, _, 53, 56, 61, 67, 59, 56, 68, 55, 49, 58, 
    53, 69, 74, 70, 69, 61, 47, 58, 54, 62, 55, 55, 59, 50, 47, 38, 40, 32, 
    36, 27, 31, 20, 30, 21, 49, 14, 21, 17, 21, 37, 21, 29, 23, 26, 36, 49, 
    46, 45, 47, 49, 51, 56, 62, 28, 44, 46, 43, 41, 53, 41, 40, 34, 53, 62, 
    48, 82, 55, 71, 67, 87, 83, 104, 109, 118, 118, 143, 138, 137, 147, 157, 
    _, 159, 150, 147, 127, 137, 130, 137, 129, 126, 121, 121, 122, 121, 110, 
    109, 111, 114, 110, 108, 111, 107, 99, _, 107, 109, 114, 117, 116, 116, 
    118, 124, 127, 139, 131, _, 177, 91, 102, 305, 271, 319, 306, 291, 282, 
    287, 290, 293, 287, 285, 285, 287, 297, 285, 285, 279, 267, 268, 278, 
    279, 282, 289, 291, 290, 293, 282, 272, 295, 290, 305, 305, 308, _, 329, 
    0, 8, 25, 112, 85, 90, 100, 106, 83, 80, 73, 64, 68, 66, 94, 107, 89, 
    101, 117, 89, 74, 67, 79, 73, 78, 82, 110, 100, 105, 100, 100, 107, 103, 
    100, 107, 107, 104, 101, 104, 103, 103, 104, 103, 108, 112, 116, 121, 
    117, 117, 120, 117, 111, 113, 107, _, 110, 108, 110, 108, 118, 110, 113, 
    112, 120, 123, 120, 124, 175, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 1, 2, 360, 356, 0, 357, 351, 346, 341, 338, 335, 335, 
    332, 330, 329, 325, 326, 322, 323, 324, 322, 323, 314, 315, 314, 312, 
    320, 321, 320, 309, 309, 298, 315, 301, 300, 307, 310, 313, 310, 312, 
    310, 322, 314, 307, 314, 308, 300, 295, 296, 305, 312, 313, 315, 312, 
    313, 311, 316, 319, 321, 321, 321, 326, 323, _, 325, 324, 328, 327, 333, 
    339, 338, 341, 342, 341, 360, 349, 352, 258, 40, 29, 3, 26, 350, 46, 56, 
    52, 50, 53, 47, 48, 43, 43, 48, 32, 36, 23, 45, 23, 11, 30, 30, 22, 42, 
    14, 63, 40, 49, 30, 44, 52, 50, 49, 63, 48, 41, 50, 77, 106, 105, 109, 
    121, 162, 161, 163, 168, 163, 163, 175, 171, 170, 183, 171, 154, 136, 
    133, 151, 149, 150, 141, 145, 151, 150, 151, 153, 156, 151, 150, 152, 
    157, 165, 163, 159, 157, 158, 151, 140, 131, 136, 127, 126, 124, 127, 
    126, 125, 116, 118, 114, 123, 128, 117, 121, 113, 114, 128, 136, 145, 
    139, 191, 201, 204, _, 109, 187, 204, 203, 186, 153, 116, 118, 144, 125, 
    132, 136, 131, 127, 133, 128, 121, 116, 111, 99, 96, 96, 93, 92, 91, _, 
    95, 85, 76, 76, 280, 352, 0, 0, 313, 322, 315, 324, 275, 278, 277, 282, 
    292, _, 302, 298, 293, 291, 287, 288, 298, 293, 290, 291, 291, 292, 288, 
    283, 285, 283, 282, 267, 278, _, 278, 286, 285, 288, 291, 288, 296, 285, 
    296, _, 294, 279, 297, 297, 299, 299, 303, 316, 311, 305, 297, 300, 311, 
    320, 314, 299, 291, 285, 282, 286, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 239, 245, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 109, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 127, 129, 128, 119, 121, 120, 108, 
    120, 116, 108, 114, 160, 168, 127, 130, 125, 112, 150, 146, 167, 174, 
    167, 162, 148, 178, _, 202, 195, 95, 125, 109, 114, 110, 116, 136, 174, 
    177, 198, 97, 102, 119, 100, 82, 93, 106, 122, 125, 119, 64, 59, 35, 75, 
    71, 77, 67, 67, 71, 72, 76, 65, 75, 74, 90, 81, 65, 85, 90, 91, 104, 101, 
    98, 96, 95, 93, 90, 89, 93, 97, 101, 95, 94, 92, 90, 97, 95, 98, 101, 
    104, 107, 108, 109, 106, 105, 108, _, 112, 117, 111, _, 107, 111, 101, 
    105, 104, 96, 103, 104, 101, 97, 92, 84, 81, 85, 82, 73, 71, 71, 65, 67, 
    63, 65, 62, 62, 56, 54, 51, 52, 53, 53, 48, 48, 51, 50, _, 53, 45, 49, 
    45, 49, 48, 44, 45, 37, 0, 64, 79, 72, 49, 292, 313, 307, 319, 307, 312, 
    309, 303, 260, 267, 253, 243, 240, 231, 237, 232, 230, 239, 233, 245, 
    251, 247, 250, 252, 256, 244, 250, 337, 303, 337, 287, 290, 332, 357, 
    350, 336, 0, 11, 222, 126, 113, 100, 288, _, 287, 289, _, 292, 294, 284, 
    _, 284, 286, 280, 286, 284, 285, 290, 289, 291, 297, 291, 292, 289, 289, 
    298, 303, 300, 298, 300, 297, 291, 292, 296, 297, 286, 282, 290, 295, 
    279, 296, 295, 308, 321, 320, 354, 20, 29, 44, 52, 38, 17, 29, 41, 30, 
    16, 24, 31, 40, 48, 48, 48, 55, 60, 54, 52, 56, 51, 58, 61, 58, 56, 62, 
    64, 58, 56, 58, 63, 56, 55, 55, 66, 72, 72, 65, 64, 65, 66, 71, 67, 68, 
    66, 63, 61, 68, 62, 56, 57, 60, 61, 64, 62, 66, 69, 71, 73, 72, 73, 65, 
    65, 61, 67, 71, 73, 326, 353, 49, 51, 41, 64, 94, 68, 60, 75, 26, 51, 73, 
    51, _, 56, _, 82, 84, 79, 76, 87, 76, 50, 81, 69, 93, 94, 70, 72, 62, 59, 
    53, 51, 52, 50, 51, 49, 49, 52, 53, 54, 55, 62, 60, 59, 56, 54, 56, 56, 
    59, 68, 68, 64, 64, 63, 67, 67, 66, 68, 70, 67, 66, 67, 74, 67, 65, 60, 
    52, 49, 56, 51, 50, 49, 50, 43, 48, 49, 47, 48, 50, 49, 47, 54, _, 43, 
    52, 55, 60, 78, 65, 66, 58, 60, 64, 68, 71, 73, 63, 60, 57, 55, 58, 57, 
    54, 52, 51, 49, 50, 45, 49, 51, 48, 50, 45, 47, 44, 45, 42, 44, 39, 37, 
    24, 27, 17, 14, 14, 28, 36, 80, 73, 76, 87, 92, 109, 70, 77, 93, 68, 69, 
    64, 61, 61, 55, 53, 20, 54, 50, 41, 50, 46, 47, 32, 24, 24, 106, 304, 2, 
    359, 2, 14, 42, 8, 10, 2, 359, 2, 1, 2, 357, _, 3, 6, 4, 1, 1, 5, _, 3, 
    349, 338, 348, 351, 355, 345, 349, 350, 358, 349, 356, 346, 347, 1, 2, 
    345, 351, 359, 27, 37, 82, 80, 94, 103, 98, 105, 87, 98, 99, 107, 107, 
    109, 114, 109, 106, 109, 113, 103, 109, 106, 106, 103, 105, 103, 105, 
    103, 103, 103, 94, 103, 89, 83, 85, 85, 92, 89, 87, 84, 88, 83, 82, 79, 
    90, 77, 84, 82, 75, 69, 72, 68, _, 70, 63, 74, 65, 52, 52, 57, 58, 52, 
    51, 47, 49, 52, 49, 47, 47, 49, 42, 48, 49, 32, 44, 42, 7, 350, 1, 5, 12, 
    10, 1, 354, 352, 348, 340, 340, 340, 353, 348, 340, 339, 335, 342, 339, 
    338, 339, 339, 337, 343, 345, 344, 342, 337, 332, 329, 330, 336, 328, 
    335, 324, 328, 334, 332, 332, 328, 332, 330, 330, 333, 330, 333, 333, 
    325, 308, 314, 321, 320, 319, 322, 326, 324, 321, 314, 313, 305, 310, 
    302, 298, 304, 302, 303, 300, 300, 292, 289, 348, 0, 358, 341, 313, 341, 
    316, 348, 327, 311, 301, 304, 309, 309, 303, _, 301, 297, 296, 304, 314, 
    317, 308, 304, 306, 304, 295, 286, 283, 277, 280, 280, 274, 266, 259, 
    273, 292, 19, 72, 69, 74, 53, 48, 61, 54, 41, 30, 39, 98, 0, 1, 8, 336, 
    19, 19, 359, 335, 347, 341, 351, 360, 353, 348, 340, 333, 318, 321, 321, 
    _, 326, 311, 310, 311, 312, 310, 306, 308, 312, 317, 321, _, 306, 302, 
    306, 304, 309, _, 303, 302, 305, 306, 304, 293, 289, 288, 298, 307, 298, 
    302, 291, 297, 309, 288, 286, 289, 288, 287, 283, 286, 288, 288, 279, 
    259, 256, 67, 279, 59, 125, 86, 99, 104, 93, 101, 142, 114, 119, 105, 
    107, 100, 93, _, 65, 63, 38, 38, 50, 59, 51, 311, 54, 47, 48, 48, 37, 37, 
    40, 38, 43, 48, 131, 112, 22, 88, 297, 295, 54, 271, 6, _, 310, 4, 359, 
    4, 18, 18, 6, 15, 17, 21, 27, 352, 1, 11, 0, 281, 244, 18, 21, 266, 102, 
    4, 8, 19, 27, 24, 23, 12, 6, 12, 13, 10, 8, 23, 16, 6, 20, 21, 7, 350, 
    352, 352, 353, 0, 1, 8, 352, 12, 25, 359, 339, 322, 5, 342, 355, 1, 11, 
    18, 12, 13, 27, 27, _, 13, 1, 334, 17, 19, 17, 26, 273, 252, 295, 25, 53, 
    25, 15, 17, 23, 14, 17, 18, _, 34, 21, 12, 13, 26, 11, 24, 20, 4, 5, 36, 
    30, 32, 1, 358, 351, 337, 346, 343, 347, 340, 347, 334, 339, 339, 338, 
    352, 350, 342, 359, 243, 14, 1, 146, 5, 16, 333, 17, 349, 359, 17, 349, 
    11, 9, _, 27, 31, 30, 27, 32, 49, 58, 52, 48, 56, 13, 6, 21, 36, 29, 21, 
    25, 33, 21, 30, 32, 320, 303, 301, 341, 295, 328, 329, 340, 305, 333, 
    336, 333, 356, 337, 349, 350, 321, 349, 326, 318, 320, 317, 305, 330, 
    312, 326, 323, 303, 297, 309, 313, 311, 315, 306, 305, 300, 305, 283, 
    289, 282, 287, 284, 280, 273, 255, 252, 243, 271, 242, 244, 247, 230, 
    243, 225, 216, 212, 187, 233, 249, 254, 257, 282, 270, 244, 279, 347, 
    325, 2, 7, 353, 296, 326, 315, 317, 321, 329, 342, 313, 318, 329, _, _, 
    _, 353, 328, 347, 327, 322, 9, 351, 51, 57, 9, 347, 335, 324, 6, 63, 64, 
    324, 22, 12, 5, 21, 27, 21, 21, 10, 346, 3, 354, 333, 338, 317, 330, 318, 
    319, 320, 326, 316, 313, 313, 313, 312, 327, 307, 290, 308, 309, 304, 
    294, 302, 298, 302, 302, 304, 304, 304, 307, 309, 309, 305, 316, 299, 
    300, 298, 306, 300, 298, 295, 293, 288, 295, 297, 300, 296, 297, 307, _, 
    304, 301, 302, 293, 306, 302, 299, 289, 289, 296, 294, 282, 282, 284, 
    289, 287, 285, 286, 276, 283, 269, 272, 281, 276, 279, 270, 270, 273, 
    266, 273, 292, 279, 275, 278, 277, 270, 283, 289, 271, 298, 318, 319, 
    315, 229, 200, 190, 199, 190, 168, 165, 148, 185, 155, 175, 163, 162, 
    162, 166, 163, 157, 164, 171, 163, 175, 169, 160, 163, 145, 122, 108, 97, 
    101, 92, 99, 106, 120, 123, 150, 147, 152, 145, 141, 109, 106, 116, 107, 
    120, 107, 110, 132, 128, _, 106, 104, 92, 93, 94, 121, 117, 114, 115, 
    122, 126, 121, 110, 119, 114, 116, 120, 119, 120, _, 86, 81, 70, 78, 60, 
    58, 67, 61, 65, 66, 68, 67, 66, 70, 69, 61, 55, 62, 59, 67, 64, 61, 60, 
    59, 57, 49, 52, 56, 58, 65, 64, 64, 67, 66, 68, 63, 65, 68, 76, 77, 78, 
    79, 85, 120, 119, 134, 128, 119, 131, 168, 180, 179, 180, 163, 180, _, 
    166, 161, 146, 185, 167, 105, 118, 133, 128, 77, 96, 54, 91, 341, 21, 24, 
    14, 7, 8, 9, 11, 15, 22, 25, 26, 352, 351, 331, 337, 347, 344, 336, _, 
    337, _, 326, 323, 321, 322, 311, 311, 312, 316, 314, 320, 314, 330, 332, 
    342, 336, 340, 341, 343, 336, 322, 315, 320, 326, 17, 336, 345, 359, 324, 
    330, 342, 350, 354, 1, 311, 320, 331, _, 6, 117, 123, 119, 120, 82, 73, 
    100, 107, 106, 106, 100, 104, 106, 110, 106, 106, 101, 101, 101, 106, 
    105, 101, 99, 97, 95, 94, 93, 90, 89, 85, 81, 76, 74, 75, 77, 82, 88, 91, 
    101, 115, 110, 101, 106, 111, 106, 100, 94, 99, 92, 90, 75, 76, 86, 69, 
    71, 74, 79, 72, 70, 84, 86, 83, 88, 88, 82, 83, 77, 73, 66, 68, _, 63, 
    59, 65, 66, 57, 53, 55, 53, 67, 67, 63, 49, 60, 88, 51, 90, 57, 14, 350, 
    34, 323, 26, 33, 20, 79, 38, 53, 44, 47, 308, 359, 144, 159, 137, 98, 89, 
    _, 97, 256, 253, 5, 308, 331, 334, 326, 332, 314, 319, 307, 298, 310, 
    325, 316, 307, 325, 314, 311, 312, 321, 318, 316, 313, 326, 318, 308, 
    301, 305, 296, 301, 304, 295, 311, 298, 309, 295, 276, 260, 255, 257, 
    244, 230, 228, 222, 198, _, 194, 151, 116, 170, 130, 133, 121, 129, 155, 
    174, 176, 157, 155, 164, 150, 146, 170, 149, 149, 142, 135, 154, 151, 
    146, 148, 132, 126, 135, 108, 83, 95, 105, 110, 112, 108, 103, 96, 89, 
    85, _, 75, 86, 92, 78, 77, 71, 67, 77, 69, 72, 74, 77, 74, 71, 67, 66, 
    66, 61, 60, 63, 64, 66, 65, 66, 74, 73, 84, 98, 94, 86, 78, _, 74, 75, 
    77, 88, 90, 105, 110, 99, 103, 101, 89, 87, 81, 81, 78, 61, 59, 59, 54, 
    53, 42, _, 47, 65, 53, 51, 54, 43, 20, 65, 87, 82, 86, 101, 102, 102, 85, 
    69, 61, 58, 60, 63, 61, 47, 33, 49, 61, 78, 100, 102, 105, 99, 99, 92, 
    91, 83, 89, 81, 71, 54, 57, 61, 63, 69, 30, 35, 42, 51, 54, 59, 61, 70, 
    45, 5, 39, 56, 53, 43, 299, 303, 265, 268, 298, 346, 210, 37, 357, 322, 
    308, 304, 295, 27, 105, 14, 13, _, 352, 343, 343, 344, 333, 335, 340, 
    338, 347, 351, 346, 360, 357, 350, 348, 344, 352, 344, 353, 348, 12, 6, 
    360, 17, 14, 9, 14, 14, 4, 359, 354, 17, 12, 26, 359, 15, 29, 44, 55, 39, 
    37, 46, 31, 35, 46, 44, 56, 45, 343, 35, 31, 354, 70, 38, 111, 134, 356, 
    339, 72, 64, 60, 97, 75, 55, 47, 63, 31, 41, 66, 118, 35, 58, 80, 106, 
    98, 103, 104, 133, 105, 103, 125, 120, 109, 110, 120, 131, 148, 114, 122, 
    115, 124, 143, 136, 114, 125, 136, 171, 151, 136, 141, 135, 76, 106, 240, 
    200, 358, 349, 28, 93, 42, 60, 83, 84, 82, 87, 81, 53, 320, 281, 219, 77, 
    2, 43, 50, 61, 66, 22, 11, 22, 31, 33, 27, 25, 20, 16, 29, 359, 5, 333, 
    310, 278, 343, 42, 358, 339, 1, 41, 35, 25, 16, 30, 35, 10, 35, 31, 26, 
    12, _, 357, 15, 341, 335, 350, 17, 11, 2, 1, 28, 21, 3, 3, 7, 1, 22, 352, 
    355, 349, 348, 348, 4, 6, 328, 344, 342, 325, 304, 343, 332, 323, 317, 
    299, 317, 290, 304, 274, 263, 305, 281, 266, 295, 280, 299, 270, 255, 
    246, 281, 279, 286, 290, 293, 288, 281, 305, 317, 354, 18, 3, 181, 166, 
    168, 152, 136, 136, 134, 134, 122, 117, 112, 120, 115, 110, 105, 301, 
    320, 314, 292, 312, 311, 318, 314, 318, 339, 321, 345, 200, 84, 83, 88, 
    127, 118, 311, 324, 351, 311, 327, 320, 305, 302, 302, 315, 349, 342, 
    305, 7, 354, 339, 318, 345, 1, 238, 312, 287, 294, _, 290, 299, 285, 291, 
    272, 276, 273, 272, 265, 269, 280, 260, 282, 277, 280, 278, 281, 262, 
    260, 269, 277, 260, 266, 271, 254, 260, 281, 282, 283, 278, 261, 257, 
    277, 271, 271, 274, 277, 272, 281, 279, 278, 277, 274, 271, 264, 263, 
    270, 256, _, 252, 253, 252, 257, 264, 261, 267, 270, 265, 305, 291, 303, 
    295, _, 329, 325, 325, 325, 328, 326, 326, 326, 320, 328, 326, 321, 324, 
    329, 337, 337, 335, 337, 343, 342, 329, 320, 336, 337, 339, 339, 339, 
    339, 334, 334, 336, 332, 334, 333, 330, 323, 325, 325, 330, 335, 333, 
    337, 332, 333, 332, 333, 334, 337, 337, 336, 335, 334, 333, 329, 331, _, 
    330, 328, 338, 330, 345, 339, 337, 342, 345, 347, 346, 342, 333, 330, 
    335, _, 299, 308, 312, 309, 306, 306, 315, 312, 305, 295, 305, 305, 307, 
    305, 316, 311, 303, 310, 305, 318, 306, 299, 310, 315, 318, 313, 318, 
    324, 324, 332, 333, 323, 317, 329, 332, 333, 328, 332, 324, 328, 328, 
    338, 342, 334, 335, 333, 330, 332, 328, 328, 336, 334, 343, 4, 348, 333, 
    332, 333, 1, 344, 326, 325, 329, 312, 16, 7, 358, 3, 357, 358, 347, 345, 
    338, 357, 347, 350, 333, 315, 313, 315, 315, 313, 315, 310, 295, 322, 
    329, 310, 308, 316, 306, 303, 297, 289, 293, 299, 299, 296, 298, 301, 
    302, 305, 307, 307, 308, 299, 303, 302, 295, 313, 300, 304, 302, 300, 
    307, 300, 299, 297, 300, 302, 308, 314, 322, 321, 324, 310, 297, 311, 
    317, 317, 321, 319, 309, 319, 320, 321, 335, 330, 337, 347, 329, 348, 
    328, 346, 353, 326, 326, 340, 316, 313, _, 318, 312, 304, 326, 300, 293, 
    271, 1, 356, 317, 8, 14, 7, 32, 45, 43, 18, 348, 314, 327, 314, 13, 16, 
    351, 349, 341, 341, 345, 350, 346, 355, 351, 351, 352, 13, 1, 348, 348, 
    357, 342, 339, 341, 338, 338, 329, 360, 2, 300, 319, 330, 342, 339, 336, 
    329, 339, 340, 352, 342, 334, 340, 335, 331, 331, 335, 357, 347, 355, 
    351, 329, 336, 330, 329, 345, 343, 334, 337, 338, 334, 12, 24, 335, 325, 
    321, 307, 310, 302, 321, 311, 306, 311, 303, 302, 302, 297, 301, 300, 
    302, 299, 299, 301, 300, 295, 291, 294, 291, 296, 291, 288, 290, 285, 
    287, 288, 304, 305, 309, 300, 298, 302, 312, 306, 310, 326, 320, 321, 
    313, 324, 313, 315, 305, 324, 333, 11, 20, 37, 9, 342, _, 347, 350, 336, 
    316, 321, 320, 321, 320, 324, 313, 305, 349, 343, 43, 32, 35, 38, 33, 
    337, 326, 321, 323, 317, 307, 175, 333, 223, 126, 344, 66, 50, 54, 59, 
    63, 62, 64, 59, 56, 62, 62, 73, 62, 51, 51, 52, 50, 57, 61, 60, 28, 57, 
    66, 56, 60, 48, 55, 58, 63, 47, 68, 57, 62, 7, 13, 341, 303, 316, 327, 
    316, 330, 322, 325, 308, 343, 317, 334, 327, 329, 352, 350, 357, 332, 
    338, 320, 333, 325, 327, 331, 330, 326, 318, 318, 321, 318, 315, 317, 
    314, 309, 317, 293, 123, 121, 116, 118, 127, 124, 131, 133, 124, 137, 
    124, 125, 125, 114, 121, 121, 123, 129, 131, 125, 128, 122, 123, 125, 
    128, 127, 120, 120, 125, 131, 132, 124, 127, 134, 140, 178, 0, 306, 319, 
    310, 344, 341, 330, 329, 334, 313, 323, 322, 328, 343, 332, 329, 332, 29, 
    31, 107, 146, 153, 152, 133, 112, 106, 113, 112, 124, 126, 116, 113, 114, 
    123, 120, 127, 130, 127, 123, 129, 132, 131, 127, 130, 117, 117, 118, 
    121, 120, 116, 118, 117, 120, 119, 121, 122, 118, 122, 122, 120, 125, 
    126, 125, 125, 131, 120, 124, 119, 119, 116, 115, 111, 110, 118, 125, 
    128, 150, 292, 325, 320, 298, 306, 110, 310, _, 0, 180, 63, 84, 84, 77, 
    135, _, 104, 108, 116, 106, 105, 108, 118, 111, 115, 115, 112, 103, 117, 
    83, 55, 359, 347, _, 304, 317, 302, 300, 303, 319, 316, 350, 281, 310, 
    313, 307, 268, 309, 312, 314, 320, 321, 320, 319, 315, 311, 281, 294, 
    111, 118, 135, 117, 132, 122, 131, 150, 139, 98, 145, 155, 146, 124, 117, 
    324, 307, 326, 338, 345, 63, 318, 327, 328, 320, 319, 6, 319, 325, 326, 
    329, 328, 330, 327, 328, 325, 330, 325, 326, 325, 323, 324, 322, 309, 
    301, 310, 321, 294, 318, 299, 318, 316, 319, 345, 330, 245, 302, 337, 
    348, 6, 20, 45, 48, 258, 352, 264, 247, 78, 106, 98, 310, 318, 293, 58, 
    54, 297, 272, 48, 334, 3, 10, 1, 338, 333, 333, 330, 318, 322, 335, 328, 
    323, 314, 302, 287, 288, 286, 262, 271, 286, 265, 248, _, 233, 234, 267, 
    239, 219, 204, 158, 169, 168, 153, 168, 144, 128, 114, 105, 114, 130, 
    120, 125, 133, 135, 87, 104, 132, 108, 113, 108, 103, 111, 97, 88, 97, 
    95, 75, 63, 95, 66, 64, 64, 74, 65, 39, 1, 346, 333, 353, 350, 322, 303, 
    344, 353, 4, 360, 346, 322, 355, 7, 15, 8, 344, 332, 331, 303, 304, 325, 
    318, 312, 315, 321, 319, 324, 309, 325, 305, 293, 294, 296, 289, 283, 
    282, 295, 277, 270, 270, 298, 297, 311, 300, 308, 306, 317, 331, 339, 
    348, 329, 321, 327, 350, 308, 293, 328, 328, 320, 312, 332, 320, 301, 
    337, 288, 268, 285, 250, 262, 288, 290, 251, 282, 293, 303, 308, 7, 334, 
    322, _, 0, 318, 307, 265, 285, 277, 271, 311, 324, 141, 229, 310, 304, 
    205, 335, 357, 120, 133, 122, 292, 126, 284, 0, 322, 123, 219, 295, 346, 
    294, 114, 302, 318, 303, 330, 315, 316, 308, 309, 305, 310, 318, 297, 
    295, 303, 309, 299, 303, 311, 314, 303, 299, 309, 304, 298, 297, 299, 
    298, 298, 300, 299, 296, 301, 297, 303, 307, 291, 308, 314, 288, 302, 
    304, 311, 300, 321, 306, 294, 295, 342, 36, 106, 112, 105, 106, 105, 102, 
    98, 87, 114, 111, 107, 91, 97, 93, 97, 97, 91, 90, 88, 87, 84, 88, 90, 
    83, 83, 89, 101, 113, 100, 112, 85, 75, 61, 74, 74, 53, 43, 46, 37, 45, 
    39, 38, 42, 52, _, 7, 12, 316, 330, 315, 330, 328, 317, 326, 310, 294, 
    293, 296, 297, 299, 303, 302, 301, 310, 315, 316, 314, 313, 315, 314, 
    321, 318, 312, 314, 320, 326, 328, 327, 329, 326, 324, 328, 327, 328, _, 
    327, 322, 323, 319, 329, 331, 328, 328, 329, 330, 330, 329, 328, 321, 
    324, 318, 317, 315, 313, 319, 309, 320, 311, 315, 316, 310, 312, 307, 
    308, 307, 309, 308, 312, 313, 316, 322, 319, 314, 304, 301, 305, 303, 
    306, 310, 311, 311, 313, 317, 320, 320, 320, 322, 316, 315, 319, 323, 
    307, 319, 317, 315, 319, 317, 316, 310, 281, 333, 0, 0, 125, 124, 0, 0, 
    130, 136, 131, 161, _, _, _, 122, 163, 137, 108, 175, 303, 324, 325, 320, 
    300, 316, 325, 329, 304, 300, 313, 307, 319, 322, 321, 316, 322, 299, 
    268, 266, 232, 215, 218, 218, 197, 178, 195, 230, 252, 264, 266, 292, 
    293, 283, 289, 293, 290, 269, 289, 303, 308, 319, 286, 310, 314, 318, 
    307, 314, 283, 275, 277, 291, 322, 309, 274, 281, 280, 293, 288, 298, 
    294, 299, 300, 305, 297, 301, 305, 308, 305, 303, 300, 306, 318, 319, 
    305, 300, 310, 312, 308, 308, 306, 312, 304, 327, 337, 331, 336, 322, 
    333, 320, 319, 327, 314, 328, 319, 326, 328, 333, 326, 333, 337, 319, 
    320, 329, 338, 329, 336, 331, 339, 326, 333, 333, _, 329, 331, 323, 9, 
    331, 331, 350, 322, 324, 322, 328, 336, 332, 321, 319, 299, 299, 291, 
    321, 318, 311, 300, 302, 292, 301, 313, 302, 307, 301, _, 302, 302, 319, 
    327, 316, 320, 321, 327, 324, 348, 331, 321, 330, 335, 328, 336, 320, 
    316, 269, 296, 318, 321, 116, 212, 181, 293, 313, 327, 333, 268, 279, 
    343, 184, 139, 208, 333, 307, 349, 281, 354, 50, 344, 324, 54, 49, 48, 
    52, 299, 337, 51, _, 63, 51, 49, 53, 55, _, 47, 302, 210, 341, 310, 326, 
    312, 189, 283, 324, 328, 322, 44, 38, 42, 47, 331, 51, 51, 57, 56, 53, 
    56, 52, 51, 47, 62, 65, 5, 53, 58, 61, 55, 48, 55, 56, 70, 65, 67, 78, 
    78, 80, 87, 82, 85, 86, 85, 83, 76, 72, 74, 78, 75, 72, 74, 88, _, 107, 
    104, 103, 105, 105, 110, 108, 108, _, 106, 107, 107, 111, 106, 107, 106, 
    104, 87, 78, 78, 62, 46, 247, 250, 284, 299, 294, 59, 64, 65, 66, 63, 72, 
    70, 70, 69, 71, 77, 96, 105, 107, 110, 103, 94, 87, 78, 86, 75, 78, 72, 
    69, 76, 73, 70, 82, 81, 89, 70, 68, 73, 70, 63, 59, 64, 56, 61, 66, 336, 
    320, 313, 111, 318, 319, 163, 285, 339, 313, 332, 10, 343, 348, 69, 1, 
    34, 55, 39, 51, 354, 357, 270, 298, 324, 333, 41, 346, 358, 10, 169, 333, 
    102, 325, 324, 321, 324, 320, 316, 309, 319, 327, 323, 333, 331, 325, 
    328, 320, _, 327, 316, 316, 305, 327, 319, 329, 224, 178, 164, 115, 147, 
    124, 131, 138, 129, 120, 124, 129, 132, 109, 106, 111, 111, 117, 119, 
    113, _, 116, 115, 112, 123, 107, 108, _, 297, 326, 297, 296, 300, 293, 
    299, 301, 319, 327, 325, 303, 302, 309, 302, 297, 294, 293, 299, 301, 
    299, 298, 301, 304, 305, 302, 303, 304, 306, 310, 307, 303, 294, 283, 
    288, 307, 310, 311, 314, 313, 313, 308, 314, 294, 305, 328, 302, _, 318, 
    329, 329, 319, 321, 309, 323, 307, 311, _, 296, 311, 330, 316, 321, 301, 
    338, 356, 321, 151, 102, 357, 120, 119, 104, 104, _, 111, 109, 122, 111, 
    113, 122, 109, 100, 97, 82, 75, 74, 74, 65, 67, 142, 96, 97, 88, 94, 106, 
    112, 107, 113, 112, 122, 107, 111, 102, 103, 97, 99, 92, 92, 96, 89, 73, 
    90, 85, 79, 74, 82, 70, 96, 88, 80, 65, 53, 60, 83, 72, 85, 54, 14, 58, 
    57, 65, 54, 55, 60, 59, 351, 284, 291, 353, 320, 320, 308, 324, 309, 313, 
    321, 322, 311, 311, 319, 319, 325, 315, 325, 325, 323, 322, 319, 321, 
    326, 326, 315, 311, 304, 308, 304, 307, 309, 308, 304, 309, 304, 305, 
    306, 310, 314, 311, 309, 310, 314, 311, 311, 313, 314, 318, 317, 318, 
    324, _, 316, 313, 307, 311, 306, 318, 303, 325, 306, _, 135, 113, 139, 
    114, 7, 4, 310, 224, 253, 266, 315, 301, 270, 273, 307, 313, 322, 317, 
    320, 302, 306, 316, 307, 315, 320, 325, 318, 313, 314, 314, 316, 266, 12, 
    116, 105, 82, 133, 137, 142, 138, 102, 101, 107, 95, 79, 67, 89, 271, 
    322, 78, 146, 130, 122, 132, 117, 140, 126, 110, 93, 83, 86, 126, 95, 90, 
    107, 90, 80, 76, 85, 93, 107, 108, 106, 101, 108, 111, 108, 100, 102, 
    101, 94, 89, 97, 104, 110, 101, 128, 111, 88, _, 115, 169, 224, 261, 290, 
    300, 298, 297, 347, 303, 317, 344, 315, 317, 321, 325, 322, 322, 318, 
    322, 315, 333, 315, 322, 322, 323, 320, 324, 307, 325, 322, 312, 69, 116, 
    162, 183, 158, 83, 88, 136, 15, 342, 337, 328, 298, 278, 302, 266, 284, 
    318, 315, 336, 332, 325, 317, 329, 324, 322, 319, 318, 313, 310, 315, 
    313, 312, 317, 315, 316, 317, 317, 314, 312, 308, 312, 309, 308, 313, 
    318, 293, 290, 276, 279, 290, 314, 281, 317, 295, 294, 286, 276, 294, 
    313, 309, 315, 320, 320, 325, 331, 326, 333, 324, 316, 295, 310, 316, 
    318, 306, 313, 315, 321, 320, 321, 318, 311, 295, 316, 281, 294, 308, 
    311, 322, 317, 319, 311, 312, 298, 316, 318, 315, 321, 328, 313, 315, 
    320, 320, 318, 314, 320, 313, 310, 311, 304, 307, 303, 308, 308, 311, 
    314, 314, 314, 315, 314, 312, 305, 314, 313, 313, 313, 329, _, 323, 327, 
    326, 326, 320, 325, 325, 323, 316, 325, 329, 329, 330, 328, 329, 317, 
    312, 321, 322, 324, 311, 213, 351, 325, 328, 327, 332, 316, 336, 282, 
    332, 144, 0, 154, 133, 128, 123, 134, 122, 118, 116, 115, 110, 109, 109, 
    111, 122, 274, 294, 302, 307, 302, 296, 292, 298, 292, 293, 296, 286, 
    278, 281, 284, _, 293, 291, 295, 296, 299, 301, 296, 319, 311, 323, 325, 
    329, 319, 315, 318, 310, 303, _, _, 310, 311, 307, 309, 313, 320, 320, 
    326, 333, 327, 324, 335, 336, 330, 332, 336, 336, 338, 347, 349, 348, 
    335, 342, 341, 332, 333, 325, 324, 331, 337, 334, 332, 331, 347, 20, 41, 
    48, 38, 30, 13, 38, 51, 352, 29, 37, 24, 30, 47, 48, 53, _, 63, 67, 84, 
    85, 94, 82, 69, 321, 276, 337, 56, 358, 57, _, 354, 32, 45, 51, 26, 15, 
    35, 354, 304, 300, 254, 244, 215, 201, 174, 182, 140, 82, 129, 149, 183, 
    210, 331, 313, _, 272, 267, 279, 293, 311, 263, 203, 212, 183, 199, 186, 
    171, 161, 151, 149, 127, 162, 164, 172, 178, 159, 163, 174, 170, 173, 
    149, 141, 175, 147, 106, 87, 95, 105, 116, _, 117, 119, 113, 107, 116, 
    108, 114, 108, 108, 125, 113, 141, 130, 129, 116, 120, 133, 125, 133, 
    136, 127, 139, 130, 126, 128, 130, 128, 124, 121, 117, 116, 119, 113, 
    117, 116, 117, _, 102, 105, 110, 113, 115, 122, 123, 126, 133, 133, 125, 
    120, 115, 117, 121, 120, 127, 120, _, 122, 116, 107, 83, 83, 102, 90, 89, 
    81, 93, 103, 105, 101, 100, 98, 100, 107, 107, 114, 114, 113, 113, 113, 
    113, 117, 111, 123, 120, 102, 114, 113, 129, 114, 113, 125, 116, 118, 
    115, 112, 115, _, 121, 112, 123, 156, 124, 95, 102, 134, 49, 118, 109, 
    119, 108, 115, 97, 93, 96, 91, 102, 107, 118, 119, 99, 103, 104, 100, 
    105, 108, 104, 117, _, 116, 115, 109, 109, 126, 118, 135, 110, 121, 139, 
    136, 124, 137, _, 181, 177, 168, 85, 138, 148, 161, 115, 142, 130, 121, 
    113, 121, 118, 109, 115, 113, 108, 110, 108, 107, 97, 97, 104, 105, 110, 
    114, 115, 115, 114, 112, 117, 109, 107, 99, 108, 30, 355, _, 316, 7, 21, 
    323, 124, 325, 116, 258, 300, 317, 233, 57, 65, 67, 74, 81, 88, 98, _, 
    100, 109, 118, 120, 115, 110, 100, 107, 102, 104, 112, 107, 109, 111, 
    112, 108, 104, 106, 94, 97, 98, 103, 100, 98, 99, 95, 97, 91, 102, 101, 
    103, 97, 94, 113, 109, 97, 93, 122, 78, 309, 319, 347, 358, 312, 312, 
    318, 325, 321, 321, 315, 313, 318, 311, 339, 323, 330, 297, 312, 310, 
    331, 59, 66, 60, 58, 57, 69, 61, 67, 70, 66, 68, 78, 71, 71, 61, _, 75, 
    80, 84, 79, 80, 71, 72, 75, 72, 81, 68, 49, 57, 53, 38, 41, 52, 360, 328, 
    353, 5, 54, 310, 12, 45, 56, 54, 199, 288, 257, 260, 227, 289, 37, 351, 
    8, 51, 64, 324, 322, 86, 224, 111, 326, 49, 42, 54, 53, 47, 332, 28, 305, 
    46, 52, 43, 324, 40, 269, 335, 278, 0, _, 339, 315, 342, 323, 322, 317, 
    324, 329, 323, 325, 324, 308, 311, 312, 313, 315, 312, 306, 311, 309, 
    314, 310, 310, 307, 305, 312, 314, 309, 316, 320, 324, 320, 315, 311, 
    327, _, 88, 112, 116, 92, 95, 114, 109, 117, 116, 112, 121, 121, 119, 
    115, 108, 108, 103, 121, 110, 121, 113, 112, 113, 106, 106, 101, 107, 
    103, 107, 111, 117, 111, 113, 105, 105, 103, 105, 109, 108, 118, 103, 
    103, 108, 111, 106, 112, 105, 108, 106, 110, 105, 107, 96, 101, 101, 99, 
    98, 100, 91, 94, 85, 86, 77, 72, 68, 84, 93, 75, 77, 67, 58, 65, 71, 67, 
    69, 73, 75, 82, 70, 72, 77, _, _, 71, _, 59, 67, 81, 83, 86, 93, 85, 92, 
    97, 89, 92, 69, 76, 82, 82, 80, 75, 79, 80, 83, 84, 86, 84, _, 86, 89, 
    87, 85, 86, 84, 82, 83, _, 82, 82, 82, 82, 82, 76, 82, 71, 75, 74, 77, 
    71, 74, 73, 67, 59, 67, 73, 63, 65, 64, 60, 64, 67, 61, 62, 63, 65, 62, 
    62, 64, 74, 77, 73, 75, 74, 71, _, 66, 69, 67, 63, 65, 64, 67, 70, 77, 
    76, 69, 64, 69, 73, 74, 80, 64, 67, 61, 206, 65, 56, 59, 59, 58, 59, 57, 
    65, 63, 70, 68, 137, 322, 308, 147, 171, 26, 11, 49, 52, 15, 28, 29, 22, 
    25, 17, 29, 34, 25, 356, 23, 14, 7, 9, 29, 4, 354, 10, 358, 343, 348, 
    353, 337, 316, 297, 306, 330, 334, 38, 35, 28, _, 21, 29, 312, 350, 351, 
    357, 346, 335, 346, 329, 330, 336, 331, 325, 330, 324, 326, _, 311, 326, 
    321, 319, 318, 322, 325, 327, 324, 319, 320, 319, 320, 319, 320, 312, 
    310, 324, 326, 314, 316, 318, 316, 309, 318, 311, 333, 329, 320, 331, 
    319, 317, 322, 315, 337, 322, 324, 328, 343, 343, 335, 334, 8, 347, 330, 
    300, 15, 324, 17, 15, 360, 5, 36, _, 347, 75, 66, 73, 65, 85, 89, 118, 
    123, 117, 148, 148, 150, 168, 152, 153, 144, _, 144, 143, 128, _, 126, 
    189, 249, 274, 276, 288, 284, 293, 293, 298, 297, 298, 295, 293, 302, _, 
    275, 285, 259, 273, 257, 231, 245, 238, 236, 204, 207, 196, 188, 205, 
    214, 194, 203, 203, 202, 184, 193, 182, 207, 165, 196, 182, 189, 150, 
    113, 136, 117, 124, 76, _, 354, 358, 1, 354, 354, _, 347, 338, 344, 354, 
    338, 353, 316, 316, 315, 318, 324, 327, 320, 316, 311, 312, 300, 308, 
    304, 308, 337, 342, 282, 289, 276, 274, 258, 257, 270, 270, 296, 280, 
    292, 288, 268, 266, 278, 316, 269, 294, 268, 261, 258, 264, 254, 254, 
    260, 257, 272, 262, 255, 238, 237, 225, 219, 215, 220, _, 250, 285, 256, 
    258, 210, 205, 199, _, 218, 219, 233, 229, 229, _, 227, 218, 234, 214, 
    217, 215, 192, 179, 108, 107, 151, 136, 131, 137, 120, 112, 119, 112, 
    109, 124, 115, 128, 122, 116, 118, 118, 110, 109, _, 110, 101, 105, 116, 
    114, 102, 101, 90, 83, 91, 84, 63, 44, 53, 36, 46, 46, 47, 51, 51, 50, 
    43, 56, 56, 66, 70, 68, 65, 73, 329, 50, 44, 40, 25, 20, 14, 13, 1, 355, 
    355, 345, 345, 333, 332, 334, 342, 340, 329, 333, 333, 335, 350, 339, 
    342, 347, 339, 336, 340, 346, 334, 339, 353, 1, 4, 22, 24, 67, 31, 22, 
    88, 71, 65, 63, 49, 99, 46, 43, 344, 114, 84, 94, 96, 102, 116, 121, 120, 
    112, 121, 114, 118, 113, 114, 129, 133, 137, 135, 140, 147, 142, 141, 
    142, 168, 155, 164, 196, 292, 265, 275, 260, 266, 297, 309, 312, 312, 
    313, 312, 310, 315, 307, 314, 316, 308, 310, 308, 331, 316, 324, 326, 
    314, 316, 356, 345, 26, _, 43, 65, 84, 60, 75, 80, 67, 67, 72, 78, 82, 
    77, 81, 100, 156, 153, 194, 198, 192, 176, 161, 205, 207, 196, 219, 230, 
    192, 205, 187, 210, 194, 190, 125, 168, 153, 143, 142, 162, 163, 177, 
    196, 177, 172, 160, 149, 146, 153, 141, 141, 141, 142, 141, 144, 140, 
    139, 144, 122, 129, 140, 139, 139, 133, 136, 136, 130, 131, 134, 130, 
    129, 126, 126, 124, 124, 128, 124, _, 128, 129, 126, 126, 126, 130, 129, 
    133, 133, 133, 131, 131, 131, 128, 117, 125, 119, 121, 124, 118, 120, 
    126, 113, 107, 102, 107, 114, 106, 86, 84, 83, 87, 93, _, 105, 116, 217, 
    294, 301, 307, 309, 318, 310, 313, 306, 309, 301, 307, 305, 297, 293, 
    308, 304, 308, 320, 360, 15, 340, 317, 6, _, 96, 105, 163, 166, 158, 161, 
    168, 169, 190, 198, 202, 203, 204, 187, 187, 181, 186, 181, 187, 181, 
    193, 195, 184, 184, 187, 176, 174, 193, 205, 239, 254, 280, 279, _, 299, 
    302, 280, 279, 275, 303, 97, 79, 121, 104, 126, 115, 133, 144, 125, 142, 
    132, 171, 157, 185, 100, 119, 113, 124, 108, 101, 107, 86, 125, 117, 76, 
    87, 75, 73, 92, 80, 118, 99, 95, 101, 110, 117, 117, 117, 119, 134, 134, 
    146, 126, 119, 145, 139, 130, 138, 125, 128, 126, 127, 122, 118, 119, 
    120, 110, 104, 94, 101, 106, 103, 87, 94, 97, 85, 88, 83, 68, 64, 61, 54, 
    56, 67, 71, 62, 57, 64, 68, 71, 64, 62, 63, 60, 64, 65, 66, 86, 71, 60, 
    60, 50, 50, 47, 51, 52, 51, 44, 52, 46, 51, 51, 56, 43, 290, 20, 16, 325, 
    304, 48, 27, 39, 34, 21, 311, 305, 294, 224, _, 325, 48, 67, 51, 353, 62, 
    64, 70, 60, 63, 60, 60, 59, 56, 57, 55, 50, 50, 46, 298, 299, 320, 334, 
    0, 21, 13, 21, 328, 354, 170, 267, 15, 169, 61, 46, 339, 43, 40, 318, 
    315, 332, 20, 26, 27, 44, 44, 51, 33, 32, 39, 28, 39, 30, 43, 31, 4, 33, 
    3, 33, 22, 19, 9, 354, 1, 10, 43, 40, 50, 40, 49, 48, 48, 60, 49, 53, 48, 
    49, 50, 52, 46, 41, 43, 39, 30, 31, 43, 40, 35, 33, 48, 36, 26, 17, 21, 
    3, 4, 359, 358, 348, 345, 339, 337, 333, 331, 326, 325, 328, 320, 316, 
    314, 311, 313, 314, 313, 308, 310, 309, 303, 306, 293, 297, 291, 301, 
    293, 289, 293, 283, 270, 260, 270, 242, 241, 233, 229, 229, 220, 210, 
    227, 216, 209, 212, 217, 227, 231, 232, 224, 257, 283, 300, _, 292, 292, 
    287, 268, 259, 264, 267, 265, 305, 341, 337, 357, 8, 20, 14, 9, 6, 1, 1, 
    7, 11, 1, 355, 3, 24, 27, 12, 11, 4, 12, 21, 13, 31, 34, 24, 13, 8, 16, 
    343, 3, 356, 3, 360, _, 7, 1, 3, 1, 19, 14, 360, 24, 355, 3, 329, 310, 
    342, 328, 314, 314, 318, _, 301, 337, 319, 321, 341, 11, 17, 7, 30, _, 
    19, 355, 352, 330, 326, 328, 340, 329, 326, 332, 328, 327, 332, 337, 334, 
    332, 332, 335, 331, 335, 340, 338, 337, 334, 322, 352, 5, 14, 25, _, _, 
    53, 43, 39, _, _, _, 55, 53, 52, _, 31, 37, 10, 54, 57, 57, 69, 67, 60, 
    49, 70, 66, 61, 65, 55, 84, 71, 83, _, 79, 54, 60, 65, 61, 51, 55, 60, 
    48, 56, 45, 45, 65, 60, 58, 61, 61, 61, 67, 82, 81, 84, 102, 98, 81, 76, 
    76, 80, 94, 95, 104, 105, 105, 100, 96, 95, 97, 100, 102, 97, 97, 102, 
    101, _, 95, 95, 99, 99, 100, 99, 103, 99, 103, 105, 107, 109, 107, 114, 
    108, 101, 115, 109, 122, 109, 115, 123, 134, 132, 119, 126, 127, 123, 
    127, 118, 104, 103, 113, 125, 120, 118, _, 115, 111, 112, 116, 116, 132, 
    137, 134, 138, 138, 125, 138, 119, 116, 112, 116, 115, 110, 114, 116, 
    109, 91, 89, 104, 115, 108, 118, 128, 143, 151, 154, 152, 135, 121, 124, 
    _, 137, 128, _, 136, 171, 194, 217, 270, 288, 291, 294, 296, 298, 304, 
    306, 316, 320, 324, 327, 333, 341, 346, 346, 351, 356, 9, 5, 2, 360, 360, 
    358, 352, 355, 353, 350, 354, 343, 343, 338, 334, 331, 333, 333, 331, 
    332, 330, 324, 334, 333, 333, _, 338, 340, 339, 339, 345, 337, _, 338, 
    338, 339, 338, 340, 342, 337, 335, 336, 336, 334, _, _, 329, 327, 328, 
    324, 325, 322, 319, 319, 318, 316, 315, 316, 316, 319, 319, 315, 316, 
    315, 314, 310, 317, 316, 312, 315, 318, _, 311, 311, 311, 310, 310, 308, 
    309, 308, 304, 306, 300, 301, 303, 299, 299, 292, 290, 289, 285, 292, 
    279, 284, 279, 268, 262, 264, 250, 241, 222, 235, 230, 222, 226, 228, 
    221, 224, _, 214, 214, 220, 225, 227, 222, 228, 230, _, 219, 224, 220, 
    212, 195, 179, 186, 162, 149, 151, 156, 153, 138, 152, 148, 129, 95, 64, 
    31, 15, 26, _, 10, 20, 22, _, 18, 28, 29, 25, 23, 15, 16, 25, 349, 309, 
    330, 4, 22, 6, 334, 335, 338, 344, 344, 356, 350, 340, 342, 346, 325, 
    323, 326, 321, 316, 309, 308, 314, 313, 313, 323, 315, 318, 309, 320, 
    319, 333, 322, 322, 321, 325, _, 332, 334, 3, 34, 24, _, 20, 20, 23, 30, 
    31, 34, 30, 35, 40, 42, 32, 19, 16, 13, 13, 6, 354, 1, 360, _, 1, 11, 10, 
    355, 4, 7, 32, 41, 37, 27, 50, 48, 33, 41, 12, 52, 32, 54, 42, 36, 61, 
    63, 64, 7, 61, 62, 57, 56, 57, 57, 50, 30, 25, 20, 45, 53, 56, 57, 48, 
    48, 49, 47, 49, 54, 53, 49, 50, 50, 46, _, 41, 36, 32, 30, 33, 33, 35, 
    40, 29, 40, 37, 36, 34, 34, 45, 29, 36, 38, 51, 59, 67, _, 66, 67, 62, 
    67, 64, 86, 85, 90, 87, 96, 86, 97, 87, 89, 98, 92, 107, 105, 104, 105, 
    103, 96, 90, 89, 94, 319, 3, 340, 342, 337, 341, 344, 331, 325, 316, 324, 
    327, 314, 308, 309, 294, 305, 307, 306, 312, 304, _, 300, 295, 291, 283, 
    283, 282, 297, 311, 306, 310, 317, 321, 311, 314, 311, 302, 301, 304, 
    304, 309, 316, 323, 298, 316, 296, 292, 290, 3, 26, 348, 342, 4, 24, 51, 
    51, 43, 45, 51, 45, 47, 41, 36, 37, 43, 39, 22, 5, 358, 11, 11, 349, 1, 
    352, 282, 311, 343, 310, 307, 301, 278, 286, 297, 302, _, _, _, _, _, _, 
    _, _, _, 295, 299, 302, 301, 311, 303, 307, 307, 298, 311, 315, 304, 319, 
    313, 311, 305, 321, 309, 291, 302, 326, 312, 321, 326, _, 338, 355, 5, 
    26, 2, 30, 71, 78, 79, 83, 82, 81, 77, 79, 80, 81, 85, 97, 104, 106, 112, 
    112, 112, 112, 111, 108, 107, 118, 117, 127, 112, 128, 120, 126, 118, 
    116, 112, 106, 104, 102, 98, 97, 90, 92, 91, 90, 88, 89, 90, 82, 63, 67, 
    49, 55, 60, 46, 49, 46, 40, 53, 51, 57, 37, 43, 39, 28, 16, 15, 11, 16, 
    3, 27, 348, 18, 56, 14, 3, 22, 21, 33, 28, 14, 25, 56, 54, 34, 24, 59, 
    85, 69, 78, 64, 71, 62, 60, 69, 61, 73, 65, 56, 45, 38, 51, 30, 26, 24, 
    15, 22, 32, 63, 62, 61, 17, 18, 10, 14, 343, 11, 6, 14, 13, 18, 11, 23, 
    11, 10, 69, 89, 89, 81, 73, 63, 51, 53, 55, 65, 72, 87, 74, 77, 84, 117, 
    113, _, 131, 98, 146, 115, 114, 106, 132, 126, 147, 122, 125, 143, 135, 
    147, 159, 148, 146, 161, 184, 160, 180, 177, 174, 108, 112, 124, 127, 
    121, 128, 138, 141, 150, 162, 152, _, 134, 126, 104, 111, 84, 87, 101, 
    93, 91, 87, 89, 78, 78, 81, 122, 99, 114, 120, 115, 119, 117, 182, 170, 
    165, 163, 151, 167, 177, 182, 208, 227, 247, 344, 331, 42, 9, _, 19, 17, 
    19, 30, 351, 19, 3, 2, 16, 12, 35, 12, 111, 11, 46, 22, 21, 44, 26, 27, 
    15, 338, 337, 351, 1, 355, 8, 20, 357, 343, 329, 302, 311, 318, _, 310, 
    322, 321, 318, 323, 320, 321, 323, 327, 335, 345, 338, 36, 47, 49, 57, 
    50, 44, 40, 40, 42, 58, 54, 50, 53, 56, 56, 52, 59, 58, 58, _, 51, 51, 
    48, 48, 49, 50, 50, 53, 50, 45, 47, 47, 55, 53, 53, 59, 55, 51, 54, 53, 
    55, 53, 128, 55, 53, 57, 53, 51, 53, 57, 64, 60, 60, 59, 56, 57, 58, 60, 
    _, _, 62, 59, 55, 51, 52, 55, 57, 54, 59, 64, 125, 102, 96, 104, 108, 
    112, 107, 118, 102, 110, 108, 103, 130, 109, 106, 94, 93, 85, 85, 69, 69, 
    64, 90, 110, 107, 105, 104, 107, 109, 109, 114, 123, 133, 138, 142, 141, 
    137, 139, 138, 136, 135, 131, 135, 138, 137, 134, 147, 146, 138, 151, 
    153, 156, 157, 157, 144, 147, 142, 141, 136, 130, 131, 133, 125, 141, 
    136, 134, 133, 130, 135, 136, 149, 147, 151, 151, 154, 156, 155, 156, 
    161, 153, 149, 149, 150, 146, 141, _, 149, 145, 146, 152, 146, 144, 143, 
    143, 140, 135, 141, 136, 134, 140, 138, 138, 134, 134, 122, 133, 132, 
    141, _, 154, 146, 156, 158, 158, 155, 170, 168, 160, 156, 150, 144, 142, 
    147, 173, 153, 147, 152, 153, 171, 172, 158, 170, 173, 170, 155, 160, 
    179, 190, 205, 199, 191, 195, 198, 196, 194, 188, 185, 176, 191, 185, 
    197, _, 137, 161, 156, 156, 129, 142, 134, 121, 104, 96, 109, 138, 139, 
    141, 146, 152, 142, 128, 129, 141, 146, 150, 134, 146, 150, 154, 157, 
    165, 184, _, 268, 256, 259, 265, 262, 257, 232, 252, 282, 296, 315, 316, 
    319, 321, 330, 329, 323, 329, 336, 347, 348, 346, 348, 349, 345, 345, 
    340, 327, 319, 321, 311, 312, 311, 318, 330, 319, 313, 320, 315, 328, 
    343, 328, 344, 348, 334, 360, 354, 11, 27, 40, 44, 48, 56, 71, 67, 59, 
    93, 151, 152, 147, 153, 151, 158, 160, 162, 161, 162, 159, 173, 177, 181, 
    187, 267, 253, 269, 278, 276, 273, 272, _, 310, 304, 311, 325, 324, 327, 
    317, 331, 324, 323, 321, 328, 324, 337, 315, 294, 307, 300, 282, 305, 
    315, 321, 330, 326, 334, 352, 18, 34, 40, 40, 47, 41, 47, 67, 72, 85, 84, 
    95, 91, 83, 88, 92, 90, 90, 88, 91, 88, 90, 91, 95, _, 103, 123, 240, 
    273, 278, 291, 291, 289, 291, 287, 269, 256, 250, 246, 241, 247, 261, 
    280, 311, 287, 311, 336, 343, 344, 345, 348, 348, 341, 339, 344, 343, 
    340, 333, 322, 332, 337, 336, 333, 334, 325, 336, 349, 341, 349, 342, 
    353, 350, 357, 355, 356, 329, 313, 296, 308, 299, 288, 284, 262, 283, 
    289, _, 290, 304, 306, 301, 303, 302, 298, 288, 290, _, 281, 282, 276, 
    284, 280, 285, _, 289, 285, 301, 285, 269, 317, 319, 325, 16, 17, 24, 9, 
    _, 23, 20, 19, 348, 329, 2, 21, 79, 69, 47, 32, 39, 33, 44, 29, 26, 22, 
    13, 17, 42, 49, 53, 46, 35, 29, 30, 2, 4, 350, 4, 44, 102, 105, 103, 101, 
    104, 124, 130, 160, 144, 144, 140, 146, 151, 154, 144, 169, 69, 64, 74, 
    79, 57, 71, 56, 58, 39, 25, 4, 1, 2, 358, 261, 270, 12, 11, 359, 3, 1, 
    359, 359, 5, 355, 352, 4, 2, 8, 3, 18, 24, 47, 32, 30, 57, 67, 83, 80, 
    93, 87, 91, 98, 99, 104, 110, 110, 107, 107, 110, 109, 109, 111, 113, 
    113, 112, 112, 110, 111, 106, 108, 106, 103, 103, 164, 144, 147, 156, 
    155, 154, 154, 157, 145, 113, 105, 102, 113, 116, 114, 111, 97, 106, 100, 
    110, 107, 106, 108, 113, 117, 114, 110, 109, 112, 109, 113, 114, 110, 
    112, 110, 103, 96, 97, 103, 103, 106, 109, 105, 101, 103, 99, 93, 93, 92, 
    94, 98, 98, 98, 97, 96, 93, _, _, 88, 87, 87, 88, 85, 82, 82, 81, 86, 88, 
    91, 91, 90, 89, 87, 87, 85, 84, 85, 85, 83, 83, 83, 82, 81, _, _, _, 80, 
    74, 74, 75, 76, 80, 81, 77, 75, 73, 71, 75, 76, 78, 81, 87, 87, 88, 89, 
    90, 90, 89, 87, 94, 93, 96, 102, 99, 96, 94, 95, 96, 95, 78, 96, 91, 74, 
    73, 78, 73, 69, 78, 91, _, 85, 61, 69, 65, 43, 42, 39, 31, 41, 47, 59, 
    55, 55, 63, 55, 53, 53, 51, 55, 56, 50, 48, 74, 83, _, 82, 87, 84, 101, 
    97, 120, 119, 93, 88, 99, 98, 107, 94, 107, 125, 127, 134, 123, 132, 125, 
    119, 121, 123, 124, 113, 117, 122, 117, 116, 114, 109, 109, 111, 112, 
    113, 112, 112, 111, 108, 108, 110, 107, 109, 114, 116, 117, _, 116, 116, 
    116, 116, 114, 113, 115, 122, 178, 105, 195, 116, 114, 111, 170, 109, 
    120, 113, 101, 97, 98, 97, 117, 153, _, 126, 115, 108, 89, 91, 114, 3, 
    357, 303, 296, 301, 293, 299, 296, 292, 292, 293, 292, 313, 301, 296, 
    306, 308, 301, 313, 300, 301, 289, 293, 297, 291, 295, 314, 305, 303, 
    279, 292, 224, 189, 148, 153, 181, 185, 176, 171, 168, 144, 221, 237, 
    236, 239, 240, 225, 231, 231, 217, 213, 221, 224, 255, 264, 281, 298, 
    281, 281, 273, 319, 60, 69, _, 68, _, 78, 81, 80, 88, 98, 98, 280, 301, 
    292, 297, 309, 308, 62, 56, 44, 45, 35, 21, 5, 357, 339, 341, 336, 330, 
    333, 334, 326, 319, 319, 314, 315, 306, 314, 311, 311, 314, 313, 317, 
    319, 319, 318, 312, 315, 308, 311, 315, _, 318, 320, 318, 317, 325, 331, 
    335, 333, 325, 327, 331, 341, 347, 345, 352, 3, 354, 16, 360, 8, 7, 24, 
    23, 21, 11, 17, 11, 24, 43, 42, 32, 39, 33, 34, 34, 28, 36, 27, 43, 48, 
    49, 50, 33, 34, 33, 34, 29, 33, 73, 82, 75, 74, 77, 86, 87, 88, 82, 85, 
    96, 98, 102, 102, 103, 102, 100, 99, 101, 96, 96, 94, 88, 81, 87, 91, 90, 
    101, 85, 97, 88, 92, 81, 94, 96, 101, 94, 100, 89, 91, 85, 73, 71, 72, 
    65, 65, 63, 63, 61, 61, 48, 49, 49, 56, 58, 62, 62, 60, 59, 60, 61, 60, 
    64, 67, 67, 70, 65, 75, 73, 64, 63, 53, 54, 52, 51, 45, 40, 34, 32, 38, 
    52, 53, 48, _, 53, 52, 54, 51, 56, 61, 42, 16, 24, 35, 37, 18, 23, 30, 
    41, 19, 20, 14, 30, 25, 39, 40, 33, 41, 48, 39, 26, 29, 57, 74, 83, 81, 
    84, 82, 80, 85, 79, 87, 96, 91, 106, 99, 104, 100, 98, 101, 94, 88, 88, 
    79, _, 64, 64, 62, 60, 59, 57, 58, 58, 56, 49, 49, 39, 35, 30, 33, 29, 
    21, 17, _, _, _, 22, 15, 16, 11, 10, 7, 10, 3, 4, 354, 357, 354, 358, 
    354, 355, 356, 1, 356, 360, 1, 360, 355, 357, 355, 2, 9, 13, 19, 10, 9, 
    33, 45, 50, 50, 42, 51, 52, 52, 37, 44, 52, 55, 47, 41, 45, 37, 35, 37, 
    39, 42, 9, 8, 36, 46, 36, 13, 3, 25, 28, 24, 36, 35, 15, 18, 16, 12, 17, 
    15, 3, 3, 4, _, 53, 56, 41, 42, 40, 38, 22, 28, 296, 53, 21, 65, 120, 
    346, 48, 15, 15, 12, 8, 29, 47, 42, 58, 33, 35, 32, 18, 18, 23, 35, 347, 
    283, 251, 318, 309, 297, 355, 27, 18, 258, 57, 78, 292, 51, 15, 28, 27, 
    26, 19, 23, 25, 5, 13, 14, 20, 28, 41, 36, 38, 53, 53, 47, 61, 28, 17, 
    14, _, 5, 15, 21, 20, 36, 50, 25, 39, 49, 68, 79, 48, 26, 44, 58, 27, 9, 
    37, 40, 41, 35, 39, 50, 35, 47, 54, 69, 70, 72, 63, 72, 92, 83, 107, 93, 
    98, 103, 116, 107, 99, 76, 54, 50, 53, 52, 46, 41, 41, 50, 46, 57, 51, 
    52, 35, 45, 48, 46, 49, _, _, _, 27, 33, 33, 45, 75, 316, 318, 325, 51, 
    51, 53, 51, 59, 346, 50, 49, 92, 152, 86, 32, 354, 340, 310, 36, 37, 42, 
    47, 47, 47, 359, 51, 65, 71, 71, 63, 55, 46, 56, 52, 57, 49, 44, 48, 48, 
    42, 44, 47, 44, 44, 48, 56, 49, 51, 45, 48, 40, 44, 34, 24, 31, 36, 39, 
    37, 29, 55, 44, 46, 41, 37, 40, 40, 44, 43, 39, 41, 45, 38, 45, 48, 47, 
    46, 49, 46, 45, 46, 51, 52, _, 41, 46, 48, 51, 55, 50, 48, 51, 51, 52, 
    51, 47, 39, 42, 47, 51, 51, 49, 337, 32, 66, 55, 325, 97, 61, 67, 76, 75, 
    68, 71, 83, 75, 76, 77, 78, 81, 76, 71, 82, 70, 64, 54, 51, 55, 60, 62, 
    57, 58, 54, 56, 63, 68, 64, 62, 63, 60, 61, 49, 57, 49, 51, 48, 54, 57, 
    59, 54, 56, 54, 54, 64, 65, 55, 61, 68, 61, 62, 65, 64, 60, 56, 58, 60, 
    56, 61, 64, 69, 60, 68, 78, 79, 142, 79, 75, 84, 77, 97, 96, 110, 111, 
    114, 108, 103, 116, 124, 92, _, 101, 104, 104, 102, 99, 107, 110, 120, 
    111, 127, 127, 127, 120, 115, 121, 115, 117, 116, 111, _, 117, 132, 110, 
    115, 111, 114, 117, 111, 113, 116, 119, 115, 115, 113, 117, 125, 120, 
    117, 117, 121, 122, 124, 118, 121, 115, 117, 130, 127, 152, 143, 146, 
    163, 147, 127, 147, 151, 142, 140, 134, 128, 132, 172, 166, 120, 117, 
    116, 132, 146, 134, 130, 136, 119, 308, 331, 321, 320, 308, 319, 306, 
    292, 358, 0, 48, 105, 118, 138, 128, 109, 109, 112, 101, 111, 121, 284, 
    301, 300, 289, 297, 297, 309, 304, 299, 295, 295, 295, 307, 303, 298, 
    309, 304, 301, 261, 247, 227, 219, 198, 213, 281, 305, 328, 319, 332, 
    337, 328, 333, 324, 336, 79, 101, 105, 109, 283, 283, 297, 293, 293, 297, 
    282, 122, 149, 135, 120, 110, _, 106, 124, 120, 111, 114, 115, 109, 118, 
    145, 133, 127, 116, 108, 107, 110, 121, 126, 114, 117, 114, 102, 90, 44, 
    18, 136, 121, 102, 93, 51, 53, 61, 55, 59, 59, 65, 70, 56, 63, 69, 67, 
    64, 58, 54, _, 56, 54, 315, 330, 286, 308, 313, 283, 288, 294, 304, 298, 
    293, 298, 298, 299, 300, 297, 306, 299, 301, 301, 310, 316, 317, 320, 
    320, 319, 314, _, 330, 359, 2, 1, 356, 1, 5, 359, 359, 345, 1, 11, 7, 10, 
    14, 90, _, 92, 112, 105, 127, 146, 154, 134, 143, 155, 143, 143, 121, 
    132, 133, 122, 120, 112, 118, 121, 131, 130, 129, 134, 344, 355, 4, 360, 
    340, 330, 330, 353, 352, 2, 6, 15, 24, 22, 24, 22, 19, 359, 9, 10, 15, 
    109, 52, 37, 33, 72, 63, 62, 61, 67, 91, 85, 104, 111, 112, 111, 116, 
    101, 93, 309, 319, 322, 331, 336, 343, 4, 27, 19, 30, 37, 12, 20, 9, 13, 
    18, 17, 22, 19, 59, 59, 54, 53, 57, 51, 51, 51, 50, 49, 46, 45, 52, 49, 
    _, 11, 6, 360, 359, 353, 347, 346, 339, 337, 338, 334, 346, 340, 333, 
    334, 333, 334, 335, 331, 331, 330, 328, 327, 325, 327, 329, 351, 352, 
    355, 353, 351, 337, 318, 335, 345, 343, 12, 27, 360, 4, 31, 16, 21, 4, 
    11, 352, 351, 1, 346, 340, 337, 352, 333, 287, 291, 325, 288, 300, 318, 
    336, 333, 330, 324, 328, 328, 326, 329, 329, 341, 319, 340, 339, 351, 
    341, 338, 333, 340, 335, 331, 317, 322, _, 313, 332, 332, 327, 330, 333, 
    324, 324, 331, 328, 334, 333, 334, 354, 350, 344, 344, 342, 341, 352, 16, 
    18, 6, 61, 75, 59, 56, 75, 91, 84, 70, 60, 58, 50, 51, 47, 49, 53, 51, _, 
    54, 56, 30, 52, 70, 53, 26, 18, _, 37, 3, 355, 5, 17, 23, 59, 61, 57, 76, 
    86, 91, 97, _, _, 104, 104, 99, 93, 88, 84, 79, 69, 71, 68, 71, 71, 100, 
    52, 59, 65, 13, 32, 20, 35, 31, 51, 13, 26, 71, 47, 6, 8, 86, 34, 15, 
    318, 344, 29, 293, 296, 31, 13, 64, 301, 323, 334, 325, 98, 5, 346, 51, 
    2, 42, 60, 111, 63, 63, 75, 78, 83, 86, 87, 86, 98, 101, 111, 98, 94, 92, 
    97, 100, 95, 95, 94, 101, 130, 103, 99, 101, 100, 104, 98, 99, 102, 103, 
    108, 107, 107, 99, 102, 107, 103, 97, 96, 99, 99, 99, 91, 97, 95, 163, 
    97, 96, 90, 73, 59, 66, 50, 51, 54, 54, 46, 28, 13, 6, 7, 1, 3, 358, 18, 
    12, 352, 353, 350, 353, 347, 345, 345, 350, 352, 339, 343, 18, 339, 338, 
    336, 335, 344, 351, 352, 346, 332, 337, 332, 330, 336, 339, 336, _, 345, 
    345, 347, 2, 1, 348, 352, 353, 5, 7, 20, 12, 21, 20, 28, 22, 4, 2, 14, 
    13, 4, 1, 349, 343, 352, 348, 351, 348, 349, 346, 356, 346, 335, 337, 
    348, 334, 334, 339, 337, 330, 329, 346, 342, 342, 343, 353, 4, 359, 29, 
    22, 26, 33, 24, 354, 355, 17, 37, 30, 339, 344, 346, 347, 335, 336, 322, 
    15, 357, 319, 351, 350, _, 358, 330, 340, 326, 325, 323, 293, 305, 320, 
    311, 329, 289, 315, 311, 319, 320, 321, 321, 321, 318, 315, 311, _, 321, 
    319, 321, 329, 329, 327, 322, 323, 325, 325, 330, 334, 331, 333, 330, 
    323, 325, 330, 330, 324, 329, 330, 330, 334, 337, 332, 336, 348, 347, 15, 
    25, 29, 328, 307, 4, 338, 344, 326, 344, 336, 327, 324, 329, 356, 33, 
    352, 324, 332, 28, 323, 51, 19, 9, 2, 346, 359, 1, 340, 351, 6, 4, 320, 
    337, 338, 321, 323, 331, 332, 328, 338, 348, 355, 343, 313, 320, 325, 
    329, 321, 315, 327, 313, 321, 321, 326, 309, 329, 333, 318, 323, 338, 
    336, 339, 342, 342, 323, 305, 303, 318, 317, 316, 320, 317, 320, 333, 
    328, 320, 331, 332, 329, 331, 323, 305, 311, 314, 329, 335, 337, 335, 
    327, 321, 322, 316, 323, 357, 357, 349, 346, 348, 339, 352, 244, 271, 32, 
    22, 195, 167, 153, 137, 124, 116, 111, 114, 110, 112, 120, _, _, 105, 
    105, 107, 107, 113, 117, 115, 109, 100, 94, 90, 95, 96, 103, 111, 95, 91, 
    95, 87, 73, 61, 63, 67, 133, 66, 84, 105, 103, 105, 59, 53, _, _, _, 55, 
    55, _, 67, 64, 69, 85, 89, 102, 105, 105, 92, 106, 103, 88, 76, 91, 99, 
    76, 68, 81, 89, 85, 65, 62, 61, 63, 73, 85, 74, 78, 78, 82, 78, 81, 68, 
    71, 73, 70, 63, 58, 59, 73, 58, 56, 48, 46, 6, 90, 118, 44, 115, 50, 53, 
    50, 49, 31, 329, 36, 28, 21, 5, 354, 352, 334, 349, 342, 349, 347, 273, 
    336, 314, 332, 344, 351, 346, 345, 325, 341, 329, 316, 345, 282, 317, 
    130, 325, 349, 21, 329, 52, 71, 350, 328, 359, 357, 97, 324, 324, 161, 
    73, 140, 71, 102, 102, 59, 92, 54, 4, 0, 0, 0, 0, 0, 0, 0, 0, 316, 318, 
    321, 317, 310, 330, 325, 340, 327, 309, 323, 319, 327, 326, 322, 328, 
    325, 314, 308, 318, 316, 302, 304, 298, 298, 296, 300, 301, 304, 316, 
    322, 321, 318, 301, 314, 319, 321, 320, 323, 318, 317, 318, 316, 333, 
    323, 321, 325, 330, 320, 334, 332, 328, 330, 330, 327, 320, 313, 305, 
    301, 303, 301, 317, 328, 337, _, 315, 323, 331, 325, 328, 323, 338, 317, 
    5, 23, 348, 326, 9, 25, 26, 318, 315, 330, 319, 326, 326, 325, 320, 26, 
    325, 317, 326, 311, 328, 296, 302, 351, 350, 304, _, 338, 334, 38, 42, 
    45, 43, 39, 40, 25, 30, 301, 303, 277, 43, 28, 360, 56, 58, _, _, _, 55, 
    52, 52, 50, 55, 65, 43, 52, 54, 58, 59, 72, 74, 88, 88, 90, 88, 92, 85, 
    92, 73, 82, 82, 86, 85, 82, 83, 85, 79, 77, 71, 66, 67, 69, 69, 75, 78, 
    79, 77, 73, 70, 74, 72, 82, 71, 66, 67, 73, 74, 66, 64, 64, 63, 58, 58, 
    58, 55, 52, 54, 53, 51, 49, 49, 46, 47, 52, 43, 54, 48, 52, 47, 48, 51, 
    58, 87, 53, 28, 24, 20, 30, 35, 41, 42, 47, 47, 48, 50, 47, 48, 48, 46, 
    44, 43, 40, 39, 38, 33, 36, 34, 9, 336, 1, 358, 22, 24, 31, 34, 42, 39, 
    323, 289, 359, 3, 359, 319, 38, 102, 344, 36, 38, 45, 49, 48, 51, 58, 53, 
    54, 60, 66, 71, 77, 83, 78, 77, 76, 71, 60, 56, 54, 50, 50, 47, 57, 62, 
    62, 70, 64, 54, 64, 69, 68, 65, 61, 59, 65, 122, _, 93, 99, 97, _, 104, 
    118, 127, 136, 75, 65, 53, 58, 82, 90, 82, 83, 82, 73, 61, 59, 320, 192, 
    11, 65, 77, 57, 350, 27, 73, 325, 20, 299, 323, 284, 295, 344, 313, 47, 
    48, 46, 51, 50, 21, 6, 48, 46, 50, 50, 50, 48, 43, 20, 2, 349, 342, 354, 
    350, 342, 340, 345, 358, 339, 343, 347, 327, 338, 337, 327, 326, 341, 
    332, 328, 4, 340, 322, 332, 333, 330, 325, 325, 326, 322, 322, 329, _, 
    335, 331, 337, 331, 337, _, 337, 337, _, 332, 333, 331, 332, 325, 329, 
    333, 332, 329, 336, 333, 326, 323, 326, 324, 325, 329, 327, 330, 338, 
    339, 330, 333, 337, 350, 342, 330, 328, 336, 336, 333, 331, 333, 322, 
    321, 321, 321, 324, 327, 323, 324, 316, 321, 321, 322, 321, 323, 319, 
    313, 315, 307, 302, 310, 311, 306, 313, 315, 316, 326, 319, 328, 329, 
    327, 326, 321, 321, 321, 320, 319, 318, 311, 310, 312, 317, 316, 315, 
    317, 318, 322, 326, 319, 322, 315, 317, 318, 321, 321, 323, 326, 322, 
    309, 307, 305, 311, 308, 314, 310, _, 307, 305, 311, 302, 306, 309, 308, 
    305, 310, 311, 307, 304, 306, 306, 303, 303, 302, 297, 304, 300, 313, 
    317, 321, 317, 312, 312, 313, 311, 314, 313, 317, 321, 317, 313, 322, 
    323, 332, 330, 313, 320, 315, 322, _, 314, 318, 319, 341, 342, 345, 351, 
    345, 329, 330, 336, 338, 319, 317, 325, 16, 105, 111, 131, 152, 139, 142, 
    141, 139, 120, 115, 113, 114, 115, 113, 115, 110, 109, 112, 108, 113, 
    114, 115, 92, 37, 331, 320, 331, 2, 332, 352, 326, 334, 340, 27, 45, 47, 
    87, 91, 86, 92, 98, 96, 99, 116, 61, 99, 2, 348, 59, 327, 330, 323, 319, 
    328, 330, 325, 320, 312, 312, 314, 307, 295, 314, 345, 318, 325, 303, 
    310, 306, 309, 324, 334, 326, 250, 260, 205, 208, 200, 205, 210, 252, 
    286, 297, 294, 291, 298, 299, 316, 321, 327, 328, 324, 326, 326, 320, 
    326, 311, 294, 304, 306, 312, 313, 321, 312, 320, 321, 322, 338, 348, 1, 
    327, 316, 317, 317, 317, 318, 309, 316, 306, 312, 313, 314, 311, 318, 
    324, 334, 339, 326, 323, 329, 330, 319, 320, 322, 335, 331, 332, 325, 
    321, 334, 331, 311, _, 318, 319, 317, 311, 312, 321, 304, 303, 298, 299, 
    303, 294, 312, 294, 307, 309, _, 312, _, 334, 333, 341, 342, 346, 340, 
    343, 329, 311, 311, 313, 320, 314, 319, 315, 317, _, _, _, _, 319, 325, 
    28, 5, 113, 104, 117, 117, 112, 113, 117, 109, 101, 97, 158, 0, 0, 103, 
    112, 115, 115, 109, 116, 116, 127, 133, 123, 115, 122, 121, 128, 123, 
    123, 119, 118, 133, 129, 104, 100, 85, 92, 104, _, 103, 106, 99, 104, 
    104, 109, 112, 110, 104, 100, 94, 96, 92, 98, 93, 93, 98, 104, 107, 111, 
    111, 112, 110, 107, 107, 102, 100, 99, 97, 90, 89, 92, 94, 101, 105, 105, 
    105, _, _, _, _, 103, 104, _, _, 108, 117, 120, 118, 123, 128, 126, 114, 
    112, 111, 114, 105, 103, 103, 98, _, 93, 99, 101, 91, 95, 98, 101, 100, 
    103, 107, _, 110, 110, 109, 107, 107, 109, 110, 107, 103, 102, 97, 96, 
    99, 98, 96, 96, 100, 100, 101, 102, 101, 101, 100, 99, 94, 104, 104, 110, 
    109, 103, 106, 105, 111, 100, 104, 105, 103, 106, 106, 112, 109, 107, 
    107, 109, 106, 103, 109, 106, 101, 95, 102, 104, 106, 108, 103, 109, 119, 
    125, 127, 130, 123, 127, 126, 116, 128, 115, 128, 136, 131, 142, 136, 
    112, 108, 106, 104, 108, 94, 97, 96, 108, 109, 101, 103, 105, 82, 82, 60, 
    54, 49, 332, 358, 51, 52, 338, 310, 46, 55, 54, 61, 64, 58, 50, 55, 59, 
    72, 74, 82, 79, 79, 78, 86, 95, 100, 101, 104, 103, 121, 112, 96, 108, 
    116, 110, 109, 107, 103, 110, 141, 125, 128, 119, 116, 117, 106, 98, 132, 
    129, 127, 157, 126, 107, 94, 87, 76, 56, 58, 52, 49, 66, 49, 52, 48, 45, 
    48, 306, 46, 333, 359, 11, 347, 355, 336, 341, 305, 296, 310, 302, 294, 
    297, 302, 309, 313, 314, 314, 318, 329, 320, 326, 321, 323, 312, 313, 
    318, 313, 317, 315, 318, 313, 300, 305, 315, 312, 304, 305, 311, 311, 
    292, 306, 303, 294, 308, 296, 299, 298, 295, 305, 295, 295, 296, 296, 
    294, 292, 294, 290, 293, 290, 293, 289, _, 292, 292, 290, 290, 291, 295, 
    295, 301, 299, 295, 298, 294, 334, 334, 325, 336, 319, 319, 326, 322, 
    324, 328, 322, 327, 335, 335, 339, 332, 342, 335, 324, 324, 335, 333, 
    341, 335, 337, 336, 330, 328, 330, 315, 332, 324, 319, 322, _, 320, 325, 
    322, 338, 345, 346, 10, 17, 345, 349, 340, 339, 332, 321, 321, 320, 324, 
    326, 322, 327, 323, 328, 340, 339, 19, 335, 77, 66, 44, 17, 25, 45, 68, 
    70, 44, 58, 98, 334, 69, 67, 62, 83, 86, 87, 77, 76, 68, 65, 61, 60, 67, 
    74, 67, 73, 67, 81, 78, 84, 79, 69, 65, 67, 87, 90, 100, 116, 101, 113, 
    150, 112, 94, _, 74, 53, 56, 59, 60, 64, 70, 76, 62, 64, 69, 69, 66, 65, 
    65, 51, 59, 63, 61, 70, 71, 92, 81, 75, _, 67, 64, 69, 68, 78, 72, 70, 
    134, 117, 125, 114, 110, 120, 126, 100, 91, 91, 93, 79, 76, 73, 81, 95, 
    91, 90, 72, 74, 72, 50, 325, 327, 13, 5, 330, 320, 329, 311, 307, 312, 
    323, 319, 308, 311, 319, 328, 318, 321, 324, 302, 315, 331, 308, 309, 
    305, 312, 317, 314, 312, 321, 314, 315, 316, 309, 310, 307, 304, 304, 
    304, 309, 307, 307, 322, 306, 296, 306, 317, 330, 309, 323, 310, 303, 
    303, 308, 308, 316, 307, 321, 287, 309, 287, 305, 289, 313, 308, 330, 
    283, 325, 322, 349, 331, 333, 17, 15, 18, 26, _, 45, 22, 12, 324, 336, 
    356, 6, 354, 358, 354, 317, 325, 6, 30, 22, 10, _, 32, 29, 36, 35, 18, 
    33, 20, 51, 242, 117, 130, 109, 101, 115, 117, 93, _, 96, 87, 105, 84, 
    70, 127, 59, 149, 133, 131, 56, 105, 32, 16, 18, 310, 342, 131, 117, 118, 
    130, 128, 119, 141, 339, 68, 138, 157, 147, 121, 119, 140, 122, 132, 146, 
    169, 142, 150, 143, 121, 81, 88, 92, 113, 119, 119, 126, 118, 117, 119, 
    119, 112, 109, 113, 115, 111, 100, 105, 107, 103, 99, 97, 97, 94, 97, 90, 
    83, 82, 84, 81, 70, 61, 53, 180, 95, 344, 286, 294, 298, 310, 298, 306, 
    289, 296, 287, 288, 290, 290, 293, 300, 298, 292, 294, 302, 294, 287, 
    289, 289, 288, 288, 288, 289, 288, 288, 294, 292, 294, 287, 304, 349, 
    323, 18, 137, 119, 124, 132, 110, 108, 119, 117, 120, 123, 120, 121, 126, 
    123, 125, 114, 115, 125, 126, 127, 111, 5, 325, 325, 351, 330, 337, 337, 
    345, 337, 331, 332, 325, 327, 326, 328, 331, 4, 353, 301, 297, 309, 309, 
    313, 302, 310, 297, 296, 301, 300, 309, 311, 302, 303, 324, 324, 329, 
    328, 309, 325, 316, 306, 304, 343, 343, 355, 26, 18, 71, 81, 67, 67, 68, 
    67, 103, _, 129, 146, 137, 128, 127, 127, 125, 127, 127, 126, 131, 135, 
    140, 144, 144, 138, 132, 123, 119, 118, 69, 66, 57, 62, 64, 70, 60, 61, 
    58, 42, 47, 40, 33, 312, 336, 334, 329, 331, 333, 331, 328, 332, 335, 
    333, 330, 322, 327, 318, 318, 308, 305, 311, _, 295, 291, 300, 300, 296, 
    296, 288, 285, 287, 283, 287, 284, 287, 282, 286, 276, 286, 275, 278, 
    277, 272, _, 279, 273, 270, 276, 279, 275, 273, 298, 278, 272, 268, 259, 
    253, 249, 246, 247, 269, 257, 253, 256, 244, 252, 235, 229, 224, 205, 
    210, 218, 218, 204, 205, 214, 299, 316, 323, 308, 312, 295, 306, 285, 
    285, 290, 292, 283, 289, 280, 279, 277, 274, 260, 255, 255, 256, 254, 
    257, 249, 244, 184, 171, 157, 142, 111, 124, 129, 122, 138, 142, 193, _, 
    260, 266, 266, 281, 290, 308, 297, 292, 283, 282, 326, 351, 346, 121, 
    111, 117, 120, 115, 114, 121, 117, 122, 106, 101, _, 114, 117, 120, 121, 
    126, 122, 129, 173, 175, 222, 348, 299, 303, 305, 301, 307, 318, 325, 
    329, 330, 22, 106, 309, 125, 115, 129, 144, 130, 138, 139, 139, 139, 127, 
    121, 113, 117, 40, 2, 291, 309, 286, 276, 269, 295, 306, 339, _, 318, 
    326, 328, _, 337, 323, 310, 299, 65, 73, 81, 80, 89, 97, 115, 116, 101, 
    115, 116, 116, 112, 117, 111, 102, _, 99, 109, 116, 114, 113, 109, 115, 
    116, _, 118, 120, 117, 115, 110, 108, 114, 112, 114, 111, 92, 100, 106, 
    94, 99, 98, 103, 103, 106, 107, _, 111, 110, 107, 104, 104, 98, 97, 104, 
    108, 104, _, 112, 113, 122, 123, 139, _, _, 143, 129, _, 122, 116, 120, 
    118, _, _, _, 314, 120, 91, 123, 142, 131, 104, 108, 116, 121, 117, 117, 
    119, 123, 115, 123, 139, 114, _, _, 115, 100, 288, 339, 336, 332, 332, 
    324, 325, 322, 301, 282, 262, 271, 187, 182, 197, 257, 250, 241, 240, 
    219, 67, 138, 134, 132, 122, 119, 130, 127, 145, 128, 96, 78, 90, 98, 
    117, 122, 258, 320, _, 290, 289, 284, 294, 294, 291, 291, 290, 285, 279, 
    281, 273, 267, 259, 254, 252, 255, 273, 268, 260, 271, 273, 276, 273, 
    286, 305, 297, 270, 240, 263, 131, _, 189, 168, 162, 120, 116, 117, 126, 
    125, 116, 113, 106, 154, 132, 115, 123, 129, 165, 277, 258, 295, 287, 
    310, 315, 319, 310, 320, 304, 301, 307, 308, 297, 302, 303, 287, 283, 
    288, 289, 288, 284, 274, 281, 285, 284, 281, 286, 298, 305, 300, 298, 
    304, 299, 301, 302, 303, 302, 300, 303, 298, 301, 303, 310, 307, 297, 
    301, 303, 299, 278, 279, 300, 306, 304, 288, 284, _, 291, 297, 283, 300, 
    290, 290, 278, 280, 277, 286, 286, 276, 281, 277, 282, 283, 286, 287, 
    283, 283, 281, 282, 293, 289, 279, 275, 266, 281, 290, 288, 275, 280, 
    284, 286, _, 246, 271, 258, 246, 246, 248, 291, 274, 266, 236, 244, 227, 
    279, 270, 269, 269, 263, 208, 239, 263, 278, 270, 262, 257, 260, 266, 
    259, 260, 272, 268, 257, 263, 262, 265, 271, 277, 264, 283, 279, 275, 
    286, 282, 282, 284, 296, 291, 271, 280, 289, 286, 277, 305, 288, 293, 
    278, 273, 280, 275, 282, 293, 275, 278, 277, 264, 264, 268, 266, 267, 
    285, 285, 290, 286, 256, 265, 258, _, _, 268, 271, 265, 249, 255, 234, 
    208, 199, 179, 180, 154, 146, 126, 130, 121, 123, 118, 175, 197, 153, 
    143, 133, 135, 106, 124, 129, 118, 133, 136, 137, 126, 132, 134, 165, 
    135, 148, 123, 221, 284, 313, 295, 287, 320, 312, 315, 295, 241, 250, 
    338, 157, 157, 144, 133, 312, 169, 61, 67, 62, 72, 77, 69, 58, 305, 9, 
    308, 204, 0, 328, 319, 328, _, 97, 181, 287, 303, 326, 266, 211, 127, 
    109, 132, 114, 115, 104, 118, 122, 120, 136, 117, 115, 108, 117, 128, 
    125, 125, 125, 125, 114, 111, 110, 122, 115, 115, 124, 118, 111, 114, 
    122, 118, 126, 125, 127, 124, _, 126, 132, 76, 77, 64, 68, 71, 67, 69, 
    65, 55, 11, 1, 57, 306, _, 272, 329, 309, 341, 302, 269, 274, 328, 309, 
    78, 94, 109, 135, _, 125, 115, 108, 82, 96, 77, 68, 74, 68, 70, 71, 70, 
    66, 65, 64, 67, 60, 62, 63, 57, 68, 82, 119, 97, 142, 137, 136, 180, 153, 
    302, 309, 320, 310, 352, 121, 214, 230, 227, 225, 221, 216, 220, 240, 
    257, 267, 267, 264, 271, 279, 282, 282, 273, 279, _, _, _, _, _, 302, 
    302, 309, 303, 311, 317, 321, 325, 170, 112, 101, 127, 135, 142, 136, 
    130, 91, 95, 82, 94, 95, 92, 97, 108, 123, 118, 130, 108, 118, 127, 118, 
    132, 136, 136, 134, 139, 139, 141, _, 118, 125, 135, 132, 155, 145, 162, 
    152, 146, 138, 127, 134, 133, 131, 123, 136, 126, 121, 122, 117, 122, 
    107, 124, 116, 113, 111, 111, 113, 115, 133, 141, 345, 126, 105, 69, 102, 
    132, 119, 124, 123, 117, 143, 168, 135, 117, 129, _, 143, 134, 343, 271, 
    240, 133, 144, 132, 143, 133, 86, 76, 77, 84, 131, 98, 113, 104, 100, 
    106, 72, 65, 339, 68, 54, 323, 256, 334, 309, 39, 210, 232, 321, 170, 
    135, 144, 134, 123, 116, 111, 136, 107, 111, 101, 94, 109, 94, 100, 93, 
    _, 90, 87, 92, 107, 107, 113, 114, _, 125, _, 103, 142, 114, 127, 135, 
    116, 103, 299, 300, 217, 91, _, 121, 115, 124, 127, 124, 120, 119, 119, 
    113, 126, 112, 109, 111, 123, 127, 122, 182, 273, 304, 307, 307, 313, 
    288, 342, 334, 323, 305, 310, 323, 304, 315, 339, 155, 320, 359, 346, 
    262, 293, 328, 197, 52, 64, 60, 65, 53, 57, 53, 55, 331, 48, 48, 47, 44, 
    41, 333, 334, 351, 12, 348, 346, 20, 53, 55, 58, 258, 28, 37, 344, 360, 
    57, 57, 51, 60, 52, 48, 49, 56, 51, 52, 55, 61, 58, 59, 67, 71, 68, 81, 
    75, 86, 91, 89, 98, 91, 92, 80, 86, 98, 99, 85, 88, 84, _, 85, 76, 81, 
    78, 88, 98, 92, 91, 89, 100, 98, 95, 73, 74, 72, 79, 80, 85, 89, 102, 91, 
    75, 89, 106, 92, 88, 93, 73, _, 92, 109, 109, 113, 116, 113, 115, 115, 
    114, 117, 112, 115, 114, 104, 100, 99, 111, 111, 98, 106, 101, 106, 103, 
    112, 111, 117, 112, 105, 107, 102, 116, 102, 111, 113, 113, 114, 68, 83, 
    63, 47, 304, 289, 318, 340, 60, 205, 315, 328, 312, 296, 301, 322, 317, 
    312, 304, 287, 280, 304, 304, 297, 313, 287, 275, 148, 223, 201, 181, 
    198, 0, 114, 108, 94, 76, 67, 93, 109, 120, 109, 107, 97, 90, 79, 70, 68, 
    _, 57, 45, 45, 48, 50, 54, 51, 59, 322, 38, 343, 346, 323, 300, 309, 316, 
    23, 312, 358, 318, 301, 305, 10, 314, 325, 328, 317, 312, 318, 320, 327, 
    323, 324, 330, 310, 311, 313, 334, 323, 334, 323, 318, 323, 321, 317, 
    321, 327, 318, 320, 324, 321, 322, 318, 317, 320, 320, 322, 320, 328, 
    329, 327, 325, 325, 332, 326, 331, 329, 327, 327, 317, 325, 329, 324, 
    316, 321, 321, 329, 326, 322, 315, 324, 321, 319, 327, 327, 328, 324, 
    326, 339, 311, 319, 328, 326, 325, 328, 322, _, 326, 325, _, 323, 325, 
    327, 329, 332, 333, 333, 325, 325, 323, 329, 329, 321, 323, 316, 325, 
    329, 329, 323, 317, 320, 301, 298, 294, 286, 301, 311, 298, 300, 296, 
    310, 305, 311, 308, 304, 288, 287, 282, 283, 273, 284, 288, 279, 284, 
    285, 281, 271, 268, 279, 284, 291, 292, 292, 301, 296, 286, 293, 274, 
    248, 221, 174, 175, 174, 159, 171, 148, 165, 215, 219, 315, 280, 310, 
    295, 318, 314, 306, 308, 316, 27, 129, 115, 140, 273, 313, 287, 278, 322, 
    302, 270, _, 269, 178, 77, 289, 189, 94, 153, 152, 143, 155, 295, 144, 
    141, 140, 145, 146, 155, 279, 190, 150, _, _, 256, 273, 287, 248, 268, 
    289, 59, 60, 69, 57, 60, 59, 68, 70, 58, 37, 64, 59, 48, 38, 47, 58, 55, 
    56, 57, 60, 58, 60, 58, 54, 53, 57, 61, 59, 67, 73, 77, 84, 84, 82, 71, 
    62, 69, 72, 75, 79, 89, 100, 107, 109, 114, 116, 116, 115, 115, 115, 112, 
    113, 113, 119, 118, 113, _, 117, 117, 125, 119, 116, 114, 112, 116, _, 
    121, 127, 128, 127, 132, 128, 134, 130, 124, 127, 129, 127, 126, 110, 
    112, 118, 141, 109, 111, 119, 155, _, 296, 319, 304, 337, 358, 350, 1, 
    360, 360, 24, 313, 301, 318, _, 332, 0, 324, 141, 332, 321, 307, 332, 
    330, 329, 31, 171, 232, 358, 30, 172, 168, 137, 165, 165, 162, 80, 109, 
    121, 127, 107, 108, 108, 118, 104, 110, 113, 107, 112, 117, _, 134, 134, 
    129, 107, 125, _, 133, 132, 152, 226, 249, 259, 283, 242, 250, 263, 252, 
    254, 253, 259, 270, 263, 297, 305, 304, 304, 281, 232, 218, 182, 120, 91, 
    105, 95, 90, 85, 86, 79, 75, 88, 90, 88, 117, 97, 108, 103, 107, 105, 
    102, 103, 99, 105, 107, 132, 132, 133, 132, 135, 122, 131, 121, 118, 114, 
    126, 129, 126, 134, 114, _, 116, 144, 146, 121, 107, 116, 124, 116, 122, 
    125, 144, 119, 118, 113, 100, 96, 94, 103, 126, 114, 116, 111, 114, 112, 
    123, 94, 106, 94, 174, 196, 256, 315, 304, 310, 314, 306, 287, 159, 175, 
    84, 80, 78, 76, 76, 87, 88, 91, 80, 99, 112, 121, 106, 114, 105, 101, 
    117, 110, 135, 145, 141, 144, 117, 117, 116, 122, 119, 115, 112, 113, 
    121, 103, 97, 92, 80, 97, 80, 71, 81, 79, 73, 68, 66, 65, 8, 240, 104, 
    129, 97, 132, 118, 119, 94, 99, 87, 83, 69, 69, 90, 106, 102, 106, 100, 
    91, 98, 83, 63, 62, 98, 77, 84, 101, 96, 95, 111, 117, 113, 116, 114, 
    112, 110, 118, 119, 126, 121, 115, 125, 134, 138, 143, 220, 313, 315, 
    304, 308, 298, 310, 304, 307, 306, 307, 306, 300, 301, 300, _, 306, 297, 
    310, 309, 308, 310, 318, 307, 305, 327, 324, 310, 325, 324, 310, 323, 
    327, 309, 313, 312, 307, 329, _, _, _, 155, 172, 65, 256, 285, 149, 185, 
    193, 115, 149, 141, 150, 167, 154, _, _, _, _, 145, 151, 144, 214, 152, 
    215, _, 255, 169, 182, 237, 292, 312, 307, 319, 113, 133, 343, 322, 320, 
    327, 294, 307, 345, 273, 0, 256, 285, 129, 149, 106, 108, 112, 112, 98, 
    88, 97, 100, 106, 105, 109, 116, 118, 116, 129, 122, 117, 121, 121, 117, 
    114, 121, 111, 113, 115, 121, 119, 127, 120, 118, 110, 108, 102, 104, 99, 
    87, 106, 305, 327, 320, 4, 344, 343, 327, 328, 328, 331, 332, 343, 335, 
    342, 348, 342, 348, 343, 342, 343, 337, 341, 343, 345, 353, 352, 346, 
    343, 348, 331, 335, 331, 323, _, 328, 317, 298, 322, 327, 318, 304, 292, 
    298, 295, 287, 279, 276, 283, 290, 285, 293, 256, 150, 125, 155, 167, 
    212, 253, 211, 203, 198, 233, 266, 276, 283, 295, 298, 299, 297, 295, 
    293, 285, 280, 278, 279, 268, 271, 270, 252, 251, 256, 232, 219, 209, 
    214, 208, 205, 198, 192, 180, 178, 168, 175, 132, 130, 150, 119, 115, 
    127, 194, 192, 165, 192, 166, 118, 149, 208, 276, 300, 306, 323, 341, 
    341, 316, 320, 7, 61, 70, 66, 73, 80, 326, 329, 332, 327, 323, 322, 321, 
    313, 297, 279, 264, 248, 295, 171, 37, 43, 26, 7, 1, 347, 355, 339, 332, 
    330, 331, 334, 327, 321, 318, 306, 298, 297, 307, 300, 286, 280, 277, 
    283, 278, 306, 311, 331, 132, 95, 95, 114, 113, 111, 119, 126, 136, 128, 
    129, 125, 128, 161, 99, 92, 101, 110, 112, 117, 104, 115, 107, 105, 115, 
    113, 110, 121, 117, 125, 115, 112, 116, 125, 123, 119, 109, 111, 104, 
    118, 114, 118, 124, 133, 131, 122, 115, 115, 132, 134, 115, 109, 114, 
    112, 114, 112, 117, 117, 113, 111, 113, 112, 112, 114, 115, 111, 114, 
    112, 112, 122, 113, 114, 120, 109, 118, 115, 114, 118, 118, 113, 111, 
    118, 110, 107, 101, 116, 116, 120, 113, 103, 105, 96, 98, 101, 110, 106, 
    106, 105, 93, 93, 88, 84, 79, 80, 82, 88, 93, 93, 99, 104, 110, 112, 113, 
    97, 99, 98, 93, 94, 88, 84, 80, 83, 78, 83, 85, 92, 88, 78, 78, _, 78, 
    67, 77, 83, 86, 88, 85, 82, 86, 94, 90, 96, 91, 88, 89, 78, 76, 80, 88, 
    97, 116, 111, 112, 117, 114, 117, 115, 118, 120, 122, 115, 123, 116, 119, 
    113, 111, 108, 119, 114, 106, 81, 82, 75, 63, 75, 90, 100, 96, 93, 105, 
    94, 111, 118, 130, 119, 138, 114, 138, 113, 96, 123, 116, 120, 127, 124, 
    134, 122, 82, 71, 70, 65, 69, 67, 71, 250, 325, 69, 129, 94, 98, 125, 
    103, 127, 130, 110, 94, 83, _, 96, 90, 107, 109, 91, 96, 79, 82, 73, 64, 
    300, 335, 24, 131, 76, 308, 300, 313, 288, 296, 284, 205, 245, 292, 307, 
    294, 301, 314, 332, 318, 20, 0, 16, 142, 139, 89, 116, 117, 139, 134, 
    131, 137, 135, 104, 109, 112, 112, 113, 115, 121, 124, 119, 120, 118, 
    116, 113, 107, 109, 114, 114, 110, 109, 104, _, 95, 91, 89, 85, 76, 75, 
    66, 68, _, 74, 70, 79, 77, 82, 87, 80, 71, 77, 69, 63, 66, 63, 63, 64, 
    59, 68, 74, 68, 70, 62, 64, 67, 64, 60, 61, 60, 61, 67, 62, 63, 68, 69, 
    73, 74, 71, 71, 72, 76, 75, 78, 78, 74, 79, 70, 55, 54, 58, 55, 59, 59, 
    57, 60, 64, 59, 54, 57, 54, 48, 45, 47, 58, 61, 51, 44, 40, 40, 41, _, 
    40, 43, _, 42, 42, 42, 46, 42, 43, 40, 38, 35, 11, 11, 350, 347, 343, 
    341, 334, 337, 325, 319, 322, 325, 334, 318, 327, 325, 320, 333, 307, 
    311, 309, 308, 318, 313, 316, 311, 314, 320, 312, 304, 297, 304, 312, 
    317, 318, 312, 317, 319, 320, 312, 302, 298, 300, 303, 299, 298, 301, 
    301, 300, 300, 310, 308, 309, 309, 295, 307, 297, 290, 311, 305, 296, 
    294, 297, 298, 310, 309, 314, 310, 315, 324, 327, 328, 330, 325, 305, 
    311, 262, 257, 234, 256, 243, 237, 251, 231, 201, 204, 149, 352, 171, 
    161, 131, 118, 139, 144, 194, 169, 162, 147, 169, 174, 180, 162, 186, 
    176, 186, 186, 170, 129, 131, 181, 169, 155, 148, 123, 115, 115, 114, 
    116, 119, 122, 125, 124, 121, 114, 116, 114, 117, 114, 114, 117, 131, 
    124, 117, 114, 114, 119, 119, 112, 115, 113, 106, 115, 118, 116, 117, 
    129, 103, 134, 123, 107, 110, 123, 128, 128, 128, 124, 130, 119, 117, 
    115, 101, 146, 117, 120, 120, 113, 121, 119, 125, 132, 105, 107, 121, 
    135, 137, 106, 134, 110, 110, 118, 110, 129, 99, 129, 110, 102, 112, 121, 
    112, 117, 107, 115, 119, 121, 113, 104, 107, 126, 158, 311, 270, 277, 
    304, 298, 304, 307, 299, 280, 199, 118, 128, 176, 191, 157, 110, 113, 
    124, 115, 140, 113, _, 103, 27, 321, 328, 340, 321, 321, 322, 343, 325, 
    333, 328, 299, 315, 360, 124, 84, 31, 66, 70, 69, 69, 66, 59, 51, 21, 
    323, 3, 337, 331, 327, 315, 307, 312, _, 286, 286, 296, 292, 295, 307, 
    314, 311, 314, 309, 309, 319, 315, 318, 330, 331, 318, 324, 339, 335, 60, 
    66, 99, 106, 71, 82, 85, 79, 102, 84, 81, 80, 81, 79, 87, 74, 70, 65, 60, 
    60, 25, 60, 56, 56, 47, 39, 23, 15, 9, 28, 36, 36, 48, 45, 51, 51, 40, 
    49, 53, 51, 49, 52, 58, 38, 55, 65, 64, 66, 66, 66, 64, 70, 67, 63, 59, 
    63, 66, 76, 90, 87, 76, 70, 73, 75, 83, 92, 86, 94, 98, 96, 92, 82, 95, 
    98, 101, 90, 93, 92, 93, 91, 83, 73, 72, _, 90, 91, 94, 92, 89, 107, 113, 
    107, 108, 132, 124, 116, 114, 136, 137, 125, 114, 118, 115, 114, 99, 92, 
    107, 102, 103, 107, 106, 106, 116, 126, 123, 128, 133, 139, 129, 116, 
    110, 161, 19, 12, 326, 315, 318, 336, 316, 330, 305, 328, 333, 335, 302, 
    315, 319, 332, 312, 298, 286, 282, 306, 310, 306, 303, 171, 120, 123, 
    119, 113, 108, 107, 127, 102, 98, 86, 80, 87, 76, 84, 91, 88, 81, 85, 88, 
    89, 84, 86, 83, 90, 90, 104, 98, 105, 113, 121, 116, 111, 110, 114, 102, 
    116, 121, 126, 128, 123, 140, 135, 124, 120, 128, 130, 130, 118, 125, 
    118, 125, _, 10, 0, 141, 34, 0, 132, 318, 345, 359, 151, 306, 110, 153, 
    99, 136, 105, 343, 310, 133, _, 132, 114, 102, 122, 117, _, 304, 92, 111, 
    97, 101, 88, 85, 81, 76, 69, 65, 70, 77, 88, 81, 84, 98, 102, 88, 85, 84, 
    79, 90, 85, 83, 84, 88, 90, 95, 99, 96, 103, 106, 117, _, 114, 113, 110, 
    113, 112, 107, 108, 108, 116, 106, 104, 112, 112, 104, 110, 95, 91, 98, 
    101, 94, 93, 103, 102, 101, 101, 104, 105, 108, 110, 117, 101, 102, 97, 
    99, 97, 97, _, 94, 105, 107, 105, 112, 116, 108, 111, 115, 122, 118, 121, 
    125, 140, 122, _, 325, 307, 15, 0, 356, 333, 322, 325, 298, 316, 0, 322, 
    316, 321, 317, _, _, _, 312, 309, 318, 325, 1, 352, 305, 326, 116, 125, 
    98, _, 125, 122, 115, 72, 72, 103, 68, 72, 75, 88, 100, 147, 131, 125, 
    116, 97, 93, 99, 113, 126, 123, 114, 119, 112, 113, 115, 108, 120, 135, 
    144, 126, 123, 125, 126, 118, 125, 137, 126, 130, 157, 138, 148, 118, 
    138, 146, 136, 147, 135, 143, 137, _, 136, 140, 133, 126, 146, 157, 157, 
    153, 154, 160, 157, 154, 168, 134, 151, 133, 121, 144, 128, 133, 151, 
    172, 140, 141, 128, 122, 123, 120, 118, 119, 132, 130, 114, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 123, 
    124, 116, 113, 128, 121, 122, 116, 116, 113, 131, 110, 115, 105, 106, 
    132, 110, 123, 100, 99, 103, 132, 126, 131, 140, 140, 145, 154, 145, 135, 
    125, 132, 127, 131, 114, 118, 120, 130, 129, 126, 121, 121, 122, 119, 
    118, 127, 133, 131, 130, 126, 134, 129, 139, 140, 134, 128, 121, 109, 
    117, 0, _, 295, 285, 285, 292, 284, 244, 224, 354, 193, 153, 114, 140, 
    134, 129, 144, 127, 115, 112, 111, 80, 65, 63, 130, 103, 309, 302, 299, 
    306, 306, 299, 292, 284, 281, 270, 270, 273, 285, 282, 280, 283, 286, 
    282, 282, 279, 279, 281, 280, 308, 307, 303, 306, 301, 303, 300, 305, 
    299, 308, 303, 304, 310, 305, 310, 307, 304, 303, 304, 308, 302, 308, 
    312, 308, _, 315, 318, 320, 317, 329, 332, 334, 331, 333, 333, 338, 332, 
    334, 331, 338, 335, 348, 358, 358, 341, 6, 9, 1, 3, 4, _, 2, 6, 16, 3, 
    14, 27, 9, 9, 23, 30, 17, 32, 17, 43, 16, 44, 27, 20, 15, 27, 46, 29, 20, 
    27, 14, 32, 36, 41, 35, 56, 47, 48, 43, 28, 46, 67, 48, 35, 49, 92, 117, 
    97, 85, 106, 292, 84, 93, 71, 112, 99, 86, 84, 84, 81, 95, 97, 131, 188, 
    153, 133, 122, 105, 178, 154, 181, 172, 177, 172, 170, 172, 170, 169, 
    188, 168, 178, 149, 142, 153, 141, 100, 106, 145, 131, 113, 110, 101, 
    115, 106, 96, 94, 89, 79, 77, _, 67, 76, 66, 69, 71, 70, 81, 93, 108, 
    115, 123, 114, 116, 113, 109, 102, 102, 96, 97, 90, 92, 86, 77, 79, 78, 
    80, 80, 77, 75, 72, 74, 69, 65, 59, 279, 337, 39, 8, 337, 332, 330, 301, 
    317, 327, 288, 285, 284, 285, 282, 278, 344, 359, 1, 31, 29, 36, 47, 41, 
    38, 38, 30, 27, 22, 7, 9, 2, 6, 9, 11, 14, 11, 1, 0, 8, 23, 9, 23, 20, 
    25, 27, 29, 28, 15, 26, 28, 25, 47, 53, 58, 49, 55, 53, 59, _, 60, 65, _, 
    45, 48, 50, 51, 48, 43, 21, 28, 24, 46, 38, 24, 24, 17, 25, 28, 38, 21, 
    32, 43, 47, 33, 28, 38, 19, 18, 15, 328, 9, 9, 20, 19, 10, 40, 28, 33, 7, 
    30, 56, 54, 47, 45, 52, 45, 35, 15, 19, 28, 36, 39, 56, 60, 90, 81, 86, 
    99, 143, 194, 229, 211, 224, 233, 338, 322, 322, 7, 51, 251, 276, 302, 
    297, _, 300, 317, 309, 325, 316, 325, 356, 352, 4, 10, 5, 4, 3, 360, 1, 
    1, 8, 21, 10, 2, 346, 337, 331, 330, 351, 5, 3, 8, 12, 38, 35, 31, 26, 
    17, 13, 15, 14, 42, 10, 10, 345, 320, 326, 305, 312, 332, 320, 330, 351, 
    11, 14, 342, 334, 324, 328, 13, 335, _, 298, 344, 307, 11, 307, 8, 2, 9, 
    329, 335, 315, 330, 327, _, 359, 12, 293, 327, 314, 318, 5, 316, 347, 9, 
    27, 31, 24, 31, 10, 37, 31, 35, 34, 36, 32, 18, 21, 10, 357, 350, 285, 
    93, 117, 188, 189, 202, 237, 262, 265, 284, 330, 342, 360, 25, 21, 14, 
    296, 288, 284, 291, 297, 295, 301, _, 296, 310, 302, 313, 259, 239, 257, 
    _, 306, 310, 303, 318, 320, 344, 348, 348, 14, 25, 23, 357, 329, 316, 
    324, 308, 311, 319, 303, 309, 311, 304, 308, 308, 298, 304, 321, 302, _, 
    304, 316, 306, 306, 299, 303, 282, 285, 303, 296, 302, 307, 317, 301, 
    304, 312, 297, 301, 301, 306, 306, 305, 305, 311, 302, 307, 307, 303, 
    314, 308, 307, 306, 304, 315, 301, 297, 298, 301, 307, 309, 304, 299, 
    304, 305, 309, _, _, _, 301, 305, 310, 296, 306, 306, 308, 304, 300, 300, 
    294, 300, 301, 308, 305, 298, 301, 301, 303, 304, 303, 301, 309, 302, 
    306, 303, 316, 316, 310, 308, 310, 311, 311, 307, 305, 313, 314, 317, 
    315, 310, 320, 320, 306, 317, 313, 315, 316, 326, 336, 357, 4, 11, 10, 
    17, 18, 20, 23, 25, 42, 49, 51, 52, 53, 58, 45, 54, 43, 51, 44, 51, 49, 
    37, 43, 42, 38, 34, 39, 36, 35, 35, 35, 29, 29, 29, 38, 14, 30, 32, 35, 
    27, 20, 360, 14, 20, 349, 4, 11, 359, 21, 21, 35, 17, 34, 51, 17, 63, 57, 
    61, 57, 56, 55, 55, 69, 105, 83, 90, 80, 19, 11, 26, 30, 35, 22, 28, 21, 
    8, 3, 332, 332, 317, 315, 320, 308, 314, 307, 311, 311, 308, 311, 301, 
    303, 305, 320, 312, 309, 326, 333, 309, 360, 32, 29, 19, 38, 10, 47, 57, 
    69, 22, 27, 21, 44, 42, 45, 55, 50, 60, 51, 49, 57, 51, 46, 48, 55, 50, 
    58, 58, 69, 76, 86, 71, 78, 83, 76, 74, 77, 69, 76, 73, 65, 62, 64, 75, 
    67, 67, 71, 63, 63, 66, 64, 64, 66, 65, 64, 64, 60, 55, 52, 52, 68, 110, 
    103, 94, 69, 75, 72, 73, 74, 97, 31, 18, 360, 319, 311, 316, 323, 316, 
    319, 324, 327, 330, 321, 341, 331, 332, 325, 343, 348, 349, 9, 283, 237, 
    122, 327, 55, 63, 65, 67, 70, 66, 71, 72, 71, 70, 74, 73, 70, 67, 72, 74, 
    71, 72, 77, 77, 75, 78, 76, 72, 88, 101, 103, 130, 166, 171, 0, 209, 237, 
    277, 237, 216, 190, 210, 185, 169, 175, 171, 170, 187, 186, 176, 177, 
    174, 176, 176, 176, 173, 182, 199, 202, 233, 237, 209, 209, 199, 185, 
    184, 197, 206, 192, 217, 212, 223, 173, 168, 181, 199, 257, 291, 354, 31, 
    116, 271, 263, 266, 277, 264, 277, 270, 286, 278, 285, 293, 291, 292, 
    287, 284, 300, 303, 306, 295, 309, 315, 311, _, _, _, _, _, 308, 306, 37, 
    54, 55, 68, 110, 207, 185, 188, 138, 138, 122, 140, 203, 161, 157, 162, 
    152, 169, 176, 164, 159, 159, 160, 156, 164, 167, 161, 156, 156, 149, 
    144, 140, 137, 156, 138, 135, 135, 136, 121, 116, 117, 114, 110, 109, 94, 
    95, 97, 99, 101, 102, 106, 126, 260, 271, 281, 285, 291, 298, 303, 300, 
    300, 286, 288, 280, 293, 293, 273, 271, 255, 262, 250, 242, 236, 236, 
    229, 232, 229, 230, 217, 211, 207, 202, 182, 200, 207, 217, 216, 217, 
    242, 238, 246, 258, 283, 291, 288, 292, 297, 296, 293, 308, 306, 317, 
    309, 315, 318, 314, 317, 317, 320, 307, 305, 298, 316, 309, 301, 303, 
    301, 311, 296, 291, 302, 300, 300, 305, 306, 297, 322, 305, 286, 281, 
    292, 266, 239, 107, 170, 179, 153, 144, 153, 148, 163, 148, 145, 131, 
    125, 119, 121, 115, 111, 109, 110, 100, 103, 111, 116, 119, 121, 123, 
    125, 130, 129, 124, 121, 120, 123, 122, 114, 113, 113, 111, 126, 304, 
    315, 311, 318, 315, 319, 325, 325, 324, 326, 325, 323, 314, 315, 314, 
    223, 117, 87, 88, 84, 87, 71, 79, 79, 80, 294, 288, 294, 309, 311, 309, 
    310, 312, 313, 318, 314, 319, 316, 314, 316, 307, 309, 290, 273, 278, 
    269, 276, 284, 301, 310, 358, 3, 14, 33, 42, 42, 48, 80, 103, 168, 172, 
    117, 209, 268, 8, 7, 325, 13, 15, 22, 24, 18, 15, 25, 13, 16, 17, 18, 46, 
    47, 35, 27, 22, 19, 11, 12, 14, 15, 349, 5, 353, 348, 345, 343, 353, 357, 
    358, 30, 33, 20, 25, 21, 17, 30, 9, 343, 326, 343, 338, 333, 358, 337, 
    13, 33, 34, 43, 28, 35, 31, 43, 49, 64, 75, 75, 81, 78, 83, 82, 87, 82, 
    118, 110, 115, 123, 117, 140, 133, 140, 133, 127, 134, 142, 143, 142, 
    146, 141, 134, 125, 117, 105, 101, 101, 100, 99, 103, 98, 99, 98, 92, 83, 
    87, 95, 87, 74, 74, 66, 74, 73, 74, 75, 74, 76, 79, 78, 72, 67, 74, 75, 
    76, 69, 69, 68, 60, 50, 44, 39, 41, 37, 34, 25, 15, 11, 13, 6, 6, 1, 1, 
    2, 360, 360, 354, 352, 355, 353, 338, 334, 326, 322, 322, 320, 333, 320, 
    332, 324, 322, 324, 320, 314, 322, 316, 317, 327, 318, 310, 308, 322, 
    312, 309, 301, 309, 296, 308, 301, 299, 303, 301, 299, 300, 291, 302, 
    303, 304, 308, 314, 315, 315, 313, 300, 304, 303, 303, 297, 293, 306, 
    312, 308, 308, 335, 314, 322, 317, 4, 346, 51, 48, 49, 48, 49, 51, 49, 
    50, 55, 51, 356, 2, 1, 2, 334, 320, 329, 314, 331, 345, 343, 335, 330, 
    330, 327, 295, 301, 325, 310, 314, 303, 317, 304, 301, 315, 294, 288, 
    307, 314, 311, 300, 301, 293, 296, 289, 279, 267, 277, 277, 286, 276, 
    276, 266, 277, 267, 273, 270, 275, 277, 284, 273, 272, 307, 319, 300, 
    297, 9, 19, 21, 12, 20, 16, 18, 10, 17, 33, 35, 39, 45, 40, 30, 26, 28, 
    14, 5, 3, 2, 2, 2, 360, 330, 351, 3, 1, 360, 335, 345, 334, 348, 317, 
    313, 319, 292, 303, 306, 297, 292, 299, 308, 318, 321, 317, 335, 319, 
    319, 315, 322, 315, 309, 295, 290, 306, 310, 308, 305, 317, 324, 336, 1, 
    19, 288, 304, 311, 304, 315, 297, 294, 297, 298, 309, 311, 309, 309, 309, 
    309, 307, 310, 304, 309, 307, 306, 299, 309, 290, 301, 305, 302, 309, 
    303, 303, 304, 330, 353, 330, 326, 325, 7, 6, 5, 2, 359, 3, 14, 10, 7, 6, 
    9, 355, 2, 4, 356, 360, 2, 360, 354, 353, 352, 360, 359, 348, 351, 3, 
    351, 355, 342, 335, 348, 347, 1, 2, 2, 354, 327, 334, 331, 333, 330, 336, 
    329, 340, 335, 335, 330, 320, 316, 320, 324, 323, 330, 326, 321, 315, 
    317, 332, 321, 317, 319, 320, 322, 325, 322, 317, 331, 337, 320, 322, 
    325, 333, 349, 341, 335, 336, 336, 343, 345, 337, 336, 334, 334, 333, 
    330, 333, 334, 337, 331, 327, 332, 323, 320, 322, 310, 335, 327, 324, 
    318, 317, 308, 308, 308, 290, 294, 290, 294, 297, 299, 309, 303, 297, 
    296, 297, 292, 289, 292, 298, 302, 307, 299, 304, 315, 341, 340, 341, 
    354, 352, 6, 6, 1, 84, 97, 99, 100, 106, 113, 230, 224, 328, 2, 353, 332, 
    358, 81, 338, 358, 352, 356, 15, 26, 30, 36, 7, 323, 71, 347, 33, 40, 
    321, 47, 38, 3, 59, 20, 5, 356, 57, 39, 48, 28, 322, 62, 56, 58, 54, 52, 
    44, 44, 45, 46, 44, 41, 45, 48, 48, 50, 53, 62, 64, 62, 73, 53, 57, 50, 
    51, 59, 55, 55, 54, 54, 53, 51, 51, 51, 47, 40, 32, 30, 26, 24, 20, 360, 
    360, 358, 324, 311, 312, 308, 297, 283, 295, 287, 307, 293, 307, 300, 
    305, 305, 295, 239, 248, 229, 199, 162, 158, 148, 158, 133, 138, 117, 
    115, 107, 100, 109, 115, 135, 113, 111, 173, 203, 210, 161, 207, 236, 
    260, 251, 239, 209, 206, 126, 219, 137, 111, 105, 101, 110, 104, 113, 
    123, 118, 127, 149, 134, 129, 111, 118, 116, 117, 114, 116, 113, 116, 
    119, 120, 124, 125, 116, 110, 113, 115, 122, 121, 121, 114, 101, 100, 
    100, 105, 101, 107, 106, 104, 106, 104, 101, 103, 105, 108, 115, 115, 
    115, 103, 109, 104, 97, 93, 94, 94, 98, 100, 106, 108, 108, 107, 107, 
    108, 107, 105, 110, 120, 115, 114, 125, 128, 116, 119, 115, 119, 115, 
    109, 70, 66, 10, 3, 1, 3, 13, 31, 38, 36, 44, 51, 55, 54, 60, 57, 63, 72, 
    75, 82, 75, 86, 94, 84, 82, 87, 84, 101, 108, 104, 106, 111, 95, 105, 
    102, 99, 99, 99, 102, 92, 96, 98, 94, 77, 80, 88, 107, 93, 85, 90, 92, 
    86, 95, 89, 94, 94, 92, 110, 107, 93, 86, 102, 84, 93, 51, 58, 69, 95, 
    86, 89, 80, 97, 74, 64, 62, 57, 52, 53, 59, 51, 63, 72, 102, 93, 88, 87, 
    97, 97, 99, 98, 115, 96, 80, 71, 91, 70, 65, 294, 32, 38, 60, 63, 70, 70, 
    63, 63, 65, 60, 62, 56, 59, 62, 64, 62, 61, 63, 60, 57, 60, 63, 61, 62, 
    67, 65, 63, 61, 63, 60, 55, 50, 53, 54, 55, 51, 52, 53, 53, 51, 53, 50, 
    53, 346, 319, 58, 348, 57, 53, 49, 53, 56, 326, 66, 57, 50, 50, 52, 52, 
    48, 53, 55, 56, 59, 61, 56, 56, 53, 53, 51, 51, 60, 61, 59, 56, 55, 51, 
    52, 54, 52, 52, 52, 49, 51, 57, 56, 59, 55, 53, 51, 49, 50, 48, 46, 47, 
    48, 49, 50, 44, 52, 49, 33, 37, 61, 110, 2, 84, 74, 115, 97, 98, 34, 58, 
    46, 357, 344, 31, 32, 30, 31, 33, 32, 49, 48, 46, 45, 45, 52, 12, 61, 
    101, 110, 115, 66, 58, 64, 58, 54, 48, 52, 51, 51, 53, 53, 51, 48, 51, 
    52, 54, 52, 53, 55, 55, 52, 55, 53, 52, 52, 54, 52, 49, 51, 50, 52, 49, 
    50, 49, 45, 359, 45, 49, 57, 54, 46, 49, 52, 52, 54, 54, 52, 53, 51, 52, 
    50, 50, 56, 56, 56, 51, 51, 51, 52, 54, 55, 54, 57, 57, 57, 57, 68, 69, 
    72, 73, 79, 81, 81, 87, 81, 93, 94, 91, 91, 112, 131, 125, 118, 126, 122, 
    107, 129, 101, 19, 50, 50, 3, 357, 1, 27, 17, 71, 65, 60, 82, 81, 105, 
    123, 113, 114, 111, 115, 117, 109, 109, 107, 102, 111, 117, 138, 149, 
    153, 153, 151, 169, 186, 176, 180, 186, 198, 187, 169, 179, 157, 195, 
    192, 180, 148, 143, 122, 124, 139, 151, 135, 119, 121, 124, 116, 126, 
    114, 160, 180, 202, 326, 332, 330, 355, 347, 349, 331, 322, 299, 325, 23, 
    33, 323, 331, 337, 335, 340, 346, 42, 24, 330, 318, 328, 332, 333, 339, 
    321, 344, 344, 347, 341, 357, 12, 2, 3, 356, 10, 5, 2, 20, 29, 23, 16, 
    23, 23, 9, 9, 9, 2, 6, 18, 18, 22, 18, 22, 24, 32, 22, 17, 26, 31, 19, 
    17, 35, 18, 22, 21, 18, 43, 51, 63, 40, 57, 51, 57, 46, 27, 9, 56, 59, 
    62, 68, 68, 74, 86, 100, 107, 103, 78, 72, 97, 81, 61, 63, 91, 88, 103, 
    55, 55, 38, 35, 47, 51, 49, 46, 43, 54, 81, 117, 122, 60, 61, 62, 70, 66, 
    60, 58, 59, 60, 60, 335, 48, 53, 56, 53, 48, 52, 56, 58, 62, 64, 72, 79, 
    77, 72, 73, 77, 72, 73, 84, 86, 92, 91, 108, 114, 109, 112, 112, 116, 
    109, 114, 130, 128, 131, 129, 131, 124, 126, 126, 122, 116, 135, 129, 
    132, 133, 145, 144, 140, 149, 152, 151, 154, 152, 151, 143, 155, 159, 
    131, 131, 128, 117, 119, 109, 106, 106, 113, 115, 135, 113, 119, 127, 
    124, 120, 102, 107, 120, 120, 122, 144, 130, 129, 127, 137, 130, 101, 
    101, 7, 104, 104, 0, 88, 138, 0, 114, 104, 179, 358, 223, 240, 239, 246, 
    254, 265, 266, 254, 265, 270, 254, 250, 261, 247, 234, 272, 286, 313, 
    277, 303, 305, 318, 318, 310, 303, 291, 305, 185, 112, 125, 112, 110, 
    151, 117, 117, 113, 133, 276, 269, 287, 295, 307, 307, 328, 323, 340, 
    350, 14, 7, 335, 351, 358, 346, 6, 360, 115, 178, 178, 129, 125, 130, 
    135, 118, 118, 114, 116, 139, 154, 153, 159, 119, 113, 104, 103, 128, 
    124, 109, 102, 122, 111, 111, 110, 126, 120, 115, 95, 111, 121, 105, 105, 
    118, 124, 119, 113, 113, 113, 115, 115, 110, 111, 113, 118, 114, 119, 
    114, 115, 118, 115, 120, 115, 122, 131, 114, 114, 126, 109, 92, 107, 111, 
    105, 125, 113, 127, 113, 133, 105, 98, 125, 118, 113, 108, 119, 115, 106, 
    327, 329, 306, 344, 1, 152, 125, 95, 119, 110, 118, 115, 123, 124, 118, 
    130, 149, 295, 290, 287, 277, 291, 286, 291, 295, 293, 277, 291, 286, 
    290, 282, 287, 290, 296, 286, 294, 285, 293, 294, 301, 301, 301, 303, 
    318, 325, 315, 325, 327, 329, 321, 322, 327, 330, 342, 327, 2, 77, 67, 
    66, 70, 70, 77, 76, 84, 132, 114, 123, 118, 114, 108, 108, 116, 115, 111, 
    106, 95, 94, 82, 72, 61, 359, 0, 0, 286, 287, 303, 310, 25, 49, 51, 52, 
    54, 56, 58, 60, 59, 63, 74, 78, 79, 92, 115, 100, 115, 125, 123, 126, 
    128, 133, 138, 143, 136, 121, 112, 121, 110, 113, 128, 137, 127, 114, 
    118, 169, 168, 168, 160, 101, 95, 0, 0, 56, 0, 0, 96, 0, 0, 0, 352, 320, 
    316, 319, 319, 296, 286, 288, 288, 298, 304, 302, 304, 309, 308, 325, 1, 
    68, 86, 110, 101, 98, 75, 61, 67, 63, 52, 60, 58, 61, 62, 61, 66, 65, 69, 
    70, 75, 71, 67, 70, 68, 74, 82, 83, 82, 84, 90, 86, 88, 88, 84, 78, 76, 
    80, 78, 80, 77, 83, 82, 80, 82, 90, 84, 79, 77, 79, 81, 74, 72, 60, 69, 
    97, 118, 137, 140, 162, 170, 166, 165, 168, 159, 159, 160, 138, 126, 129, 
    123, 132, 139, 134, 130, 126, 136, 124, 124, 114, 116, 168, 186, 200, 
    196, 188, 169, 175, 159, 191, 171, 175, 116, 230, 116, 68, 52, 191, 93, 
    95, 104, 103, 92, 90, 98, 84, 92, 93, 90, 73, 91, 88, 86, 86, 82, 79, 91, 
    85, 86, 91, 86, 81, 79, 77, 73, 69, 61, 67, 65, 55, 51, 49, 48, 53, 52, 
    46, 41, 44, 324, 333, 332, 328, 299, 290, 287, 286, 274, 255, 282, 231, 
    208, 178, 172, 155, 129, 129, 161, 155, 112, 101, 109, 114, 103, 116, 
    115, 115, 111, 124, 114, 120, 109, 120, 119, 117, 117, 113, 115, 120, 
    111, 116, 114, 115, 121, 117, 121, 122, 123, 125, 126, 121, 120, 118, 
    116, 122, 115, 127, 119, 125, 114, 115, 125, 123, 114, 119, 123, 124, 
    125, 131, 122, 140, 151, 139, 121, 118, 124, 134, 139, 132, 132, 121, 
    110, 93, 85, 90, 99, 113, 119, 110, 109, 108, 108, 106, 105, 109, 110, 
    108, 110, 110, 111, 108, 104, 103, 98, 97, 96, 97, 98, 99, 98, 90, 90, 
    96, 95, 95, 97, 94, 91, 96, 107, 109, 111, 115, 118, 120, 119, 119, 128, 
    122, 203, 215, 356, 223, 96, 107, 118, 121, 121, 91, 138, 116, 332, 356, 
    344, 335, 333, 105, 41, 108, 123, 123, 109, 105, 127, 127, 137, 108, 102, 
    86, 89, 96, 93, 92, 91, 96, 85, 91, 75, 70, 66, 65, 62, 63, 69, 68, 70, 
    66, 72, 76, 77, 76, 87, 75, 72, 71, 77, 74, 69, 61, 73, 86, 79, 87, 80, 
    72, 68, 69, 73, 79, 82, 87, 82, 95, 101, 103, 105, 108, 101, 94, 104, 96, 
    95, 99, 101, 99, 94, 96, 95, 93, 92, 91, 92, 83, 79, 90, 99, 94, 88, 88, 
    90, 89, 88, 83, 83, 83, 82, 84, 81, 79, 78, 74, 78, 85, 91, 84, 89, 90, 
    89, 89, 89, 84, 83, 88, 100, 90, 90, 94, 93, 90, 91, 94, 100, 102, 90, 
    85, 88, 91, 90, 86, 84, 92, 92, 94, 92, 93, 96, 95, 93, 97, 96, 99, 102, 
    115, 119, 116, 116, 114, 115, 115, 114, 116, 121, 123, 122, 125, 121, 
    122, 128, 124, 125, 120, 118, 117, 116, 124, 123, 120, 116, 120, 113, 
    114, 111, 107, 104, 115, 122, 122, 122, 119, 116, 119, 122, 125, 122, 
    121, 114, 109, 103, 110, 121, 121, 121, 117, 107, 98, 97, 108, 116, 108, 
    110, 104, 109, 113, 116, 110, 106, 104, 106, 112, 109, 106, 100, 98, 102, 
    98, 98, 94, 96, 96, 95, 95, 94, 97, 99, 100, 100, 104, 100, 95, 93, 91, 
    100, 90, 93, 89, 94, 93, 90, 99, 96, 103, 94, 92, 93, 88, 88, 91, 84, 80, 
    80, 77, 78, 96, 105, 105, 101, 91, 86, 82, 84, 83, 82, 78, 79, 83, 85, 
    76, 70, 70, 87, 77, 70, 67, 60, 76, 74, 84, 80, 69, 67, 69, 68, 80, 77, 
    69, 73, 82, 78, 82, 84, 98, 107, 111, 122, 120, 120, 117, 113, 108, 107, 
    108, 109, 108, 115, 108, 108, 108, 102, 95, 97, 95, 100, 101, 94, 103, 
    102, 113, 115, 114, 115, 115, 102, 115, 116, 107, 108, 125, 119, 123, 
    123, 136, 127, 105, 102, 101, 88, 100, 94, 107, 110, 126, 128, 136, 133, 
    109, 108, 102, 100, 109, 112, 116, 127, 118, 188, 170, 175, 167, 174, 
    179, 175, 180, 178, 185, 192, 178, 121, 136, 123, 160, 110, 155, 76, 109, 
    112, 164, 104, 128, 179, 93, 110, 92, 112, 112, 145, 151, 146, 113, 136, 
    110, 135, 127, 128, 225, 227, 244, 254, 227, 213, 209, 197, 209, 216, 
    209, 205, 237, 8, 4, 314, 314, 315, 316, 337, 335, 4, 68, 67, 66, 72, 72, 
    80, 99, 92, 120, 147, 148, 128, 169, 172, 163, 163, 157, 152, 145, 151, 
    161, 181, 104, 153, 143, 123, 111, 98, 81, 85, 84, 82, 92, 77, 82, 83, 
    85, 65, 52, 53, 54, 60, 71, 68, 61, 66, 48, 51, 49, 44, 42, 50, 49, 51, 
    51, 52, 53, 61, 61, 58, 67, 66, 54, 51, 52, 45, 40, 46, 50, 55, 67, 60, 
    60, 61, 72, 66, 56, 55, 50, 38, 49, 44, 41, 42, 44, 39, 42, 43, 34, 31, 
    15, 21, 5, 342, 338, 344, 353, 348, 344, 342, 346, 345, 343, 341, 339, 
    333, 336, 341, 347, 15, 22, 9, 350, 14, 40, 52, 88, 91, 90, 115, 91, 80, 
    77, 78, 99, 110, 139, 226, 300, 294, 297, 295, 302, 308, 309, 322, 342, 
    335, 334, 335, 344, 331, 332, 330, 330, 329, 320, 317, 330, 327, 329, 
    326, 322, 322, 327, 328, 328, 325, 326, 326, 326, 327, 324, 320, 318, 
    316, 317, 317, 310, 319, 317, 320, 317, 312, 319, 319, 311, 325, 330, 
    327, 319, 318, 315, 315, 316, 319, 321, 321, 318, 323, 321, 346, 343, 
    344, 353, 5, 23, 15, 84, 342, 81, 65, 63, 65, 62, 58, 53, 51, 61, 59, 60, 
    62, 78, 91, 95, 105, 112, 132, 125, 128, 134, 130, 129, 130, 135, 135, 
    135, _, _, _, _, _, _, 316, 321, 313, 315, 316, 320, 318, 324, 321, 327, 
    324, 319, 331, 325, 319, 332, 332, 334, 1, 356, 353, 61, 81, 114, 96, 89, 
    206, 206, 212, 210, 187, 162, 149, 154, 141, 132, 126, 129, 146, 168, 
    224, 232, 222, 104, 93, 114, 124, 117, 116, 119, 121, 114, 118, 115, 110, 
    111, 111, 108, 103, 95, 105, 104, 110, 100, 108, 104, 107, 100, 93, 90, 
    88, 89, 96, 97, 93, 93, 92, 88, 92, 105, 106, 99, 96, 96, 91, 88, 83, 87, 
    88, 85, 78, 77, 80, 80, 81, 77, 78, 86, 81, 82, 77, 82, 72, 78, 86, 96, 
    96, 80, 90, 102, 84, 89, 93, 87, 90, 89, 94, 85, 85, 78, 79, 73, 78, 77, 
    83, 80, 76, 79, 85, 87, 79, 86, 80, 77, 69, 57, 69, 65, 57, 48, 32, 14, 
    28, 57, 11, 24, 40, 33, 29, 23, 27, 25, 8, 35, 43, 38, 41, 44, 21, 336, 
    4, 358, 4, 17, 9, 2, 345, 340, 339, 336, 339, 334, 315, 319, 322, 324, 
    323, 321, 302, 304, 303, 310, 313, 309, 325, 331, 321, 328, 332, 339, 
    337, 339, 341, 332, 335, 340, 342, 336, 334, 337, 337, 335, 328, 325, 
    325, 322, 325, 323, 322, 324, 332, 325, 327, 321, 321, 321, 323, 328, 
    324, 331, 337, 343, 318, 335, 339, 341, 343, 357, 1, 343, 345, 359, 344, 
    355, 358, 5, 349, 343, 346, 355, 7, 8, 2, 4, 2, 355, 2, 357, 351, 352, 
    360, 27, 15, 360, 341, 332, 329, 326, 330, 329, 321, 325, 320, 319, 312, 
    319, 321, 326, 334, 335, 334, 332, 335, 334, 328, 328, 330, 329, 332, 
    329, 326, 325, 327, 327, 322, 322, 324, 313, 316, 317, 318, 320, 319, 
    319, 316, 320, 317, 312, 305, 313, 313, 312, 316, 323, 323, 322, 324, 
    318, 324, 323, 324, 325, 322, 320, 320, 322, 317, 324, 319, 314, 322, 
    318, 323, 317, 316, 316, 317, 316, 321, 331, 331, 329, 330, 331, 326, 
    328, 331, 329, 332, 318, 317, 318, 322, 320, 320, 316, 317, 318, 323, 
    325, 325, 325, 330, 324, 333, 330, 325, 324, 320, 320, 325, 326, 322, 
    321, 323, 319, 331, 317, 321, 326, 327, 314, 316, 321, 323, 311, 329, 
    319, 311, 318, 332, 331, 338, 334, 337, 328, 334, 325, 316, 318, 311, 
    323, 347, 360, 352, 346, 350, 347, 336, 335, 338, 333, 334, 329, 329, 
    336, 346, 335, 8, 25, 14, 353, 8, 15, 74, 85, 278, 2, 2, 328, 60, 61, 53, 
    66, 62, 42, 33, 353, 18, 2, 8, 4, 344, 339, 32, 347, 8, 359, 347, 336, 
    319, 344, 330, 333, 322, 329, 307, 328, 319, 354, 277, 292, 353, 9, 360, 
    343, 335, 346, 359, 339, 355, 344, 336, 355, 349, 345, 349, 337, 335, 
    334, 318, 318, 328, 313, 288, 259, 241, 285, 267, 259, 257, 253, 250, 
    245, 253, 252, 255, 252, 249, 245, 255, 245, 245, 244, 250, 246, 245, 
    247, 242, 241, 232, 236, 236, 243, 243, 245, 250, 255, 257, 301, 287, 
    312, 328, 325, 320, 306, 298, 288, 322, 318, 316, 311, 307, 313, 294, 
    311, 320, 326, 315, 300, 309, 316, 311, 316, 311, 311, 308, 303, 306, 
    311, 331, 329, 334, 334, 333, 334, 336, 328, 329, 336, 348, 326, 327, 
    328, 360, 7, 360, 27, 72, 112, 89, 55, 8, 15, 36, 65, 128, 136, 142, 138, 
    142, 143, 138, 134, 141, 130, 127, 121, 121, 118, 107, 112, 112, 111, 
    154, 307, 319, 321, 286, 293, 280, 278, 277, 264, 253, 246, 248, 286, 
    300, 301, 308, 292, 307, 331, 324, 327, 319, 324, 324, 323, 323, 324, 
    325, 325, 320, 315, 318, 312, 316, 308, 310, 309, 314, 322, 322, 317, 
    322, 324, 313, 313, 323, 323, 325, 328, 321, 322, 325, 316, 306, 292, 
    304, 298, 315, 323, 332, 329, 322, 321, 318, 318, 317, 324, 323, 323, 
    322, 321, 320, 320, 315, 315, 314, 314, 317, 318, 319, 319, 311, 310, 
    313, 313, 315, 321, 321, 325, 323, 321, 328, 320, 313, 318, 315, 309, 
    310, 312, 322, 317, 314, 314, 317, 301, 299, 307, 305, 311, 329, 326, 
    319, 319, 316, 315, 310, 313, 309, 310, 318, 316, 321, 321, 317, 321, 
    323, 319, 318, 320, 317, 313, 331, 331, 329, 326, 324, 321, 327, 328, 
    325, 320, 292, 292, 298, 305, 301, 302, 296, 290, 291, 270, 255, 276, 
    257, 249, 254, 269, 273, 252, 253, 292, 291, 266, 253, 239, 258, 251, 
    262, 255, 258, 236, 230, 252, 258, 232, 226, 229, 223, 237, 248, 265, 
    257, 257, 245, 269, 267, 259, 356, 4, 2, 276, 15, 351, 327, 336, 353, 
    335, 328, 327, 330, 351, 336, 325, 325, 326, 322, 323, 332, 327, 333, 
    327, 330, 324, 333, 334, 329, 332, 331, 331, 329, 329, 330, 329, 330, 
    332, 335, 334, 343, 330, 340, 343, 355, 346, 350, 352, 348, 342, 342, 
    347, 359, 355, 347, 343, 335, 335, 321, 323, 329, 333, 329, 334, 330, 
    331, 350, 3, 2, 356, 349, 345, 349, 348, 343, 347, 354, 4, 10, 344, 323, 
    322, 324, 36, 53, 87, 102, 110, 146, 143, 141, 136, 151, 151, 136, 131, 
    137, 140, 143, 132, 141, 126, 101, 281, 344, 319, 311, 324, 322, 324, 
    321, 325, 17, 55, 58, 57, 49, 60, 56, 60, 55, 56, 56, 50, 53, 47, 51, 52, 
    45, 61, 353, 3, 13, 319, 322, 330, 329, 325, 324, 307, 23, 19, 26, 12, 
    19, 338, 330, 337, 340, 347, 19, 177, 308, 339, 325, 328, 314, 304, 324, 
    326, 327, 5, 90, 58, 56, 60, 60, 335, 2, 3, 360, 349, 339, 316, 320, 326, 
    320, 313, 318, 318, 331, 325, 331, 322, 320, 324, 334, 335, 331, 333, 
    331, 336, 339, 340, 320, 308, 309, 312, 1, 351, 344, 332, 319, 317, 320, 
    333, 324, 329, 334, 334, 337, 340, 344, 350, 1, 350, 342, 346, 343, 332, 
    333, 338, 313, 336, 336, 279, 235, 246, 217, 197, 203, 204, 248, 253, 
    289, 276, 288, 285, 313, 303, 311, 312, 310, 296, 310, 316, 316, 309, 
    304, 280, 206, 121, 109, 170, 163, 153, 156, 170, 170, 179, 134, 124, 
    114, 121, 94, 124, 100, 111, 102, 102, 102, 97, 100, 121, 113, 110, 112, 
    109, 100, 86, 81, 60, 78, 100, 99, 109, 109, 104, 102, 99, 94, 80, 75, 
    62, 54, 55, 58, 65, 54, 42, 326, 312, 288, 294, 305, 288, 293, 298, 297, 
    292, 293, 297, 296, 302, 301, 291, 300, 296, 304, 295, 292, 289, 291, 
    301, 294, 289, 292, 291, 293, 288, 287, 253, 251, 246, 256, 271, 263, 
    265, 249, 275, 284, 279, 270, 291, 285, 277, 278, 277, 293, 292, 289, 
    293, 302, 286, 286, 301, 285, 283, 297, 293, 292, 302, 291, 290, 289, 
    294, 293, 299, 292, 290, 290, 286, 285, 284, 279, 278, 281, 274, 276, 
    277, 272, 279, 289, 316, 328, 351, 38, 79, 78, 109, 130, 254, 269, 274, 
    273, 267, 274, 298, 315, 318, 310, 319, 315, 321, 320, 305, 306, 304, 
    300, 298, 300, 314, 301, 301, 299, 312, 315, 319, 312, 310, 313, 306, 
    308, 306, 309, 310, 314, 312, 313, 315, 317, 315, 317, 314, 320, 316, 
    294, 318, 307, 314, 305, 317, 312, 313, 318, 301, 307, 304, 314, 311, 
    324, 324, 307, 325, 318, 316, 325, 329, 315, 309, 309, 313, 313, 309, 
    311, 307, 304, 303, 301, 300, 290, 296, 300, 306, 311, 317, 325, 322, 
    319, 320, 309, 311, 299, 299, 306, 312, 310, 314, 308, 311, 314, 313, 
    306, 300, 299, 294, 303, 294, 305, 304, 305, 297, 295, 296, 299, 320, 
    317, 311, 305, 303, 300, 312, 313, 312, 309, 305, 307, 305, 305, 306, 
    304, 303, 302, 299, 295, 295, 299, 307, 309, 300, 303, 303, 312, 299, 
    298, 310, 299, 330, 325, 323, 331, 360, 4, 16, 27, 8, 53, 56, 50, 54, 87, 
    73, 81, 95, 106, 63, 48, 13, 347, 24, 3, 28, 337, 335, 323, 324, 319, 
    325, 323, 318, 325, 305, 309, 320, 311, 303, 303, 308, 306, 315, 320, 
    326, 326, 329, 330, 330, 331, 336, 332, 349, 358, 356, 350, 356, 357, 
    353, 352, 345, 343, 345, 355, 347, 349, 352, 356, 351, 351, 359, 360, 1, 
    357, 8, 9, 32, 31, 37, 32, 38, 37, 41, 35, 41, 44, 42, 49, 42, 35, 14, 
    31, 42, 38, 29, 33, 26, 27, 27, 42, 39, 32, 21, 16, 13, 3, 14, 33, 36, 
    38, 27, 21, 356, 28, 16, 16, 16, 15, 25, 21, 15, 3, 346, 7, 1, 1, 351, 7, 
    353, 353, 353, 345, 338, 338, 330, 330, 322, 320, 316, 309, 324, 334, 
    327, 324, 329, 325, 325, 331, 327, 322, 328, 329, 320, 315, 322, 322, 
    330, 336, 334, 336, 336, 336, 330, 320, 312, 331, 304, 308, 312, 320, 
    307, 312, 302, 316, 305, 326, 323, 316, 331, 321, 320, 296, 327, 334, 
    346, 355, 300, 271, 105, 84, 117, 118, 119, 121, 121, 138, 134, 134, 121, 
    128, 131, 133, 125, 122, 120, 132, 115, 115, 127, 110, 108, 115, 109, 
    111, 111, 113, 107, 119, 105, 117, 120, 124, 112, 123, 113, 108, 121, 
    132, 126, 133, 124, 52, 6, 157, 102, 119, 126, 117, 115, 115, 128, 122, 
    119, 116, 121, 119, 130, 121, 126, 134, 114, 114, 119, 115, 116, 117, 
    105, 133, 150, 266, 279, 293, 274, 281, 284, 285, 290, 290, 290, 280, 
    285, 270, 285, 281, 264, 283, 270, 277, 291, 321, 353, 280, 309, 314, 
    320, 326, 324, 332, 286, 281, 272, 270, 281, 296, 285, 290, 349, 325, 
    325, 326, 323, 312, 310, 325, 308, 297, 294, 296, 306, 304, 312, 274, 
    246, 238, 260, 303, 283, 289, 296, 300, 304, 293, 284, 265, 262, 258, 
    270, 237, 290, 278, 249, 284, 275, 269, 268, 265, 256, 303, 277, 251, 
    310, 301, 341, 331, 328, 21, 24, 33, 33, 24, 35, 13, 2, 8, 16, 19, 20, 
    35, 48, 52, 45, 47, 42, 18, 23, 33, 18, 42, 220, 27, 17, 11, 348, 349, 
    353, 304, 328, 35, 34, 23, 330, 330, 328, 344, 1, 13, 306, 332, 335, 337, 
    3, 310, 320, 332, 10, 357, 6, 7, 2, 2, 357, 11, 324, 317, 310, 300, 323, 
    309, 305, 308, 311, 331, 354, 354, 348, 347, 341, 335, 317, 323, 333, 
    312, 314, 310, 313, 308, 292, 281, 302, 302, 306, 302, 297, 296, 296, 
    297, 306, 305, 266, 312, 293, 310, 245, 250, 201, 173, 186, 78, 112, 60, 
    43, 75, 97, 108, 113, 125, 152, 154, 132, 126, 135, 153, 140, 128, 134, 
    116, 113, 115, 106, 109, 109, 117, 120, 121, 150, 148, 152, 149, 154, 
    151, 152, 153, 166, 163, 235, 255, 259, 257, 272, 280, 298, 305, 304, 
    306, 309, 320, 310, 307, 317, 315, 314, 314, 311, 307, 300, 307, 297, 
    295, 302, 302, 285, 290, 300, 293, 297, 288, 269, 284, 287, 300, 316, 
    303, 261, 276, 286, 276, 287, 300, 331, 324, 316, 319, 346, 33, 122, 102, 
    117, 157, 161, 170, 174, 183, 204, 159, 217, 311, 305, 296, 295, 327, 
    282, 284, 273, 274, 279, 259, 249, 248, 248, 252, 238, 237, 223, 216, 
    216, 265, 274, 251, 252, 247, 252, 243, 235, 235, 240, 281, 277, 276, 
    281, 290, 286, 290, 291, 299, 301, 292, 298, 294, 285, 285, 284, 279, 
    291, 295, 285, 281, 276, 281, 276, 288, 298, 313, 301, 298, 297, 290, 
    288, 288, 289, 286, 297, 282, 285, 293, 284, 299, 289, 303, 286, 281, 
    295, 297, 294, 294, 297, 293, 292, 288, 303, 325, 310, 313, 314, 309, 
    310, 309, 313, 333, 325, 345, 327, 330, 329, 329, 331, 337, 326, 329, 
    326, 317, 316, 317, 326, 326, 317, 321, 321, 321, 322, 314, 309, 315, 
    310, 314, 317, 317, 320, 315, 317, 320, 320, 321, 328, 328, 323, 325, 
    320, 319, 323, 324, 321, 324, 325, 318, 321, 322, 321, 313, 310, 317, 
    320, 314, 322, 318, 320, 323, 325, 309, 314, 320, 311, 319, 312, 314, 
    307, 320, 306, 268, 108, 88, 89, 127, 181, 152, 161, 126, 138, 143, 144, 
    127, 133, 127, 122, 128, 111, 96, 101, 102, 122, 119, 122, 112, 110, 108, 
    94, 181, 147, 77, 317, 320, 300, 281, 265, 247, 259, 255, 285, 290, 302, 
    303, 310, 331, 307, 310, 327, 318, 329, 316, 264, 278, 291, 356, 0, 128, 
    136, 125, 115, 124, 114, 139, 130, 158, 243, 0, 142, 106, 125, 119, 108, 
    120, 129, 112, 127, 121, 115, 117, 126, 128, 120, 133, 135, 142, 353, 
    300, 323, 310, 308, 304, 320, 321, 346, 318, 321, 132, 114, 314, 325, 
    318, 321, 324, 324, 324, 309, 322, 329, 333, 331, 302, 308, 314, 301, 
    286, 285, 274, 304, 310, 311, 329, 331, 316, 300, 284, 281, 318, 300, 
    305, 301, 298, 323, 320, 308, 320, 299, 304, 279, 291, 296, 280, 290, 
    279, 285, 293, 287, 307, 293, 295, 312, 298, 304, 299, 331, 288, 300, 
    343, 252, 227, 141, 136, 117, 120, 123, 143, 126, 116, 104, 102, 97, 107, 
    108, 101, 101, 100, 145, 59, 273, 277, 290, 307, 323, 302, 304, 291, 289, 
    294, 296, 296, 300, 305, 306, 307, 303, 299, 284, 304, 322, 300, 302, 
    296, 300, 303, 329, 303, 311, 310, 331, 323, 259, 352, 360, 90, 142, 139, 
    139, 135, 132, 118, 113, 115, 126, 134, 144, 161, 166, 175, 167, 160, 
    152, 130, 129, 137, 133, 134, 135, 127, 118, 112, 112, 113, 115, 115, 
    116, 114, 112, 109, 105, 102, 112, 98, 89, 279, 263, 306, 323, 308, 301, 
    308, 345, 310, 318, 320, 320, 334, 314, 326, 312, 309, 309, 312, 314, 
    320, 277, 6, 228, 184, 99, 141, 124, 125, 116, 116, 124, 121, 114, 114, 
    118, 126, 124, 121, 116, 118, 116, 115, 116, 131, 134, 131, 132, 123, 
    113, 113, 114, 115, 113, 123, 118, 116, 221, 313, 310, 321, 317, 302, 
    305, 287, 284, 278, 279, 280, 288, 282, 282, 281, 296, 296, 287, 297, 
    308, 309, 311, 309, 297, 317, 293, 315, 296, 7, 287, 319, 37, 40, 103, 
    118, 113, 105, 99, 105, 58, 59, 57, 52, 61, 56, 49, 37, 8, 18, 327, 320, 
    6, 327, 323, 321, 328, 330, 316, 315, 317, 296, 314, 291, 298, 305, 305, 
    323, 273, 284, 303, 249, 353, 87, 105, 187, 163, 154, 157, 148, 131, 167, 
    190, 128, 256, 286, 302, 296, 309, 298, 314, 310, 320, 315, 312, 306, 
    299, 300, 292, 291, 288, 289, 267, 279, 272, 264, 257, 258, 253, 260, 
    258, 260, 264, 264, 277, 222, 239, 174, 180, 185, 200, 210, 237, 244, 
    247, 242, 238, 321, 307, 290, 282, 272, 280, 271, 264, 255, 224, 246, 
    241, 212, 220, 237, 207, 198, 178, 240, 248, 247, 324, 69, 47, 48, 16, 
    55, 36, 355, 350, 344, 326, 321, 325, 5, 5, 360, 33, 36, 36, 35, 27, 31, 
    19, 25, 26, 30, 35, 27, 285, 337, 17, 14, 327, 60, 55, 57, 63, 65, 102, 
    89, 100, 98, 103, 128, 111, 125, 112, 103, 109, 108, 120, 119, 96, 98, 
    102, 101, 98, 92, 96, 90, 85, 78, 87, 82, 77, 70, 70, 64, 62, 25, 31, 23, 
    10, 24, 4, 4, 349, 356, 349, 346, 346, 343, 341, 339, 336, 334, 328, 326, 
    335, 330, 330, 317, 319, 336, 329, 320, 319, 318, 312, 307, 306, 303, 
    300, 300, 295, 297, 294, 291, 292, 293, 289, 288, 282, 290, 290, 290, 
    272, 292, 296, 304, 298, 289, 298, 307, 300, 311, 302, 311, 317, 323, 
    323, 319, 316, 317, 308, 308, 320, 321, 330, 329, 330, 335, 319, 322, 
    330, 318, 316, 307, 313, 312, 323, 327, 313, 312, 307, 299, 310, 311, 
    312, 322, 315, 318, 317, 317, 310, 309, 331, 325, 318, 316, 330, 353, 
    317, 329, 340, 321, 316, 315, 320, 315, 317, 315, 332, 320, 317, 328, 
    332, 331, 325, 319, 316, 315, 312, 313, 299, 300, 305, 283, 305, 289, 
    284, 291, 286, 287, 283, 294, 295, 302, 275, 280, 287, 314, 317, 329, 
    335, 339, 308, 298, 300, 322, 322, 329, 326, 327, 317, 332, 329, 323, 
    328, 317, 321, 325, 310, 311, 321, 300, 0, 360, 1, 94, 116, 117, 120, 
    295, 300, 311, 287, 302, 317, 351, 322, 323, 321, 314, 233, 305, 286, 
    309, 0, 331, 321, 355, 38, 70, 360, 355, 5, 360, 0, 125, 119, 152, 129, 
    84, 73, 66, 60, 69, 76, 77, 79, 87, 94, 129, 147, 146, 149, 134, 131, 96, 
    155, 83, 85, 132, 185, 163, 144, 114, 134, 112, 95, 131, 131, 111, 124, 
    116, 130, 114, 76, 125, 146, 145, 139, 120, 115, 159, 150, 125, 126, 116, 
    106, 116, 109, 118, 122, 129, 122, 124, 130, 153, 135, 128, 127, 170, 
    140, 131, 150, 165, 152, 140, 175, 128, 123, 151, 119, 119, 116, 119, 
    118, 119, 119, 121, 130, 121, 120, 128, 128, 123, 118, 121, 119, 118, 
    123, 127, 86, 77, 73, 59, 56, 58, 61, 58, 51, 51, 56, 60, 68, 81, 106, 
    105, 104, 111, 109, 111, 113, 110, 110, 111, 115, 116, 112, 111, 110, 
    110, 107, 106, 104, 103, 105, 105, 106, 103, 104, 104, 105, 104, 101, 
    101, 101, 100, 95, 95, 98, 72, 17, 314, 314, 325, 313, 276, 282, 127, 
    307, 3, 280, 163, 355, 30, 186, 194, 140, 145, 159, 141, 140, 140, 136, 
    137, 137, 137, 138, 135, 139, 135, 132, 143, 138, 141, 135, 141, 145, 
    146, 134, 129, 98, 133, 133, 139, 123, 130, 135, 125, 129, 147, 132, 127, 
    135, 136, 143, 129, 132, 221, 273, 284, 287, 310, 317, 316, 311, 307, 
    286, 297, 299, 289, 280, 277, 272, 272, 271, 274, 283, 275, 275, 276, 
    257, 265, 282, 282, 277, 278, 302, 312, 323, 233, 12, 131, 149, 144, 91, 
    103, 109, 65, 129, 98, 118, 143, 133, 132, 120, 124, 132, 141, 143, 114, 
    116, 117, 126, 114, 115, 123, 345, 320, 297, 302, 313, 312, 317, 312, 
    315, 309, 294, 308, 316, 317, 315, 323, 342, 328, 320, 318, 323, 326, 
    317, 324, 327, 319, 329, 319, 320, 307, 313, 318, 331, 327, 321, 317, 
    313, 324, 328, 305, 314, 310, 307, 312, 308, 309, 318, 24, 127, 122, 108, 
    129, 119, 129, 118, 121, 119, 116, 120, 122, 121, 118, 117, 115, 117, 
    126, 125, 121, 343, 315, 20, 143, 164, 307, 321, 339, 325, 344, 341, 335, 
    333, 298, 359, 97, 135, 120, 72, 77, 81, 88, 85, 90, 87, 95, 120, 155, 
    272, 320, 317, 321, 315, 319, 324, 324, 319, 328, 315, 318, 321, 324, 
    324, 269, 279, 303, 282, 271, 191, 43, 90, 118, 319, 313, 332, 184, 294, 
    322, 320, 303, 301, 305, 306, 300, 295, 293, 287, 281, 293, 286, 285, 
    271, 267, 276, 273, 279, 281, 289, 293, 291, 280, 277, 280, 280, 279, 
    277, 283, 286, 285, 284, 282, 283, 283, 284, 282, 280, 282, 280, 285, 
    280, 282, 284, 285, 283, 281, 283, 288, 279, 279, 276, 277, 281, 287, 
    284, 284, 286, 287, 286, 286, 285, 285, 291, 294, 293, 293, 288, 301, 
    305, 303, 310, 316, 306, 314, 287, 290, 316, 312, 279, 267, 244, 251, 
    206, 179, 141, 152, 129, 114, 118, 122, 118, 119, 121, 115, 111, 122, 
    117, 118, 119, 120, 118, 120, 126, 120, 118, 123, 118, 117, 120, 124, 
    118, 121, 121, 121, 122, 122, 128, 121, 127, 134, 117, 114, 116, 122, 
    116, 123, 123, 126, 116, 121, 187, 220, 17, 323, 316, 315, 303, 311, 317, 
    312, 305, 307, 314, 306, 316, 312, 302, 313, 326, 319, 302, 61, 359, 339, 
    130, 185, 149, 146, 117, 136, 130, 122, 124, 114, 117, 136, 124, 130, 
    146, 145, 153, 175, 254, 155, 137, 134, 140, 130, 143, 112, 101, 108, 
    120, 113, 116, 118, 126, 259, 325, 332, 324, 326, 339, 321, 312, 196, 
    138, 67, 238, 270, 310, 308, 329, 321, 97, 109, 115, 128, 120, 118, 116, 
    118, 123, 116, 145, 136, 124, 280, 299, 334, 330, 328, 314, 331, 329, 
    329, 309, 315, 311, 305, 310, 305, 306, 297, 301, 304, 296, 302, 286, 
    276, 272, 276, 287, 289, 311, 309, 313, 294, 146, 152, 109, 130, 127, 
    121, 123, 120, 116, 116, 124, 119, 118, 120, 116, 115, 112, 112, 110, 
    114, 115, 116, 115, 117, 116, 110, 121, 137, 122, 135, 133, 125, 101, 
    322, 93, 81, 45, 328, 343, 118, 94, 37, 132, 316, 257, 159, 323, 311, 
    345, 311, 304, 351, 252, 172, 288, 267, 314, 309, 315, 349, 327, 329, 
    322, 314, 317, 320, 323, 316, 318, 318, 318, 324, 306, 317, 298, 314, 
    316, 305, 290, 289, 309, 314, 315, 322, 322, 316, 307, 296, 186, 151, 
    115, 109, 137, 131, 120, 115, 117, 107, 113, 116, 115, 117, 114, 114, 
    118, 120, 132, 172, 275, 279, 306, 320, 321, 331, 315, 319, 334, 317, 
    316, 319, 323, 313, 317, 312, 319, 307, 312, 304, 300, 314, 312, 324, 
    318, 323, 317, 312, 315, 313, 310, 325, 321, 317, 326, 316, 305, 319, 
    315, 305, 301, 303, 323, 319, 321, 318, 320, 314, 313, 316, 322, 321, 
    323, 311, 314, 309, 299, 308, 316, 300, 296, 292, 286, 277, 303, 302, 
    291, 299, 295, 291, 283, 284, 288, 278, 266, 282, 267, 257, 261, 250, 
    251, 263, 269, 264, 264, 262, 252, 245, 249, 246, 248, 245, 245, 238, 
    237, 232, 227, 214, 215, 210, 204, 193, 200, 191, 201, 185, 184, 183, 
    180, 185, 174, 171, 161, 154, 164, 156, 152, 156, 357, 156, 219, 265, 
    314, 316, 322, 327, 316, 301, 299, 304, 299, 284, 266, 259, 282, 268, 
    256, 231, 222, 225, 224, 223, 239, 251, 259, 265, 274, 277, 285, 291, 
    293, _, _, 287, 285, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 288, 278, _, 296, 308, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, 311, 327, 323, 319, 322, _, _, _, 311, _, 315, 329, 316, 308, 
    295, 298, 300, 300, 300, 310, 307, 297, 300, 297, 310, 300, 303, 297, 
    303, 303, 305, 328, 315, 316, 310, 315, 320, 340, 347, 354, 355, 359, 
    338, 326, 325, 330, 320, 315, 315, 311, 315, 308, 324, 320, 320, 302, 
    291, 299, 304, 312, 317, 314, 318, 320, 315, 310, 305, 302, 289, 291, 
    284, 283, 283, 289, 291, 289, 291, 285, 295, 302, 303, 299, _, _, _, _, 
    _, _, 284, 287, 291, _, 295, _, 292, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 317, 313, _, 303, 325, 354, _, _, _, _, _, 203, 164, 146, 150, 
    167, 281, 325, 135, 266, 145, _, _, _, _, _, _, _, _, 146, 161, _, 128, 
    111, _, 127, 123, 136, 134, _, _, 139, 146, _, _, 101, 140, 124, 112, 
    128, _, 177, 153, _, _, _, _, 18, 24, 323, 322, 320, 317, 316, 310, 310, 
    334, _, 325, 326, 317, 320, 329, 322, 315, 314, 314, 313, 313, 312, 311, 
    311, 310, 309, 312, 316, 286, 302, 317, 308, 312, 315, 323, 321, 321, 
    324, 325, 325, 324, 327, 306, 300, 305, 299, 297, 328, 311, 313, 300, 
    305, 301, 304, 315, 318, 321, 322, 322, 330, 325, 319, 318, 305, 315, 
    311, 316, 328, 331, 322, _, 335, 327, 319, 313, 341, 337, 331, 330, 337, 
    _, _, _, 330, 313, 331, 323, 331, 319, 322, 326, _, _, _, _, 325, 326, 
    327, 323, 335, 322, 318, 334, 319, 317, 327, 315, 316, 313, 324, 327, 
    322, 312, 308, 309, 312, 313, 313, 312, 313, 316, 314, _, 310, 312, 311, 
    306, _, _, 312, 306, 306, _, 303, 305, 304, 300, 307, 307, 307, 303, 313, 
    _, 320, 319, 325, 321, 325, 329, _, _, 310, 318, _, _, _, _, _, _, _, _, 
    _, 316, 317, 311, 312, 318, 324, 316, 315, 317, 315, 315, 299, 304, 302, 
    302, 314, 300, _, _, _, _, _, _, _, 305, 302, _, _, 298, 295, 295, 306, 
    _, 315, 316, 321, 309, _, 327, 314, 314, 311, _, _, 319, 322, 316, 314, 
    300, 298, 292, 303, _, 304, 304, 304, 308, _, 309, 306, 306, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 292, 293, 295, 299, 302, 309, 312, 310, 319, 
    318, 316, _, _, _, _, _, 321, 319, _, 319, 319, 323, 333, 331, _, _, 337, 
    327, 316, 304, 309, 307, _, 302, _, _, _, _, _, _, _, _, 282, 290, 291, 
    _, 301, 307, 307, 302, _, 296, _, _, 294, 293, 294, 293, 293, 290, 289, 
    285, _, _, _, 281, 285, 320, 311, 312, 307, 314, _, _, _, 298, 309, 323, 
    298, 304, 301, 300, 300, 300, _, _, 300, 300, 300, 312, 349, 350, 0, 300, 
    0, _, 300, 300, 300, 300, 139, 143, 137, 143, _, 153, 160, 148, 127, 128, 
    133, 137, 138, _, _, _, _, _, 79, 97, 83, 86, 78, 79, 90, 93, 102, 96, 
    108, _, _, 107, _, 108, 110, 110, 106, 105, 106, 108, _, 109, 109, 105, 
    114, 117, 117, 113, 118, _, 118, 112, 117, 112, 111, 111, 110, 112, 116, 
    116, 114, 114, 113, 124, 124, 124, 124, 131, 148, 135, 121, 138, 324, 
    275, 340, 316, 297, 302, 271, 263, 229, 255, 218, 261, 275, 239, 277, 
    264, 259, 266, 271, 269, 278, 273, 271, 275, 276, 278, 286, 282, 281, 
    275, 271, 270, 260, 290, 232, 118, 119, 134, 111, 126, 113, 122, 125, 
    122, 136, 134, 294, 285, 261, 231, 261, 248, 256, 259, 257, 255, 254, 
    270, 291, 291, 290, 309, 320, 322, 301, 284, 284, 301, 284, 280, 276, 
    279, 283, 286, 288, 283, 282, 282, 288, 293, 311, 296, 310, 297, 316, 
    310, 303, 326, 326, 320, 319, 341, 305, 336, 325, 334, 320, 306, 18, 337, 
    302, 80, 76, 151, 56, 79, 87, 96, 104, 112, 111, 110, 96, 111, 96, 83, 
    76, 75, 80, 144, 207, 256, 318, 302, 317, 286, 303, 270, 313, 320, 320, 
    140, 130, 140, 110, 120, 190, 100, 60, 51, 53, 55, 56, 59, 44, 91, 85, 
    111, 106, 101, 97, 92, 87, 82, 78, 73, 68, 77, 88, 87, 70, 68, 39, 78, 
    57, 35, 14, 11, 85, 106, 122, 108, 113, 128, _, _, _, _, _, _, 124, 113, 
    112, 116, 112, 117, 111, 111, _, _, _, _, _, 114, 116, 116, 115, 115, 
    114, 114, _, _, _, _, 115, 115, 117, 52, 293, 308, 308, 317, 320, _, _, 
    _, _, _, _, 311, 308, 303, 311, 308, 308, 300, 296, _, _, _, _, 309, 302, 
    305, 308, 301, 308, 308, 289, _, 285, 285, 297, 302, 296, 300, 294, 265, 
    _, _, 240, 234, 227, 237, 180, 157, 130, 160, _, _, 106, 106, 106, 100, 
    109, 92, 83, 66, _, 46, 44, 49, 48, 38, 34, 21, 13, _, _, _, _, _, _, 
    353, 360, _, 337, 305, _, 324, 308, 319, 339, 320, 331, 342, 22, 30, 33, 
    332, _, _, _, _, _, _, _, _, 339, 53, 254, 20, 181, 104, 0, 75, _, 317, 
    302, 319, 292, 326, 309, 302, 311, _, _, _, _, 314, 322, 316, 307, 321, 
    317, 320, 329, _, 333, 331, 321, 315, 264, 257, 101, 112, _, _, _, 108, 
    110, 114, 103, 101, 99, 94, 103, _, _, _, 121, 117, 116, 123, 110, 117, 
    118, 114, 112, _, _, _, 105, 108, 111, 106, 114, 104, 125, 110, _, 120, 
    115, 70, 244, 288, 289, 286, 291, 287, 290, 287, 290, 293, 295, 294, _, 
    _, _, 286, 291, 291, 297, 308, 321, 305, 311, _, 301, 321, 317, 313, 305, 
    305, 304, 292, 301, 288, _, _, _, _, 101, 112, 110, 110, 115, 113, 116, 
    112, _, _, _, 112, 114, 111, 106, 112, 117, 125, 118, _, _, _, 115, 119, 
    115, 112, 121, 125, 115, 114, 117, _, _, _, 101, 132, 122, 131, 312, 322, 
    299, 314, _, _, _, 226, 215, 204, 220, 222, 224, 231, 229, _, _, _, 262, 
    262, 246, 276, 280, 281, 276, 279, _, _, _, _, _, _, _, _, 218, 210, 197, 
    197, 196, 193, 190, 187, _, _, 140, 120, 110, 60, 45, 51, 52, 49, _, _, 
    _, _, _, _, _, _, _, _, 52, 65, 56, _, _, _, 345, 13, 1, _, 356, _, _, 
    355, _, 292, _, _, _, 340, 6, 8, 357, _, _, 36, _, _, 43, 43, _, 27, 25, 
    _, _, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, 26, 25, 24, 57, 180, 
    155, _, _, _, _, _, 193, 156, _, 142, 142, 135, 143, 153, _, _, 159, 154, 
    147, _, 143, 141, 148, 159, _, _, 154, 147, 137, 140, 132, 144, 119, _, 
    117, 115, 123, 144, 154, 139, 139, 150, _, 119, _, 128, 128, 127, 125, 
    126, 125, 127, 131, 121, 133, 122, 117, 117, 127, _, _, 134, 128, _, _, 
    133, 117, 119, 118, _, _, 120, 120, 116, 111, 117, 101, 94, 87, 88, _, _, 
    _, 71, 71, 62, _, _, _, 60, 69, 65, 70, 61, 58, 56, _, 56, 51, 44, 42, 
    45, 44, 43, 181, _, _, _, 0, 324, 299, _, 352, 315, 325, 333, 326, 333, 
    336, _, 323, _, 332, _, _, _, _, _, 320, 322, _, 314, _, 310, _, 308, 
    310, _, 307, 300, 299, 301, _, _, _, _, _, _, 300, _, 300, _, 295, _, 
    296, _, _, _, 298, 293, 295, 295, 319, 322, 316, 318, _, 323, 331, 332, 
    _, 323, 327, 325, 323, _, _, 308, 306, 312, 306, 309, 302, 291, _, 296, 
    _, _, _, 304, 311, 317, 292, 329, 257, 230, 238, _, _, 187, _, _, 212, 
    287, 288, _, 274, _, _, _, _, _, _, _, _, 245, 244, 240, 241, 240, 226, 
    228, _, 239, 243, 125, 124, 109, 103, 123, _, _, _, _, 95, 84, _, 69, 76, 
    _, 77, 76, 76, 71, _, 68, _, 45, 47, 45, 293, _, _, 145, 139, 21, _, _, 
    _, 252, 252, 250, 251, 260, 267, 279, 288, _, 291, _, 317, _, _, 324, _, 
    _, _, 0, 307, 327, 108, 338, 18, 354, 284, 49, _, 58, _, 63, _, 71, 71, 
    72, 80, _, _, _, 91, 91, 99, 105, 113, 138, 114, 116, _, _, _, _, _, _, 
    _, _, _, _, 116, 118, 123, 125, 115, 100, 81, 76, _, _, 85, _, 301, 311, 
    _, 305, 304, _, _, _, _, 273, _, 267, 260, 265, 271, _, _, 278, _, _, 
    267, _, 273, 275, 277, 276, 276, 281, _, _, _, 289, _, _, _, 303, 311, 
    316, 319, 324, 324, 327, 327, 331, _, _, _, _, 337, 333, 331, 336, 346, 
    337, 339, 360, _, 15, 11, 1, 10, 10, 14, 24, 32, 326, 38, 39, 37, 41, 52, 
    63, 59, 61, _, _, _, _, 62, 63, _, 75, 77, 97, 155, 153, 165, 160, 143, 
    _, _, _, _, 162, 153, 150, 153, 161, 172, 133, 139, _, _, 251, 281, 317, 
    318, 321, 314, 324, 315, _, _, 302, 301, 309, 297, 293, 295, 299, 304, _, 
    _, 287, 285, 303, 299, 304, 294, 318, 317, _, _, 316, 321, 320, 329, 325, 
    333, 335, 328, _, _, 360, 339, 334, 327, 316, 301, 311, 321, _, _, _, _, 
    316, 334, 322, 313, 315, 321, _, _, 327, 310, 323, 306, 312, 314, 325, 
    324, _, _, 319, 324, 321, 324, 302, 303, _, 317, 316, _, _, 320, 320, 
    333, 328, 328, 313, 312, 317, _, _, _, _, 320, 332, 332, 343, 339, 333, 
    338, 320, _, _, _, 327, 322, 325, 323, 324, 323, 325, 331, 327, _, _, 
    309, 315, 312, 319, 308, 303, 293, 303, _, 294, 300, 295, 296, 302, 301, 
    315, 321, _, _, _, _, _, 296, 303, 294, 319, 324, 326, 335, 338, _, _, 
    328, 346, _, 327, 307, 334, 344, 10, _, _, _, 359, 336, 48, 16, 8, 55, 
    54, 55, _, _, 79, 75, 67, 85, 107, 127, 132, 183, 194, _, _, 183, 29, 
    216, 289, 283, 306, 308, 300, _, _, _, _, 334, 332, 324, 326, 330, 331, 
    329, 328, _, _, _, _, _, _, _, _, _, 15, 12, 17, 21, 22, 20, 20, 25, 13, 
    325, 311, 317, 331, 346, 339, 341, _, _, _, _, _, _, 320, 316, 310, 356, 
    327, 10, 319, 308, _, _, 325, 324, 318, 322, 322, 327, 6, 351, _, _, 321, 
    317, 317, 313, 317, 313, 319, 310, 322, 54, 52, 62, 73, 90, 106, _, 153, 
    156, 149, 139, 126, 120, _, _, _, _, _, _, 112, 117, 112, 121, 119, 117, 
    118, 112, _, _, _, _, _, 129, 121, 126, 123, 119, 124, 120, 122, _, _, _, 
    _, _, _, _, _, _, 124, 124, 121, 124, 127, 120, 124, 126, _, _, _, 111, 
    111, 110, 115, 114, 113, 113, 120, _, _, _, _, 118, 118, 117, 117, 117, 
    117, 118, 118, _, _, 118, 121, 124, 127, 128, 124, 123, 123, _, _, _, _, 
    112, 117, 122, 124, 122, 120, 120, _, _, _, 124, 125, 123, 120, 121, 121, 
    125, 125, _, _, _, 123, 122, 118, 116, 114, 109, 112, 113, _, _, 105, 
    100, 100, 100, 96, 96, 95, 94, _, _, _, 87, 85, 85, 85, 85, 86, 85, 89, 
    _, _, _, _, 87, 91, 84, 75, 77, 80, 87, 82, _, _, _, _, _, 76, 70, 72, 
    70, _, 77, 73, 76, 80, 84, 86, 79, 85, 85, 81, _, 83, 87, 102, 92, 80, 
    73, 74, _, _, _, _, _, _, _, _, 82, 85, 97, 93, 94, 91, 95, 91, 87, 75, 
    80, 85, 80, 85, 74, 80, 58, 52, 46, 40, 33, 20, 33, 45, 41, 43, 35, 26, 
    40, 32, 36, 34, 22, 25, 35, 45, 41, 34, 264, 243, 73, 99, 102, 100, 91, 
    111, 93, 101, 112, 117, 98, 107, 108, 124, 124, 118, 110, 115, 115, 113, 
    181, 186, 193, 210, 265, 273, 291, 311, 311, 331, 332, 325, 324, 339, 
    342, 344, 348, 22, 41, 14, 7, 11, 13, 15, 13, 41, 23, 38, 20, 16, 20, 8, 
    6, 15, 11, 14, 5, 5, 321, 330, 334, 338, 334, 327, 325, 318, 323, 342, 
    329, 334, 337, 331, 325, 327, 313, 321, 308, 320, 308, 327, 308, 312, 
    322, 319, 321, 331, 342, 341, 342, 343, 345, 344, 345, 340, 340, 339, 
    332, 339, 338, 345, 350, 346, 4, 4, 356, 2, 2, 356, 5, 9, 26, 55, 346, 
    343, 358, 47, 89, 85, 89, 97, 100, 106, 105, 111, 106, 102, 109, 114, 
    111, 111, 100, 90, 78, 78, 81, 75, 103, 100, 125, 73, 36, 331, 48, 22, 9, 
    350, 4, 1, 2, 16, 7, 335, 319, 317, 318, 317, 312, 316, 312, 313, 322, 
    316, 317, 320, 334, 314, 324, 325, 327, 342, 335, 334, 343, 350, 341, 4, 
    354, 346, 3, 18, 92, 84, 87, 95, 76, 71, 64, 86, 81, 71, 54, 59, 55, 54, 
    57, 55, 60, 62, 61, 53, 58, 55, 55, 57, 57, 55, 57, 57, 55, 53, 50, 43, 
    38, 37, 39, 37, 19, 4, 355, 348, 346, 346, 347, 348, 352, 345, 343, 341, 
    338, 343, 335, 324, 326, 326, 322, 322, 325, 320, 320, 328, 319, 336, 
    335, 323, 311, 308, 312, 312, 316, 333, 334, 334, 329, 318, 314, 312, 
    318, 314, 314, 312, 311, 304, 291, 307, 292, 286, 286, 292, 310, 312, 
    311, 309, 322, 315, 316, 315, 309, 309, 305, 305, 303, 307, 307, 311, 
    313, 310, 304, 302, 294, 319, 317, 305, 309, 306, 323, 315, 320, 325, 
    326, 319, 308, 302, 310, 306, 305, 294, 298, 302, 309, 307, 303, 297, 
    299, 298, 298, 307, 309, 306, 308, 320, 326, 296, 288, 295, 299, 309, 
    316, 313, 306, 305, 303, 334, 325, 318, 317, 324, 330, 320, 313, 302, 
    311, 317, 325, 315, 302, 306, 307, 312, 308, 304, 318, 320, 324, 321, 
    325, 324, 326, 330, 314, 284, 292, 310, 358, 90, 118, 129, 119, 115, 118, 
    112, 117, 118, 113, 116, 117, 111, 117, 134, 255, 296, 307, 309, 316, 
    300, 299, 296, 297, 295, 290, 292, 289, 284, 303, 304, 305, 320, 317, 
    315, 311, 308, 314, 324, 324, 287, 298, 296, 294, 302, 325, 326, 315, 
    331, 328, 332, 325, 316, 332, 18, 24, 78, 72, 96, 81, 112, 110, 105, 83, 
    70, 74, 76, 72, 66, 69, 66, 66, 62, 62, 62, 54, 55, 74, 80, 74, 79, 89, 
    84, 144, 121, 131, 140, 133, 119, 115, 247, 284, 302, 302, 325, 320, 316, 
    327, 322, 329, 334, 336, 329, 320, 320, 327, 322, 326, 325, 308, 307, 
    314, 318, 312, 315, 331, 304, 306, 324, 327, 297, 307, 298, 301, 278, 
    315, 326, 330, 335, 326, 330, 331, 328, 336, 325, 332, 325, 342, 337, 
    318, 329, 111, 111, 109, 117, 120, 119, 112, 102, 81, 89, 87, 88, 87, 86, 
    79, 87, 86, 85, 90, 85, 87, 85, 87, 91, 89, 92, 95, 96, 97, 100, 101, 
    106, 113, 118, 123, 120, 121, 121, 119, 130, 123, 122, 119, 118, 114, 
    115, 155, 49, 0, 298, 305, 329, 329, 340, 336, 352, 280, 125, 125, 112, 
    139, 208, 202, 126, 303, 207, 110, 118, 113, 115, 124, 113, 104, 143, 
    292, 302, 310, 321, 318, 316, 314, 316, 317, 303, 307, 310, 299, 301, 
    302, 305, 305, 304, 302, 302, 317, 318, 323, 325, 322, 317, 322, 338, 
    334, 339, 321, 310, 307, 308, 333, 323, 125, 334, 139, 107, 134, 117, 92, 
    109, 92, 86, 92, 94, 95, 110, 105, 109, 102, 110, 105, 110, 105, 105, 
    105, 109, 98, 92, 93, 102, 91, 94, 82, 78, 76, 93, 92, 91, 94, 93, 91, 
    95, 96, 104, 105, 107, 114, 118, 117, 112, 111, 115, 112, 111, 114, 112, 
    109, 112, 113, 115, 121, 134, 139, 294, 309, 317, 315, 310, 324, 325, 
    329, 334, 329, 329, 328, 327, 332, 330, 327, 330, 324, 316, 314, 316, 
    320, 313, 319, 304, 306, 304, 308, 316, 319, 315, 319, 328, 333, 344, 
    343, 324, 346, 341, 324, 315, 359, 7, 51, 87, 89, 95, 113, 121, 114, 123, 
    96, 113, 114, 111, 111, 112, 113, 113, 113, 116, 114, 115, 112, 114, 114, 
    118, 115, 116, 115, 112, 109, 101, 96, 96, 99, 106, 116, 116, 106, 113, 
    115, 120, 118, 115, 113, 112, 114, 114, 115, 110, 108, 111, 97, 97, 94, 
    98, 95, 84, 85, 89, 89, 85, 75, 81, 74, 73, 79, 75, 78, 79, 74, 70, 63, 
    60, 65, 67, 68, 67, 80, 66, 76, 67, 74, 67, 65, 58, 62, 63, 73, 80, 80, 
    72, 75, 77, 62, 77, 70, 59, 62, 58, 61, 51, 46, 42, 39, 40, 44, 44, 333, 
    37, 33, 24, 5, 348, 344, 314, 314, 312, 316, 313, 321, 316, 323, 324, 
    328, 315, 310, 318, 323, 331, 346, 335, 337, 350, 17, 334, 101, 57, 66, 
    83, 95, 0, 54, 108, 90, 94, 106, 107, 105, 107, 102, 63, 99, 90, 81, 79, 
    80, 69, 60, 57, 53, 54, 54, 56, 50, 61, 47, 43, 43, 45, 57, 61, 65, 65, 
    63, 67, 69, 67, 56, 58, 59, 58, 59, 61, 62, 61, 60, 62, 63, 65, 64, 54, 
    40, 45, 49, 49, 46, 54, 54, 50, 50, 52, 47, 44, 44, 46, 43, 50, 44, 28, 
    41, 20, 15, 360, 355, 3, 1, 349, 4, 350, 335, 331, 334, 322, 315, 297, 
    288, 286, 278, 264, 237, 239, 235, 200, 110, 102, 105, 115, 118, 124, 94, 
    122, 105, 107, 103, 102, 101, 96, 90, 96, 91, 93, 95, 94, 102, 106, 81, 
    75, 72, 75, 83, 85, 77, 60, 64, 62, 59, 61, 59, 59, 64, 56, 49, 56, 56, 
    55, 47, 55, 51, 55, 52, 47, 53, 50, 46, 48, 46, 40, 37, 39, 43, 41, 46, 
    51, 54, 54, 57, 60, 57, 59, 57, 64, 66, 69, 67, 64, 68, 90, 99, 104, 85, 
    110, 95, 101, 119, 118, 132, 125, 132, 148, 125, 114, 112, 116, 119, 121, 
    122, 118, 121, 118, 118, 120, 118, 121, 118, 111, 119, 117, 115, 118, 
    122, 122, 124, 125, 119, 114, 110, 102, 111, 103, 130, 121, 119, 116, 
    106, 100, 104, 118, 101, 97, 91, 85, 75, 68, 69, 57, 52, 58, 78, 74, 92, 
    79, 82, 84, 92, 86, 87, 85, 85, 77, 79, 78, 77, 75, 79, 83, 77, 77, 73, 
    70, 68, 66, 61, 55, 57, 59, 55, 61, 61, 83, 97, 114, 94, 91, 112, 120, 
    100, 89, 90, 104, 108, 99, 84, 91, 129, 119, 115, 130, 119, 119, 114, 
    114, 130, 140, 184, 170, 156, 168, 168, 167, 167, 166, 225, 218, 226, 
    247, 125, 172, 192, 190, 240, 264, 270, 278, 298, 321, 356, 331, 318, 
    333, 360, 12, 341, 118, 101, 132, 277, 96, 298, 63, 129, 116, 93, 91, 76, 
    89, 126, 4, 2, 360, 319, 11, 276, 330, 336, 5, 319, 316, 317, 315, 322, 
    317, 315, 305, 316, 296, 316, 315, 329, 327, 310, 320, 317, 319, 320, 
    327, 323, 322, 320, 323, 325, 323, 322, 320, 320, 324, 319, 324, 327, 
    320, 317, 318, 317, 323, 317, 324, 317, 315, 327, 334, 329, 322, 329, 
    328, 320, 331, 330, 322, 316, 316, 323, 333, 322, 324, 331, 317, 330, 
    338, 330, 322, 333, 309, 312, 323, 329, 321, 333, 331, 323, 330, 329, 
    325, 319, 325, 324, 323, 311, 322, 328, 311, 312, 313, 318, 313, 315, 
    322, 320, 338, 337, 325, 350, 321, 323, 346, 346, 314, 316, 318, 322, 
    347, 342, 348, 351, 359, 350, 323, 328, 322, 335, 324, 326, 321, 316, 
    321, 330, 321, 327, 335, 348, 338, 329, 327, 325, 333, 336, 303, 326, 
    329, 336, 330, 329, 325, 325, 295, 331, 304, 309, 312, 310, 308, 306, 
    316, 318, 312, 313, 306, 322, 328, 318, 310, 305, 304, 315, 317, 330, 
    342, 332, 323, 311, 311, 311, 310, 304, 309, 342, 318, 295, 316, 330, 
    318, 309, 309, 319, 318, 330, 337, 320, 315, 300, 299, 302, 304, 307, 
    304, 318, 307, 303, 294, 296, 299, 310, 311, 308, 319, 311, 306, 310, 
    331, 329, 336, 316, 323, 348, 307, 332, 311, 287, 285, 319, 334, 329, 84, 
    85, 86, 69, 79, 84, 94, 120, 69, 69, 73, 73, 72, 71, 67, 61, 62, 56, 64, 
    64, 66, 63, 61, 47, 56, 56, 60, 56, 58, 57, 55, 55, 53, 51, 50, 51, 51, 
    51, 49, 50, 49, 50, 49, 51, 51, 52, 51, 52, 51, 48, 48, 48, 51, 61, 64, 
    62, 66, 57, 55, 57, 62, 53, 60, 65, 70, 68, 61, 66, 74, 79, 81, 81, 89, 
    81, 81, 80, 71, 70, 69, 68, 71, 74, 73, 81, 81, 76, 80, 84, 82, 83, 88, 
    92, 94, 94, 99, 98, 93, 94, 90, 92, 87, 85, 84, 83, 79, 82, 82, 86, 83, 
    82, 87, 88, 87, 91, 89, 87, 83, 80, 93, 101, 104, 102, 98, 98, 91, 88, 
    91, 88, 88, 86, 87, 89, 92, 93, 93, 92, 91, 90, 92, 92, 94, 98, 99, 103, 
    100, 101, 100, 95, 97, 93, 92, 91, 90, 94, 95, 92, 89, 74, 70, 64, 56, 
    57, 71, 65, 62, 64, 62, 64, 67, 63, 59, 56, 65, 65, 67, 84, 76, 82, 77, 
    77, 94, 116, 108, 103, 107, 116, 120, 118, 120, 118, 108, 127, 120, 352, 
    316, 299, 294, 289, 315, 316, 292, 305, 322, 325, 325, 320, 317, 314, 
    310, 303, 314, 356, 9, 8, 118, 95, 104, 104, 90, 93, 91, 78, 85, 75, 78, 
    82, 86, 72, 77, 83, 87, 98, 104, 103, 108, 113, 112, 111, 117, 120, 120, 
    113, 117, 115, 118, 119, 119, 118, 118, 117, 109, 108, 107, 109, 110, 
    113, 113, 117, 123, 135, 160, 170, 174, 98, 113, 122, 133, 72, 346, 281, 
    138, 304, 340, 93, 102, 103, 120, 119, 121, 117, 115, 111, 119, 119, 127, 
    113, 111, 110, 112, 120, 115, 115, 126, 124, 123, 121, 115, 118, 116, 
    116, 115, 113, 113, 137, 128, 123, 102, 119, 103, 89, 118, 64, 48, 48, 
    51, 56, 54, 52, 52, 52, 51, 54, 55, 55, 66, 54, 59, 59, 62, 63, 64, 64, 
    70, 69, 77, 81, 93, 119, 103, 109, 115, 115, 116, 117, 117, 119, 128, 
    127, 120, 119, 116, 114, 120, 111, 112, 89, 128, 78, 333, 294, 119, 107, 
    11, 317, 315, 316, 311, 310, 342, 1, 344, 87, 314, 51, 340, 55, 52, 36, 
    42, 48, 50, 41, 53, 203, 54, 66, 54, 51, 52, 56, 58, 66, 53, 56, 161, 4, 
    138, 134, 57, 8, 323, 62, 63, 62, 61, 56, 60, 59, 56, 53, 56, 57, 55, 52, 
    355, 356, 46, 104, 29, 55, 55, 28, 67, 62, 297, 321, 358, 303, 301, 199, 
    317, 320, 8, 0, 131, 66, 320, 330, 354, 1, 360, 21, 127, 118, 46, 39, 47, 
    39, 307, 8, 8, 32, 27, 25, 21, 45, 25, 19, 25, 228, 306, 357, 4, 11, 28, 
    24, 331, 102, 18, 310, 28, 19, 358, 348, 348, 346, 350, 358, 352, 346, 
    348, 2, 350, 355, 2, 5, 8, 359, 2, 347, 14, 337, 305, 15, 93, 124, 135, 
    119, 105, 143, 137, 139, 138, 131, 112, 115, 131, 138, 124, 111, 271, 
    277, 330, 305, 352, 6, 17, 353, 350, 359, 1, 326, 317, 335, 351, 110, 99, 
    96, 103, 102, 116, 113, 109, 106, 105, 105, 98, 97, 95, 85, 72, 70, 74, 
    73, 74, 68, 52, 44, 29, 303, 314, 91, 36, 11, 55, 36, 52, 52, 55, 48, 51, 
    49, 359, 96, 10, 50, 281, 41, 89, 82, 88, 91, 100, 107, 96, 106, 107, 
    115, 110, 114, 107, 111, 106, 107, 113, 110, 109, 112, 110, 117, 109, 
    116, 118, 109, 117, 121, 120, 112, 112, 117, 130, 128, 123, 136, 153, 
    104, 105, 185, 188, 184, 122, 112, 108, 122, 165, 164, 170, 185, 184, 
    186, 188, 184, 170, 167, 181, 160, 127, 120, 137, 126, 97, 43, 119, 112, 
    299, 320, 255, 325, 332, 87, 53, 60, 56, 45, 54, 50, 48, 41, 47, 49, 46, 
    43, 31, 48, 305, 95, 22, 248, 0, 27, 16, 32, 31, 4, 233, 19, 42, 22, 50, 
    30, 23, 42, 7, 3, 358, 111, 73, 50, 21, 50, 51, 52, 53, 51, 52, 54, 50, 
    49, 43, 47, 47, 49, 49, 49, 46, 54, 50, 44, 50, 44, 48, 45, 160, 134, 
    360, 338, 242, 288, 332, 335, 340, 8, 266, 4, 2, 360, 48, 43, 26, 66, 74, 
    129, 18, 20, 35, 30, 29, 42, 24, 246, 260, 360, 26, 339, 9, 360, 333, 
    300, 266, 12, 321, 5, 7, 8, 328, 343, 344, 317, 323, 322, 326, 326, 329, 
    320, 297, 16, 17, 17, 51, 27, 111, 43, 15, 41, 50, 46, 51, 60, 66, 65, 
    66, 66, 73, 77, 74, 90, 67, 82, 74, 96, 100, 114, 128, 138, 128, 113, 
    110, 111, 119, 109, 115, 107, 107, 99, 104, 97, 113, 113, 105, 109, 100, 
    105, 110, 115, 120, 123, 110, 109, 119, 91, 129, 62, 39, 12, 64, 92, 73, 
    49, 11, 33, 25, 26, 65, 31, 55, 316, 155, 69, 133, 115, 58, 61, 59, 54, 
    56, 64, 56, 61, 59, 77, 72, 72, 64, 67, 58, 57, 53, 53, 55, 33, 50, 56, 
    55, 55, 49, 53, 60, 53, 53, 54, 55, 56, 55, 53, 56, 54, 54, 54, 55, 49, 
    52, 55, 52, 50, 51, 53, 62, 64, 66, 72, 70, 71, 69, 72, 77, _, _, 87, 91, 
    92, 105, 93, 88, 86, 99, 106, 106, 114, 117, 114, 115, 116, 111, 124, 
    137, 139, 142, 148, 148, 148, 150, 144, 142, 137, 128, 122, 124, 124, 
    121, 129, 134, 140, 143, 145, 145, 146, 144, 145, 144, 139, 139, 137, 
    133, 128, 127, 125, 128, 130, 126, 128, 128, 126, 126, 131, 136, 147, 
    143, 140, 139, 132, 124, 116, 300, 307, 305, 324, 319, 308, 304, 305, 
    306, 317, 309, 313, 317, _, 321, 323, _, _, 318, _, 309, 308, 309, _, 
    307, _, 308, 307, 310, 305, 306, _, 295, 297, 324, 334, 329, 321, 7, 19, 
    14, 356, 302, 7, _, 333, _, 328, 329, 324, 328, 324, 316, 320, 327, 327, 
    327, 326, 323, 328, 322, 322, 322, 320, 320, 319, 321, 321, 317, 317, 
    319, 311, 307, 308, 307, 319, 305, 305, 304, 307, 314, 316, 310, 314, 
    324, 320, 319, 320, 316, 318, 332, 332, 333, 324, 323, 330, 329, 324, 
    323, 334, 337, 332, 344, 330, 341, 324, 353, 339, 324, 331, 7, 353, 347, 
    9, 8, 9, 6, 14, 20, 14, 6, 6, 9, 14, 25, 25, 32, 10, 14, 15, 19, 10, 9, 
    20, 37, 45, 36, 12, 10, 14, 1, 327, 13, 5, 1, 2, 11, 9, 2, 359, 349, 348, 
    351, 352, 359, 358, 354, 348, 299, 350, 6, 36, 3, 70, 78, 21, 21, 19, 
    345, 317, 358, 331, 17, 51, 342, 347, 358, 310, 307, 355, 324, 301, 319, 
    326, 347, 342, 350, 333, 335, 333, 333, 344, 334, 337, 324, 324, 328, 
    331, 331, 332, 321, 331, 334, 348, 5, 3, 342, 328, 332, 320, 89, 60, 328, 
    327, 328, 341, 338, 347, 357, 3, 6, 3, 360, 30, 91, 97, 102, 94, 105, 
    105, 105, 106, 93, 89, 81, 77, 81, 82, 81, 82, 79, 80, 74, 71, 69, 65, 
    63, 66, 73, 97, 119, 112, 114, 103, 118, 120, 120, 151, 157, 119, 104, 
    130, 131, 143, 88, 160, 169, 118, 164, 149, 103, 116, 110, 100, 118, 115, 
    114, 70, 71, 71, 184, 17, 36, 325, 320, 113, 318, 346, 313, 309, 312, 
    319, 317, 315, 312, 305, 308, 319, 317, 303, 303, 310, 313, 318, 320, 
    317, 316, 306, 316, 314, 313, 292, 310, 308, 310, 312, 309, 308, 293, 
    296, 296, 297, 300, 294, 291, 285, 255, 254, 258, 256, 255, 256, 252, 
    278, 292, 307, 310, 327, 300, 302, 298, 303, 309, 311, 307, 306, 319, 
    303, 326, 307, 310, 313, 317, 309, 309, 282, 285, 279, 305, 279, 350, 
    291, 254, 259, 254, 249, 250, 221, 228, 215, 200, 199, 206, 184, 115, 43, 
    101, 105, 181, 216, 149, 32, 52, 75, 71, 62, 25, 14, 41, 43, 15, 22, 329, 
    334, 332, 319, 315, 313, 310, 309, 310, 314, 326, 299, 276, 324, 328, 
    257, 253, 275, 231, 251, 265, 21, 13, 12, 15, 33, 13, 17, 8, 15, 12, 8, 
    354, 4, 12, 15, 18, 16, 13, 12, 13, 18, 16, 23, 9, 85, 321, 23, 25, 315, 
    134, 351, 35, 2, 334, 84, 68, 343, 48, 356, 341, 14, 58, 54, 53, 54, 54, 
    54, 54, 61, 61, 56, 57, 53, 47, 55, 53, 55, 53, 55, 55, 58, 54, 54, 51, 
    51, 50, 50, 51, 22, 257, 311, 301, 315, 359, 2, 8, 355, 330, 306, 307, 
    306, 284, 293, 295, 303, 305, 294, 303, 303, 295, 294, 292, 301, 305, 
    314, 313, 317, 297, 296, 295, 308, 314, 306, 328, 303, 330, 327, 350, 
    344, 10, 312, 337, 97, 327, 321, 325, 90, 89, 126, 40, 1, 75, 340, 7, 46, 
    327, 351, 328, 314, 33, 50, 8, 322, 20, 334, 44, 55, 64, 65, 82, 46, 43, 
    48, 120, 78, 79, 69, 60, 55, 54, 53, 54, 56, 50, 56, 63, 70, 64, 55, 55, 
    53, 54, 55, 57, 58, 55, 56, 56, 57, 57, 60, 57, 61, 61, 63, 70, 69, 71, 
    65, 73, 68, 66, 66, 68, 64, 76, 67, 70, 70, 70, 70, 72, 71, 76, 78, 79, 
    80, 81, 77, 79, 85, 89, 95, 96, 99, 103, 100, 102, 104, 104, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 124, 114, 124, 117, 116, 117, 109, 109, 
    106, 103, 106, 110, 124, 149, 163, 182, 180, 188, 186, 184, 193, 191, 
    175, 177, 168, 154, 159, 174, 238, 289, 305, 269, 273, 266, 265, 260, 
    266, 269, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 337, 347, 323, 348, 353, 351, 342, 345, 
    347, 340, 331, 329, 334, 331, 314, 309, 318, 329, 325, 328, 339, 320, 
    338, 349, 341, 336, 347, 348, 359, 354, 350, 351, 342, 341, 326, 346, 
    336, 325, 334, 334, 336, 338, 335, 338, 332, 319, 319, 311, 311, 312, 
    313, 310, 312, 315, 318, 318, 324, 325, 325, 322, 319, 316, 311, 309, 
    310, 318, 314, 314, 307, 309, 306, 309, 307, 322, 317, 316, 315, 313, 
    311, 312, 314, 314, 314, 313, 321, 318, 333, 352, 344, 352, 353, 346, 
    357, 358, 336, 340, 333, 313, 315, 323, 316, 317, 321, 324, 334, 330, 69, 
    74, _, 63, _, _, 64, 66, 354, 56, 288, 358, _, 345, 356, _, 7, 332, _, 
    351, 1, _, _, _, _, 0, 355, _, 352, _, 335, 331, 330, 346, 328, 336, 335, 
    337, 339, 339, 330, 331, 319, 318, 323, 322, 327, 317, 315, 305, 312, 
    308, 315, 310, 319, 319, 315, 323, 315, 316, 320, 314, 318, 311, 318, 
    326, 332, 336, 345, 348, 328, 308, 325, 322, 318, 320, 322, 332, 144, 
    103, 102, 128, 124, 135, 135, 142, 144, 140, 135, 131, 130, 127, 119, 
    117, 116, 111, 109, 110, 122, 115, 112, 140, 173, 143, 118, 123, 106, 
    114, 127, 119, 126, 114, 141, 198, 199, 95, 254, 107, 108, 120, 107, 145, 
    125, 120, 105, 123, 115, 107, 116, _, _, _, 124, 149, 119, 105, 114, 114, 
    123, 123, 108, 100, 90, 94, 59, 57, 57, 65, 66, 72, 72, 77, 79, 59, 54, 
    55, 53, 49, 51, 51, 51, 50, 48, 49, 51, 51, 318, 297, 284, 30, 44, 326, 
    342, 76, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 47, 50, 51, 49, 54, 54, 57, 59, _, 55, 54, 52, 52, 57, _, 
    _, 55, 52, 53, 51, 50, 49, 49, 47, _, 47, 41, 43, 45, _, 44, 31, 31, 18, 
    2, 0, 359, 336, 354, 338, 330, 324, 333, 348, 342, 331, 339, 335, 333, 
    328, 330, 330, 328, 329, 323, 323, 324, 327, 323, 325, 319, 319, 317, 
    319, 312, 313, 311, 309, 309, 303, 296, 297, 297, 306, 307, 308, 309, 
    302, 298, 300, 297, 300, 295, 298, 305, 305, 297, 304, 307, 301, 301, 
    301, 303, 305, 320, 315, _, 326, 323, 327, 331, 325, 324, 324, 332, 336, 
    334, 332, 323, 329, 326, 325, 322, 313, 319, 314, 327, 324, 330, 343, 3, 
    110, 119, 129, 140, 100, 103, 109, 115, 111, 108, 105, 100, 100, 102, 90, 
    105, 97, 80, 95, 82, 94, 91, 89, 85, 78, 83, 85, 97, 100, 89, 74, 74, 67, 
    62, 71, 70, 80, 57, 46, 53, 54, 69, 76, 57, 54, 50, 59, 61, 62, 64, 74, 
    71, 82, 81, 90, 94, 101, 97, 84, 89, 81, 92, 97, 89, _, 93, 96, 106, 101, 
    98, 98, 53, 76, 62, 58, 56, 49, 53, 55, 58, 55, 58, 57, 46, 50, 43, 43, 
    43, 23, 129, 6, 315, 352, 326, 342, 323, 324, 326, 346, 334, 322, 309, 
    305, 306, 304, 312, 311, 317, 314, 316, 343, 339, 342, 333, 335, 5, 354, 
    316, 33, 32, 23, 13, 20, 346, 328, 334, 46, 52, 65, 60, 81, 87, 71, 68, 
    65, 63, 71, 75, 72, 66, 65, 64, 61, 55, 45, 43, 29, 57, 305, 84, 323, 
    349, 10, 318, 0, 355, 355, 321, 339, 339, 328, 325, 322, 320, 320, 323, 
    307, 307, 302, 310, 318, 312, 309, 306, 308, 317, 310, 310, 313, 304, 
    305, 296, 289, 293, 303, 304, 317, 321, 327, 323, 317, 308, 295, 327, 
    333, 335, 347, 354, 358, 0, 52, 30, 58, 66, 92, 94, 74, 116, 127, 130, 
    122, 143, 138, 125, 138, 131, 132, 129, 105, 98, 102, 97, 101, 99, 98, 
    95, 96, 100, 98, 89, 86, 88, 89, 96, 99, 110, 114, 119, 117, 122, 116, 
    128, 153, 132, 134, 121, 114, 114, 109, 111, 104, 123, 132, 124, 100, 89, 
    86, 81, 111, 118, 114, 114, 116, 130, 129, 125, 126, 125, 126, 127, 129, 
    130, 127, 126, 126, 122, 122, 124, 123, 123, 125, 136, 140, 143, 156, 
    271, 306, 289, 307, 306, 319, 261, 153, 147, 185, 221, 276, 291, 357, 
    323, 99, 75, 74, 85, 96, 120, 123, 100, 95, 88, 93, 90, 101, 113, 113, 
    96, 84, 63, 46, 328, 353, 322, 327, 328, 329, 329, 334, 317, 318, 329, 
    311, 322, 321, 311, 315, 309, 314, 308, 308, 307, 306, 303, 299, 320, 
    341, 357, 2, 10, 15, 228, 221, 218, 214, 198, 195, 216, 219, 343, 336, 
    342, 345, 333, 343, 283, 310, 307, 306, 338, 326, 296, 312, 304, 316, 
    293, 300, 290, 250, 244, 255, 215, 206, 200, 196, 195, 178, 118, 107, 
    113, 132, 126, 129, 127, 129, 117, 111, 122, 122, 32, 15, 18, 4, 14, 13, 
    359, 186, 287, 54, 63, 52, 61, 58, 58, 63, 59, 64, 67, 68, 67, 62, 66, 
    65, 48, 64, 45, 67, 79, 350, 279, 314, 7, 324, 346, 335, 335, 327, 331, 
    326, 330, 332, 330, 324, 328, 333, 329, 319, 310, 306, 317, 316, 314, 
    295, 298, 301, 296, 308, 301, 301, 299, 304, 308, 304, 310, 316, 318, 
    316, 320, 331, 332, 326, 320, 334, 332, 330, 333, 330, 330, 332, 334, 
    337, 342, 338, 335, 336, 347, 346, 341, 333, 341, 325, 339, 339, 330, 
    342, 344, 328, 335, 334, 332, 336, 330, 332, 340, 341, 324, 334, 334, 
    333, 334, 326, 328, 324, 333, 336, 331, 332, 337, 319, 318, 320, 317, 
    329, 337, 325, 331, 341, 335, 335, 335, 329, 5, 319, 328, 321, 322, 337, 
    325, 323, 294, 32, 357, 31, 30, 27, 32, 12, 14, 351, 334, 13, 24, 17, 
    327, 319, 22, 330, 329, 347, 325, 304, 332, 359, 53, 354, 80, 83, 97, 
    116, 85, 103, 100, 89, 123, 69, 55, 41, 304, 85, 110, 320, 59, 101, 100, 
    100, 86, 60, 346, 344, 317, 55, 59, 49, 51, 19, 333, 2, 323, 328, 89, 
    305, 323, 324, 305, 307, 311, 275, 276, 281, 297, 312, 306, 312, 320, 
    321, 311, 313, 302, 242, 233, 234, 273, 273, 296, 281, 322, 318, 327, 
    340, 67, 83, 118, 112, 97, 103, 104, 101, 80, 89, 66, 75, 70, 75, 71, 72, 
    64, 63, 65, 64, 62, 64, 59, 64, 62, 74, 77, 69, 31, 32, 68, 64, 56, 51, 
    54, 46, 39, 35, 30, 17, 5, 8, 3, 3, 351, 349, 348, 351, 350, 349, 343, 
    345, 345, 341, 343, 343, 346, 336, 330, 329, 328, 330, 332, 333, 334, 
    336, 338, 340, 343, 348, 1, 9, 10, 306, 334, 339, 353, 14, 27, 221, 318, 
    314, 306, 49, 23, 14, 10, 14, 321, 328, 326, 41, 303, 334, 326, 311, 114, 
    108, 112, 94, 105, 114, 91, 88, 84, 83, 78, 72, 74, 89, 62, 56, 53, 277, 
    357, 156, 87, 81, 71, 59, 54, 39, 331, 323, 29, 351, 353, 352, 19, 340, 
    350, 341, 348, 354, 333, 344, 346, 2, 349, 11, 25, 25, 26, 341, 16, 302, 
    291, 266, 31, 15, 351, 2, 2, 335, 5, 350, 5, 3, 0, 354, 349, 356, 7, 29, 
    18, 14, 29, 21, 17, 17, 13, 2, 2, 7, 356, 356, 10, 356, 5, 10, 353, 356, 
    17, 25, 19, 6, 19, 24, 1, 3, 356, 1, 7, 1, 1, 343, 323, 338, 358, 14, 15, 
    322, 14, 149, 287, 11, 322, 349, 115, 132, 169, 161, 142, 145, 143, 136, 
    139, 137, 127, 137, 119, 122, 133, 123, 116, 114, 129, 131, 119, 120, 
    130, 115, 121, 128, 127, 115, 118, 147, 132, 124, 122, 135, 123, 121, 
    129, 115, 135, 109, 108, 116, 111, 113, 120, 130, 116, 118, 107, 101, 
    109, 110, 125, 113, 121, 345, 285, 284, 289, 277, 307, 310, 315, 325, 
    319, 313, 298, 322, 314, 306, 301, 308, 317, 343, 328, 329, 318, 340, 
    300, 337, 326, 328, 327, 326, 324, 340, 341, 316, 2, 109, 132, 137, 137, 
    138, 127, 126, 111, 95, 84, 89, 88, 92, 100, 106, 106, 114, 117, 120, 
    129, 138, 123, 126, 122, 124, 132, 126, 124, 117, 109, 93, 101, 112, 112, 
    113, 111, 112, 108, 119, 110, 119, 116, 131, 133, 131, 122, 117, 109, 95, 
    91, 80, 68, 41, 41, 318, 35, 49, 279, 155, 42, 50, 3, 58, 40, 53, 58, 56, 
    59, 76, 56, 53, 54, 48, 22, 324, 266, 254, 263, 326, 47, 52, 38, 54, 69, 
    60, 66, 57, 63, 58, 46, 51, 45, 340, 29, 247, 357, 323, 293, 289, 270, 
    282, 282, 286, 308, 320, 325, 311, 310, 302, 296, 294, 300, 296, 298, 
    300, 304, 301, 301, 300, 301, 303, 294, 301, 301, 302, 297, 296, 291, 
    298, 310, 314, 301, 309, 335, 320, 315, 317, 320, 315, 318, 335, 327, 
    334, 353, 338, 322, 321, 357, 355, 345, 331, 17, 344, 347, 352, 321, 312, 
    314, 316, 321, 307, 322, 309, 311, 320, 315, 312, 298, 305, 309, 314, 
    320, 355, 319, 305, 302, 300, 294, 299, 301, 306, 321, 330, 356, 321, 
    305, 337, 349, 334, 340, 337, 326, 319, 323, 321, 333, 330, 335, 307, 
    318, 350, 353, 22, 0, 347, 335, 330, 324, 324, _, 311, _, _, _, 327, 328, 
    321, 327, 324, 322, 322, 320, 273, 255, 295, 57, 55, 49, 63, 328, 49, 
    111, 124, 109, 115, 124, 100, 105, 120, 104, 101, _, 107, 118, 105, 110, 
    _, 55, _, _, 65, 64, 65, 63, 77, 60, 57, 78, 50, 63, _, 62, 51, 306, 5, 
    _, 322, 347, 310, 304, _, 13, 357, 23, _, _, 14, _, 4, 358, 2, 351, 336, 
    333, 329, 329, 331, 328, 327, 321, 323, _, 311, _, 311, 314, 314, 317, _, 
    307, _, 306, 305, 308, 307, 303, _, 299, 293, 287, 294, 295, 297, 297, 
    297, 300, 300, 286, 284, 283, 289, 297, 303, 313, 318, 328, 331, 338, 
    321, 344, 19, 325, 331, 336, 342, 354, 346, 348, 2, 2, 358, 357, 360, 
    358, 351, 349, _, _, 356, 344, _, 357, 338, 327, 331, 329, 324, 324, 329, 
    343, 353, 358, 355, 348, 345, 339, 345, 343, 340, 342, 343, 336, 343, 
    337, 340, 340, 331, 346, 331, 322, 327, 333, 322, 328, 321, 327, 326, 
    330, 323, 337, 319, 314, 11, 348, 332, 329, 316, 320, 324, 326, 322, 324, 
    323, 318, 309, 304, 303, 311, 314, 314, 308, 303, 303, 309, 326, 330, 
    322, 319, _, 318, 311, 313, 315, 321, 322, 323, 318, 318, 313, 307, 311, 
    311, 319, 319, 310, 325, 323, 319, 313, 312, 318, _, 306, 308, 303, 289, 
    302, 298, 292, 281, 260, 262, 299, 296, 304, 290, 279, 281, 291, 296, 
    306, 285, 291, 284, 279, 289, 272, 278, 266, 286, 291, 299, 219, 86, 127, 
    139, 138, 59, 108, 126, 133, 122, 115, 124, 118, 115, 114, 113, 116, 119, 
    120, 128, 127, 124, 114, 117, 120, 136, 127, 123, 124, 122, 136, 132, 
    136, 143, 137, 136, 131, 126, 123, 123, 114, _, 114, 113, 108, 105, 108, 
    105, 105, 98, 91, 87, 85, 89, 86, 87, 79, 89, 85, 64, 60, 43, 35, 52, 96, 
    57, 36, 302, 310, 349, 279, 287, 310, 307, 58, 39, 14, 18, 351, 9, 4, 
    353, 341, 343, 340, 344, 334, 336, 334, 341, 350, _, 9, 12, 4, 1, 1, 10, 
    6, 2, 358, 354, 355, 3, 4, 4, 6, 7, 7, 4, 15, 16, 18, 36, 41, 51, 52, 46, 
    47, 49, 57, 57, 61, 54, 52, 41, 31, 35, 39, 32, 39, 39, 43, 50, 51, 55, 
    61, 58, 58, 55, 50, 55, 58, 58, 73, 259, 75, 158, 27, 77, 88, 77, 73, 80, 
    79, 74, 72, 77, 86, 84, 82, 80, 75, _, 303, 276, 55, 78, 71, 91, 84, 88, 
    81, 51, 271, 187, 336, 301, 107, 343, 359, 339, 338, 352, 318, 324, 352, 
    16, 349, 317, 322, 346, 325, 336, 343, 337, 342, 316, 315, 342, 316, 315, 
    321, 321, 315, 311, 319, 321, 328, 327, 324, 329, 325, 325, 329, 322, 
    325, 325, 329, 329, 328, 335, 337, 332, 328, 332, 326, 319, 326, 325, 
    322, 327, 325, 318, 318, _, 312, 321, 325, 322, 325, 327, 327, 318, 318, 
    312, 308, 315, 321, 324, 322, 320, 310, 310, 314, 312, 314, 321, 318, 
    316, 317, 312, 325, 321, 326, 326, 326, 323, 324, 323, 329, 327, 347, 
    339, 339, 337, 336, 318, 310, 324, 309, 321, 324, 324, 326, 322, 322, 
    323, 324, 323, 349, 322, 329, 318, 324, 340, 39, 151, 169, 226, 239, 285, 
    0, 335, 148, 130, 144, 156, 294, 331, 290, 145, 331, 186, 274, 323, 294, 
    318, 326, 323, 312, 303, 310, 311, 322, 304, 301, 280, 238, 280, 269, 
    244, 245, 266, 189, 323, 339, 325, 160, 234, 184, 177, 207, 246, 255, 
    242, 306, 282, 277, 310, 265, 313, 298, 283, 299, 292, 267, 173, 319, 
    301, 305, 316, 319, 303, 314, 299, 290, 284, 1, 159, 194, 229, 257, 136, 
    163, 162, 156, 154, 181, 175, _, 159, 140, 111, 110, 132, 140, 130, 110, 
    119, 146, 138, 134, 122, 114, 111, 132, 129, 116, 126, 130, 121, 105, 71, 
    72, 110, 260, 53, 55, 299, 40, 205, 242, 291, 317, 326, 300, 307, 294, 
    314, 286, 304, 316, 327, 83, 30, 99, 293, 284, 281, 54, 54, 57, 50, 50, 
    257, 210, 88, 99, 46, 45, 282, 354, 321, 333, 326, 311, 324, 326, 347, 
    332, 326, _, 339, 342, 346, 354, 327, 331, 326, 329, 320, 322, 320, 323, 
    326, 318, 325, 316, 284, 235, 296, 256, 209, 67, 64, 65, 228, 271, 335, 
    197, 15, 352, 50, 59, 57, 56, 24, 110, 243, 125, 30, 32, 325, 337, 343, 
    321, 310, 319, _, 315, 307, 314, 319, 315, 326, 324, 321, 334, 331, 320, 
    316, 324, 315, 315, 330, 321, 323, 311, 289, 288, 293, 305, 308, 308, 
    309, _, 314, 317, 309, 307, 318, 326, 326, 329, 329, 335, 344, 334, 5, 
    326, 325, 326, 325, 335, 327, 302, 299, 309, _, 320, 320, 321, 322, 322, 
    300, 301, 312, 296, 271, 273, 354, 332, 317, 315, 324, 317, 256, 205, 
    194, 148, 183, 223, 283, 260, 15, 257, 297, 163, 116, 107, 120, 126, 122, 
    143, 87, 351, 252, 354, 296, 272, 176, 140, _, 136, 118, 108, 143, 159, 
    112, 217, 292, 309, 310, 318, 318, 316, 321, 323, 355, 342, 349, 329, 
    328, 322, 324, 333, 315, 322, 320, 322, 322, 318, 317, 317, 311, 308, 
    319, 329, 330, 329, 324, 325, 328, 327, 329, 327, 327, 321, 320, 319, 
    327, 317, 315, 317, 316, 318, 322, 309, 319, 332, 321, 316, 318, 321, 
    349, 318, 305, 331, 312, 311, 328, 323, 314, 360, _, 297, 303, 318, 324, 
    328, 330, 322, 318, 319, 320, 320, 321, 317, 318, 315, 315, 312, 318, 
    315, 302, 316, 320, 319, 309, 308, 307, 320, 319, 320, 324, 319, 326, 
    323, 319, 326, 329, 331, 327, 328, 329, 329, 331, 319, 313, 327, 319, 
    327, 314, 359, 320, 301, 7, 285, _, 330, 272, 318, 333, 324, 323, _, 60, 
    353, 317, 255, 342, 320, 336, 321, _, _, _, 19, _, 335, 323, 335, 320, 
    322, 321, _, _, 322, _, 312, 317, 317, 318, 327, _, 331, _, 327, _, _, 
    313, 316, 307, 323, _, 325, _, 325, 339, 331, _, 311, 325, 329, _, 331, 
    330, 333, _, 323, 333, _, 309, 314, 320, 327, 330, 311, 316, 318, 316, 
    314, _, _, _, _, 302, 299, _, 312, 317, 324, 318, 314, 318, 322, 313, 
    303, 311, 304, 313, 311, _, _, 318, _, 320, 318, 312, 315, 329, 325, 313, 
    324, 318, 313, 298, 288, 308, 302, 314, 301, 320, 314, 317, 309, 319, 
    321, 310, 317, 319, 319, 320, 312, 324, 333, 324, 323, 305, 306, 313, 
    306, 302, 308, 316, 294, 313, _, 310, 320, 319, 317, 321, _, 316, 312, _, 
    324, 318, 314, 319, 325, 305, _, 312, 316, 305, 304, 312, 316, 307, 306, 
    308, 304, 299, 305, 306, 304, 306, 314, 317, 317, 326, 320, 325, 319, 
    317, 313, 306, 301, 294, 290, 298, 307, 326, 324, 330, 335, 332, 340, 
    343, 360, 354, 2, 345, 329, 327, 334, 324, 324, 327, 322, 8, 21, 30, 8, 
    355, 326, 322, 299, 310, 297, 323, 312, 277, 288, 279, 312, 42, 291, 343, 
    _, 333, 335, 322, 319, 344, 360, 345, 334, 357, 27, 29, 211, 342, 341, 
    340, 328, 331, 329, 325, 324, 317, 324, 333, 341, 9, 12, 12, 351, 16, 14, 
    9, 308, 26, 330, 256, 231, 321, 333, 298, 357, 37, 33, 40, 239, 283, 308, 
    49, 55, 49, 11, 245, 344, 273, 328, 305, 328, 326, 324, 327, 328, 325, 
    323, 282, 274, 72, 38, 40, 251, 323, 320, 306, 320, 22, 17, 14, 9, 285, 
    348, 305, 346, 309, 332, 213, 119, 55, 322, 311, 301, 315, 309, 318, 328, 
    311, 310, 316, 314, 301, 321, 318, 324, 319, 317, 308, 321, 326, 315, 
    304, 324, 306, 297, 311, 317, 322, 328, 324, 325, 330, _, 325, 321, 324, 
    332, 324, 321, 327, 321, 326, 328, 330, 329, 323, 326, 335, 326, 329, 
    333, 332, 331, 328, 329, 326, 326, 328, 330, 325, 324, 334, 331, 332, 
    289, 291, 353, 330, 338, 293, 348, _, 312, 40, _, _, 42, _, _, 44, 46, _, 
    45, 48, 49, _, _, 71, 65, 76, 83, 90, 100, 94, 97, _, 112, 116, 118, 132, 
    130, _, 132, 121, _, 115, 113, 111, 116, 108, 120, 116, 99, 88, 93, 92, 
    83, 83, 74, 62, 67, 72, _, 88, 102, 98, 105, _, 119, 130, 127, 140, 113, 
    115, _, 125, 120, _, 112, _, _, 113, 121, _, 122, 122, 117, 138, 122, 
    120, 118, 136, 125, 130, 124, _, 141, 139, _, 88, 68, 114, 117, 115, 141, 
    119, 99, _, _, 111, _, 83, 93, 79, 106, 139, _, 87, 101, 82, _, _, 85, _, 
    63, 55, 52, 67, 61, 57, 54, 54, 55, 66, 63, 57, 58, 59, 65, 72, 70, 67, 
    71, 72, 82, 75, 80, 84, 72, _, 72, 78, 83, 81, 75, 80, 70, 73, 72, 71, 
    69, 73, 81, 81, 83, 87, 95, 94, 81, 74, 83, 89, 89, 83, 74, 60, 56, _, 
    69, _, _, 53, _, 51, 53, _, 59, _, 63, 59, _, 52, _, 53, 319, 317, _, _, 
    _, _, _, _, 54, 48, 58, _, 47, 58, 51, _, 56, 58, 4, _, _, 345, _, 69, 
    352, 320, 302, 49, 91, 191, 340, 246, 108, 219, 333, _, 308, _, 73, 197, 
    185, _, 330, 291, _, _, _, 133, _, _, _, _, _, 50, 26, 35, 341, 293, 347, 
    352, 37, _, 71, 304, 66, 339, 262, _, 314, 281, 318, _, 288, 327, 284, 
    349, 327, _, 217, 316, _, _, _, 42, _, _, 55, 56, 65, 88, 81, 71, _, 79, 
    _, _, 73, 81, 99, _, 92, 100, 107, _, _, 118, _, 127, 122, 118, _, 125, 
    128, 115, 121, 128, 113, 148, _, 123, 123, _, 108, 101, 105, 110, 97, 98, 
    93, 99, 95, 96, 89, 93, 105, 106, 112, 110, 108, 108, 115, 119, 110, 110, 
    111, 108, 113, 103, 117, 102, 109, 103, 103, 112, 115, 117, 119, 114, 98, 
    106, 135, 117, 137, 108, 128, 309, 329, 292, 317, 322, 311, 305, _, 325, 
    314, 316, 317, 300, 334, 311, 332, 336, 61, 25, 174, 83, 57, 48, 94, _, 
    354, 3, 85, 177, 93, 197, 219, 179, 183, 84, 293, 294, 56, 49, 68, 69, 
    65, 67, 69, 73, 76, 77, 79, 78, 95, 89, 85, 83, 76, 76, 85, 72, 70, 72, 
    76, 82, 83, 103, 81, 91, 104, 87, 94, 99, 109, 115, 94, 94, 94, 99, 91, 
    91, 102, 114, 113, 111, 110, 115, 136, 135, 130, 146, 115, 132, 109, 113, 
    105, 110, 106, 107, 104, 108, 122, 120, 138, 137, 118, 103, 103, 111, 
    111, 114, 131, 136, 123, 109, 112, 105, 103, 105, 112, 112, 106, 107, 
    105, 110, 111, 106, 105, 101, 96, 90, 88, 113, 78, 64, 267, 330, 261, 2, 
    158, 12, 14, 1, 239, 25, 17, 343, 319, 331, 339, 328, 318, 307, 305, 312, 
    328, 332, 336, 330, 323, 314, 312, 335, 327, 325, 323, 322, 326, 330, 
    333, 327, 329, 340, 329, 318, 326, 326, 326, 327, 334, 322, 331, 327, 
    308, 311, 310, 304, 314, 313, 320, 349, 321, 150, 162, 121, 112, 114, 
    113, 97, 114, 145, 157, 168, 151, 165, 161, 181, 174, 183, 186, 181, 181, 
    163, 157, 163, 146, 165, 131, 110, 123, 128, 108, 109, 134, 135, 94, 104, 
    109, 142, 145, 85, 174, 159, 167, 133, 139, 126, 123, 111, 116, 115, 110, 
    106, 122, 111, 119, 110, 124, 116, 119, 112, 112, 115, 113, 110, 117, 
    118, 117, 108, 100, 106, 107, 117, 110, 22, 102, 344, 319, 323, 322, 321, 
    308, 337, 329, 327, 324, 327, 315, 286, 325, 37, 131, 123, 122, 119, 104, 
    114, 93, 134, 110, 115, 112, 125, 129, 103, 126, 114, 108, 126, 136, 110, 
    107, 149, 117, 133, 148, 146, 235, 294, 308, 312, 328, 310, 320, 303, 
    314, 317, 304, 302, 290, 300, 277, 276, 310, 300, 316, 285, 280, 293, 
    309, 307, 299, 305, 310, 305, 304, 305, 300, 303, 306, 296, 296, 295, 
    298, 293, 296, 298, 299, 299, 311, 311, 309, 314, 322, 310, 308, 316, 
    314, 317, 315, 313, 311, 304, 296, 292, 290, 303, 298, 315, 311, 311, 
    311, 314, 304, 291, 311, 308, 305, 325, 286, 274, 326, 345, 302, 351, 
    102, 181, 108, 71, 76, 82, 92, 117, 105, 109, 103, 86, 84, 68, 64, 76, 
    80, 79, 79, 81, 66, 63, 66, 65, 43, 20, 257, 8, 270, 270, 212, 347, 200, 
    235, 315, 91, 341, 138, 139, 325, 132, 23, 38, 105, 355, 232, 109, 43, 
    349, 323, 337, 331, 334, 333, 332, 315, 322, 328, 337, 317, 333, 323, 
    312, 322, 327, 321, 321, 325, 331, 331, 326, 319, 319, 318, 325, 324, 
    326, 327, 321, 314, 315, 326, 329, 318, 321, 319, 321, 312, 316, 320, 
    325, 318, 309, 306, 312, 309, 310, 303, 300, 304, 307, 306, 311, 307, 
    300, 296, 291, 286, 291, 299, 295, 292, 293, 296, 301, 310, 305, 293, 
    303, 299, 315, 302, 293, 294, 324, 336, 341, 346, 311, 242, 230, 227, 
    235, 222, 209, 209, 212, 204, 181, 181, 160, 156, 154, 161, 143, 144, 
    138, 128, 117, 118, 118, 164, 145, 131, 131, 115, 125, 137, 155, 144, 
    156, 179, 264, 320, 317, 321, 324, 326, 321, 326, 326, 335, 355, 336, 
    356, 8, 353, 2, 3, 359, 345, 357, 177, 20, 41, 32, 2, 3, 357, 323, 262, 
    257, 39, 21, 345, 355, 11, 36, 41, 17, 12, 20, 28, 13, 12, 31, 26, 6, 6, 
    294, 273, 263, 17, 9, 4, 10, 8, 9, 4, 360, 359, 1, 356, 352, 351, _, 348, 
    347, 340, 337, 339, 340, 341, 337, 337, 334, 332, 332, 336, 332, 334, 
    332, 328, 331, 325, 326, 328, 321, 322, 318, 319, 324, 317, 318, 323, 
    322, 328, 329, 327, 325, 331, 330, 334, 331, 331, 330, 331, 333, 330, 
    332, 332, 326, 324, 337, 338, 338, 335, 334, 336, 330, 322, 320, 324, 
    331, 327, 332, _, 317, _, 319, 316, 316, 321, 313, 314, 326, 325, 320, 
    305, 311, 314, 314, 308, 310, 324, 310, 318, 311, 311, _, 315, 308, 305, 
    302, 298, 304, 313, 306, 307, 292, 300, 292, 291, 288, 287, 293, 301, 
    285, 268, 258, 292, 297, 316, 312, 293, 262, 232, 4, _, 227, 230, 221, 
    233, 228, 61, 94, 68, 109, 108, 109, 118, 114, 112, 122, 122, 130, 151, 
    143, 125, 123, _, 99, 87, 87, 113, 136, 150, 144, 141, 138, 138, 127, 
    117, 100, 111, 105, 107, 106, 107, 115, 123, _, 120, 118, 111, 110, 111, 
    110, 104, 108, 125, 119, 112, 107, 107, 120, 136, 138, 262, 257, 253, 
    260, 264, 271, 265, 266, 272, 277, 286, 286, 297, 286, 283, 280, 283, 
    285, 289, 290, 289, 290, 288, 293, 291, 283, 287, _, 292, 285, 281, _, 
    295, 299, _, 290, 287, 282, 278, 296, 284, 265, 217, 176, 146, 156, 155, 
    144, 140, 143, 138, 143, 181, 204, 229, 276, 271, 269, 273, 286, 286, 
    300, 306, 295, 304, 310, 314, 306, 317, 282, 33, 101, 100, 90, 98, 109, 
    108, 83, 76, 65, 84, 84, 96, 101, 96, 96, 109, 136, 122, 122, 118, 106, 
    278, 297, 315, 311, 301, 306, 279, 241, 186, 179, 177, 159, _, 114, _, 
    102, 99, 110, 95, 85, 92, 84, 84, 85, 141, 0, 287, 322, 323, 314, 307, 
    314, 334, 237, 212, 130, 208, 184, 346, 22, 126, 99, 117, 115, 118, 114, 
    122, 122, 115, 117, 115, 112, 108, 100, 106, 115, 116, 114, 108, 113, 
    118, 110, 123, 123, 137, 120, 60, 316, 318, 313, _, 312, 311, 312, 310, 
    306, 319, 324, 316, 317, 309, 318, 321, 301, _, 352, 39, 7, 347, 76, 97, 
    103, 109, 102, 106, 115, 100, 109, 113, 156, 138, 143, 132, 139, 125, 
    121, 127, 131, 124, 136, 130, 129, 134, 126, _, 138, 141, 169, 148, 100, 
    81, 129, 54, 323, 296, 312, 306, 313, 319, 325, 326, 298, 115, 245, 97, 
    27, 343, 238, 253, 292, 326, 323, 311, 316, 316, 303, 314, 327, 311, 320, 
    315, 339, 122, 29, 92, 129, _, 84, 74, 79, 89, 75, 71, 75, 79, 116, 119, 
    100, 107, 118, 131, 132, 127, 122, 124, 124, 141, 133, 140, 145, _, 139, 
    146, 145, 130, 127, 123, 131, 133, 151, 157, 164, 174, 138, 235, 82, 144, 
    98, 95, 92, 89, 108, 98, 52, 15, 317, 332, 346, 327, 306, 294, 290, 287, 
    287, _, 265, 270, 285, 289, 287, 289, 290, 294, 289, 303, 305, 293, 277, 
    _, 89, 97, 104, 114, 120, 118, 113, 110, 120, 112, 109, 113, 120, 127, 
    119, 142, 132, 127, 134, 131, 134, 130, 135, 132, 131, 117, 129, 114, 
    131, 111, 117, 114, 125, 119, 114, 17, 293, 294, 314, 318, 315, 314, 316, 
    332, 323, 330, 335, 333, 332, 331, 338, 339, 333, 111, 1, 26, 296, 177, 
    303, 57, 47, 60, 52, 48, 55, 47, 62, 52, 341, 285, _, 284, 11, _, 321, 
    316, 352, 0, 332, 321, 308, 321, 318, 323, 313, 320, 316, 323, 3, 2, 340, 
    346, 336, _, _, _, _, _, _, _, 340, 335, 337, 333, 342, 341, 338, 345, 
    347, 349, 345, 352, 336, 349, 353, 353, 349, 342, _, 324, 320, 323, 337, 
    314, 311, 315, 321, 308, 295, 298, 324, 309, 257, 255, 284, 256, 216, 
    182, _, 155, 161, 162, 164, 177, 182, 178, 161, 149, 148, 141, 125, 129, 
    140, 123, 108, 113, 115, 117, 119, 159, 148, 122, 126, 124, 129, 139, 
    124, 118, 122, 122, 139, 168, 181, 176, 103, 118, 117, 123, 105, 124, 
    120, 127, 110, 115, 88, 74, 75, 117, 113, 108, 115, 120, 117, 111, 105, 
    97, 95, 96, 99, 92, 95, 104, 111, 159, 261, 269, 271, 271, 274, 274, _, 
    264, 268, 266, 266, _, 276, 277, 279, 280, 283, 284, 284, 277, 284, 276, 
    277, 279, 274, 272, 282, 287, 296, 303, 294, 298, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 306, 317, 318, 322, 313, 314, 316, 314, 318, 311, 
    313, 299, 314, 315, 328, 333, 340, 351, 353, 355, 11, 9, 6, 325, 80, 344, 
    90, 70, 78, 74, 80, _, 95, 93, 146, 121, 117, 108, 123, 127, 132, 148, 
    141, 132, 125, 128, 122, 109, 112, 110, 113, 102, 104, 105, 104, 109, 
    112, 111, 115, 119, 111, 126, 118, 108, 108, 114, 107, 114, 115, 119, 
    116, 116, 119, 115, 115, 112, 117, 120, 116, 112, 115, 122, 121, 155, 
    161, 142, 124, 107, 115, 111, 109, 109, 115, 116, 120, 123, 120, 120, 
    128, 136, 142, 117, 124, _, 123, 127, 132, 135, _, 140, 163, 150, 142, 
    129, 142, 136, 133, 138, 161, 166, 145, 143, 130, 119, 112, 118, 136, 
    125, 100, 98, 123, 97, 103, 83, 86, 102, 103, 105, 105, 100, 105, 114, 
    118, 121, 111, 102, 99, 109, 109, 105, 103, 98, 97, 76, 71, 69, 70, 78, 
    76, 67, 61, 58, 58, 56, 59, 61, 67, 70, 65, 65, 71, 73, 65, 71, 88, _, 
    92, 95, 76, 83, 78, 73, 77, 65, 76, 56, 60, 71, 78, 70, 76, 64, 77, 85, 
    77, 85, 77, 70, 94, 86, 87, 79, 85, 93, 81, 100, 83, 75, 67, 76, 76, 83, 
    97, 102, 101, 105, 93, 82, 98, 109, 119, 118, 114, 110, 118, 115, 109, 
    119, 106, 100, 102, 107, 121, 116, 121, 113, 101, 101, 92, 94, 102, 101, 
    96, 90, 92, 93, 90, 90, 85, 82, 82, 83, 84, 88, 96, 96, 103, 105, 107, 
    104, 105, 103, 101, 101, 96, 96, 91, 87, 90, 90, 91, 93, 88, 86, 77, 65, 
    60, 71, 73, 38, 59, 61, 65, 64, 69, 77, 80, 66, 82, 84, 82, 71, 63, 75, 
    81, 89, 86, 84, 99, 134, 147, 176, 243, 319, 316, 344, 342, 322, 37, 20, 
    67, 96, 108, 103, 115, 126, 118, 159, 144, 135, 117, _, _, 145, 130, 135, 
    130, 138, _, 114, 105, _, 115, 128, 194, 200, 277, 287, 338, 312, 318, 
    338, 330, 349, 338, 342, 338, 337, 337, 332, 324, 321, 320, 315, 327, 
    324, 325, 327, 324, 320, 319, 318, 318, 304, 305, 283, 303, 297, 299, 
    296, 300, 293, 311, 323, 304, 359, 5, 23, 22, 32, 42, 51, 57, 13, 31, 25, 
    33, 23, 22, 14, 30, 25, 24, 30, 32, 35, 34, 51, 55, 59, 81, 73, 78, 71, 
    81, 76, 79, 80, 69, 88, 86, 75, 73, 73, 70, 77, 63, 68, 79, 73, 66, 60, 
    62, 63, 75, 79, 84, 81, 77, 72, 75, 77, 79, 88, 84, 92, 88, 81, 74, 82, 
    _, 84, 84, 87, 69, 64, 68, 68, 79, 73, 71, 70, 66, 67, 66, 61, 63, 61, 
    102, 74, 89, 76, 80, 83, 93, 95, 90, 94, 75, 78, 74, 65, 65, 61, 63, 68, 
    109, 96, 81, 73, 60, 63, 66, 59, 49, 42, 38, 27, 20, 8, 5, 353, 341, 334, 
    340, 334, 333, 335, 334, 336, 334, 326, 331, 329, 330, 332, 330, 334, 
    338, 329, 328, 327, 330, 326, 333, 325, 323, _, 323, 316, 318, 314, 315, 
    339, 323, 327, 4, 21, 15, 24, 65, 88, 69, 77, 85, 83, 6, 299, 305, 307, 
    309, 311, 300, 294, 304, 311, 308, 295, 306, 311, 307, 317, 306, 303, 
    303, 314, 313, 316, 317, 306, 306, 304, 297, 302, 303, 304, 306, 300, 
    307, 306, 303, 308, 302, 306, 311, 308, 311, 311, 294, 305, 300, 293, 
    302, 305, 311, 319, 301, 327, 315, 316, 356, 31, 59, 71, 66, 62, 67, 82, 
    82, 91, 94, 88, 91, 92, 84, 85, 83, 81, 79, 85, 90, 89, 93, 101, 107, 
    114, 114, 110, 111, 114, 118, 115, 112, 112, 116, 114, 106, 107, 112, 
    103, 120, 118, 121, 110, 115, 114, 116, 110, 120, 111, 120, 105, 122, 
    121, 121, 114, 109, 111, 110, 119, 135, 125, 121, 109, 111, 112, 112, 
    116, 115, _, 111, 112, 111, 103, 96, 123, 47, 18, 299, 341, 303, 345, 
    336, 56, 54, 50, 47, 32, 308, 339, 119, _, 329, 330, 7, 330, 332, 335, 
    338, 335, 334, 334, 333, 334, 340, 341, 338, 337, 346, 340, 347, 2, 2, 1, 
    2, 3, 353, 4, 337, 337, 342, 331, 331, 338, 336, 342, 339, 337, _, 328, 
    334, 331, 314, 320, 322, 324, 319, 326, 313, 315, 320, 317, 322, 325, 
    322, 327, 336, _, 320, 318, 308, 312, 295, 304, 311, 318, 312, 311, 318, 
    65, 104, 109, 241, 309, 289, 289, 296, 286, 273, 234, 240, 240, 281, 295, 
    273, 292, 279, 286, 254, 233, 223, 224, 223, 233, 236, 241, 285, 287, 
    280, 4, 82, 232, 235, 241, 239, 243, 248, 240, 238, 231, 214, 212, 207, 
    180, 186, 180, 174, 190, 166, 152, 161, 165, 179, 194, 186, 185, 182, 
    176, 174, 161, 169, 158, 153, 156, 146, 129, 128, 137, 133, 128, 125, 
    116, 123, _, 124, _, 125, 123, 124, 121, 122, 130, 132, 137, 128, 122, 
    132, 139, 139, 128, 123, 128, 139, 133, 130, 122, 130, 126, 132, 124, 
    123, 120, 115, 132, 116, 109, 113, 119, 116, 115, 117, 116, 119, 122, 
    121, 124, 124, 125, 125, 118, 124, 117, 119, 121, 114, 116, 118, 121, 
    123, 121, 121, _, 125, 125, 127, 126, 126, 129, 132, 134, 137, 138, 141, 
    139, 137, _, 130, 132, 132, 137, 137, 137, 136, 135, 134, 139, 136, 135, 
    134, 134, 133, 132, 132, 134, 134, 133, 140, 137, 137, 138, 134, 128, 
    128, 130, 128, 134, 139, 138, 139, 141, 143, 140, 144, 143, 125, 120, 
    121, 124, 125, _, 121, 126, 121, 120, 119, 106, 114, 111, 106, 96, 86, 
    99, 100, 86, 80, 73, 77, 77, 90, 92, 89, 86, 82, 81, 94, 90, 94, _, 87, 
    98, 90, 80, 82, 86, 85, 82, 80, 83, 78, 76, 72, 75, 77, 75, 71, 74, 71, 
    75, 78, 79, 81, 91, 95, 101, 101, 97, _, 105, 113, 107, 107, 107, 112, 
    110, 107, 100, 105, 101, 111, 108, 105, _, 95, _, 95, 97, 95, 92, 94, 93, 
    94, 95, 103, 100, 106, 104, 106, 130, 130, 125, 137, 142, 136, 142, 142, 
    144, 162, 147, 150, _, 148, 153, 183, 171, 180, 181, 170, 106, 105, 133, 
    228, 284, 298, 292, 298, 290, 293, 295, 293, 300, 288, 283, 290, 284, 
    269, 284, 278, 296, 284, 263, 256, 243, 251, 230, 264, 265, 263, 290, 
    296, 288, 335, 310, 305, _, 331, 339, 333, 336, 337, 335, 335, 328, 332, 
    337, 334, 332, 323, 136, 64, 63, 29, 351, 354, 336, 314, 314, 307, 267, 
    263, 257, 260, 255, 259, 259, 264, 265, 261, 261, 265, 259, 264, 268, 
    256, 261, 261, 255, 244, 252, 242, 245, 253, 259, 265, 262, 262, 260, 
    260, 283, 276, 274, 288, 311, 28, 32, 27, 47, 61, 64, 65, 74, 69, 61, 89, 
    213, 184, 162, 164, 163, _, 140, 134, 127, 125, 285, 285, 283, 279, 274, 
    272, 251, 238, 208, 204, 183, 191, 167, 147, 99, _, 33, 5, 3, 1, 337, 45, 
    47, 30, 2, 22, 344, 4, 7, 20, 316, 311, 315, 323, 322, 318, 316, 314, 
    323, 315, 320, 342, 3, 11, 360, 23, 344, 16, 10, 13, 19, 23, 31, 26, 42, 
    45, 62, 77, 53, 53, 50, 48, 41, 29, 41, 54, 53, 50, 63, 57, 66, 99, 104, 
    108, 111, 117, 121, 129, 129, 122, 108, 99, 102, 120, 119, 123, 122, _, 
    114, 111, 100, 95, _, 92, 83, 88, 84, 77, 85, _, 90, 88, 92, 85, 87, 83, 
    74, 77, 74, 71, 68, 69, 59, 44, 42, 34, 39, 49, 57, 43, 31, 33, 35, 28, 
    29, 31, 38, 39, 38, 36, 45, 41, 37, 35, 26, 35, 38, 45, 38, 35, 34, 40, 
    34, 38, 48, 45, 53, 52, 36, 43, 27, 37, 39, 20, 29, 40, 38, 38, 22, _, 
    43, 44, 39, 45, 50, 51, 51, 51, 51, 47, 48, _, 49, 52, 52, 58, 65, 69, 
    70, 70, 73, 76, 78, 77, 85, 91, 82, _, 94, 97, 90, 96, 85, _, 81, 89, 94, 
    89, _, 86, _, 87, 82, 75, _, _, 78, 73, 80, 79, 82, 81, _, _, 97, _, 105, 
    101, 102, 108, 109, _, 117, 124, 123, 123, 118, 118, 111, 112, 111, 109, 
    _, 114, 113, 105, _, 106, _, _, 113, 114, 109, 107, 102, _, 98, 94, 92, 
    86, _, _, _, 89, 88, 88, 85, 87, 95, 103, 106, 107, 106, 113, 105, 101, 
    96, 95, 93, 92, 96, 99, 93, 83, 83, 87, 91, 93, 98, 94, 96, 98, 93, 92, 
    89, 84, 84, 92, 92, 86, 81, 82, 81, 74, 72, 69, 71, 73, 88, 94, 83, 83, 
    90, 85, 83, 81, 73, 75, _, 70, 69, 66, 69, 69, 69, 67, 46, 40, 42, 26, 
    43, 43, 44, 46, 45, 47, 44, 44, 44, 41, 31, 330, 2, 67, 64, 60, _, 42, 
    42, 44, 40, 43, 40, 41, 37, 31, 7, 11, 14, 5, 6, 2, 9, 3, 6, 27, 19, 10, 
    15, 11, 6, 5, 16, 6, 10, 1, 1, 21, 12, 12, 13, 20, 355, 9, 356, 22, 21, 
    22, 2, 28, _, 11, 31, 34, 35, 34, 26, _, 32, 37, 19, 45, 64, 320, 24, 27, 
    21, 355, 12, 332, 353, 346, 317, 326, 318, 316, 320, 306, 305, 314, 311, 
    314, 319, 312, 320, 287, 304, 352, 17, 24, 45, 60, 83, 81, 69, 71, 68, 
    66, 68, 68, 75, 76, 78, 80, 83, 87, 87, 79, 79, 86, 56, 53, 51, 45, 39, 
    14, 10, 342, 342, 308, 303, 299, 315, 316, 319, 309, 324, 317, 321, _, 
    304, 322, 317, 314, 310, 314, 313, 318, 313, 315, 312, 310, 304, 318, 
    315, 307, 308, 304, 318, 313, 316, 318, 311, 308, 307, 307, 310, 319, 
    305, 303, 296, 301, 332, 356, 348, 358, 321, 311, 322, 325, 322, 328, 
    303, 46, 25, 32, 27, 27, 40, 45, 54, 46, 39, 40, 52, 44, 42, 27, 13, 38, 
    42, 33, 34, 41, 43, 42, 39, 45, 33, 34, 22, 19, 5, 352, 344, 339, 339, 
    350, 353, 355, _, 3, 3, _, 4, 6, 7, 6, 5, 2, _, 2, _, 358, 351, _, 356, 
    351, _, 355, _, _, 2, _, 2, 357, 351, 356, 351, 355, _, 354, 357, 354, 
    357, 344, 358, 353, 6, 254, 312, 27, 56, 296, 354, 29, 39, 77, 29, 32, 
    32, 37, 48, 70, 20, 62, 81, 152, 100, 82, 95, 90, 76, 77, 79, 76, 68, 66, 
    70, 78, 72, 71, 71, 71, 70, 63, 72, 74, 66, 58, 65, 64, 63, 56, 50, 61, 
    72, 76, 70, 71, 73, 72, 73, 72, 69, 72, 69, 72, 71, 73, 74, 80, 81, 75, 
    74, 73, 75, 76, 77, 75, 75, 73, 69, 69, 90, 83, 81, 82, 81, 75, 67, 70, 
    64, 66, 74, 77, 73, 69, 80, 77, 73, 80, 75, 75, 77, 83, 80, 78, 85, 79, 
    75, 69, 69, 64, 58, 54, 55, 54, 52, 47, 42, 40, 30, 26, _, 23, _, _, _, 
    18, _, _, 3, _, 354, 354, 349, 342, 347, _, _, 342, 332, 342, 334, 316, 
    _, _, 315, 311, _, _, 310, _, _, _, 310, 319, 319, _, 317, _, 312, 305, 
    324, _, _, _, _, 28, 43, 65, 65, _, 70, 81, 73, 79, _, 82, _, _, 116, 
    129, 136, 140, 129, 123, _, 123, _, 108, 93, _, _, 30, 32, 32, 22, 24, 
    23, 22, 17, 16, 20, _, 15, 15, 15, 17, 16, 11, 22, 18, 19, 22, 13, 14, 
    12, 3, 359, 338, 334, _, 320, 307, 301, 295, 301, 308, 309, 312, 295, 
    294, 299, 302, 302, 308, _, 305, 319, 323, _, 324, 321, 324, 324, _, 316, 
    311, 315, _, _, 313, _, 313, 313, 308, 304, 307, 309, _, _, 304, 305, 
    302, _, 299, 298, _, _, 298, 313, _, 4, 17, 46, 69, _, 93, 107, _, 105, 
    _, 86, _, 73, 83, 81, 58, 71, 80, 91, 90, 101, 100, 108, _, 111, 121, 
    112, 116, 110, _, 114, 120, 120, 116, _, 116, 114, 118, 125, 124, 122, 
    121, 118, 121, 119, 125, 127, _, 115, 144, _, 136, 141, 139, 140, 137, 
    136, 136, 131, _, _, 136, 135, _, 115, 110, 121, 124, _, _, 112, 116, 
    117, 65, 117, 116, 114, 127, 133, 118, 107, 109, 137, 142, 107, 170, _, 
    120, _, _, 107, 96, 132, 113, 117, 107, 105, _, _, _, 116, 116, _, 117, 
    126, 147, _, 157, _, 165, _, 133, 164, 192, 151, 149, _, _, 134, 132, _, 
    152, _, _, _, 187, _, _, _, 311, 296, _, 281, _, _, 322, 114, 124, 117, 
    114, 120, 121, 152, _, 128, 134, 143, _, _, 142, 145, _, _, 156, _, 163, 
    _, _, 175, _, 182, 180, 188, _, _, 119, 140, 113, 34, 18, 358, 341, 330, 
    272, 301, 304, 295, 323, 327, _, 315, _, 311, _, 326, 340, 5, _, 11, 13, 
    79, _, 87, 89, 119, _, _, _, _, _, _, _, 172, 240, 208, 50, 25, 114, 71, 
    357, 43, 13, 16, 356, _, 343, 350, 342, 359, 1, 3, 6, 11, 11, 3, 357, 
    337, 28, 22, 31, 20, 18, 17, 10, 13, 10, 22, 19, 344, 17, 16, 15, 17, 23, 
    8, 44, 42, 46, 53, 50, 47, 52, 59, 53, 37, 38, 47, 44, 45, 42, 43, 45, 
    46, 48, 51, 46, 38, 33, 25, 19, 24, 30, 38, 42, 49, 46, 43, 45, 46, 48, 
    49, 42, 54, 35, 29, 27, 28, 28, 33, 39, 40, 42, 43, 40, 32, 30, 27, 22, 
    18, 15, 12, 20, 25, 24, 36, 21, 20, 18, 18, 20, 23, 23, 34, 44, 55, 56, 
    53, 45, 48, 51, 66, 69, 79, 74, 87, 86, 93, 99, 106, 98, 87, 99, 102, 88, 
    91, 83, 86, 77, 83, 80, 79, 84, 85, 83, 78, 77, 79, 81, 84, 70, 49, 29, 
    22, 16, 10, 13, 18, 12, _, 16, 11, 360, 2, 2, 358, 358, 337, 322, 328, 
    327, 323, 325, 311, 309, 317, 317, 313, 314, 312, 308, 312, 309, 308, 
    304, _, 310, 313, 305, 302, 305, 288, 284, 274, 273, 268, 273, 283, 275, 
    271, 271, 269, 268, 252, 223, 222, 229, 224, 222, 289, 321, 344, 8, 31, 
    29, 38, 39, 50, 64, 64, 54, 51, 69, 67, 62, 346, 5, 7, 347, 357, 12, 14, 
    13, 16, 23, 31, 42, 58, 61, 58, 57, 53, 54, 54, 56, 56, 58, 59, 62, 73, 
    71, 73, 81, 86, 97, 99, 100, 99, 95, 94, 96, 97, 97, 92, 92, 93, 80, 107, 
    88, 79, 103, 108, 106, 102, 89, 99, 101, 105, 100, 95, 100, 109, 108, 97, 
    94, 97, 111, _, 113, 113, 112, 121, 107, 99, 108, 102, 107, 112, 104, 92, 
    93, 105, 111, 111, 114, 113, 113, 110, 118, 113, 117, 117, 120, 117, 119, 
    106, 108, 103, 105, 100, 107, 105, 102, 112, _, _, 123, 122, 117, 110, 
    101, 99, 103, 108, 108, 116, 116, 125, 111, 107, 97, 95, 102, 105, 113, 
    113, 113, 107, 113, 111, 112, 116, 112, 120, 138, 151, 145, 123, 148, 
    176, 175, 234, 103, 85, 76, 7, 26, 86, 100, 99, 123, 118, 114, 101, 113, 
    125, 136, 106, 96, 92, 111, 125, 158, 117, 118, 100, 178, 137, 115, 124, 
    106, 103, 107, 116, 109, 103, 104, 94, 94, 96, 93, 157, 235, 304, 357, 4, 
    29, 115, 145, 91, 105, 119, 102, 119, 110, 83, 78, 66, 73, 78, 67, 84, 
    95, 121, 106, 110, 125, 116, 115, 116, 112, 110, 107, 116, 113, 116, 117, 
    118, 113, 119, 126, 122, 118, 139, 117, 132, 138, 131, 126, 121, 126, 
    132, 146, 144, 146, 148, 143, 143, _, 148, 157, 148, 144, 141, 139, 140, 
    142, 145, 141, 141, 138, 139, 139, 137, 143, 138, 139, 139, 138, 140, 
    138, 134, 135, 136, 128, 126, 131, 126, 124, 120, 106, 111, 121, 116, 
    111, 104, 101, 96, 78, 78, 69, 63, 61, 61, 62, 56, 56, 67, 58, 52, 43, 
    46, 53, 60, 60, 60, 58, 53, 54, 60, 68, 63, 85, 77, 84, 75, 86, 84, 77, 
    77, 75, 73, 69, 78, 72, 71, 66, 57, 65, 60, 64, 61, 60, 61, 57, 59, 52, 
    55, 54, 53, 56, 57, 66, 65, 57, 49, 47, 50, 54, 52, 61, 63, 64, 65, 63, 
    61, 62, 67, 67, 65, 70, 79, 86, 94, 110, 99, 94, 82, 68, 69, 64, 56, 57, 
    64, 63, 66, 73, 67, 59, 55, 53, _, 62, 62, 59, 59, 58, 59, 58, 53, 46, 
    39, _, 30, 15, 9, 20, 13, 19, 26, 35, 34, 39, 44, 52, 52, 50, 46, 40, 45, 
    34, 40, 43, 43, 43, 52, 53, 62, 66, 59, 50, 47, 48, 54, 54, 52, 54, 49, 
    51, 47, 45, 47, 50, 48, 45, 43, 44, 48, 47, 40, 44, 51, 45, 48, 42, 36, 
    35, 45, 48, 43, 59, 62, 64, 58, 51, 42, 40, 35, 40, 34, 32, 39, 43, 44, 
    _, 40, 41, 37, 40, 38, 39, 38, 30, 27, 34, 32, 26, 26, 38, 39, 52, 52, 
    53, 57, 57, 60, 61, 62, 58, 314, 32, 33, 43, 46, 44, 44, 49, 285, 360, 
    38, 34, 29, 356, 14, 5, 1, 339, 358, 349, 347, 358, 5, 349, 359, 3, 359, 
    359, 342, 360, 341, 338, 342, 342, 342, 2, _, 4, 33, 19, 46, 42, 53, 55, 
    56, 40, 8, 36, 23, 60, 28, 53, 55, 58, 64, 72, 51, 28, 22, 4, 13, 17, 9, 
    26, 26, 29, 36, 38, 85, _, 58, 47, 56, 25, 43, 43, 13, 1, 16, 16, 10, 11, 
    6, 17, 19, 12, 17, 9, _, 43, 26, 67, 60, 45, 43, 57, 67, 62, 61, 56, 25, 
    25, 48, 59, 41, 56, 43, 50, 40, 51, 47, 44, 51, 50, 47, 47, 47, 40, 36, 
    _, 19, 29, 27, 44, 54, 53, 48, 40, 29, _, 28, 20, 17, 19, 16, 3, 349, 
    354, 358, _, 2, 3, 2, 3, 5, 8, 5, 4, 339, 340, 350, 340, 349, 347, 336, 
    331, 317, 309, 297, 294, 282, 277, 281, 273, 276, 264, 262, 257, 243, 
    242, 239, 236, 246, 267, 242, 253, 251, 242, 237, 224, 221, 200, 180, 
    184, 179, 194, 197, 220, 202, 209, 204, _, 197, 217, 215, 212, 198, 200, 
    201, 217, 231, 230, 232, 234, 44, 18, 273, 234, 229, 235, 261, 253, 250, 
    249, 244, 225, 218, 168, 183, 176, 182, 227, 201, 217, 231, 237, 233, 
    236, 225, 209, 240, 237, 263, 263, 271, 262, 262, 260, 263, 254, 260, 
    262, 257, 232, 224, 187, 151, 139, 131, 134, 113, 103, 115, 101, 96, 102, 
    112, 117, 125, 124, 117, 114, 112, 112, 114, 110, 100, 95, 96, 104, 104, 
    93, 87, 82, 82, 85, 84, 88, 90, 86, 86, 84, 88, 95, 97, 98, 99, 100, 99, 
    98, 99, 96, 98, 99, 101, 100, 92, 94, 90, 88, 88, 87, 90, 94, 93, 93, 96, 
    104, 97, 98, 98, 96, 93, 97, 95, 99, 100, _, 84, 82, 91, 95, 83, 82, 75, 
    65, 52, 71, 82, 98, 99, 84, 88, 81, 62, 53, 55, 93, 99, 114, 137, 123, 
    102, 118, 130, 119, 105, 99, 101, 93, 92, 86, 89, 103, 101, 100, 100, 
    102, 99, 116, 115, 115, 117, 101, 86, 90, 85, 84, 87, 92, 86, 88, 92, 89, 
    81, 77, 82, 84, 86, 92, 96, 103, 109, 111, 132, 128, 124, 130, 136, _, 
    129, 123, 122, 113, 90, 86, 104, 93, 106, 117, 107, 108, 112, 110, 117, 
    108, 124, 137, 122, 111, 108, 111, 124, 147, 125, 133, 163, 121, 151, 
    126, 112, 102, 94, 118, 103, 82, 22, 63, 57, 61, 61, 74, 81, 79, 78, 80, 
    69, 62, 70, 74, 78, 94, 104, 106, 104, 103, 101, 109, 106, 109, 106, 106, 
    107, 110, 103, 107, 99, 103, 99, 99, 90, _, 70, 59, 55, 55, 59, 79, 91, 
    100, 64, 74, _, 75, 71, 76, 80, 89, 92, 85, 77, 79, 67, 60, 48, 47, 44, 
    60, 60, 48, 42, 37, 36, 37, 30, 21, 34, 25, 19, 5, 12, 16, 6, 1, 360, 5, 
    1, 17, 44, 14, 8, 20, 12, 29, 36, 12, 4, 20, 49, _, 28, 15, 28, 28, 22, 
    12, 2, 24, 28, 19, 11, 22, 13, 16, 13, 26, 13, 23, 13, 18, 38, 26, 19, 
    28, _, 25, 21, _, 18, 18, 22, 30, 25, 29, 35, 16, 92, 69, 30, 66, 62, 51, 
    48, 44, 78, 59, 52, 32, 44, 360, 29, 62, 54, 58, 53, 50, 51, 50, 53, 54, 
    52, 54, 54, 48, 51, 59, 51, 52, 53, 52, 52, 52, 62, 50, 10, 34, 29, 26, 
    42, 23, 54, 49, 27, 44, 65, 56, 53, 55, 58, 58, 59, 58, 61, 59, 57, 57, 
    63, 68, 96, 110, 99, 96, 106, 84, 83, 80, 87, 87, 80, 79, 81, 97, 121, 
    110, 99, 112, 101, 97, 88, 90, 91, 88, 88, 93, 93, 92, 103, 98, 91, 89, 
    117, 115, 107, 107, 106, 105, 104, 98, 97, 105, 109, 106, 109, 112, 116, 
    115, 117, 117, 122, 122, 120, 117, 118, 115, 110, 111, 104, 104, 109, 
    113, 113, 114, 115, 114, 117, 116, 118, 116, 115, 114, 108, 112, 114, 
    112, 116, 121, 123, 126, 127, 128, 126, 124, 125, 122, 119, 119, 118, 
    120, 124, 125, 120, 116, 107, 106, 103, 100, 92, 85, 92, 96, 101, 96, 89, 
    94, 98, 97, 106, 118, 112, 155, 188, 198, 192, 193, 184, 181, 65, 156, 
    130, 140, 142, 141, 5, 90, 0, 316, 267, 288, 310, 248, 217, 274, 13, 128, 
    110, 157, 145, 166, 199, 208, 254, 329, 324, 328, 349, 347, 340, 331, 
    311, 317, 330, 336, 17, _, 44, 81, 88, 103, 95, 175, 134, 155, 154, 155, 
    164, 132, 137, 139, 127, 148, 124, 125, 117, 108, 105, 96, 94, 81, 83, 
    91, 97, 106, 108, 111, 115, 94, 96, 77, 74, 64, 61, 64, 78, 112, 110, 82, 
    67, 64, 54, 56, 50, 51, 58, 60, 61, 81, 102, 88, 76, 60, 61, 58, 64, 55, 
    59, 74, 90, 95, 88, 85, 81, 87, 80, 87, 66, 61, 55, 44, 34, 48, 39, 8, 
    348, 145, 12, 355, 303, 353, 10, 3, 238, 50, 96, 107, 115, 98, 104, 118, 
    115, 119, 116, 119, 136, 124, 123, 116, 139, 143, 143, 129, 126, 127, 
    118, 119, 120, 121, 124, 119, 124, 137, 138, 129, 126, _, 131, 128, 131, 
    125, 131, 129, _, 135, 143, 136, 131, _, 127, 138, 134, 131, 107, 193, 
    174, 159, 157, 112, 117, 127, 113, 142, 141, 139, 120, 121, 119, 113, 
    114, 124, 125, 130, 137, 146, 163, 153, 180, 203, 190, 184, 119, 109, 
    127, 267, 292, 308, 300, 294, 300, 289, 294, 296, 298, 286, 287, 292, 
    290, 295, 323, 90, 97, 111, 108, 100, 97, 76, 67, 69, 63, 55, 33, 23, 13, 
    359, 353, 339, 332, 330, 329, 316, 319, 326, 317, 315, 306, 321, 322, 
    314, 314, 315, 313, 312, 309, 319, 317, _, 308, 306, 309, 309, 310, 312, 
    309, 311, 306, 307, 307, 309, 305, 313, 322, 322, 315, 322, 317, 318, 
    315, 316, 327, 325, 323, 319, 317, 321, 317, 317, 319, 320, 333, 311, 
    318, 313, 310, 311, 322, 318, 320, 332, 336, 336, 342, _, 341, 337, 344, 
    1, 2, 351, 3, 2, 357, 352, 351, 354, 340, _, 349, 337, 332, 334, 335, 
    326, 323, 322, 323, 321, 322, 344, 341, 345, 340, 4, 3, 345, 4, 32, 31, 
    23, 21, 18, 12, 12, 9, 20, 29, 13, 2, 2, 1, 9, 8, 8, 1, 355, 343, 350, 
    349, 349, 351, 343, 338, 321, 305, 310, 304, 301, 300, 311, 305, 309, 
    305, 302, 303, _, 304, 309, 311, 307, 306, 300, 304, 306, 299, 307, 308, 
    307, 307, 308, 298, 294, 300, 296, 293, 283, 286, 287, 299, 292, 295, 
    297, 290, 288, 307, 339, 330, 284, 337, 2, 33, 27, 13, 9, 20, 7, 6, 17, 
    14, 8, 3, 14, 1, 360, 11, 1, 20, 30, 22, 4, 350, 40, 56, 66, 63, 44, 26, 
    63, 45, 46, 44, 54, 54, 46, 28, 53, 52, _, 61, 53, 55, 55, 83, 83, 96, 
    97, 97, 67, 45, 48, 36, 42, 44, 29, 9, 62, 82, 5, 323, 37, 44, 53, 61, 
    62, 85, _, 110, 103, 106, 102, 102, 88, 94, 94, 93, 96, 102, 103, 105, 
    106, 105, 104, 113, 119, 117, 118, 123, 116, 117, 106, 88, 311, 110, 88, 
    74, _, 90, 82, 73, 92, 87, 101, 89, 87, 98, 87, 85, 70, 73, _, 62, 64, 
    64, 65, 63, 71, 83, 77, 78, 82, 69, 82, 82, 90, 90, 86, 82, 79, 81, 79, 
    79, 81, 79, 82, 85, 83, 81, 77, 74, 75, 73, 69, _, 70, 74, 75, 70, 69, 
    81, 85, 84, 78, 75, 74, 77, 76, 77, 71, 72, 74, 79, 63, 78, _, 69, 70, 
    82, 154, 159, 165, 125, 119, 113, 112, 99, 110, 98, 82, 76, 67, 73, 55, 
    53, 50, 32, 17, 357, 355, 350, 353, 359, 350, _, 18, 14, 1, 1, 359, 357, 
    359, 2, 356, 348, 360, 349, 355, 355, 359, 359, 355, 360, 345, 336, 337, 
    _, 323, 327, 330, 336, 338, _, 329, 322, 323, 326, 320, 322, 320, 316, 
    314, 321, 319, 316, 319, 326, 324, 323, 344, 354, 334, 296, 300, 302, 
    306, 308, 312, 313, 307, 343, 353, 358, 26, 98, 112, 86, _, 93, 118, 163, 
    151, 160, 147, 160, 173, _, 104, 109, 106, 100, 99, 114, 114, 120, 120, 
    111, 112, 107, 119, 104, 122, 124, 112, 111, 109, 118, 112, _, 112, 131, 
    111, 209, 215, 184, 233, 270, 24, 301, 337, 329, _, 345, 2, 331, 335, 24, 
    324, 321, 315, 325, 320, 326, 325, 77, 58, 60, 59, 56, 59, 53, 55, 57, 
    54, 52, 52, 51, 52, 52, 61, _, 64, 62, 72, 72, 72, 97, 72, 72, 75, 68, 
    69, 63, 77, 70, 306, 11, 354, 345, 15, 3, 5, 90, 90, 78, 103, 106, 123, 
    163, 141, 211, 259, 357, 56, 138, 117, 86, 104, 115, 120, 108, 115, _, 
    124, 120, 121, 120, 116, 119, 127, 129, 125, _, 136, 171, 172, 219, 198, 
    255, 273, 290, 305, 327, 351, _, 299, 315, 336, 353, 18, 23, 24, 36, 291, 
    303, 334, 246, 68, 67, 69, 74, 75, 81, 94, 86, 105, 124, 127, 117, 163, 
    167, 162, 146, 138, 184, 130, 166, 126, 144, 133, 156, 177, 154, 200, 
    190, 211, 227, 226, 4, 341, 343, 350, 355, 340, 348, 318, 322, 317, 328, 
    321, 314, 314, 313, 308, 302, 297, 314, 299, 300, 326, 317, 302, 326, 
    325, 324, 323, 321, 313, 307, 317, 304, 303, 303, 311, 306, 308, 305, 
    311, 307, 311, 312, 311, 306, 305, 313, 330, 345, 346, 348, 352, 349, 
    348, 346, 347, 346, 342, 350, 354, 351, 351, 351, 346, 350, 346, 355, 
    345, 339, 338, 348, 342, 336, 336, 334, 333, 339, 339, 340, 338, 338, 
    340, 329, 336, 333, 339, 350, 337, 351, 344, 345, 344, 347, 338, 341, 
    344, 342, 340, 345, 347, 334, 334, 343, 334, 349, 333, 333, 347, _, _, 
    343, 342, 349, 335, 334, 341, 339, 334, 334, 321, 347, 339, 343, 352, 
    358, 358, 343, 343, 335, 337, 340, 332, 345, 333, 335, 334, 321, 333, 
    329, 332, 334, 338, _, 353, 336, 337, 337, 337, 337, 340, 335, 336, 334, 
    329, 336, 337, 331, 334, 332, 337, 338, 318, 336, 334, 342, 333, 339, 
    341, 1, 3, _, 359, 358, 2, 359, 354, 359, 1, 7, 1, _, _, 337, 320, 316, 
    317, 17, 8, 331, 8, 7, 357, 357, 21, 337, 14, 8, 8, 5, 1, 7, 353, 8, 8, 
    21, 360, 345, 316, 324, 2, 326, 333, 337, 337, 327, 332, 33, 30, 17, 1, 
    355, 340, 333, 330, 329, 326, 325, 326, 322, 319, 314, 314, 317, 319, 
    307, 312, 5, 336, 325, 323, 316, 312, _, 310, 318, 303, 300, 304, 304, 
    301, 308, 295, 293, _, 282, 283, _, 287, 282, 287, 287, 300, 284, 288, 
    302, 308, 307, 285, 284, 282, 280, 276, 281, 280, 283, 310, 301, 309, 
    307, 306, 306, 306, 318, 311, 312, 323, 320, 308, 331, 351, 3, 359, 19, 
    360, 44, 59, 80, 49, 49, 55, 56, 52, 55, 65, 67, 69, 67, 73, 82, 69, 74, 
    75, 80, 75, _, 82, 92, 95, 93, 107, 80, 80, 87, 76, 60, _, 28, 52, _, 
    354, 338, 334, 328, 315, 318, 337, 352, 339, 329, 335, 338, 333, 329, 
    324, 319, 312, 331, 322, 328, 324, 325, 326, 325, 332, 331, 325, 333, 
    326, 318, 325, 321, 321, 328, 326, 325, 321, 324, 322, 318, 314, 312, 
    312, 309, 303, 307, 295, 305, 308, 303, 289, 305, 303, 303, 306, 312, 
    307, _, 312, 319, 311, 327, 338, 352, 4, 18, 41, 70, _, 104, 119, 189, 
    182, 170, 149, 175, 144, 140, 133, 112, 97, 82, 71, 66, 51, 52, 55, 64, 
    67, 55, 339, 64, 38, 51, 327, 40, 338, 343, 335, 327, 26, 342, 343, 76, 
    _, 92, 13, 58, 5, 2, 324, 104, 1, 341, 347, 0, 133, 6, 330, 355, 123, 
    121, 153, 115, 132, 359, 325, 294, 296, _, 319, 321, 312, 308, 313, 306, 
    311, 309, 314, 318, 302, 314, 326, 319, 333, 335, 27, 357, 51, 107, 170, 
    132, 123, _, 243, 268, 295, 296, 329, 354, 285, 281, 332, 325, 360, 79, 
    110, 113, 129, 152, 148, 125, 131, 122, 127, 134, 148, 140, 140, 146, 
    166, 159, 185, 212, 313, 320, 204, 149, 105, 133, 21, 294, 316, 326, 320, 
    303, 300, 297, 293, 305, 300, 294, 308, 300, 316, 314, 318, 319, 329, 
    337, 314, 322, 315, 328, 313, 317, 323, 320, 325, 343, 348, 2, 8, 17, 12, 
    _, 13, 15, 22, 27, 33, 13, 19, 38, 26, 35, 40, 60, 22, 23, 322, 313, 299, 
    322, 308, 330, 319, 336, 312, 348, 332, 342, 334, 305, 348, 5, 356, 358, 
    15, 2, 352, 339, 351, 331, 357, 345, 7, 29, 68, 81, 112, 132, 118, 110, 
    109, 106, 100, 102, 102, 107, 106, 105, 106, 102, 103, _, 98, 94, 97, 87, 
    110, 120, 123, 117, 111, 112, 110, _, 114, 115, 114, 92, 78, 77, 70, 85, 
    94, 102, 111, 105, 96, 96, 82, 85, 92, 82, 70, 73, 61, 63, 64, 63, 67, 
    61, 59, 59, 58, 51, 50, 48, 52, 65, 105, 97, 96, 82, 73, 67, 65, 59, 54, 
    56, 57, 56, 64, 67, 84, 77, 69, 80, 79, 91, 92, 93, 95, 97, 94, _, 94, 
    96, 99, 98, 91, 86, 87, 86, 90, 92, 97, 101, 74, 80, 67, 69, 74, 79, 90, 
    84, 82, 92, 89, 89, 95, 110, 101, 109, 107, 111, 112, 112, 111, 112, 107, 
    99, 88, 91, 101, 98, 110, 120, 135, 120, 114, 120, 118, 116, 105, 109, 
    107, 122, 119, 112, 110, 102, 114, 106, _, 106, 103, 103, 104, 100, 106, 
    116, 130, 112, 112, 114, 110, 118, 118, 113, 105, 107, 100, 100, 98, 88, 
    87, 82, 85, 85, 81, 84, 82, 69, 62, 74, 83, 87, 90, 89, 90, 98, 96, 98, 
    102, 106, 101, 102, 104, 97, 97, 97, 98, 99, 97, 98, 99, 99, 108, 106, 
    107, 103, 103, 109, 111, 112, 110, 110, 108, 109, 111, 114, 114, 118, 
    117, 115, 112, 114, 109, 110, 110, 111, 110, 111, 107, 105, 103, 102, 99, 
    99, 98, 98, 90, 91, 87, 89, 88, 89, 87, 87, 86, 86, 78, 77, 80, 80, 80, 
    80, 81, 80, 80, 79, 80, 83, 78, 85, 88, 91, 96, 88, 89, 90, 91, 83, 75, 
    59, 72, 88, 104, 96, 105, 110, 70, 42, 24, 57, 59, 64, 65, 53, 55, 54, 
    50, 44, 41, 285, 319, 8, 34, 291, 317, 310, 52, 40, 37, 100, 130, 50, 60, 
    186, 247, 335, 360, 45, 49, 41, 54, 31, 50, 54, 318, 304, 293, 234, 20, 
    51, 16, 34, 57, 63, 54, 43, 41, 39, 52, 59, 27, 44, 43, 9, 19, 38, 50, 
    37, 7, 360, 347, 8, 352, 359, 18, 17, 25, 3, 351, 359, 5, 3, 1, 351, 352, 
    360, 344, 342, 356, 5, 341, 356, 340, 349, 333, 359, 331, 333, 335, 320, 
    307, 270, 265, 275, 268, 353, 333, 314, 293, 272, 250, 335, 330, 327, 
    324, 303, 298, 301, 311, 310, 312, 310, 315, 308, 304, 304, 291, 292, 
    296, 308, 287, 289, 277, 254, 240, 119, 149, 201, 106, 108, 115, 109, 
    115, 113, 114, 99, 128, 102, 115, 91, 83, 121, 114, 119, 120, 112, 126, 
    116, 106, 114, 118, 119, 118, 109, 92, 86, 110, 96, 99, 112, 104, 101, 
    81, 68, 63, 60, 64, 64, 71, 70, 78, 77, 79, 102, 109, 106, 116, 103, 89, 
    99, 103, 99, 67, 56, 58, 60, 62, 62, 74, 27, 57, 43, 40, 36, 46, 61, 63, 
    63, 59, 60, 64, 64, 66, 67, 70, 71, 53, 50, 48, 52, 55, 281, 305, 294, 
    316, 14, 346, 343, 355, 13, 1, 5, 356, 344, 331, 339, 335, 350, 351, 319, 
    328, 318, 322, 324, 322, 320, 324, 327, 358, 12, 317, 21, 57, 122, 78, 
    114, 110, 117, 105, 109, 121, 118, 113, 117, 129, 119, 114, 116, 119, 
    117, 106, 108, 109, 110, 110, 98, 105, 102, 103, 101, 99, 98, 91, 94, 96, 
    106, 110, 117, 115, 115, 118, 119, 117, 114, 120, 110, 109, 128, 148, 
    264, 314, 307, 319, 296, 287, 293, 300, 315, 321, 305, 309, 309, 318, 
    330, 334, 342, 335, 342, 3, 310, 336, 300, 324, 305, 326, 286, 309, 307, 
    254, 249, 313, 319, 338, 337, 119, 107, 139, 125, 129, 138, 129, 129, 
    126, 130, 151, 147, 145, 157, 163, 159, 167, 163, 137, 145, 130, 123, 
    121, 120, 118, 123, 117, 121, 124, 120, 120, 126, 136, 131, 117, 117, 
    119, 118, 122, 131, 126, 121, 122, 121, 119, 124, 130, 159, 315, 318, 
    268, 52, 50, 48, 47, 49, 44, 39, 35, 29, 17, 25, 93, 336, 325, 342, 344, 
    325, 335, 336, 326, 308, 306, 298, 298, 311, 306, 314, 285, 300, 276, 
    282, 286, 275, 292, 301, 309, 308, 307, 301, 295, 304, 311, 316, 312, 
    299, 301, 305, 307, 314, 312, 310, 310, 312, 315, 314, 309, 310, _, 314, 
    314, 315, 315, 315, 311, 309, 307, 311, 307, 310, 312, 314, 316, 315, 
    307, 306, 304, 303, 304, 305, 302, 307, 313, 310, 313, 315, 316, 314, 
    316, 313, 316, 312, _, _, 313, 316, 320, 312, 310, 316, 316, 315, 316, 
    315, 317, 318, 318, 315, 315, 309, 314, 311, 304, 306, 323, 315, 319, 
    319, 308, 329, 321, 309, 304, _, 303, 314, 311, _, 305, 300, 289, 291, 
    285, 303, 289, _, 292, 293, 287, 291, _, 307, 301, 294, 287, _, 290, 289, 
    288, 298, _, 301, 300, 299, 310, _, 307, 304, 309, 304, _, 310, 316, 324, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 302, _, 298, 302, 302, 310, 
    314, 311, 305, 298, 292, 290, 275, _, 274, 274, 277, 277, _, 266, 267, 
    279, 271, _, 283, 281, 280, 280, _, 286, 288, 287, 284, _, _, 287, 287, 
    _, _, 291, 288, _, _, _, _, 275, _, 279, _, 278, 281, 274, 244, _, 268, 
    _, 256, 271, _, 286, _, _, 295, _, _, 293, _, 304, 313, 319, 313, 310, _, 
    312, 316, 312, 305, 302, _, _, 311, _, 319, 318, 313, 310, 308, 306, _, 
    _, 315, 307, _, 304, 299, _, 279, 272, 285, 274, _, _, _, _, 228, _, 220, 
    _, 235, 240, _, _, 232, _, 237, _, 126, _, 134, 115, _, 124, 115, 122, 
    131, _, 121, 125, 126, 119, _, 119, 121, _, 123, _, 120, 121, 117, 118, 
    123, 122, 152, 151, 139, 125, 117, 139, 124, _, 117, 116, 90, 125, 338, 
    _, 220, _, _, 42, 303, 62, 24, 327, 308, _, 45, _, 51, 45, _, 50, _, 57, 
    57, 59, 61, _, 75, 62, _, 75, _, 83, 109, 108, _, _, 104, _, 102, 96, _, 
    100, 98, 101, 108, _, 109, 109, 109, 113, _, 117, 117, 114, 111, 107, 
    103, 105, 109, 115, 121, 125, 119, 121, 114, 120, 117, 122, 119, 110, 
    118, 114, 119, 113, 106, 116, 114, _, 125, 133, 122, 119, _, 126, 118, 
    119, 118, _, 119, 120, 108, 112, _, 90, 83, _, 42, _, 321, 347, 109, 329, 
    _, 302, 300, 297, 283, _, 283, 276, 273, 278, _, 273, 270, 268, 273, _, 
    272, 276, 275, 278, _, _, 276, 277, 268, 247, 255, _, 266, 253, 240, 227, 
    224, 235, 241, 264, 273, 295, _, _, 295, 114, _, 137, 130, 121, 126, _, 
    113, 130, 90, 355, _, 47, 27, 16, 313, _, 311, 290, 305, 281, _, 276, 
    292, 308, 326, _, 308, 322, 297, 305, _, 293, 351, 71, 110, 137, 109, 
    126, _, 138, _, 127, 136, 124, 119, _, 128, 130, 124, 119, 128, 116, _, 
    119, 120, 101, 94, 95, 92, 90, 92, 109, 127, 125, 116, 105, 102, _, 106, 
    110, 116, 117, 124, 120, 318, 327, 315, 329, 321, 329, 321, 144, 125, 
    121, 119, 120, 101, 112, 119, 134, 112, 120, 126, 118, 115, 128, 142, 
    191, 304, 32, 131, 315, 321, 313, 325, 82, 266, 183, 4, 260, 255, 268, 
    286, 304, 288, 291, 291, 305, 314, 301, 302, 284, 216, 216, 57, 105, 100, 
    132, 17, 106, 125, 119, 123, 120, 133, 143, 133, 133, 137, 131, 122, 134, 
    133, 133, 127, 124, 116, 120, 118, 118, 115, 112, 119, 122, 116, 115, 
    115, 120, 116, 123, 112, 123, 134, 86, 204, 357, 323, 317, 325, 334, 329, 
    322, 323, 323, 323, 321, 302, 280, 263, 291, 285, 302, 321, 322, 321, 
    299, 304, 321, 304, 317, 314, 301, 294, 317, 288, 314, 310, 276, 0, 130, 
    136, 120, 122, 127, 123, 133, 132, 127, 121, 120, 114, 120, 119, 128, 
    131, 149, 135, 125, 127, 117, 117, 126, 140, 133, 149, 144, 143, 163, _, 
    80, 91, 92, 139, 144, 142, 135, 135, 142, 152, 155, 157, 172, 169, 160, 
    149, 213, 295, 304, 315, 319, 327, 330, 324, 330, 324, 23, 24, 351, 323, 
    319, 314, 317, 311, 317, 289, 323, 319, 324, 155, 126, 128, 116, 112, 
    112, 110, 130, 126, 116, 133, 118, 113, 141, 127, 142, 155, 138, 143, 
    134, 136, 82, 128, 54, 89, 87, 97, 86, 72, 68, 62, 64, 46, 63, 68, 65, 
    60, 57, _, 347, _, _, _, _, _, _, _, _, _, _, 297, _, _, _, _, _, _, _, 
    _, _, 146, 134, 204, 211, 237, 252, 288, 275, 296, 284, 315, 315, 300, 
    306, 312, 322, 318, 329, 332, 315, 277, 292, 279, 273, 255, 229, 234, 
    224, 226, 221, 249, 269, 275, 264, 273, 295, 298, 292, 300, 317, 302, 
    305, 318, 328, 314, 311, 311, 319, 333, 329, 289, 282, 292, 324, 4, 272, 
    203, _, 259, 286, 353, 148, 187, 158, 116, 358, 315, 333, 125, 171, 250, 
    323, 290, 339, 304, 306, _, 315, 327, 189, 161, 275, 311, 149, 259, 293, 
    325, 323, 330, 335, 328, 294, 235, 264, 270, 230, 268, 245, 242, 275, 
    291, 211, 231, 255, 245, 281, 298, 152, 301, 295, 322, 339, 294, 46, 355, 
    322, 326, 4, 317, 302, 333, 332, 342, 316, 312, 319, 326, 323, 328, 323, 
    350, 352, 346, 345, 132, 146, 273, 258, 158, 171, _, 234, 197, 317, 65, 
    47, 79, 355, 316, 333, 320, 310, _, 347, 6, 56, 305, 57, 263, 202, 279, 
    227, 267, 63, 297, 312, 58, 57, 59, 54, 55, 58, 57, 58, 55, 52, 62, 56, 
    60, 49, 53, 54, 56, 52, 42, 49, 48, 52, 48, 54, 265, 273, 50, 50, 50, 47, 
    47, 329, 214, 304, 46, 323, 48, 46, 57, 52, 54, 52, 57, 56, 57, 51, 47, 
    291, 249, 351, 294, 293, 254, 196, 323, 327, 328, 339, 200, 282, 274, 
    311, 305, 319, 216, 327, 311, 267, 250, 281, 307, 281, 257, 289, 236, 
    272, 259, 285, 348, 284, 318, 353, 196, 353, 46, 237, 289, 125, 250, 73, 
    77, 39, 317, 203, 291, 333, 276, 64, 68, 76, 84, 88, 87, 82, 85, 75, 79, 
    76, 70, 60, 61, 61, 61, 328, 303, 352, 338, 163, 320, 299, 309, 301, 18, 
    110, 142, 304, 308, 332, 348, 310, 319, 318, 313, _, 304, 298, 305, 318, 
    317, 321, 324, 322, 325, 324, 324, 354, 356, 312, 163, 151, 276, 310, 
    276, 113, 334, 291, 231, 223, 305, 287, 283, 290, 265, 280, 335, 271, 
    307, 264, 329, 347, 279, 254, 301, 303, 315, 46, 52, 62, 55, 51, 54, 48, 
    343, 42, 54, 55, 54, 49, 53, 56, 53, 55, 56, 54, 53, 54, 311, 99, _, 77, 
    83, 77, 74, 70, 77, 66, 71, 85, 87, 100, 106, 104, _, 106, 112, 113, 112, 
    110, 112, 112, 110, 113, 113, 100, 80, 73, 67, 66, 65, 61, 308, 335, 304, 
    1, 311, 330, 345, 329, 321, 309, 297, 301, 303, 307, 346, 294, 298, 283, 
    275, 277, 283, 294, 292, 279, 274, 284, 289, 298, 318, 311, 307, 310, 
    312, 313, 312, 304, 296, 302, 308, 306, 306, 309, 309, 322, 312, 331, 
    320, _, 291, 314, 302, 324, 326, 303, _, 322, 304, 320, 327, 320, 328, 
    335, 320, 306, 291, 281, 308, 286, 241, 160, 163, 144, 149, 158, 147, 
    145, 144, 172, 332, 319, 143, 337, 178, 108, 130, 105, 112, 103, 88, 164, 
    301, 313, 257, 318, 352, 352, 296, 350, 330, 328, 326, 329, 319, 327, 
    333, 327, 318, 320, 329, 319, 326, 331, 324, 326, 312, 309, 308, 324, 
    323, 326, 323, 315, 317, 302, 303, 315, 316, 320, 328, 331, 322, 324, 
    329, 325, 327, 324, 325, 333, 335, 335, 336, 338, 332, 315, 316, 316, 
    322, 336, 341, 326, 322, 321, 327, 323, 344, 266, 234, 188, 152, 184, 
    178, 182, 176, 168, 158, 241, 115, 127, 153, 106, 131, 138, 97, 103, 128, 
    112, 136, 134, 130, 145, 137, 139, 140, 140, 115, 140, 135, 142, 128, 
    115, 127, 118, 146, 131, 130, 126, 143, 197, 166, 237, 279, 275, 254, 
    210, 189, 100, 195, 274, 332, 302, 289, 307, 315, 301, 303, 290, 273, 
    281, 279, 270, 247, 226, 248, 231, 167, 133, 179, 91, 322, 307, 336, 317, 
    329, 322, 302, 324, 323, 242, 193, 166, 123, 203, 281, 294, 313, 318, 
    333, 313, 3, 316, 316, 315, 329, 334, 340, 325, 328, 319, _, 332, 321, 
    341, 327, 305, 321, 298, 331, 328, 325, 322, 320, 310, 308, 312, 322, 
    320, 297, 300, 302, 344, 335, 317, 327, 329, 326, 335, 343, 333, 329, 
    329, 317, _, 307, 304, 299, 301, 297, 302, 307, 240, 310, 295, 331, 331, 
    322, 334, 337, 333, 287, 240, 145, 92, _, 128, 120, 303, _, 323, 332, 
    314, 322, 310, 329, 296, 287, 296, 299, 291, 252, 251, _, 279, 249, 254, 
    239, 237, 238, 229, 193, 168, 164, 118, 156, 112, 123, 125, 128, 144, 
    140, 135, 155, 148, 140, 137, 130, 100, 134, 127, 106, 77, 142, 142, 143, 
    147, 126, 242, 161, 134, 141, 145, 180, 151, 177, 173, 151, 168, 189, 
    165, 173, 153, 124, 150, 123, 46, 350, 353, 309, 287, 319, 355, 310, 337, 
    322, 332, 335, 313, 312, 291, 312, 317, 316, 348, 341, 329, 337, 324, 
    323, 278, 173, 111, 82, 95, 120, 117, 106, 108, 113, 101, 89, 97, 101, 
    102, 99, 87, 123, 114, 113, 111, 111, 113, 116, 113, 111, 114, 118, 115, 
    114, 105, 106, 104, 99, 92, 96, 99, 98, 91, 98, 91, 109, 132, 122, 145, 
    313, 300, 296, 300, 300, 2, 4, 317, 343, 222, 235, 254, 281, 258, 340, 
    314, 359, 283, 327, 330, 337, 311, 320, 359, 329, 329, 327, 328, 334, 
    329, 332, 334, 333, 331, 338, 329, 332, 335, 348, 348, 321, 338, 334, 
    327, 346, 335, 334, 331, 330, 325, 334, 341, 330, 330, 326, 327, 316, 
    325, 310, 306, 326, 322, 296, 286, 282, 289, 290, 292, 292, 292, 302, 
    292, 298, 303, 332, 314, 286, 284, 294, 285, 289, 292, 298, 280, 254, 
    218, 173, 143, 142, 172, 153, 141, 149, 136, 147, 157, 163, 142, 132, 
    135, 121, 107, 71, 26, 340, 359, 323, 334, 322, 319, 316, 233, 179, 249, 
    315, 325, 265, 297, 322, 316, 315, 323, 313, 288, 3, 53, 99, 99, 114, 
    117, 121, 119, 121, 124, 138, 151, 150, 152, 147, 141, 157, 152, 148, 
    142, 178, 211, 219, 259, 292, 310, 290, 316, 284, 291, 290, 267, 269, 
    262, 282, 237, 229, 220, 237, 223, 209, 214, 199, 183, 178, 174, 172, 
    117, 124, 134, 120, 117, 106, 135, 110, 61, 102, 189, 164, 176, 165, 164, 
    161, 159, 173, 187, 202, 162, 97, 117, 127, 141, 134, 118, 118, 107, 133, 
    115, 116, 111, 110, 99, 115, 111, 112, 114, 116, 116, 114, 115, 113, 104, 
    105, 108, 102, 101, 70, 340, 330, 339, 323, 322, 323, 335, 317, 323, 319, 
    312, 298, 308, 330, 151, 137, 100, 115, 118, 112, 130, 120, 115, 119, 
    125, 126, 113, 120, 97, 105, 67, 322, 337, 312, 309, 92, 168, 111, 146, 
    84, 108, 105, 99, 125, 98, 112, 115, 115, 115, 102, 108, 119, 137, 120, 
    144, 117, 358, 327, 333, 358, 167, 166, 54, 55, 56, 54, 60, 76, 97, 94, 
    96, 100, 105, 108, 114, 119, 122, 128, 120, 139, 176, 41, 268, 286, 308, 
    268, 275, 283, 275, 279, 292, 303, 295, 292, 287, 282, 302, 299, 291, 
    291, 301, 308, 292, 289, 302, 300, 292, 321, 323, 322, 1, 94, 114, 109, 
    115, 113, 131, 200, 268, 277, 329, 314, 296, 293, 290, 291, 280, 275, 
    276, 278, 282, 275, 281, 281, 283, 285, 278, 287, 280, 280, 281, 280, 
    282, 282, 283, 285, 289, 288, 288, 287, 283, 275, 256, 237, 203, 205, 
    207, 201, 198, 200, 192, 196, 238, 287, 274, 301, 290, 300, 283, 295, 
    307, 290, 295, 294, 309, 318, 327, 323, 327, 333, 330, 318, 318, 319, 
    312, 311, 307, 297, 316, 318, 310, 315, 317, 317, 312, 314, 320, 322, 
    326, 344, 352, 356, 339, 347, 336, 342, 337, 336, 330, 328, 326, 326, 
    324, 321, 335, 325, 324, _, 318, 310, 313, 315, 312, 314, 309, 309, 309, 
    305, 312, 314, 310, 306, 309, 302, 300, 293, 290, 292, 290, 296, _, 302, 
    315, 316, 313, 311, 307, 309, 304, 303, 304, 302, 298, 294, 295, 287, 
    290, 289, 285, 267, 256, 232, 216, 219, 230, 231, 246, 256, 257, 262, 
    258, 262, 264, 272, 275, 280, 296, 303, 332, 333, 329, 337, 342, 327, 
    336, 347, 339, 347, 336, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, 276, 282, 242, 266, 213, 221, _, 200, 180, 199, 181, 174, 170, 155, 
    128, 146, 138, 116, 98, 82, 79, 65, 52, _, 249, 288, 345, 328, 332, 332, 
    61, 336, 137, 115, 118, 100, 115, 119, 112, 102, 86, 71, _, 321, _, 335, 
    328, 317, 315, 318, 319, 323, 311, 318, 316, _, _, 329, _, 330, 328, 307, 
    281, 280, 274, 272, 262, 246, 242, 242, 244, 246, 230, 210, 200, 206, 
    200, 184, _, 153, 116, 120, 108, 126, 155, 153, 187, 185, 243, 6, 95, 12, 
    195, 24, 19, 23, 30, 32, 46, 54, 53, _, 58, 54, 58, 53, 56, 56, 49, 52, 
    48, 52, 50, 46, 32, 3, 1, 304, 335, 347, 344, 340, 335, 336, 341, 333, 
    327, 324, _, 317, 325, 338, 322, 314, 301, 316, 319, 312, 317, 326, 309, 
    348, 345, 348, 8, 360, 0, 80, 96, _, 144, 145, 151, 143, 134, 142, 142, 
    137, 153, 144, 145, 148, 153, 146, 152, 149, 142, 127, 148, 145, 152, 
    148, 142, 140, 122, _, 110, 112, 114, 120, 115, 119, 113, 96, 99, 101, 
    108, 112, 109, 116, 127, 209, 239, 329, 291, 324, 324, 296, 313, 329, 
    313, 317, 321, 313, 333, 356, 343, 335, 323, 314, 320, 325, 345, 310, 
    335, 317, 99, 99, 42, 182, 340, 137, 189, 17, 6, 114, 78, 60, 18, 26, 
    277, 314, 358, 321, 340, 356, 352, 339, 331, 330, 339, 344, 344, 346, 
    350, 344, 340, 330, 339, 360, 339, 348, 352, 360, 321, 326, 324, 341, 
    309, 309, 306, 324, 303, 300, 15, 331, 329, 327, 323, 324, 122, 313, 311, 
    332, 310, 332, 318, 332, 345, 341, 350, 301, 327, 351, 50, 11, 185, _, 
    297, 55, 57, 60, 267, 68, 278, 332, 128, 244, 309, 316, 270, 327, 318, 
    330, 334, 330, 335, 329, 328, 316, 312, 305, 314, 324, 319, 317, 311, 
    320, 317, 316, 319, 315, 317, 330, 324, 315, 320, 309, 306, 353, 9, 95, 
    96, 103, 117, 118, 110, 114, 129, 122, 108, 110, 115, 119, 113, 113, 109, 
    104, 100, 107, 108, 118, 111, 117, 128, 110, 125, 115, 131, 134, 128, 
    130, 123, 120, 114, 129, 126, 123, 120, 117, 248, 326, 333, 323, 301, 
    293, 295, 300, 331, 318, 306, 304, 300, 298, 310, 314, 307, 301, 303, 
    303, 296, 298, 295, 300, 306, 319, 323, 324, 325, 342, 349, 2, 19, 122, 
    103, 168, 151, 127, 130, 112, 138, _, 130, 124, 128, 131, 128, 134, 130, 
    129, 120, 122, 115, 114, 112, 126, 121, 120, 121, 119, 121, 121, 122, 
    118, 119, 119, 121, 130, _, 127, 122, 125, 123, 118, 110, 108, 111, 109, 
    123, 123, 119, 115, 119, 118, 119, 123, 128, 110, 106, 112, 121, 119, 
    120, 130, 131, 138, 145, 157, 178, 189, 201, 189, 205, 234, 242, 270, 
    297, 297, 322, 321, 318, 320, 324, 321, 320, 309, 299, 292, 296, 289, 
    292, 289, 299, 299, 305, 262, 296, 313, 306, 302, 318, 19, 98, 110, 116, 
    104, 104, 105, 106, 107, 101, 96, 101, 88, 87, 89, 108, 116, 114, 110, 
    105, 102, 102, 107, 111, 139, 145, 145, 181, 213, 209, 222, 262, 195, 
    268, 294, 303, 312, 293, 334, 315, 295, 334, 153, 82, 98, 106, 98, 122, 
    144, 160, 204, 281, 307, 291, 283, 290, 291, 290, 292, 301, 320, 332, 
    343, 67, 143, 157, 141, 122, 113, 121, 126, 131, 129, 123, 114, 101, 122, 
    94, 97, 327, 328, 345, 22, 22, 22, 356, 326, 122, 38, 52, 53, 51, 53, 60, 
    60, 75, 79, 68, 72, 70, 69, 72, 65, 66, 243, 276, 317, 335, 303, 308, 
    347, 14, 156, 2, 330, 332, _, 300, 277, 322, 337, 239, 277, _, 332, 87, 
    116, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 112, 109, 110, 113, 135, 115, 
    118, 111, 123, 122, 107, 113, 114, 117, 120, 119, 121, 115, 125, 114, 
    130, 128, 137, 131, 138, 166, 138, 137, 167, 100, 347, _, 348, 329, 6, 
    356, 33, 2, 351, 326, 323, 331, 333, 335, 339, 343, 345, 345, 7, _, 13, 
    22, 34, 31, 28, 31, 29, 34, 27, 30, 27, 23, 19, 30, 36, 39, 43, 45, 49, 
    60, 66, 72, 84, 96, 93, 100, 100, 99, 93, 91, 106, 103, 105, 103, 101, 
    100, 90, 65, 70, 66, 65, 67, 57, 76, 86, 92, 90, 82, 78, 81, 79, 77, 77, 
    80, 83, 82, 74, 61, 70, 72, 73, 70, 69, 69, 71, 70, 72, 75, 76, 71, 72, 
    73, 70, 73, 74, 84, 83, 80, 79, 69, 72, 73, 72, 69, 71, 83, 79, 75, 281, 
    300, 300, 302, 306, 303, _, 295, 302, 299, 298, 296, 292, 287, 286, 276, 
    274, 283, 281, 290, 289, 289, 292, 289, 284, 280, 267, 226, 229, 192, 
    193, 175, 151, 154, 156, 157, 152, 146, 143, 130, 124, 118, 118, 112, 
    114, 129, 112, 109, 110, 116, 124, 110, 111, 115, 120, _, 114, 117, 117, 
    110, 119, 116, 22, 301, 322, 319, 316, 275, 287, 302, 302, 308, 310, 309, 
    308, 305, 324, 329, 320, 318, 316, 308, 345, 86, 108, 111, 115, 119, 141, 
    132, 125, 123, 125, 117, 113, 115, 104, 121, 118, 122, 112, 116, 112, 
    114, 131, 196, 194, 217, 311, 12, 338, 314, 288, 293, 275, 275, 275, 280, 
    276, 279, 280, 282, 280, 288, 284, 281, 281, _, 293, 297, 294, 297, 294, 
    291, 307, 204, 192, 199, 222, 247, 264, 291, 288, 279, 276, 290, 291, 
    283, 247, 242, 46, 99, 98, 81, 84, 100, 104, 97, 92, 108, 110, 113, 121, 
    120, 109, 111, 89, 97, 112, 109, 112, 106, 108, 103, 107, 131, 113, 113, 
    124, 114, 113, 110, 319, 333, 313, 331, 309, 314, 319, 305, 302, 290, 
    286, 292, 294, 285, 299, 53, 64, 81, 137, 91, 61, 57, 55, 52, 52, 51, 14, 
    50, 294, 319, 339, 331, 335, 331, 311, 290, 277, 292, 312, 311, 311, 306, 
    308, 314, 312, 303, 301, 312, 310, 308, 305, 306, 304, 317, 326, 330, 
    341, 348, 356, 2, 8, 356, 52, _, 283, 276, 224, 79, 141, 202, 217, 211, 
    172, 164, 167, 175, 168, 152, 107, 107, 109, 97, 93, 101, 91, 94, 96, 
    102, 120, 111, 120, 119, 118, 112, 116, 112, 113, 116, 132, 109, 95, 110, 
    115, 121, 282, 328, 327, 360, 314, 180, 87, 125, 80, 69, 326, 313, 303, 
    292, 265, 252, 249, 261, 257, 258, 265, 269, 292, 285, 290, 288, 290, 
    288, 294, 289, 290, 295, 293, 295, 291, 288, 289, 294, 300, 301, 311, 
    304, 310, 293, 298, 299, 298, 295, 294, 308, 357, 110, 223, 232, 239, 
    218, 213, 213, 209, 217, 216, 162, 147, 115, 117, 106, 103, 95, 101, 93, 
    85, 115, 121, _, 134, 119, 114, 111, 104, 142, 0, 0, 0, 0, 0, 0, 0, 0, 
    141, 122, 135, 127, 122, 121, 122, 121, 113, 120, 104, 123, 117, 108, 
    130, 105, 129, 119, 127, 121, 133, 125, 136, 129, 115, _, 117, 121, 120, 
    123, 127, 112, 115, 111, 110, 109, 121, 116, 114, 104, 111, 113, 100, 
    117, 113, 109, 104, 100, 122, 111, 114, 115, 121, 121, _, _, _, _, 140, 
    188, 175, 166, 167, 159, 190, 188, 213, 194, 204, 157, 113, 290, 334, 
    315, 353, 296, 309, 307, 306, 301, 303, 310, 311, 309, 307, 309, 306, 
    309, 306, 307, 306, 307, 305, 305, 305, 306, 295, _, 303, 295, 320, 331, 
    19, 71, 68, 77, 67, 72, 99, 108, 102, 104, 111, 107, 105, 100, 91, 90, 
    93, 97, 95, 91, 72, 95, 122, 114, 114, 116, 42, 351, 150, 336, 117, 124, 
    116, 125, 122, 127, 123, 123, 123, 125, 137, 100, 130, 125, 97, 45, 112, 
    126, 122, 112, 129, 131, 131, 113, 106, 126, 113, 117, 111, 83, 78, 73, 
    80, 97, 87, 86, 85, 82, 79, 84, 89, 82, 77, 71, 71, 67, 65, 67, 61, 62, 
    61, 59, 61, 59, 62, 62, 72, 106, 129, 119, 118, 120, 96, 91, 102, 114, 
    108, 121, 108, 117, 113, 121, 109, 111, 121, 120, 106, 105, 107, 102, 99, 
    _, 100, 106, 109, 108, 94, 97, 92, 88, 81, 72, 74, 65, 57, 49, 58, 52, 
    54, 51, 49, 55, 56, 53, 47, 50, 52, 52, 49, 36, 33, 29, 32, 42, 47, 58, 
    60, 62, 50, 51, 51, 49, 49, 52, 43, 56, 58, 48, 49, 59, 55, 50, _, 64, 
    49, 46, 45, 44, 317, 358, 326, 335, 16, 48, 45, 40, 44, 323, 333, 23, 21, 
    28, 30, 34, 29, 37, 15, 0, 49, 14, 18, 42, 29, 33, 24, 18, 39, 38, 30, 
    12, 79, 49, 9, 348, 14, 45, _, 66, 61, 55, 47, 66, 325, 65, 101, 97, 29, 
    42, 35, 47, 36, 41, 48, 51, 51, 75, 80, 75, 71, 74, 77, 86, 97, 95, 102, 
    105, 104, 118, 114, 116, 115, 113, 112, 122, 132, 126, 123, 122, 109, 
    103, 103, 109, 115, 103, 103, 114, 131, 118, 116, 119, 149, 148, 126, 95, 
    _, 109, 114, 121, 128, 136, 128, 121, 129, 125, 129, 130, 136, 123, 118, 
    135, 160, 171, 157, 165, 176, 162, 159, 157, 154, 152, 146, 146, 142, 
    144, 165, 159, 156, 152, 142, 129, 150, 143, 147, 113, _, 114, 120, 154, 
    154, 137, 126, 127, 180, 181, 198, 208, 360, 309, 312, 324, 328, 334, 
    334, 338, 340, 343, 348, 360, 7, 22, 29, 21, 32, 53, 65, 60, 108, 100, 
    118, 128, 154, 144, 147, 156, 161, 158, 148, 159, 161, 162, 159, 158, 
    156, 155, 148, 148, 152, 155, 151, 154, 149, 140, 125, 120, _, 121, 118, 
    135, 135, 131, 152, 138, 143, 151, 158, 162, 172, 167, 175, 168, 166, 
    162, 167, 165, 171, 166, 166, 176, 183, 190, 201, 209, 266, 279, 268, 
    269, 249, 258, 239, 262, 269, 268, 263, 275, 263, 278, 276, 278, 277, 
    275, 277, 276, 280, 283, 285, 286, 286, 285, 291, 283, 293, 289, 288, 
    294, 304, 300, 299, 294, 288, 291, 282, 281, 288, 290, 281, 282, 290, 
    291, 292, 304, 26, 180, 97, 4, 245, 261, 247, 253, 227, 28, 116, 243, 
    347, 81, 111, 124, 108, 111, 131, 128, 145, 94, 123, 102, 104, 104, 110, 
    115, 114, 111, 109, 107, 108, 111, 115, 123, 123, 113, 114, 117, 117, 
    117, 113, 114, 113, 112, 114, 114, 112, 109, 110, 109, 104, 110, 110, 
    105, 101, 100, 93, 90, 98, 96, 99, 97, 98, 102, 95, 91, 89, 87, 83, _, 
    84, 91, 98, 103, 116, 105, 95, 106, 103, 109, 113, 119, 120, 132, 143, 
    144, 140, 138, 131, 136, 138, 120, 122, 115, 118, 122, 129, 121, 119, 
    123, 113, 118, 121, 121, 120, 117, 116, 113, 115, 113, 116, 121, 126, 
    126, 133, 139, 137, 146, 149, 146, 149, 142, 143, 144, 139, 144, 148, 
    150, 140, 152, 153, 142, 139, 130, 127, 126, 119, 117, 114, 108, 108, 99, 
    101, 96, 101, 98, 100, 106, 104, 108, 107, 107, 106, 107, 104, 102, 100, 
    110, 111, 110, 118, 125, 127, 130, 134, 142, 148, 150, 129, 139, 118, 
    118, 107, 133, 129, 134, 130, 127, 131, 130, 126, 128, 125, 125, 127, 
    125, 124, 128, 135, 132, 122, 122, 118, 115, _, 99, 96, 105, 110, 110, 
    121, 114, 115, 106, 103, 87, 90, 107, 97, 97, 102, 100, 93, 100, _, 91, 
    72, 87, 86, 84, 76, 66, 50, 50, 60, 64, 58, 62, 59, 71, 57, 56, 54, 47, 
    317, 54, 60, 62, 61, 56, 55, 53, 60, 60, 75, 73, 55, 49, 41, 45, 40, 50, 
    49, 52, 56, 48, _, 286, 45, 26, 22, 92, 78, 69, 56, 67, _, 19, 12, 16, 
    23, 344, 58, 75, 61, 35, 52, 11, 10, 347, 14, 5, 10, 3, 19, 15, 23, 38, 
    26, 330, 31, 59, 43, 54, 62, 55, 42, 52, 49, 55, 56, 53, 52, 56, 52, 54, 
    55, 52, 55, 62, 54, 45, 38, 60, 37, 48, 49, 47, 43, 58, 51, 54, 52, 51, 
    33, 40, 74, 246, 10, 307, 275, 326, 4, 51, 51, 43, 34, 60, _, 58, 19, 58, 
    59, 93, 87, 74, 77, 56, 80, 19, 12, 17, 17, 360, 352, 324, _, 344, _, 
    348, 355, 349, 346, 343, 337, 18, 18, 3, 358, 357, 355, 2, 12, 10, 2, 
    355, 352, 345, 352, 342, 14, 348, 353, 346, 340, 8, 4, 16, 5, 35, 32, 40, 
    29, 40, 32, 26, 24, 12, 21, 19, 40, 44, 40, 30, 31, 28, 18, 19, 14, 24, 
    23, 21, 13, 23, 22, 23, 21, 6, 331, 325, 321, 334, 322, 335, 15, 33, 38, 
    53, 63, 56, 57, 51, 55, 53, 55, 66, 49, 45, 50, 93, 116, 87, 92, 92, 95, 
    85, 81, _, 71, 81, 71, 81, 51, 57, 64, 67, 58, 62, 69, 65, 61, 73, 55, 
    38, 37, 36, 38, 28, 38, 62, 83, 76, 70, 69, 48, 48, 44, 39, 25, 43, 38, 
    35, 40, 37, 45, 47, 39, 28, 46, 32, 29, 39, 40, 35, 41, 35, 30, 39, 46, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 213, 224, 212, 213, 192, 213, 232, 254, 253, 271, 231, 228, 218, 
    209, 212, 208, 240, 241, 241, 229, 222, 231, 230, 223, 225, 205, 197, 
    204, 231, 204, 216, 208, 211, 243, 257, 259, 260, 246, 282, 299, 338, 
    329, 337, 351, 351, 1, 2, 23, 5, 13, 22, 29, 41, 47, 47, 50, 50, 51, 52, 
    52, 48, 49, 39, 42, 16, 355, 341, 335, 326, 322, 327, 320, 287, 296, 303, 
    296, 312, 296, 297, 298, 283, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 161, 158, 158, 153, 160, 163, 159, 153, 154, 153, 
    149, 150, 152, 142, 143, 140, 143, 155, 174, 187, 273, 301, 279, 317, _, 
    313, 321, 321, 334, 336, 5, 53, 346, 104, 69, 112, 354, 9, 271, 34, 58, 
    59, 62, 62, 60, 65, 60, _, 52, 48, 46, 50, 56, 61, 54, 55, 52, 43, 49, 
    54, 60, 64, 67, 76, 77, 109, 118, 117, 121, 120, 116, 117, 115, 117, 124, 
    126, 121, 114, 110, 110, 112, 106, 110, 113, 116, 120, 118, 119, 109, 
    109, 114, 113, 112, 118, 116, 115, _, 115, 116, 114, 113, 118, 129, 123, 
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 119, 109, 
    102, 96, 91, 86, 93, 100, 102, 121, 141, 171, 244, 247, 239, 242, 235, 
    242, 239, 326, 255, 316, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 
    101, 105, 102, 95, 109, 123, 135, 133, 142, 141, 145, 137, 143, 138, 130, 
    _, 135, 135, 135, 139, 132, 127, 146, 161, 148, 165, 120, _, 115, _, 108, 
    123, 116, 114, 108, 105, 70, 60, 44, 44, 50, 51, 59, 71, 72, 72, 88, 89, 
    89, 90, 89, 82, 80, 84, 75, 77, 74, 70, 64, 80, 89, 125, 112, 121, 108, 
    97, 89, 99, 101, 81, 83, 81, 86, 281, 119, 75, 331, 59, 46, 49, 60, 49, 
    63, 54, 42, 36, 57, _, 115, _, 91, 103, 104, 90, 97, 87, 59, 43, 66, _, 
    76, _, 69, 89, 83, 96, 89, 70, 70, 83, 82, 75, 73, 78, 69, 65, 72, 76, 
    68, 58, 49, 54, 55, 57, 59, 57, 56, 75, 76, 78, 74, 70, 74, 80, 68, 62, 
    59, 62, 59, 54, 45, 34, 27, 23, 24, 21, 26, 23, 50, 45, 48, 51, 53, 59, 
    55, 63, 64, 337, 82, 70, 64, 53, 60, 56, 67, 56, 58, 66, 66, 62, 54, 66, 
    89, 92, 96, 102, 100, 96, 101, 102, 97, 92, 93, 99, 98, 98, 93, 91, 96, 
    90, 93, 96, 91, 86, 91, 89, 82, 86, 82, 79, 68, 70, 66, 66, 70, 75, 59, 
    68, 74, 72, 62, 60, 68, 70, 68, 70, 59, 62, 56, 61, 65, 67, 62, 67, 80, 
    75, 66, 56, 59, 52, 60, _, 40, _, 33, 21, 29, 30, 28, 32, 38, 41, 30, 27, 
    18, _, 28, 26, 14, 9, 35, 26, 21, 10, 16, 39, 336, 18, 27, 10, 31, 29, 
    29, _, 23, 42, 20, 44, 46, 62, 68, 76, 64, 73, 69, 73, 60, _, 74, 87, 83, 
    85, 82, 75, 79, 79, 84, 89, 88, 91, 101, 105, 103, 98, 116, 118, 135, 
    118, 116, 119, 119, 121, 132, 131, 131, 136, 140, 141, 138, 137, 146, 
    149, 153, 150, 153, 153, 158, _, 153, _, 164, 172, 168, 162, 173, 179, 
    183, 175, 178, 181, 194, 202, 207, 208, 208, 215, 211, 215, 212, 212, 
    206, 199, 221, 204, 213, 192, 199, 191, 209, 208, 224, 250, 251, 248, 3, 
    28, 39, 55, 67, _, 62, 62, 91, 84, 122, 152, 145, 140, 133, 131, 127, 
    145, 130, _, 111, 116, 107, 89, 62, 24, 22, 351, 327, 334, 338, 335, 337, 
    338, 339, _, 5, 3, 5, 6, 18, 4, 11, 10, 18, 11, 20, 10, 27, 22, 4, 357, 
    356, 356, 357, 355, 330, 321, 317, 314, 307, 316, 321, 305, 313, 298, 
    309, 305, 314, 311, 321, 282, 302, 311, 308, 9, 344, _, 317, 322, 1, 334, 
    301, 291, 289, 351, 335, 330, 325, 311, 306, 291, 313, 322, 338, _, _, 
    325, 353, 336, 337, 352, 336, 341, 350, 333, 346, 341, 349, 343, 330, 
    336, 336, 330, 335, 324, 332, 324, 315, 314, 315, 329, 328, 324, 321, 
    312, 313, 305, 302, 296, 298, 297, 295, 294, 289, 289, 283, 281, 279, 
    275, 266, 264, 261, 253, 249, 242, 249, 243, 228, 184, 268, 2, 8, 266, 
    290, 278, 295, 298, 354, 6, 5, 13, 6, 15, 4, 4, 13, 5, 20, 24, 14, 40, 
    45, 60, 60, 40, 43, 28, 54, 48, 45, 42, 47, 32, 46, 29, 44, 45, 56, 55, 
    70, 356, 108, 155, 206, 240, 213, 319, 312, 307, 286, 289, 285, 291, 293, 
    283, 292, 293, 273, 270, 273, 297, 298, 333, 19, 29, 33, 49, 44, 38, 35, 
    36, 39, 46, 44, 47, 39, 33, 23, 29, 8, 23, 17, 24, 38, 30, 35, 30, 35, _, 
    46, 41, 28, 29, 357, 358, 350, 340, 337, 335, 300, 310, 306, 277, 268, 
    265, 268, 270, 245, 291, 284, 285, 275, 281, 294, 247, 198, 166, 180, 
    151, 142, 142, 134, 131, 134, 133, 130, 136, 138, 140, 137, 132, 132, 
    132, 129, 135, 139, 149, 182, 186, 193, 173, 171, _, 166, 153, 159, 159, 
    162, 182, 179, 164, 171, 205, 215, 217, 244, 246, 269, 261, 267, 266, 
    263, 269, 263, 267, 256, 268, 266, 253, 234, 229, 230, 232, 229, 236, 
    229, 231, 263, 253, 275, 268, 278, 283, 285, 290, 287, 284, 268, 238, 
    225, 209, 222, 210, 235, 184, 176, 214, 224, 235, 233, 270, 265, 265, 
    259, 253, 255, 242, 238, 251, 239, 245, 251, 258, 261, 266, 261, 281, 
    277, 291, 289, 301, 308, 312, 309, 289, 275, 322, 315, 307, 295, 322, 
    312, 310, 319, 314, 321, 319, 311, 360, 13, 13, 20, 14, 16, 11, 11, 18, 
    21, 16, 8, 13, 4, 17, 33, 33, 35, 47, 47, 62, 41, 358, 312, 319, 324, 
    328, 317, 312, 1, 14, 30, 47, 80, 73, 75, 85, 90, 85, 82, 86, 95, 108, 
    137, 141, 150, 145, 151, 159, 154, 163, 160, 150, 152, 160, 162, 155, 
    163, 165, 163, 182, 169, 176, 178, 188, 188, 192, 185, _, _, 161, 161, 
    156, 160, 174, 175, 174, 170, 170, 172, 178, 178, 171, 186, 284, 276, 
    276, 271, 280, 281, 290, 293, 299, 313, 307, 311, 317, 322, 326, 333, 
    323, 336, 356, 349, 351, 350, 344, 343, 350, 349, 345, 346, 339, 343, 
    339, 321, 328, 314, 319, 319, 315, _, 311, 309, 298, 305, 306, 306, 305, 
    301, 294, 296, 299, 297, 298, 288, 292, 285, 291, 293, 284, 289, 292, 
    290, 284, 285, 289, 281, 284, 286, 292, 290, 290, 294, 297, 307, 300, 
    302, 318, 322, 310, 312, 300, 297, 293, 293, 316, 299, 287, 309, 322, 
    297, 278, 280, 277, 273, 278, 273, 278, 280, 280, 286, 296, 296, 280, 
    294, 293, 281, 282, 282, 297, 288, 283, 289, _, 288, 290, 302, 293, 286, 
    288, 302, 296, 303, 300, 309, 296, 298, 310, 305, 294, 297, 300, 308, 
    307, 314, 303, 303, 294, 296, 297, 294, 292, 293, 342, 36, 49, 20, 50, 
    56, 48, 70, 337, 322, 319, 306, 300, 335, 345, 13, 5, 327, 339, 335, 326, 
    320, 302, 298, 298, 302, 297, 302, 300, 298, 289, 292, 291, 291, 287, 
    292, 289, 300, 294, 306, 298, 295, 295, 295, 300, 301, 294, 290, 313, 
    311, 314, 295, 292, 268, 244, 295, 178, 142, 134, 123, 154, 159, 158, 
    151, 148, 145, 151, 157, 152, 151, 150, 155, 161, 162, 152, 146, 151, 
    147, 144, 142, 142, 140, 140, 139, 142, 143, 145, 144, 146, 139, 137, 
    142, 141, 142, 143, 140, 142, 138, 134, 132, 132, 130, 131, 131, 137, 
    139, 138, 139, 139, 140, 138, 144, 146, 139, _, 100, 91, 336, 359, 354, 
    345, 344, 345, 349, 349, 28, 52, 85, 68, 101, 110, 123, 131, _, 151, 148, 
    _, 143, 153, 151, 144, 116, 104, 104, 109, 110, 117, 112, 113, 122, 138, 
    325, 315, 315, 323, 306, 333, 336, 235, 106, 69, 86, 13, 330, 331, 137, 
    96, 78, 94, 110, 112, 123, 109, 118, 142, 127, 111, 118, 108, 127, 113, 
    147, 121, 136, 137, 106, 160, 198, 123, 90, 113, 207, 243, 86, 239, 246, 
    279, 286, 312, 293, 291, 290, 292, 295, 300, _, 295, 285, 296, 292, 300, 
    304, 293, 288, 328, 38, 115, 112, 113, 120, 128, 121, 112, 108, 114, 110, 
    110, 118, 100, 127, 93, 97, 114, 107, 116, 120, 131, 110, 141, 279, 152, 
    246, 240, 243, 269, 281, 278, 293, 294, 292, 309, 286, 311, 296, 323, 
    196, 114, 84, 109, 113, 103, 102, 132, 128, 112, 142, 120, 126, 126, 134, 
    136, 134, 155, 142, 158, 179, 195, 192, 213, 206, 178, 182, 90, 143, 105, 
    205, 135, 125, 119, 129, 119, 131, 195, 206, 145, 185, 167, 165, 111, 
    114, 186, 75, 119, 106, 127, 133, 105, 100, 342, 314, 16, 4, 339, 338, 
    334, 332, 335, 340, 330, 325, 325, 324, 337, 329, 329, 335, 339, 324, 
    319, 331, 328, 321, 335, 330, 318, 319, 322, 317, 315, _, 318, 315, 318, 
    302, 298, 314, 304, 312, 308, 306, 301, 300, 298, 298, 300, 295, 298, 
    293, 292, 297, 301, 299, 301, 302, 312, 310, 297, 289, 303, 329, 338, 1, 
    11, 25, 21, 15, 13, 13, 10, 8, 4, 360, 348, 345, 342, 343, 341, 319, 302, 
    299, 306, 324, 324, 318, 297, 291, 299, 296, 293, 302, 300, 291, 307, 
    304, 298, 312, 300, 297, 299, 298, 294, 292, 290, 304, 291, 302, 291, 
    294, 295, 296, 292, 289, 298, 311, 289, 300, 345, 343, 331, 329, 324, 
    323, 334, 316, 313, 322, 347, 331, 352, 342, 316, 331, 310, 290, 308, 
    314, 287, 284, 291, 289, 280, 289, 276, 281, 300, 283, 301, 291, 302, 9, 
    33, 25, 45, 50, 59, 66, 64, 59, 55, 63, 74, 78, 148, 142, 142, 125, 118, 
    113, 111, 105, 101, 102, 102, 100, 99, 94, 93, 85, 74, 75, 85, 85, 89, 
    88, 88, 102, 93, 90, 81, 81, 82, 81, 72, 74, 83, 84, 80, 73, 74, 75, 75, 
    73, 74, 77, 72, 69, 68, 64, 64, 70, 66, 65, 65, 68, 72, 58, 41, 33, 32, 
    35, 35, 27, 29, 26, 16, 23, 24, 23, 20, 20, 24, 30, 21, 17, 11, 15, 45, 
    18, 17, 79, 54, 51, 48, 50, 52, 52, 52, 46, 46, 46, 45, 49, 42, 41, 33, 
    35, 37, 54, 50, 51, 53, 55, 51, 50, 48, 44, 46, 44, 46, 88, 37, 32, 20, 
    19, 25, 21, 14, 16, 16, 10, 357, 3, 7, 1, 356, 7, 18, 14, 18, 20, 4, 21, 
    358, 360, 352, 346, 351, 350, 346, 353, 348, 340, 336, 330, 340, 345, 
    330, 309, 298, 307, 308, 309, 309, 314, 327, 322, 308, 329, 330, 318, 
    315, 321, 322, 325, 313, 304, 305, 312, 315, 316, 316, 360, 356, 350, 
    338, 292, 302, 292, 292, 295, 293, 300, 304, 319, 329, 319, 336, 337, 
    356, 292, 295, 293, 312, 313, 320, 313, 328, 321, 327, 330, 318, 317, 
    323, 335, 332, 360, 7, 5, 3, 352, 348, 1, 19, 5, 2, 1, 355, 351, 2, 348, 
    3, 8, 9, 359, 340, 337, 332, 19, 355, 355, 357, 343, 340, 336, 325, 328, 
    331, 331, 330, 347, 351, 340, 333, 340, 4, 3, 15, 23, 19, 2, 15, 18, 7, 
    4, 22, 60, 52, 351, 77, 85, 100, 129, 114, 117, 109, 117, 92, 79, 80, 71, 
    67, 69, 72, 71, 59, 58, 59, 55, 53, 54, 54, 49, 51, 46, 48, 50, 57, 87, 
    93, 80, 68, 65, 77, 79, 89, 101, 93, 88, 94, 90, 82, 92, 96, 99, 95, 93, 
    95, 97, 96, 85, 81, 90, 105, 90, 84, 84, 88, 102, 92, 97, 104, 101, 101, 
    101, 108, 102, 107, 104, 103, 103, 103, 108, 106, 102, 102, 88, 105, 105, 
    105, 107, 114, 119, 150, 289, 286, 278, 293, 291, 290, 289, 287, 288, 
    289, 287, 289, 288, 293, 293, 287, 288, 287, 288, 287, 289, 285, 286, 
    287, 285, 286, 287, 285, 285, 284, 291, 292, 292, 289, 295, 291, 296, 
    288, 302, 301, 305, 304, 306, 308, 306, 304, 310, 298, 296, 3, 14, 42, 
    45, 70, 61, 75, 123, 116, 114, 76, 89, 71, 76, 83, 104, 92, 107, 114, 
    111, 137, 169, 282, 345, 42, 69, 32, 18, 15, 32, 37, 13, 347, 344, 347, 
    328, 307, 337, 335, 343, 359, 337, 352, 5, 354, 7, 22, 15, 60, 14, 18, 
    25, 19, 28, 32, 60, 80, 108, 112, 121, 119, 102, 119, 120, 112, 103, 99, 
    88, 83, 71, 70, 61, 63, 62, 68, 52, 43, 38, 356, 347, 66, 203, 310, 309, 
    300, 297, 295, 295, 290, 289, 287, 282, 280, 280, 285, 338, 347, 352, 
    355, 360, 2, 6, 18, 25, 26, 26, 12, 15, 27, 25, 20, 20, 323, 315, 315, 
    310, 311, 315, 307, 308, 305, 305, 308, 304, 314, 329, 331, 315, 334, 
    314, 300, 66, 104, 110, 156, 164, 159, 173, 154, 177, 175, 185, 186, 213, 
    225, 300, 307, 303, 306, 322, 307, 315, 339, 343, 343, 351, 2, 4, 329, 
    327, 94, 88, 83, 58, 59, 59, 65, 63, 63, 68, 66, 63, 74, 82, 88, 78, 74, 
    88, 97, 98, 103, 102, 97, 93, 91, 90, 89, 92, 100, 109, 124, 141, 299, 
    296, 291, 295, 300, 302, 302, 301, 309, 304, 308, 317, 316, 314, 316, 
    318, 313, 323, 324, 322, 322, 321, 317, 319, 315, 311, 313, 311, 312, 
    310, 308, 306, 305, 307, 307, 311, 309, 307, 309, 312, 316, 315, 309, 
    310, 310, 307, 305, 308, 309, 308, 312, 301, 296, 293, 293, 294, 292, 
    285, 285, 286, 285, 282, 281, 287, 288, 290, 291, 287, 299, 301, 307, 
    289, 297, 297, 296, 292, 297, 294, 299, 293, 290, 284, 285, 284, 283, 
    284, 292, 288, 291, 282, 278, 294, 304, 319, 331, 308, 310, 311, 311, 
    320, 340, 331, 329, 325, 323, 320, 324, 325, 332, 338, 333, 310, 312, 
    315, 315, 314, 311, 306, 302, 301, 307, 314, 310, 305, 293, 286, 283, 
    280, 270, 270, 280, 284, 289, 289, 287, 289, 284, 284, 284, 278, 298, 
    308, 300, 293, 293, 306, 298, 314, 328, 352, 5, 8, 1, 350, 360, 6, 333, 
    299, 339, 291, 326, 330, 48, 11, 329, 349, 349, 360, 8, 42, 317, 38, 12, 
    54, 51, 49, 49, 50, 51, 47, 46, 50, 53, 55, 56, 53, 59, 61, 65, 69, 67, 
    73, 78, 91, 109, 264, 260, 282, 293, 278, 303, 289, 282, 283, 300, 296, 
    298, 290, 285, 280, 280, 311, 290, 284, 293, 293, 274, 275, 275, 273, 
    273, 272, 275, 268, 280, 290, 293, 279, 285, 281, 279, 285, 288, 291, 
    281, 281, 283, 287, 291, 310, 306, 308, 299, 309, 334, 331, 316, 320, 
    336, 342, 320, 333, 352, 344, 34, 334, 328, 331, 334, 325, 326, 323, 333, 
    326, 323, 322, 321, 308, 307, 309, 304, 308, 311, 313, 304, 301, 303, 
    306, 304, 300, 300, 299, 302, 303, 302, 299, 297, 302, 306, 307, 307, 
    311, 303, 313, 321, 327, 324, 323, 323, 313, 322, 326, 320, 329, 328, 
    326, 326, 308, 304, 303, 307, 306, 306, 305, 305, 305, 303, 306, 305, 
    310, 305, 310, 300, 307, 309, 315, 311, 311, 316, 310, 304, 302, 300, 
    302, 290, 290, 288, 298, 295, 300, 306, 306, 310, 307, 309, 302, 311, 
    310, 336, 354, 331, 334, 352, 314, 294, 313, 333, 327, 329, 332, 306, 
    308, 310, 309, 307, 308, 317, 335, 327, 318, 307, 313, 300, 305, 305, 
    303, 304, 307, 301, 307, 308, 305, 312, 325, 325, 322, 315, 321, 315, 
    305, 309, 308, 302, 310, 327, 321, 334, 320, 319, 325, 322, 314, 317, 
    313, 314, 308, 304, 303, 302, 307, 307, 301, 300, 304, 296, 296, 314, 
    309, 278, 279, 301, 301, 314, 306, 308, 300, 306, 311, 319, 312, 312, 
    310, 309, 267, 285, 271, 284, 332, 333, 332, 351, 303, 320, 340, 18, 13, 
    45, 82, 9, 353, 359, 339, 344, 323, 333, 324, 321, 11, 326, 5, 360, 331, 
    3, 6, 16, 3, 10, 334, 339, 348, 346, 350, 337, 336, 333, 332, 328, 330, 
    335, 340, 340, 332, 312, 329, 329, 360, 76, 69, 67, 70, 71, 88, 72, 100, 
    195, 287, 300, 257, 54, 348, 320, 318, 317, 325, 360, 54, 61, 57, 60, 42, 
    13, 35, 48, 54, 360, 334, 238, 54, 35, 12, 350, 93, 107, 104, 113, 119, 
    124, 78, 72, 64, 57, 63, 59, 59, 7, 359, 255, 67, 68, 61, 63, 57, 53, 60, 
    71, 67, 106, 87, 141, 142, 97, 112, 110, 100, 123, 108, 104, 107, 111, 
    115, 110, 130, 120, 112, 86, 89, 89, 84, 80, 68, 89, 93, 95, 114, 114, 
    121, 120, 115, 121, 119, 121, 126, 121, 117, 109, 121, 114, 122, 104, 
    109, 110, 110, 109, 111, 110, 112, 116, 113, 122, 120, 115, 108, 120, 93, 
    107, 107, 105, 111, 110, 105, 113, 94, 88, 88, 68, 82, 76, 92, 77, 88, 
    81, 74, 74, 69, 71, 84, 76, 63, 72, 67, 65, 56, 52, 56, 51, 51, 334, 330, 
    326, 44, 42, 54, 341, 55, 33, 322, 317, 341, 358, 313, 314, 303, 333, 52, 
    57, 52, 54, 56, 60, 67, 30, 0, 0, 322, 0, 0, 319, 317, 317, 0, 137, 129, 
    133, 131, 133, 122, 120, 117, 128, 149, 0, 32, 325, 304, 312, 317, 322, 
    360, 0, 0, 0, 317, 315, 305, 311, 326, 313, 280, 296, 24, 121, 102, 310, 
    314, 302, 301, 323, 323, 304, 302, 309, 310, 319, 309, 309, 297, 297, 
    306, 311, 312, 301, 304, 306, 301, 315, 310, 306, 306, 336, 302, 306, 
    310, 312, 319, 318, 316, 324, 323, 304, 303, 304, 307, 303, 310, 316, 
    316, 312, 310, 314, 314, 317, 320, 320, 320, 324, 330, 329, 328, 326, 
    323, 328, 330, 326, 331, 328, 328, 329, 326, 324, 326, 326, 330, 332, 
    332, 327, 328, 328, 325, 324, 329, 328, 329, 325, 329, 323, 322, 322, 
    314, 320, 330, 314, 317, 311, 305, 316, 43, 30, 45, 41, 41, 45, 313, 297, 
    360, 327, 341, 200, 192, 343, 318, 324, 325, 322, 310, 309, 341, 341, 3, 
    305, 33, 2, 351, 329, 1, 53, 58, 59, 56, 66, 110, 111, 113, 132, 112, 
    123, 144, 68, 55, 51, 62, 64, 61, 59, 57, 57, 54, 59, 60, 59, 60, 57, 58, 
    58, 56, 58, 59, 58, 49, 56, 57, 56, 58, 58, 59, 56, 58, 61, 54, 50, 41, 
    40, 35, 44, 54, 54, 44, 42, 40, 30, 15, 16, 23, 287, 304, 34, 6, 343, 17, 
    2, 7, 357, 25, 25, 35, 37, 26, 25, 352, 349, 344, 341, 340, 4, 322, 328, 
    328, 316, 322, 326, 330, 326, 324, 327, 332, 335, 335, 340, 341, 334, 
    332, 338, 336, 336, 338, 328, 340, 341, 334, 330, 337, 317, 322, 311, 
    317, 310, 313, 307, 315, 311, 309, 297, 302, 290, 305, 315, 306, 299, 
    291, 286, 294, 293, 298, 300, 307, 290, 304, 311, 309, 304, 297, 300, 
    300, 295, 313, 312, 324, 308, 297, 289, 287, 282, 286, 291, 299, 335, 
    333, 290, 296, 286, 286, 278, 280, 285, 285, 278, 281, 291, 284, 286, 
    294, 294, 314, 323, 320, 319, 317, 319, 337, 323, 321, 320, 331, 324, 
    314, 322, 277, 267, 277, 267, 272, 257, 268, 239, 231, 256, 199, 172, 
    150, 149, 157, 140, 135, 147, 157, 188, 225, 283, 289, 285, 282, 283, 
    284, 301, 298, 302, 304, 305, 307, 316, 319, 340, 8, 67, 114, 114, 103, 
    113, 105, 113, 104, 112, 107, 108, 106, 100, 82, 96, 104, 92, 102, 116, 
    114, 0, 353, 291, 334, 0, 120, 99, 252, 273, 297, 298, 315, 316, 326, 
    321, 327, 325, 309, 311, 320, 318, 308, 313, 313, 312, 298, 301, 298, 
    299, 312, 301, 294, 293, 295, 282, 287, 283, 277, 271, 261, 261, 281, 
    253, 251, 226, 210, 173, 191, 177, 158, 148, 154, 138, 141, 134, 133, 
    132, 130, 129, 126, 122, 125, 132, 132, 137, 136, 135, 133, 130, 126, 
    125, 127, 130, 138, 140, 149, 155, 169, 144, 302, 307, 305, 305, 308, 
    302, 310, 294, 301, 289, 291, 294, 284, 290, 294, 293, 291, 296, 300, 
    293, 300, 299, 297, 297, 306, 309, 310, 301, 304, 295, 295, 358, 29, 112, 
    125, 130, 121, 111, 110, 102, 108, 111, 110, 106, 88, 85, 60, 57, 50, 50, 
    50, 52, 291, 104, 340, 31, 292, 6, 27, 25, 28, 11, 347, 342, 352, 355, 
    344, 334, 324, 330, 324, 325, 332, 323, 319, 320, 314, 326, 324, 316, 
    314, 316, 324, 325, 316, 316, 318, 314, 313, 312, 305, 315, 315, 316, 
    321, 314, 322, 319, 309, 307, 307, 308, 308, 326, 324, 327, 321, 319, 
    331, 333, 329, 329, 328, 328, 333, 332, 326, 329, 330, 331, 331, 330, 
    326, 326, 330, 331, 333, 330, 328, 326, 326, 325, 324, 336, 332, 328, 
    321, 316, 326, 323, 317, 328, 326, 329, 321, 314, 323, 327, 319, 324, 
    315, 316, 330, 333, 319, 321, 328, 313, 333, 328, 326, 317, 324, 326, 
    328, 313, 323, 333, 320, 326, 329, 319, 322, 326, 328, 330, 335, 330, 
    328, 334, 337, 329, 327, 323, 332, 330, 331, 342, 334, 335, 332, 337, 
    340, 345, 350, 345, 337, 347, 341, 326, 332, 342, 333, 335, 350, 340, 
    347, 322, 330, 308, 324, 337, 321, 330, 335, 338, 349, 0, 331, 346, 323, 
    319, 331, 323, 329, 321, 328, 308, 324, 325, 328, 76, 81, 68, 76, 107, 
    62, 299, 319, 9, 316, 0, 264, 114, 57, 79, 108, 153, 197, 206, 174, 175, 
    133, 155, 125, 147, 142, 157, 130, 140, 152, 138, 146, 151, 153, 137, 
    126, 159, 155, 182, 182, 172, 156, 176, 132, 121, 113, 170, 140, 114, 
    107, 113, 102, 116, 115, 114, 120, 114, 122, 111, 117, 121, 125, 133, 
    131, 116, 120, 124, 129, 110, 128, 129, 114, 105, 112, 119, 120, 118, 
    111, 118, 115, 115, 131, 117, 116, 114, 115, 129, 163, 151, 156, 164, 
    214, 264, 304, 299, 294, 294, 297, 308, 301, 307, 301, 299, 311, 295, 
    293, 279, 279, 278, 280, 279, 288, 301, 299, 294, 298, 300, 296, 309, 
    305, 307, 305, 310, 306, 306, 302, 300, 294, 283, 295, 303, 298, 302, 
    329, 337, 332, 327, 314, 333, 322, 336, 330, 331, 339, 332, 323, 348, 
    335, 339, 330, 323, 341, 338, 319, 333, 326, 324, 333, 337, 326, 324, 
    331, 326, 335, 355, 332, 351, 350, 349, 11, 346, 321, 340, 2, 335, 328, 
    320, 321, 332, 315, 318, 315, 338, 348, 337, 320, 356, 345, 333, 351, 
    347, 313, 359, 329, 344, 13, 347, 3, 360, 328, 315, 327, 298, 295, 338, 
    86, 108, 140, 113, 146, 131, 119, 118, 115, 120, 116, 122, 119, 121, 122, 
    121, 123, 155, 146, 131, 137, 123, 133, 110, 97, 116, 117, 114, 115, 94, 
    100, 112, 116, 118, 117, 117, 115, 114, 121, 138, 120, 119, 221, 316, 
    309, 316, 328, 329, 319, 319, 308, 311, 305, 300, 299, 304, 308, 315, 
    297, 327, 341, 327, 274, 314, 298, 324, 284, 291, 289, 298, 310, 337, 
    319, 319, 309, 299, 290, 295, 300, 301, 302, 307, 309, 309, 297, 299, 
    301, 359, 358, 331, 327, 344, 321, 359, 335, 339, 332, 324, 322, 322, 
    326, 329, 316, 302, 323, 325, 22, 3, 350, 331, 327, 345, 333, 313, 306, 
    317, 319, 305, 308, 301, 294, 282, 288, 287, 280, 280, 279, 283, 286, 
    286, 292, 288, 300, 306, 302, 293, 304, 293, 290, 283, 284, 289, 298, 
    287, 277, 274, 271, 273, 254, 261, 289, 278, 264, 278, 264, 244, 249, 
    236, 250, 283, 259, 347, 338, 337, 278, 0, 0, 360, 266, 280, 314, 22, 17, 
    356, 340, 336, 326, 319, 336, 341, 331, 356, 345, 49, 46, 58, 42, 30, 29, 
    38, 43, 27, 22, 16, 1, 342, 27, 18, 360, 336, 339, 335, 335, 338, 327, 
    322, 332, 330, 320, 317, 326, 336, 330, 341, 352, 338, 358, 2, 7, 352, 7, 
    17, 12, 359, 358, 349, 357, 2, 10, 12, 24, 23, 28, 34, 25, 27, 32, 30, 
    36, 37, 14, 33, 39, 34, 24, 45, 44, 47, 45, 41, 38, 32, 39, 42, 43, 40, 
    40, 316, 328, 40, 32, 298, 85, 58, 289, 341, 360, 15, 299, 299, 292, 294, 
    345, 8, 26, 42, 49, 52, 44, 360, 346, 334, 18, 13, 20, 25, 17, 29, 36, 
    31, 251, 45, 60, 64, 349, 34, 64, 28, 355, 29, 25, 23, 17, 51, 45, 40, 
    352, 74, 58, 318, 140, 9, 2, 347, 347, 306, 284, 267, 150, 146, 133, 151, 
    127, 129, 125, 136, 110, 158, 144, 141, 132, 145, 160, 159, 153, 129, 
    152, 154, 126, 137, 131, 140, 131, 173, 124, 115, 127, 135, 128, 155, 
    118, 96, 90, 120, 128, 114, 162, 193, 201, 180, 107, 70, 72, 63, 60, 59, 
    60, 133, 113, 135, 158, 174, 128, 108, 110, 162, 132, 110, 124, 117, 120, 
    104, 146, 115, 136, 140, 146, 144, 150, 138, 147, 207, 175, 150, 265, 
    280, 250, 123, 124, 130, 292, 355, 0, 143, 287, 57, 66, 67, 76, 60, 75, 
    61, 69, 64, 67, 63, 60, 61, 61, 101, 110, 64, 78, 81, 91, 86, 95, 98, 94, 
    124, 134, 114, 65, 90, 84, 85, 135, 149, 151, 305, 286, 135, 8, 323, 326, 
    319, 316, 315, 320, 325, 330, 338, 350, 319, 322, 26, 30, 2, 340, 343, 
    322, 308, 305, 313, 302, 302, 287, 301, 328, 280, 248, 285, 264, 313, 
    284, 298, 305, 309, 321, 317, 314, 336, 332, 322, 318, 320, 320, 320, 
    314, 315, 307, 302, 318, 323, 323, 297, 308, 319, 307, 312, 313, 301, 
    312, 316, 312, 324, 322, 314, 317, 326, 327, 345, 330, 332, 346, 343, 1, 
    282, 133, 90, 116, 66, 303, 310, 312, 306, 306, 309, 314, 314, 314, 313, 
    311, 312, 319, 311, 315, 318, 312, 313, 302, 322, 320, 330, 317, 305, 
    312, 319, 325, 322, 311, 306, 310, 315, 320, 316, 313, 360, 1, 339, 334, 
    328, 329, 330, 326, 326, 329, 325, 323, 333, 335, 339, 335, 334, 317, 
    325, 322, 329, 319, 316, 316, 298, 319, 318, 295, 302, 310, 316, 312, 
    313, 317, 317, 315, 314, 310, 309, 312, 308, 304, 302, 299, 323, 323, 
    320, 328, 335, 347, 357, 41, 314, 63, 77, 69, 93, 90, 76, 95, 100, 110, 
    105, 117, 105, 121, 125, 136, 132, 140, 154, 113, 115, 120, 110, 141, 
    124, 138, 129, 127, 119, 109, 121, 122, 125, 129, 163, 133, 54, 75, 60, 
    60, 55, 73, 229, 300, 342, 322, 312, 305, 303, 309, 296, 293, 282, 284, 
    297, 287, 304, 300, 283, 289, 294, 292, 293, 291, 292, 289, 295, 288, 
    300, 287, 297, 303, 309, 303, 310, 293, 308, 320, 304, 299, 312, 306, 
    299, 287, 299, 306, 314, 284, 296, 306, 282, 291, 300, 302, 299, 303, 
    297, 298, 300, 295, 297, 301, 302, 306, 299, 302, 296, 298, 321, 327, 
    306, 314, 318, 311, 310, 306, 292, 256, 300, 284, 276, 308, 299, 295, 
    287, 285, 281, 280, 292, 292, 295, 296, 306, 302, 312, 313, 302, 285, 
    306, 306, 263, 249, 254, 276, 295, 294, 265, 262, 268, 280, 258, 266, 
    286, 271, 246, 249, 273, 272, 261, 277, 267, 286, 265, 266, 270, 278, 
    276, 280, 282, 281, 280, 281, 293, 294, 290, 282, 275, 284, 274, 267, 
    270, 269, 265, 263, 280, 243, 244, 258, 272, 271, 274, 273, 278, 271, 
    266, 264, 272, 274, 276, 255, 262, 249, 261, 284, 285, 262, 244, 267, 
    257, 257, 272, 275, 254, 223, 236, 238, 238, 245, 253, 288, 289, 294, 
    292, 286, 295, 305, 302, 305, 305, 305, 294, 326, 334, 315, 316, 307, 
    321, 320, 313, 335, 305, 312, 315, 322, 317, 315, 298, 304, 304, 300, 
    307, 315, 301, 303, 307, 307, 310, 306, 289, 250, 235, 256, 257, 0, 0, 
    156, 173, 156, 161, 140, 137, 135, 130, 126, 122, 110, 125, 125, 122, 
    125, 123, 125, 130, 125, 125, 137, 122, 143, 117, 139, 129, 125, 118, 
    121, 130, 131, 131, 130, 124, 121, 135, 136, 133, 127, 110, 118, 120, 
    123, 112, 117, 129, 124, 107, 112, 117, 120, 118, 120, 118, 120, 120, 
    119, 122, 129, 118, 117, 117, 114, 115, 120, 112, 113, 110, 115, 123, 
    120, 113, 107, 107, 105, 107, 105, 105, 102, 102, 92, 102, 101, 105, 99, 
    93, 93, 108, 93, 126, 135, 156, 285, 302, 310, 302, 294, 297, 291, 285, 
    284, 284, 289, 287, 286, 295, 298, 290, 287, 288, 286, 285, 283, 287, 
    274, 269, 275, 270, 274, 270, 270, 268, 288, 275, 297, 311, 307, 324, 
    307, 300, 298, 295, 280, 279, 287, 288, 282, 279, 276, 300, 325, 313, 
    304, 296, 295, 293, 312, 313, 308, 300, 290, 293, 344, 323, 325, 337, 
    348, 330, 259, 275, 300, 264, 306, 302, 302, 287, 298, 290, 287, 275, 
    308, 271, 303, 291, 296, 312, 294, 266, 327, 212, 156, 153, 165, 135, 
    137, 139, 134, 134, 137, 143, 134, 136, 133, 135, 135, 132, 128, 125, 
    122, 120, 124, 119, 113, 112, 101, 121, 109, 70, 83, 74, 77, 86, 88, 80, 
    87, 70, 78, 74, 63, 86, 83, 87, 111, 135, 170, 157, 150, 141, 129, 131, 
    144, 149, 156, 155, 161, 180, 203, 188, 139, 136, 129, 130, 117, 141, 
    134, 135, 9, 124, 0, 160, 137, 150, 137, 127, 128, 125, 130, 129, 129, 
    176, 159, 355, 284, 130, 170, 178, 281, 140, 100, 68, 210, 131, 81, 134, 
    316, 97, 93, 9, 360, 320, 215, 261, 272, 244, 225, 186, 246, 201, 251, 
    177, 28, 13, 339, 11, 357, 339, 334, 335, 348, 330, 327, 330, 330, 316, 
    309, 306, 310, 304, 297, 292, 290, 286, 285, 280, 280, 284, 287, 283, 
    279, 280, 270, 270, 271, 267, 254, 252, 253, 256, 252, 259, 264, 267, 
    260, 246, 262, 279, 289, 267, 297, 290, 301, 285, 333, 337, 236, 297, 
    310, 331, 249, 71, 136, 170, 122, 171, 174, 141, 163, 158, 122, 122, 133, 
    144, 117, 200, 276, 279, 324, 319, 227, 200, 153, 135, 129, 128, 123, 
    130, 127, 129, 123, 129, 125, 120, 122, 124, 114, 118, 126, 120, 113, 
    115, 122, 133, 122, 123, 116, 125, 113, 117, 131, 134, 133, 130, 141, 
    144, 146, 145, 153, 141, 150, 159, 149, 159, 166, 148, 149, 151, 102, 
    281, 271, 228, 310, 280, 310, 314, 274, 282, 320, 245, 339, 55, 57, 60, 
    62, 60, 56, 61, 66, 62, 84, 77, 87, 114, 130, 203, 302, 316, 311, 85, 
    130, 141, 137, 137, 130, 163, 158, 138, 159, 190, 167, 168, 144, 139, 
    143, 128, 129, 177, 115, 120, 131, 166, 328, 245, 341, 343, 353, 130, 96, 
    137, 79, 75, 85, 83, 98, 113, 127, 106, 137, 134, 129, 136, 106, 128, 
    136, 113, 119, 99, 75, 62, 59, 61, 62, 58, 67, 72, 82, 91, 85, 111, 123, 
    125, 131, 122, 122, 123, 120, 125, 127, 116, 124, 118, 116, 116, 116, 
    123, 106, 110, 105, 109, 106, 109, 109, 103, 82, 124, 91, 93, 100, 107, 
    119, 133, 130, 125, 128, 139, 136, 150, 135, 127, 137, 128, 92, 318, 304, 
    284, 340, 327, 292, 305, 317, 323, 307, 280, 91, 55, 43, 49, 45, 30, 324, 
    226, 2, 10, 68, 74, 77, 285, 240, 308, 100, 133, 201, 303, 310, 302, 310, 
    322, 322, 324, 322, 318, 271, 300, 330, 151, 130, 131, 130, 128, 129, 
    126, 118, 113, 109, 111, 119, 118, 107, 112, 111, 110, 115, 123, 122, 
    141, 146, 175, 145, 268, 313, 321, 15, 12, 14, 19, 14, 11, 1, 326, 307, 
    316, 319, 328, 337, 26, 97, 124, 131, 112, 107, 117, 121, 119, 120, 119, 
    116, 116, 115, 119, 115, 118, 117, 120, 122, 116, 120, 128, 135, 115, 
    118, 136, 223, 39, 238, 280, 321, 325, 251, 265, 282, 243, 245, 160, 276, 
    289, 320, 304, 317, 301, 293, 341, 348, 167, 126, 140, 128, 129, 136, 
    125, 141, 149, 154, 151, 162, 169, 166, 163, 160, 157, 145, 177, 160, 
    150, 161, 176, 155, 350, 345, 356, 359, 357, 352, 359, 358, 3, 360, 349, 
    359, 358, 352, 159, 275, 314, 353, 4, 0, 320, 347, 0, 0, 0, 0, 0, 0, 228, 
    216, 225, 214, 190, 188, 176, 148, 184, 175, 173, 170, 173, 176, 169, 
    142, 141, 138, 128, 147, 162, 153, 156, 156, 158, 156, 142, 109, 128, 
    113, 113, 134, 132, 132, 157, 163, 149, 152, 127, 151, 158, 143, 172, 
    161, 176, 184, 175, 176, 331, 359, 354, 357, 352, 352, 356, 359, 2, 359, 
    360, 355, 5, 359, 3, 11, 359, 1, 360, 7, 6, 5, 358, 358, 356, 348, 354, 
    358, 357, 347, 349, 349, 337, 337, 355, 357, 349, 346, 359, 351, 359, 
    358, 355, 352, 357, 354, 357, 1, 352, 343, 342, 341, 346, 354, 343, 328, 
    346, 336, 336, 340, 337, 331, 328, 334, 337, 351, 6, 6, 357, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 17, 336, 0, 0, 327, 358, 177, 174, 344, 236, 212, 0, 358, 357, 358, 
    7, 354, 358, 357, 350, 360, 338, 340, 332, 347, 352, 351, 333, 331, 334, 
    340, 340, 342, 351, 350, 333, 341, 357, 358, 346, 344, 31, 352, 283, 0, 
    0, 0, 360, 244, 0, 15, 213, 322, 317, 14, 12, 358, 1, 20, 360, 0, 360, 9, 
    341, 3, 346, 350, 5, 20, 5, 359, 354, 338, 342, 5, 11, 9, 351, 13, 11, 2, 
    349, 349, 13, 8, 16, 40, 356, 242, 277, 0, 337, 0, 0, 0, 11, 358, 309, 
    199, 198, 359, 355, 346, 350, 355, 349, 348, 359, 1, 356, 353, 354, 342, 
    3, 354, 11, 13, 18, 355, 296, 307, 355, 351, 359, 311, 51, 149, 157, 155, 
    170, 159, 151, 160, 164, 159, 155, 169, 161, 163, 154, 149, 150, 153, 
    160, 155, 154, 158, 161, 169, 163, 163, 153, 153, 167, 161, 167, 161, 
    158, 160, 161, 161, 157, 157, 159, 162, 156, 159, 163, 156, 167, 170, 
    172, 0, 7, 322, 360, 1, 4, 341, 2, 15, 339, 321, 7, 8, 21, 360, 0, 0, 
    358, 174, 104, 213, 184, 162, 155, 152, 128, 122, 112, 125, 111, 167, 
    140, 137, 142, 153, 157, 154, 144, 145, 157, 142, 141, 152, 147, 143, 
    154, 134, 148, 152, 153, 154, 152, 158, 155, 156, 157, 158, 159, 160, 
    159, 160, 159, 158, 157, 148, 141, 143, 139, 136, 145, 149, 149, 145, 
    144, 137, 144, 142, 142, 140, 132, 131, 136, 126, 123, 124, 137, 137, 
    138, 141, 133, 125, 134, 126, 128, 130, 135, 138, 137, 133, 132, 139, 
    143, 138, 141, 143, 147, 120, 118, 106, 134, 100, 112, 117, 151, 149, 
    124, 128, 102, 106, 104, 100, 95, 105, 108, 107, 106, 105, 106, 105, 103, 
    102, 101, 100, 106, 107, 103, 103, 100, 103, 107, 106, 99, 95, 94, 91, 
    87, 95, 91, 101, 102, 94, 85, 74, 332, 75, 354, 0, 0, 0, 331, 16, 10, 1, 
    3, 7, 6, 2, 360, 358, 359, 354, 355, 348, 346, 347, 341, 339, 353, 340, 
    342, 334, 344, 336, 3, 1, 348, 335, 329, 349, 341, 359, 350, 320, 314, 
    360, 5, 6, 7, 1, 332, 336, 322, 327, 328, 323, 321, 318, 307, 306, 307, 
    290, 281, 274, 275, 276, 273, 278, 296, 301, 305, 319, 325, 328, 329, 
    332, 333, 341, 336, 333, 335, 328, 329, 332, 330, 331, 331, 325, 324, 
    332, 331, 348, 350, 342, 7, 342, 335, 321, 320, 334, 335, 332, 332, 329, 
    330, 333, 328, 330, 333, 328, 325, 324, 324, 306, 305, 309, 310, 317, 
    317, 324, 333, 331, 0, 315, 315, 314, 327, 332, 340, 335, 335, 343, 339, 
    327, 344, 350, 356, 316, 337, 331, 325, 321, 321, 321, 321, 330, 332, 
    344, 351, 332, 318, 319, 329, 348, 341, 338, 342, 320, 319, 325, 327, 
    346, 340, 348, 322, 339, 345, 345, 339, 326, 318, 325, 320, 321, 323, 
    337, 333, 340, 343, 9, 6, 11, 3, 4, 5, 356, 7, 357, 348, 349, 360, 4, 
    340, 343, 356, 339, 337, 343, 354, 332, 331, 5, 11, 360, 343, 147, 160, 
    162, 167, 151, 26, 0, 0, 350, 343, 358, 360, 0, 148, 147, 39, 151, 163, 
    155, 162, 169, 168, 166, 169, 172, 164, 168, 166, 178, 170, 166, 134, 
    147, 138, 138, 143, 133, 143, 150, 146, 150, 155, 156, 156, 157, 149, 
    157, 165, 159, 155, 152, 152, 157, 154, 156, 156, 158, 154, 151, 152, 
    154, 154, 152, 147, 150, 153, 154, 150, 147, 150, 148, 142, 143, 143, 
    143, 139, 141, 139, 144, 152, 112, 148, 188, 167, 1, 323, 349, 4, 3, 358, 
    352, 340, 341, 293, 343, 0, 0, 241, 265, 255, 240, 213, 183, 170, 169, 
    181, 170, 157, 158, 151, 156, 154, 139, 155, 131, 146, 146, 159, 153, 
    139, 133, 146, 149, 155, 156, 160, 161, 154, 155, 157, 157, 153, 146, 
    141, 150, 144, 126, 115, 149, 169, 162, 169, 157, 145, 135, 147, 156, 
    152, 163, 158, 160, 155, 154, 160, 156, 153, 146, 137, 155, 138, 130, 
    127, 119, 126, 113, 101, 100, 108, 115, 117, 118, 117, 130, 125, 122, 
    119, 163, 165, 0, 356, 1, 347, 360, 1, 2, 360, 359, 357, 358, 359, 358, 
    356, 357, 350, 353, 351, 358, 354, 357, 354, 354, 355, 353, 357, 3, 360, 
    3, 353, 343, 339, 346, 354, 348, 354, 349, 354, 2, 3, 4, 5, 352, 349, 
    350, 354, 4, 0, 69, 175, 167, 141, 143, 129, 162, 134, 130, 127, 120, 
    117, 123, 127, 124, 144, 146, 149, 148, 154, 153, 135, 140, 141, 143, 
    145, 140, 136, 138, 142, 151, 147, 157, 155, 156, 155, 155, 154, 149, 
    151, 149, 147, 142, 141, 139, 138, 138, 137, 148, 144, 149, 143, 144, 
    150, 153, 148, 180, 204, 19, 0, 310, 358, 5, 357, 335, 310, 304, 339, 
    350, 300, 268, 280, 288, 305, 332, 334, 330, 335, 331, 327, 331, 335, 
    337, 343, 345, 334, 336, 337, 339, 329, 349, 336, 347, 349, 351, 353, 
    350, 9, 8, 68, 39, 3, 123, 138, 151, 160, 160, 170, 156, 141, 126, 111, 
    115, 124, 121, 124, 123, 145, 144, 147, 135, 130, 136, 126, 134, 148, 
    150, 153, 151, 157, 149, 150, 146, 146, 149, 147, 148, 149, 145, 141, 
    141, 139, 135, 130, 127, 126, 129, 130, 133, 134, 131, 129, 129, 127, 
    129, 131, 130, 124, 132, 139, 141, 139, 141, 145, 149, 150, 148, 150, 
    149, 156, 154, 159, 152, 158, 150, 164, 156, 146, 156, 162, 164, 167, 
    156, 157, 157, 160, 158, 159, 156, 160, 151, 159, 165, 161, 159, 156, 
    157, 155, 158, 153, 160, 160, 159, 156, 157, 158, 154, 155, 155, 157, 
    155, 155, 156, 156, 156, 154, 154, 156, 154, 157, 158, 157, 160, 154, 
    156, 154, 153, 155, 152, 152, 151, 151, 151, 150, 147, 149, 147, 146, 
    143, 142, 143, 147, 146, 149, 149, 144, 148, 153, 155, 153, 139, 140, 
    135, 133, 148, 147, 147, 147, 143, 146, 132, 125, 114, 106, 113, 127, 
    133, 144, 138, 147, 136, 129, 126, 126, 150, 151, 137, 146, 145, 145, 
    145, 136, 133, 137, 144, 138, 142, 138, 141, 141, 150, 145, 142, 146, 
    152, 160, 113, 115, 100, 110, 117, 42, 100, 156, 166, 177, 178, 158, 0, 
    359, 5, 342, 7, 358, 15, 356, 80, 0, 0, 2, 3, 0, 0, 0, 0, 0, 5, 0, 1, 0, 
    0, 0, 165, 72, 359, 1, 142, 141, 143, 139, 147, 142, 159, 158, 165, 159, 
    176, 162, 167, 176, 161, 167, 164, 165, 161, 169, 155, 158, 160, 151, 
    153, 150, 152, 163, 153, 155, 164, 159, 160, 162, 158, 154, 152, 153, 
    154, 149, 152, 152, 160, 167, 176, 140, 146, 10, 0, 0, 0, 2, 21, 0, 137, 
    157, 155, 155, 161, 153, 156, 159, 170, 154, 155, 154, 150, 155, 162, 
    181, 165, 167, 166, 156, 178, 143, 151, 136, 152, 158, 166, 159, 3, 25, 
    9, 355, 19, 1, 344, 347, 338, 334, 330, 332, 331, 320, 323, 317, 320, 
    320, 327, 329, 333, 326, 330, 328, 335, 321, 325, 318, 327, 329, 328, 
    318, 316, 320, 320, 317, 315, 316, 315, 306, 294, 275, 253, 245, 228, 
    217, 209, 208, 237, 252, 259, 308, 335, 343, 347, 337, 330, 333, 342, 
    342, 335, 345, 334, 3, 360, 341, 346, 353, 3, 144, 146, 149, 187, 179, 
    175, 167, 173, 171, 169, 170, 160, 164, 156, 156, 153, 155, 155, 149, 
    153, 147, 140, 131, _, _, _, _, _, _, _, 129, 152, 132, 163, 151, 155, 
    155, 149, 150, 156, 136, 162, 169, 172, 146, 174, 0, 0, 5, 354, 350, 5, 
    359, 350, 358, 3, 1, 342, 349, 345, 346, 336, 328, 326, 328, 314, 332, 
    286, 297, 311, 339, 267, 200, 171, 192, 170, 185, 161, 150, 155, 147, 
    152, 151, 153, 152, 153, 153, 153, 156, 153, 153, 162, 152, 153, 160, 
    164, 178, 147, 159, 186, 174, 149, 327, 162, 114, 44, 0, 20, 41, 54, 6, 
    158, 0, 1, 7, 321, 7, 7, 146, 151, 161, 208, 164, 161, 164, 163, 0, 3, 
    342, 8, 1, 1, 355, 347, 352, 348, 309, 326, 354, 279, 241, 238, 237, 235, 
    200, 183, 163, 155, 150, 158, 154, 166, 240, 6, 0, 0, 156, 238, 6, 129, 
    243, 208, 179, 201, 194, 171, 237, 2, 141, 134, 205, 169, 166, 276, 176, 
    160, 159, 169, 174, 154, 169, 160, 157, 165, 159, 154, 163, 163, 163, 
    165, 171, 156, 153, 269, 22, 169, 358, 196, 206, 78, 18, 8, 4, 4, 12, 3, 
    353, 0, 0, 0, 0, 176, 156, 173, 178, 149, 150, 165, 163, 162, 165, 151, 
    148, 167, 164, 152, 148, 145, 142, 156, 158, 154, 156, 157, 164, 156, 
    167, 151, 157, 154, 161, 153, 161, 152, 154, 150, 156, 158, 167, 173, 
    175, 162, 155, 152, 157, 160, 161, 157, 160, 157, 157, 157, 156, 157, 
    156, 155, 156, 159, 158, 156, 158, 161, 155, 160, 161, 161, 162, 156, 
    158, 162, 155, 150, 139, 115, 110, 111, 110, 114, 115, 116, 0, 4, 360, 8, 
    163, 0, 0, 1, 359, 360, 360, 25, 1, 360, 5, 356, 35, 33, 351, 49, 49, 38, 
    33, 31, 30, 36, 18, 20, 36, 31, 23, 27, 24, 29, 19, 10, 5, 16, 23, 24, 
    20, 18, 32, 28, 30, 30, 19, 18, 18, 29, 37, 22, 37, 36, 12, 3, 4, 8, 5, 
    10, 12, 16, 7, 2, 356, 352, 352, 349, 360, 8, 20, 22, 19, 10, 8, 355, 
    360, 360, 7, 358, 11, 10, 9, 6, 10, 13, 13, 12, 14, 14, 10, 13, 15, 17, 
    14, 18, 26, 29, 46, 28, 19, 17, 7, 351, 30, 11, 54, 37, 35, 40, 41, 33, 
    46, 1, 360, 0, 35, 24, 41, 0, 0, 31, 221, 203, 223, 163, 140, 139, 160, 
    150, 149, 150, 148, 119, 113, 112, 108, 137, 153, 149, 149, 152, 0, 4, 
    17, 20, 25, 0, 105, 131, 163, 175, 159, 149, 152, 153, 162, 150, 152, 
    156, 157, 132, 164, 156, 7, 0, 0, 352, 11, 353, 92, 0, 0, 154, 182, 141, 
    166, 154, 163, 152, 156, 151, 158, 154, 185, 154, 150, 153, 155, 151, 
    150, 158, 156, 151, 153, 152, 158, 150, 150, 140, 155, 158, 172, 198, 
    157, 155, 158, 154, 153, 147, 140, 135, 139, 129, 122, 115, 110, 106, 
    105, 122, 115, 109, 125, 123, 121, 126, 130, 118, 120, 125, 130, 131, 
    131, 128, 134, 128, 135, 136, 132, 133, 134, 134, 130, 125, 136, 132, 
    134, 136, 140, 141, 138, 138, 138, 142, 141, 144, 143, 141, 139, 139, 
    135, 131, 126, 120, 116, 130, 126, 127, 124, 128, 130, 130, 130, 130, 
    126, 121, 127, 128, 128, 130, 126, 126, 125, 125, 125, 123, 122, 123, 
    125, 125, 124, 124, 124, 123, 125, 119, 120, 121, 125, 133, 128, 127, 
    129, 127, 129, 128, 130, 129, 126, 122, 116, 121, 117, 118, 120, 121, 
    127, 128, 134, 127, 130, 128, 129, 127, 123, 130, 130, 134, 129, 133, 
    140, 138, 139, 134, 135, 126, 128, 134, 131, 125, 139, 144, 124, 137, 
    133, 121, 119, 108, 105, 106, 99, 86, 85, 84, 92, 90, 76, 80, 85, 91, 68, 
    66, 62, 75, 54, 82, 66, 66, 66, 30, 35, 55, 63, 76, 82, 78, 69, 59, 67, 
    52, 65, 45, 24, 44, 62, 72, 74, 76, 65, 76, 42, 73, 50, 65, 68, 64, 57, 
    50, 52, 55, 52, 77, 71, 37, 47, 84, 103, 41, 68, 97, 124, 108, 0, 133, 
    132, 152, 159, 152, 145, 158, 176, 173, 173, 153, 163, 159, 174, 161, 
    169, 169, 189, 180, 194, 185, 187, 200, 183, 193, 185, 186, 188, 169, 
    176, 174, 159, 160, 159, 152, 146, 145, 134, 140, 162, 154, 156, 155, 
    145, 150, 163, 164, 360, 1, 3, 349, 360, 2, 1, 353, 360, 352, 347, 340, 
    334, 333, 328, 320, 329, 321, 324, 327, 328, 333, 341, 333, 327, 322, 
    336, 329, 328, 315, 311, 321, 321, 340, 330, 333, 342, 340, 338, 346, 
    328, 337, 354, 335, 360, 4, 358, 341, 2, 8, 348, 18, 17, 360, 356, 359, 
    347, 351, 28, 355, 37, 340, 331, 359, 346, 357, 360, 87, 108, 104, 105, 
    106, 112, 118, 133, 142, 139, 152, 166, 176, 172, 160, 153, 155, 142, 
    135, 137, 132, 120, 118, 122, 122, 116, 112, 109, 105, 103, 103, 98, 92, 
    89, 76, 74, 87, 75, 66, 67, 59, 61, 55, 51, 48, 42, 39, 38, 33, 33, 35, 
    38, 35, 37, 38, 37, 35, 34, 32, 26, 28, 28, 32, 39, 41, 38, 38, 36, 32, 
    29, 31, 32, 31, 31, 26, 28, 31, 20, 22, 16, 20, 20, 26, 59, 71, 72, 63, 
    54, 51, 42, 45, 49, 44, 44, 43, 40, 38, 37, 44, 50, 52, 47, 44, 35, 30, 
    28, 25, 19, 18, 18, 18, 20, 22, 18, 21, 26, 85, 90, 77, 16, 96, 92, 91, 
    86, 82, 36, 48, 38, 40, 358, 2, 4, 4, 14, 359, 346, 12, 329, 335, 325, 
    306, 297, 290, 289, 287, 284, 283, 278, 270, 283, 283, 277, 269, 270, 
    253, 251, 238, 240, 260, 251, 262, 258, 314, 244, 308, 222, 11, 321, 5, 
    129, 154, 175, 121, 146, 145, 147, 145, 119, 83, 97, 107, 114, 0, 83, 92, 
    87, 87, 84, 94, 102, 106, 116, 116, 119, 131, 125, 117, 117, 108, 106, 
    105, 95, 86, 87, 88, 89, 94, 92, 90, 87, 88, 88, 87, 90, 95, 98, 97, 100, 
    104, 107, 102, 105, 89, 91, 74, 73, 71, 59, 41, 45, 53, 64, 48, 42, 45, 
    48, 49, 55, 16, 343, 331, 330, 40, 340, 348, 16, 120, 97, 0, 77, 47, 45, 
    44, 50, 81, 83, 294, 0, 83, 72, 73, 80, 89, 85, 90, 94, 92, 90, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 105, 1, 100, 107, 25, 54, 68, 53, 48, 71, 0, 0, 70, 
    65, 60, 78, 66, 62, 60, 55, 72, 80, 82, 82, 82, 93, 92, 92, 85, 90, 92, 
    94, 84, 105, 123, 34, 85, 87, 90, 94, 100, 101, 101, 100, 101, 110, 101, 
    96, 97, 99, 97, 105, 97, 107, 113, 131, 133, 134, 120, 101, 116, 123, 
    124, 109, 101, 110, 109, 109, 113, 119, 110, 123, 110, 112, 112, 93, 93, 
    79, 88, 100, 111, 133, 132, 126, 130, 129, 124, 120, 117, 115, 122, 118, 
    114, 115, 116, 112, 98, 92, 90, 94, 97, 103, 101, 106, 106, 104, 102, 
    100, 102, 105, 103, 108, 110, 106, 107, 110, 99, 95, 98, 103, 102, 105, 
    107, 101, 100, 103, 102, 102, 101, 101, 100, 93, 91, 89, 89, 94, 95, 92, 
    100, 110, 112, 115, 105, 109, 110, 110, 111, 107, 103, 89, 99, 106, 131, 
    148, 152, 160, 152, 165, 151, 156, 157, 151, 157, 149, 152, 147, 149, 
    146, 138, 129, 124, 100, 102, 120, 136, 137, 118, 113, 115, 117, 132, 
    138, 140, 154, 133, 146, 140, 123, 113, 117, 119, 146, 145, 139, 145, 
    142, 140, 130, 127, 120, 127, 117, 120, 124, 117, 102, 104, 100, 96, 120, 
    150, 138, 131, 124, 121, 120, 114, 113, 112, 109, 111, 107, 107, 104, 
    107, 93, 79, 98, 110, 106, 115, 124, 119, 117, 123, 114, 125, 123, 117, 
    126, 119, 122, 113, 115, 100, 108, 100, 98, 91, 81, 87, 102, 99, 94, 91, 
    92, 100, 97, 95, 110, 104, 106, 109, 111, 118, 123, 113, 101, 101, 100, 
    97, 105, 106, 99, 99, 117, 109, 117, 103, 95, 108, 97, 91, 82, 85, 98, 
    80, 76, 62, 69, 78, 57, 60, 76, 64, 68, 66, 67, 64, 61, 62, 66, 65, 70, 
    73, 76, 68, 74, 73, 68, 66, 73, 59, 62, 77, 75, 74, 73, 72, 80, 87, 86, 
    86, 88, 84, 88, 78, 82, 79, 78, 91, 115, 109, 90, 80, 79, 70, 65, 88, 
    110, 100, 100, 97, 98, 94, 94, 88, 80, 81, 79, 80, 75, 73, 76, 75, 82, 
    83, 81, 60, 48, 77, 80, 98, 86, 79, 81, 80, 85, 88, 95, 93, 94, 99, 112, 
    38, 70, 76, 75, 90, 76, 78, 73, 76, 78, 90, 88, 86, 92, 82, 90, 98, 106, 
    104, 101, 104, 107, 112, 111, 114, 97, 101, 91, 108, 115, 138, 151, 122, 
    131, 124, 122, 142, 131, 115, 98, 145, 133, 134, 139, 149, 154, 136, 138, 
    134, 136, 137, 150, 159, 149, 125, 128, 127, 130, 132, 133, 143, 141, 
    145, 127, 142, 155, 127, 124, 140, 180, 224, 242, 230, 256, 252, 226, 
    237, 242, 247, 222, 230, 223, 253, 253, 234, 260, 254, 256, 258, 240, 
    286, 256, 235, 214, 248, 107, 263, 247, 221, 202, 209, 228, 241, 308, 
    283, 267, 249, 30, 19, 6, 26, 45, 51, 39, 41, 46, 13, 43, 43, 48, 34, 31, 
    25, 21, 15, 26, 31, 6, 75, 81, 81, 67, 58, 51, 38, 26, 33, 21, 18, 34, 
    46, 43, 41, 16, 91, 92, 96, 92, 85, 78, 83, 73, 70, 55, 53, 60, 58, 55, 
    50, 52, 44, 48, 58, 37, 42, 41, 36, 55, 56, 51, 70, 90, 109, 80, 118, 70, 
    63, 86, 81, 85, 85, 86, 87, 90, 107, 82, 87, 69, 67, 346, 96, 109, 127, 
    117, 108, 102, 96, 106, 97, 100, 104, 100, 101, 100, 106, 103, 109, 113, 
    120, 124, 114, 111, 99, 105, 124, 124, 118, 117, 122, 117, 115, 110, 104, 
    99, 96, 93, 123, 151, 150, 150, 153, 168, 156, 167, 156, 155, 155, 154, 
    147, 143, 133, 125, 131, 132, 125, 123, 122, 120, 117, 121, 123, 127, 
    124, 124, 122, 121, 115, 114, 113, 111, 111, 111, 113, 107, 103, 101, 
    102, 102, 99, 95, 105, 104, 106, 107, 103, 100, 101, 93, 92, 97, _, 82, 
    91, 89, 85, 88, 91, 88, 86, 85, 88, 88, 90, 87, 86, 85, 87, 81, 84, 84, 
    79, 74, 62, 62, 67, 67, 51, 60, 52, 59, 59, 66, 71, 86, 79, 79, 82, 74, 
    72, 80, 85, 78, 78, 83, 65, 85, 85, 83, 84, 94, 97, 95, 93, 96, 95, 91, 
    91, 92, 99, 93, 91, 94, 90, 91, 93, 96, 96, 95, 90, 95, 93, 90, 90, 91, 
    92, 88, 87, 85, 82, 89, 95, 94, 95, 89, 88, 83, 97, 110, 114, 123, 122, 
    120, 120, 123, 110, 100, 103, 106, 103, 103, 103, 105, 105, 100, 100, 
    107, 105, 109, 103, 103, 104, 110, 116, 117, 115, 115, 115, 108, 110, 
    107, 111, 103, 111, 111, 110, 108, 99, 100, 106, 109, 107, 121, 110, 110, 
    111, 105, 104, 106, 102, 106, 113, 124, 118, 111, 99, 106, 90, 93, 98, 
    89, 92, 94, 104, 137, 128, 129, 132, 129, 131, 124, 119, 115, 118, 121, 
    125, 129, 130, 123, 123, 120, 107, 102, 98, 95, 90, 98, 96, 95, 88, 112, 
    116, 116, 114, 110, 104, 105, 111, 114, 113, 113, 113, 115, 121, 122, 
    102, 104, 112, 115, 106, 97, 116, 119, 99, 106, 106, 103, 96, 91, 94, 91, 
    92, 88, 87, 89, 27, 84, 81, 68, 88, 86, 84, 88, 94, 82, 91, 88, 87, 90, 
    95, 112, 133, 140, 138, 136, 123, 112, 107, 101, 91, 105, 104, 102, 100, 
    94, 90, 87, 86, 82, 81, 81, 78, 23, 20, 337, 347, 11, 49, 46, 48, 44, 50, 
    55, 62, 51, 71, 66, 64, 75, 75, 81, 80, 325, 35, 17, 331, 338, 31, 2, 67, 
    77, 300, 302, 353, 14, 356, 87, 84, 84, 85, 88, 86, 87, 88, 88, 86, 84, 
    87, 88, 88, 89, 89, 87, 83, 90, 87, 87, 84, 85, 84, 85, 87, 88, 90, 91, 
    94, 97, 97, 97, 98, 103, 98, 99, 97, 102, 104, 91, 95, 98, 97, 104, 102, 
    101, 97, 96, 97, 99, 103, 104, 112, 126, 127, 130, 131, 140, 146, 139, 
    142, 146, 152, 141, 151, 152, 149, 148, 152, 178, 196, 192, 169, 160, 
    169, 157, 150, 146, 164, 155, 150, 150, 162, 157, 150, 163, 194, 155, 
    152, 159, 148, 149, 147, 143, 149, 140, 153, 149, 146, 144, 142, 136, 
    134, 130, 129, 127, 123, 124, 126, 132, 136, 142, 125, 124, 127, 128, 
    127, 126, 124, 124, 121, 118, 113, 109, 111, 114, 122, 139, 134, 130, 
    121, 127, 125, 123, 118, 112, 109, 116, 114, 109, 96, 88, 88, 93, 95, 
    114, 104, 91, 95, 101, 105, 107, 107, 108, 105, 109, 113, 99, 83, 78, 61, 
    77, 86, 91, 101, 110, 96, 95, 94, 96, 120, 122, 123, 126, 124, 118, 131, 
    134, 137, 136, 119, 124, 123, 117, 121, 123, 110, 106, 120, 109, 25, 12, 
    106, 53, 0, 72, 67, 75, 46, 40, 29, 54, 346, 352, 54, 46, 39, 47, 42, 37, 
    37, 40, 43, 34, 37, 47, 51, 47, 65, 69, 62, 59, 46, 59, 83, 83, 97, 76, 
    90, 325, 324, 332, 83, 76, 60, 43, 39, 47, 37, 33, 30, 35, 41, 53, 46, 
    39, 45, 34, 37, 34, 17, 16, 16, 1, 354, 357, 350, 352, 348, 6, 6, 1, 359, 
    3, 14, 13, 32, 28, 13, 25, 18, 15, 13, 19, 25, 13, 16, 16, 17, 23, 15, 
    19, 12, 8, 14, 17, 16, 21, 39, 89, 147, 168, 175, 166, 179, 184, 208, 
    239, 250, 304, 265, 256, 49, 100, 177, 150, 140, 126, 130, 137, 131, 339, 
    143, 128, 136, 117, 126, 85, 83, 84, 79, 57, 31, 20, 6, 6, 7, 1, 354, 
    353, 349, 1, 355, 352, 349, 349, 349, 349, 348, 349, 347, 349, 351, 352, 
    354, 350, 349, 349, 346, 334, 349, 354, 349, 359, 7, 9, 5, 14, 6, 5, 14, 
    4, 15, 17, 17, 27, 13, 20, 18, 17, 10, 8, 15, 17, 8, 8, 10, 19, 25, 14, 
    17, 29, 41, 33, 1, 40, 21, 34, 64, 90, 147, 40, 8, 38, 2, 9, 0, 50, 87, 
    45, 55, 82, 352, 87, 83, 91, 104, 108, 35, 23, 4, 70, 11, 77, 62, 49, 53, 
    17, 21, 23, 49, 15, 50, 53, 45, 40, 30, 27, 26, 20, 19, 11, 15, 14, 14, 
    11, 9, 8, 5, 17, 11, 13, 9, 14, 12, 11, 10, 10, 11, 11, 14, 12, 10, 8, 6, 
    4, 3, 359, 7, 6, 5, 360, 2, 2, 3, 7, 12, 25, 8, 339, 355, 6, 17, 14, 12, 
    15, 2, 15, 18, 23, 29, 38, 39, 37, 26, 26, 36, 38, 15, 343, 7, 11, 12, 7, 
    19, 16, 14, 15, 37, 39, 30, 35, 342, 3, 4, 8, 25, 8, 20, 0, 0, 0, 334, 
    327, 28, 80, 83, 83, 88, 89, 85, 95, 100, 99, 96, 94, 119, 140, 147, 137, 
    135, 125, 124, 119, 130, 127, 127, 147, 160, 112, 115, 105, 88, 76, 84, 
    94, 104, 104, 92, 95, 88, 94, 95, 94, 89, 95, 97, 103, 104, 111, 101, 96, 
    96, 92, 90, 88, 86, 85, 81, 81, 81, 87, 87, 82, 78, 90, 92, 86, 102, 109, 
    61, 141, 145, 155, 139, 138, 144, 141, 156, 158, 146, 152, 151, 151, 144, 
    151, 170, 171, 207, 215, 193, 178, 176, 175, 188, 187, 190, 193, 200, 
    193, 206, 196, 200, 202, 192, 193, 200, 187, 193, 187, 189, 182, 185, 
    181, 204, 202, 220, 203, 192, 192, 208, 207, 187, 161, 147, 175, 156, 98, 
    12, 356, 0, 159, 298, 280, 278, 284, 325, 337, 302, 303, 329, 14, 21, 13, 
    100, 157, 357, 28, 359, 160, 160, 0, 2, 0, 0, 93, 94, 94, 100, 101, 108, 
    117, 115, 138, 144, 359, 360, 346, 324, 329, 12, 107, 114, 120, 130, 137, 
    144, 140, 140, 149, 149, 150, 152, 156, 155, 158, 158, 155, 182, 137, 
    186, 206, 235, 242, 236, 217, 234, 108, 242, 341, 351, 8, 351, 333, 312, 
    301, 289, 297, 296, 344, 318, 186, 318, 328, 330, 323, 360, 4, 358, 26, 
    187, 116, 128, 119, 108, 99, 94, 93, 91, 91, 92, 89, 94, 94, 92, 88, 88, 
    91, 92, 93, 92, 93, 88, 90, 95, 94, 102, 101, 103, 94, 97, 106, 100, 116, 
    119, 105, 97, 106, 106, 105, 102, 105, 105, 109, 111, 108, 110, 106, 107, 
    109, 104, 105, 97, 91, 90, 93, 93, 90, 84, 81, 83, 85, 85, 85, 87, 88, 
    89, 87, 88, 87, 85, 87, 86, 83, 84, 90, 98, 104, 105, 96, 96, 88, 89, 92, 
    96, 99, 90, 103, 117, 120, 128, 137, 143, 148, 143, 147, 145, 142, 146, 
    146, 148, 148, 147, 142, 154, 150, 146, 137, 133, 131, 109, 121, 134, 
    133, 121, 115, 98, 96, 94, 102, 106, 109, 104, 99, 103, 105, 106, 95, 95, 
    101, 110, 121, 123, 134, 127, 109, 99, 104, 133, 137, 159, 160, 198, 227, 
    216, 172, 157, 156, 159, 173, 182, 171, 161, 150, 135, 124, 134, 152, 
    161, 170, 145, 135, 113, 116, 135, 150, 154, 147, 144, 143, 150, 152, 
    151, 139, 138, 139, 137, 135, 135, 137, 140, 137, 145, 146, 144, 143, 
    140, 138, 140, 140, 141, 138, 133, 133, 117, 129, 142, 134, 151, 151, 
    150, 143, 145, 136, 137, 128, 132, 142, 136, 132, 135, 135, 135, 134, 
    136, 138, 137, 127, 118, 115, 107, 106, 103, 97, 93, 91, 130, 125, 116, 
    127, 127, 124, 126, 112, 112, 104, 97, 98, 99, 3, 89, 89, 86, 87, 85, 92, 
    86, 86, 86, 84, 86, 85, 84, 89, 86, 83, 76, 72, 92, 80, 54, 54, 55, 40, 
    33, 33, 21, 23, 25, 19, 21, 21, 18, 26, 19, 17, 15, 14, 17, 14, 17, 16, 
    22, 16, 14, 16, 20, 20, 5, 28, 19, 25, 24, 28, 29, 33, 33, 334, 14, 40, 
    22, 25, 36, 36, 9, 10, 133, 91, 147, 149, 80, 86, 89, 87, 88, 89, 106, 
    98, 94, 85, 85, 73, 77, 86, 94, 112, 97, 65, 46, 128, 110, 90, 98, 81, 
    78, 71, 103, 111, 74, 92, 109, 94, 50, 70, 54, 13, 128, 125, 51, 47, 57, 
    128, 131, 131, 133, 144, 138, 13, 79, 129, 149, 166, 192, 193, 141, 226, 
    321, 269, 0, 153, 117, 134, 142, 132, 123, 121, 95, 142, 142, 0, 120, 
    174, 168, 149, 144, 161, 90, 88, 14, 12, 37, 32, 37, 35, 47, 32, 50, 0, 
    47, 41, 43, 4, 76, 105, 81, 71, 94, 77, 65, 47, 41, 358, 139, 118, 102, 
    99, 87, 84, 101, 94, 84, 87, 87, 102, 126, 129, 127, 151, 167, 150, 139, 
    134, 140, 141, 157, 156, 151, 154, 150, 142, 143, 141, 140, 150, 151, 
    142, 143, 140, 137, 143, 150, 147, 142, 154, 159, 154, 170, 144, 140, 
    130, 139, 133, 124, 130, 141, 137, 142, 142, 130, 120, 132, 134, 136, 
    143, 145, 144, 157, 159, 154, 149, 151, 142, 146, 157, 156, 166, 163, 
    168, 168, 168, 170, 168, 165, 174, 169, 176, 191, 169, 169, 165, 176, 
    167, 164, 175, 171, 172, 182, 194, 200, 201, 200, 195, 200, 213, 211, 
    205, 220, 229, 238, 244, 265, 270, 273, 285, 280, 289, 276, 295, 291, 
    297, 305, 297, 306, 303, 321, 316, 311, 311, 302, 295, 358, 147, 149, 
    145, 135, 129, 143, 182, 304, 4, 5, 17, 131, 128, 131, 126, 109, 86, 89, 
    96, 98, 101, 108, 114, 138, 150, 150, 147, 150, 169, 167, 170, 164, 153, 
    186, 185, 182, 178, 168, 148, 139, 159, 144, 172, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 158, 137, 143, 134, 133, 129, 122, 
    126, 128, 127, 125, 124, 128, 131, 130, 142, 154, 155, 168, 184, 190, 
    184, 182, 187, 180, 178, 181, 175, 167, 169, 168, 178, 187, 185, 195, 
    208, 166, 0, 309, 337, 318, 285, 315, 291, 299, 297, 306, 323, 354, 5, 
    152, 268, 251, 241, 258, 263, 278, 283, 274, 264, 295, 309, 300, 281, 
    276, 289, 302, 306, 295, 297, 263, 262, 262, 266, 292, 273, 278, 268, 
    276, 271, 333, 320, 319, 313, 328, 354, 349, 322, 360, 25, 16, 20, 26, 
    37, 41, 31, 46, 35, 17, 25, 28, 51, 36, 39, 32, 36, 36, 28, 25, 22, 40, 
    56, 12, 39, 72, 25, 88, 64, 46, 35, 55, 52, 47, 50, 79, 78, 37, 87, 100, 
    72, 89, 120, 130, 134, 21, 128, 147, 153, 134, 121, 127, 142, 165, 167, 
    169, 168, 175, 161, 146, 160, 148, 122, 111, 112, 113, 106, 105, 106, 
    101, 100, 95, 92, 84, 90, 89, 88, 97, 95, 95, 97, 101, 103, 104, 101, 
    102, 104, 99, 104, 103, 105, 113, 140, 135, 145, 154, 148, 143, 143, 150, 
    135, 134, 121, 117, 119, 136, 126, 71, 22, 101, 144, 135, 133, 134, 132, 
    128, 128, 125, 123, 118, 121, 107, 110, 112, 117, 112, 95, 85, 61, 112, 
    107, 110, 111, 108, 112, 139, 138, 136, 131, 100, 101, 97, 95, 95, 96, 
    100, 108, 114, 105, 101, 95, 97, 101, 108, 113, 114, 119, 123, 118, 116, 
    123, 118, 118, 118, 114, 113, 112, 114, 107, 106, 97, 106, 103, 107, 103, 
    111, 108, 105, 107, 108, 104, 105, 109, 107, 107, 110, 106, 99, 104, 105, 
    100, 106, 101, 105, 109, 117, 113, 111, 113, 113, 116, 117, 122, 117, 
    121, 126, 136, 121, 120, 120, 124, 129, 140, 143, 146, 144, 145, 134, 
    138, 133, 149, 155, 145, 144, 144, 152, 154, 156, 158, 155, 158, 152, 
    145, 146, 153, 152, 152, 149, 148, 147, 143, 144, 145, 146, 146, 142, 
    144, 145, 148, 156, 154, 161, 163, 164, 169, 168, 170, 156, 147, 156, 
    155, 153, 157, 156, 158, 158, 161, 163, 162, 161, 166, 167, 171, 175, 
    169, 169, 170, 171, 175, 178, 182, 178, 176, 184, 170, 162, 165, 169, 
    156, 171, 152, 148, 172, 156, 153, 146, 200, 226, 244, 189, 137, 357, 
    187, 173, 159, 157, 157, 202, 206, 210, 220, 233, 240, 251, 235, 244, 
    230, 238, 253, 262, 360, 6, 356, 5, 4, 360, 5, 28, 18, 18, 15, 15, 1, 5, 
    359, 355, 352, 342, 347, 340, 338, 340, 334, 336, 332, 346, 350, 352, 
    351, 350, 351, 360, 356, 347, 359, 359, 355, 348, 355, 349, 357, 350, 
    347, 346, 350, 352, 352, 352, 350, 342, 351, 346, 348, 352, 346, 341, 
    343, 346, 347, 346, 347, 347, 349, 353, 350, 348, 347, 351, 347, 354, 
    358, 355, 352, 355, 351, 360, 9, 13, 5, 11, 360, 30, 26, 37, 41, 44, 64, 
    53, 55, 74, 67, 63, 50, 48, 47, 51, 67, 54, 50, 55, 71, 89, 93, 94, 85, 
    84, 70, 56, 70, 77, 67, 77, 60, 55, 335, 355, 359, 45, 62, 63, 65, 71, 
    69, 65, 62, 58, 62, 64, 63, 205, 56, 64, 76, 76, 80, 58, 45, 50, 57, 60, 
    62, 62, 55, 50, 48, 75, 54, 49, 47, 60, 54, 59, 69, 66, 64, 72, 85, 79, 
    82, 356, 93, 9, 90, 104, 88, 95, 90, 81, 86, 93, 96, 99, 87, 108, 122, 
    114, 109, 118, 120, 134, 125, 138, 129, 118, 119, 123, 140, 123, 141, 
    140, 159, 155, 155, 157, 161, 141, 118, 122, 125, 146, 166, 156, 171, 
    162, 134, 157, 159, 141, 150, 157, 138, 140, 145, 160, 167, 145, 160, 
    157, 177, 191, 165, 148, 160, 163, 166, 154, 158, 161, 166, 159, 163, 
    150, 157, 151, 150, 149, 148, 158, 150, 165, 150, 148, 165, 161, 153, 
    149, 142, 147, 154, 152, 152, 153, 148, 156, 143, 158, 170, 166, 163, 
    163, 162, 160, 157, 137, 120, 116, 15, 41, 74, 1, 130, 91, 92, 91, 92, 
    93, 84, 82, 66, 152, 152, 153, 135, 111, 144, 134, 131, 149, 110, 108, 0, 
    65, 336, 88, 88, 94, 96, 90, 85, 106, 95, 70, 89, 62, 72, 53, 69, 26, 45, 
    32, 1, 312, 311, 307, 319, 42, 32, 45, 16, 51, 56, 48, 50, 64, 57, 52, 
    56, 45, 43, 22, 49, 65, 66, 43, 52, 119, 170, 177, 146, 134, 156, 145, 
    98, 193, 175, 141, 160, 181, 180, 156, 118, 110, 111, 125, 153, 116, 146, 
    126, 121, 125, 131, 124, 138, 137, 158, 144, 140, 137, 181, 160, 145, 
    148, 178, 166, 148, 150, 143, 152, 146, 147, 152, 160, 135, 159, 151, 
    170, 164, 56, 169, 19, 136, 43, 1, 95, 100, 110, 105, 149, 113, 104, 112, 
    113, 112, 112, 120, 137, 138, 138, 140, 136, 132, 130, 130, 136, 131, 
    129, 126, 129, 123, 120, 125, 132, 132, 125, 127, 134, 132, 135, 141, 
    141, 139, 138, 136, 135, 137, 136, 131, 129, 129, 124, 122, 118, 122, 
    118, 109, 114, 111, 108, 104, 111, 112, 114, 113, 110, 105, 100, 94, 96, 
    94, 92, 92, 90, 91, 95, 96, 96, 93, 96, 99, 104, 96, 329, 86, 83, 81, 70, 
    68, 68, 44, 48, 62, 60, 59, 59, 55, 77, 56, 53, 51, 62, 62, 55, 64, 67, 
    99, 84, 86, 92, 96, 98, 100, 99, 96, 89, 103, 85, 63, 61, 84, 82, 84, 
    107, 108, 99, 108, 89, 48, 52, 58, 61, 50, 48, 48, 59, 62, 61, 47, 42, 
    33, 292, 295, 290, 289, 288, 280, 336, 349, 354, 352, 359, 357, 356, 356, 
    357, 356, 352, 356, 359, 9, 16, 39, 16, 9, 5, 8, 7, 358, 6, 13, 17, 21, 
    14, 24, 24, 25, 25, 27, 23, 28, 12, 12, 25, 25, 28, 36, 31, 36, 37, 38, 
    25, 40, 29, 25, 24, 32, 26, 26, 28, 28, 26, 28, 28, 30, 31, 35, 35, 38, 
    35, 32, 33, 35, 41, 38, 42, 41, 41, 37, 41, 42, 39, 40, 42, 32, 36, 33, 
    34, 29, 29, 26, 30, 28, 28, 25, 28, 23, 22, 11, 12, 5, 9, 2, 356, 349, 
    337, 337, 345, 1, 8, 7, 14, 15, 15, 14, 14, 11, 10, 10, 9, 13, 5, 341, 
    329, 327, 349, 1, 3, 14, 14, 33, 34, 45, 40, 44, 42, 20, 24, 346, 338, 
    322, 344, 337, 348, 7, 14, 22, 321, 342, 332, 359, 342, 7, 18, 14, 31, 
    58, 23, 39, 65, 94, 16, 59, 62, 33, 29, 57, 46, 57, 64, 53, 79, 94, 44, 
    62, 64, 57, 8, 22, 0, 0, 55, 40, 44, 360, 337, 14, 30, 18, 16, 14, 359, 
    5, 19, 18, 13, 8, 19, 12, 27, 43, 33, 147, 158, 146, 155, 235, 11, 38, 
    65, 57, 50, 61, 77, 71, 119, 0, 0, 357, 10, 19, 32, 68, 71, 142, 74, 50, 
    20, 60, 94, 78, 75, 63, 27, 82, 0, 37, 83, 65, 68, 71, 61, 70, 87, 86, 
    85, 82, 75, 21, 75, 42, 73, 92, 77, 70, 75, 32, 1, 355, 349, 55, 55, 53, 
    62, 342, 10, 21, 31, 31, 10, 357, 38, 5, 50, 76, 69, 52, 57, 52, 40, 40, 
    47, 52, 46, 56, 27, 36, 40, 50, 64, 90, 100, 139, 99, 81, 15, 58, 53, 49, 
    52, 57, 76, 109, 90, 74, 103, 152, 57, 86, 27, 50, 83, 74, 83, 75, 87, 
    86, 84, 83, 85, 87, 85, 44, 349, 2, 10, 359, 29, 79, 75, 72, 62, 73, 70, 
    68, 42, 50, 56, 30, 22, 96, 16, 2, 230, 22, 20, 0, 0, 57, 39, 126, 94, 
    75, 109, 109, 121, 116, 108, 67, 122, 21, 74, 57, 0, 0, 0, 120, 59, 0, 
    116, 107, 115, 20, 0, 19, 113, 66, 118, 123, 103, 10, 0, 114, 0, 12, 80, 
    74, 359, 353, 56, 53, 60, 61, 57, 54, 60, 62, 346, 3, 323, 101, 45, 44, 
    44, 44, 35, 37, 26, 24, 1, 359, 360, 358, 12, 11, 17, 19, 19, 25, 16, 17, 
    16, 12, 9, 2, 6, 18, 27, 59, 21, 0, 140, 178, 121, 327, 330, 341, 336, 
    347, 339, 331, 359, 355, 350, 2, 342, 359, 349, 328, 13, 41, 23, 11, 95, 
    134, 165, 151, 152, 153, 159, 188, 147, 152, 146, 154, 159, 154, 151, 
    147, 146, 144, 139, 131, 149, 107, 120, 132, 110, 102, 337, 3, 5, 345, 
    344, 328, 343, 345, 339, 340, 338, 338, 354, 5, 4, 7, 9, 6, 241, 217, 
    178, 185, 216, 263, 281, 0, 0, 49, 45, 43, 128, 137, 137, 123, 112, 110, 
    110, 112, 122, 121, 133, 120, 134, 159, 143, 156, 153, 144, 137, 154, 
    169, 168, 163, 182, 183, 174, 174, 169, 165, 158, 143, 142, 146, 145, 
    156, 136, 359, 3, 349, 358, 328, 326, 328, 329, 317, 313, 313, 314, 327, 
    317, 347, 354, 352, 350, 351, 351, 350, 351, 358, 360, 352, 348, 356, 2, 
    358, 341, 340, 338, 336, 351, 357, 346, 353, 354, 360, 6, 21, 27, 79, 0, 
    23, 73, 56, 45, 51, 56, 58, 65, 67, 116, 26, 0, 109, 162, 225, 164, 153, 
    173, 152, 140, 140, 138, 144, 150, 141, 139, 142, 148, 146, 139, 140, 
    150, 146, 150, 165, 155, 130, 131, 122, 130, 122, 131, 143, 151, 147, 
    149, 148, 120, 116, 142, 127, 140, 163, 153, 354, 321, 323, 327, 328, 
    333, 323, 321, 318, 323, 316, 317, 320, 354, 3, 7, 1, 359, 356, 357, 356, 
    351, 343, 344, 345, 348, 355, 356, 350, 8, 9, 7, 9, 10, 12, 15, 12, 10, 
    10, 4, 357, 341, 345, 348, 360, 9, 360, 6, 5, 5, 2, 1, 1, 1, 357, 360, 1, 
    359, 356, 355, 357, 356, 351, 347, 340, 345, 7, 340, 341, 338, 349, 335, 
    342, 349, 351, 2, 360, 2, 6, 10, 7, 19, 5, 2, 16, 28, 34, 28, 28, 39, 33, 
    48, 48, 67, 78, 25, 90, 133, 185, 166, 158, 172, 148, 158, 149, 146, 124, 
    109, 113, 106, 102, 101, 93, 90, 88, 81, 88, 85, 88, 86, 83, 85, 84, 73, 
    347, 359, 3, 332, 4, 20, 29, 29, 47, 25, 0, 0, 303, 274, 263, 294, 300, 
    30, 32, 34, 27, 31, 24, 22, 30, 42, 2, 5, 331, 351, 340, 338, 349, 13, 
    27, 26, 37, 45, 42, 47, 40, 59, 57, 52, 55, 58, 65, 65, 52, 0, 356, 51, 
    64, 58, 62, 85, 110, 83, 72, 75, 75, 68, 71, 66, 59, 58, 64, 80, 81, 81, 
    81, 89, 61, 95, 90, 107, 68, 80, 114, 83, 90, 78, 4, 47, 55, 23, 90, 60, 
    97, 93, 63, 83, 3, 18, 0, 62, 130, 150, 185, 180, 166, 226, 240, 251, 
    271, 8, 29, 29, 26, 39, 49, 53, 51, 37, 29, 20, 11, 28, 55, 0, 122, 87, 
    69, 97, 62, 10, 0, 0, 0, 0, 0, 111, 125, 108, 4, 89, 91, 112, 124, 135, 
    135, 130, 126, 130, 132, 135, 145, 145, 145, 159, 151, 183, 188, 180, 
    156, 156, 162, 143, 139, 146, 152, 154, 143, 146, 130, 148, 136, 17, 0, 
    0, 0, 0, 0, 0, 0, 358, 346, 20, 13, 22, 28, 8, 16, 10, 42, 30, 29, 33, 1, 
    354, 3, 360, 7, 8, 337, 346, 355, 357, 352, 351, 360, 354, 357, 3, 1, 6, 
    8, 4, 4, 2, 4, 5, 3, 3, 3, 1, 1, 360, 358, 349, 2, 6, 10, 6, 351, 354, 8, 
    9, 348, 3, 20, 359, 11, 134, 124, 165, 135, 158, 156, 172, 160, 177, 200, 
    190, 203, 184, 180, 183, 176, 171, 173, 171, 170, 181, 146, 143, 155, 
    143, 176, 153, 151, 151, 164, 157, 163, 155, 156, 155, 152, 159, 150, 
    156, 177, 186, 194, 190, 192, 188, 185, 184, 188, 178, 182, 170, 163, 
    163, 169, 157, 161, 162, 161, 158, 149, 150, 146, 154, 154, 150, 147, 
    150, 148, 149, 156, 155, 166, 151, 156, 143, 153, 157, 155, 150, 144, 
    152, 160, 167, 159, 161, 160, 160, 153, 155, 156, 161, 150, 154, 156, 
    152, 151, 153, 153, 152, 154, 155, 158, 160, 153, 143, 140, 135, 136, 
    133, 128, 127, 132, 126, 123, 126, 126, 128, 133, 130, 128, 128, 127, 
    129, 125, 121, 125, 120, 117, 101, 316, 355, 333, 329, 330, 336, 336, 
    357, 313, 337, 169, 164, 155, 140, 138, 155, 155, 143, 151, 151, 147, 
    161, 154, 155, 152, 143, 149, 142, 150, 153, 139, 140, 137, 145, 154, 
    148, 137, 128, 117, 101, 61, 16, 346, 353, 10, 10, 313, 311, 331, 312, 
    338, 355, 177, 124, 99, 106, 121, 104, 112, 109, 105, 106, 106, 98, 99, 
    100, 100, 103, 104, 102, 105, 101, 104, 102, 108, 107, 109, 114, 111, 
    111, 117, 120, 123, 137, 188, 257, 326, 324, 295, 311, 336, 337, 327, 
    340, 308, 296, 304, 271, 350, 360, 191, 147, 118, 103, 114, 137, 135, 
    111, 100, 89, 92, 93, 81, 70, 45, 41, 26, 16, 14, 11, 9, 7, 2, 1, 4, 360, 
    358, 358, 353, 356, 9, 360, 3, 6, 1, 16, 17, 3, 5, 5, 49, 78, 145, 132, 
    139, 144, 128, 127, 132, 133, 110, 121, 113, 112, 110, 103, 90, 86, 83, 
    84, 74, 39, 39, 31, 32, 42, 35, 49, 47, 50, 64, 84, 3, 142, 191, 193, 
    193, 192, 194, 203, 207, 207, 205, 181, 222, 213, 213, 197, 214, 209, 
    237, 237, 243, 236, 252, 256, 250, 251, 261, 257, 253, 187, 39, 45, 148, 
    130, 138, 163, 117, 134, 115, 109, 95, 98, 102, 98, 95, 93, 98, 98, 95, 
    103, 113, 114, 109, 111, 111, 114, 112, 113, 114, 123, 121, 120, 125, 
    128, 124, 125, 129, 134, 135, 128, 120, 120, 116, 114, 116, 117, 120, 
    125, 126, 124, 125, 122, 119, 121, 114, 102, 105, 103, 102, 106, 105, 
    106, 102, 113, 115, 115, 118, 107, 98, 95, 109, 108, 122, 135, 134, 118, 
    116, 96, 95, 95, 101, 99, 110, 113, 108, 111, 107, 116, 111, 100, 105, 
    103, 95, 86, 85, 94, 100, 102, 92, 102, 105, 98, 98, 90, 90, 91, 100, 
    103, 107, 111, 112, 107, 109, 114, 114, 104, 24, 58, 62, 5, 98, 97, 95, 
    96, 93, 162, 323, 207, 228, 115, 82, 85, 53, 46, 36, 36, 30, 19, 36, 11, 
    16, 18, 30, 31, 20, 8, 334, 305, 287, 293, 0, 0, 0, 165, 169, 165, 150, 
    127, 132, 120, 132, 193, 169, 193, 188, 176, 179, 177, 187, 209, 232, 
    240, 257, 251, 295, 310, 315, 352, 348, 348, 349, 342, 322, 351, 295, 
    259, 271, 332, 317, 277, 277, 260, 279, 277, 280, 279, 242, 164, 152, 
    158, 151, 151, 153, 150, 139, 132, 132, 134, 153, 141, 130, 122, 124, 
    121, 118, 114, 126, 156, 141, 143, 134, 138, 133, 133, 113, 130, 142, 
    214, 337, 351, 352, 343, 345, 347, 343, 351, 357, 360, 337, 337, 331, 
    358, 4, 9, 4, 340, 1, 6, 4, 7, 359, 360, 5, 1, 355, 358, 357, 342, 342, 
    341, 349, 337, 329, 328, 313, 314, 316, 318, 335, 329, 322, 332, 331, 
    326, 328, 329, 333, 316, 319, 303, 294, 254, 196, 184, 148, 152, 150, 
    151, 133, 132, 133, 106, 105, 106, 109, 113, 104, 102, 102, 120, 135, 
    124, 120, 118, 111, 104, 97, 102, 106, 111, 113, 112, 100, 100, 105, 137, 
    136, 130, 141, 118, 127, 147, 141, 130, 129, 163, 131, 120, 116, 134, 
    359, 130, 30, 2, 165, 42, 206, 356, 214, 21, 233, 0, 0, 58, 11, 338, 355, 
    340, 285, 346, 19, 358, 273, 172, 160, 155, 151, 144, 146, 168, 150, 144, 
    161, 172, 196, 170, 153, 147, 132, 128, 153, 148, 155, 161, 154, 148, 
    152, 158, 148, 144, 140, 137, 138, 134, 135, 130, 132, 132, 134, 139, 
    139, 131, 127, 127, 126, 125, 121, 131, 131, 131, 131, 123, 119, 120, 
    122, 121, 132, 146, 154, 153, 152, 142, 142, 143, 149, 146, 148, 148, 
    155, 157, 159, 155, 157, 158, 158, 155, 151, 148, 147, 137, 124, 116, 95, 
    98, 107, 105, 115, 118, 120, 124, 127, 131, 137, 142, 143, 142, 120, 110, 
    108, 106, 103, 98, 98, 107, 116, 110, 116, 117, 119, 123, 112, 135, 128, 
    117, 121, 122, 118, 82, 91, 94, 98, 95, 86, 93, 80, 88, 82, 62, 58, 20, 
    4, 30, 25, 24, 26, 22, 29, 28, 24, 19, 20, 10, 22, 11, 13, 8, 19, 8, 10, 
    11, 12, 12, 8, 9, 12, 11, 8, 16, 23, 15, 19, 15, 15, 13, 16, 15, 20, 18, 
    14, 18, 17, 16, 16, 34, 29, 20, 19, 28, 22, 11, 11, 11, 18, 12, 10, 9, 
    11, 4, 2, 351, 358, 356, 354, 350, 347, 341, 341, 337, 336, 339, 343, 
    342, 343, 344, 342, 340, 335, 333, 332, 331, 328, 332, 341, 328, 320, 
    323, 326, 326, 327, 318, 336, 328, 327, 325, 324, 317, 320, 328, 325, 
    315, 310, 306, 314, 321, 313, 327, 331, 4, 341, 351, 340, 334, 332, 342, 
    340, 335, 333, 333, 332, 340, 340, 347, 347, 339, 335, 335, 348, 348, 
    353, 3, 355, 351, 15, 21, 11, 360, 356, 358, 11, 9, 27, 9, 354, 5, 12, 
    20, 9, 14, 14, 6, 11, 9, 11, 3, 7, 8, 8, 2, 4, 357, 8, 3, 1, 353, 360, 
    359, 360, 359, 5, 6, 6, 7, 9, 4, 67, 80, 46, 2, 84, 34, 349, 41, 30, 22, 
    25, 9, 9, 9, 5, 355, 9, 5, 359, 90, 359, 63, 21, 347, 351, 87, 88, 357, 
    345, 0, 354, 122, 354, 76, 101, 86, 62, 72, 85, 91, 90, 90, 96, 82, 104, 
    128, 149, 155, 154, 153, 150, 153, 159, 146, 150, 151, 154, 156, 151, 
    159, 160, 166, 154, 152, 144, 131, 130, 134, 141, 152, 156, 166, 161, 
    161, 147, 163, 157, 161, 155, 163, 150, 145, 108, 108, 120, 109, 111, 
    107, 120, 130, 136, 126, 128, 131, 122, 116, 120, 116, 111, 113, 120, 
    122, 123, 120, 109, 111, 107, 110, 120, 126, 123, 123, 126, 126, 131, 
    132, 124, 130, 131, 117, 113, 118, 117, 110, 112, 124, 125, 124, 138, 
    143, 138, 138, 137, 142, 145, 153, 147, 145, 151, 159, 156, 154, 358, 
    156, 354, 337, 186, 0, 10, 358, 347, 339, 319, 311, 360, 344, 10, 0, 183, 
    194, 158, 164, 178, 152, 156, 152, 132, 119, 125, 119, 129, 137, 124, 
    128, 140, 130, 123, 124, 125, 131, 126, 131, 123, 121, 115, 109, 104, 
    104, 106, 108, 108, 111, 113, 120, 123, 112, 133, 113, 119, 120, 136, 
    145, 155, 154, 153, 150, 151, 157, 155, 154, 157, 106, 350, 5, 8, 350, 3, 
    333, 340, 354, 353, 358, 0, 0, 352, 342, 7, 1, 4, 174, 353, 181, 176, 0, 
    0, 0, 0, 0, 0, 2, 347, 0, 167, 146, 330, 195, 189, 300, 325, 356, 169, 
    15, 9, 302, 0, 360, 96, 111, 132, 133, 128, 130, 143, 12, 95, 10, 351, 
    348, 162, 358, 348, 344, 310, 343, 358, 331, 12, 338, 323, 173, 30, 54, 
    28, 1, 8, 248, 94, 92, 30, 246, 337, 43, 349, 70, 12, 84, 90, 106, 100, 
    102, 96, 94, 90, 92, 88, 88, 87, 87, 88, 303, 291, 353, 69, 312, 87, 64, 
    323, 4, 4, 360, 356, 7, 15, 14, 356, 339, 298, 340, 60, 0, 260, 30, 3, 
    360, 318, 0, 358, 357, 8, 347, 9, 5, 355, 352, 355, 265, 229, 204, 234, 
    166, 143, 145, 129, 157, 15, 343, 3, 353, 359, 14, 359, 354, 6, 6, 350, 
    2, 2, 26, 5, 360, 2, 360, 359, 359, 346, 344, 341, 347, 355, 350, 350, 
    338, 346, 345, 348, 360, 4, 355, 1, 355, 353, 350, 348, 346, 344, 340, 
    337, 337, 340, 341, 348, 341, 343, 346, 343, 343, 335, 331, 337, 338, 
    337, 342, 353, 347, 347, 340, 335, 334, 336, 341, 334, 335, 340, 340, 
    341, 341, 340, 344, 342, 346, 353, 346, 356, 356, 354, 351, 346, 347, 
    340, 336, 337, 331, 333, 334, 337, 340, 341, 320, 320, 319, 313, 312, 
    313, 304, 305, 302, 303, 309, 311, 313, 324, 321, 315, 310, 319, 330, 
    323, 314, 325, 319, 323, 324, 316, 329, 330, 335, 347, 335, 334, 338, 
    338, 338, 342, 341, 341, 340, 335, 346, 345, 338, 341, 317, 325, 321, 
    322, 326, 323, 323, 322, 320, 314, 318, 321, 330, 339, 338, 334, 339, 
    344, 344, 344, 339, 334, 341, 337, 342, 337, 331, 333, 340, 333, 352, 
    345, 342, 344, 346, 341, 350, 350, 346, 11, 15, 357, 360, 2, 4, 357, 346, 
    359, 354, 336, 339, 341, 356, 355, 346, 1, 353, 351, 330, 1, 356, 344, 
    351, 358, 319, 50, 354, 326, 339, 320, 317, 340, 351, 320, 0, 358, 321, 
    355, 182, 143, 163, 159, 161, 159, 153, 159, 149, 150, 176, 178, 121, 
    345, 353, 338, 322, 13, 181, 121, 120, 153, 171, 126, 121, 128, 148, 124, 
    124, 117, 132, 154, 159, 147, 126, 138, 147, 145, 147, 153, 158, 151, 
    147, 146, 143, 145, 141, 140, 138, 137, 142, 137, 140, 151, 157, 162, 
    157, 155, 159, 157, 142, 146, 147, 148, 148, 148, 151, 151, 147, 157, 
    152, 152, 165, 151, 144, 146, 150, 155, 159, 160, 145, 150, 165, 148, 
    143, 153, 162, 167, 169, 327, 1, 337, 334, 132, 141, 164, 150, 139, 151, 
    151, 157, 151, 158, 153, 153, 161, 172, 178, 167, 149, 150, 168, 160, 
    155, 145, 148, 142, 163, 136, 241, 217, 174, 146, 146, 136, 142, 162, 
    175, 338, 314, 6, 6, 7, 360, 352, 359, 328, 272, 199, 185, 151, 176, 194, 
    321, 356, 55, 51, 187, 336, 5, 166, 165, 101, 97, 110, 122, 120, 116, 
    117, 112, 110, 133, 143, 151, 151, 154, 157, 151, 159, 149, 160, 169, 
    149, 12, 287, 1, 345, 359, 316, 327, 315, 329, 308, 278, 279, 306, 304, 
    272, 311, 306, 326, 316, 343, 39, 351, 161, 148, 155, 147, 152, 151, 162, 
    160, 157, 154, 152, 159, 131, 131, 122, 141, 133, 132, 170, 330, 334, 
    358, 15, 17, 358, 1, 354, 341, 2, 357, 355, 356, 349, 343, 341, 230, 174, 
    118, 102, 100, 101, 102, 102, 103, 105, 109, 105, 99, 102, 100, 96, 102, 
    103, 101, 99, 114, 148, 152, 153, 175, 178, 189, 337, 342, 346, 347, 358, 
    347, 348, 347, 341, 351, 341, 345, 349, 348, 350, 3, 13, 18, 9, 7, 359, 
    12, 354, 7, 344, 330, 328, 206, 200, 196, 186, 179, 175, 206, 180, 185, 
    239, 298, 355, 6, 23, 346, 253, 305, 343, 318, 292, 247, 226, 193, 183, 
    176, 172, 189, 170, 168, 154, 150, 150, 150, 151, 153, 152, 156, 158, 
    152, 155, 161, 148, 144, 163, 154, 149, 157, 158, 168, 152, 127, 130, 
    138, 119, 118, 131, 143, 144, 138, 144, 144, 148, 151, 153, 153, 166, 
    149, 214, 203, 218, 232, 171, 155, 192, 166, 160, 148, 146, 174, 158, 
    185, 154, 150, 138, 205, 168, 107, 166, 13, 357, 233, 354, 347, 2, 22, 
    351, 8, 12, 12, 5, 360, 0, 352, 329, 4, 33, 2, 337, 304, 345, 16, 355, 9, 
    327, 348, 239, 105, 119, 130, 144, 123, 141, 120, 107, 124, 106, 103, 
    110, 108, 111, 106, 146, 273, 100, 91, 81, 82, 266, 342, 89, 85, 76, 81, 
    81, 100, 236, 142, 81, 345, 12, 167, 358, 98, 354, 327, 341, 356, 321, 0, 
    227, 20, 10, 0, 357, 243, 99, 110, 111, 120, 130, 134, 145, 145, 144, 
    155, 153, 167, 163, 166, 159, 277, 330, 335, 309, 315, 328, 347, 14, 3, 
    20, 37, 223, 178, 169, 160, 122, 123, 118, 123, 113, 111, 125, 123, 123, 
    117, 139, 131, 133, 154, 150, 153, 158, 166, 166, 161, 218, 139, 176, 
    216, 200, 130, 360, 10, 24, 27, 24, 7, 156, 138, 124, 130, 216, 145, 190, 
    180, 196, 240, 342, 304, 291, 285, 319, 319, 237, 172, 172, 156, 145, 
    139, 155, 152, 164, 150, 164, 147, 153, 156, 155, 171, 202, 177, 196, 
    176, 153, 156, 180, 107, 12, 19, 3, 26, 4, 2, 338, 6, 360, 335, 8, 12, 6, 
    22, 111, 257, 59, 190, 22, 289, 300, 331, 329, 332, 333, 331, 328, 334, 
    333, 321, 318, 323, 329, 328, 334, 332, 340, 339, 336, 338, 44, 341, 8, 
    242, 345, 189, 165, 162, 151, 153, 154, 180, 167, 170, 177, 185, 175, 
    171, 154, 156, 158, 178, 175, 169, 158, 153, 167, 158, 147, 143, 141, 
    144, 140, 139, 149, 149, 147, 162, 168, 159, 156, 176, 138, 182, 339, 1, 
    15, 347, 33, 348, 319, 357, 1, 355, 85, 87, 86, 86, 60, 98, 91, 83, 90, 
    93, 91, 100, 125, 100, 98, 93, 97, 94, 100, 116, 121, 121, 122, 124, 133, 
    144, 159, 142, 152, 147, 154, 157, 152, 152, 149, 155, 143, 153, 149, 
    148, 148, 152, 154, 166, 158, 168, 164, 168, 169, 164, 155, 151, 170, 
    169, 165, 160, 150, 151, 161, 154, 148, 148, 153, 157, 145, 158, 143, 
    141, 149, 194, 220, 226, 314, 314, 346, 340, 306, 219, 152, 3, 79, 90, 
    83, 89, 91, 90, 91, 48, 58, 21, 31, 6, 358, 7, 5, 19, 355, 47, 13, 6, 12, 
    352, 7, 10, 8, 8, 5, 3, 3, 9, 353, 5, 349, 7, 360, 9, 11, 8, 4, 14, 19, 
    18, 6, 8, 358, 3, 357, 358, 354, 1, 6, 6, 356, 5, 4, 7, 10, 7, 4, 4, 2, 
    2, 6, 9, 4, 350, 14, 174, 315, 81, 337, 333, 157, 40, 76, 299, 30, 360, 
    344, 25, 29, 38, 46, 50, 67, 7, 18, 14, 346, 15, 15, 16, 13, 16, 13, 28, 
    7, 10, 2, 4, 359, 360, 345, 343, 9, 324, 315, 337, 309, 304, 227, 211, 
    204, 201, 197, 238, 259, 319, 6, 346, 346, 355, 354, 9, 358, 347, 347, 3, 
    14, 4, 16, 24, 10, 7, 9, 8, 12, 7, 3, 3, 5, 16, 9, 5, 7, 10, 7, 9, 10, 
    11, 10, 9, 8, 9, 9, 9, 11, 11, 7, 2, 10, 5, 27, 322, 1, 351, 4, 10, 12, 
    10, 11, 9, 5, 5, 5, 7, 7, 8, 8, 4, 9, 7, 9, 9, 12, 2, 7, 16, 8, 15, 359, 
    350, 4, 6, 7, 8, 6, 6, 7, 6, 5, 3, 2, 360, 355, 356, 358, 2, 1, 6, 3, 
    358, 1, 358, 356, 353, 356, 352, 354, 3, 355, 355, 356, 357, 1, 1, 360, 
    2, 8, 5, 4, 2, 3, 7, 9, 8, 5, 13, 4, 12, 49, 356, 353, 356, 20, 43, 36, 
    356, 5, 6, 30, 5, 1, 315, 52, 50, 14, 357, 360, 119, 116, 357, 309, 206, 
    63, 93, 354, 342, 352, 2, 1, 121, 295, 235, 334, 147, 223, 307, 333, 247, 
    17, 89, 41, 16, 23, 97, 96, 103, 96, 109, 134, 150, 198, 98, 94, 107, 
    144, 147, 145, 145, 160, 156, 163, 159, 153, 152, 143, 144, 124, 135, 
    144, 142, 99, 100, 101, 101, 100, 98, 95, 91, 97, 101, 103, 108, 111, 
    121, 150, 156, 154, 146, 137, 129, 129, 124, 129, 123, 125, 118, 103, 
    106, 99, 103, 109, 116, 117, 114, 125, 124, 125, 129, 135, 143, 137, 127, 
    126, 123, 116, 106, 91, 94, 98, 106, 107, 115, 117, 103, 107, 100, 90, 
    96, 90, 85, 86, 83, 78, 77, 79, 78, 76, 70, 61, 60, 48, 33, 23, 21, 20, 
    19, 16, 15, 17, 13, 9, 10, 10, 5, 360, 359, 352, 350, 347, 345, 344, 343, 
    343, 341, 337, 332, 333, 333, 330, 330, 326, 324, 336, 334, 326, 334, 
    328, 311, 305, 309, 306, 315, 351, 270, 263, 282, 260, 254, 283, 320, 
    328, 250, 215, 269, 0, 0, 351, 151, 350, 326, 3, 343, 6, 352, 356, 355, 
    356, 360, 11, 21, 9, 3, 11, 16, 17, 12, 4, 1, 5, 8, 355, 360, 351, 355, 
    357, 8, 360, 3, 360, 358, 360, 4, 7, 8, 7, 3, 3, 3, 5, 360, 6, 3, 10, 10, 
    1, 8, 12, 11, 15, 16, 12, 8, 25, 38, 44, 36, 43, 41, 29, 331, 33, 41, 25, 
    30, 37, 18, 18, 22, 23, 13, 14, 13, 10, 13, 6, 4, 7, 5, 355, 343, 344, 
    338, 341, 341, 332, 348, 346, 348, 347, 360, 15, 17, 289, 264, 255, 244, 
    223, 230, 283, 109, 0, 234, 195, 107, 114, 11, 5, 0, 8, 84, 21, 0, 43, 
    88, 87, 92, 84, 23, 11, 360, 28, 5, 4, 7, 355, 2, 57, 319, 0, 267, 110, 
    144, 312, 263, 267, 290, 135, 154, 163, 147, 145, 154, 152, 152, 155, 
    165, 157, 155, 171, 187, 162, 188, 181, 170, 170, 160, 156, 147, 157, 
    150, 148, 147, 135, 134, 132, 130, 117, 120, 121, 117, 117, 133, 129, 
    160, 150, 144, 145, 132, 139, 149, 153, 173, 159, 149, 147, 119, 146, 
    156, 143, 161, 183, 162, 216, 242, 256, 235, 257, 288, 284, 278, 291, 
    289, 285, 300, 314, 312, 307, 308, 307, 309, 318, 309, 307, 324, 315, 
    321, 318, 259, 234, 225, 215, 122, 134, 125, 117, 113, 126, 120, 111, 
    107, 109, 108, 127, 145, 156, 157, 156, 163, 151, 159, 155, 138, 127, 
    148, 136, 133, 128, 150, 155, 170, 166, 156, 182, 176, 145, 134, 161, 
    200, 265, 273, 273, 263, 269, 286, 263, 318, 337, 213, 295, 9, 13, 89, 
    81, 21, 30, 17, 19, 17, 12, 15, 11, 8, 6, 6, 10, 349, 10, 3, 321, 333, 
    20, 342, 338, 321, 318, 357, 13, 285, 29, 152, 165, 165, 161, 222, 246, 
    254, 277, 287, 352, 315, 332, 299, 11, 182, 163, 163, 155, 156, 171, 167, 
    152, 146, 155, 146, 152, 155, 167, 170, 181, 100, 88, 98, 0, 6, 344, 7, 
    358, 333, 332, 343, 351, 352, 341, 350, 338, 338, 327, 332, 334, 308, 
    304, 327, 331, 335, 335, 334, 345, 338, 315, 309, 263, 234, 255, 222, 
    206, 220, 226, 213, 191, 153, 143, 98, 6, 51, 5, 0, 0, 296, 242, 274, 
    266, 280, 0, 183, 222, 202, 182, 163, 144, 154, 147, 146, 159, 157, 159, 
    156, 160, 153, 152, 155, 166, 174, 340, 45, 0, 84, 21, 219, 212, 122, 
    190, 266, 274, 307, 304, 330, 323, 308, 337, 334, 328, 332, 338, 340, 
    344, 348, 342, 4, 9, 3, 1, 14, 34, 16, 358, 6, 357, 4, 0, 236, 329, 85, 
    3, 0, 281, 105, 116, 100, 91, 90, 86, 91, 115, 156, 150, 138, 149, 136, 
    115, 131, 124, 156, 161, 140, 141, 141, 147, 143, 129, 117, 120, 117, 
    108, 146, 134, 106, 118, 114, 113, 107, 93, 90, 76, 65, 77, 70, 62, 65, 
    45, 40, 34, 6, 358, 346, 359, 345, 348, 336, 329, 329, 325, 319, 321, 
    319, 323, 318, 318, 315, 316, 325, 318, 342, 329, 329, 330, 336, 346, 
    336, 321, 328, 340, 309, 307, 319, 332, 314, 344, 340, 339, 336, 333, 
    332, 335, 328, 333, 345, 353, 346, 343, 332, 335, 0, 115, 123, 115, 123, 
    112, 106, 106, 108, 116, 117, 117, 117, 119, 114, 111, 99, 100, 129, 114, 
    117, 118, 125, 123, 122, 124, 127, 128, 125, 119, 106, 108, 118, 117, 
    103, 101, 101, 106, 116, 100, 98, 95, 100, 111, 106, 106, 91, 74, 88, 90, 
    106, 110, 111, 108, 118, 108, 95, 83, 89, 57, 52, 69, 56, 24, 23, 14, 51, 
    71, 65, 63, 63, 55, 26, 29, 10, 49, 28, 66, 54, 57, 41, 42, 83, 25, 61, 
    65, 51, 65, 47, 23, 28, 321, 284, 328, 318, 3, 34, 35, 39, 35, 28, 31, 
    34, 11, 334, 55, 87, 11, 13, 341, 2, 355, 16, 20, 16, 5, 15, 249, 57, 38, 
    54, 44, 40, 47, 35, 52, 48, 60, 64, 32, 30, 18, 33, 20, 10, 9, 6, 314, 
    50, 71, 41, 43, 38, 62, 44, 61, 40, 35, 47, 53, 52, 51, 41, 47, 50, 52, 
    61, 50, 64, 59, 57, 43, 37, 54, 33, 40, 49, 51, 40, 42, 45, 48, 60, 61, 
    51, 59, 59, 64, 65, 57, 54, 48, 40, 42, 47, 64, 68, 76, 73, 65, 64, 60, 
    60, 68, 58, 57, 62, 60, 60, 70, 66, 74, 84, 88, 83, 91, 81, 83, 91, 83, 
    84, 87, 88, 90, 98, 105, 107, 104, 100, 96, 105, 116, 111, 110, 103, 99, 
    95, 101, 98, 103, 96, 94, 92, 106, 96, 101, 119, 110, 117, 113, 114, 115, 
    115, 118, 124, 123, 125, 125, 131, 136, 132, 126, 132, 127, 129, 128, 
    126, 120, 108, 104, 117, 5, 4, 307, 310, 303, 313, 312, 320, 326, 321, 
    327, 327, 331, 336, 335, 345, 331, 337, 344, 348, 344, 349, 343, 346, 
    347, 345, 347, 347, 355, 343, 355, 343, 341, 338, 344, 337, 328, 325, 
    313, 308, 303, 302, 295, 286, 280, 291, 279, 282, 289, 284, 269, 271, 
    265, 261, 269, 256, 263, 259, 267, 273, 277, 286, 252, 245, 258, 262, 
    148, 123, 196, 195, 163, 202, 191, 203, 208, 184, 220, 205, 206, 199, 
    200, 143, 142, 141, 192, 188, 143, 125, 117, 110, 106, 104, 81, 76, 80, 
    73, 60, 45, 49, 41, 35, 37, 40, 28, 359, 358, 345, 345, 337, 326, 329, 
    345, 352, 348, 346, 358, 341, 333, 343, 343, 350, 346, 344, 356, 355, 
    352, 351, 354, 342, 345, 351, 355, 354, 351, 350, 349, 348, 344, 340, 1, 
    359, 6, 7, 5, 3, 5, 5, 5, 11, 8, 16, 16, 16, 15, 9, 8, 10, 21, 20, 30, 
    15, 17, 16, 19, 9, 12, 15, 20, 28, 14, 21, 23, 22, 21, 16, 26, 27, 18, 
    16, 20, 25, 31, 27, 19, 18, 18, 18, 17, 23, 22, 30, 21, 17, 15, 8, 9, 11, 
    7, 7, 10, 10, 26, 35, 28, 14, 1, 20, 34, 15, 20, 19, 358, 40, 4, 4, 2, 
    345, 353, 348, 347, 4, 360, 311, 279, 265, 261, 245, 255, 210, 206, 203, 
    198, 188, 181, 166, 150, 153, 160, 147, 136, 151, 151, 145, 138, 143, 
    134, 135, 133, 122, 121, 144, 133, 122, 121, 124, 127, 125, 102, 97, 82, 
    85, 86, 76, 72, 64, 59, 46, 40, 33, 24, 26, 22, 22, 18, 16, 19, 10, 14, 
    12, 10, 13, 12, 12, 14, 10, 5, 3, 355, 351, 343, 345, 346, 349, 340, 350, 
    340, 342, 345, 332, 322, 322, 327, 330, 330, 325, 315, 307, 330, 330, 
    332, 345, 346, 323, 266, 241, 147, 220, 233, 251, 252, 232, 227, 222, 
    221, 210, 202, 198, 162, 148, 182, 125, 159, 164, 155, 188, 156, 170, 
    136, 136, 122, 104, 75, 42, 13, 40, 46, 34, 26, 351, 342, 339, 340, 341, 
    342, 342, 336, 342, 343, 340, 349, 346, 339, 344, 347, 350, 350, 348, 
    350, 350, 347, 353, 349, 350, 348, 351, 352, 354, 359, 359, 2, 360, 358, 
    349, 345, 351, 358, 23, 53, 123, 191, 228, 195, 160, 174, 176, 168, 172, 
    185, 175, 190, 183, 229, 260, 275, 85, 14, 32, 35, 50, 64, 37, 50, 125, 
    131, 117, 111, 108, 113, 120, 124, 135, 134, 151, 146, 147, 156, 168, 
    146, 151, 154, 157, 149, 147, 146, 146, 145, 141, 138, 132, 133, 133, 
    132, 134, 133, 137, 133, 132, 130, 128, 130, 133, 126, 124, 125, 127, 
    130, 131, 127, 126, 122, 120, 116, 116, 128, 131, 127, 124, 123, 121, 
    121, 124, 131, 123, 118, 125, 119, 110, 121, 127, 111, 124, 120, 129, 
    132, 125, 129, 129, 133, 133, 130, 134, 129, 136, 126, 130, 131, 134, 
    122, 108, 104, 113, 117, 126, 139, 109, 117, 115, 110, 107, 99, 90, 90, 
    93, 98, 101, 98, 96, 99, 109, 112, 118, 133, 123, 149, 132, 128, 123, 
    128, 132, 134, 143, 137, 122, 139, 123, 116, 104, 102, 101, 94, 107, 104, 
    100, 117, 149, 152, 147, 165, 171, 170, 170, 118, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, 152, 161, 166, 157, 158, 153, 146, 145, 148, 149, 146, 139, 136, 
    131, 126, 124, 122, 121, 117, 117, 114, 121, 122, 123, 121, 120, 123, 
    126, 129, 130, 128, 117, 119, 118, 117, 119, 116, 112, 110, 111, 111, 
    114, 114, 113, 122, 123, 117, 132, 119, 116, 115, 101, 102, 90, 89, 85, 
    68, 73, 95, 79, 109, 84, 106, 98, 78, 69, 76, 68, 73, 77, 79, 73, 70, 55, 
    349, 7, 360, 359, 25, 56, 68, 66, 70, 71, 68, 61, 62, 71, 67, 64, 59, 57, 
    58, 58, 65, 63, 67, 66, 60, 58, 68, 77, 70, 69, 75, 84, 62, 66, 53, 50, 
    58, 54, 58, 64, 63, 57, 60, 57, 57, 43, 45, 46, 40, 48, 34, 35, 37, 26, 
    19, 9, 4, 1, 359, 352, 347, 345, 360, 4, 358, 360, 8, 8, 7, 15, 13, 4, 5, 
    5, 360, 355, 1, 352, 1, 354, 353, 360, 354, 354, 359, 357, 356, 360, 356, 
    358, 355, 348, 352, 359, 352, 2, 354, 343, 355, 17, 89, 77, 89, 110, 123, 
    112, 112, 108, 107, 141, 195, 164, 160, 173, 162, 159, 159, 158, 152, 
    145, 138, 133, 132, 146, 162, 163, 154, 161, 153, 158, 153, 159, 158, 
    171, 160, 150, 0, 0, 336, 325, 320, 328, 320, 314, 335, 353, 349, 353, 
    343, 360, 349, 1, 358, 350, 334, 6, 338, 281, 273, 274, 102, 125, 127, 
    138, 133, 135, 162, 154, 144, 157, 158, 163, 161, 161, 164, 159, 157, 
    168, 170, 176, 168, 169, 173, 195, 267, 331, 360, 347, 360, 27, 30, 17, 
    13, 5, 1, 351, 359, 15, 20, 10, 23, 31, 18, 41, 360, 324, 340, 347, 313, 
    311, 315, 323, 255, 259, 342, 338, 344, 343, 341, 357, 354, 2, 356, 350, 
    2, 356, 6, 4, 347, 340, 360, 349, 5, 4, 23, 28, 6, 52, 95, 106, 113, 53, 
    54, 27, 139, 78, 118, 154, 132, 132, 124, 124, 126, 152, 141, 113, 105, 
    106, 116, 145, 139, 133, 151, 159, 126, 115, 117, 122, 133, 129, 131, 
    144, 120, 127, 120, 115, 113, 107, 92, 100, 99, 106, 103, 102, 106, 102, 
    101, 84, 84, 71, 54, 60, 56, 54, 51, 45, 41, 42, 26, 51, 61, 60, 60, 62, 
    54, 51, 49, 64, 60, 58, 58, 65, 62, 65, 70, 62, 66, 59, 64, 63, 47, 47, 
    77, 74, 73, 65, 55, 50, 74, 62, 65, 87, 90, 116, 121, 117, 116, 110, 126, 
    118, 128, 105, 103, 109, 121, 127, 125, 123, 130, 134, 138, 142, 145, 
    146, 148, 151, 151, 161, 160, 163, 167, 173, 168, 175, 168, 177, 183, 
    188, 181, 181, 183, 198, 193, 196, 200, 199, 199, 205, 201, 202, 205, 
    204, 217, 218, 217, 216, 211, 208, 212, 213, 216, 218, 219, 215, 219, 
    219, 217, 224, 219, 219, 227, 225, 220, 208, 200, 168, 182, 154, 152, 
    150, 155, 153, 159, 136, 139, 121, 116, 108, 102, 102, 102, 102, 97, 95, 
    90, 87, 85, 91, 92, 92, 91, 90, 91, 85, 81, 84, 90, 99, 130, 150, 118, 
    112, 134, 134, 134, 336, 331, 330, 306, 323, 312, 305, 295, 287, 286, 
    295, 288, 284, 287, 287, 281, 287, 285, 298, 292, 337, 338, 347, 345, 
    339, 10, 356, 13, 9, 359, 4, 6, 9, 13, 5, 359, 3, 355, 354, 2, 3, 354, 4, 
    353, 10, 8, 356, 20, 358, 28, 45, 59, 43, 44, 341, 290, 72, 351, 77, 120, 
    148, 174, 168, 166, 170, 188, 190, 218, 222, 232, 225, 221, 220, 221, 
    218, 220, 219, 237, 258, 274, 291, 23, 18, 9, 10, 12, 6, 356, 339, 344, 
    344, 347, 344, 354, 358, 2, 10, 20, 7, 3, 10, 8, 356, 2, 1, 354, 359, 3, 
    357, 358, 7, 7, 11, 31, 35, 80, 101, 142, 126, 119, 115, 117, 116, 114, 
    122, 111, 128, 293, 270, 242, 249, 287, 281, 291, 292, 321, 309, 202, 
    246, 275, 286, 269, 270, 272, 279, 245, 223, 224, 222, 226, 224, 215, 
    207, 201, 220, 225, 224, 221, 234, 239, 120, 210, 106, 330, 279, 286, 
    295, 2, 3, 228, 148, 153, 94, 99, 91, 88, 86, 84, 87, 88, 88, 42, 102, 
    168, 309, 308, 305, 46, 65, 41, 34, 27, 17, 5, 4, 351, 357, 350, 345, 
    347, 351, 347, 346, 343, 345, 348, 349, 342, 354, 348, 354, 358, 350, 
    346, 350, 352, 343, 356, 345, 342, 350, 347, 351, 352, 344, 347, 353, 
    351, 350, 349, 350, 358, 351, 356, 360, 355, 360, 355, 2, 4, 8, 12, 359, 
    356, 357, 10, 355, 9, 7, 6, 20, 38, 23, 14, 23, 21, 53, 62, 81, 90, 91, 
    86, 91, 97, 124, 131, 111, 109, 118, 118, 125, 131, 107, 100, 83, 57, 64, 
    58, 38, 50, 67, 59, 48, 52, 43, 31, 35, 37, 40, 54, 51, 68, 64, 57, 55, 
    49, 51, 51, 46, 70, 76, 64, 61, 59, 60, 57, 44, 46, 47, 53, 54, 53, 81, 
    88, 97, 85, 74, 80, 55, 53, 79, 82, 68, 60, 58, 57, 64, 59, 54, 55, 60, 
    58, 54, 52, 34, 50, 56, 57, 55, 65, 68, 69, 82, 78, 90, 79, 65, 93, 132, 
    131, 107, 113, 127, 135, 133, 112, 94, 44, 41, 41, 43, 45, 59, 54, 65, 
    80, 108, 110, 107, 100, 108, 112, 116, 134, 122, 116, 116, 122, 131, 137, 
    134, 135, 137, 145, 128, 117, 122, 122, 122, 128, 128, 128, 130, 137, 
    135, 133, 130, 126, 136, 127, 123, 120, 119, 109, 110, 115, 113, 114, 
    110, 109, 108, 103, 103, 102, 100, 90, 102, 99, 92, 71, 115, 109, 104, 
    95, 106, 96, 102, 96, 94, 104, 102, 105, 107, 92, 94, 102, 104, 102, 100, 
    106, 106, 103, 107, 103, 109, 109, 111, 112, 103, 105, 112, 103, 115, 
    110, 107, 106, 100, 107, 104, 106, 103, 105, 110, 112, 114, 110, 105, 
    105, 107, 102, 98, 99, 97, 98, 97, 95, 93, 87, 90, 95, 82, 82, 94, 94, 
    95, 98, 95, 97, 97, 94, 97, 89, 75, 73, 64, 60, 40, 30, 17, 27, 27, 26, 
    20, 25, 21, 15, 17, 15, 18, 24, 22, 33, 34, 34, 37, 48, 60, 67, 83, 82, 
    55, 68, 83, 89, 85, 86, 85, 88, 90, 97, 109, 114, 121, 119, 107, 98, 92, 
    92, 91, 87, 88, 94, 96, 100, 92, 97, 96, 102, 99, 107, 109, 121, 129, 
    114, 134, 130, 125, 121, 115, 137, 138, 144, 155, 150, 150, 153, 153, 
    156, 156, 154, 155, 152, 151, 151, 153, 147, 147, 154, 163, 159, 177, 
    150, 158, 160, 149, 141, 154, 164, 161, 161, 150, 133, 116, 100, 100, 
    126, 130, 123, 109, 103, 104, 109, 112, 101, 105, 106, 106, 99, 97, 98, 
    97, 112, 108, 106, 98, 91, 91, 96, 99, 95, 99, 75, 85, 87, 82, 74, 78, 
    78, 55, 46, 58, 58, 55, 57, 60, 72, 76, 79, 66, 74, 66, 71, 56, 66, 67, 
    61, 34, 51, 36, 37, 359, 347, 333, 348, 347, 348, 349, 341, 334, 344, 
    350, 346, 346, 341, 343, 341, 335, 330, 324, 320, 314, 325, 324, 334, 
    334, 334, 341, 329, 315, 327, 323, 331, 332, 325, 321, 323, 337, 330, 
    328, 333, 320, 321, 311, 271, 273, 280, 284, 283, 287, 342, 309, 289, 
    290, 303, 325, 326, 359, 259, 256, 227, 233, 239, 249, 258, 274, 278, 
    320, 333, 330, 330, 333, 332, 335, 331, 332, 334, 325, 328, 329, 337, 
    336, 327, 327, 325, 323, 322, 320, 285, 280, 200, 195, 166, 218, 219, 
    208, 183, 151, 137, 150, 149, 142, 126, 127, 110, 102, 92, 101, 96, 92, 
    94, 94, 96, 94, 94, 99, 106, 114, 107, 113, 105, 106, 99, 95, 92, 90, 81, 
    84, 85, 92, 94, 106, 109, 130, 190, 186, 181, 202, 221, 229, 224, 237, 
    243, 255, 264, 146, 110, 114, 134, 119, 136, 144, 132, 132, 135, 141, 
    112, 113, 108, 110, 103, 109, 157, 112, 149, 150, 148, 146, 151, 157, 
    327, 324, 328, 326, 320, 315, 310, 307, 308, 310, 306, 296, 298, 299, 
    294, 300, 297, 297, 294, 294, 300, 304, 315, 318, 328, 332, 333, 334, 
    338, 336, 352, 342, 345, 339, 340, 345, 357, 352, 347, 355, 356, 357, 
    354, 3, 357, 344, 340, 357, 360, 333, 352, 342, 341, 340, 306, 311, 338, 
    320, 321, 348, 79, 331, 71, 119, 119, 117, 143, 149, 154, 158, 157, 164, 
    160, 158, 151, 149, 210, 231, 206, 223, 213, 227, 233, 265, 331, 334, 
    323, 319, 298, 308, 302, 310, 298, 311, 301, 308, 305, 319, 320, 328, 
    327, 326, 328, 335, 340, 335, 343, 356, 360, 1, 346, 4, 37, 69, 120, 93, 
    128, 122, 112, 111, 119, 121, 127, 146, 149, 165, 180, 175, 175, 157, 
    155, 166, 150, 154, 157, 150, 157, 137, 167, 146, 150, 186, 161, 144, 
    153, 191, 175, 253, 6, 6, 20, 54, 1, 102, 87, 91, 90, 90, 85, 85, 74, 85, 
    87, 90, 150, 152, 172, 183, 196, 25, 20, 15, 11, 360, 356, 349, 345, 346, 
    343, 343, 345, 339, 339, 345, 345, 347, 338, 338, 330, 332, 335, 332, 
    325, 326, 325, 327, 327, 325, 327, 78, 263, 261, 267, 283, 287, 299, 276, 
    26, 47, 54, 63, 61, 60, 55, 43, 46, 39, 44, 40, 43, 45, 43, 51, 54, 52, 
    52, 50, 48, 46, 46, 44, 47, 45, 50, 62, 50, 69, 62, 57, 49, 48, 42, 48, 
    46, 45, 50, 52, 52, 48, 38, 32, 36, 18, 16, 15, 13, 7, 3, 2, 7, 9, 12, 
    10, 4, 2, 351, 350, 347, 346, 1, 356, 352, 348, 347, 350, 349, 352, 350, 
    360, 342, 347, 355, 338, 349, 343, 344, 350, 323, 331, 322, 319, 318, 
    320, 322, 318, 329, 326, 315, 324, 320, 326, 22, 59, 69, 61, 71, 94, 313, 
    328, 332, 339, 343, 337, 23, 15, 11, 359, 360, 6, 355, 353, 344, 355, 
    348, 342, 336, 349, 333, 333, 321, 341, 344, 339, 344, 340, 343, 346, 
    339, 346, 340, 336, 333, 337, 338, 348, 341, 347, 330, 325, 326, 328, 
    328, 335, 335, 325, 321, 315, 338, 340, 346, 346, 337, 352, 353, 326, 
    337, 331, 325, 326, 327, 333, 321, 325, 334, 348, 340, 332, 333, 354, 
    340, 328, 326, 327, 332, 329, 336, 344, 344, 349, 348, 339, 337, 333, 
    342, 338, 343, 350, 341, 336, 354, 348, 347, 342, 351, 351, 354, 338, 
    351, 353, 354, 352, 352, 351, 353, 352, 353, 342, 348, 357, 342, 354, 
    355, 355, 1, 359, 4, 325, 317, 336, 20, 89, 89, 127, 127, 128, 169, 175, 
    170, 180, 182, 177, 180, 187, 193, 193, 197, 199, 210, 214, 214, 223, 
    243, 244, 249, 244, 237, 240, 240, 275, 294, 310, 315, 309, 1, 343, 352, 
    348, 4, 350, 5, 10, 18, 13, 12, 358, 357, 358, 350, 353, 346, 358, 7, 8, 
    5, 4, 4, 359, 360, 8, 3, 15, 7, 14, 34, 81, 68, 103, 79, 284, 47, 47, 69, 
    70, 64, 62, 68, 89, 67, 132, 137, 104, 100, 19, 256, 81, 263, 258, 93, 
    99, 100, 129, 78, 127, 132, 131, 129, 129, 124, 133, 120, 121, 99, 98, 
    103, 100, 99, 100, 89, 87, 88, 86, 87, 88, 93, 93, 98, 113, 131, 64, 107, 
    97, 98, 95, 87, 25, 69, 52, 81, 83, 57, 86, 81, 73, 89, 83, 110, 123, 
    124, 157, 65, 81, 127, 109, 119, 115, 113, 134, 158, 163, 154, 150, 152, 
    146, 148, 145, 141, 143, 143, 143, 141, 138, 140, 142, 140, 138, 132, 
    129, 123, 121, 125, 120, 117, 116, 112, 115, 112, 102, 95, 99, 94, 94, 
    91, 94, 93, 95, 98, 98, 97, 97, 94, 91, 84, 72, 41, 54, 61, 62, 65, 70, 
    71, 70, 67, 66, 66, 66, 69, 69, 73, 67, 74, 74, 55, 60, 62, 58, 64, 66, 
    64, 49, 43, 58, 48, 10, 34, 37, 33, 48, 52, 53, 54, 18, 36, 58, 74, 72, 
    69, 60, 62, 63, 65, 27, 347, 16, 69, 323, 332, 85, 86, 84, 77, 81, 85, 
    100, 69, 320, 305, 320, 336, 358, 66, 53, 55, 48, 40, 33, 47, 81, 80, 83, 
    66, 64, 52, 60, 61, 57, 55, 53, 69, 78, 68, 5, 290, 41, 85, 72, 329, 88, 
    87, 57, 63, 67, 62, 57, 58, 58, 67, 61, 73, 75, 74, 91, 93, 91, 97, 85, 
    85, 85, 79, 87, 78, 75, 73, 79, 78, 76, 69, 72, 65, 71, 69, 53, 93, 67, 
    74, 77, 78, 80, 80, 100, 169, 76, 82, 330, 338, 68, 62, 59, 70, 71, 74, 
    67, 65, 61, 57, 72, 67, 76, 77, 81, 86, 72, 60, 55, 60, 54, 111, 67, 63, 
    57, 56, 65, 64, 67, 57, 54, 55, 59, 63, 50, 58, 60, 70, 73, 73, 61, 74, 
    68, 85, _, 53, 51, 44, 46, 41, 48, 47, 47, 22, 41, 40, 37, 56, 44, 44, 
    47, 44, 44, 62, 48, 49, 50, 49, 41, 37, 40, _, 38, _, 20, 11, 30, 34, 33, 
    47, 16, 23, 20, 21, 19, 25, 25, 22, 17, _, 16, 13, 14, 16, 22, 16, 24, 
    32, 39, 36, 38, 37, 36, 29, 33, 29, 35, 32, 36, 20, 22, 20, 17, 11, 11, 
    12, 41, 41, 40, 49, 58, 44, 35, 38, 38, 50, 60, 37, 45, 43, 40, 52, 51, 
    53, 40, 52, 56, 55, 53, 80, 77, 79, 73, 55, 87, 65, 42, 67, 51, 67, 64, 
    72, 116, 68, 66, 64, 79, 125, 113, 133, 144, 143, 134, 137, 139, 137, 
    136, 144, 98, 124, 63, 123, 125, 43, 126, 143, 160, 144, 152, 165, 178, 
    253, 231, 118, 245, 255, 243, 248, 250, 233, 159, 208, 145, 189, 125, 
    131, 194, 150, 218, 202, 148, 155, 153, 162, 153, 153, 144, 155, 150, 
    146, 155, 154, 155, 166, 156, 160, 164, 156, 155, 169, 175, 4, 15, 21, 
    25, 134, 97, 91, 98, 99, 100, 105, 110, 119, 125, 144, 146, 159, 151, 
    153, 152, 156, 159, 160, 169, 159, 168, 150, 159, 155, 152, 153, 150, 
    151, 162, 155, 159, 157, 148, 154, 146, 154, 151, 149, 155, 154, 156, 
    168, 155, 147, 150, 149, 159, 156, 159, 153, 156, 150, 151, 139, 138, 
    136, 136, 139, 139, 131, 133, 134, 137, 128, 116, 115, 118, 119, 108, 
    103, 99, 107, 119, _, 149, 137, 149, 137, 124, _, 131, 144, 146, 141, 
    139, 141, 143, 141, 138, 132, 131, 130, 139, 137, 141, 141, 145, 150, 
    150, 153, 142, 142, 142, 146, 148, 143, 151, 148, 154, 155, 153, 146, 
    150, 151, 157, 153, 153, 157, 157, 160, 161, 165, 168, 167, 172, 173, 
    173, 172, 173, 173, 178, 176, 172, 167, 165, 167, 171, 174, 173, 179, 
    182, 184, 181, 178, 182, 186, 181, 185, 175, 184, 156, 170, 180, 189, 
    185, 182, 182, 184, 161, 175, 167, 182, 167, 152, 172, 176, 181, 188, 
    178, 162, 154, 178, 176, 167, 171, 155, 153, 150, 156, 159, 152, 158, 
    162, 169, 169, 166, 170, 171, 167, 169, 170, 170, 176, 175, 176, 182, 
    184, 188, 183, 185, 183, 188, 188, 184, 185, 188, 183, 186, 192, 186, 
    184, 191, 191, 189, 186, 181, 184, 178, 188, 183, 190, 189, 200, 195, 
    192, 194, 191, 194, 195, 192, 190, 199, 197, 201, 200, 204, 206, 203, 
    202, 204, 196, 206, 204, 206, 203, 214, 202, 206, 203, 192, 160, 160, 
    159, 158, 153, 159, 141, 138, 143, 142, 145, 143, 139, 182, 145, 146, 
    148, 156, 138, 138, 143, 152, 143, 151, 155, 156, 162, 161, 160, 152, 
    132, 143, 170, 140, 138, 132, 125, 131, 136, 140, 128, 116, 106, 114, 
    102, 100, 88, 97, 87, 88, 81, 77, 82, 89, 86, 90, 92, 93, 90, 98, 84, 86, 
    81, 84, 79, 71, 66, 61, 64, 67, 69, 70, 79, 81, 79, 63, 53, 50, 45, 52, 
    57, 53, 44, 56, 56, 61, 71, 78, 79, 80, 79, 80, 83, 88, 91, 89, 87, 91, 
    92, 89, 90, 91, 89, 84, 85, 91, 86, 90, 93, 92, 97, 100, 92, 96, 100, 
    112, 107, 126, 160, 187, 104, 106, 289, 326, 358, 8, 200, 138, 155, 151, 
    170, 6, 2, 6, 8, 3, 4, 4, 6, 359, 358, 7, 9, 360, 360, 359, 2, 360, 2, 3, 
    358, 7, 360, 349, 10, 351, 360, 355, 3, 3, 31, 22, 4, 311, 308, 285, 4, 
    5, 1, 355, 30, 32, 358, 84, 161, 0, 321, 22, 310, 335, 261, 261, 249, 
    256, 253, 223, 225, 230, 237, 252, 253, 245, 231, 237, 244, 226, 237, 
    235, 246, 246, 261, 279, 275, 274, 272, 292, 339, 28, 28, 18, 17, 6, 51, 
    49, 63, 51, 64, 69, 87, 70, 65, 74, 63, 62, 60, 36, 34, 57, 43, 59, 39, 
    59, 41, 28, 19, 28, 36, 19, 38, 5, 94, 87, 124, 141, 127, 94, 357, 348, 
    360, 352, 357, 356, 5, 359, 14, 18, 7, 2, 342, 352, 2, 11, 19, 343, 336, 
    324, 345, 353, 352, 357, 356, 357, 354, 352, 355, 353, 2, 6, 4, 357, 349, 
    353, 355, 357, 3, 355, 360, 359, 359, 354, 351, 357, 352, 349, 353, 355, 
    1, 351, 352, 358, 360, 7, 9, 30, 23, 19, 31, 34, 39, 25, 30, 26, 26, 18, 
    31, 36, 28, 24, 15, 351, 359, 2, 7, 6, 1, 2, 2, 5, 10, 9, 4, 4, 1, 4, 8, 
    10, 337, 333, 328, 337, 323, 324, 325, 322, 326, 6, 2, 1, 360, 3, 360, 1, 
    4, 7, 360, 358, 343, 319, 326, 327, 327, 322, 328, 310, 304, 286, 290, 
    295, 298, 300, 296, 300, 310, 310, 312, 324, 294, 278, 282, 287, 360, 
    148, 208, 189, 191, 159, 159, 157, 167, 176, 163, 172, 181, 196, 202, 
    217, 243, 252, 254, 279, 319, 334, 357, 351, 2, 11, 10, 356, 6, 360, 94, 
    87, 56, 67, 0, 357, 8, 169, 133, 0, 292, 331, 352, 26, 128, 13, 20, 35, 
    29, 40, 39, 12, 43, 34, 47, 355, 33, 344, 355, 13, 18, 11, 6, 83, 59, 80, 
    58, 32, 87, 360, 53, 51, 42, 35, 19, 15, 16, 3, 11, 7, 8, 4, 6, 360, 359, 
    358, 354, 2, 350, 355, 340, 345, 335, 334, 337, 343, 344, 341, 342, 347, 
    336, 334, 337, 359, 352, 342, 347, 337, 332, 336, 330, 332, 330, 330, 
    328, 328, 328, 320, 320, 324, 346, 340, 11, 8, 9, 8, 16, 27, 19, 7, 15, 
    20, 18, 15, 23, 12, 10, 8, 12, 11, 5, 5, 4, 7, 12, 2, 350, 348, 346, 359, 
    355, 352, 350, 357, 348, 346, 352, 359, 351, 360, 359, 2, 7, 8, 9, 7, 16, 
    16, 16, 18, 23, 22, 20, 28, 21, 22, 16, 12, 22, 25, 27, 18, 18, 15, 30, 
    9, 336, 338, 1, 340, _, 338, 326, 348, 345, 332, 335, 334, 341, 339, 338, 
    340, 341, 333, 340, 341, 347, 347, 347, 351, 350, 353, 354 ;

 relative_humidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, -1, -1, -1, -1, -1, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, _, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, _, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -1, -1, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -1, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, _, -1, -1, _, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    _, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, _, _, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, _, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, _, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.87, 0.87, 0.89, 0.9, 0.89, -1, 0.93, 0.93, 0.94, 0.95, 0.95, 0.94, 
    0.95, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.95, 0.95, 0.94, 0.93, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.94, 0.95, 0.96, 0.97, 0.96, 0.94, _, _, _, _, _, _, 0.79, 0.79, 0.81, 
    0.85, 0.89, 0.94, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.96, 0.98, 0.95, 
    0.93, 0.93, 0.93, 0.9, 0.88, 0.87, 0.87, 0.87, 0.87, 0.88, 0.88, 0.87, 
    0.88, 0.89, 0.9, 0.91, 0.9, 0.92, 0.92, 0.92, 0.93, 0.94, 0.94, 0.94, 
    0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.93, 0.93, 0.93, 0.92, 
    0.92, 0.92, 0.92, 0.96, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.97, 0.97, 0.97, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.91, 0.91, 
    0.92, 0.92, 0.92, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 0.94, 0.93, 
    0.92, 0.92, 0.92, 0.95, 0.94, 0.95, 0.97, 0.97, 0.95, 0.93, 0.93, 0.92, 
    0.89, 0.89, 0.96, 0.97, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.95, 0.98, 
    0.98, 0.96, 0.95, 0.96, 0.96, 0.95, 0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 
    0.94, 0.94, 0.96, 0.96, 0.96, 0.97, 0.95, 0.94, 0.94, 0.94, 0.93, 0.94, 
    0.94, 0.93, 0.91, 0.91, 0.87, 0.8, 0.78, 0.81, 0.88, 0.92, 0.93, 0.93, 
    0.94, 0.93, 0.92, 0.89, 0.92, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.93, 
    0.93, 0.92, 0.93, 0.92, 0.93, 0.94, 0.95, 0.96, 0.97, 0.96, 0.97, 0.95, 
    0.96, 0.96, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.95, 
    0.94, 0.93, 0.92, 0.95, 0.93, 0.92, 0.92, 0.92, 0.91, 0.9, 0.9, 0.89, 
    0.87, 0.86, 0.87, 0.89, 0.91, 0.92, 0.93, 0.94, 0.94, 0.95, 0.94, 0.94, 
    0.94, 0.94, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 
    0.93, 0.93, 0.93, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 
    0.94, 0.94, 0.93, 0.93, 0.91, 0.91, 0.9, 0.89, 0.88, 0.87, 0.86, 0.86, 
    0.86, 0.86, 0.86, 0.82, 0.81, 0.81, 0.81, 0.81, 0.82, 0.82, 0.83, 0.84, 
    0.84, 0.82, 0.8, 0.81, 0.81, 0.81, 0.82, 0.83, 0.83, 0.84, 0.84, 0.85, 
    0.86, 0.88, 0.88, 0.88, 0.89, 0.9, 0.91, 0.92, 0.93, 0.93, 0.94, 0.94, 
    0.93, 0.93, 0.94, 0.91, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.91, 0.92, 
    0.92, 0.92, 0.93, 0.94, 0.95, 0.95, 0.96, 0.95, 0.94, 0.94, 0.94, 0.93, 
    0.93, 0.92, 0.9, 0.9, 0.88, 0.87, 0.85, 0.84, 0.84, 0.85, 0.86, 0.85, 
    0.86, 0.9, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.92, 0.93, 0.94, 0.94, 
    0.95, 0.95, 0.93, 0.93, 0.93, 0.94, 0.93, 0.93, 0.93, 0.91, 0.89, 0.89, 
    0.9, 0.92, 0.94, 0.94, 0.91, 0.9, 0.91, 0.92, 0.93, 0.93, 0.94, 0.92, 
    0.93, 0.97, 0.99, 0.98, 0.97, 0.94, 0.94, 0.93, 0.96, 0.96, 0.96, 0.95, 
    0.87, 0.85, 0.87, 0.9, 0.92, 0.94, 0.95, 0.95, 0.95, 0.95, 0.96, 0.97, 
    0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.95, 0.96, 0.96, 0.96, 0.97, 0.97, 0.95, 0.93, 0.97, 0.96, 
    0.97, 0.96, 0.91, 0.92, 0.93, 0.94, 0.93, 0.92, 0.9, 0.9, 0.92, 0.93, 
    0.94, 0.94, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.94, 0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.94, 0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 
    0.94, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 
    0.92, 0.93, 0.93, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.95, 0.96, 0.95, 
    0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.94, 
    0.93, 0.92, 0.95, 0.95, 0.94, 0.94, 0.94, 0.92, 0.91, 0.96, 0.97, 0.97, 
    0.96, 0.96, 0.95, 0.97, 0.97, 0.96, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 
    0.97, 0.96, 0.97, 0.97, 0.96, 0.94, 0.95, 0.95, 0.96, 0.97, 0.97, 0.98, 
    0.97, 0.94, 0.92, 0.92, 0.93, 0.95, 0.96, 0.97, 0.98, 0.97, 0.96, 0.96, 
    0.97, 0.97, 0.96, 0.95, 0.94, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.95, 
    0.95, 0.95, 0.93, 0.93, 0.92, 0.93, 0.93, 0.93, 0.93, 0.91, 0.91, 0.91, 
    0.91, 0.92, 0.9, 0.89, 0.9, 0.9, 0.91, 0.92, 0.92, 0.91, 0.91, 0.91, 
    0.93, 0.94, 0.96, 0.96, 0.95, 0.93, 0.92, 0.91, 0.9, 0.9, 0.88, 0.87, 
    0.86, 0.87, 0.91, 0.92, 0.92, 0.91, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 
    0.92, 0.92, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 0.91, 0.91, 0.89, 
    0.88, 0.88, 0.9, 0.91, 0.88, 0.88, 0.89, 0.9, 0.9, 0.89, 0.89, 0.9, 0.91, 
    0.92, 0.8, 0.81, 0.82, 0.84, 0.87, 0.9, 0.91, 0.9, 0.86, 0.82, 0.82, 
    0.83, 0.75, 0.77, 0.8, 0.85, 0.89, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.92, 0.9, 0.89, 0.91, 0.94, 0.95, 0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 
    0.95, 0.96, 0.97, 0.96, 0.95, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 
    0.96, 0.98, 0.98, 0.98, 0.98, 0.97, 0.98, 0.97, 0.97, 0.97, 0.96, 0.96, 
    0.95, 0.96, 0.91, 0.88, 0.88, 0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 0.87, 
    0.87, 0.87, 0.87, 0.88, 0.91, 0.93, 0.92, 0.92, 0.93, 0.92, 0.91, 0.93, 
    0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 
    0.96, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.98, 0.98, 0.97, 0.96, 0.95, 0.93, 0.92, 0.92, 0.92, 0.92, 
    0.91, 0.92, 0.92, 0.92, 0.95, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.96, 
    0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.95, 0.95, 0.95, 
    0.96, 0.96, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 
    0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.95, 0.93, 0.93, 
    0.93, 0.9, 0.89, 0.89, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.91, 0.92, 0.92, 
    0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 
    0.95, 0.94, 0.94, 0.93, 0.93, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.92, 
    0.91, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.91, 0.91, 
    0.89, 0.89, 0.91, 0.91, 0.92, 0.94, 0.93, 0.92, 0.93, 0.93, 0.93, 0.94, 
    0.94, 0.95, 0.97, 0.98, 0.96, 0.94, 0.94, 0.93, 0.91, 0.91, 0.91, 0.92, 
    0.94, 0.94, 0.91, 0.85, 0.85, 0.85, 0.87, 0.89, 0.9, 0.91, 0.93, 0.95, 
    0.93, 0.92, 0.89, 0.86, 0.84, 0.85, 0.87, 0.89, 0.9, 0.91, 0.9, 0.9, 0.9, 
    0.9, 0.9, 0.9, 0.9, 0.9, 0.91, 0.91, 0.9, 0.9, 0.9, 0.89, 0.87, 0.87, 
    0.88, 0.88, 0.88, 0.88, 0.89, 0.89, 0.88, 0.87, 0.85, 0.84, 0.83, 0.81, 
    0.8, 0.79, 0.79, 0.81, 0.84, 0.88, 0.91, 0.91, 0.92, 0.94, 0.93, 0.93, 
    0.93, 0.94, 0.94, 0.94, 0.95, 0.97, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 
    0.94, 0.93, 0.93, 0.93, 0.93, 0.92, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.95, 0.94, 0.9, 0.87, 0.9, 0.89, 
    0.89, 0.9, 0.88, 0.86, 0.84, 0.84, 0.86, 0.88, 0.9, 0.9, 0.9, 0.9, 0.91, 
    0.92, 0.94, 0.95, 0.94, 0.93, 0.92, 0.93, 0.91, 0.91, 0.9, 0.91, 0.9, 
    0.9, 0.88, 0.88, 0.89, 0.89, 0.88, 0.88, 0.87, 0.87, 0.9, 0.91, 0.91, 
    0.91, 0.91, 0.9, 0.91, 0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 0.92, 
    0.91, 0.9, 0.89, 0.89, 0.9, 0.91, 0.92, 0.93, 0.94, 0.93, 0.94, 0.95, 
    0.95, 0.94, 0.94, 0.94, 0.94, 0.93, 0.93, 0.94, 0.94, 0.95, 0.94, 0.93, 
    0.93, 0.92, 0.92, 0.93, 0.92, 0.93, 0.93, 0.95, 0.95, 0.96, 0.95, 0.94, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.89, 0.87, 0.85, 0.84, 
    0.85, 0.87, 0.89, 0.91, 0.92, 0.93, 0.95, 0.96, 0.95, 0.93, 0.92, 0.92, 
    0.91, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 0.9, 0.89, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 0.87, 0.88, 0.9, 0.93, 0.94, 
    0.91, 0.91, 0.92, 0.93, 0.94, 0.94, 0.96, 0.96, 0.95, 0.94, 0.95, 0.94, 
    0.94, 0.95, 0.94, 0.92, 0.91, 0.91, 0.92, 0.94, 0.94, 0.96, 0.95, 0.94, 
    0.96, 0.97, 0.97, 0.96, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 
    0.94, 0.95, 0.96, 0.96, 0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 
    0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.95, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 0.97, 0.96, 0.95, 0.93, 0.91, 0.9, 
    0.88, 0.87, 0.87, 0.85, 0.82, 0.81, 0.8, 0.8, 0.8, 0.78, 0.79, 0.8, 0.82, 
    0.82, 0.82, 0.82, 0.83, 0.84, 0.85, 0.86, 0.87, 0.85, 0.85, 0.85, 0.84, 
    0.82, 0.82, 0.81, 0.81, 0.82, 0.82, 0.83, 0.84, 0.88, 0.88, 0.88, 0.91, 
    0.89, 0.85, 0.83, 0.8, 0.8, 0.8, 0.79, 0.8, 0.82, 0.81, 0.8, 0.81, 0.8, 
    0.79, 0.79, 0.78, 0.78, 0.79, 0.79, 0.8, 0.88, 0.88, 0.88, 0.88, 0.89, 
    0.9, 0.93, 0.91, 0.93, 0.91, 0.88, 0.83, 0.85, 0.85, 0.83, 0.82, 0.82, 
    0.84, 0.86, 0.87, 0.87, 0.88, 0.89, 0.89, 0.88, 0.87, 0.88, 0.9, 0.91, 
    0.91, 0.92, 0.91, 0.89, 0.9, 0.91, 0.91, 0.92, 0.93, 0.91, 0.88, 0.87, 
    0.87, 0.83, 0.79, 0.78, 0.8, 0.81, 0.82, 0.84, 0.85, 0.86, 0.86, 0.86, 
    0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.87, 0.84, 0.84, 0.85, 0.85, 0.85, 
    0.84, 0.84, 0.85, 0.86, 0.88, 0.88, 0.87, 0.88, 0.89, 0.9, 0.91, 0.92, 
    0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 0.94, 0.94, 0.94, 0.93, 0.92, 0.91, 
    0.91, 0.93, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.95, 0.93, 0.92, 0.92, 0.91, 0.89, 0.91, 0.92, 0.93, 0.94, 0.94, 
    0.92, 0.92, 0.92, 0.93, 0.94, 0.95, 0.95, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.98, 0.99, 0.98, 0.96, 0.87, 0.88, 0.85, 0.8, 0.8, 0.8, 0.81, 
    0.81, 0.82, 0.81, 0.81, 0.82, 0.85, 0.86, 0.79, 0.84, 0.88, 0.87, 0.89, 
    0.85, 0.85, 0.86, 0.88, 0.9, 0.92, 0.87, 0.81, 0.85, 0.87, 0.89, 0.88, 
    0.87, 0.87, 0.88, 0.89, 0.9, 0.9, 0.91, 0.92, 0.91, 0.92, 0.92, 0.9, 0.9, 
    0.9, 0.9, 0.9, 0.92, 0.91, 0.91, 0.77, 0.78, 0.79, 0.79, 0.8, 0.82, 0.84, 
    0.87, 0.89, 0.9, 0.92, 0.94, 0.95, 0.93, 0.92, 0.92, 0.91, 0.92, 0.92, 
    0.92, 0.92, 0.92, 0.91, 0.85, 0.83, 0.82, 0.83, 0.83, 0.83, 0.83, 0.83, 
    0.84, 0.85, 0.87, 0.9, 0.92, 0.85, 0.86, 0.82, 0.81, 0.84, 0.87, 0.86, 
    0.83, 0.8, 0.78, 0.77, 0.77, 0.76, 0.73, 0.71, 0.71, 0.71, 0.74, 0.75, 
    0.78, 0.81, 0.86, 0.9, 0.92, 0.82, 0.87, 0.9, 0.92, 0.94, 0.95, 0.94, 
    0.94, 0.94, 0.94, 0.95, 0.95, 0.93, 0.92, 0.9, 0.86, 0.82, 0.79, 0.77, 
    0.76, 0.74, 0.73, 0.74, 0.77, 0.92, 0.93, 0.95, 0.97, 0.96, 0.93, 0.94, 
    0.94, 0.93, 0.91, 0.9, 0.87, 0.77, 0.74, 0.73, 0.72, 0.73, 0.74, 0.77, 
    0.78, 0.8, 0.84, 0.88, 0.9, 0.8, 0.81, 0.79, 0.77, 0.76, 0.75, 0.76, 
    0.77, 0.77, 0.75, 0.72, 0.71, 0.72, 0.72, 0.73, 0.75, 0.76, 0.76, 0.76, 
    0.75, 0.7, 0.72, 0.74, 0.73, 0.76, 0.76, 0.78, 0.78, 0.78, 0.79, 0.83, 
    0.86, 0.85, 0.86, 0.86, 0.84, 0.83, 0.83, 0.85, 0.87, 0.88, 0.88, 0.91, 
    0.93, 0.95, 0.95, 0.94, 0.95, 0.99, 0.98, 0.99, 0.97, 0.95, 0.95, 0.96, 
    0.96, 0.98, 0.98, 0.98, 0.98, 0.93, 0.92, 0.95, 0.96, 0.97, 0.97, 0.98, 
    0.97, 0.97, 0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 
    0.96, 0.97, 0.97, 0.98, 0.98, 0.99, 0.97, 0.99, 0.98, 0.96, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 0.95, 0.96, 
    0.97, 0.98, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.97, 0.98, 0.97, 0.95, 0.93, 0.92, 0.92, 0.91, 
    0.91, 0.91, 0.91, 0.91, 0.93, 0.99, 0.99, 0.99, 1, 1, 0.97, 0.96, 0.98, 
    0.98, 0.95, 0.95, 0.95, 0.93, 0.92, 0.9, 0.9, 0.91, 0.93, 0.93, 0.92, 
    0.94, 0.96, 0.98, 0.98, 0.98, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 0.97, 0.97, 0.98, 0.98, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.97, 0.96, 0.96, 0.95, 
    0.95, 0.96, 0.97, 0.97, 0.96, 0.94, 0.94, 0.96, 0.98, 0.97, 0.97, 0.98, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.95, 0.95, 0.95, 0.95, 0.97, 0.96, 0.95, 0.93, 0.93, 0.93, 0.94, 0.95, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.95, 0.96, 0.95, 0.94, 0.93, 0.93, 0.94, 0.91, 
    0.9, 0.91, 0.92, 0.93, _, _, _, _, _, _, _, _, _, _, _, _, 0.79, 0.78, 
    0.81, 0.83, 0.87, 0.91, 0.92, 0.92, 0.93, 0.93, 0.95, 0.96, 0.93, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.95, 0.96, 0.95, 0.95, 0.95, 0.95, 0.93, 0.93, 
    0.92, 0.92, 0.91, 0.9, 0.89, 0.89, 0.89, 0.89, 0.89, 0.9, 0.91, 0.92, 
    0.93, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.92, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.92, 0.92, 0.9, 0.9, 0.91, 
    0.91, 0.91, 0.91, 0.95, 0.97, 0.98, 0.99, 0.99, 0.96, 0.95, 0.86, 0.85, 
    0.84, 0.83, 0.83, 0.84, 0.85, 0.88, 0.91, 0.92, 0.92, 0.96, 0.96, 0.98, 
    0.97, 0.95, 0.91, 0.91, 0.91, 0.9, 0.92, 0.93, 0.9, 0.87, 0.94, 0.9, 
    0.89, 0.87, 0.88, 0.89, 0.88, 0.9, 0.91, 0.93, 0.94, 0.95, 0.95, 0.96, 
    0.92, 0.95, 0.94, 0.95, 0.97, 0.95, 0.93, 0.92, 0.93, 0.93, 0.94, 0.93, 
    0.92, 0.92, 0.92, 0.93, 0.94, 0.95, 0.95, 0.97, 0.97, 0.98, 0.96, 0.96, 
    0.95, 0.95, 0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.96, 
    0.94, 0.96, 0.95, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 
    0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.93, 0.94, 0.95, 0.93, 
    0.93, 0.93, 0.92, 0.9, 0.92, 0.94, 0.93, 0.94, 0.95, 0.94, 0.96, 0.95, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 0.96, 0.95, 0.96, 
    0.96, 0.94, 0.95, 0.96, 0.94, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.95, 
    0.94, 0.94, 0.93, 0.94, 0.95, 0.94, 0.96, 0.96, 0.95, 0.94, 0.95, 0.93, 
    0.91, 0.93, 0.94, 0.92, 0.92, 0.92, 0.92, 0.92, 0.89, 0.88, 0.93, 0.94, 
    0.92, 0.91, 0.91, 0.92, 0.9, 0.9, 0.91, 0.91, 0.92, 0.93, 0.92, 0.91, 
    0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 0.92, 0.92, 0.92, 0.92, 0.8, 0.79, 
    0.81, 0.81, 0.81, 0.82, 0.83, 0.8, 0.77, 0.76, 0.75, 0.77, 0.73, 0.75, 
    0.75, 0.75, 0.75, 0.73, 0.72, 0.79, 0.82, 0.85, 0.87, 0.89, 0.89, 0.9, 
    0.9, 0.88, 0.88, 0.89, 0.89, 0.9, 0.9, 0.9, 0.9, 0.88, 0.91, 0.91, 0.9, 
    0.89, 0.89, 0.89, 0.89, 0.9, 0.9, 0.91, 0.91, 0.91, 0.94, 0.93, 0.92, 
    0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.94, 0.95, 0.95, 0.96, 0.94, 
    0.93, 0.92, 0.91, 0.91, 0.92, 0.92, 0.93, 0.92, 0.92, 0.9, 0.89, 0.88, 
    0.88, 0.86, 0.85, 0.86, 0.8, 0.8, 0.78, 0.79, 0.81, 0.77, 0.76, 0.77, 
    0.78, 0.8, 0.82, 0.81, 0.79, 0.77, 0.75, 0.75, 0.75, 0.73, 0.7, 0.7, 
    0.71, 0.72, 0.71, 0.72, 0.73, 0.73, 0.71, 0.69, 0.7, 0.72, 0.74, 0.71, 
    0.65, 0.62, 0.6, 0.58, 0.58, 0.58, 0.59, 0.6, 0.61, 0.97, 0.97, 0.97, 
    0.97, 0.93, 0.84, 0.72, 0.66, 0.67, 0.7, 0.75, 0.79, 0.69, 0.66, 0.65, 
    0.64, 0.66, 0.68, 0.71, 0.75, 0.77, 0.8, 0.83, 0.85, 0.89, 0.92, 0.95, 
    0.93, 0.88, 0.83, 0.81, 0.79, 0.78, 0.76, 0.75, 0.74, 0.65, 0.65, 0.6, 
    0.61, 0.61, 0.59, 0.59, 0.58, 0.57, 0.58, 0.59, 0.61, 0.68, 0.65, 0.64, 
    0.66, 0.68, 0.69, 0.7, 0.7, 0.72, 0.73, 0.78, 0.81, 0.83, 0.83, 0.83, 
    0.84, 0.84, 0.81, 0.8, 0.8, 0.8, 0.79, 0.78, 0.79, 0.83, 0.85, 0.88, 
    0.91, 0.93, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.93, 0.88, 
    0.86, 0.82, 0.79, 0.79, 0.78, 0.79, 0.8, 0.74, 0.7, 0.75, 0.69, 0.67, 
    0.67, 0.67, 0.67, 0.66, 0.67, 0.7, 0.71, 0.72, 0.73, 0.79, 0.79, 0.8, 
    0.8, 0.81, 0.85, 0.87, 0.87, 0.79, 0.84, 0.86, 0.89, 0.89, 0.9, 0.88, 
    0.86, 0.85, 0.85, 0.87, 0.89, 0.9, 0.9, 0.89, 0.87, 0.84, 0.84, 0.84, 
    0.81, 0.82, 0.83, 0.82, 0.82, 0.83, 0.88, 0.89, 0.91, 0.92, 0.93, 0.92, 
    0.91, 0.87, 0.84, 0.83, 0.82, 0.83, 0.85, 0.88, 0.91, 0.88, 0.9, 0.91, 
    0.92, 0.92, 0.91, 0.92, 0.91, 0.92, 0.95, 0.96, 0.96, 0.94, 0.94, 0.96, 
    0.97, 0.98, 0.99, 0.98, 0.99, 0.99, 0.99, 0.98, 0.99, 0.98, 0.98, 0.98, 
    0.97, 0.96, 0.96, 0.99, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.97, 0.97, 0.98, 0.99, 0.98, 
    0.97, 0.98, 0.98, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.95, 0.95, 0.94, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.96, 0.95, 0.96, 0.96, 0.95, 0.93, 
    0.91, 0.89, 0.88, 0.88, 0.88, 0.89, 0.85, 0.82, 0.8, 0.76, 0.75, 0.74, 
    0.73, 0.73, 0.73, 0.72, 0.71, 0.71, 0.7, 0.7, 0.69, 0.96, 0.96, 0.96, 
    0.96, 0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 0.95, 0.94, 0.93, 0.91, 0.9, 
    0.91, 0.9, 0.89, 0.87, 0.87, 0.87, 0.88, 0.88, 0.87, 0.85, 0.85, 0.86, 
    0.86, 0.88, 0.88, 0.9, 0.92, 0.93, 0.84, 0.81, 0.79, 0.85, 0.85, 0.83, 
    0.81, 0.8, 0.77, 0.74, 0.73, 0.72, 0.72, 0.72, 0.72, 0.71, 0.7, 0.7, 0.7, 
    0.69, 0.69, 0.69, 0.7, 0.7, 0.69, 0.68, 0.68, 0.68, 0.67, 0.66, 0.66, 
    0.65, 0.64, 0.63, 0.63, 0.62, 0.61, 0.6, 0.6, 0.59, 0.59, 0.59, 0.59, 
    0.59, 0.58, 0.6, 0.62, 0.62, 0.62, 0.63, 0.62, 0.73, 0.75, 0.76, 0.78, 
    0.8, 0.82, 0.81, 0.78, 0.78, 0.78, 0.8, 0.81, 0.67, 0.66, 0.64, 0.64, 
    0.66, 0.67, 0.7, 0.72, 0.73, 0.72, 0.72, 0.7, 0.68, 0.69, 0.7, 0.7, 0.73, 
    0.79, 0.81, 0.87, 0.87, 0.86, 0.86, 0.86, 0.88, 0.9, 0.92, 0.92, 0.93, 
    0.93, 0.94, 0.97, 0.98, 0.97, 0.96, 0.95, 0.98, 0.97, 0.96, 0.97, 0.96, 
    0.97, 0.97, 0.98, 0.97, 0.97, 0.95, 0.97, 0.97, 0.94, 0.96, 0.96, 0.95, 
    0.96, 0.95, 0.95, 0.93, 0.9, 0.91, 0.93, 0.97, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.96, 0.99, 0.99, 0.99, 1, 0.99, 0.98, 0.99, 0.98, 0.99, 
    0.98, 0.98, 1, 0.91, 0.83, 0.82, 0.81, 0.78, 0.76, 0.75, 0.75, 0.75, 
    0.77, 0.75, 0.73, 0.71, 0.71, 0.7, 0.68, 0.7, 0.69, 0.7, 0.72, 0.76, 
    0.81, 0.85, 0.88, 0.88, 0.88, 0.89, 0.86, 0.79, 0.8, 0.82, 0.82, 0.79, 
    0.77, 0.73, 0.73, 0.76, 0.79, 0.81, 0.83, 0.84, 0.84, 0.83, 0.81, 0.78, 
    0.73, 0.73, 0.86, 0.87, 0.89, 0.87, 0.87, 0.87, 0.87, 0.86, 0.89, 0.89, 
    0.85, 0.84, 0.84, 0.85, 0.84, 0.85, 0.89, 0.86, 0.9, 0.94, 0.96, 0.98, 
    0.98, 1, 0.98, 0.97, 0.97, 0.97, 0.99, 0.96, 0.92, 0.93, 0.96, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.98, 0.99, 0.98, 0.97, 0.95, 
    0.96, 0.97, 0.96, 0.9, 0.86, 0.83, 0.82, 0.88, 0.86, 0.87, 0.89, 0.89, 
    0.92, 0.94, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.9, 0.9, 0.95, 0.98, 
    0.97, 0.93, 0.9, 0.9, 0.9, 0.89, 0.89, 0.88, 0.9, 0.9, 0.89, 0.85, 0.84, 
    0.84, 0.84, 0.86, 0.87, 0.9, 0.92, 0.93, 0.92, 0.93, 0.94, 0.94, 0.94, 
    0.95, 0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.97, 
    0.95, 0.93, 0.95, 0.96, 0.97, 0.96, 0.92, 0.91, 0.91, 0.91, 0.9, 0.89, 
    0.89, 0.88, 0.89, 0.9, 0.9, 0.92, 0.92, 0.93, 0.94, 0.93, 0.92, 0.92, 
    0.94, 0.95, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 
    0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.96, 0.95, 0.94, 0.94, 
    0.94, 0.93, 0.93, 0.94, 0.94, 0.94, 0.92, 0.93, 0.93, 0.93, 0.94, 0.94, 
    0.95, 0.94, 0.94, 0.92, 0.92, 0.91, 0.9, 0.92, 0.95, 0.93, 0.91, 0.89, 
    0.89, 0.92, 0.93, 0.88, 0.83, 0.87, 0.65, 0.65, 0.66, 0.65, 0.65, 0.67, 
    0.68, 0.71, 0.74, 0.77, 0.79, 0.8, 0.94, 0.93, 0.9, 0.87, 0.86, 0.86, 
    0.86, 0.86, 0.88, 0.88, 0.89, 0.89, 0.7, 0.74, 0.77, 0.79, 0.81, 0.83, 
    0.85, 0.86, 0.88, 0.88, 0.87, 0.85, 0.91, 0.91, 0.91, 0.91, 0.9, 0.87, 
    0.85, 0.86, 0.9, 0.94, 0.91, 0.86, 0.8, 0.79, 0.78, 0.78, 0.79, 0.78, 
    0.78, 0.79, 0.8, 0.79, 0.79, 0.8, 0.78, 0.78, 0.79, 0.8, 0.79, 0.78, 
    0.79, 0.79, 0.78, 0.77, 0.77, 0.76, 0.71, 0.71, 0.71, 0.71, 0.71, 0.71, 
    0.7, 0.71, 0.71, 0.71, 0.71, 0.72, 0.66, 0.64, 0.6, 0.59, 0.61, 0.59, 
    0.61, 0.63, 0.65, 0.66, 0.66, 0.66, 0.52, 0.54, 0.57, 0.61, 0.65, 0.66, 
    0.77, 0.83, 0.86, 0.87, 0.88, 0.88, 0.87, 0.89, 0.89, 0.88, 0.9, 0.85, 
    0.82, 0.88, 0.91, 0.89, 0.9, 0.9, 0.93, 0.93, 0.89, 0.91, 0.91, 0.9, 
    0.86, 0.84, 0.85, 0.88, 0.92, 0.92, 0.76, 0.78, 0.81, 0.87, 0.88, 0.91, 
    0.91, 0.91, 0.91, 0.94, 0.96, 0.94, 0.91, 0.92, 0.92, 0.86, 0.88, 0.93, 
    0.92, 0.83, 0.77, 0.76, 0.77, 0.79, 0.72, 0.77, 0.84, 0.86, 0.84, 0.88, 
    0.91, 0.91, 0.91, 0.89, 0.89, 0.92, 0.91, 0.92, 0.87, 0.89, 0.88, 0.86, 
    0.84, 0.82, 0.81, 0.82, 0.85, 0.86, 0.87, 0.84, 0.8, 0.79, 0.8, 0.8, 0.8, 
    0.83, 0.83, 0.85, 0.86, 0.85, 0.83, 0.83, 0.83, 0.82, 0.83, 0.82, 0.81, 
    0.8, 0.78, 0.77, 0.79, 0.81, _, _, _, _, 0.91, 0.9, 0.88, 0.88, 0.89, 
    0.89, 0.92, 0.91, 0.87, 0.85, 0.88, 0.89, 0.89, 0.88, 0.86, 0.83, 0.85, 
    0.87, 0.87, 0.89, 0.96, 0.97, 0.97, 0.96, 0.97, 0.97, 0.94, 0.94, 0.96, 
    0.95, 0.96, 0.92, 0.86, 0.85, 0.87, 0.9, 0.9, 0.85, 0.81, 0.82, 0.85, 
    0.85, 0.82, 0.81, 0.93, 0.96, 0.98, 0.98, 0.99, 1, 0.99, 0.99, 0.98, 
    0.98, 0.96, 0.94, 0.89, 0.92, 0.92, 0.91, 0.91, 0.86, 0.82, 0.85, 0.88, 
    0.89, 0.88, 0.85, 0.8, 0.8, 0.8, 0.81, 0.82, 0.82, 0.82, 0.83, 0.84, 
    0.85, 0.85, 0.85, 0.83, 0.84, 0.85, 0.86, 0.87, 0.88, 0.89, 0.89, 0.9, 
    0.92, 0.94, 0.95, 0.92, 0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.92, 0.92, 0.93, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.97, 0.98, 
    0.98, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.98, 0.96, 0.94, 0.96, 0.96, 0.95, 0.97, 0.97, 0.98, 0.97, 0.95, 
    0.9, 0.84, 0.82, 0.8, 0.8, 0.8, 0.8, 0.79, 0.78, 0.79, 0.79, 0.8, 0.79, 
    0.79, 0.79, 0.78, 0.79, 0.8, 0.81, 0.81, 0.82, 0.83, 0.84, 0.85, 0.85, 
    0.85, 0.86, 0.86, 0.87, 0.87, 0.88, 0.88, 0.87, 0.87, 0.86, 0.85, 0.85, 
    0.83, 0.83, 0.83, 0.83, 0.82, 0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.8, 
    0.8, 0.8, 0.83, 0.83, 0.83, 0.83, 0.83, 0.84, 0.83, 0.84, 0.84, 0.84, 
    0.83, 0.83, 0.85, 0.85, 0.85, 0.86, 0.85, 0.86, 0.86, 0.86, 0.85, 0.86, 
    0.86, 0.86, 0.87, 0.87, 0.87, 0.87, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 
    0.86, 0.86, 0.85, 0.85, 0.85, 0.86, 0.86, 0.86, 0.86, 0.85, 0.86, 0.86, 
    0.85, 0.85, 0.86, 0.86, 0.86, 0.85, 0.84, 0.84, 0.83, 0.82, 0.8, 0.79, 
    0.78, 0.77, 0.74, 0.72, 0.7, 0.68, 0.66, 0.65, 0.64, 0.65, 0.66, 0.7, 
    0.69, 0.69, 0.68, 0.67, 0.68, 0.69, 0.7, 0.71, 0.72, 0.72, 0.72, 0.71, 
    0.68, 0.66, 0.7, 0.66, 0.64, 0.65, 0.67, 0.63, 0.65, 0.69, 0.71, 0.73, 
    0.72, 0.73, 0.74, 0.78, 0.81, 0.84, 0.88, 0.93, 0.95, 0.95, 0.95, 0.94, 
    0.91, 0.89, 0.82, 0.81, 0.81, 0.81, 0.81, 0.8, 0.8, 0.81, 0.81, 0.82, 
    0.83, 0.83, 0.84, 0.84, 0.86, 0.87, 0.87, 0.88, 0.89, 0.9, 0.9, 0.91, 
    0.93, 0.95, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 0.99, 0.97, 0.95, 0.93, 
    0.92, 0.9, 0.89, 0.89, 0.88, 0.88, 0.88, 0.85, 0.85, 0.84, 0.83, 0.81, 
    0.8, 0.81, 0.8, 0.81, 0.81, 0.83, 0.84, 0.85, 0.86, 0.87, 0.9, 0.92, 
    0.93, 0.93, 0.94, 0.94, 0.95, 0.95, 0.94, 0.93, 0.92, 0.92, 0.91, 0.91, 
    0.89, 0.87, 0.86, 0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.83, 0.84, 
    0.86, 0.81, 0.8, 0.8, 0.8, 0.81, 0.83, 0.84, 0.87, 0.91, 0.92, 0.93, 
    0.96, 0.92, 0.9, 0.9, 0.92, 0.92, 0.92, 0.9, 0.9, 0.88, 0.85, 0.85, 0.85, 
    0.81, 0.77, 0.76, 0.75, 0.74, 0.74, 0.76, 0.77, 0.79, 0.8, 0.81, 0.81, 
    0.79, 0.72, 0.75, 0.77, 0.77, 0.76, 0.75, 0.76, 0.76, 0.77, 0.77, 0.76, 
    0.65, 0.64, 0.65, 0.65, 0.67, 0.66, 0.67, 0.7, 0.72, 0.73, 0.72, 0.7, 
    0.93, 0.93, 0.93, 0.97, 0.98, 0.97, 0.93, 0.92, 0.91, 0.91, 0.91, 0.91, 
    0.89, 0.86, 0.84, 0.82, 0.8, 0.79, 0.79, 0.75, 0.72, 0.69, 0.69, 0.69, 
    0.75, 0.79, 0.82, 0.84, 0.86, 0.89, 0.93, 0.91, 0.85, 0.86, 0.9, 0.88, 
    0.84, 0.78, 0.77, 0.78, 0.79, 0.8, 0.79, 0.78, 0.78, 0.77, 0.75, 0.73, 
    0.69, 0.69, 0.68, 0.67, 0.66, 0.69, 0.72, 0.74, 0.75, 0.76, 0.77, 0.78, 
    0.76, 0.79, 0.81, 0.79, 0.78, 0.78, 0.78, 0.75, 0.74, 0.75, 0.76, 0.73, 
    0.72, 0.7, 0.7, 0.72, 0.73, 0.76, 0.76, 0.76, 0.75, 0.75, 0.74, 0.73, 
    0.77, 0.78, 0.78, 0.78, 0.76, 0.75, 0.75, 0.77, 0.78, 0.79, 0.79, 0.78, 
    0.82, 0.8, 0.79, 0.78, 0.75, 0.73, 0.69, 0.7, 0.75, 0.77, 0.73, 0.72, 
    0.67, 0.66, 0.63, 0.67, 0.7, 0.7, 0.7, 0.7, 0.71, 0.71, 0.73, 0.72, _, _, 
    _, _, _, _, _, _, _, _, _, _, 0.76, 0.76, 0.76, 0.76, 0.77, 0.77, 0.77, 
    0.77, 0.77, 0.77, 0.76, 0.76, 0.77, 0.78, 0.78, 0.79, 0.8, 0.82, 0.85, 
    0.88, 0.91, 0.92, 0.94, 0.95, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.96, 
    0.95, 0.94, 0.93, 0.92, 0.9, 0.84, 0.83, 0.82, 0.81, 0.8, 0.79, 0.79, 
    0.79, 0.78, 0.78, 0.78, 0.78, 0.68, 0.66, 0.65, 0.65, 0.63, 0.64, 0.65, 
    0.69, 0.73, 0.76, 0.77, 0.78, 0.74, 0.76, 0.79, 0.8, 0.83, 0.85, 0.85, 
    0.87, 0.89, 0.91, 0.9, 0.89, 0.89, 0.9, 0.91, 0.92, 0.94, 0.93, 0.91, 
    0.88, 0.83, 0.79, 0.8, 0.81, 0.86, 0.88, 0.89, 0.9, 0.89, 0.85, 0.82, 
    0.81, 0.79, 0.78, 0.78, 0.79, 0.81, 0.82, 0.82, 0.82, 0.81, 0.82, 0.83, 
    0.85, 0.87, 0.9, 0.92, 0.91, 0.87, 0.88, 0.89, 0.89, 0.86, 0.82, 0.8, 
    0.79, 0.78, 0.78, 0.78, 0.78, 0.8, 0.81, 0.81, 0.79, 0.78, 0.78, 0.81, 
    0.83, 0.84, 0.85, 0.86, 0.86, 0.89, 0.9, 0.91, 0.93, 0.94, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.93, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.96, 0.95, 0.95, 0.87, 0.91, 0.95, 0.96, 0.96, 0.97, 0.98, 
    0.98, 0.97, 0.95, 0.93, 0.9, 0.84, 0.81, 0.81, 0.82, 0.82, 0.82, 0.82, 
    0.84, 0.85, 0.87, 0.89, 0.91, 0.8, 0.83, 0.85, 0.87, 0.89, 0.9, 0.94, 
    0.95, 0.96, 0.98, 0.98, 0.98, 0.84, 0.83, 0.85, 0.9, 0.92, 0.94, 0.96, 
    0.98, 0.99, 0.99, 0.99, 0.97, 0.94, 0.96, 0.99, 0.99, 0.99, 0.97, 0.95, 
    0.95, 0.98, 0.99, 0.92, 0.86, 0.91, 0.9, 0.91, 0.93, 0.94, 0.96, 0.98, 
    0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.98, 0.96, 0.84, 0.78, 0.83, 
    0.92, 0.96, 0.97, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.94, 0.85, 0.84, 
    0.82, 0.77, 0.73, 0.7, 0.68, 0.76, 0.79, 0.79, 0.82, 0.83, 0.82, 0.83, 
    0.83, 0.82, 0.81, 0.79, 0.77, 0.77, 0.77, 0.79, 0.82, 0.83, 0.81, 0.81, 
    0.8, 0.81, 0.82, 0.81, 0.81, 0.79, 0.79, 0.8, 0.81, 0.81, 0.8, 0.79, 0.8, 
    0.78, 0.78, 0.77, 0.77, 0.81, 0.8, 0.79, 0.78, 0.78, 0.78, 0.8, 0.81, 
    0.82, 0.83, 0.84, 0.84, 0.87, 0.86, 0.86, 0.85, 0.84, 0.84, 0.83, 0.82, 
    0.82, 0.82, 0.83, 0.82, 0.83, 0.81, 0.81, 0.81, 0.82, 0.82, 0.82, 0.83, 
    0.83, 0.85, 0.87, 0.86, 0.84, 0.84, 0.85, 0.85, 0.86, 0.86, 0.86, 0.86, 
    0.87, 0.88, 0.9, 0.91, 0.88, 0.89, 0.88, 0.88, 0.89, 0.92, 0.96, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.96, 0.96, 
    0.96, 0.97, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.99, 1, 1, 
    0.99, 0.98, 0.99, 0.98, 0.97, 0.96, 0.95, 0.93, 0.92, 0.93, 0.94, 0.93, 
    0.93, 0.93, 0.94, _, _, _, _, _, _, _, _, _, _, _, _, 0.93, 0.95, 0.95, 
    0.95, 0.95, 0.93, 0.91, 0.9, 0.92, 0.89, 0.91, 0.95, 0.96, 0.95, 0.96, 
    0.96, 0.94, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 0.88, 0.88, 0.87, 
    0.87, 0.89, 0.91, 0.92, 0.92, 0.93, 0.94, 0.94, 0.93, 0.88, 0.88, 0.89, 
    0.9, 0.9, 0.91, 0.92, 0.91, 0.91, 0.93, 0.93, 0.92, 0.9, 0.91, 0.91, 
    0.91, 0.91, 0.91, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 
    0.95, 0.96, 0.95, 0.96, 0.93, 0.87, 0.9, 0.92, 0.91, 0.88, 0.9, 0.92, 
    0.94, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 0.98, 0.95, 0.95, 0.95, 0.94, 
    0.93, 0.92, 0.92, 0.9, 0.91, 0.92, 0.92, 0.91, 0.9, 0.88, 0.88, 0.89, 
    0.89, 0.89, 0.9, 0.9, 0.94, 0.96, 0.99, 0.99, 0.98, 0.97, 0.95, 0.95, 
    0.92, 0.97, 0.99, 0.99, 0.96, 0.93, 0.91, 0.91, 0.9, 0.89, 0.9, 0.91, 
    0.91, 0.91, 0.93, 0.9, 0.93, 0.92, 0.93, 0.94, 0.94, 0.94, 0.96, 0.91, 
    0.84, 0.87, 0.85, 0.86, 0.83, 0.87, 0.85, 0.83, 0.82, 0.8, 0.79, 0.78, 
    0.77, 0.77, 0.77, 0.76, 0.75, 0.75, 0.74, 0.75, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.75, 0.75, 0.74, 0.74, 0.72, 0.71, 0.71, 0.72, 0.7, 0.71, 0.7, 
    0.7, 0.69, 0.68, 0.68, 0.67, 0.67, 0.65, 0.64, 0.63, 0.64, 0.64, 0.62, 
    0.61, 0.6, 0.6, 0.6, 0.6, 0.61, 0.64, 0.65, 0.64, 0.64, 0.63, 0.64, 0.66, 
    0.69, 0.69, 0.7, 0.72, 0.73, 0.73, 0.74, 0.76, 0.8, 0.78, 0.83, 0.79, 
    0.85, 0.8, 0.81, 0.81, 0.79, 0.8, 0.82, 0.81, 0.78, 0.78, 0.75, 0.73, 
    0.72, 0.74, 0.76, 0.77, 0.74, 0.73, 0.71, 0.7, 0.69, 0.68, 0.66, 0.65, 
    0.64, 0.67, 0.69, 0.7, 0.73, 0.75, 0.8, 0.81, 0.78, 0.78, 0.8, 0.79, 
    0.79, 0.8, 0.81, 0.82, 0.82, 0.82, 0.84, 0.85, 0.82, 0.82, 0.85, 0.86, 
    0.85, 0.83, 0.82, 0.8, 0.79, 0.8, 0.81, 0.82, 0.9, 0.95, 0.82, 0.86, 0.8, 
    0.8, 0.8, 0.77, 0.72, 0.73, 0.71, 0.68, 0.64, 0.6, 0.58, 0.61, 0.66, 0.7, 
    0.71, 0.66, 0.71, 0.76, 0.71, 0.72, 0.75, 0.76, 0.77, 0.78, 0.81, 0.81, 
    0.81, 0.83, 0.83, 0.82, 0.82, 0.82, 0.8, 0.79, 0.77, 0.76, 0.75, 0.73, 
    0.73, 0.72, 0.71, 0.71, 0.7, 0.7, 0.67, 0.67, 0.67, 0.66, 0.66, 0.64, 
    0.62, 0.6, 0.58, 0.58, 0.58, 0.6, 0.78, 0.75, 0.74, 0.76, 0.73, 0.69, 
    0.69, 0.69, 0.7, 0.67, 0.67, 0.66, 0.66, 0.67, 0.68, 0.68, 0.64, 0.66, 
    0.63, 0.64, 0.63, 0.62, 0.59, 0.6, 0.59, 0.56, 0.56, 0.56, 0.56, 0.57, 
    0.6, 0.63, 0.68, 0.72, 0.71, 0.7, 0.69, 0.69, 0.71, 0.77, 0.8, 0.81, 
    0.83, 0.81, 0.81, 0.8, 0.79, 0.77, 0.72, 0.71, 0.67, 0.64, 0.65, 0.66, 
    0.68, 0.7, 0.7, 0.7, 0.73, 0.79, 0.82, 0.83, 0.92, 0.87, 0.86, 0.82, 
    0.74, 0.71, 0.71, 0.71, 0.71, 0.72, 0.7, 0.69, 0.72, 0.73, 0.74, 0.76, 
    0.81, 0.85, 0.84, 0.83, 0.83, 0.83, 0.88, 0.9, 0.84, 0.64, 0.6, 0.7, 
    0.78, 0.83, 0.83, 0.85, 0.86, 0.86, 0.94, 0.95, 0.96, 0.96, 0.97, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.95, 0.9, 0.93, 0.94, 0.95, 0.93, 0.92, 0.91, 0.92, 0.87, 0.89, 
    0.89, 0.9, 0.89, 0.89, 0.88, 0.88, 0.87, 0.87, 0.84, 0.85, 0.85, 0.86, 
    0.86, 0.87, 0.87, 0.87, 0.88, 0.86, 0.72, 0.68, 0.67, 0.63, 0.62, 0.63, 
    0.69, 0.75, 0.8, 0.84, 0.86, 0.85, 0.91, 0.91, 0.9, 0.88, 0.87, 0.86, 
    0.87, 0.9, 0.93, 0.96, 0.97, 0.97, 0.88, 0.89, 0.89, 0.89, 0.89, 0.84, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.83, 0.83, 0.84, 0.84, 0.84, 0.85, 0.82, 0.83, 0.83, 0.84, 0.85, 0.85, 
    0.86, 0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 0.87, 0.86, 0.86, 0.85, 0.86, 
    0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 0.88, 0.88, 0.88, 0.88, 0.89, 0.89, 
    0.9, 0.89, 0.89, 0.89, 0.9, 0.9, 0.91, 0.91, 0.92, 0.92, 0.91, 0.9, 0.88, 
    0.87, 0.86, 0.87, 0.88, 0.88, 0.87, 0.86, 0.84, 0.85, 0.84, 0.81, 0.79, 
    0.78, 0.78, 0.78, 0.78, 0.78, 0.83, 0.84, 0.84, 0.82, 0.81, 0.79, 0.81, 
    0.81, 0.83, 0.81, 0.78, 0.76, 0.74, 0.74, 0.74, 0.74, 0.73, 0.75, 0.77, 
    0.76, 0.75, 0.75, 0.74, 0.73, 0.8, 0.8, 0.81, 0.79, 0.79, 0.8, 0.79, 
    0.79, 0.76, 0.75, 0.75, 0.76, 0.86, 0.84, 0.84, 0.84, 0.84, 0.84, 0.82, 
    0.81, 0.79, 0.76, 0.75, 0.73, 0.82, 0.82, 0.81, 0.81, 0.81, 0.82, 0.8, 
    0.76, 0.76, 0.78, 0.79, 0.8, 0.79, 0.76, 0.78, 0.82, 0.83, 0.86, 0.87, 
    0.87, 0.88, 0.89, 0.9, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 
    0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 0.94, 0.95, 0.96, 0.95, 0.93, 
    0.93, 0.93, 0.94, 0.96, 0.97, 0.95, 0.95, 0.98, 0.99, 0.99, 0.99, 1, 1, 
    0.96, 0.87, 0.85, 0.85, 0.98, 0.99, 0.98, 0.98, 0.98, 0.99, 0.96, 0.88, 
    0.82, 0.8, 0.8, 0.79, 0.77, 0.74, 0.73, 0.72, 0.73, 0.74, 0.75, 0.74, 
    0.76, 0.75, 0.74, 0.73, 0.72, 0.71, 0.7, 0.69, 0.68, 0.67, 0.67, 0.67, 
    0.67, 0.63, 0.66, 0.7, 0.69, 0.73, 0.75, 0.78, 0.81, 0.85, 0.86, 0.88, 
    0.88, 0.91, 0.91, 0.9, 0.89, 0.89, 0.89, 0.89, 0.88, 0.86, 0.84, 0.82, 
    0.75, 0.79, 0.81, 0.83, 0.84, 0.83, 0.83, 0.85, 0.88, 0.92, 0.94, 0.95, 
    0.93, 0.92, 0.9, 0.88, 0.89, 0.89, 0.9, 0.76, 0.75, 0.74, 0.76, 0.79, 
    0.83, 0.82, 0.82, 0.79, 0.77, 0.72, 0.7, 0.74, 0.72, 0.7, 0.69, 0.69, 
    0.68, 0.69, 0.69, 0.69, 0.7, 0.7, 0.72, 0.73, 0.75, 0.76, 0.78, 0.77, 
    0.76, 0.76, 0.75, 0.75, 0.75, 0.75, 0.74, 0.73, 0.74, 0.74, 0.74, 0.73, 
    0.73, 0.73, 0.73, 0.74, 0.74, 0.73, 0.73, 0.72, 0.71, 0.69, 0.69, 0.68, 
    0.67, 0.7, 0.69, 0.67, 0.67, 0.67, 0.68, 0.68, 0.69, 0.69, 0.69, 0.69, 
    0.68, 0.67, 0.68, 0.71, 0.69, 0.71, 0.72, 0.71, 0.7, 0.68, 0.67, 0.66, 
    0.68, 0.7, 0.72, 0.72, 0.8, 0.79, 0.78, 0.77, 0.76, 0.76, 0.77, 0.76, 
    0.76, 0.75, 0.75, 0.75, 0.73, 0.72, 0.72, 0.72, 0.71, 0.71, 0.71, 0.71, 
    0.7, 0.7, 0.69, 0.67, 0.67, 0.66, 0.63, 0.61, 0.59, 0.61, 0.64, 0.64, 
    0.63, 0.64, 0.65, 0.68, 0.77, 0.84, 0.84, 0.83, 0.82, 0.82, 0.8, 0.77, 
    0.76, 0.76, 0.75, 0.78, 0.81, 0.81, 0.83, 0.85, 0.85, 0.85, 0.85, 0.85, 
    0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 
    0.84, 0.84, 0.85, 0.86, 0.85, 0.85, 0.85, 0.84, 0.83, 0.83, 0.83, 0.83, 
    0.84, 0.84, 0.84, 0.83, 0.84, 0.85, 0.84, 0.84, 0.84, 0.85, 0.86, 0.85, 
    0.85, 0.84, 0.83, 0.81, 0.81, 0.8, 0.78, 0.78, 0.77, 0.76, 0.77, 0.78, 
    0.77, 0.77, 0.76, 0.74, 0.76, 0.75, 0.75, 0.75, 0.75, 0.75, 0.76, 0.77, 
    0.77, 0.77, 0.76, 0.76, 0.75, 0.76, 0.76, 0.76, 0.76, 0.75, 0.74, 0.73, 
    0.72, 0.72, 0.73, 0.75, 0.76, 0.79, 0.82, 0.86, 0.86, 0.85, 0.85, 0.84, 
    0.86, 0.87, 0.87, 0.86, 0.85, 0.84, 0.84, 0.84, 0.83, 0.81, 0.81, 0.81, 
    0.81, 0.8, 0.8, 0.8, 0.82, 0.81, 0.8, 0.79, 0.78, 0.78, 0.77, 0.77, 0.77, 
    0.78, 0.78, 0.79, 0.77, 0.75, 0.75, 0.75, 0.74, 0.74, 0.74, 0.74, 0.73, 
    0.74, 0.74, 0.73, 0.72, 0.72, 0.73, 0.73, 0.74, 0.74, 0.74, 0.74, 0.75, 
    0.76, 0.76, 0.77, 0.79, 0.8, 0.81, 0.8, 0.81, 0.82, 0.82, 0.83, 0.83, 
    0.83, 0.8, 0.82, 0.84, 0.84, 0.85, 0.85, 0.85, 0.86, 0.84, 0.82, 0.79, 
    0.78, 0.79, 0.79, 0.85, 0.85, 0.86, 0.87, 0.83, 0.83, 0.83, 0.83, 0.81, 
    0.8, 0.81, 0.81, 0.85, 0.85, 0.85, 0.85, 0.86, 0.85, 0.85, 0.81, 0.74, 
    0.72, 0.7, 0.74, 0.75, 0.76, 0.78, 0.8, 0.81, 0.82, 0.82, 0.83, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.84, 0.85, 0.86, 0.86, 0.87, 0.88, 0.87, 0.86, 
    0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 0.85, 0.86, 0.87, 0.86, 0.84, 
    0.85, 0.86, 0.86, 0.82, 0.82, 0.83, 0.84, 0.84, 0.85, 0.86, 0.85, 0.84, 
    0.83, 0.84, 0.85, 0.87, 0.86, 0.87, 0.87, 0.86, 0.85, 0.86, 0.86, 0.86, 
    0.87, 0.88, 0.88, 0.85, 0.84, 0.83, 0.82, 0.83, 0.84, 0.83, 0.84, 0.82, 
    0.83, 0.84, 0.85, 0.8, 0.8, 0.81, 0.82, 0.82, 0.83, 0.82, 0.82, 0.82, 
    0.82, 0.83, 0.83, 0.74, 0.74, 0.75, 0.76, 0.76, 0.78, 0.79, 0.79, 0.79, 
    0.8, 0.79, 0.79, 0.72, 0.74, 0.75, 0.75, 0.75, 0.76, 0.76, 0.75, 0.73, 
    0.74, 0.76, 0.75, 0.7, 0.7, 0.71, 0.72, 0.71, 0.71, 0.71, 0.71, 0.72, 
    0.72, 0.75, 0.74, 0.69, 0.68, 0.68, 0.67, 0.67, 0.66, 0.66, 0.66, 0.67, 
    0.69, 0.71, 0.73, 0.7, 0.72, 0.73, 0.74, 0.76, 0.78, 0.8, 0.83, 0.84, 
    0.85, 0.86, 0.86, 0.86, 0.86, 0.87, 0.86, 0.86, 0.86, 0.86, 0.86, 0.87, 
    0.9, 0.93, 0.94, 0.88, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.9, 0.9, 0.9, 
    0.9, 0.9, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.87, 0.86, 
    0.86, 0.86, 0.85, 0.84, 0.85, 0.85, 0.85, 0.86, 0.85, 0.85, 0.84, 0.85, 
    0.86, 0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 0.84, 
    0.83, 0.83, 0.78, 0.78, 0.77, 0.77, 0.77, 0.77, 0.76, 0.76, 0.74, 0.72, 
    0.72, 0.71, 0.82, 0.82, 0.82, 0.82, 0.82, 0.81, 0.81, 0.81, 0.8, 0.8, 
    0.81, 0.82, 0.88, 0.89, 0.9, 0.92, 0.93, 0.94, 0.95, 0.95, 0.96, 0.97, 
    0.99, 0.99, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.98, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 
    0.95, 0.94, 0.92, 0.92, 0.91, 0.92, 0.92, 0.93, 0.93, 0.93, 0.92, 0.92, 
    0.91, 0.91, 0.91, 0.92, 0.91, 0.92, 0.9, 0.9, 0.9, 0.89, 0.89, 0.88, 
    0.88, 0.88, 0.9, 0.89, 0.89, 0.93, 0.91, 0.9, 0.9, 0.91, 0.9, 0.9, 0.9, 
    0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.93, 0.93, 
    0.94, 0.92, 0.91, 0.92, 0.91, 0.91, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 
    0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 
    0.88, 0.88, 0.88, 0.89, 0.89, 0.9, 0.9, 0.89, 0.9, 0.9, 0.9, 0.9, 0.88, 
    0.88, 0.89, 0.89, 0.9, 0.9, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.91, 
    0.89, 0.89, 0.9, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.92, 0.92, 0.91, 0.91, 
    0.91, 0.92, 0.93, 0.94, 0.94, 0.95, 0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.97, 0.93, 0.94, 0.94, 0.94, 0.96, 0.96, 
    0.95, 0.94, 0.93, 0.92, 0.92, 0.94, 0.94, 0.92, 0.92, 0.92, 0.91, 0.91, 
    0.9, 0.89, 0.9, 0.83, 0.78, 0.77, 0.81, 0.82, 0.78, 0.75, 0.78, 0.78, 
    0.78, 0.79, 0.8, 0.8, 0.8, 0.79, 0.77, 0.78, 0.81, 0.82, 0.86, 0.87, 
    0.89, 0.89, 0.87, 0.86, 0.87, 0.88, 0.89, 0.89, 0.88, 0.87, 0.89, 0.89, 
    0.89, 0.88, 0.87, 0.86, 0.86, 0.87, 0.89, 0.92, 0.92, 0.92, 0.93, 0.94, 
    0.92, 0.93, 0.95, 0.95, 0.92, 0.93, 0.93, 0.94, 0.94, 0.93, 0.92, 0.91, 
    0.91, 0.92, 0.92, 0.93, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.91, 
    0.91, 0.93, 0.94, 0.94, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.93, 0.94, 
    0.93, 0.92, 0.92, 0.92, 0.92, 0.9, 0.9, 0.91, 0.91, 0.91, 0.92, 0.92, 
    0.93, 0.93, 0.93, 0.94, 0.94, 0.95, 0.94, 0.93, 0.95, 0.94, 0.83, 0.79, 
    0.77, 0.77, 0.77, 0.8, 0.74, 0.73, 0.73, 0.73, 0.76, 0.76, 0.76, 0.77, 
    0.78, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.8, 0.75, 0.75, 
    0.76, 0.76, 0.77, 0.79, 0.8, 0.83, 0.85, 0.85, 0.86, 0.86, 0.8, 0.82, 
    0.84, 0.86, 0.89, 0.87, 0.86, 0.87, 0.89, 0.89, 0.87, 0.87, 0.85, 0.86, 
    0.85, 0.85, 0.86, 0.87, 0.87, 0.87, 0.88, 0.9, 0.88, 0.8, 0.9, 0.9, 0.87, 
    0.83, 0.8, 0.81, 0.82, 0.82, 0.83, 0.82, 0.83, 0.83, 0.83, 0.84, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.87, 0.88, 0.88, 0.85, 0.83, 0.81, 
    0.8, 0.81, 0.82, 0.83, 0.83, 0.86, 0.89, 0.91, 0.9, 0.85, 0.84, 0.77, 
    0.75, 0.79, 0.86, 0.84, 0.84, 0.86, 0.88, 0.88, 0.88, 0.88, 0.89, 0.87, 
    0.86, 0.83, 0.81, 0.83, 0.82, 0.82, 0.84, 0.87, 0.88, 0.89, 0.87, 0.89, 
    0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.81, 0.78, 0.78, 0.79, 
    0.81, 0.82, 0.81, 0.8, 0.81, 0.82, 0.83, 0.83, 0.86, 0.85, 0.86, 0.85, 
    0.86, 0.87, 0.87, 0.86, 0.86, 0.87, 0.87, 0.86, 0.86, 0.84, 0.84, 0.85, 
    0.84, 0.82, 0.83, 0.81, 0.78, 0.78, 0.77, 0.76, 0.75, 0.74, 0.72, 0.71, 
    0.7, 0.7, 0.71, 0.71, 0.71, 0.7, 0.72, 0.73, 0.7, 0.72, 0.74, 0.75, 0.76, 
    0.78, 0.83, 0.75, 0.73, 0.72, 0.69, 0.69, 0.66, 0.66, 0.67, 0.69, 0.71, 
    0.73, 0.78, 0.81, 0.83, 0.82, 0.83, 0.83, 0.73, 0.74, 0.74, 0.76, 0.78, 
    0.77, 0.77, 0.77, 0.78, 0.79, 0.81, 0.84, 0.69, 0.7, 0.73, 0.77, 0.81, 
    0.8, 0.81, 0.83, 0.85, 0.88, 0.88, 0.88, 0.72, 0.7, 0.69, 0.68, 0.67, 
    0.69, 0.66, 0.67, 0.67, 0.66, 0.66, 0.65, 0.61, 0.63, 0.64, 0.65, 0.66, 
    0.66, 0.66, 0.67, 0.67, 0.67, 0.68, 0.67, 0.63, 0.63, 0.62, 0.62, 0.63, 
    0.69, 0.67, 0.72, 0.68, 0.66, 0.66, 0.69, 0.67, 0.65, 0.65, 0.66, 0.66, 
    0.66, 0.65, 0.66, 0.67, 0.67, 0.67, 0.67, 0.66, 0.66, 0.66, 0.66, 0.66, 
    0.65, 0.64, 0.63, 0.63, 0.75, 0.68, 0.67, 0.66, 0.66, 0.65, 0.65, 0.65, 
    0.65, 0.66, 0.66, 0.67, 0.68, 0.68, 0.68, 0.69, 0.69, 0.69, 0.68, 0.68, 
    0.68, 0.69, 0.69, 0.68, 0.68, 0.69, 0.69, 0.69, 0.7, 0.7, 0.7, 0.7, 0.71, 
    0.71, 0.73, 0.73, 0.74, 0.74, 0.74, 0.69, 0.7, 0.7, 0.7, 0.71, 0.71, 0.7, 
    0.69, 0.69, 0.69, 0.7, 0.7, 0.66, 0.66, 0.67, 0.66, 0.66, 0.67, 0.67, 
    0.67, 0.68, 0.69, 0.7, 0.7, 0.61, 0.61, 0.62, 0.63, 0.64, 0.65, 0.65, 
    0.64, 0.64, 0.64, 0.63, 0.64, 0.65, 0.65, 0.65, 0.66, 0.66, 0.68, 0.68, 
    0.7, 0.71, 0.71, 0.72, 0.73, 0.72, 0.72, 0.72, 0.73, 0.73, 0.73, 0.73, 
    0.72, 0.72, 0.74, 0.75, 0.78, 0.84, 0.85, 0.85, 0.83, 0.84, 0.86, 0.85, 
    0.84, 0.83, 0.82, 0.82, 0.82, 0.83, 0.84, 0.84, 0.83, 0.83, 0.83, 0.84, 
    0.84, 0.84, 0.84, 0.84, 0.86, 0.85, 0.86, 0.87, 0.87, 0.89, 0.88, 0.87, 
    0.89, 0.87, 0.88, 0.89, 0.87, 0.88, 0.89, 0.88, 0.89, 0.89, 0.89, 0.89, 
    0.89, 0.89, 0.89, 0.89, 0.89, 0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 0.85, 
    0.85, 0.86, 0.87, 0.87, 0.88, 0.85, 0.86, 0.86, 0.87, 0.88, 0.89, 0.89, 
    0.89, 0.89, 0.89, 0.89, 0.89, 0.86, 0.87, 0.87, 0.86, 0.86, 0.87, 0.86, 
    0.87, 0.87, 0.86, 0.83, 0.82, 0.8, 0.81, 0.81, 0.8, 0.79, 0.79, 0.77, 
    0.77, 0.78, 0.75, 0.76, 0.77, 0.72, 0.69, 0.7, 0.71, 0.71, 0.71, 0.7, 
    0.71, 0.7, 0.7, 0.7, 0.7, 0.66, 0.66, 0.65, 0.66, 0.66, 0.67, 0.71, 0.73, 
    0.74, 0.76, 0.77, 0.74, 0.64, 0.64, 0.65, 0.66, 0.68, 0.71, 0.73, 0.76, 
    0.79, 0.82, 0.83, 0.84, 0.82, 0.83, 0.83, 0.82, 0.82, 0.81, 0.81, 0.81, 
    0.82, 0.82, 0.82, 0.82, 0.79, 0.79, 0.79, 0.79, 0.79, 0.8, 0.8, 0.81, 
    0.82, 0.82, 0.83, 0.83, 0.77, 0.77, 0.77, 0.77, 0.77, 0.77, 0.77, 0.76, 
    0.76, 0.76, 0.75, 0.75, 0.73, 0.73, 0.73, 0.72, 0.72, 0.72, 0.72, 0.71, 
    0.71, 0.7, 0.7, 0.71, 0.71, 0.71, 0.71, 0.71, 0.7, 0.7, 0.71, 0.71, 0.72, 
    0.73, 0.74, 0.74, 0.79, 0.79, 0.79, 0.8, 0.79, 0.8, 0.8, 0.81, 0.81, 
    0.81, 0.81, 0.81, 0.78, 0.78, 0.79, 0.79, 0.79, 0.8, 0.8, 0.8, 0.8, 0.81, 
    0.8, 0.8, 0.78, 0.79, 0.79, 0.79, 0.78, 0.77, 0.76, 0.75, 0.74, 0.73, 
    0.7, 0.69, 0.67, 0.66, 0.67, 0.69, 0.69, 0.7, 0.72, 0.74, 0.77, 0.79, 
    0.8, 0.81, 0.74, 0.75, 0.76, 0.76, 0.76, 0.76, 0.77, 0.77, 0.76, 0.77, 
    0.77, 0.76, 0.72, 0.72, 0.72, 0.71, 0.72, 0.71, 0.71, 0.71, 0.71, 0.69, 
    0.67, 0.65, 0.59, 0.59, 0.63, 0.58, 0.59, 0.6, 0.62, 0.62, 0.65, 0.69, 
    0.7, 0.73, 0.7, 0.7, 0.72, 0.73, 0.72, 0.73, 0.73, 0.73, 0.75, 0.75, 
    0.76, 0.76, 0.77, 0.78, 0.79, 0.79, 0.79, 0.79, 0.78, 0.75, 0.74, 0.71, 
    0.7, 0.7, 0.72, 0.71, 0.71, 0.7, 0.7, 0.71, 0.71, 0.72, 0.73, 0.71, 0.73, 
    0.75, 0.72, 0.71, 0.73, 0.75, 0.77, 0.79, 0.81, 0.83, 0.84, 0.85, 0.85, 
    0.84, 0.81, 0.81, 0.82, 0.81, 0.82, 0.83, 0.84, 0.85, 0.85, 0.85, 0.87, 
    0.86, 0.93, 0.92, 0.92, 0.91, 0.91, 0.92, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 
    0.89, 0.89, 0.89, 0.89, 0.9, 0.9, 0.91, 0.91, 0.91, 0.9, 0.9, 0.89, 0.86, 
    0.85, 0.84, 0.82, 0.81, 0.8, 0.8, 0.8, 0.81, 0.81, 0.81, 0.82, 0.77, 
    0.78, 0.78, 0.77, 0.77, 0.77, 0.78, 0.78, 0.79, 0.8, 0.8, 0.81, 0.77, 
    0.77, 0.77, 0.77, 0.78, 0.78, 0.78, 0.79, 0.8, 0.81, 0.81, 0.81, 0.81, 
    0.81, 0.79, 0.78, 0.78, 0.77, 0.78, 0.78, 0.78, 0.76, 0.75, 0.74, 0.75, 
    0.74, 0.72, 0.71, 0.71, 0.71, 0.71, 0.7, 0.68, 0.66, 0.66, 0.66, 0.64, 
    0.63, 0.62, 0.62, 0.62, 0.62, 0.62, 0.62, 0.62, 0.62, 0.62, 0.62, 0.59, 
    0.6, 0.6, 0.61, 0.63, 0.65, 0.68, 0.74, 0.75, 0.76, 0.79, 0.8, 0.84, 
    0.83, 0.82, 0.78, 0.79, 0.77, 0.74, 0.76, 0.79, 0.79, 0.8, 0.82, 0.81, 
    0.81, 0.83, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.83, 0.82, 0.8, 
    0.8, 0.81, 0.81, 0.8, 0.8, 0.8, 0.8, 0.79, 0.79, 0.79, 0.79, 0.76, 0.76, 
    0.75, 0.75, 0.75, 0.75, 0.75, 0.75, 0.75, 0.75, 0.76, 0.76, 0.75, 0.75, 
    0.75, 0.75, 0.75, 0.75, 0.74, 0.74, 0.74, 0.74, 0.74, 0.74, 0.74, 0.74, 
    0.74, 0.75, 0.75, 0.75, 0.76, 0.77, 0.78, 0.78, 0.78, 0.78, 0.81, 0.82, 
    0.84, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.85, 0.84, 0.85, 0.85, 0.85, 
    0.85, 0.85, 0.84, 0.84, 0.84, 0.83, 0.82, 0.81, 0.81, 0.8, 0.8, 0.81, 
    0.82, 0.82, 0.82, 0.82, 0.81, 0.81, 0.81, 0.82, 0.84, 0.84, 0.81, 0.79, 
    0.79, 0.79, 0.8, 0.8, 0.8, 0.8, 0.79, 0.79, 0.78, 0.81, 0.82, 0.84, 0.85, 
    0.87, 0.89, 0.91, 0.91, 0.92, 0.89, 0.88, 0.89, 0.89, 0.88, 0.87, 0.86, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.87, 0.87, 0.85, 0.84, 0.84, 
    0.84, 0.84, 0.84, 0.85, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 
    0.84, 0.83, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.8, 0.8, 0.79, 
    0.78, 0.77, 0.77, 0.76, 0.75, 0.75, 0.75, 0.75, 0.77, 0.77, 0.78, 0.8, 
    0.81, 0.82, 0.82, 0.83, 0.84, 0.83, 0.83, 0.84, 0.84, 0.83, 0.84, 0.83, 
    0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.85, 0.85, 
    0.84, 0.84, 0.85, 0.86, 0.86, 0.85, 0.84, 0.84, 0.83, 0.84, 0.84, 0.84, 
    0.84, 0.84, 0.83, 0.82, 0.82, 0.82, 0.82, 0.83, 0.84, 0.84, 0.83, 0.83, 
    0.83, 0.83, 0.83, 0.82, 0.82, 0.85, 0.86, 0.86, 0.89, 0.89, 0.89, 0.89, 
    0.89, 0.89, 0.88, 0.88, 0.88, 0.87, 0.88, 0.89, 0.89, 0.9, 0.89, 0.87, 
    0.86, 0.86, 0.87, 0.88, 0.88, 0.89, 0.89, 0.89, 0.91, 0.89, 0.89, 0.87, 
    0.83, 0.82, 0.82, 0.83, 0.83, 0.83, 0.79, 0.75, 0.72, 0.78, 0.79, 0.81, 
    0.84, 0.87, 0.88, 0.89, 0.88, 0.88, 0.87, 0.86, 0.86, 0.84, 0.84, 0.81, 
    0.81, 0.81, 0.8, 0.8, 0.81, 0.8, 0.8, 0.8, 0.8, 0.82, 0.82, 0.81, 0.82, 
    0.82, 0.82, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.83, 0.83, 
    0.83, 0.83, 0.84, 0.84, 0.84, 0.85, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 
    0.86, 0.85, 0.85, 0.85, 0.86, 0.86, 0.86, 0.85, 0.87, 0.86, 0.83, 0.82, 
    0.82, 0.83, 0.85, 0.85, 0.83, 0.83, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 
    0.83, 0.83, 0.82, 0.82, 0.82, 0.82, 0.82, 0.83, 0.8, 0.8, 0.81, 0.81, 
    0.81, 0.82, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.82, 0.82, 0.83, 0.84, 
    0.84, 0.84, 0.84, 0.84, 0.85, 0.85, 0.85, 0.85, 0.83, 0.82, 0.82, 0.81, 
    0.81, 0.82, 0.83, 0.83, 0.84, 0.85, 0.85, 0.85, 0.83, 0.82, 0.83, 0.84, 
    0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.85, 0.86, 0.84, 0.84, 0.86, 0.87, 
    0.84, 0.82, 0.82, 0.82, 0.82, 0.82, 0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 
    0.83, 0.86, 0.87, 0.88, 0.88, 0.88, 0.89, 0.88, 0.87, 0.87, 0.87, 0.88, 
    0.88, 0.89, 0.88, 0.88, 0.88, 0.86, 0.86, 0.85, 0.89, 0.88, 0.88, 0.86, 
    0.84, 0.82, 0.8, 0.8, 0.8, 0.79, 0.79, 0.8, 0.85, 0.86, 0.87, 0.87, 0.87, 
    0.87, 0.88, 0.88, 0.87, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.84, 0.83, 
    0.82, 0.83, 0.82, 0.82, 0.82, 0.82, 0.83, 0.85, 0.86, 0.87, 0.87, 0.86, 
    0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 0.85, 0.84, 0.83, 0.83, 0.83, 0.83, 
    0.83, 0.83, 0.82, 0.82, 0.83, 0.83, 0.84, 0.83, 0.84, 0.86, 0.87, 0.87, 
    0.85, 0.85, 0.84, 0.82, 0.78, 0.76, 0.76, 0.78, 0.8, 0.81, 0.82, 0.82, 
    0.8, 0.81, 0.81, 0.81, 0.82, 0.83, 0.84, 0.86, 0.86, 0.87, 0.87, 0.88, 
    0.86, 0.84, 0.83, 0.83, 0.83, 0.83, 0.83, 0.82, 0.83, 0.84, 0.85, 0.86, 
    0.87, 0.87, 0.88, 0.88, 0.88, 0.88, 0.87, 0.87, 0.86, 0.86, 0.85, 0.84, 
    0.83, 0.83, 0.82, 0.83, 0.83, 0.84, 0.84, 0.73, 0.75, 0.76, 0.77, 0.79, 
    0.84, 0.86, 0.85, 0.84, 0.84, 0.83, 0.83, 0.84, 0.83, 0.83, 0.83, 0.84, 
    0.85, 0.79, 0.79, 0.8, 0.8, 0.81, 0.81, 0.79, 0.81, 0.82, 0.84, 0.84, 
    0.8, 0.8, 0.8, 0.81, 0.82, 0.82, 0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 
    0.82, 0.82, 0.82, 0.81, 0.8, 0.77, 0.76, 0.75, 0.75, 0.76, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.75, 0.79, 0.8, 0.8, 0.8, 0.79, 
    0.77, 0.75, 0.75, 0.75, 0.74, 0.74, 0.75, 0.75, 0.77, 0.78, 0.78, 0.78, 
    0.79, 0.79, 0.8, 0.82, 0.82, 0.83, 0.83, 0.83, 0.84, 0.85, 0.85, 0.86, 
    0.86, 0.84, 0.83, 0.83, 0.84, 0.85, 0.85, 0.79, 0.81, 0.83, 0.84, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.81, 0.83, 0.84, 0.85, 0.85, 
    0.81, 0.77, 0.77, 0.77, 0.77, 0.77, 0.77, 0.78, 0.79, 0.8, 0.81, 0.81, 
    0.81, 0.82, 0.82, 0.82, 0.82, 0.83, 0.83, 0.79, 0.78, 0.77, 0.78, 0.77, 
    0.78, 0.76, 0.76, 0.75, 0.76, 0.76, 0.74, 0.73, 0.76, 0.78, 0.8, 0.79, 
    0.8, 0.8, 0.81, 0.82, 0.83, 0.84, 0.83, 0.8, 0.82, 0.82, 0.83, 0.82, 
    0.79, 0.77, 0.76, 0.75, 0.74, 0.74, 0.75, 0.81, 0.83, 0.84, 0.85, 0.85, 
    0.86, 0.87, 0.87, 0.86, 0.86, 0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.86, 
    0.87, 0.87, 0.87, 0.86, 0.85, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 
    0.88, 0.88, 0.89, 0.89, 0.89, 0.89, 0.9, 0.91, 0.92, 0.92, 0.92, 0.92, 
    0.92, 0.92, 0.92, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 0.9, 0.91, 0.92, 
    0.92, 0.93, 0.94, 0.94, 0.95, 0.96, 0.97, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.93, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.95, 0.96, 0.95, 0.95, 0.95, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.94, 0.93, 
    0.94, 0.94, 0.95, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.94, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.93, 
    0.93, 0.94, 0.94, 0.93, 0.92, 0.92, 0.91, 0.91, 0.89, 0.87, 0.87, 0.85, 
    0.84, 0.86, 0.88, 0.85, 0.87, 0.89, 0.89, 0.89, 0.88, 0.84, 0.82, 0.82, 
    0.83, 0.82, 0.82, 0.82, 0.84, 0.86, 0.86, 0.87, 0.87, 0.88, 0.88, 0.88, 
    0.89, 0.9, 0.92, 0.91, 0.91, 0.91, 0.9, 0.9, 0.9, 0.89, 0.89, 0.91, 0.91, 
    0.92, 0.91, 0.91, 0.91, 0.9, 0.84, 0.83, 0.87, 0.9, 0.91, 0.91, 0.91, 
    0.93, 0.94, 0.95, 0.94, 0.95, 0.93, 0.91, 0.89, 0.85, 0.84, 0.84, 0.87, 
    0.91, 0.89, 0.89, 0.93, 0.92, 0.94, 0.84, 0.85, 0.88, 0.91, 0.93, 0.94, 
    0.95, 0.94, 0.92, 0.9, 0.9, 0.9, 0.94, 0.95, 0.96, 0.93, 0.9, 0.87, 0.87, 
    0.86, 0.84, 0.83, 0.84, 0.84, 0.83, 0.85, 0.86, 0.86, 0.87, 0.88, 0.88, 
    0.88, 0.87, 0.88, 0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 0.86, 0.86, 0.86, 
    0.87, 0.87, 0.87, 0.87, 0.87, 0.86, 0.87, 0.88, 0.87, 0.87, 0.87, 0.87, 
    0.86, 0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 0.84, 0.84, 0.85, 0.85, 0.85, 
    0.85, 0.85, 0.86, 0.87, 0.87, 0.88, 0.89, 0.9, 0.91, 0.92, 0.93, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.93, 0.91, 0.9, 0.9, 0.89, 0.89, 0.88, 0.87, 
    0.86, 0.87, 0.89, 0.91, 0.92, 0.8, 0.82, 0.83, 0.81, 0.8, 0.78, 0.77, 
    0.77, 0.76, 0.78, 0.77, 0.78, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.79, 0.78, 
    0.77, 0.77, 0.77, 0.77, 0.77, 0.76, 0.75, 0.76, 0.75, 0.76, 0.75, 0.74, 
    0.76, 0.76, 0.76, 0.76, 0.75, 0.75, 0.74, 0.74, 0.74, 0.73, 0.75, 0.76, 
    0.77, 0.77, 0.78, 0.78, 0.81, 0.84, 0.86, 0.87, 0.89, 0.89, 0.89, 0.88, 
    0.88, 0.89, 0.9, 0.89, 0.85, 0.85, 0.84, 0.82, 0.79, 0.8, 0.82, 0.84, 
    0.86, 0.87, 0.87, 0.88, 0.86, 0.88, 0.89, 0.9, 0.9, 0.9, 0.9, 0.89, 0.88, 
    0.86, 0.84, 0.8, 0.83, 0.81, 0.8, 0.77, 0.75, 0.75, 0.75, 0.75, 0.75, 
    0.74, 0.74, 0.75, 0.83, 0.82, 0.81, 0.79, 0.77, 0.77, 0.79, 0.8, 0.79, 
    0.8, 0.79, 0.78, 0.9, 0.89, 0.89, 0.88, 0.87, 0.87, 0.87, 0.87, 0.88, 
    0.88, 0.89, 0.91, 0.89, 0.9, 0.9, 0.91, 0.91, 0.92, 0.93, 0.91, 0.89, 
    0.9, 0.9, 0.92, 0.88, 0.86, 0.85, 0.86, 0.88, 0.9, 0.91, 0.91, 0.91, 
    0.91, 0.92, 0.92, 0.9, 0.9, 0.92, 0.94, 0.94, 0.95, 0.95, 0.95, 0.94, 
    0.93, 0.92, 0.92, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.93, 0.92, 0.92, 0.9, 0.89, 0.9, 0.91, 0.9, 0.9, 0.9, 0.89, 0.87, 0.87, 
    0.84, 0.83, 0.78, 0.74, 0.72, 0.74, 0.73, 0.76, 0.77, 0.75, 0.78, 0.88, 
    0.91, 0.9, 0.88, 0.87, 0.86, 0.86, 0.85, 0.85, 0.86, 0.89, 0.9, 0.88, 
    0.83, 0.82, 0.81, 0.79, 0.78, 0.77, 0.77, 0.78, 0.79, 0.79, 0.77, 0.78, 
    0.79, 0.79, 0.79, 0.79, 0.78, 0.79, 0.78, 0.77, 0.77, 0.76, 0.76, 0.75, 
    0.75, 0.75, 0.82, 0.82, 0.82, 0.82, 0.81, 0.8, 0.8, 0.79, 0.79, 0.8, 0.8, 
    0.8, 0.81, 0.82, 0.84, 0.86, 0.86, 0.87, 0.87, 0.87, 0.87, 0.86, 0.85, 
    0.84, 0.84, 0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 0.84, 0.83, 0.82, 0.81, 
    0.8, 0.79, 0.79, 0.78, 0.77, 0.76, 0.76, 0.75, 0.73, 0.72, 0.69, 0.69, 
    0.69, 0.69, 0.68, 0.68, 0.67, 0.67, 0.68, 0.69, 0.69, 0.69, 0.69, 0.69, 
    0.71, 0.75, 0.78, 0.81, 0.82, 0.84, 0.86, 0.85, 0.84, 0.83, 0.83, 0.83, 
    0.84, 0.81, 0.84, 0.84, 0.82, 0.79, 0.81, 0.83, 0.84, 0.84, 0.86, 0.87, 
    0.89, 0.88, 0.9, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 
    0.9, 0.9, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.91, 0.91, 0.91, 0.94, 
    0.94, 0.95, 0.97, 0.96, 0.96, 0.95, 0.95, 0.94, 0.93, 0.91, 0.91, 0.9, 
    0.89, 0.88, 0.87, 0.87, 0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 0.85, 0.82, 
    0.82, 0.82, 0.82, 0.83, 0.84, 0.86, 0.87, 0.87, 0.87, 0.89, 0.92, 0.95, 
    0.91, 0.87, 0.88, 0.88, 0.89, 0.91, 0.92, 0.92, 0.93, 0.93, 0.94, 0.93, 
    0.93, 0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.94, 0.94, 
    0.93, 0.93, 0.91, 0.89, 0.88, 0.87, 0.85, 0.82, 0.81, 0.79, 0.78, 0.77, 
    0.76, 0.75, 0.72, 0.72, 0.75, 0.76, 0.77, 0.79, 0.78, 0.78, 0.78, 0.7, 
    0.71, 0.74, 0.74, 0.75, 0.74, 0.74, 0.76, 0.78, 0.79, 0.77, 0.76, 0.73, 
    0.72, 0.72, 0.73, 0.74, 0.76, 0.75, 0.76, 0.76, 0.76, 0.76, 0.76, 0.71, 
    0.73, 0.75, 0.75, 0.74, 0.76, 0.78, 0.8, 0.83, 0.85, 0.86, 0.88, 0.87, 
    0.88, 0.89, 0.9, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.93, 0.92, 0.9, 
    0.9, 0.91, 0.91, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.92, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 0.91, 0.89, 0.89, 0.87, 0.85, 0.83, 
    0.81, 0.8, 0.77, 0.76, 0.77, 0.76, 0.76, 0.74, 0.75, 0.75, 0.76, 0.76, 
    0.77, 0.78, 0.78, 0.8, 0.8, 0.81, 0.81, 0.82, 0.81, 0.8, 0.8, 0.78, 0.79, 
    0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.82, 0.82, 0.82, 0.81, 0.82, 
    0.82, 0.82, 0.81, 0.77, 0.73, 0.75, 0.78, 0.79, 0.8, 0.8, 0.78, 0.74, 
    0.71, 0.71, 0.74, 0.77, 0.79, 0.78, 0.74, 0.73, 0.74, 0.76, 0.83, 0.83, 
    0.85, 0.88, 0.88, 0.85, 0.84, 0.85, 0.87, 0.88, 0.88, 0.87, 0.86, 0.86, 
    0.86, 0.85, 0.82, 0.8, 0.81, 0.82, 0.83, 0.85, 0.86, 0.88, 0.89, 0.9, 
    0.9, 0.9, 0.91, 0.93, 0.95, 0.95, 0.92, 0.91, 0.95, 0.94, 0.92, 0.93, 
    0.92, 0.93, 0.88, 0.87, 0.88, 0.85, 0.89, 0.91, 0.9, 0.89, 0.89, 0.88, 
    0.9, 0.94, 0.94, 0.94, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.94, 0.94, 
    0.94, 0.95, 0.95, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.92, 0.86, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.87, 0.87, 0.91, 0.92, 
    0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 0.93, 0.93, 
    0.93, 0.92, 0.9, 0.88, 0.86, 0.85, 0.85, 0.86, 0.86, 0.86, 0.86, 0.87, 
    0.88, 0.88, 0.88, 0.89, 0.9, 0.92, 0.93, 0.92, 0.91, 0.9, 0.83, 0.84, 
    0.87, 0.89, 0.9, 0.88, 0.88, 0.87, 0.89, 0.91, 0.93, 0.94, 0.91, 0.93, 
    0.94, 0.95, 0.95, 0.94, 0.93, 0.93, 0.94, 0.94, 0.93, 0.93, 0.92, 0.91, 
    0.91, 0.91, 0.91, 0.93, 0.94, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.95, 0.96, 0.96, 0.95, 0.96, 0.97, 0.96, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.93, 0.92, 0.91, 0.91, 0.93, 0.94, 
    0.95, 0.92, 0.93, 0.94, 0.96, 0.97, 0.97, 0.97, 0.95, 0.94, 0.94, 0.93, 
    0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.95, 0.95, 0.94, 0.93, 
    0.92, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.91, 0.92, 0.92, 0.9, 
    0.9, 0.9, 0.95, 0.97, 0.96, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.97, 0.97, 0.96, 0.97, 0.96, 0.97, 0.97, 0.96, 0.97, 0.96, 0.97, 0.95, 
    0.93, 0.88, 0.86, 0.89, 0.85, 0.81, 0.79, 0.8, 0.8, 0.83, 0.83, 0.82, 
    0.81, 0.82, 0.83, 0.84, 0.84, 0.83, 0.82, 0.79, 0.77, 0.78, 0.81, 0.82, 
    0.83, 0.84, 0.85, 0.85, 0.83, 0.84, 0.85, 0.87, 0.89, 0.91, 0.89, 0.87, 
    0.89, 0.91, 0.91, 0.92, 0.94, 0.95, 0.96, 0.96, 0.96, 0.96, 0.94, 0.94, 
    0.94, 0.94, 0.93, 0.91, 0.91, 0.92, 0.93, 0.94, 0.93, 0.89, 0.8, 0.82, 
    0.85, 0.88, 0.9, 0.9, 0.9, 0.9, 0.89, 0.88, 0.88, 0.89, 0.9, 0.9, 0.89, 
    0.89, 0.89, 0.91, 0.92, 0.93, 0.93, 0.93, 0.92, 0.91, 0.92, 0.93, 0.93, 
    0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 0.93, 0.92, 0.92, 0.91, 0.91, 0.9, 
    0.9, 0.9, 0.9, 0.9, 0.89, 0.89, 0.9, 0.9, 0.9, 0.88, 0.89, 0.91, 0.91, 
    0.9, 0.9, 0.91, 0.91, 0.91, 0.9, 0.9, 0.86, 0.85, 0.86, 0.86, 0.86, 0.86, 
    0.87, 0.88, 0.88, 0.89, 0.9, 0.87, 0.87, 0.89, 0.9, 0.9, 0.9, 0.91, 0.91, 
    0.92, 0.91, 0.91, 0.92, 0.92, 0.92, 0.9, 0.9, 0.88, 0.84, 0.82, 0.82, 
    0.83, 0.84, 0.86, 0.88, 0.9, 0.9, 0.92, 0.93, 0.92, 0.91, 0.92, 0.93, 
    0.94, 0.94, 0.94, 0.95, 0.94, 0.92, 0.91, 0.89, 0.89, 0.9, 0.9, 0.9, 
    0.91, 0.89, 0.88, 0.88, 0.89, 0.9, 0.91, 0.92, 0.92, 0.9, 0.87, 0.89, 
    0.91, 0.91, 0.91, 0.91, 0.9, 0.89, 0.89, 0.86, 0.85, 0.84, 0.84, 0.85, 
    0.84, 0.85, 0.87, 0.88, 0.89, 0.89, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 
    0.92, 0.92, 0.91, 0.9, 0.9, 0.89, 0.87, 0.86, 0.86, 0.87, 0.88, 0.87, 
    0.85, 0.85, 0.86, 0.88, 0.88, 0.88, 0.88, 0.9, 0.89, 0.88, 0.9, 0.91, 
    0.92, 0.92, 0.93, 0.93, 0.94, 0.94, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 
    0.93, 0.93, 0.94, 0.94, 0.95, 0.95, 0.95, 0.96, 0.96, 0.95, 0.96, 0.96, 
    0.95, 0.96, 0.95, 0.94, 0.93, 0.93, 0.92, 0.9, 0.9, 0.94, 0.96, 0.96, 
    0.96, 0.95, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.94, 0.93, 0.93, 0.92, 0.94, 0.96, 0.95, 0.95, 0.96, 0.97, 0.97, 
    0.97, 0.97, 0.96, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.95, 0.95, 0.94, 0.94, 0.93, 0.92, 
    0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 0.93, 0.94, 0.94, 0.95, 0.95, 0.95, 
    0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 0.96, 0.95, 0.94, 0.95, 0.95, 0.95, 
    0.95, 0.96, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.95, 0.96, 0.97, 0.97, 0.96, 0.96, 0.94, 0.94, 0.95, 0.98, 
    0.98, 0.93, 0.89, 0.89, 0.89, 0.88, 0.92, 0.91, 0.92, 0.92, 0.91, 0.91, 
    0.91, 0.91, 0.89, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.91, 0.91, 0.92, 
    0.92, 0.92, 0.92, 0.91, 0.89, 0.87, 0.9, 0.9, 0.9, 0.89, 0.9, 0.95, 0.96, 
    0.96, 0.97, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.93, 0.94, 0.94, 0.93, 0.93, 0.92, 0.92, 0.92, 
    0.93, 0.92, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.94, 0.94, 0.95, 0.94, 
    0.96, 0.97, 0.96, 0.96, 0.95, 0.96, 0.95, 0.95, 0.95, 0.94, 0.94, 0.95, 
    0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.96, 0.97, 
    0.96, 0.97, 0.95, 0.92, 0.92, 0.92, 0.91, 0.92, 0.92, 0.92, 0.92, 0.92, 
    0.93, 0.93, 0.94, 0.93, 0.94, 0.93, 0.94, 0.95, 0.96, 0.97, 0.98, 0.97, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.94, 0.95, 
    0.95, 0.95, 0.95, 0.94, 0.93, 0.92, 0.92, 0.93, 0.94, 0.93, 0.94, 0.95, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 
    0.97, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.94, 0.94, 0.94, 0.92, 0.91, 0.97, 0.96, 0.94, 0.91, 0.93, 0.94, 0.95, 
    0.94, 0.94, 0.93, 0.92, 0.91, 0.93, 0.92, 0.91, 0.9, 0.89, 0.88, 0.87, 
    0.85, 0.83, 0.83, 0.84, 0.83, 0.88, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 
    0.92, 0.93, 0.92, 0.91, 0.9, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 
    0.93, 0.94, 0.96, 0.96, 0.95, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.96, 0.95, 0.94, 0.93, 0.92, 
    0.91, 0.91, 0.94, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.95, 0.95, 0.95, 0.92, 0.94, 0.95, 0.95, 0.94, 0.94, 0.93, 0.92, 0.91, 
    0.94, 0.95, 0.95, 0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 
    0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.94, 0.93, 0.93, 0.92, 0.94, 0.94, 
    0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 0.97, 
    0.97, 0.96, 0.95, 0.96, 0.95, 0.91, 0.91, 0.92, 0.91, 0.89, 0.89, 0.91, 
    0.89, 0.87, 0.87, 0.87, 0.86, 0.92, 0.94, 0.94, 0.93, 0.94, 0.94, 0.95, 
    0.95, 0.96, 0.95, 0.96, 0.96, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.92, 
    0.92, 0.91, 0.91, 0.91, 0.92, 0.97, 0.96, 0.95, 0.95, 0.95, 0.95, 0.96, 
    0.97, 0.97, 0.96, 0.95, 0.94, 0.94, 0.93, 0.91, 0.89, 0.89, 0.9, 0.91, 
    0.9, 0.9, 0.9, 0.91, 0.92, 0.91, 0.92, 0.93, 0.93, 0.94, 0.93, 0.94, 
    0.93, 0.91, 0.91, 0.91, 0.92, 0.9, 0.89, 0.89, 0.87, 0.88, 0.89, 0.89, 
    0.89, 0.89, 0.9, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 
    0.91, 0.91, 0.91, 0.9, 0.89, 0.86, 0.83, 0.81, 0.79, 0.77, 0.76, 0.75, 
    0.76, 0.76, 0.78, 0.88, 0.93, 0.87, 0.85, 0.83, 0.83, 0.84, 0.84, 0.84, 
    0.85, 0.86, 0.86, 0.86, 0.86, 0.84, 0.84, 0.85, 0.86, 0.86, 0.85, 0.84, 
    0.84, 0.85, 0.84, 0.85, 0.86, 0.89, 0.89, 0.88, 0.87, 0.88, 0.87, 0.87, 
    0.87, 0.86, 0.86, 0.85, 0.85, 0.86, 0.84, 0.84, 0.85, 0.86, 0.87, 0.88, 
    0.88, 0.89, 0.89, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 0.91, 0.91, 
    0.91, 0.91, 0.91, 0.9, 0.89, 0.91, 0.91, 0.9, 0.88, 0.87, 0.88, 0.88, 
    0.89, 0.9, 0.92, 0.93, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 0.94, 
    0.94, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.9, 0.89, 0.89, 0.89, 0.89, 
    0.89, 0.89, 0.89, 0.9, 0.91, 0.93, 0.93, 0.93, 0.93, 0.92, 0.93, 0.92, 
    0.92, 0.91, 0.92, 0.92, 0.9, 0.87, 0.83, 0.82, 0.83, 0.83, 0.84, 0.85, 
    0.85, 0.85, 0.86, 0.88, 0.89, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.95, 0.97, 0.97, 0.92, 0.93, 0.92, 0.93, 0.93, 0.95, 0.95, 
    0.94, 0.94, 0.95, 0.94, 0.94, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.95, 
    0.95, 0.96, 0.97, 0.97, 0.95, 0.93, 0.93, 0.92, 0.91, 0.91, 0.91, 0.91, 
    0.92, 0.91, 0.91, 0.91, 0.91, 0.95, 0.95, 0.94, 0.95, 0.94, 0.95, 0.95, 
    0.95, 0.95, 0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 
    0.92, 0.94, 0.94, 0.95, 0.94, 0.95, 0.97, 0.98, 0.98, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.96, 0.97, 0.96, 0.96, 
    0.95, 0.94, 0.93, 0.94, 0.95, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 
    0.93, 0.92, 0.92, 0.91, 0.91, 0.92, 0.93, 0.93, 0.94, 0.95, 0.95, 0.95, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.93, 0.91, 0.89, 0.87, 0.85, 0.84, 
    0.85, 0.86, 0.87, 0.86, 0.83, 0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 0.92, 
    0.9, 0.89, 0.89, 0.87, 0.85, 0.92, 0.92, 0.92, 0.93, 0.93, 0.92, 0.91, 
    0.91, 0.91, 0.91, 0.91, 0.92, 0.95, 0.95, 0.95, 0.96, 0.96, 0.97, 0.96, 
    0.95, 0.95, 0.96, 0.96, 0.96, 0.91, 0.91, 0.91, 0.9, 0.9, 0.88, 0.87, 
    0.87, 0.88, 0.88, 0.9, 0.91, 0.94, 0.95, 0.96, 0.97, 0.96, 0.95, 0.94, 
    0.94, 0.94, 0.93, 0.93, 0.93, 0.96, 0.95, 0.95, 0.95, 0.93, 0.92, 0.9, 
    0.9, 0.92, 0.93, 0.92, 0.9, 0.93, 0.92, 0.91, 0.9, 0.89, 0.89, 0.89, 0.9, 
    0.89, 0.86, 0.87, 0.88, 0.9, 0.91, 0.93, 0.94, 0.94, 0.94, 0.93, 0.92, 
    0.91, 0.93, 0.94, 0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.96, 0.96, 0.95, 0.96, 0.95, 0.95, 0.95, 0.93, 0.93, 0.93, 0.94, 
    0.94, 0.95, 0.95, 0.95, 0.92, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 
    0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.92, 0.92, 0.94, 0.92, 0.92, 0.95, 
    0.95, 0.94, 0.93, 0.94, 0.93, 0.95, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.96, 0.95, 0.93, 0.93, 0.94, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.93, 0.95, 0.96, 0.96, 0.95, 0.95, 
    0.95, 0.94, 0.91, 0.9, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.89, 0.89, 0.91, 
    0.93, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 
    0.95, 0.94, 0.94, 0.92, 0.94, 0.95, 0.96, 0.95, 0.95, 0.95, 0.96, 0.96, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 
    0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.92, 0.93, 0.92, 0.92, 0.91, 0.91, 0.9, 0.89, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.88, 0.77, 0.76, 0.75, 0.74, 0.74, 0.75, 0.78, 0.78, 0.79, 
    0.79, 0.76, 0.74, 0.74, 0.74, 0.73, 0.74, 0.74, 0.74, 0.74, 0.74, 0.74, 
    0.76, 0.78, 0.81, 0.8, 0.82, 0.87, 0.91, 0.94, 0.96, 0.98, 0.99, 0.96, 
    0.92, 0.88, 0.86, _, 0.81, 0.81, 0.81, 0.8, 0.79, 0.79, 0.79, 0.8, 0.82, 
    0.82, 0.83, _, 0.79, 0.78, 0.77, 0.77, 0.76, 0.73, 0.71, 0.7, 0.7, 0.7, 
    0.69, 0.67, 0.68, 0.69, 0.72, 0.75, 0.74, 0.72, 0.74, 0.77, 0.78, 0.79, 
    0.81, 0.82, 0.84, 0.88, 0.93, 0.96, 0.96, 0.98, 0.98, 0.97, 0.97, 0.95, 
    0.91, 0.94, 0.94, 0.94, 0.95, 0.94, 0.93, 0.93, 0.94, 0.95, 0.95, 0.95, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 
    0.93, 0.84, 0.83, 0.82, 0.78, 0.75, 0.73, 0.72, 0.7, 0.69, 0.71, 0.71, 
    0.73, 0.74, 0.75, 0.77, 0.78, 0.79, 0.79, 0.8, 0.78, 0.78, 0.78, 0.78, 
    0.78, 0.74, 0.71, 0.68, 0.68, 0.69, 0.66, 0.67, 0.69, 0.72, 0.7, 0.71, 
    0.72, 0.81, 0.82, 0.83, 0.84, 0.83, 0.79, 0.76, 0.72, 0.71, 0.71, 0.72, 
    0.73, 0.78, 0.79, 0.83, 0.83, 0.84, 0.85, 0.77, 0.77, 0.79, 0.76, 0.74, 
    0.74, 0.72, 0.8, 0.81, 0.85, 0.85, 0.81, 0.82, 0.79, 0.8, 0.79, 0.82, 
    0.85, 0.76, 0.76, 0.74, 0.71, 0.71, 0.69, 0.68, 0.67, 0.72, 0.75, 0.75, 
    0.74, 0.79, 0.8, 0.81, 0.83, 0.84, 0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 
    0.88, 0.87, 0.88, 0.88, 0.88, 0.89, 0.88, 0.86, 0.84, 0.82, 0.81, 0.8, 
    0.81, 0.94, 0.95, 0.95, 0.96, 0.95, 0.95, 0.97, 0.93, 0.89, 0.87, 0.84, 
    0.81, 0.85, 0.85, 0.84, 0.83, 0.8, 0.78, 0.76, 0.77, 0.8, 0.84, 0.87, 
    0.86, 0.86, 0.87, 0.88, 0.87, 0.88, 0.87, 0.86, 0.85, 0.83, 0.8, 0.82, 
    0.84, 0.8, 0.78, 0.77, 0.77, 0.77, 0.77, 0.76, 0.76, 0.74, 0.76, 0.86, 
    0.84, 0.86, 0.87, 0.92, 0.93, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 
    0.95, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 
    0.95, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.97, 0.96, 0.97, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 
    0.97, 0.97, 0.95, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 
    0.97, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.97, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 
    0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.94, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.97, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 
    0.97, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.91, 0.9, 0.9, 0.92, 0.94, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.95, 0.94, 
    0.93, 0.96, 0.95, 0.92, 0.91, 0.89, 0.86, 0.88, 0.9, 0.92, 0.91, 0.92, 
    0.94, 0.92, 0.93, 0.96, 0.97, 0.98, 0.97, 0.94, 0.9, 0.88, 0.85, 0.8, 
    0.75, 0.81, 0.8, 0.79, 0.79, 0.79, 0.8, 0.81, 0.82, 0.84, 0.86, 0.89, 
    0.92, 0.94, 0.93, 0.9, 0.87, 0.86, 0.88, 0.88, 0.88, 0.92, 0.94, 0.94, 
    0.97, 0.91, 0.9, 0.91, 0.89, 0.91, 0.91, 0.93, 0.92, 0.91, 0.93, 0.94, 
    0.93, 0.96, 0.95, 0.9, 0.87, 0.87, 0.83, 0.84, 0.88, 0.91, 0.9, 0.88, 
    0.88, 0.89, 0.89, 0.9, 0.91, 0.92, 0.92, 0.93, 0.95, 0.96, 0.97, 0.97, 
    0.97, 0.97, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 
    0.95, 0.94, 0.93, 0.93, 0.92, 0.92, 0.91, 0.91, 0.9, 0.9, 0.89, 0.89, 
    0.9, 0.91, 0.92, 0.92, 0.91, 0.89, 0.87, 0.85, 0.85, 0.87, 0.89, 0.9, 
    0.9, 0.89, 0.9, 0.91, 0.91, 0.92, 0.93, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.97, 0.97, 0.96, 
    0.95, 0.92, 0.89, 0.85, 0.85, 0.88, 0.88, 0.88, 0.88, 0.89, 0.89, 0.89, 
    0.9, 0.94, 0.93, 0.92, 0.91, 0.92, 0.92, 0.93, 0.94, 0.94, 0.94, 0.93, 
    0.92, 0.89, 0.89, 0.89, 0.89, 0.87, 0.86, 0.84, 0.84, 0.87, 0.88, 0.88, 
    0.86, 0.84, 0.86, 0.87, 0.89, 0.86, 0.86, 0.87, 0.86, 0.84, 0.85, 0.87, 
    0.87, 0.87, 0.88, 0.88, 0.88, 0.89, 0.89, 0.9, 0.9, 0.91, 0.92, 0.92, 
    0.92, 0.94, 0.94, 0.94, 0.93, 0.93, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 
    0.89, 0.87, 0.85, 0.82, 0.81, 0.8, 0.8, 0.8, 0.8, 0.78, 0.77, 0.78, 0.79, 
    0.84, 0.84, 0.86, 0.89, 0.89, 0.9, 0.89, 0.89, 0.89, 0.89, 0.88, 0.87, 
    0.88, 0.89, 0.9, 0.94, 0.96, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.95, 
    0.96, 0.98, 0.97, 0.96, 0.99, 0.98, 0.98, 0.97, 0.96, 0.95, 0.94, 0.93, 
    0.89, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.93, 0.94, 0.91, 0.92, 0.93, 
    0.96, 0.97, 0.96, 0.96, 0.97, 0.96, 0.98, 0.99, 0.98, 0.94, 0.94, 0.94, 
    0.96, 0.95, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 
    0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.97, 0.97, 0.96, 0.96, 0.94, 0.94, 0.93, 0.93, 
    0.98, 0.99, 0.99, 1, 0.99, 0.98, 0.98, 0.97, 0.98, 0.98, 0.97, 0.97, 
    0.95, 0.95, 0.94, 0.95, 0.95, 0.94, 0.94, 0.95, 0.96, 0.97, 0.96, 0.96, 
    0.96, 0.94, 0.95, 0.96, 0.98, 1, 0.99, 0.99, 0.98, 0.96, 0.95, 0.94, 
    0.93, 0.93, 0.93, 0.92, 0.93, 0.88, 0.86, 0.82, 0.8, 0.87, 0.87, 0.8, 
    0.78, 0.83, 0.87, 0.88, 0.88, 0.88, 0.89, 0.92, 0.94, 0.96, 0.96, 0.97, 
    0.98, 0.96, 0.94, 0.94, 0.92, 0.9, 0.88, 0.86, 0.84, 0.83, 0.91, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.96, 0.95, 0.96, 0.98, 0.99, 1, 1, 1, 1, 0.99, 
    0.97, 0.95, 0.95, 0.97, 0.98, 0.96, 0.93, 0.92, 0.91, 0.94, 0.77, 0.73, 
    0.74, 0.8, 0.8, 0.82, 0.81, 0.83, 0.84, 0.85, 0.87, 0.88, 0.85, 0.84, 
    0.81, 0.78, 0.75, 0.71, 0.67, 0.68, 0.69, 0.68, 0.67, 0.67, 0.74, 0.78, 
    0.85, 0.88, 0.9, 0.83, 0.83, 0.84, 0.84, 0.72, 0.71, 0.72, 0.83, 0.83, 
    0.84, 0.84, 0.85, 0.86, 0.86, 0.88, 0.88, 0.88, 0.89, 0.89, 0.88, 0.89, 
    0.87, 0.88, 0.88, 0.89, 0.86, 0.87, 0.86, 0.86, 0.87, 0.88, 0.78, 0.76, 
    0.76, 0.75, 0.74, 0.74, 0.75, 0.76, 0.81, 0.84, 0.87, 0.88, 0.87, 0.86, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.89, 0.91, 0.89, 0.86, 0.81, 0.8, 
    0.8, 0.81, 0.82, 0.83, 0.78, 0.76, 0.78, 0.79, 0.82, 0.82, 0.87, 0.87, 
    0.88, 0.86, 0.9, 0.92, 0.95, 0.94, 0.92, 0.92, 0.92, 0.92, 0.95, 0.96, 
    0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.97, 0.99, 0.98, 
    0.98, 0.99, 0.99, 0.98, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 0.97, 0.97, 0.96, 0.94, 0.96, 0.96, 
    0.95, 0.98, 0.98, 0.98, 0.97, 0.95, 0.93, 0.9, 0.9, 0.9, 0.85, 0.83, 
    0.82, 0.82, 0.8, 0.82, 0.85, 0.89, 0.88, 0.88, 0.87, 0.9, 0.95, 0.96, 
    0.96, 0.91, 0.88, 0.83, 0.82, 0.82, 0.82, 0.83, 0.86, 0.86, 0.85, 0.86, 
    0.88, 0.9, 0.92, 0.94, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 
    0.94, 0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 0.95, 
    0.95, 0.94, 0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.95, 0.95, 
    0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 0.94, 0.93, 
    0.93, 0.93, 0.93, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.97, 0.94, 0.93, 
    0.92, 0.92, 0.92, 0.92, 0.93, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.91, 
    0.91, 0.9, 0.88, 0.86, 0.83, 0.8, 0.79, 0.8, 0.8, 0.81, 0.72, 0.71, 0.72, 
    0.73, 0.73, 0.75, 0.76, 0.79, 0.79, 0.82, 0.87, 0.93, 0.83, 0.81, 0.86, 
    0.82, 0.84, 0.85, 0.83, 0.85, 0.86, 0.86, 0.88, 0.89, 0.96, 0.95, 0.95, 
    0.93, 0.87, 0.88, 0.9, 0.9, 0.88, 0.88, 0.89, 0.9, 0.84, 0.84, 0.83, 
    0.83, 0.82, 0.82, 0.82, 0.8, 0.81, 0.89, 0.94, 0.93, 0.97, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.93, 0.95, 0.93, 0.91, 
    0.9, 0.91, 0.91, 0.92, 0.94, 0.95, 0.97, 0.99, 0.99, 0.97, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.98, 0.97, 
    0.96, 0.95, 0.94, 0.92, 0.89, 0.87, 0.85, 0.84, 0.83, 0.99, 0.97, 0.97, 
    0.97, 0.96, 0.94, 0.91, 0.89, 0.87, 0.85, 0.8, 0.69, 0.79, 0.8, 0.82, 
    0.84, 0.77, 0.69, 0.69, 0.7, 0.75, 0.83, 0.88, 0.9, 0.97, 0.96, 0.97, 
    0.96, 0.94, 0.96, 0.95, 0.97, 0.99, 0.89, 0.85, 0.88, 0.92, 0.9, 0.9, 
    0.92, 0.95, 0.97, 0.98, 0.98, 0.99, 0.99, 0.98, 0.96, 0.99, 0.99, 0.99, 
    0.98, 0.98, 0.98, 0.98, 0.98, 1, 1, 0.98, 0.98, 0.94, 1, 0.94, 0.98, 
    0.96, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.98, 0.97, 0.98, 
    0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.99, 0.99, 0.99, 
    0.98, 0.94, 0.95, 0.99, 0.97, 0.96, 0.98, 0.97, 0.99, 0.99, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.99, 0.98, 0.96, 0.98, 0.97, 0.96, 
    0.96, 0.96, 0.95, 0.97, 0.96, 0.97, 0.98, 0.97, 0.96, 0.96, 0.94, 0.93, 
    0.91, 0.9, 0.93, 0.93, 0.93, 0.93, 0.92, 0.93, 0.93, 0.92, 0.91, 0.92, 
    0.92, 0.92, 0.9, 0.92, 0.93, 0.98, 0.98, 0.97, 0.96, 0.96, 0.98, 0.98, 
    0.98, 0.98, 0.99, 0.99, 0.98, 0.92, 0.93, 0.84, 0.8, 0.79, 0.8, 0.8, 
    0.85, 0.92, 0.94, 0.94, 0.94, 0.93, 0.94, 0.93, 0.94, 0.95, 0.99, 0.99, 
    0.97, 0.95, 0.93, 0.89, 0.86, 0.93, 0.98, 1, 0.81, 0.84, 0.76, 0.72, 
    0.72, 0.76, 0.79, 0.79, 0.81, 0.79, 0.78, 0.81, 0.8, 0.78, 0.8, 0.81, 
    0.82, 0.87, 0.79, 0.77, 0.77, 0.76, 0.76, 0.77, 0.78, 0.77, 0.77, 0.77, 
    0.78, 0.79, 0.79, 0.78, 0.79, 0.79, 0.79, 0.8, 0.8, 0.81, 0.81, 0.81, 
    0.81, 0.82, 0.82, 0.83, 0.84, 0.84, 0.86, 0.83, 0.78, 0.85, 0.81, 0.83, 
    0.83, 0.82, 0.8, 0.8, 0.8, 0.78, 0.78, 0.78, 0.79, 0.78, 0.77, 0.77, 
    0.76, 0.76, 0.75, 0.74, 0.71, 0.67, 0.66, 0.65, 0.64, 0.64, 0.64, 0.64, 
    0.63, 0.62, 0.62, 0.63, 0.62, 0.61, 0.61, 0.61, 0.61, 0.61, 0.6, 0.61, 
    0.61, 0.61, 0.62, 0.61, 0.61, 0.62, 0.63, 0.63, 0.6, 0.61, 0.61, 0.61, 
    0.59, 0.59, 0.58, 0.57, 0.57, 0.58, 0.58, 0.58, 0.61, 0.61, 0.6, 0.6, 
    0.59, 0.57, 0.55, 0.55, 0.55, 0.54, 0.54, 0.54, 0.76, 0.77, 0.77, 0.75, 
    0.76, 0.76, 0.78, 0.79, 0.8, 0.8, 0.79, 0.77, 0.71, 0.68, 0.66, 0.67, 
    0.67, 0.72, 0.74, 0.75, 0.74, 0.73, 0.77, 0.81, 0.75, 0.75, 0.73, 0.75, 
    0.76, 0.74, 0.74, 0.77, 0.81, 0.78, 0.78, 0.82, 0.89, 0.9, 0.91, 0.92, 
    0.91, 0.91, 0.91, 0.93, 0.93, 0.91, 0.91, 0.93, 0.95, 0.95, 0.97, 0.99, 
    0.99, 0.97, 0.95, 0.96, 0.96, 0.97, 0.97, 0.96, 0.94, 0.93, 0.94, 0.95, 
    0.95, 0.94, 0.94, 0.91, 0.88, 0.87, 0.86, 0.85, 0.86, 0.83, 0.83, 0.84, 
    0.86, 0.87, 0.86, 0.86, 0.86, 0.87, 0.89, 0.89, 0.88, 0.89, 0.88, 0.88, 
    0.88, 0.88, 0.89, 0.88, 0.86, 0.86, 0.86, 0.87, 0.89, 0.89, 0.88, 0.87, 
    0.86, 0.85, 0.84, 0.84, 0.83, 0.8, 0.75, 0.75, 0.73, 0.71, 0.71, 0.72, 
    0.72, 0.73, 0.72, 0.73, 0.7, 0.73, 0.81, 0.78, 0.85, 0.84, 0.85, 0.86, 
    0.87, 0.86, 0.87, 0.84, 0.79, 0.74, 0.76, 0.74, 0.85, 0.86, 0.87, 0.9, 
    0.93, 0.95, 0.95, 0.96, 0.97, 0.97, 0.89, 0.87, 0.76, 0.75, 0.75, 0.77, 
    0.81, 0.84, 0.86, 0.87, 0.84, 0.8, 0.82, 0.81, 0.81, 0.8, 0.79, 0.79, 
    0.77, 0.79, 0.81, 0.84, 0.83, 0.81, 0.79, 0.76, 0.81, 0.82, 0.81, 0.77, 
    0.78, 0.79, 0.77, 0.74, 0.72, 0.7, 0.68, 0.65, 0.7, 0.72, 0.73, 0.75, 
    0.76, 0.77, 0.77, 0.75, 0.76, 0.83, 0.85, 0.85, 0.77, 0.83, 0.86, 0.86, 
    0.85, 0.81, 0.79, 0.77, 0.71, 0.75, 0.79, 0.77, 0.75, 0.7, 0.68, 0.68, 
    0.7, 0.77, 0.77, 0.74, 0.71, 0.69, 0.68, 0.69, 0.68, 0.69, 0.72, 0.74, 
    0.77, 0.79, 0.81, 0.8, 0.8, 0.78, 0.75, 0.77, 0.85, 0.88, 0.9, 0.96, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.95, 0.97, 
    0.99, 0.95, 0.94, 0.94, 0.93, 0.91, 0.91, 0.93, 0.76, 0.74, 0.74, 0.73, 
    0.69, 0.68, 0.67, 0.66, 0.66, 0.66, 0.67, 0.67, 0.65, 0.67, 0.67, 0.69, 
    0.69, 0.68, 0.68, 0.69, 0.69, 0.7, 0.71, 0.71, 0.68, 0.68, 0.67, 0.67, 
    0.67, 0.66, 0.66, 0.66, 0.65, 0.65, 0.65, 0.66, 0.62, 0.63, 0.63, 0.65, 
    0.66, 0.67, 0.68, 0.69, 0.69, 0.7, 0.7, 0.71, 0.71, 0.71, 0.72, 0.71, 
    0.72, 0.71, 0.72, 0.68, 0.66, 0.71, 0.78, 0.8, 0.72, 0.77, 0.81, 0.81, 
    0.82, 0.82, 0.79, 0.76, 0.8, 0.75, 0.73, 0.75, 0.81, 0.83, 0.81, 0.79, 
    0.75, 0.72, 0.72, 0.73, 0.74, 0.74, 0.73, 0.73, 0.71, 0.72, 0.72, 0.75, 
    0.76, 0.76, 0.77, 0.78, 0.76, 0.78, 0.76, 0.75, 0.74, 0.72, 0.71, 0.71, 
    0.72, 0.75, 0.78, 0.77, 0.74, 0.71, 0.71, 0.7, 0.68, 0.68, 0.68, 0.68, 
    0.68, 0.66, 0.67, 0.67, 0.66, 0.66, 0.67, 0.66, 0.67, 0.67, 0.67, 0.67, 
    0.68, 0.67, 0.67, 0.68, 0.68, 0.68, 0.69, 0.69, 0.71, 0.71, 0.71, 0.7, 
    0.7, 0.7, 0.69, 0.67, 0.67, 0.66, 0.67, 0.67, 0.67, 0.68, 0.67, 0.68, 
    0.68, 0.69, 0.7, 0.7, 0.71, 0.7, 0.7, 0.7, 0.73, 0.71, 0.72, 0.71, 0.71, 
    0.72, 0.72, 0.72, 0.73, 0.74, 0.74, 0.74, 0.75, 0.74, 0.74, 0.72, 0.72, 
    0.74, 0.75, 0.73, 0.72, 0.72, 0.72, 0.71, 0.73, 0.73, 0.74, 0.75, 0.77, 
    0.78, 0.78, 0.78, 0.77, 0.78, 0.78, 0.79, 0.78, 0.77, 0.77, 0.77, 0.77, 
    0.77, 0.75, 0.75, 0.76, 0.77, 0.75, 0.73, 0.72, 0.73, 0.74, 0.77, 0.79, 
    0.81, 0.83, 0.83, 0.84, 0.85, 0.86, 0.88, 0.88, 0.9, 0.91, 0.93, 0.92, 
    0.92, 0.93, 0.94, 0.94, 0.94, 0.93, 0.93, 0.88, 0.89, 0.9, 0.91, 0.93, 
    0.95, 0.96, 0.96, 0.96, 0.95, 0.94, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.89, 0.89, 0.89, 0.89, 0.87, 
    0.87, 0.87, 0.87, 0.88, 0.88, 0.9, 0.92, 0.78, 0.78, 0.78, 0.78, 0.77, 
    0.8, 0.82, 0.82, 0.83, 0.83, 0.83, 0.84, 0.71, 0.69, 0.69, 0.69, 0.71, 
    0.72, 0.72, 0.7, 0.72, 0.73, 0.77, 0.76, 0.77, 0.77, 0.73, 0.76, 0.83, 
    0.86, 0.83, 0.79, 0.75, 0.74, 0.74, 0.75, 0.77, 0.78, 0.78, 0.78, 0.78, 
    0.78, 0.77, 0.77, 0.76, 0.75, 0.75, 0.74, 0.74, 0.74, 0.73, 0.72, 0.71, 
    0.7, 0.7, 0.7, 0.69, 0.69, 0.7, 0.7, 0.7, 0.7, 0.71, 0.73, 0.73, 0.7, 
    0.67, 0.66, 0.65, 0.64, 0.63, 0.63, 0.63, 0.61, 0.61, 0.61, 0.6, 0.6, 
    0.63, 0.64, 0.65, 0.68, 0.7, 0.68, 0.67, 0.68, 0.68, 0.69, 0.69, 0.72, 
    0.72, 0.72, 0.72, 0.74, 0.76, 0.77, 0.76, 0.77, 0.76, 0.77, 0.76, 0.77, 
    0.77, 0.8, 0.81, 0.81, 0.82, 0.83, 0.85, 0.85, 0.87, 0.87, 0.88, 0.93, 
    0.94, 0.94, 0.94, 0.93, 0.93, 0.94, 0.89, 0.92, 0.93, 0.92, 0.93, 0.94, 
    0.9, 0.87, 0.86, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.82, 0.85, 0.86, 
    0.86, 0.86, 0.86, 0.87, 0.86, 0.86, 0.84, 0.83, 0.82, 0.82, 0.83, 0.83, 
    0.82, 0.82, 0.81, 0.8, 0.81, 0.8, 0.81, 0.83, 0.85, 0.86, 0.86, 0.87, 
    0.88, 0.9, 0.93, 0.93, 0.95, 0.94, 0.96, 0.96, 0.96, 0.97, 0.98, 0.98, 
    0.95, 0.95, 0.96, 0.97, 0.88, 0.79, 0.91, 0.89, 0.89, 0.8, 0.8, 0.82, 
    0.77, 0.79, 0.81, 0.81, 0.79, 0.72, 0.73, 0.74, 0.73, 0.76, 0.79, 0.81, 
    0.77, 0.73, 0.72, 0.71, 0.69, 0.66, 0.66, 0.71, 0.69, 0.67, 0.67, 0.64, 
    0.66, 0.66, 0.64, 0.66, 0.65, 0.65, 0.64, 0.63, 0.6, 0.63, 0.7, 0.8, 
    0.85, 0.86, 0.81, 0.77, 0.74, 0.73, 0.71, 0.7, 0.71, 0.74, 0.73, 0.74, 
    0.74, 0.76, 0.76, 0.77, 0.78, 0.77, 0.76, 0.74, 0.74, 0.73, 0.71, 0.69, 
    0.68, 0.66, 0.65, 0.64, 0.65, 0.65, 0.63, 0.65, 0.67, 0.69, 0.71, 0.71, 
    0.71, 0.69, 0.68, 0.67, 0.68, 0.7, 0.64, 0.65, 0.68, 0.69, 0.73, 0.74, 
    0.73, 0.76, 0.76, 0.75, 0.72, 0.74, 0.74, 0.72, 0.74, 0.75, 0.76, 0.77, 
    0.78, 0.79, 0.81, 0.82, 0.84, 0.85, 0.82, 0.81, 0.79, 0.79, 0.82, 0.88, 
    0.88, 0.9, 0.91, 0.92, 0.93, 0.95, 0.96, 0.97, 0.98, 0.99, 0.92, 0.9, 
    0.88, 0.86, 0.84, 0.84, 0.83, 0.81, 0.84, 0.8, 0.8, 0.78, 0.76, 0.74, 
    0.73, 0.72, 0.71, 0.69, 0.7, 0.68, 0.67, 0.64, 0.62, 0.62, 0.62, 0.62, 
    0.64, 0.64, 0.63, 0.63, 0.64, 0.65, 0.68, 0.69, 0.67, 0.7, 0.71, 0.67, 
    0.65, 0.68, 0.74, 0.79, 0.77, 0.77, 0.82, 0.82, 0.79, 0.78, 0.8, 0.8, 
    0.8, 0.79, 0.79, 0.79, 0.79, 0.8, 0.8, 0.8, 0.8, 0.78, 0.78, 0.79, 0.79, 
    0.79, 0.78, 0.77, 0.75, 0.74, 0.77, 0.76, 0.75, 0.74, 0.73, 0.72, 0.71, 
    0.69, 0.69, 0.68, 0.67, 0.65, 0.66, 0.67, 0.66, 0.68, 0.73, 0.76, 0.77, 
    0.77, 0.78, 0.78, 0.77, 0.78, 0.81, 0.8, 0.8, 0.8, 0.79, 0.82, 0.83, 
    0.83, 0.82, 0.83, 0.84, 0.85, 0.85, 0.85, 0.88, 0.92, 0.94, 0.94, 0.95, 
    0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.95, 0.91, 0.89, 0.89, 0.89, 0.89, 
    0.89, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 0.94, 0.98, 0.98, 0.98, 
    0.95, 0.93, 0.92, 0.93, 0.94, 0.92, 0.91, 0.91, 0.91, 0.92, 0.91, 0.89, 
    0.9, 0.89, 0.87, 0.87, 0.86, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.83, 
    0.83, 0.83, 0.83, 0.84, 0.85, 0.83, 0.84, 0.87, 0.87, 0.86, 0.85, 0.85, 
    0.85, 0.84, 0.85, 0.88, 0.89, 0.82, 0.81, 0.81, 0.83, 0.82, 0.83, 0.83, 
    0.84, 0.83, 0.81, 0.81, 0.82, 0.85, 0.83, 0.86, 0.86, 0.88, 0.9, 0.92, 
    0.95, 0.98, 0.97, 0.98, 0.98, 0.85, 0.87, 0.81, 0.79, 0.75, 0.71, 0.7, 
    0.69, 0.68, 0.68, 0.68, 0.68, 0.66, 0.65, 0.65, 0.65, 0.65, 0.65, 0.65, 
    0.65, 0.64, 0.64, 0.63, 0.64, 0.63, 0.63, 0.64, 0.63, 0.62, 0.61, 0.61, 
    0.62, 0.63, 0.64, 0.66, 0.68, 0.71, 0.73, 0.73, 0.7, 0.64, 0.64, 0.66, 
    0.73, 0.78, 0.81, 0.83, 0.83, 0.85, 0.91, 0.92, 0.85, 0.83, 0.83, 0.82, 
    0.83, 0.85, 0.83, 0.82, 0.81, 0.89, 0.88, 0.85, 0.84, 0.84, 0.86, 0.87, 
    0.87, 0.86, 0.85, 0.83, 0.83, 0.86, 0.86, 0.87, 0.87, 0.89, 0.89, 0.88, 
    0.9, 0.9, 0.91, 0.9, 0.89, 0.89, 0.89, 0.88, 0.88, 0.88, 0.88, 0.9, 0.9, 
    0.89, 0.88, 0.88, 0.87, 0.89, 0.88, 0.87, 0.88, 0.87, 0.86, 0.86, 0.86, 
    0.86, 0.87, 0.88, 0.87, 0.86, 0.85, 0.85, 0.84, 0.83, 0.81, 0.8, 0.79, 
    0.78, 0.76, 0.76, 0.78, 0.78, 0.77, 0.77, 0.79, 0.77, 0.75, 0.74, 0.75, 
    0.75, 0.75, 0.75, 0.74, 0.75, 0.74, 0.74, 0.75, 0.75, 0.75, 0.75, 0.75, 
    0.74, 0.74, 0.75, 0.75, 0.75, 0.74, 0.74, 0.74, 0.74, 0.73, 0.73, 0.73, 
    0.73, 0.72, 0.72, 0.71, 0.7, 0.7, 0.7, 0.69, 0.7, 0.69, 0.69, 0.69, 0.69, 
    0.69, 0.69, 0.68, 0.7, 0.7, 0.7, 0.69, 0.69, 0.69, 0.69, 0.69, 0.7, 0.68, 
    0.67, 0.67, 0.68, 0.68, 0.69, 0.69, 0.68, 0.67, 0.68, 0.68, 0.67, 0.67, 
    0.67, 0.68, 0.71, 0.68, 0.68, 0.68, 0.67, 0.67, 0.68, 0.68, 0.69, 0.7, 
    0.7, 0.7, 0.71, 0.71, 0.71, 0.71, 0.7, 0.7, 0.7, 0.71, 0.64, 0.66, 0.72, 
    0.63, 0.75, 0.74, 0.67, 0.76, 0.78, 0.73, 0.74, 0.79, 0.78, 0.64, 0.78, 
    0.7, 0.71, 0.57, 0.75, 0.81, 0.61, 0.7, 0.83, 0.8, 0.79, 0.81, 0.75, 
    0.68, 0.67, 0.74, 0.63, 0.63, 0.59, 0.76, 0.6, 0.57, 0.72, 0.75, 0.73, 
    0.72, 0.7, 0.72, 0.57, 0.57, 0.66, 0.75, 0.64, 0.76, 0.71, 0.69, 0.71, 
    0.72, 0.72, 0.77, 0.78, 0.78, 0.78, 0.79, 0.79, 0.79, 0.73, 0.78, 0.83, 
    0.83, 0.81, 0.75, 0.8, 0.72, 0.81, 0.79, 0.78, 0.77, 0.79, 0.79, 0.76, 
    0.66, 0.71, 0.75, 0.73, 0.8, 0.8, 0.74, 0.78, 0.75, 0.77, 0.76, 0.78, 
    0.72, 0.74, 0.8, 0.78, 0.82, 0.77, 0.79, 0.79, 0.78, 0.79, 0.79, 0.8, 
    0.81, 0.73, 0.69, 0.72, 0.75, 0.78, 0.7, 0.69, 0.7, 0.67, 0.7, 0.7, 0.67, 
    0.67, 0.71, 0.8, 0.71, 0.7, 0.73, 0.71, 0.7, 0.7, 0.73, 0.74, 0.72, 0.79, 
    0.76, 0.71, 0.75, 0.78, 0.77, 0.78, 0.77, 0.79, 0.76, 0.71, 0.68, 0.76, 
    0.72, 0.76, 0.75, 0.77, 0.77, 0.77, 0.75, 0.74, 0.76, 0.77, 0.76, 0.74, 
    0.73, 0.74, 0.76, 0.77, 0.77, 0.78, 0.79, 0.8, 0.79, 0.81, 0.83, 0.81, 
    0.78, 0.83, 0.8, 0.82, 0.84, 0.85, 0.83, 0.81, 0.81, 0.81, 0.81, 0.85, 
    0.84, 0.85, 0.84, 0.83, 0.83, 0.83, 0.8, 0.81, 0.8, 0.81, 0.81, 0.81, 
    0.81, 0.81, 0.8, 0.81, 0.79, 0.81, 0.81, 0.81, 0.83, 0.81, 0.81, 0.81, 
    0.86, 0.8, 0.8, 0.82, 0.81, 0.83, 0.82, 0.79, 0.77, 0.77, 0.79, 0.81, 
    0.82, 0.81, 0.8, 0.81, 0.82, 0.83, 0.84, 0.85, 0.85, 0.85, 0.86, 0.87, 
    0.86, 0.84, 0.84, 0.86, 0.85, 0.86, 0.86, 0.85, 0.84, 0.84, 0.83, 0.83, 
    0.84, 0.85, 0.85, 0.84, 0.84, 0.81, 0.84, 0.82, 0.81, 0.82, 0.79, 0.82, 
    0.8, 0.81, 0.8, 0.82, 0.82, 0.78, 0.79, 0.76, 0.79, 0.78, 0.79, 0.8, 
    0.84, 0.84, 0.83, 0.79, 0.8, 0.78, 0.75, 0.79, 0.73, 0.75, 0.83, 0.78, 
    0.8, 0.84, 0.87, 0.89, 0.91, 0.88, 0.89, 0.86, 0.82, 0.84, 0.83, 0.84, 
    0.9, 0.82, 0.82, 0.8, 0.84, 0.78, 0.72, 0.64, 0.73, 0.75, 0.7, 0.62, 
    0.65, 0.56, 0.64, 0.52, 0.65, 0.65, 0.7, 0.76, 0.84, 0.84, 0.88, 0.89, 
    0.8, 0.81, 0.77, 0.85, 0.84, 0.86, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 
    0.83, 0.83, 0.83, 0.83, 0.85, 0.86, 0.88, 0.91, 0.91, 0.9, 0.9, 0.87, 
    0.86, 0.82, 0.8, 0.82, 0.87, 0.88, 0.88, 0.87, 0.85, 0.8, 0.76, 0.72, 
    0.8, 0.74, 0.69, 0.69, 0.69, 0.7, 0.74, 0.74, 0.78, 0.83, 0.85, 0.82, 
    0.83, 0.82, 0.82, 0.82, 0.81, 0.79, 0.82, 0.79, 0.79, 0.77, 0.77, 0.76, 
    0.79, 0.77, 0.78, 0.75, 0.75, 0.78, 0.78, 0.79, 0.82, 0.85, 0.87, 0.89, 
    0.9, 0.9, 0.89, 0.9, 0.92, 0.9, 0.9, 0.89, 0.9, 0.89, 0.89, 0.9, 0.84, 
    0.86, 0.88, 0.8, 0.85, 0.87, 0.88, 0.89, 0.86, 0.82, 0.81, 0.85, 0.89, 
    0.89, 0.92, 0.93, 0.92, 0.91, 0.89, 0.87, 0.93, 0.93, 0.92, 0.93, 0.92, 
    0.92, 0.9, 0.9, 0.92, 0.9, 0.92, 0.94, 0.95, 0.95, 0.95, 0.94, 0.93, 
    0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 0.97, 0.96, 0.95, 0.95, 
    0.95, 0.95, 0.94, 0.95, 0.96, 0.95, 0.97, 0.97, 0.97, 0.95, 0.96, 0.97, 
    0.96, 0.96, 0.94, 0.93, 0.94, 0.94, 0.94, 0.96, 0.96, 0.96, 0.93, 0.93, 
    0.97, 0.97, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.96, 0.92, 0.92, 
    0.89, 0.88, 0.89, 0.9, 0.87, 0.82, 0.76, 0.76, 0.81, 0.87, 0.89, 0.88, 
    0.72, 0.68, 0.76, 0.74, 0.79, 0.86, 0.89, 0.89, 0.88, 0.91, 0.85, 0.86, 
    0.89, 0.89, 0.81, 0.82, 0.89, 0.9, 0.9, 0.92, 0.93, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.91, 0.92, 0.92, 0.93, 0.89, 0.95, 0.96, 0.96, 0.94, 0.95, 
    0.95, 0.95, 0.9, 0.9, 0.88, 0.89, 0.85, 0.79, 0.89, 0.9, 0.9, 0.88, 0.9, 
    0.87, 0.85, 0.88, 0.86, 0.85, 0.85, 0.86, 0.87, 0.86, 0.86, 0.83, 0.84, 
    0.81, 0.82, 0.87, 0.89, 0.88, 0.89, 0.88, 0.83, 0.89, 0.84, 0.82, 0.87, 
    0.89, 0.9, 0.87, 0.85, 0.88, 0.87, 0.89, 0.85, 0.86, 0.84, 0.85, 0.82, 
    0.85, 0.87, 0.87, 0.88, 0.87, 0.84, 0.84, 0.84, 0.85, 0.86, 0.85, 0.86, 
    0.87, 0.84, 0.85, 0.84, 0.84, 0.86, 0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 
    0.85, 0.85, 0.84, 0.85, 0.85, 0.84, 0.83, 0.83, 0.84, 0.84, 0.84, 0.81, 
    0.82, 0.82, 0.81, 0.78, 0.77, 0.74, 0.74, 0.78, 0.78, 0.78, 0.77, 0.8, 
    0.8, 0.81, 0.76, 0.79, 0.78, 0.76, 0.74, 0.77, 0.8, 0.71, 0.77, 0.8, 
    0.77, 0.79, 0.82, 0.82, 0.83, 0.85, 0.85, 0.84, 0.83, 0.82, 0.8, 0.82, 
    0.8, 0.81, 0.82, 0.84, 0.84, 0.85, 0.84, 0.83, 0.82, 0.83, 0.83, 0.83, 
    0.78, 0.78, 0.75, 0.74, 0.8, 0.81, 0.81, 0.81, 0.8, 0.79, 0.82, 0.8, 0.8, 
    0.72, 0.79, 0.81, 0.84, 0.82, 0.81, 0.76, 0.61, 0.52, 0.57, 0.61, 0.66, 
    0.76, 0.85, 0.88, 0.88, 0.89, 0.88, 0.8, 0.85, 0.83, 0.81, 0.86, 0.8, 
    0.79, 0.8, 0.78, 0.78, 0.72, 0.72, 0.74, 0.73, 0.72, 0.73, 0.76, 0.78, 
    0.8, 0.83, 0.85, 0.86, 0.85, 0.84, 0.84, 0.83, 0.83, 0.82, 0.83, 0.84, 
    0.83, 0.83, 0.83, 0.82, 0.84, 0.8, 0.82, 0.78, 0.81, 0.8, 0.83, 0.81, 
    0.74, 0.69, 0.7, 0.74, 0.74, 0.71, 0.7, 0.7, 0.69, 0.72, 0.78, 0.82, 
    0.78, 0.77, 0.8, 0.72, 0.82, 0.79, 0.75, 0.8, 0.8, 0.79, 0.76, 0.78, 
    0.79, 0.8, 0.84, 0.83, 0.83, 0.83, 0.8, 0.78, 0.77, 0.77, 0.77, 0.75, 
    0.76, 0.76, 0.79, 0.81, 0.76, 0.73, 0.75, 0.8, 0.72, 0.72, 0.67, 0.65, 
    0.63, 0.6, 0.64, 0.63, 0.65, 0.68, 0.69, 0.71, 0.73, 0.74, 0.74, 0.77, 
    0.8, 0.8, 0.81, 0.82, 0.84, 0.85, 0.86, 0.86, 0.87, 0.87, 0.88, 0.83, 
    0.79, 0.79, 0.76, 0.76, 0.79, 0.79, 0.79, 0.82, 0.82, 0.82, 0.77, 0.8, 
    0.78, 0.83, 0.85, 0.86, 0.87, 0.88, 0.88, 0.88, 0.9, 0.91, 0.93, 0.93, 
    0.94, 0.93, 0.94, 0.92, 0.89, 0.89, 0.9, 0.89, 0.9, 0.89, 0.87, 0.87, 
    0.87, 0.88, 0.89, 0.9, 0.95, 0.96, 0.94, 0.93, 0.94, 0.94, 0.94, 0.92, 
    0.91, 0.91, 0.92, 0.91, 0.92, 0.92, 0.91, 0.89, 0.9, 0.88, 0.85, 0.84, 
    0.86, 0.81, 0.84, 0.8, 0.85, 0.84, 0.83, 0.77, 0.79, 0.78, 0.84, 0.86, 
    0.84, 0.85, 0.83, 0.86, 0.83, 0.83, 0.83, 0.82, 0.84, 0.85, 0.85, 0.85, 
    0.87, 0.86, 0.87, 0.85, 0.85, 0.78, 0.8, 0.8, 0.81, 0.79, 0.84, 0.83, 
    0.82, 0.81, 0.81, 0.79, 0.77, 0.77, 0.77, 0.77, 0.76, 0.76, 0.75, 0.74, 
    0.71, 0.74, 0.72, 0.74, 0.74, 0.74, 0.74, 0.77, 0.69, 0.71, 0.78, 0.75, 
    0.76, 0.73, 0.72, 0.74, 0.72, 0.76, 0.74, 0.69, 0.79, 0.78, 0.82, 0.79, 
    0.74, 0.75, 0.74, 0.77, 0.77, 0.81, 0.81, 0.8, 0.8, 0.79, 0.81, 0.81, 
    0.8, 0.8, 0.81, 0.79, 0.8, 0.79, 0.82, 0.82, 0.82, 0.78, 0.78, 0.71, 
    0.69, 0.75, 0.78, 0.8, 0.81, 0.81, 0.81, 0.85, 0.85, 0.85, 0.86, 0.84, 
    0.83, 0.78, 0.8, 0.81, 0.81, 0.8, 0.78, 0.77, 0.71, 0.67, 0.7, 0.75, 
    0.79, 0.82, 0.81, 0.8, 0.8, 0.8, 0.8, 0.79, 0.77, 0.77, 0.77, 0.79, 0.81, 
    0.82, 0.83, 0.83, 0.83, 0.84, 0.84, 0.85, 0.86, 0.86, 0.85, 0.85, 0.85, 
    0.85, 0.85, 0.85, 0.86, 0.87, 0.87, 0.87, 0.88, 0.89, 0.89, 0.9, 0.91, 
    0.91, 0.91, 0.9, 0.91, 0.9, 0.9, 0.89, 0.88, 0.89, 0.89, 0.9, 0.91, 0.92, 
    0.93, 0.93, 0.94, 0.94, 0.95, 0.96, 0.97, 0.96, 0.96, 0.95, 0.95, 0.96, 
    0.95, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.94, 0.95, 0.94, 
    0.93, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.95, 0.93, 0.94, 0.92, 
    0.88, 0.91, 0.94, 0.87, 0.84, 0.83, 0.88, 0.87, 0.85, 0.85, 0.84, 0.85, 
    0.84, 0.84, 0.85, 0.82, 0.83, 0.87, 0.85, 0.83, 0.85, 0.83, 0.78, 0.77, 
    0.79, 0.82, 0.77, 0.83, 0.87, 0.82, 0.8, 0.77, 0.83, 0.86, 0.85, 0.77, 
    0.73, 0.72, 0.68, 0.84, 0.83, 0.79, 0.81, 0.83, 0.82, 0.79, 0.78, 0.76, 
    0.77, 0.78, 0.73, 0.74, 0.74, 0.73, 0.72, 0.72, 0.73, 0.7, 0.69, 0.67, 
    0.65, 0.69, 0.77, 0.8, 0.77, 0.82, 0.82, 0.85, 0.81, 0.79, 0.79, 0.82, 
    0.85, 0.9, 0.92, 0.92, 0.92, 0.91, 0.91, 0.92, 0.9, 0.89, 0.81, 0.84, 
    0.83, 0.87, 0.88, 0.9, 0.9, 0.87, 0.87, 0.87, 0.88, 0.79, 0.85, 0.96, 
    0.95, 0.94, 0.93, 0.93, 0.94, 0.94, 0.94, 0.88, 0.89, 0.91, 0.91, 0.88, 
    0.87, 0.89, 0.91, 0.91, 0.9, 0.91, 0.92, 0.93, 0.93, 0.94, 0.95, 0.94, 
    0.93, 0.92, 0.91, 0.89, 0.9, 0.9, 0.92, 0.91, 0.93, 0.91, 0.91, 0.9, 
    0.93, 0.9, 0.87, 0.89, 0.89, 0.88, 0.91, 0.91, 0.91, 0.93, 0.96, 0.96, 
    0.96, 0.97, 0.94, 0.82, 0.79, 0.8, 0.86, 0.86, 0.87, 0.87, 0.88, 0.89, 
    0.89, 0.88, 0.93, 0.87, 0.81, 0.77, 0.82, 0.79, 0.76, 0.79, 0.78, 0.81, 
    0.81, 0.82, 0.8, 0.77, 0.83, 0.8, 0.76, 0.74, 0.74, 0.79, 0.78, 0.8, 
    0.83, 0.88, 0.91, 0.93, 0.93, 0.93, 0.91, 0.91, 0.9, 0.92, 0.92, 0.92, 
    0.93, 0.91, 0.89, 0.89, 0.88, 0.9, 0.88, 0.9, 0.92, 0.94, 0.93, 0.93, 
    0.94, 0.92, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 0.92, 0.91, 0.91, 
    0.89, 0.89, 0.89, 0.89, 0.85, 0.84, 0.91, 0.94, 0.92, 0.88, 0.91, 0.9, 
    0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 0.84, 0.84, 0.85, 0.85, 0.87, 0.87, 
    0.87, 0.87, 0.89, 0.89, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 
    0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 
    0.98, 0.98, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.98, 0.99, 0.98, 0.97, 0.96, 0.93, 0.91, 0.89, 0.88, 0.88, 
    0.9, 0.9, 0.91, 0.92, 0.93, 0.91, 0.89, 0.88, 0.9, 0.9, 0.95, 0.92, 0.92, 
    0.87, 0.86, 0.82, 0.86, 0.86, 0.86, 0.89, 0.87, 0.89, 0.91, 0.9, 0.88, 
    0.88, 0.87, 0.87, 0.87, 0.87, 0.87, 0.89, 0.89, 0.91, 0.9, 0.9, 0.91, 
    0.9, 0.91, 0.89, 0.89, 0.89, 0.88, 0.88, 0.88, 0.87, 0.87, 0.87, 0.86, 
    0.86, 0.86, 0.86, 0.85, 0.86, 0.86, 0.87, 0.9, 0.92, 0.92, 0.92, 0.91, 
    0.92, 0.95, 0.97, 0.97, 0.96, 0.95, 0.9, 0.85, 0.85, 0.81, 0.81, 0.8, 
    0.85, 0.86, 0.87, 0.87, 0.89, 0.87, 0.85, 0.86, 0.85, 0.87, 0.86, 0.89, 
    0.9, 0.91, 0.91, 0.86, 0.84, 0.88, 0.9, 0.91, 0.91, 0.91, 0.92, 0.93, 
    0.93, 0.94, 0.93, 0.94, 0.94, 0.94, 0.95, 0.96, 0.96, 0.95, 0.93, 0.94, 
    0.78, 0.78, 0.76, 0.73, 0.72, 0.73, 0.76, 0.84, 0.89, 0.84, 0.77, 0.73, 
    0.76, 0.81, 0.78, 0.74, 0.71, 0.78, 0.82, 0.84, 0.86, 0.86, 0.86, 0.87, 
    0.89, 0.9, 0.9, 0.9, 0.87, 0.85, 0.86, 0.87, 0.86, 0.85, 0.86, 0.87, 
    0.86, 0.89, 0.91, 0.9, 0.92, 0.92, 0.9, 0.92, 0.88, 0.89, 0.89, 0.89, 
    0.89, 0.93, 0.94, 0.96, 0.95, 0.93, 0.97, 0.96, 0.95, 0.94, 0.94, 0.93, 
    0.89, 0.89, 0.94, 0.94, 0.96, 0.93, 0.91, 0.87, 0.87, 0.86, 0.86, 0.85, 
    0.85, 0.85, 0.86, 0.86, 0.86, 0.84, 0.84, 0.85, 0.86, 0.82, 0.82, 0.86, 
    0.85, 0.85, 0.86, 0.87, 0.89, 0.9, 0.89, 0.87, 0.87, 0.85, 0.89, 0.88, 
    0.84, 0.91, 0.92, 0.94, 0.96, 0.95, 0.95, 0.95, 0.91, 0.91, 0.84, 0.83, 
    0.82, 0.88, 0.94, 0.86, 0.79, 0.8, 0.88, 0.84, 0.9, 0.88, 0.88, 0.9, 
    0.88, 0.91, 0.9, 0.9, 0.87, 0.88, 0.91, 0.93, 0.9, 0.91, 0.9, 0.89, 0.92, 
    0.91, 0.91, 0.91, 0.89, 0.9, 0.9, 0.9, 0.89, 0.89, 0.89, 0.88, 0.88, 
    0.89, 0.91, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 0.95, 
    0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.98, 0.97, 
    0.97, 0.97, 0.96, 0.95, 0.94, 0.96, 0.96, 0.96, 0.98, 0.98, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.97, 0.92, 0.9, 0.89, 0.9, 0.91, 0.89, 0.86, 0.88, 
    0.86, 0.87, 0.85, 0.82, 0.82, 0.84, 0.9, 0.89, 0.89, 0.9, 0.88, 0.89, 
    0.92, 0.94, 0.95, 0.96, 0.94, 0.93, 0.91, 0.9, 0.9, 0.92, 0.92, 0.91, 
    0.93, 0.93, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 
    0.92, 0.93, 0.92, 0.92, 0.96, 0.96, 0.92, 0.93, 0.93, 0.92, 0.9, 0.84, 
    0.87, 0.82, 0.86, 0.84, 0.88, 0.9, 0.94, 0.94, 0.94, 0.91, 0.91, 0.9, 
    0.9, 0.93, 0.93, 0.94, 0.94, 0.92, 0.92, 0.87, 0.85, 0.88, 0.9, 0.91, 
    0.92, 0.91, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.91, 0.91, 
    0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 0.95, 
    0.92, 0.92, 0.93, 0.94, 0.93, 0.94, 0.94, 0.93, 0.92, 0.93, 0.92, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.95, 0.95, 0.97, 0.96, 0.96, 0.96, 0.96, 0.95, 
    0.95, 0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.95, 
    0.94, 0.95, 0.94, 0.94, 0.94, 0.94, 0.95, 0.96, 0.97, 0.99, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.97, 0.99, 0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.96, 0.92, 0.94, 0.9, 
    0.93, 0.96, 0.97, 0.98, 0.94, 0.94, 0.93, 0.89, 0.89, 0.89, 0.93, 0.89, 
    0.87, 0.9, 0.89, 0.82, 0.8, 0.76, 0.81, 0.79, 0.86, 0.77, 0.9, 0.89, 
    0.81, 0.8, 0.86, 0.81, 0.84, 0.79, 0.89, 0.91, 0.91, 0.85, 0.91, 0.91, 
    0.91, 0.92, 0.92, 0.9, 0.87, 0.9, 0.89, 0.85, 0.88, 0.88, 0.85, 0.86, 
    0.87, 0.9, 0.9, 0.92, 0.91, 0.9, 0.92, 0.91, 0.89, 0.9, 0.91, 0.91, 0.9, 
    0.89, 0.9, 0.92, 0.92, 0.92, 0.95, 0.95, 0.95, 0.93, 0.93, 0.92, 0.92, 
    0.92, 0.92, 0.91, 0.93, 0.93, 0.93, 0.92, 0.89, 0.93, 0.94, 0.93, 0.93, 
    0.94, 0.95, 0.93, 0.95, 0.94, 0.96, 0.95, 0.94, 0.94, 0.94, 0.93, 0.94, 
    0.94, 0.96, 0.96, 0.98, 0.98, 0.96, 0.91, 0.93, 0.96, 0.97, 0.97, 0.97, 
    0.97, 0.96, 0.93, 0.91, 0.9, 0.91, 0.91, 0.9, 0.88, 0.86, 0.86, 0.83, 
    0.86, 0.86, 0.89, 0.9, 0.88, 0.9, 0.88, 0.9, 0.87, 0.84, 0.81, 0.77, 
    0.82, 0.79, 0.85, 0.85, 0.82, 0.82, 0.8, 0.77, 0.77, 0.68, 0.71, 0.7, 
    0.72, 0.74, 0.66, 0.74, 0.75, 0.66, 0.71, 0.82, 0.92, 0.93, 0.81, 0.74, 
    0.72, 0.73, 0.7, 0.66, 0.69, 0.79, 0.81, 0.85, 0.84, 0.9, 0.67, 0.74, 
    0.83, 0.81, 0.7, 0.76, 0.79, 0.81, 0.82, 0.83, 0.89, 0.82, 0.83, 0.82, 
    0.81, 0.84, 0.84, 0.84, 0.8, 0.81, 0.83, 0.86, 0.85, 0.86, 0.84, 0.83, 
    0.79, 0.8, 0.85, 0.83, 0.82, 0.87, 0.88, 0.86, 0.85, 0.86, 0.89, 0.89, 
    0.9, 0.76, 0.75, 0.76, 0.77, 0.84, 0.78, 0.81, 0.77, 0.83, 0.86, 0.84, 
    0.86, 0.89, 0.91, 0.94, 0.93, 0.91, 0.88, 0.85, 0.87, 0.86, 0.87, 0.83, 
    0.87, 0.9, 0.9, 0.92, 0.92, 0.92, 0.91, 0.89, 0.87, 0.93, 0.92, 0.89, 
    0.89, 0.89, 0.87, 0.85, 0.87, 0.85, 0.9, 0.92, 0.96, 0.93, 0.96, 0.93, 
    0.88, 0.87, 0.87, 0.85, 0.87, 0.88, 0.89, 0.87, 0.9, 0.88, 0.82, 0.87, 
    0.85, 0.86, 0.86, 0.87, 0.88, 0.89, 0.87, 0.89, 0.88, 0.84, 0.86, 0.86, 
    0.85, 0.84, 0.84, 0.86, 0.88, 0.88, 0.88, 0.86, 0.91, 0.92, 0.9, 0.87, 
    0.86, 0.85, 0.85, 0.84, 0.86, 0.87, 0.9, 0.91, 0.92, 0.93, 0.91, 0.91, 
    0.9, 0.89, 0.86, 0.86, 0.89, 0.91, 0.88, 0.9, 0.91, 0.91, 0.88, 0.86, 
    0.86, 0.85, 0.85, 0.85, 0.84, 0.86, 0.86, 0.87, 0.92, 0.93, 0.93, 0.93, 
    0.94, 0.94, 0.94, 0.93, 0.91, 0.91, 0.92, 0.92, 0.91, 0.9, 0.88, 0.89, 
    0.88, 0.88, 0.88, 0.88, 0.88, 0.87, 0.87, 0.87, 0.88, 0.88, 0.88, 0.87, 
    0.88, 0.87, 0.87, 0.87, 0.89, 0.91, 0.91, 0.91, 0.84, 0.85, 0.84, 0.86, 
    0.89, 0.88, 0.88, 0.85, 0.86, 0.85, 0.84, 0.82, 0.83, 0.82, 0.82, 0.81, 
    0.8, 0.79, 0.8, 0.8, 0.79, 0.78, 0.8, 0.79, 0.79, 0.78, 0.78, 0.78, 0.78, 
    0.8, 0.75, 0.74, 0.77, 0.77, 0.75, 0.75, 0.76, 0.75, 0.73, 0.76, 0.7, 
    0.74, 0.76, 0.75, 0.74, 0.74, 0.77, 0.84, 0.84, 0.83, 0.82, 0.74, 0.73, 
    0.73, 0.75, 0.74, 0.77, 0.77, 0.77, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 
    0.77, 0.79, 0.76, 0.72, 0.77, 0.78, 0.78, 0.79, 0.8, 0.82, 0.81, 0.82, 
    0.82, 0.82, 0.81, 0.83, 0.81, 0.83, 0.82, 0.81, 0.84, 0.88, 0.88, 0.9, 
    0.9, 0.89, 0.88, 0.93, 0.92, 0.94, 0.91, 0.93, 0.94, 0.95, 0.89, 0.9, 
    0.9, 0.91, 0.95, 0.94, 0.92, 0.91, 0.89, 0.88, 0.87, 0.86, 0.86, 0.86, 
    0.84, 0.84, 0.85, 0.83, 0.83, 0.84, 0.82, 0.81, 0.81, 0.81, 0.83, 0.83, 
    0.81, 0.78, 0.81, 0.82, 0.83, 0.83, 0.85, 0.78, 0.8, 0.79, 0.78, 0.78, 
    0.76, 0.75, 0.81, 0.86, 0.92, 0.94, 0.95, 0.92, 0.88, 0.83, 0.87, 0.83, 
    0.88, 0.89, 0.88, 0.85, 0.86, 0.86, 0.88, 0.87, 0.88, 0.9, 0.92, 0.89, 
    0.85, 0.86, 0.94, 0.93, 0.92, 0.93, 0.93, 0.95, 0.92, 0.9, 0.91, 0.9, 
    0.92, 0.93, 0.94, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.97, 0.96, 
    0.95, 0.95, 0.95, 0.94, 0.94, 0.93, 0.94, 0.94, 0.94, 0.94, 0.93, 0.94, 
    0.94, 0.94, 0.93, 0.94, 0.94, 0.95, 0.95, 0.97, 0.96, 0.95, 0.96, 0.97, 
    0.98, 0.99, 0.98, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.96, 0.95, 
    0.94, 0.93, 0.91, 0.91, 0.88, 0.86, 0.84, 0.82, 0.81, 0.8, 0.81, 0.86, 
    0.88, 0.87, 0.87, 0.84, 0.82, 0.82, 0.81, 0.8, 0.81, 0.79, 0.86, 0.78, 
    0.82, 0.81, 0.79, 0.78, 0.76, 0.75, 0.77, 0.78, 0.82, 0.76, 0.76, 0.79, 
    0.81, 0.8, 0.79, 0.79, 0.77, 0.77, 0.78, 0.8, 0.81, 0.8, 0.77, 0.8, 0.83, 
    0.8, 0.78, 0.75, 0.81, 0.79, 0.75, 0.83, 0.83, 0.76, 0.77, 0.79, 0.8, 
    0.86, 0.8, 0.78, 0.8, 0.83, 0.81, 0.81, 0.81, 0.82, 0.8, 0.8, 0.81, 0.82, 
    0.83, 0.83, 0.81, 0.84, 0.83, 0.83, 0.83, 0.83, 0.84, 0.8, 0.79, 0.81, 
    0.8, 0.81, 0.82, 0.79, 0.82, 0.8, 0.81, 0.8, 0.83, 0.83, 0.84, 0.83, 
    0.83, 0.82, 0.82, 0.83, 0.82, 0.82, 0.81, 0.79, 0.83, 0.82, 0.83, 0.83, 
    0.81, 0.7, 0.59, 0.59, 0.64, 0.69, 0.74, 0.75, 0.68, 0.7, 0.71, 0.73, 
    0.74, 0.7, 0.68, 0.69, 0.73, 0.78, 0.79, 0.79, 0.81, 0.82, 0.85, 0.87, 
    0.75, 0.76, 0.76, 0.83, 0.81, 0.81, 0.8, 0.79, 0.78, 0.8, 0.78, 0.79, 
    0.81, 0.82, 0.82, 0.82, 0.82, 0.81, 0.81, 0.81, 0.81, 0.8, 0.8, 0.81, 
    0.8, 0.79, 0.8, 0.78, 0.79, 0.77, 0.77, 0.78, 0.79, 0.81, 0.82, 0.82, 
    0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 
    0.82, 0.82, 0.82, 0.82, 0.81, 0.81, 0.8, 0.79, 0.8, 0.8, 0.79, 0.79, 
    0.79, 0.77, 0.79, 0.8, 0.8, 0.81, 0.8, 0.8, 0.82, 0.82, 0.84, 0.82, 0.81, 
    0.8, 0.79, 0.79, 0.8, 0.83, 0.74, 0.75, 0.77, 0.79, 0.74, 0.78, 0.82, 
    0.84, 0.8, 0.82, 0.84, 0.83, 0.83, 0.83, 0.84, 0.84, 0.83, 0.85, 0.86, 
    0.85, 0.84, 0.85, 0.86, 0.85, 0.86, 0.86, 0.85, 0.86, 0.86, 0.87, 0.86, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.85, 0.85, 0.83, 0.84, 0.85, 
    0.85, 0.84, 0.85, 0.85, 0.85, 0.86, 0.85, 0.86, 0.85, 0.82, 0.83, 0.84, 
    0.83, 0.85, 0.85, 0.84, 0.84, 0.84, 0.83, 0.84, 0.83, 0.82, 0.81, 0.81, 
    0.81, 0.78, 0.78, 0.8, 0.81, 0.82, 0.83, 0.84, 0.84, 0.83, 0.83, 0.8, 
    0.83, 0.87, 0.85, 0.83, 0.82, 0.78, 0.81, 0.86, 0.86, 0.83, 0.82, 0.77, 
    0.76, 0.78, 0.75, 0.79, 0.79, 0.81, 0.78, 0.76, 0.81, 0.82, 0.84, 0.82, 
    0.8, 0.83, 0.81, 0.83, 0.82, 0.81, 0.82, 0.81, 0.85, 0.82, 0.82, 0.8, 
    0.79, 0.8, 0.77, 0.81, 0.79, 0.79, 0.83, 0.82, 0.84, 0.82, 0.82, 0.83, 
    0.85, 0.84, 0.81, 0.78, 0.8, 0.81, 0.8, 0.78, 0.77, 0.79, 0.8, 0.8, 0.8, 
    0.79, 0.78, 0.76, 0.76, 0.78, 0.78, 0.8, 0.81, 0.83, 0.85, 0.82, 0.82, 
    0.81, 0.8, 0.8, 0.81, 0.81, 0.83, 0.83, 0.85, 0.84, 0.84, 0.84, 0.83, 
    0.85, 0.85, 0.84, 0.86, 0.86, 0.87, 0.88, 0.87, 0.87, 0.86, 0.86, 0.84, 
    0.84, 0.87, 0.85, 0.85, 0.86, 0.82, 0.83, 0.86, 0.82, 0.82, 0.86, 0.83, 
    0.83, 0.81, 0.81, 0.8, 0.77, 0.78, 0.81, 0.81, 0.83, 0.83, 0.84, 0.84, 
    0.84, 0.82, 0.83, 0.85, 0.83, 0.84, 0.84, 0.85, 0.85, 0.85, 0.84, 0.82, 
    0.84, 0.84, 0.84, 0.84, 0.83, 0.85, 0.86, 0.86, 0.84, 0.84, 0.87, 0.86, 
    0.86, 0.85, 0.85, 0.86, 0.86, 0.87, 0.87, 0.88, 0.88, 0.79, 0.77, 0.77, 
    0.76, 0.78, 0.81, 0.81, 0.81, 0.81, 0.8, 0.84, 0.87, 0.85, 0.88, 0.9, 
    0.9, 0.91, 0.92, 0.92, 0.93, 0.94, 0.95, 0.95, 0.96, 0.94, 0.94, 0.93, 
    0.91, 0.82, 0.88, 0.85, 0.86, 0.81, 0.83, 0.89, 0.88, 0.87, 0.86, 0.87, 
    0.89, 0.9, 0.91, 0.89, 0.86, 0.86, 0.85, 0.84, 0.83, 0.82, 0.83, 0.84, 
    0.83, 0.83, 0.82, 0.79, 0.81, 0.83, 0.83, 0.81, 0.82, 0.82, 0.8, 0.8, 
    0.82, 0.82, 0.82, 0.83, 0.82, 0.83, 0.84, 0.82, 0.81, 0.79, 0.77, 0.78, 
    0.79, 0.79, 0.77, 0.7, 0.75, 0.82, 0.81, 0.79, 0.78, 0.76, 0.78, 0.76, 
    0.77, 0.75, 0.75, 0.76, 0.76, 0.76, 0.77, 0.75, 0.72, 0.75, 0.74, 0.73, 
    0.72, 0.7, 0.7, 0.7, 0.7, 0.72, 0.77, 0.78, 0.79, 0.8, 0.78, 0.81, 0.81, 
    0.79, 0.8, 0.8, 0.74, 0.75, 0.75, 0.74, 0.74, 0.75, 0.77, 0.79, 0.81, 
    0.81, 0.79, 0.79, 0.81, 0.79, 0.78, 0.8, 0.83, 0.79, 0.78, 0.77, 0.73, 
    0.74, 0.77, 0.78, 0.77, 0.76, 0.78, 0.77, 0.77, 0.77, 0.79, 0.78, 0.78, 
    0.78, 0.78, 0.78, 0.78, 0.78, 0.77, 0.79, 0.79, 0.81, 0.81, 0.82, 0.82, 
    0.82, 0.82, 0.82, 0.83, 0.83, 0.83, 0.81, 0.81, 0.77, 0.79, 0.79, 0.77, 
    0.78, 0.82, 0.84, 0.81, 0.78, 0.81, 0.78, 0.76, 0.81, 0.79, 0.78, 0.81, 
    0.81, 0.78, 0.77, 0.8, 0.78, 0.78, 0.76, 0.77, 0.78, 0.78, 0.76, 0.72, 
    0.72, 0.71, 0.74, 0.77, 0.73, 0.78, 0.81, 0.84, 0.83, 0.81, 0.8, 0.76, 
    0.83, 0.84, 0.82, 0.8, 0.74, 0.77, 0.79, 0.77, 0.78, 0.8, 0.79, 0.78, 
    0.76, 0.79, 0.77, 0.75, 0.82, 0.83, 0.82, 0.83, 0.81, 0.81, 0.82, 0.82, 
    0.84, 0.84, 0.83, 0.85, 0.84, 0.83, 0.83, 0.82, 0.81, 0.82, 0.82, 0.81, 
    0.81, 0.81, 0.8, 0.81, 0.81, 0.81, 0.81, 0.8, 0.81, 0.81, 0.78, 0.77, 
    0.78, 0.79, 0.78, 0.8, 0.8, 0.79, 0.78, 0.79, 0.8, 0.78, 0.79, 0.79, 
    0.79, 0.77, 0.78, 0.8, 0.8, 0.8, 0.81, 0.81, 0.78, 0.79, 0.8, 0.8, 0.79, 
    0.79, 0.79, 0.79, 0.79, 0.78, 0.75, 0.76, 0.79, 0.76, 0.71, 0.64, 0.67, 
    0.69, 0.76, 0.79, 0.84, 0.85, 0.83, 0.82, 0.84, 0.85, 0.88, 0.87, 0.88, 
    0.89, 0.88, 0.88, 0.89, 0.89, 0.88, 0.9, 0.89, 0.89, 0.85, 0.86, 0.82, 
    0.83, 0.83, 0.84, 0.84, 0.85, 0.86, 0.81, 0.82, 0.8, 0.82, 0.84, 0.82, 
    0.83, 0.84, 0.85, 0.86, 0.82, 0.84, 0.83, 0.82, 0.83, 0.81, 0.82, 0.82, 
    0.81, 0.84, 0.87, 0.84, 0.85, 0.81, 0.79, 0.77, 0.8, 0.79, 0.77, 0.76, 
    0.77, 0.75, 0.77, 0.75, 0.76, 0.77, 0.77, 0.72, 0.68, 0.74, 0.71, 0.73, 
    0.73, 0.7, 0.7, 0.74, 0.74, 0.68, 0.77, 0.81, 0.7, 0.7, 0.77, 0.78, 0.78, 
    0.83, 0.78, 0.78, 0.79, 0.78, 0.77, 0.77, 0.77, 0.78, 0.76, 0.75, 0.76, 
    0.77, 0.76, 0.76, 0.78, 0.79, 0.79, 0.79, 0.79, 0.8, 0.8, 0.79, 0.79, 
    0.8, 0.78, 0.8, 0.79, 0.79, 0.78, 0.76, 0.74, 0.73, 0.75, 0.75, 0.74, 
    0.73, 0.73, 0.68, 0.68, 0.71, 0.69, 0.67, 0.72, 0.73, 0.79, 0.78, 0.8, 
    0.82, 0.81, 0.81, 0.75, 0.76, 0.75, 0.76, 0.76, 0.77, 0.75, 0.71, 0.69, 
    0.67, 0.75, 0.78, 0.81, 0.8, 0.8, 0.78, 0.78, 0.76, 0.78, 0.79, 0.79, 
    0.81, 0.79, 0.82, 0.81, 0.82, 0.82, 0.84, 0.8, 0.77, 0.77, 0.75, 0.72, 
    0.73, 0.76, 0.76, 0.72, 0.77, 0.74, 0.79, 0.82, 0.85, 0.87, 0.88, 0.88, 
    0.89, 0.93, 0.9, 0.84, 0.78, 0.87, 0.85, 0.87, 0.86, 0.84, 0.82, 0.86, 
    0.86, 0.7, 0.81, 0.86, 0.89, 0.9, 0.92, 0.94, 0.95, 0.96, 0.96, 0.96, 
    0.95, 0.95, 0.94, 0.93, 0.92, 0.92, 0.91, 0.9, 0.9, 0.92, 0.94, 0.91, 
    0.95, 0.97, 0.98, 0.98, 0.93, 0.9, 0.89, 0.86, 0.86, 0.86, 0.85, 0.85, 
    0.83, 0.83, 0.82, 0.82, 0.81, 0.8, 0.79, 0.79, 0.78, 0.76, 0.74, 0.76, 
    0.78, 0.75, 0.78, 0.76, 0.77, 0.76, 0.79, 0.77, 0.79, 0.79, 0.78, 0.8, 
    0.82, 0.81, 0.84, 0.82, 0.75, 0.77, 0.73, 0.75, 0.74, 0.73, 0.7, 0.74, 
    0.73, 0.74, 0.74, 0.77, 0.76, 0.81, 0.82, 0.8, 0.8, 0.79, 0.84, 0.84, 
    0.79, 0.75, 0.73, 0.75, 0.78, 0.79, 0.8, 0.79, 0.79, 0.78, 0.79, 0.77, 
    0.76, 0.77, 0.75, 0.76, 0.75, 0.76, 0.76, 0.74, 0.74, 0.76, 0.77, 0.79, 
    0.8, 0.75, 0.74, 0.75, 0.78, 0.77, 0.8, 0.69, 0.67, 0.71, 0.71, 0.7, 
    0.72, 0.71, 0.73, 0.81, 0.81, 0.8, 0.81, 0.82, 0.83, 0.82, 0.79, 0.81, 
    0.82, 0.82, 0.81, 0.81, 0.8, 0.8, 0.82, 0.76, 0.76, 0.76, 0.77, 0.75, 
    0.74, 0.77, 0.74, 0.8, 0.8, 0.8, 0.79, 0.79, 0.81, 0.8, 0.8, 0.81, 0.82, 
    0.82, 0.82, 0.82, 0.81, 0.81, 0.82, 0.81, 0.81, 0.8, 0.79, 0.8, 0.78, 
    0.79, 0.81, 0.81, 0.84, 0.83, 0.85, 0.85, 0.86, 0.86, 0.85, 0.86, 0.86, 
    0.84, 0.83, 0.83, 0.82, 0.8, 0.81, 0.79, 0.74, 0.73, 0.76, 0.79, 0.79, 
    0.81, 0.83, 0.83, 0.83, 0.84, 0.85, 0.84, 0.86, 0.85, 0.84, 0.84, 0.83, 
    0.83, 0.83, 0.83, 0.83, 0.82, 0.82, 0.82, 0.83, 0.84, 0.83, 0.78, 0.81, 
    0.81, 0.81, 0.8, 0.83, 0.83, 0.83, 0.83, 0.84, 0.85, 0.85, 0.86, 0.85, 
    0.85, 0.84, 0.83, 0.83, 0.85, 0.84, 0.84, 0.8, 0.81, 0.81, 0.8, 0.8, 
    0.81, 0.81, 0.79, 0.79, 0.82, 0.82, 0.82, 0.83, 0.84, 0.85, 0.83, 0.85, 
    0.82, 0.84, 0.82, 0.85, 0.84, 0.84, 0.84, 0.84, 0.8, 0.83, 0.82, 0.81, 
    0.77, 0.71, 0.67, 0.67, 0.64, 0.68, 0.78, 0.77, 0.75, 0.8, 0.79, 0.8, 
    0.79, 0.78, 0.76, 0.74, 0.73, 0.76, 0.71, 0.7, 0.69, 0.73, 0.74, 0.77, 
    0.77, 0.78, 0.8, 0.83, 0.85, 0.86, 0.86, 0.83, 0.86, 0.85, 0.85, 0.86, 
    0.85, 0.87, 0.85, 0.85, 0.85, 0.84, 0.83, 0.83, 0.83, 0.84, 0.84, 0.86, 
    0.83, 0.82, 0.82, 0.85, 0.82, 0.82, 0.84, 0.84, 0.86, 0.86, 0.87, 0.84, 
    0.84, 0.83, 0.83, 0.82, 0.83, 0.83, 0.82, 0.82, 0.82, 0.81, 0.77, 0.75, 
    0.79, 0.8, 0.79, 0.78, 0.79, 0.78, 0.79, 0.79, 0.81, 0.79, 0.77, 0.74, 
    0.73, 0.72, 0.76, 0.77, 0.78, 0.78, 0.76, 0.76, 0.74, 0.76, 0.77, 0.77, 
    0.75, 0.73, 0.71, 0.75, 0.76, 0.78, 0.78, 0.75, 0.77, 0.8, 0.79, 0.77, 
    0.81, 0.78, 0.77, 0.76, 0.75, 0.74, 0.72, 0.74, 0.72, 0.73, 0.75, 0.76, 
    0.76, 0.73, 0.75, 0.76, 0.78, 0.79, 0.81, 0.83, 0.83, 0.85, 0.85, 0.85, 
    0.83, 0.83, 0.84, 0.83, 0.84, 0.82, 0.81, 0.82, 0.82, 0.82, 0.82, 0.83, 
    0.83, 0.82, 0.83, 0.85, 0.86, 0.85, 0.87, 0.86, 0.87, 0.86, 0.86, 0.86, 
    0.86, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.82, 0.83, 0.83, 0.83, 0.82, 
    0.82, 0.82, 0.82, 0.84, 0.85, 0.84, 0.86, 0.86, 0.87, 0.87, 0.88, 0.87, 
    0.87, 0.86, 0.85, 0.83, 0.77, 0.8, 0.82, 0.77, 0.72, 0.74, 0.77, 0.75, 
    0.75, 0.78, 0.79, 0.81, 0.79, 0.79, 0.8, 0.8, 0.82, 0.85, 0.88, 0.87, 
    0.84, 0.84, 0.84, 0.84, 0.81, 0.81, 0.8, 0.81, 0.78, 0.79, 0.82, 0.82, 
    0.84, 0.86, 0.85, 0.84, 0.88, 0.82, 0.88, 0.88, 0.83, 0.85, 0.85, 0.87, 
    0.86, 0.88, 0.81, 0.79, 0.86, 0.78, 0.77, 0.75, 0.75, 0.83, 0.87, 0.84, 
    0.83, 0.84, 0.85, 0.87, 0.88, 0.87, 0.86, 0.89, 0.9, 0.91, 0.92, 0.9, 
    0.9, 0.92, 0.95, 0.71, 0.68, 0.68, 0.71, 0.75, 0.77, 0.75, 0.76, 0.78, 
    0.78, 0.79, 0.78, 0.76, 0.77, 0.8, 0.81, 0.84, 0.84, 0.82, 0.83, 0.81, 
    0.79, 0.84, 0.84, 0.8, 0.75, 0.71, 0.71, 0.7, 0.67, 0.64, 0.62, 0.58, 
    0.62, 0.66, 0.67, 0.68, 0.69, 0.73, 0.74, 0.78, 0.78, 0.77, 0.76, 0.77, 
    0.77, 0.82, 0.85, 0.77, 0.69, 0.76, 0.69, 0.66, 0.68, 0.66, 0.75, 0.78, 
    0.67, 0.74, 0.76, 0.7, 0.71, 0.73, 0.68, 0.74, 0.78, 0.79, 0.73, 0.71, 
    0.7, 0.7, 0.72, 0.72, 0.7, 0.67, 0.64, 0.63, 0.6, 0.59, 0.56, 0.57, 0.61, 
    0.61, 0.64, 0.68, 0.72, 0.76, 0.76, 0.75, 0.77, 0.76, 0.76, 0.81, 0.84, 
    0.83, 0.83, 0.82, 0.8, 0.76, 0.78, 0.78, 0.77, 0.76, 0.76, 0.75, 0.74, 
    0.73, 0.71, 0.72, 0.72, 0.72, 0.75, 0.73, 0.72, 0.72, 0.72, 0.7, 0.68, 
    0.71, 0.7, 0.69, 0.72, 0.73, 0.78, 0.71, 0.68, 0.61, 0.59, 0.59, 0.58, 
    0.57, 0.59, 0.61, 0.69, 0.76, 0.77, 0.75, 0.74, 0.67, 0.69, 0.75, 0.81, 
    0.85, 0.79, 0.81, 0.79, 0.77, 0.83, 0.77, 0.81, 0.8, 0.83, 0.79, 0.81, 
    0.78, 0.8, 0.79, 0.79, 0.8, 0.85, 0.83, 0.84, 0.85, 0.85, 0.82, 0.82, 
    0.79, 0.8, 0.84, 0.87, 0.86, 0.82, 0.76, 0.75, 0.71, 0.74, 0.73, 0.72, 
    0.71, 0.72, 0.77, 0.76, 0.77, 0.75, 0.77, 0.77, 0.8, 0.82, 0.82, 0.82, 
    0.79, 0.76, 0.75, 0.71, 0.83, 0.82, 0.86, 0.83, 0.83, 0.84, 0.84, 0.88, 
    0.87, 0.85, 0.84, 0.88, 0.85, 0.89, 0.92, 0.94, 0.96, 0.95, 0.96, 0.96, 
    0.94, 0.95, 0.93, 0.93, 0.94, 0.93, 0.93, 0.94, 0.94, 0.9, 0.86, 0.82, 
    0.82, 0.84, 0.85, 0.84, 0.87, 0.88, 0.87, 0.87, 0.88, 0.89, 0.88, 0.88, 
    0.87, 0.85, 0.85, 0.85, 0.83, 0.84, 0.83, 0.8, 0.78, 0.8, 0.79, 0.85, 
    0.84, 0.83, 0.83, 0.81, 0.82, 0.82, 0.84, 0.86, 0.79, 0.84, 0.83, 0.82, 
    0.85, 0.83, 0.81, 0.82, 0.79, 0.8, 0.81, 0.81, 0.78, 0.76, 0.72, 0.79, 
    0.71, 0.73, 0.83, 0.86, 0.81, 0.87, 0.88, 0.87, 0.84, 0.85, 0.87, 0.87, 
    0.84, 0.84, 0.87, 0.83, 0.84, 0.77, 0.74, 0.71, 0.72, 0.7, 0.73, 0.71, 
    0.73, 0.77, 0.77, 0.85, 0.88, 0.9, 0.9, 0.91, 0.88, 0.85, 0.84, 0.85, 
    0.84, 0.83, 0.87, 0.87, 0.87, 0.83, 0.78, 0.86, 0.8, 0.86, 0.77, 0.84, 
    0.78, 0.84, 0.86, 0.84, 0.86, 0.82, 0.83, 0.88, 0.89, 0.87, 0.89, 0.87, 
    0.82, 0.86, 0.86, 0.88, 0.83, 0.85, 0.83, 0.83, 0.84, 0.85, 0.81, 0.8, 
    0.72, 0.76, 0.81, 0.8, 0.83, 0.84, 0.82, 0.82, 0.84, 0.86, 0.85, 0.86, 
    0.85, 0.92, 0.88, 0.84, 0.84, 0.86, 0.84, 0.83, 0.84, 0.82, 0.78, 0.79, 
    0.8, 0.79, 0.75, 0.74, 0.76, 0.76, 0.78, 0.78, 0.88, 0.88, 0.91, 0.86, 
    0.84, 0.85, 0.84, 0.85, 0.82, 0.82, 0.79, 0.77, 0.75, 0.78, 0.77, 0.81, 
    0.81, 0.82, 0.79, 0.8, 0.78, 0.82, 0.82, 0.84, 0.85, 0.88, 0.89, 0.9, 
    0.9, 0.89, 0.89, 0.88, 0.87, 0.84, 0.82, 0.78, 0.8, 0.83, 0.79, 0.79, 
    0.8, 0.81, 0.79, 0.8, 0.8, 0.8, 0.83, 0.81, 0.83, 0.84, 0.87, 0.89, 0.87, 
    0.88, 0.88, 0.87, 0.85, 0.84, 0.84, 0.86, 0.87, 0.87, 0.88, 0.88, 0.88, 
    0.9, 0.92, 0.91, 0.92, 0.92, 0.92, 0.91, 0.9, 0.9, 0.92, 0.9, 0.9, 0.91, 
    0.91, 0.9, 0.89, 0.9, 0.9, 0.92, 0.92, 0.93, 0.94, 0.95, 0.93, 0.9, 0.88, 
    0.85, 0.89, 0.87, 0.89, 0.88, 0.86, 0.82, 0.74, 0.88, 0.85, 0.82, 0.84, 
    0.84, 0.87, 0.89, 0.92, 0.83, 0.84, 0.85, 0.85, 0.85, 0.85, 0.86, 0.87, 
    0.86, 0.9, 0.89, 0.88, 0.91, 0.9, 0.88, 0.89, 0.89, 0.85, 0.79, 0.87, 
    0.88, 0.87, 0.88, 0.88, 0.87, 0.82, 0.85, 0.83, 0.8, 0.74, 0.88, 0.84, 
    0.89, 0.88, 0.88, 0.89, 0.9, 0.9, 0.94, 0.95, 0.91, 0.85, 0.91, 0.89, 
    0.87, 0.9, 0.87, 0.9, 0.8, 0.89, 0.91, 0.92, 0.94, 0.94, 0.93, 0.93, 
    0.87, 0.87, 0.93, 0.9, 0.94, 0.93, 0.93, 0.95, 0.96, 0.95, 0.94, 0.94, 
    0.93, 0.93, 0.89, 0.86, 0.88, 0.88, 0.82, 0.82, 0.88, 0.9, 0.91, 0.92, 
    0.92, 0.93, 0.94, 0.91, 0.91, 0.91, 0.91, 0.9, 0.92, 0.88, 0.89, 0.89, 
    0.92, 0.9, 0.88, 0.82, 0.84, 0.83, 0.84, 0.86, 0.87, 0.88, 0.91, 0.91, 
    0.83, 0.84, 0.89, 0.87, 0.9, 0.89, 0.87, 0.9, 0.9, 0.91, 0.92, 0.94, 
    0.93, 0.93, 0.91, 0.89, 0.86, 0.8, 0.73, 0.8, 0.84, 0.86, 0.86, 0.85, 
    0.86, 0.89, 0.92, 0.93, 0.95, 0.96, 0.94, 0.92, 0.92, 0.91, 0.89, 0.82, 
    0.86, 0.82, 0.86, 0.89, 0.83, 0.82, 0.9, 0.9, 0.87, 0.87, 0.89, 0.9, 0.9, 
    0.92, 0.91, 0.91, 0.92, 0.92, 0.91, 0.89, 0.94, 0.91, 0.9, 0.9, 0.88, 
    0.86, 0.84, 0.82, 0.79, 0.78, 0.76, 0.77, 0.77, 0.72, 0.72, 0.73, 0.76, 
    0.81, 0.83, 0.82, 0.83, 0.84, 0.84, 0.88, 0.91, 0.92, 0.91, 0.92, 0.89, 
    0.85, 0.84, 0.8, 0.81, 0.86, 0.9, 0.94, 0.97, 0.97, 0.97, 0.97, 0.96, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.95, 0.94, 
    0.92, 0.88, 0.86, 0.87, 0.94, 0.95, 0.95, 0.95, 0.94, 0.94, 0.93, 0.9, 
    0.9, 0.91, 0.92, 0.92, 0.91, 0.97, 0.97, 0.97, 0.93, 0.87, 0.82, 0.79, 
    0.7, 0.77, 0.78, 0.72, 0.78, 0.81, 0.89, 0.89, 0.95, 0.96, 0.97, 0.97, 
    0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 
    0.99, 0.98, 0.97, 0.97, 0.93, 0.89, 0.92, 0.88, 0.88, 0.9, 0.91, 0.91, 
    0.87, 0.84, 0.83, 0.85, 0.86, 0.86, 0.88, 0.87, 0.89, 0.88, 0.87, 0.87, 
    0.84, 0.85, 0.84, 0.83, 0.83, 0.84, 0.84, 0.83, 0.82, 0.81, 0.82, 0.83, 
    0.84, 0.84, 0.86, 0.83, 0.83, 0.81, 0.85, 0.83, 0.84, 0.84, 0.84, 0.83, 
    0.84, 0.89, 0.93, 0.87, 0.93, 0.93, 0.93, 0.93, 0.93, 0.87, 0.88, 0.88, 
    0.85, 0.8, 0.82, 0.84, 0.85, 0.86, 0.88, 0.85, 0.86, 0.87, 0.88, 0.91, 
    0.89, 0.9, 0.92, 0.95, 0.97, 0.95, 0.98, 0.98, 0.97, 0.96, 0.96, 0.89, 
    0.92, 0.92, 0.93, 0.88, 0.85, 0.83, 0.86, 0.84, 0.86, 0.91, 0.89, 0.9, 
    0.9, 0.92, 0.93, 0.94, 0.92, 0.91, 0.9, 0.87, 0.83, 0.87, 0.89, 0.89, 
    0.91, 0.91, 0.94, 0.9, 0.84, 0.8, 0.73, 0.71, 0.81, 0.83, 0.81, 0.83, 
    0.94, 0.95, 0.92, 0.92, 0.93, 0.94, 0.96, 0.93, 0.9, 0.9, 0.85, 0.84, 
    0.84, 0.81, 0.79, 0.83, 0.87, 0.87, 0.89, 0.89, 0.88, 0.88, 0.89, 0.93, 
    0.92, 0.91, 0.89, 0.84, 0.87, 0.79, 0.78, 0.81, 0.82, 0.78, 0.8, 0.81, 
    0.86, 0.9, 0.91, 0.9, 0.81, 0.8, 0.86, 0.83, 0.84, 0.84, 0.84, 0.82, 
    0.81, 0.81, 0.8, 0.79, 0.79, 0.79, 0.76, 0.85, 0.78, 0.83, 0.79, 0.71, 
    0.74, 0.76, 0.72, 0.7, 0.74, 0.74, 0.76, 0.75, 0.82, 0.85, 0.85, 0.86, 
    0.86, 0.81, 0.77, 0.8, 0.79, 0.78, 0.82, 0.88, 0.9, 0.93, 0.93, 0.94, 
    0.94, 0.91, 0.89, 0.91, 0.88, 0.88, 0.87, 0.85, 0.85, 0.83, 0.81, 0.8, 
    0.74, 0.79, 0.78, 0.78, 0.76, 0.81, 0.81, 0.86, 0.87, 0.85, 0.9, 0.9, 
    0.9, 0.91, 0.91, 0.91, 0.91, 0.92, 0.93, 0.91, 0.92, 0.92, 0.92, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 
    0.91, 0.91, 0.91, 0.89, 0.89, 0.9, 0.9, 0.88, 0.88, 0.87, 0.87, 0.88, 
    0.86, 0.87, 0.88, 0.89, 0.91, 0.89, 0.88, 0.86, 0.85, 0.84, 0.81, 0.81, 
    0.8, 0.86, 0.83, 0.88, 0.91, 0.92, 0.92, 0.93, 0.92, 0.9, 0.92, 0.93, 
    0.88, 0.9, 0.89, 0.9, 0.95, 0.94, 0.91, 0.91, 0.93, 0.87, 0.86, 0.84, 
    0.88, 0.83, 0.84, 0.85, 0.85, 0.87, 0.87, 0.84, 0.88, 0.87, 0.89, 0.9, 
    0.84, 0.89, 0.9, 0.92, 0.91, 0.9, 0.9, 0.92, 0.92, 0.93, 0.94, 0.92, 
    0.92, 0.92, 0.9, 0.89, 0.9, 0.89, 0.89, 0.91, 0.9, 0.9, 0.88, 0.91, 0.92, 
    0.88, 0.92, 0.92, 0.9, 0.94, 0.95, 0.94, 0.9, 0.92, 0.92, 0.81, 0.88, 
    0.84, 0.87, 0.84, 0.78, 0.79, 0.78, 0.84, 0.85, 0.88, 0.91, 0.89, 0.89, 
    0.84, 0.83, 0.89, 0.89, 0.93, 0.93, 0.94, 0.94, 0.92, 0.92, 0.94, 0.92, 
    0.88, 0.9, 0.89, 0.9, 0.91, 0.9, 0.89, 0.89, 0.89, 0.89, 0.88, 0.94, 
    0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 
    0.96, 0.96, 0.96, 0.95, 0.94, 0.95, 0.95, 0.92, 0.93, 0.95, 0.93, 0.93, 
    0.89, 0.89, 0.89, 0.88, 0.87, 0.89, 0.9, 0.92, 0.88, 0.91, 0.93, 0.86, 
    0.82, 0.84, 0.87, 0.79, 0.78, 0.8, 0.8, 0.81, 0.83, 0.85, 0.93, 0.94, 
    0.92, 0.94, 0.91, 0.79, 0.9, 0.81, 0.77, 0.88, 0.91, 0.83, 0.87, 0.88, 
    0.84, 0.82, 0.79, 0.81, 0.81, 0.81, 0.81, 0.83, 0.85, 0.88, 0.92, 0.92, 
    0.94, 0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.93, 0.93, 0.92, 
    0.93, 0.94, 0.96, 0.95, 0.96, 0.97, 0.95, 0.94, 0.95, 0.95, 0.96, 0.96, 
    0.95, 0.96, 0.97, 0.97, 0.97, 0.98, 0.97, 0.97, 0.97, 0.94, 0.93, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.93, 0.92, 0.95, 0.96, 0.96, 0.91, 
    0.9, 0.91, 0.91, 0.87, 0.91, 0.93, 0.95, 0.9, 0.95, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.96, 0.97, 0.97, 0.97, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.96, 0.96, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.94, 0.9, 0.87, 0.92, 0.92, 0.91, 
    0.92, 0.9, 0.91, 0.88, 0.92, 0.87, 0.91, 0.94, 0.9, 0.94, 0.96, 0.97, 
    0.97, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.96, 0.93, 0.96, 
    0.93, 0.9, 0.92, 0.93, 0.94, 0.93, 0.93, 0.95, 0.97, 0.97, 0.96, 0.92, 
    0.87, 0.95, 0.98, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.96, 
    0.95, 0.97, 0.97, 0.98, 0.97, 0.96, 0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 
    0.96, 0.9, 0.87, 0.88, 0.91, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.93, 
    0.94, 0.91, 0.93, 0.94, 0.94, 0.92, 0.94, 0.92, 0.92, 0.9, 0.93, 0.91, 
    0.86, 0.94, 0.93, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.95, 0.94, 
    0.92, 0.93, 0.94, 0.92, 0.94, 0.93, 0.96, 0.96, 0.97, 0.98, 0.97, 0.96, 
    0.96, 0.97, 0.98, 0.97, 0.93, 0.94, 0.96, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.96, 0.93, 0.92, 0.93, 0.96, 0.96, 0.97, 0.96, 0.91, 0.95, 0.97, 0.92, 
    0.92, 0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 
    0.95, 0.95, 0.94, 0.96, 0.93, 0.91, 0.96, 0.91, 0.91, 0.93, 0.96, 0.97, 
    0.98, 0.98, 0.99, 0.97, 0.97, 0.96, 0.92, 0.93, 0.94, 0.95, 0.97, 0.98, 
    0.98, 0.97, 0.97, 0.97, 0.97, 0.95, 0.93, 0.94, 0.93, 0.89, 0.94, 0.95, 
    0.93, 0.93, 0.95, 0.95, 0.93, 0.88, 0.87, 0.76, 0.78, 0.73, 0.73, 0.74, 
    0.77, 0.82, 0.8, 0.89, 0.81, 0.91, 0.82, 0.83, 0.88, 0.9, 0.92, 0.95, 
    0.94, 0.94, 0.94, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.97, 0.96, 0.95, 0.94, 0.93, 0.96, 0.98, 0.95, 0.94, 0.94, 
    0.94, 0.92, 0.96, 0.97, 0.98, 0.99, 0.93, 0.97, 0.97, 0.98, 0.99, 0.99, 
    0.98, 0.98, 0.95, 0.96, 0.96, 0.97, 0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.95, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.96, 0.96, 0.96, 0.97, 0.96, 0.96, 0.98, 0.98, 0.98, 0.97, 0.97, 
    0.95, 0.95, 0.95, 0.95, 0.96, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 
    0.97, 0.98, 0.98, 0.97, 0.98, 0.97, 0.97, 0.97, 0.97, 0.96, 0.97, 0.97, 
    0.98, 0.98, 0.93, 0.92, 0.92, 0.93, 0.94, 0.95, 0.92, 0.89, 0.91, 0.91, 
    0.9, 0.9, 0.94, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.96, 0.96, 0.97, 
    0.94, 0.93, 0.94, 0.94, 0.95, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.97, 0.97, 0.95, 
    0.96, 0.93, 0.94, 0.95, 0.96, 0.94, 0.92, 0.95, 0.95, 0.94, 0.94, 0.97, 
    0.95, 0.97, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.96, 0.98, 0.99, 0.98, 0.96, 0.96, 0.97, 0.95, 0.97, 0.98, 0.98, 
    0.97, 0.96, 0.9, 0.93, 0.92, 0.9, 0.93, 0.93, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.93, 0.93, 0.93, 0.92, 0.92, 0.9, 0.85, 0.84, 0.82, 0.88, 0.88, 
    0.82, 0.83, 0.88, 0.87, 0.84, 0.85, 0.83, 0.85, 0.85, 0.87, 0.9, 0.9, 
    0.88, 0.88, 0.89, 0.87, 0.89, 0.89, 0.93, 0.92, 0.94, 0.97, 0.98, 0.99, 
    0.97, 0.96, 0.9, 0.86, 0.87, 0.91, 0.92, 0.96, 0.98, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.97, 0.98, 0.97, 0.99, 0.99, 0.99, 0.99, 0.98, 0.96, 0.94, 
    0.94, 0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 0.92, 0.96, 0.97, 0.98, 0.98, 
    0.97, 0.95, 0.94, 0.94, 0.97, 0.98, 0.99, 0.98, 0.98, 0.98, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.98, 0.99, 0.96, 0.98, 0.95, 0.99, 0.96, 0.95, 0.98, 0.91, 
    0.94, 0.94, 0.91, 0.87, 0.92, 0.94, 0.93, 0.92, 0.88, 0.94, 0.95, 0.92, 
    0.96, 0.97, 0.97, 0.96, 0.98, 0.94, 0.99, 0.98, 0.98, 0.96, 0.94, 0.98, 
    0.97, 0.98, 0.98, 0.97, 0.97, 0.93, 0.93, 0.93, 0.95, 0.92, 0.96, 0.96, 
    0.97, 0.96, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.95, 
    0.93, 0.86, 0.87, 0.97, 0.95, 0.94, 0.94, 0.96, 0.96, 0.98, 0.97, 0.98, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 
    0.98, 0.98, 0.96, 0.94, 0.94, 0.94, 0.97, 0.98, 0.99, 0.98, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.96, 0.97, 0.96, 0.96, 
    0.96, 0.93, 0.92, 0.93, 0.93, 0.94, 0.93, 0.94, 0.95, 0.96, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.96, 0.94, 0.95, 
    0.93, 0.96, 0.94, 0.96, 0.94, 0.88, 0.91, 0.93, 0.91, 0.95, 0.94, 0.93, 
    0.93, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 0.95, 
    0.91, 0.85, 0.88, 0.92, 0.89, 0.88, 0.89, 0.92, 0.92, 0.88, 0.87, 0.87, 
    0.85, 0.81, 0.79, 0.81, 0.85, 0.9, 0.89, 0.91, 0.89, 0.88, 0.9, 0.96, 
    0.88, 0.9, 0.92, 0.94, 0.92, 0.9, 0.9, 0.92, 0.89, 0.88, 0.89, 0.93, 
    0.92, 0.92, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.94, 0.94, 0.99, 0.99, 0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.95, 0.95, 0.95, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 0.93, 0.91, 0.89, 0.9, 
    0.97, 0.98, 0.89, 0.97, 0.96, 0.9, 0.91, 0.92, 0.92, 0.92, 0.93, 0.93, 
    0.94, 0.94, 0.95, 0.95, 0.95, 0.96, 0.96, 0.95, 0.94, 0.94, 0.9, 0.9, 
    0.99, 0.99, 0.99, 0.97, 0.96, 0.94, 0.93, 0.91, 0.91, 0.91, 0.91, 0.91, 
    0.93, 0.98, 0.99, 0.99, 0.98, 0.95, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.95, 0.95, 0.96, 0.97, 0.91, 0.89, 0.9, 0.89, 0.9, 
    0.84, 0.83, 0.88, 0.89, 0.92, 0.9, 0.91, 0.89, 0.88, 0.87, 0.92, 0.86, 
    0.85, 0.84, 0.9, 0.92, 0.87, 0.87, 0.89, 0.92, 0.93, 0.95, 0.94, 0.94, 
    0.97, 0.95, 0.93, 0.92, 0.94, 0.95, 0.96, 0.96, 0.95, 0.95, 0.93, 0.94, 
    0.94, 0.93, 0.9, 0.9, 0.91, 0.92, 0.91, 0.91, 0.9, 0.9, 0.91, 0.95, 0.95, 
    0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.93, 0.91, 0.9, 0.94, 
    0.93, 0.93, 0.92, 0.92, 0.93, 0.92, 0.92, 0.92, 0.92, 0.94, 0.94, 0.94, 
    1, 0.99, 0.98, 0.97, 0.96, 0.95, 0.88, 0.87, 0.95, 0.94, 0.93, 0.88, 
    0.88, 0.87, 0.83, 0.85, 0.87, 0.91, 0.88, 0.94, 0.91, 0.95, 0.96, 0.96, 
    0.97, 0.96, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 
    0.97, 0.96, 0.95, 0.95, 0.96, 0.96, 0.96, 0.93, 0.9, 0.87, 0.85, 0.85, 
    0.87, 0.88, 0.89, 0.89, 0.89, 0.91, 0.91, 0.88, 0.87, 0.87, 0.88, 0.93, 
    0.97, 0.93, 0.9, 0.96, 0.94, 0.94, 0.96, 0.95, 0.95, 0.95, 0.96, 0.98, 
    0.97, 0.92, 0.94, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.99, 0.97, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 0.99, 0.99, 1, 0.99, 1, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.98, 
    0.97, 0.96, 0.96, 0.96, 0.96, 0.92, 0.89, 0.96, 0.98, 0.97, 0.96, 0.96, 
    0.99, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.96, 0.89, 
    0.88, 0.93, 0.95, 0.96, 0.89, 0.91, 0.93, 0.97, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 1, 0.99, 0.99, 0.95, 0.95, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.95, 0.91, 0.92, 0.98, 0.98, 0.98, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.99, 
    0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.98, 0.98, 0.98, 0.99, 0.98, 
    0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 
    0.97, 0.99, 0.99, 0.99, 0.98, 0.99, 0.98, 0.98, 0.97, 0.97, 0.98, 0.95, 
    0.9, 0.94, 0.95, 0.96, 0.96, 0.94, 0.95, 0.95, 0.96, 0.97, 0.97, 0.97, 
    0.98, 0.97, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 
    0.94, 0.93, 0.93, 0.94, 0.95, 0.93, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.96, 0.95, 0.94, 0.93, 0.96, 0.93, 0.94, 0.93, 0.93, 0.93, 0.92, 
    0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.95, 
    0.94, 0.95, 0.95, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 
    0.99, 0.98, 0.99, 0.99, 0.9, 0.92, 0.95, 0.98, 0.98, 0.98, 0.97, 0.97, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.97, 0.98, 0.98, 0.97, 0.97, 
    0.96, 0.96, 0.96, 0.95, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 
    0.97, 0.96, 0.96, 0.96, 0.95, 0.95, 0.94, 0.93, 0.93, 0.94, 0.95, 0.97, 
    0.96, 0.95, 0.94, 0.95, 0.96, 0.98, 0.98, 0.97, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 
    0.94, 0.94, 0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.91, 0.91, 0.94, 
    0.96, 0.96, 0.9, 0.92, 0.95, 0.95, 0.91, 0.94, 0.92, 0.94, 0.9, 0.95, 
    0.94, 0.93, 0.92, 0.96, 0.96, 0.96, 0.95, 0.95, 0.9, 0.9, 0.98, 0.98, 
    0.97, 0.92, 0.91, 0.9, 0.89, 0.9, 0.89, 0.92, 0.91, 0.91, 0.91, 0.94, 
    0.94, 0.95, 0.95, 0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 0.98, 0.97, 0.97, 
    0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 0.97, 0.98, 0.98, 0.98, 
    0.99, 0.99, 1, 1, 0.99, 0.97, 1, 1, 0.97, 1, 1, 0.97, 0.97, 1, 0.99, 
    0.99, 0.96, 1, 0.93, 0.85, 0.85, 0.93, 0.9, 0.85, 0.83, 0.85, 0.84, 0.87, 
    0.87, 0.95, 0.93, 0.95, 0.98, 0.94, 0.95, 0.95, 0.93, 0.92, 0.93, 0.92, 
    0.93, 0.9, 0.92, 0.91, 0.91, 0.91, 0.94, 0.91, 0.89, 0.88, 0.87, 0.87, 
    0.86, 0.78, 0.76, 0.85, 0.86, 0.84, 0.81, 0.81, 0.81, 0.84, 0.86, 0.96, 
    0.99, 0.96, 0.94, 0.93, 0.94, 0.92, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 
    0.97, 0.95, 0.94, 0.96, 0.96, 0.94, 0.94, 0.97, 0.97, 0.95, 0.92, 0.91, 
    0.93, 0.94, 0.93, 0.93, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.93, 0.89, 
    0.92, 0.92, 0.95, 0.93, 0.93, 0.95, 0.92, 0.92, 0.93, 0.92, 0.94, 0.94, 
    0.93, 0.93, 0.92, 0.89, 0.85, 0.84, 0.87, 0.81, 0.87, 0.91, 0.93, 0.95, 
    0.96, 0.95, 0.9, 0.93, 0.92, 0.92, 0.9, 0.92, 0.93, 0.94, 0.97, 0.93, 
    0.89, 0.87, 0.82, 0.8, 0.88, 0.95, 0.95, 0.94, 0.9, 0.91, 0.9, 0.93, 
    0.93, 0.92, 0.93, 0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 
    0.91, 0.91, 0.91, 0.91, 0.88, 0.89, 0.87, 0.87, 0.79, 0.81, 0.83, 0.85, 
    0.88, 0.88, 0.87, 0.88, 0.89, 0.91, 0.94, 0.95, 0.97, 0.97, 0.95, 0.93, 
    0.92, 0.9, 0.88, 0.81, 0.84, 0.88, 0.92, 0.93, 0.97, 0.98, 0.96, 0.96, 
    0.95, 0.96, 0.96, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.99, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 
    0.98, 0.99, 0.99, 1, 0.99, 0.99, 1, 1, 1, 0.98, 0.96, 0.94, 0.91, 0.91, 
    0.9, 0.9, 0.9, 0.9, 0.92, 0.92, 0.91, 0.89, 0.91, 0.9, 0.89, 0.88, 0.88, 
    0.89, 0.86, 0.86, 0.86, 0.89, 0.87, 0.86, 0.82, 0.83, 0.92, 0.91, 0.89, 
    0.89, 0.87, 0.84, 0.82, 0.84, 0.86, 0.9, 0.92, 0.93, 0.93, 0.92, 0.91, 
    0.93, 0.92, 0.9, 0.86, 0.85, 0.85, 0.86, 0.86, 0.83, 0.84, 0.92, 0.87, 
    0.86, 0.87, 0.87, 0.89, 0.92, 0.91, 0.87, 0.85, 0.84, 0.82, 0.79, 0.83, 
    0.85, 0.95, 0.94, 0.95, 0.94, 0.93, 0.94, 0.95, 0.93, 0.92, 0.95, 0.96, 
    0.97, 0.97, 0.98, 0.98, 0.99, 0.99, 0.97, 0.88, 0.9, 0.88, 0.87, 0.87, 
    0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.91, 0.91, 0.83, 0.84, 0.8, 0.83, 
    0.87, 0.91, 0.92, 0.91, 0.89, 0.88, 0.85, 0.87, 0.9, 0.94, 0.91, 0.93, 
    0.94, 0.92, 0.92, 0.96, 0.96, 0.96, 0.96, 0.96, 0.95, 0.95, 0.96, 0.96, 
    0.96, 0.96, 0.95, 0.92, 0.9, 0.9, 0.93, 0.94, 0.95, 0.95, 0.81, 0.9, 
    0.88, 0.87, 0.89, 0.92, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0.98, 0.98, 0.98, 1, 1, 1, 1, 1, 0.98, 0.99, 0.99, 
    1, 0.99, 0.99, 0.99, 0.99, 0.98, 0.92, 0.93, 0.87, 0.88, 0.87, 0.88, 
    0.86, 0.88, 0.87, 0.89, 0.9, 0.91, 0.9, 0.91, 0.93, 0.95, 0.98, 0.97, 
    0.96, 0.99, 0.98, 0.99, 0.99, 0.98, 0.97, 0.96, 0.94, 0.92, 0.93, 0.94, 
    0.95, 0.95, 0.93, 0.92, 0.93, 0.83, 0.82, 0.93, 0.94, 0.88, 0.84, 0.86, 
    0.91, 0.94, 0.97, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 1, 0.97, 
    0.98, 0.98, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.95, 0.98, 0.98, 0.94, 0.93, 
    0.92, 0.93, 0.96, 0.92, 0.95, 0.96, 0.93, 0.85, 0.81, 0.76, 0.75, 0.92, 
    0.88, 0.91, 0.92, 0.83, 0.9, 0.89, 0.85, 0.85, 0.86, 0.92, 0.94, 0.94, 
    0.93, 0.9, 0.91, 0.9, 0.9, 0.85, 0.84, 0.86, 0.86, 0.87, 0.86, 0.95, 
    0.95, 0.95, 0.95, 0.96, 0.96, 0.95, 0.96, 0.94, 0.93, 0.92, 0.91, 0.9, 
    0.9, 0.88, 0.88, 0.88, 0.84, 0.82, 0.82, 0.91, 0.91, 0.91, 0.92, 0.92, 
    0.92, 0.93, 0.93, 0.86, 0.87, 0.89, 0.87, 0.87, 0.89, 0.87, 0.87, 0.83, 
    0.86, 0.87, 0.88, 0.87, 0.86, 0.86, 0.88, 0.9, 0.91, 0.92, 0.9, 0.89, 
    0.87, 0.85, 0.9, 0.89, 0.88, 0.87, 0.87, 0.86, 0.86, 0.84, 0.84, 0.85, 
    0.84, 0.84, 0.9, 0.89, 0.89, 0.9, 0.9, 0.89, 0.91, 0.89, 0.89, 0.88, 
    0.92, 0.92, 0.93, 0.93, 0.93, 0.73, 0.74, 0.8, 0.84, 0.79, 0.83, 0.84, 
    0.85, 0.9, 0.89, 0.88, 0.88, 0.89, 0.76, 0.77, 0.79, 0.82, 0.82, 0.79, 
    0.79, 0.79, 0.79, 0.8, 0.82, 0.84, 0.85, 0.85, 0.86, 0.85, 0.86, 0.87, 
    0.88, 0.89, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.91, 0.91, 0.92, 0.9, 
    0.9, 0.9, 0.89, 0.89, 0.89, 0.88, 0.87, 0.86, 0.86, 0.86, 0.86, 0.85, 
    0.86, 0.87, 0.89, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 0.93, 0.94, 
    0.94, 0.93, 0.91, 0.89, 0.88, 0.84, 0.83, 0.84, 0.86, 0.88, 0.91, 0.89, 
    0.86, 0.87, 0.89, 0.91, 0.93, 0.93, 0.93, 0.96, 0.94, 0.95, 0.96, 0.95, 
    0.96, 0.95, 0.98, 0.98, 0.98, 0.98, 0.96, 0.94, 0.94, 0.97, 0.94, 0.91, 
    0.89, 0.93, 0.95, 0.91, 0.92, 0.93, 0.91, 0.91, 0.94, 0.92, 0.92, 0.91, 
    0.97, 0.94, 0.92, 0.98, 0.97, 0.95, 0.98, 0.99, 0.98, 0.97, 0.97, 0.96, 
    0.96, 0.96, 0.93, 0.94, 0.93, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.95, 
    0.94, 0.94, 0.95, 0.95, 0.94, 0.94, 0.93, 0.93, 0.93, 0.9, 0.9, 0.9, 0.9, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 0.94, 0.86, 0.94, 0.93, 
    0.91, 0.88, 0.91, 0.92, 0.91, 0.89, 0.89, 0.87, 0.85, 0.81, 0.81, 0.83, 
    0.85, 0.86, 0.87, 0.9, 0.89, 0.87, 0.86, 0.85, 0.84, 0.85, 0.85, 0.88, 
    0.88, 0.89, 0.89, 0.88, 0.76, 0.82, 0.79, 0.78, 0.82, 0.76, 0.79, 0.74, 
    0.8, 0.74, 0.77, 0.81, 0.83, 0.84, 0.85, 0.86, 0.87, 0.8, 0.8, 0.8, 0.8, 
    0.86, 0.86, 0.86, 0.86, 0.86, 0.85, 0.8, 0.8, 0.77, 0.76, 0.78, 0.78, 
    0.81, 0.82, 0.81, 0.79, 0.8, 0.89, 0.86, 0.82, 0.83, 0.84, 0.85, 0.92, 
    0.92, 0.86, 0.87, 0.88, 0.89, 0.9, 0.89, 0.9, 0.92, 0.94, 0.94, 0.94, 
    0.94, 0.93, 0.93, 0.94, 0.92, 0.9, 0.94, 0.95, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.93, 0.97, 0.96, 0.96, 0.95, 0.94, 0.92, 0.95, 0.94, 0.94, 0.94, 
    0.94, 0.92, 0.91, 0.92, 0.92, 0.93, 0.93, 0.91, 0.94, 0.94, 0.95, 0.94, 
    0.87, 0.87, 0.86, 0.87, 0.9, 0.92, 0.93, 0.94, 0.93, 0.92, 0.9, 0.88, 
    0.89, 0.83, 0.91, 0.92, 0.94, 0.91, 0.93, 0.97, 0.98, 0.95, 0.97, 0.96, 
    0.99, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    1, 1, 0.98, 0.94, 0.93, 0.93, 0.92, 0.92, 0.92, 0.94, 0.95, 0.95, 0.95, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.95, 0.95, 0.93, 0.92, 0.94, 0.96, 0.96, 
    0.96, 0.97, 0.95, 0.93, 0.91, 0.89, 0.88, 0.87, 0.88, 0.9, 0.86, 0.87, 
    0.89, 0.91, 0.89, 0.9, 0.87, 0.93, 0.94, 0.94, 0.88, 0.95, 0.95, 0.95, 
    0.93, 0.94, 0.93, 0.93, 0.94, 0.92, 0.91, 0.9, 0.89, 0.89, 0.88, 0.87, 
    0.88, 0.9, 0.9, 0.91, 0.92, 0.9, 0.87, 0.86, 0.85, 0.84, 0.77, 0.78, 
    0.81, 0.84, 0.8, 0.8, 0.8, 0.73, 0.73, 0.75, 0.74, 0.77, 0.72, 0.73, 
    0.75, 0.76, 0.83, 0.81, 0.79, 0.79, 0.78, 0.8, 0.83, 0.84, 0.85, 0.8, 
    0.79, 0.78, 0.8, 0.83, 0.85, 0.9, 0.92, 0.87, 0.89, 0.91, 0.93, 0.93, 
    0.92, 0.93, 0.96, 0.96, 0.97, 0.98, 0.98, 0.97, 0.96, 0.95, 0.94, 0.93, 
    0.89, 0.9, 0.89, 0.88, 0.88, 0.91, 0.91, 0.91, 0.89, 0.89, 0.9, 0.9, 
    0.89, 0.88, 0.87, 0.9, 0.88, 0.87, 0.89, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.87, 0.86, 0.87, 0.88, 0.85, 0.85, 0.84, 0.83, 0.82, 0.82, 0.83, 
    0.84, 0.85, 0.84, 0.86, 0.83, 0.84, 0.85, 0.83, 0.83, 0.86, 0.87, 0.88, 
    0.87, 0.87, 0.81, 0.79, 0.79, 0.8, 0.8, 0.8, 0.79, 0.86, 0.88, 0.88, 
    0.87, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.9, 0.92, 0.87, 0.88, 0.88, 0.86, 
    0.86, 0.88, 0.88, 0.87, 0.88, 0.89, 0.89, 0.89, 0.87, 0.87, 0.87, 0.86, 
    0.86, 0.88, 0.88, 0.85, 0.86, 0.85, 0.84, 0.85, 0.85, 0.88, 0.89, 0.87, 
    0.89, 0.88, 0.87, 0.87, 0.87, 0.86, 0.86, 0.86, 0.86, 0.87, 0.88, 0.88, 
    0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.91, 0.89, 0.89, 0.9, 0.9, 0.9, 0.9, 
    0.9, 0.9, 0.9, 0.91, 0.91, 0.84, 0.84, 0.84, 0.9, 0.9, 0.9, 0.89, 0.9, 
    0.91, 0.9, 0.9, 0.89, 0.89, 0.9, 0.91, 0.89, 0.9, 0.91, 0.92, 0.91, 0.91, 
    0.91, 0.91, 0.85, 0.9, 0.9, 0.9, 0.91, 0.91, 0.9, 0.92, 0.9, 0.86, 0.87, 
    0.9, 0.92, 0.93, 0.93, 0.95, 0.96, 0.94, 0.94, 0.91, 0.9, 0.9, 0.89, 
    0.89, 0.88, 0.88, 0.87, 0.88, 0.87, 0.86, 0.87, 0.87, 0.87, 0.87, 0.86, 
    0.86, 0.87, 0.87, 0.87, 0.87, 0.87, 0.87, 0.88, 0.88, 0.91, 0.91, 0.83, 
    0.86, 0.86, 0.86, 0.86, 0.84, 0.83, 0.82, 0.79, 0.8, 0.8, 0.84, 0.84, 
    0.85, 0.83, 0.85, 0.91, 0.89, 0.88, 0.83, 0.83, 0.85, 0.86, 0.87, 0.87, 
    0.87, 0.87, 0.91, 0.91, 0.9, 0.92, 0.84, 0.88, 0.8, 0.9, 0.82, 0.84, 
    0.86, 0.88, 0.9, 0.9, 0.9, 0.91, 0.9, 0.91, 0.91, 0.92, 0.94, 0.95, 0.94, 
    0.94, 0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.88, 0.93, 0.91, 0.96, 0.98, 
    0.98, 0.97, 0.96, 0.95, 0.96, 0.95, 0.93, 0.92, 0.91, 0.98, 0.94, 0.94, 
    0.94, 0.88, 0.87, 0.86, 0.87, 0.89, 0.92, 0.95, 0.94, 0.91, 0.91, 0.94, 
    0.95, 0.95, 0.91, 0.91, 0.91, 0.91, 0.9, 0.92, 0.91, 0.9, 0.89, 0.88, 
    0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.94, 0.85, 0.86, 0.87, 0.88, 0.88, 
    0.88, 0.9, 0.91, 0.93, 0.93, 0.95, 0.92, 0.92, 0.92, 0.93, 0.97, 0.97, 
    0.95, 0.96, 0.96, 0.96, 0.97, 0.96, 0.95, 0.95, 0.94, 0.96, 0.96, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 
    0.95, 0.95, 0.95, 0.95, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.95, 0.97, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.95, 0.97, 0.97, 0.98, 0.96, 0.96, 0.93, 0.91, 0.93, 0.93, 0.93, 0.93, 
    0.93, 0.91, 0.92, 0.92, 0.92, 0.94, 0.94, 0.95, 0.95, 0.93, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.94, 0.93, 0.93, 0.93, 
    0.93, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.9, 0.9, 0.9, 0.92, 
    0.92, 0.88, 0.86, 0.89, 0.89, 0.89, 0.89, 0.88, 0.88, 0.89, 0.88, 0.89, 
    0.86, 0.81, 0.83, 0.85, 0.85, 0.8, 0.77, 0.79, 0.84, 0.82, 0.81, 0.8, 
    0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.77, 0.77, 0.77, 0.75, 0.77, 0.74, 
    0.74, 0.74, 0.76, 0.77, 0.78, 0.76, 0.77, 0.76, 0.74, 0.75, 0.71, 0.75, 
    0.75, 0.76, 0.78, 0.75, 0.79, 0.82, 0.81, 0.8, 0.78, 0.76, 0.71, 0.76, 
    0.71, 0.73, 0.72, 0.75, 0.7, 0.72, 0.74, 0.75, 0.75, 0.84, 0.87, 0.87, 
    0.85, 0.82, 0.8, 0.84, 0.8, 0.8, 0.79, 0.82, 0.81, 0.85, 0.85, 0.81, 0.8, 
    0.81, 0.81, 0.86, 0.9, 0.91, 0.92, 0.93, 0.9, 0.84, 0.92, 0.9, 0.93, 
    0.89, 0.9, 0.9, 0.9, 0.89, 0.86, 0.87, 0.87, 0.86, 0.85, 0.79, 0.74, 
    0.73, 0.76, 0.78, 0.77, 0.78, 0.79, 0.8, 0.76, 0.79, 0.78, 0.8, 0.8, 
    0.79, 0.84, 0.83, 0.79, 0.78, 0.79, 0.79, 0.78, 0.81, 0.76, 0.77, 0.75, 
    0.78, 0.8, 0.8, 0.82, 0.84, 0.83, 0.83, 0.83, 0.83, 0.84, 0.84, 0.84, 
    0.84, 0.85, 0.85, 0.76, 0.77, 0.81, 0.8, 0.8, 0.83, 0.83, 0.84, 0.82, 
    0.83, 0.84, 0.83, 0.82, 0.82, 0.82, 0.81, 0.83, 0.83, 0.82, 0.82, 0.8, 
    0.79, 0.82, 0.79, 0.81, 0.81, 0.81, 0.81, 0.77, 0.79, 0.79, 0.81, 0.78, 
    0.73, 0.68, 0.68, 0.66, 0.66, 0.61, 0.68, 0.74, 0.82, 0.81, 0.83, 0.82, 
    0.8, 0.8, 0.81, 0.82, 0.83, 0.84, 0.84, 0.86, 0.85, 0.84, 0.82, 0.81, 
    0.82, 0.82, 0.83, 0.83, 0.85, 0.84, 0.85, 0.87, 0.77, 0.78, 0.78, 0.78, 
    0.75, 0.81, 0.75, 0.76, 0.76, 0.79, 0.79, 0.81, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.81, 0.81, 0.81, 0.82, 0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 
    0.81, 0.82, 0.82, 0.82, 0.82, 0.83, 0.83, 0.83, 0.83, 0.83, 0.84, 0.84, 
    0.84, 0.84, 0.83, 0.82, 0.83, 0.83, 0.82, 0.82, 0.82, 0.83, 0.83, 0.84, 
    0.85, 0.85, 0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 0.88, 0.89, 0.89, 0.89, 
    0.89, 0.9, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 0.89, 
    0.89, 0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 0.86, 0.86, 0.85, 0.84, 0.85, 
    0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.82, 0.83, 0.82, 0.82, 0.82, 0.82, 
    0.82, 0.84, 0.83, 0.83, 0.83, 0.82, 0.81, 0.81, 0.82, 0.82, 0.82, 0.81, 
    0.83, 0.82, 0.82, 0.84, 0.83, 0.82, 0.84, 0.83, 0.84, 0.83, 0.82, 0.83, 
    0.84, 0.83, 0.82, 0.82, 0.83, 0.83, 0.83, 0.83, 0.83, 0.84, 0.83, 0.83, 
    0.83, 0.83, 0.83, 0.82, 0.82, 0.82, 0.81, 0.81, 0.82, 0.81, 0.81, 0.82, 
    0.82, 0.83, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.83, 0.82, 0.84, 0.82, 
    0.82, 0.83, 0.82, 0.83, 0.83, 0.83, 0.82, 0.82, 0.83, 0.83, 0.86, 0.84, 
    0.85, 0.84, 0.85, 0.85, 0.85, 0.85, 0.86, 0.86, 0.86, 0.85, 0.86, 0.85, 
    0.86, 0.86, 0.86, 0.86, 0.85, 0.86, 0.86, 0.86, 0.85, 0.86, 0.86, 0.86, 
    0.85, 0.85, 0.86, 0.85, 0.85, 0.85, 0.85, 0.86, 0.85, 0.84, 0.83, 0.83, 
    0.83, 0.83, 0.84, 0.85, 0.86, 0.86, 0.86, 0.87, 0.81, 0.8, 0.82, 0.81, 
    0.83, 0.85, 0.85, 0.86, 0.87, 0.88, 0.9, 0.91, 0.92, 0.93, 0.94, 0.94, 
    0.94, 0.95, 0.96, 0.96, 0.92, 0.88, 0.85, 0.85, 0.84, 0.82, 0.82, 0.77, 
    0.82, 0.83, 0.84, 0.82, 0.83, 0.85, 0.84, 0.83, 0.82, 0.82, 0.8, 0.82, 
    0.82, 0.82, 0.83, 0.85, 0.87, 0.83, 0.84, 0.87, 0.85, 0.85, 0.83, 0.82, 
    0.83, 0.84, 0.84, 0.84, 0.82, 0.79, 0.79, 0.79, 0.72, 0.7, 0.8, 0.81, 
    0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.85, 0.84, 0.84, 0.84, 0.84, 0.83, 
    0.83, 0.83, 0.82, 0.81, 0.8, 0.82, 0.81, 0.82, 0.82, 0.8, 0.8, 0.81, 
    0.78, 0.84, 0.84, 0.84, 0.84, 0.85, 0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 
    0.87, 0.87, 0.86, 0.86, 0.84, 0.83, 0.85, 0.85, 0.84, 0.82, 0.81, 0.81, 
    0.79, 0.81, 0.79, 0.8, 0.81, 0.77, 0.78, 0.77, 0.78, 0.76, 0.76, 0.77, 
    0.77, 0.76, 0.78, 0.75, 0.76, 0.78, 0.77, 0.77, 0.75, 0.76, 0.75, 0.75, 
    0.76, 0.75, 0.78, 0.78, 0.8, 0.77, 0.78, 0.8, 0.8, 0.82, 0.82, 0.8, 0.79, 
    0.82, 0.81, 0.81, 0.81, 0.81, 0.8, 0.81, 0.81, 0.81, 0.81, 0.81, 0.83, 
    0.82, 0.83, 0.84, 0.84, 0.84, 0.84, 0.83, 0.82, 0.77, 0.74, 0.78, 0.82, 
    0.84, 0.85, 0.87, 0.88, 0.89, 0.9, 0.91, 0.91, 0.93, 0.94, 0.95, 0.96, 
    0.96, 0.95, 0.95, 0.96, 0.98, 0.98, 0.97, 0.97, 0.96, 0.96, 0.96, 0.94, 
    0.93, 0.92, 0.92, 0.91, 0.93, 0.97, 0.96, 0.95, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.96, 0.96, 0.94, 0.91, 0.9, 0.9, 0.9, 0.92, 0.95, 0.94, 
    0.91, 0.88, 0.84, 0.83, 0.8, 0.81, 0.82, 0.82, 0.82, 0.81, 0.79, 0.77, 
    0.81, 0.78, 0.77, 0.76, 0.8, 0.82, 0.83, 0.83, 0.82, 0.82, 0.8, 0.81, 
    0.81, 0.8, 0.76, 0.74, 0.77, 0.82, 0.83, 0.83, 0.8, 0.69, 0.7, 0.81, 
    0.85, 0.83, 0.81, 0.81, 0.82, 0.81, 0.8, 0.78, 0.78, 0.8, 0.89, 0.9, 
    0.89, 0.9, 0.9, 0.9, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 0.9, 
    0.9, 0.89, 0.89, 0.9, 0.9, 0.9, 0.92, 0.91, 0.92, 0.92, 0.93, 0.94, 0.95, 
    0.95, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.99, 
    0.99, 0.99, 1, 0.99, 1, 0.99, 1, 1, 0.99, 0.97, 0.94, 0.97, 0.94, 0.92, 
    0.9, 0.91, 0.92, 0.91, 0.9, 0.89, 0.89, 0.89, 0.87, 0.88, 0.9, 0.88, 
    0.89, 0.88, 0.87, 0.87, 0.87, 0.88, 0.87, 0.86, 0.86, 0.86, 0.86, 0.85, 
    0.85, 0.86, 0.85, 0.86, 0.86, 0.85, 0.85, 0.84, 0.83, 0.82, 0.82, 0.8, 
    0.81, 0.68, 0.63, 0.72, 0.85, 0.85, 0.88, 0.87, 0.86, 0.85, 0.87, 0.88, 
    0.87, 0.87, 0.88, 0.87, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.87, 
    0.87, 0.87, 0.89, 0.91, 0.9, 0.91, 0.92, 0.93, 0.93, 0.9, 0.91, 0.92, 
    0.92, 0.93, 0.92, 0.92, 0.92, 0.93, 0.94, 0.95, 0.92, 0.94, 0.94, 0.91, 
    0.92, 0.91, 0.88, 0.89, 0.88, 0.83, 0.6, 0.59, 0.58, 0.61, 0.73, 0.78, 
    0.81, 0.78, 0.82, 0.83, 0.81, 0.7, 0.68, 0.69, 0.69, 0.68, 0.66, 0.64, 
    0.66, 0.65, 0.78, 0.78, 0.8, 0.82, 0.83, 0.81, 0.82, 0.82, 0.83, 0.82, 
    0.82, 0.82, 0.82, 0.82, 0.83, 0.84, 0.84, 0.83, 0.84, 0.85, 0.85, 0.84, 
    0.83, 0.83, 0.84, 0.83, 0.83, 0.81, 0.81, 0.78, 0.77, 0.77, 0.78, 0.74, 
    0.72, 0.79, 0.79, 0.86, 0.86, 0.86, 0.85, 0.85, 0.85, 0.83, 0.85, 0.85, 
    0.83, 0.85, 0.84, 0.84, 0.83, 0.84, 0.86, 0.87, 0.87, 0.87, 0.86, 0.86, 
    0.85, 0.86, 0.84, 0.87, 0.79, 0.87, 0.87, 0.88, 0.87, 0.87, 0.88, 0.87, 
    0.87, 0.87, 0.86, 0.85, 0.86, 0.86, 0.86, 0.85, 0.84, 0.85, 0.86, 0.87, 
    0.86, 0.86, 0.85, 0.85, 0.85, 0.84, 0.85, 0.86, 0.87, 0.89, 0.9, 0.89, 
    0.9, 0.9, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 0.92, 
    0.92, 0.92, 0.91, 0.92, 0.92, 0.92, 0.91, 0.9, 0.9, 0.89, 0.89, 0.88, 
    0.87, 0.85, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 0.82, 0.82, 
    0.83, 0.83, 0.82, 0.82, 0.8, 0.81, 0.78, 0.79, 0.81, 0.8, 0.79, 0.82, 
    0.85, 0.86, 0.86, 0.87, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 0.89, 0.89, 0.89, 
    0.88, 0.88, 0.85, 0.83, 0.83, 0.84, 0.83, 0.77, 0.81, 0.83, 0.82, 0.85, 
    0.82, 0.8, 0.79, 0.8, 0.79, 0.78, 0.79, 0.82, 0.83, 0.85, 0.82, 0.76, 
    0.77, 0.79, 0.79, 0.81, 0.76, 0.73, 0.72, 0.74, 0.72, 0.76, 0.77, 0.79, 
    0.81, 0.81, 0.83, 0.84, 0.8, 0.86, 0.84, 0.86, 0.86, 0.86, 0.88, 0.86, 
    0.87, 0.86, 0.84, 0.87, 0.87, 0.86, 0.83, 0.84, 0.81, 0.82, 0.86, 0.89, 
    0.89, 0.9, 0.89, 0.91, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 
    0.94, 0.94, 0.95, 0.93, 0.92, 0.91, 0.92, 0.9, 0.95, 0.94, 0.99, 0.93, 
    0.91, 0.96, 0.96, 0.95, 0.9, 0.9, 0.87, 0.85, 0.88, 0.88, 0.87, 0.88, 
    0.89, 0.87, 0.85, 0.86, 0.88, 0.92, 0.9, 0.91, 0.91, 0.91, 0.86, 0.87, 
    0.91, 0.91, 0.87, 0.84, 0.85, 0.87, 0.86, 0.83, 0.83, 0.8, 0.8, 0.85, 
    0.89, 0.93, 0.85, 0.78, 0.76, 0.78, 0.76, 0.76, 0.92, 0.86, 0.78, 0.77, 
    0.74, 0.76, 0.78, 0.76, 0.82, 0.84, 0.89, 0.94, 0.96, 0.94, 0.9, 0.91, 
    0.9, 0.81, 0.8, 0.8, 0.82, 0.82, 0.82, 0.8, 0.76, 0.74, 0.8, 0.82, 0.81, 
    0.82, 0.87, 0.88, 0.85, 0.84, 0.85, 0.85, 0.86, 0.88, 0.88, 0.89, 0.91, 
    0.9, 0.92, 0.91, 0.86, 0.89, 0.86, 0.87, 0.86, 0.82, 0.76, 0.76, 0.82, 
    0.78, 0.77, 0.79, 0.79, 0.84, 0.86, 0.86, 0.91, 0.81, 0.84, 0.79, 0.82, 
    0.82, 0.82, 0.82, 0.81, 0.84, 0.82, 0.85, 0.9, 0.91, 0.92, 0.82, 0.77, 
    0.84, 0.75, 0.86, 0.83, 0.83, 0.82, 0.86, 0.84, 0.85, 0.87, 0.88, 0.88, 
    0.87, 0.88, 0.89, 0.88, 0.89, 0.9, 0.9, 0.91, 0.89, 0.9, 0.89, 0.92, 0.9, 
    0.83, 0.89, 0.89, 0.9, 0.86, 0.83, 0.77, 0.79, 0.93, 0.73, 0.8, 0.86, 
    0.84, 0.84, 0.85, 0.89, 0.86, 0.87, 0.86, 0.86, 0.86, 0.87, 0.87, 0.88, 
    0.89, 0.89, 0.9, 0.9, 0.88, 0.87, 0.88, 0.88, 0.88, 0.88, 0.87, 0.87, 
    0.87, 0.86, 0.86, 0.86, 0.85, 0.85, 0.86, 0.86, 0.85, 0.84, 0.84, 0.83, 
    0.83, 0.83, 0.84, 0.83, 0.82, 0.82, 0.83, 0.82, 0.83, 0.82, 0.82, 0.81, 
    0.8, 0.81, 0.82, 0.81, 0.8, 0.81, 0.8, 0.8, 0.81, 0.8, 0.81, 0.81, 0.8, 
    0.81, 0.81, 0.8, 0.81, 0.8, 0.79, 0.84, 0.83, 0.83, 0.82, 0.82, 0.82, 
    0.83, 0.82, 0.82, 0.83, 0.83, 0.82, 0.82, 0.82, 0.81, 0.82, 0.82, 0.83, 
    0.82, 0.82, 0.82, 0.82, 0.82, 0.83, 0.83, 0.81, 0.8, 0.79, 0.8, 0.8, 
    0.78, 0.79, 0.78, 0.8, 0.8, 0.79, 0.8, 0.8, 0.8, 0.79, 0.79, 0.79, 0.79, 
    0.78, 0.78, 0.78, 0.78, 0.8, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 
    0.78, 0.78, 0.78, 0.77, 0.77, 0.76, 0.77, 0.78, 0.77, 0.78, 0.77, 0.77, 
    0.76, 0.77, 0.76, 0.77, 0.77, 0.77, 0.77, 0.77, 0.77, 0.77, 0.76, 0.78, 
    0.79, 0.77, 0.77, 0.77, 0.78, 0.77, 0.78, 0.78, 0.78, 0.78, 0.79, 0.79, 
    0.79, 0.79, 0.8, 0.8, 0.8, 0.79, 0.79, 0.79, 0.79, 0.8, 0.8, 0.8, 0.79, 
    0.78, 0.79, 0.78, 0.79, 0.77, 0.78, 0.78, 0.78, 0.78, 0.77, 0.78, 0.76, 
    0.75, 0.75, 0.77, 0.78, 0.78, 0.78, 0.78, 0.77, 0.77, 0.76, 0.77, 0.77, 
    0.77, 0.77, 0.76, 0.77, 0.78, 0.78, 0.78, 0.79, 0.77, 0.76, 0.75, 0.75, 
    0.76, 0.76, 0.77, 0.76, 0.76, 0.75, 0.77, 0.77, 0.77, 0.76, 0.77, 0.76, 
    0.78, 0.8, 0.8, 0.8, 0.79, 0.8, 0.78, 0.78, 0.79, 0.8, 0.79, 0.79, 0.79, 
    0.79, 0.79, 0.79, 0.78, 0.77, 0.78, 0.79, 0.77, 0.77, 0.73, 0.75, 0.77, 
    0.78, 0.78, 0.78, 0.78, 0.78, 0.77, 0.77, 0.75, 0.73, 0.72, 0.71, 0.71, 
    0.78, 0.8, 0.79, 0.8, 0.79, 0.79, 0.79, 0.8, 0.8, 0.8, 0.81, 0.82, 0.82, 
    0.81, 0.83, 0.83, 0.84, 0.86, 0.88, 0.9, 0.9, 0.92, 0.92, 0.91, 0.92, 
    0.93, 0.94, 0.93, 0.93, 0.94, 0.93, 0.94, 0.95, 0.94, 0.93, 0.92, 0.92, 
    0.91, 0.9, 0.9, 0.91, 0.9, 0.91, 0.91, 0.92, 0.93, 0.92, 0.93, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.94, 0.93, 0.94, 0.94, 
    0.93, 0.94, 0.94, 0.93, 0.94, 0.94, 0.93, 0.93, 0.93, 0.94, 0.95, 0.94, 
    0.94, 0.93, 0.93, 0.92, 0.93, 0.92, 0.92, 0.92, 0.91, 0.92, 0.92, 0.92, 
    0.93, 0.92, 0.91, 0.9, 0.9, 0.89, 0.89, 0.9, 0.9, 0.9, 0.9, 0.88, 0.87, 
    0.86, 0.85, 0.85, 0.87, 0.87, 0.89, 0.87, 0.86, 0.85, 0.85, 0.86, 0.86, 
    0.81, 0.85, 0.84, 0.84, 0.84, 0.83, 0.85, 0.87, 0.85, 0.84, 0.83, 0.86, 
    0.85, 0.87, 0.87, 0.88, 0.89, 0.89, 0.87, 0.85, 0.84, 0.83, 0.84, 0.84, 
    0.85, 0.87, 0.88, 0.86, 0.87, 0.89, 0.91, 0.92, 0.92, 0.93, 0.93, 0.93, 
    0.92, 0.86, 0.86, 0.85, 0.88, 0.87, 0.89, 0.82, 0.86, 0.83, 0.84, 0.85, 
    0.85, 0.84, 0.84, 0.85, 0.85, 0.79, 0.76, 0.81, 0.85, 0.86, 0.84, 0.83, 
    0.84, 0.84, 0.83, 0.85, 0.85, 0.87, 0.9, 0.9, 0.92, 0.92, 0.93, 0.93, 
    0.92, 0.92, 0.94, 0.93, 0.94, 0.93, 0.93, 0.93, 0.93, 0.92, 0.91, 0.92, 
    0.91, 0.91, 0.91, 0.91, 0.9, 0.9, 0.9, 0.87, 0.85, 0.84, 0.85, 0.84, 0.9, 
    0.9, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.98, 
    0.97, 0.97, 0.97, 0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.96, 0.94, 0.96, 
    0.93, 0.9, 0.88, 0.89, 0.89, 0.87, 0.88, 0.89, 0.91, 0.9, 0.91, 0.91, 
    0.9, 0.92, 0.94, 0.93, 0.93, 0.94, 0.93, 0.93, 0.93, 0.94, 0.93, 0.92, 
    0.91, 0.91, 0.91, 0.9, 0.91, 0.9, 0.89, 0.88, 0.85, 0.83, 0.91, 0.92, 
    0.88, 0.89, 0.86, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.83, 0.85, 0.84, 
    0.81, 0.76, 0.8, 0.82, 0.81, 0.81, 0.8, 0.78, 0.75, 0.73, 0.72, 0.83, 
    0.87, 0.87, 0.86, 0.85, 0.84, 0.84, 0.83, 0.86, 0.83, 0.83, 0.83, 0.85, 
    0.84, 0.83, 0.85, 0.84, 0.85, 0.86, 0.89, 0.91, 0.9, 0.88, 0.92, 0.93, 
    0.92, 0.92, 0.92, 0.94, 0.94, 0.92, 0.88, 0.86, 0.77, 0.78, 0.89, 0.82, 
    0.88, 0.86, 0.84, 0.83, 0.83, 0.85, 0.82, 0.87, 0.83, 0.88, 0.85, 0.84, 
    0.86, 0.85, 0.87, 0.85, 0.81, 0.83, 0.86, 0.86, 0.57, 0.51, 0.64, 0.63, 
    0.61, 0.65, 0.75, 0.75, 0.72, 0.72, 0.75, 0.72, 0.72, 0.7, 0.68, 0.68, 
    0.7, 0.7, 0.7, 0.71, 0.75, 0.73, 0.81, 0.82, 0.76, 0.81, 0.75, 0.79, 
    0.75, 0.77, 0.83, 0.78, 0.84, 0.9, 0.87, 0.84, 0.89, 0.86, 0.84, 0.85, 
    0.84, 0.85, 0.86, 0.86, 0.86, 0.85, 0.82, 0.82, 0.84, 0.78, 0.76, 0.73, 
    0.7, 0.74, 0.77, 0.73, 0.77, 0.72, 0.72, 0.76, 0.73, 0.72, 0.76, 0.69, 
    0.64, 0.7, 0.7, 0.71, 0.69, 0.7, 0.66, 0.69, 0.61, 0.63, 0.66, 0.59, 
    0.75, 0.77, 0.77, 0.75, 0.75, 0.74, 0.75, 0.75, 0.76, 0.76, 0.74, 0.75, 
    0.76, 0.78, 0.78, 0.78, 0.75, 0.73, 0.7, 0.78, 0.76, 0.8, 0.83, 0.79, 
    0.82, 0.8, 0.81, 0.74, 0.79, 0.8, 0.81, 0.82, 0.83, 0.87, 0.83, 0.83, 
    0.83, 0.85, 0.82, 0.88, 0.83, 0.87, 0.85, 0.83, 0.8, 0.78, 0.79, 0.78, 
    0.74, 0.74, 0.69, 0.69, 0.65, 0.74, 0.6, 0.6, 0.8, 0.8, 0.79, 0.81, 0.82, 
    0.82, 0.81, 0.81, 0.82, 0.83, 0.83, 0.85, 0.83, 0.83, 0.83, 0.83, 0.85, 
    0.84, 0.84, 0.84, 0.83, 0.87, 0.87, 0.85, 0.87, 0.82, 0.85, 0.81, 0.82, 
    0.81, 0.81, 0.81, 0.83, 0.8, 0.78, 0.74, 0.74, 0.72, 0.64, 0.69, 0.57, 
    0.68, 0.64, 0.58, 0.58, 0.59, 0.6, 0.59, 0.58, 0.66, 0.71, 0.78, 0.8, 
    0.8, 0.81, 0.83, 0.85, 0.88, 0.88, 0.9, 0.9, 0.92, 0.92, 0.92, 0.93, 
    0.92, 0.91, 0.92, 0.93, 0.95, 0.96, 0.96, 0.98, 0.99, 0.98, 0.97, 0.95, 
    0.94, 0.93, 0.94, 0.93, 0.94, 0.95, 0.95, 0.93, 0.91, 0.92, 0.91, 0.91, 
    0.9, 0.9, 0.9, 0.89, 0.89, 0.9, 0.91, 0.89, 0.88, 0.88, 0.88, 0.88, 0.87, 
    0.87, 0.89, 0.94, 0.95, 0.89, 0.89, 0.93, 0.94, 0.95, 0.95, 0.94, 0.96, 
    0.93, 0.9, 0.9, 0.91, 0.88, 0.89, 0.89, 0.85, 0.81, 0.75, 0.74, 0.78, 
    0.72, 0.75, 0.78, 0.77, 0.86, 0.86, 0.72, 0.68, 0.67, 0.65, 0.63, 0.66, 
    0.59, 0.58, 0.63, 0.62, 0.55, 0.55, 0.56, 0.56, 0.55, 0.59, 0.59, 0.6, 
    0.67, 0.6, 0.61, 0.73, 0.74, 0.71, 0.73, 0.72, 0.75, 0.73, 0.7, 0.6, 
    0.67, 0.75, 0.67, 0.67, 0.68, 0.68, 0.69, 0.76, 0.74, 0.74, 0.79, 0.78, 
    0.8, 0.81, 0.81, 0.8, 0.8, 0.8, 0.79, 0.79, 0.79, 0.78, 0.75, 0.65, 0.68, 
    0.67, 0.65, 0.63, 0.67, 0.7, 0.7, 0.71, 0.73, 0.73, 0.73, 0.71, 0.7, 
    0.69, 0.7, 0.69, 0.7, 0.72, 0.75, 0.77, 0.66, 0.67, 0.66, 0.66, 0.67, 
    0.69, 0.72, 0.68, 0.7, 0.78, 0.77, 0.77, 0.78, 0.77, 0.78, 0.78, 0.79, 
    0.78, 0.78, 0.78, 0.77, 0.75, 0.71, 0.71, 0.72, 0.71, 0.71, 0.72, 0.71, 
    0.68, 0.69, 0.69, 0.73, 0.73, 0.71, 0.68, 0.7, 0.73, 0.77, 0.72, 0.77, 
    0.79, 0.77, 0.78, 0.76, 0.76, 0.76, 0.77, 0.77, 0.76, 0.75, 0.76, 0.76, 
    0.75, 0.71, 0.65, 0.63, 0.64, 0.62, 0.66, 0.71, 0.66, 0.72, 0.64, 0.65, 
    0.78, 0.61, 0.66, 0.65, 0.65, 0.66, 0.67, 0.68, 0.74, 0.66, 0.59, 0.66, 
    0.62, 0.58, 0.58, 0.69, 0.54, 0.7, 0.76, 0.8, 0.76, 0.81, 0.81, 0.77, 
    0.78, 0.74, 0.78, 0.78, 0.76, 0.72, 0.74, 0.72, 0.66, 0.69, 0.69, 0.7, 
    0.76, 0.76, 0.77, 0.76, 0.74, 0.76, 0.77, 0.75, 0.74, 0.74, 0.75, 0.74, 
    0.72, 0.76, 0.76, 0.72, 0.76, 0.72, 0.72, 0.77, 0.75, 0.71, 0.67, 0.71, 
    0.73, 0.73, 0.73, 0.73, 0.73, 0.7, 0.72, 0.74, 0.76, 0.73, 0.74, 0.71, 
    0.71, 0.71, 0.77, 0.79, 0.75, 0.7, 0.71, 0.73, 0.75, 0.71, 0.76, 0.75, 
    0.73, 0.72, 0.72, 0.72, 0.73, 0.73, 0.66, 0.69, 0.72, 0.75, 0.71, 0.68, 
    0.84, 0.83, 0.82, 0.83, 0.84, 0.85, 0.86, 0.85, 0.87, 0.86, 0.85, 0.83, 
    0.82, 0.8, 0.83, 0.84, 0.83, 0.82, 0.8, 0.8, 0.81, 0.85, 0.85, 0.84, 
    0.85, 0.89, 0.88, 0.93, 0.94, 0.94, 0.94, 0.93, 0.92, 0.93, 0.93, 0.95, 
    0.93, 0.95, 0.96, 0.97, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 
    0.98, 0.98, 0.97, 0.95, 0.94, 0.92, 0.91, 0.9, 0.9, 0.89, 0.92, 0.91, 
    0.9, 0.9, 0.89, 0.89, 0.89, 0.9, 0.89, 0.88, 0.89, 0.88, 0.87, 0.87, 
    0.87, 0.86, 0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 0.86, 0.86, 0.87, 0.87, 
    0.87, 0.88, 0.88, 0.89, 0.89, 0.89, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 
    0.89, 0.89, 0.9, 0.89, 0.9, 0.9, 0.89, 0.88, 0.87, 0.87, 0.87, 0.87, 
    0.87, 0.87, 0.88, 0.87, 0.86, 0.86, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 
    0.84, 0.84, 0.84, 0.84, 0.83, 0.84, 0.83, 0.84, 0.85, 0.85, 0.84, 0.83, 
    0.84, 0.84, 0.85, 0.84, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 
    0.84, 0.84, 0.83, 0.83, 0.83, 0.84, 0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 
    0.83, 0.83, 0.83, 0.83, 0.82, 0.82, 0.83, 0.83, 0.82, 0.82, 0.83, 0.84, 
    0.83, 0.84, 0.84, 0.82, 0.82, 0.82, 0.83, 0.83, 0.82, 0.81, 0.81, 0.82, 
    0.82, 0.81, 0.81, 0.81, 0.8, 0.8, 0.8, 0.8, 0.8, 0.79, 0.78, 0.79, 0.8, 
    0.8, 0.8, 0.8, 0.78, 0.79, 0.79, 0.8, 0.79, 0.79, 0.8, 0.79, 0.79, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.81, 0.81, 0.81, 0.81, 0.82, 0.82, 0.83, 
    0.83, 0.83, 0.84, 0.84, 0.84, 0.83, 0.84, 0.84, 0.85, 0.83, 0.83, 0.84, 
    0.84, 0.84, 0.84, 0.84, 0.86, 0.84, 0.82, 0.83, 0.82, 0.81, 0.81, 0.8, 
    0.8, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.8, 
    0.79, 0.79, 0.79, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.81, 0.81, 0.81, 
    0.81, 0.81, 0.81, 0.82, 0.8, 0.79, 0.79, 0.78, 0.78, 0.78, 0.78, 0.78, 
    0.78, 0.79, 0.8, 0.81, 0.8, 0.81, 0.81, 0.81, 0.82, 0.82, 0.83, 0.83, 
    0.83, 0.84, 0.84, 0.85, 0.85, 0.86, 0.86, 0.88, 0.89, 0.9, 0.91, 0.91, 
    0.92, 0.93, 0.95, 0.97, 0.97, 0.98, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.96, 0.96, 
    0.95, 0.96, 0.96, 0.95, 0.94, 0.97, 0.97, 0.94, 0.94, 0.95, 0.97, 0.96, 
    0.97, 0.97, 0.97, 0.96, 0.97, 0.95, 0.96, 0.95, 0.93, 0.91, 0.91, 0.9, 
    0.9, 0.88, 0.87, 0.87, 0.85, 0.85, 0.84, 0.83, 0.83, 0.84, 0.85, 0.84, 
    0.84, 0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 0.82, 0.82, 0.83, 0.84, 0.83, 
    0.81, 0.81, 0.8, 0.79, 0.78, 0.77, 0.79, 0.83, 0.86, 0.86, 0.86, 0.86, 
    0.87, 0.87, 0.87, 0.86, 0.86, 0.86, 0.85, 0.85, 0.83, 0.83, 0.84, 0.82, 
    0.83, 0.83, 0.81, 0.83, 0.83, 0.79, 0.83, 0.82, 0.82, 0.82, 0.82, 0.82, 
    0.82, 0.83, 0.83, 0.84, 0.84, 0.83, 0.83, 0.84, 0.84, 0.82, 0.81, 0.83, 
    0.82, 0.79, 0.82, 0.81, 0.79, 0.78, 0.77, 0.79, 0.77, 0.78, 0.77, 0.79, 
    0.77, 0.77, 0.78, 0.8, 0.78, 0.82, 0.79, 0.79, 0.79, 0.76, 0.75, 0.81, 
    0.78, 0.79, 0.75, 0.81, 0.81, 0.81, 0.81, 0.81, 0.8, 0.8, 0.81, 0.8, 
    0.82, 0.84, 0.8, 0.82, 0.82, 0.83, 0.81, 0.83, 0.83, 0.81, 0.81, 0.82, 
    0.82, 0.81, 0.81, 0.82, 0.78, 0.79, 0.78, 0.79, 0.79, 0.79, 0.76, 0.74, 
    0.76, 0.78, 0.81, 0.79, 0.79, 0.79, 0.79, 0.8, 0.81, 0.78, 0.81, 0.69, 
    0.69, 0.72, 0.68, 0.71, 0.68, 0.69, 0.68, 0.66, 0.69, 0.8, 0.81, 0.74, 
    0.8, 0.69, 0.85, 0.91, 0.88, 0.87, 0.88, 0.87, 0.88, 0.89, 0.89, 0.9, 
    0.88, 0.89, 0.88, 0.88, 0.89, 0.88, 0.88, 0.88, 0.88, 0.89, 0.89, 0.88, 
    0.88, 0.87, 0.86, 0.86, 0.85, 0.83, 0.82, 0.82, 0.83, 0.89, 0.81, 0.84, 
    0.82, 0.82, 0.82, 0.85, 0.86, 0.87, 0.88, 0.87, 0.89, 0.88, 0.87, 0.85, 
    0.86, 0.86, 0.84, 0.85, 0.83, 0.83, 0.84, 0.81, 0.82, 0.83, 0.83, 0.83, 
    0.84, 0.83, 0.83, 0.81, 0.82, 0.83, 0.86, 0.85, 0.85, 0.84, 0.85, 0.84, 
    0.8, 0.72, 0.62, 0.77, 0.82, 0.88, 0.87, 0.87, 0.88, 0.86, 0.84, 0.84, 
    0.81, 0.77, 0.69, 0.77, 0.69, 0.72, 0.74, 0.62, 0.62, 0.71, 0.79, 0.82, 
    0.82, 0.87, 0.85, 0.83, 0.82, 0.82, 0.85, 0.81, 0.83, 0.84, 0.83, 0.85, 
    0.85, 0.86, 0.84, 0.83, 0.83, 0.82, 0.83, 0.83, 0.83, 0.85, 0.84, 0.86, 
    0.85, 0.83, 0.72, 0.69, 0.69, 0.73, 0.81, 0.8, 0.81, 0.82, 0.8, 0.82, 
    0.8, 0.83, 0.82, 0.83, 0.84, 0.85, 0.85, 0.86, 0.86, 0.85, 0.86, 0.87, 
    0.86, 0.86, 0.87, 0.87, 0.89, 0.89, 0.9, 0.9, 0.91, 0.91, 0.91, 0.92, 
    0.92, 0.92, 0.93, 0.93, 0.94, 0.94, 0.95, 0.95, 0.96, 0.97, 0.98, 0.98, 
    0.99, 0.98, 0.98, 0.99, 0.99, 0.97, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.98, 0.97, 0.97, 0.96, 0.96, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.95, 0.94, 0.94, 0.91, 0.91, 0.92, 0.94, 0.95, 0.93, 0.93, 0.93, 0.93, 
    0.92, 0.92, 0.91, 0.91, 0.91, 0.9, 0.89, 0.88, 0.87, 0.87, 0.89, 0.88, 
    0.87, 0.89, 0.92, 0.92, 0.93, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.95, 
    0.95, 0.95, 0.95, 0.95, 0.95, 0.94, 0.95, 0.95, 0.95, 0.96, 0.94, 0.94, 
    0.95, 0.93, 0.93, 0.93, 0.94, 0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.95, 
    0.96, 0.95, 0.94, 0.92, 0.92, 0.92, 0.92, 0.91, 0.91, 0.91, 0.91, 0.91, 
    0.91, 0.92, 0.94, 0.94, 0.95, 0.96, 0.97, 0.97, 0.96, 0.94, 0.95, 0.95, 
    0.95, 0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.91, 0.91, 
    0.92, 0.92, 0.93, 0.94, 0.94, 0.95, 0.95, 0.95, 0.97, 0.97, 0.94, 0.94, 
    0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.93, 0.94, 0.95, 0.95, 0.94, 0.95, 0.93, 0.92, 0.92, 
    0.92, 0.91, 0.91, 0.87, 0.87, 0.85, 0.83, 0.85, 0.86, 0.82, 0.83, 0.81, 
    0.81, 0.79, 0.77, 0.76, 0.76, 0.76, 0.75, 0.75, 0.76, 0.77, 0.77, 0.78, 
    0.78, 0.76, 0.76, 0.76, 0.76, 0.75, 0.75, 0.74, 0.74, 0.76, 0.76, 0.76, 
    0.77, 0.77, 0.76, 0.76, 0.75, 0.76, 0.79, 0.82, 0.87, 0.85, 0.87, 0.87, 
    0.86, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 0.85, 0.83, 0.82, 
    0.81, 0.8, 0.8, 0.79, 0.79, 0.8, 0.82, 0.83, 0.84, 0.82, 0.82, 0.83, 
    0.84, 0.83, 0.83, 0.84, 0.83, 0.83, 0.84, 0.83, 0.83, 0.79, 0.79, 0.79, 
    0.79, 0.81, 0.8, 0.79, 0.8, 0.84, 0.85, 0.86, 0.78, 0.79, 0.84, 0.85, 
    0.86, 0.86, 0.86, 0.87, 0.9, 0.92, 0.93, 0.96, 0.98, 0.96, 0.95, 0.93, 
    0.91, 0.86, 0.81, 0.81, 0.84, 0.82, 0.83, 0.82, 0.85, 0.9, 0.96, 0.98, 
    0.99, 0.98, 0.87, 0.85, 0.86, 0.89, 0.87, 0.88, 0.83, 0.86, 0.8, 0.8, 
    0.81, 0.81, 0.8, 0.8, 0.79, 0.79, 0.79, 0.79, 0.8, 0.79, 0.79, 0.79, 
    0.78, 0.77, 0.76, 0.75, 0.77, 0.75, 0.75, 0.76, 0.77, 0.74, 0.75, 0.75, 
    0.76, 0.8, 0.81, 0.81, 0.81, 0.85, 0.85, 0.87, 0.85, 0.85, 0.86, 0.85, 
    0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.85, 0.85, 0.85, 0.83, 0.83, 
    0.82, 0.79, 0.81, 0.8, 0.8, 0.81, 0.81, 0.8, 0.78, 0.78, 0.79, 0.79, 0.8, 
    0.8, 0.81, 0.82, 0.8, 0.8, 0.8, 0.8, 0.79, 0.79, 0.78, 0.79, 0.79, 0.8, 
    0.8, 0.79, 0.8, 0.79, 0.78, 0.78, 0.78, 0.77, 0.76, 0.76, 0.77, 0.78, 
    0.78, 0.79, 0.78, 0.78, 0.78, 0.78, 0.78, 0.78, 0.78, 0.78, 0.79, 0.8, 
    0.79, 0.79, 0.81, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 
    0.82, 0.82, 0.82, 0.81, 0.82, 0.8, 0.8, 0.79, 0.79, 0.79, 0.8, 0.79, 
    0.79, 0.8, 0.8, 0.82, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.83, 0.83, 
    0.83, 0.84, 0.82, 0.84, 0.78, 0.74, 0.83, 0.84, 0.84, 0.84, 0.83, 0.84, 
    0.73, 0.79, 0.76, 0.74, 0.77, 0.86, 0.7, 0.83, 0.82, 0.72, 0.72, 0.73, 
    0.74, 0.8, 0.78, 0.8, 0.8, 0.77, 0.79, 0.81, 0.8, 0.8, 0.79, 0.79, 0.81, 
    0.82, 0.83, 0.82, 0.84, 0.83, 0.83, 0.83, 0.82, 0.81, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.77, 0.78, 0.78, 0.77, 0.78, 0.77, 0.78, 0.78, 0.79, 
    0.79, 0.79, 0.8, 0.79, 0.78, 0.78, 0.77, 0.8, 0.8, 0.8, 0.81, 0.79, 0.79, 
    0.79, 0.79, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.84, 0.85, 0.85, 0.85, 
    0.85, 0.85, 0.86, 0.86, 0.86, 0.87, 0.88, 0.89, 0.9, 0.91, 0.92, 0.92, 
    0.93, 0.94, 0.94, 0.94, 0.94, 0.95, 0.96, 0.96, 0.97, 0.96, 0.95, 0.96, 
    0.96, 0.94, 0.94, 0.95, 0.93, 0.94, 0.95, 0.94, 0.92, 0.9, 0.91, 0.92, 
    0.91, 0.9, 0.9, 0.92, 0.92, 0.95, 0.95, 0.95, 0.97, 0.98, 0.97, 0.93, 
    0.94, 0.92, 0.89, 0.84, 0.86, 0.85, 0.83, 0.83, 0.91, 0.89, 0.91, 0.91, 
    0.88, 0.85, 0.87, 0.89, 0.9, 0.9, 0.88, 0.89, 0.88, 0.87, 0.87, 0.87, 
    0.87, 0.87, 0.88, 0.87, 0.85, 0.84, 0.83, 0.83, 0.81, 0.75, 0.76, 0.75, 
    0.73, 0.69, 0.82, 0.81, 0.8, 0.8, 0.81, 0.81, 0.82, 0.83, 0.84, 0.82, 
    0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.85, 0.85, 0.84, 0.83, 0.84, 0.82, 
    0.82, 0.8, 0.8, 0.8, 0.78, 0.78, 0.78, 0.79, 0.81, 0.83, 0.83, 0.85, 
    0.81, 0.84, 0.85, 0.84, 0.85, 0.86, 0.8, 0.8, 0.86, 0.85, 0.83, 0.81, 
    0.81, 0.8, 0.81, 0.82, 0.81, 0.81, 0.8, 0.81, 0.82, 0.8, 0.8, 0.8, 0.8, 
    0.82, 0.8, 0.79, 0.8, 0.83, 0.81, 0.82, 0.83, 0.82, 0.83, 0.82, 0.83, 
    0.85, 0.85, 0.84, 0.84, 0.85, 0.85, 0.85, 0.84, 0.84, 0.85, 0.85, 0.86, 
    0.86, 0.86, 0.87, 0.87, 0.87, 0.86, 0.85, 0.85, 0.86, 0.86, 0.86, 0.85, 
    0.85, 0.83, 0.83, 0.83, 0.81, 0.81, 0.81, 0.81, 0.81, 0.83, 0.81, 0.81, 
    0.81, 0.8, 0.8, 0.8, 0.79, 0.8, 0.8, 0.79, 0.78, 0.77, 0.78, 0.78, 0.76, 
    0.76, 0.76, 0.8, 0.77, 0.77, 0.78, 0.78, 0.79, 0.8, 0.79, 0.73, 0.73, 
    0.74, 0.75, 0.75, 0.76, 0.76, 0.76, 0.73, 0.73, 0.76, 0.73, 0.74, 0.7, 
    0.63, 0.62, 0.63, 0.74, 0.76, 0.79, 0.77, 0.76, 0.7, 0.79, 0.78, 0.74, 
    0.73, 0.77, 0.73, 0.83, 0.84, 0.85, 0.81, 0.8, 0.8, 0.78, 0.79, 0.75, 
    0.72, 0.75, 0.75, 0.76, 0.8, 0.79, 0.65, 0.64, 0.68, 0.69, 0.74, 0.66, 
    0.77, 0.86, 0.85, 0.83, 0.82, 0.84, 0.84, 0.84, 0.87, 0.89, 0.87, 0.86, 
    0.87, 0.89, 0.89, 0.92, 0.9, 0.93, 0.93, 0.91, 0.92, 0.92, 0.93, 0.93, 
    0.92, 0.93, 0.92, 0.93, 0.93, 0.93, 0.92, 0.96, 0.91, 0.91, 0.91, 0.93, 
    0.92, 0.91, 0.9, 0.92, 0.93, 0.93, 0.92, 0.9, 0.91, 0.92, 0.92, 0.91, 
    0.91, 0.9, 0.9, 0.91, 0.89, 0.86, 0.86, 0.81, 0.91, 0.93, 0.91, 0.93, 
    0.94, 0.94, 0.93, 0.93, 0.93, 0.92, 0.91, 0.94, 0.95, 0.94, 0.94, 0.94, 
    0.93, 0.93, 0.93, 0.93, 0.94, 0.93, 0.93, 0.94, 0.94, 0.93, 0.9, 0.9, 
    0.91, 0.85, 0.8, 0.85, 0.88, 0.85, 0.89, 0.89, 0.91, 0.87, 0.88, 0.94, 
    0.93, 0.93, 0.93, 0.92, 0.94, 0.94, 0.89, 0.91, 0.91, 0.91, 0.88, 0.87, 
    0.86, 0.89, 0.89, 0.9, 0.89, 0.84, 0.86, 0.9, 0.94, 0.89, 0.88, 0.87, 
    0.91, 0.92, 0.94, 0.92, 0.92, 0.91, 0.91, 0.92, 0.91, 0.91, 0.91, 0.89, 
    0.91, 0.9, 0.9, 0.92, 0.92, 0.91, 0.9, 0.91, 0.91, 0.9, 0.9, 0.95, 0.94, 
    0.93, 0.92, 0.92, 0.89, 0.88, 0.9, 0.89, 0.9, 0.87, 0.85, 0.85, 0.85, 
    0.85, 0.85, 0.86, 0.88, 0.9, 0.91, 0.89, 0.9, 0.86, 0.85, 0.79, 0.78, 
    0.79, 0.81, 0.8, 0.8, 0.8, 0.8, 0.81, 0.83, 0.81, 0.82, 0.82, 0.83, 0.84, 
    0.85, 0.84, 0.85, 0.8, 0.83, 0.86, 0.87, 0.88, 0.89, 0.88, 0.88, 0.88, 
    0.9, 0.91, 0.92, 0.92, 0.92, 0.91, 0.9, 0.92, 0.95, 0.95, 0.95, 0.94, 
    0.94, 0.94, 0.93, 0.95, 0.94, 0.95, 0.95, 0.96, 0.97, 0.96, 0.97, 0.97, 
    0.97, 0.95, 0.95, 0.94, 0.92, 0.89, 0.89, 0.79, 0.79, 0.81, 0.84, 0.77, 
    0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.94, 0.93, 
    0.93, 0.92, 0.92, 0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 0.97, 0.95, 0.93, 
    0.89, 0.86, 0.81, 0.85, 0.86, 0.86, 0.86, 0.85, 0.86, 0.84, 0.84, 0.82, 
    0.81, 0.79, 0.83, 0.85, 0.83, 0.86, 0.91, 0.85, 0.8, 0.82, 0.91, 0.95, 
    0.95, 0.97, 0.97, 0.98, 0.95, 0.92, 0.89, 0.87, 0.9, 0.9, 0.96, 0.96, 
    0.94, 0.93, 0.93, 0.92, 0.9, 0.89, 0.88, 0.85, 0.81, 0.75, 0.73, 0.66, 
    0.73, 0.67, 0.7, 0.76, 0.75, 0.77, 0.72, 0.76, 0.79, 0.79, 0.78, 0.73, 
    0.77, 0.74, 0.73, 0.67, 0.69, 0.63, 0.63, 0.68, 0.69, 0.8, 0.73, 0.78, 
    0.78, 0.75, 0.73, 0.8, 0.75, 0.81, 0.72, 0.7, 0.71, 0.64, 0.77, 0.77, 
    0.74, 0.74, 0.77, 0.75, 0.77, 0.76, 0.68, 0.74, 0.68, 0.65, 0.74, 0.75, 
    0.68, 0.76, 0.79, 0.85, 0.73, 0.77, 0.78, 0.76, 0.78, 0.77, 0.76, 0.77, 
    0.73, 0.72, 0.67, 0.69, 0.71, 0.72, 0.81, 0.83, 0.84, 0.83, 0.81, 0.83, 
    0.84, 0.84, 0.85, 0.86, 0.86, 0.87, 0.87, 0.89, 0.9, 0.89, 0.89, 0.88, 
    0.87, 0.87, 0.83, 0.85, 0.78, 0.76, 0.69, 0.74, 0.63, 0.79, 0.78, 0.82, 
    0.84, 0.86, 0.87, 0.88, 0.89, 0.89, 0.88, 0.88, 0.87, 0.85, 0.85, 0.86, 
    0.83, 0.84, 0.85, 0.85, 0.85, 0.84, 0.85, 0.9, 0.89, 0.88, 0.86, 0.85, 
    0.84, 0.85, 0.82, 0.82, 0.82, 0.83, 0.86, 0.86, 0.85, 0.86, 0.87, 0.86, 
    0.83, 0.86, 0.86, 0.84, 0.83, 0.84, 0.83, 0.82, 0.85, 0.86, 0.85, 0.85, 
    0.85, 0.88, 0.86, 0.85, 0.83, 0.83, 0.85, 0.84, 0.84, 0.86, 0.85, 0.84, 
    0.85, 0.85, 0.85, 0.85, 0.83, 0.84, 0.86, 0.85, 0.86, 0.86, 0.86, 0.84, 
    0.82, 0.82, 0.83, 0.84, 0.84, 0.84, 0.85, 0.85, 0.84, 0.84, 0.85, 0.87, 
    0.87, 0.88, 0.88, 0.88, 0.87, 0.87, 0.86, 0.85, 0.86, 0.85, 0.83, 0.83, 
    0.84, 0.83, 0.74, 0.77, 0.79, 0.82, 0.78, 0.77, 0.81, 0.8, 0.82, 0.77, 
    0.83, 0.79, 0.77, 0.79, 0.76, 0.72, 0.75, 0.77, 0.82, 0.78, 0.77, 0.71, 
    0.77, 0.77, 0.73, 0.85, 0.81, 0.78, 0.72, 0.74, 0.75, 0.68, 0.78, 0.73, 
    0.75, 0.9, 0.83, 0.84, 0.84, 0.84, 0.85, 0.87, 0.82, 0.84, 0.86, 0.84, 
    0.83, 0.82, 0.81, 0.81, 0.79, 0.8, 0.81, 0.84, 0.86, 0.8, 0.85, 0.82, 
    0.87, 0.79, 0.78, 0.75, 0.75, 0.65, 0.73, 0.71, 0.61, 0.77, 0.67, 0.87, 
    0.93, 0.93, 0.92, 0.92, 0.87, 0.9, 0.88, 0.88, 0.86, 0.83, 0.82, 0.79, 
    0.79, 0.79, 0.75, 0.76, 0.78, 0.78, 0.78, 0.78, 0.75, 0.77, 0.78, 0.75, 
    0.84, 0.85, 0.84, 0.82, 0.74, 0.77, 0.84, 0.83, 0.81, 0.83, 0.82, 0.82, 
    0.79, 0.76, 0.78, 0.8, 0.79, 0.8, 0.78, 0.79, 0.81, 0.82, 0.83, 0.84, 
    0.84, 0.88, 0.88, 0.9, 0.92, 0.92, 0.87, 0.84, 0.79, 0.77, 0.75, 0.78, 
    0.84, 0.82, 0.82, 0.79, 0.78, 0.78, 0.76, 0.79, 0.82, 0.83, 0.84, 0.85, 
    0.87, 0.86, 0.85, 0.87, 0.87, 0.88, 0.9, 0.9, 0.9, 0.89, 0.87, 0.86, 
    0.86, 0.87, 0.87, 0.88, 0.87, 0.88, 0.87, 0.88, 0.88, 0.89, 0.89, 0.89, 
    0.89, 0.89, 0.87, 0.82, 0.81, 0.8, 0.81, 0.82, 0.78, 0.75, 0.7, 0.65, 
    0.71, 0.73, 0.72, 0.7, 0.75, 0.78, 0.79, 0.69, 0.74, 0.76, 0.79, 0.81, 
    0.82, 0.9, 0.87, 0.87, 0.92, 0.9, 0.85, 0.82, 0.83, 0.85, 0.83, 0.82, 
    0.81, 0.83, 0.82, 0.81, 0.77, 0.84, 0.85, 0.86, 0.86, 0.83, 0.81, 0.83, 
    0.84, 0.84, 0.84, 0.83, 0.82, 0.81, 0.78, 0.68, 0.7, 0.7, 0.73, 0.73, 
    0.72, 0.73, 0.73, 0.76, 0.78, 0.75, 0.76, 0.76, 0.75, 0.77, 0.78, 0.77, 
    0.77, 0.76, 0.74, 0.72, 0.69, 0.72, 0.74, 0.75, 0.73, 0.74, 0.8, 0.77, 
    0.75, 0.75, 0.75, 0.77, 0.76, 0.79, 0.79, 0.8, 0.8, 0.79, 0.74, 0.74, 
    0.73, 0.74, 0.7, 0.71, 0.71, 0.72, 0.72, 0.71, 0.69, 0.7, 0.73, 0.7, 
    0.67, 0.73, 0.75, 0.72, 0.74, 0.76, 0.75, 0.77, 0.78, 0.79, 0.78, 0.77, 
    0.77, 0.75, 0.76, 0.78, 0.77, 0.75, 0.79, 0.8, 0.8, 0.78, 0.75, 0.76, 
    0.76, 0.75, 0.76, 0.72, 0.71, 0.79, 0.8, 0.8, 0.83, 0.83, 0.84, 0.85, 
    0.86, 0.86, 0.87, 0.87, 0.86, 0.86, 0.86, 0.86, 0.84, 0.84, 0.82, 0.84, 
    0.85, 0.85, 0.85, 0.85, 0.87, 0.89, 0.9, 0.92, 0.92, 0.92, 0.93, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 
    0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.95, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.97, 0.97, 0.89, 0.87, 0.9, 0.88, 0.86, 0.85, 0.84, 
    0.81, 0.84, 0.84, 0.84, 0.83, 0.85, 0.85, 0.83, 0.85, 0.83, 0.85, 0.86, 
    0.86, 0.87, 0.86, 0.85, 0.86, 0.83, 0.84, 0.79, 0.76, 0.76, 0.75, 0.75, 
    0.74, 0.8, 0.8, 0.79, 0.84, 0.82, 0.83, 0.87, 0.88, 0.86, 0.85, 0.86, 
    0.88, 0.9, 0.9, 0.92, 0.93, 0.94, 0.97, 0.97, 0.97, 0.96, 0.93, 0.93, 
    0.93, 0.94, 0.97, 0.97, 0.96, 0.96, 0.95, 0.97, 0.97, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.98, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.97, 
    0.98, 0.96, 0.95, 0.9, 0.93, 0.91, 0.94, 0.87, 0.9, 0.88, 0.94, 0.92, 
    0.91, 0.93, 0.91, 0.89, 0.9, 0.88, 0.92, 0.92, 0.91, 0.9, 0.9, 0.91, 
    0.93, 0.9, 0.91, 0.89, 0.87, 0.92, 0.89, 0.92, 0.91, 0.92, 0.91, 0.94, 
    0.92, 0.9, 0.96, 0.92, 0.92, 0.95, 0.95, 0.96, 0.92, 0.94, 0.97, 0.96, 
    0.94, 0.94, 0.95, 0.97, 0.97, 0.97, 0.94, 0.93, 0.93, 0.93, 0.92, 0.92, 
    0.91, 0.9, 0.9, 0.88, 0.87, 0.86, 0.85, 0.83, 0.83, 0.83, 0.83, 0.84, 
    0.82, 0.83, 0.86, 0.87, 0.86, 0.85, 0.87, 0.86, 0.87, 0.88, 0.89, 0.9, 
    0.9, 0.9, 0.87, 0.81, 0.79, 0.8, 0.81, 0.81, 0.83, 0.84, 0.85, 0.86, 
    0.91, 0.93, 0.94, 0.93, 0.93, 0.93, 0.94, 0.95, 0.93, 0.95, 0.93, 0.88, 
    0.87, 0.9, 0.91, 0.95, 0.9, 0.91, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.95, 0.95, 0.94, 0.91, 0.88, 0.85, 0.82, 0.9, 0.87, 0.88, 0.88, 0.9, 
    0.92, 0.93, 0.9, 0.9, 0.82, 0.82, 0.94, 0.85, 0.88, 0.84, 0.85, 0.84, 
    0.82, 0.84, 0.84, 0.87, 0.86, 0.88, 0.92, 0.92, 0.85, 0.83, 0.78, 0.82, 
    0.79, 0.84, 0.8, 0.87, 0.93, 0.91, 0.91, 0.91, 0.91, 0.88, 0.9, 0.9, 
    0.91, 0.93, 0.92, 0.91, 0.89, 0.87, 0.81, 0.78, 0.75, 0.77, 0.69, 0.74, 
    0.78, 0.67, 0.62, 0.78, 0.84, 0.86, 0.87, 0.91, 0.94, 0.92, 0.92, 0.93, 
    0.93, 0.94, 0.93, 0.92, 0.93, 0.92, 0.92, 0.86, 0.81, 0.83, 0.87, 0.9, 
    0.91, 0.88, 0.83, 0.86, 0.88, 0.85, 0.81, 0.85, 0.81, 0.83, 0.84, 0.84, 
    0.82, 0.83, 0.81, 0.79, 0.76, 0.78, 0.79, 0.8, 0.81, 0.82, 0.85, 0.86, 
    0.87, 0.88, 0.88, 0.88, 0.87, 0.88, 0.89, 0.93, 0.93, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.92, 0.9, 0.91, 
    0.92, 0.91, 0.91, 0.92, 0.91, 0.91, 0.92, 0.93, 0.93, 0.91, 0.94, 0.92, 
    0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.93, 0.96, 0.97, 
    0.97, 0.98, 0.97, 0.97, 0.97, 0.97, 0.96, 0.84, 0.92, 0.95, 0.95, 0.93, 
    0.9, 0.92, 0.9, 0.86, 0.85, 0.88, 0.85, 0.86, 0.86, 0.9, 0.9, 0.91, 0.92, 
    0.92, 0.91, 0.9, 0.89, 0.92, 0.94, 0.95, 0.94, 0.96, 0.95, 0.94, 0.92, 
    0.91, 0.9, 0.92, 0.91, 0.92, 0.93, 0.91, 0.93, 0.93, 0.91, 0.92, 0.95, 
    0.93, 0.94, 0.93, 0.93, 0.94, 0.93, 0.96, 0.97, 0.97, 0.97, 0.96, 0.96, 
    0.96, 0.96, 0.95, 0.93, 0.93, 0.92, 0.93, 0.93, 0.86, 0.93, 0.97, 0.97, 
    0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.97, 0.97, 
    0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.96, 0.96, 
    0.95, 0.96, 0.97, 0.97, 0.98, 0.97, 0.96, 0.97, 0.97, 0.96, 0.95, 0.95, 
    0.96, 0.94, 0.96, 0.93, 0.93, 0.93, 0.94, 0.94, 0.91, 0.91, 0.92, 0.91, 
    0.92, 0.93, 0.88, 0.93, 0.91, 0.96, 0.95, 0.95, 0.96, 0.91, 0.88, 0.89, 
    0.92, 0.92, 0.9, 0.91, 0.89, 0.88, 0.84, 0.82, 0.87, 0.86, 0.82, 0.84, 
    0.86, 0.85, 0.84, 0.84, 0.83, 0.79, 0.86, 0.88, 0.86, 0.82, 0.85, 0.85, 
    0.83, 0.77, 0.73, 0.76, 0.8, 0.76, 0.78, 0.86, 0.89, 0.94, 0.97, 0.98, 
    0.98, 0.97, 0.93, 0.92, 0.94, 0.97, 0.98, 0.98, 0.96, 0.96, 0.98, 0.98, 
    0.98, 0.98, 0.96, 0.96, 0.96, 0.96, 0.96, 0.94, 0.92, 0.9, 0.88, 0.89, 
    0.91, 0.96, 0.96, 0.98, 0.99, 0.99, 0.98, 0.98, 0.92, 0.93, 0.89, 0.88, 
    0.82, 0.74, 0.74, 0.8, 0.79, 0.73, 0.66, 0.76, 0.82, 0.88, 0.86, 0.95, 
    0.95, 0.9, 0.96, 0.98, 0.93, 0.95, 0.84, 0.77, 0.85, 0.89, 0.88, 0.85, 
    0.88, 0.91, 0.93, 0.92, 0.93, 0.93, 0.95, 0.93, 0.95, 0.96, 0.95, 0.94, 
    0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.92, 0.92, 0.9, 
    0.92, 0.9, 0.86, 0.88, 0.87, 0.87, 0.87, 0.9, 0.88, 0.89, 0.88, 0.9, 
    0.91, 0.92, 0.95, 0.93, 0.91, 0.92, 0.9, 0.87, 0.86, 0.84, 0.82, 0.8, 
    0.79, 0.78, 0.79, 0.81, 0.82, 0.85, 0.84, 0.86, 0.89, 0.89, 0.9, 0.9, 
    0.91, 0.91, 0.95, 0.95, 0.94, 0.97, 0.93, 0.93, 0.96, 0.94, 0.96, 0.92, 
    0.9, 0.92, 0.91, 0.91, 0.9, 0.91, 0.89, 0.92, 0.9, 0.94, 0.92, 0.91, 
    0.89, 0.89, 0.93, 0.94, 0.94, 0.95, 0.94, 0.97, 0.97, 0.92, 0.93, 0.92, 
    0.95, 0.92, 0.92, 0.95, 0.89, 0.89, 0.91, 0.85, 0.93, 0.98, 0.91, 0.89, 
    0.94, 0.97, 0.98, 0.99, 0.99, 0.99, 1, 0.99, 0.97, 0.98, 0.99, 0.96, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.95, 0.97, 0.97, 0.99, 
    0.99, 0.99, 0.99, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.97, 
    0.97, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.97, 0.95, 0.95, 0.93, 0.93, 0.93, 0.95, 0.95, 0.92, 0.93, 0.95, 0.96, 
    0.98, 0.98, 0.97, 0.99, 0.97, 0.98, 0.97, 0.95, 0.95, 0.91, 0.88, 0.92, 
    0.95, 0.94, 0.93, 0.91, 0.91, 0.9, 0.73, 0.86, 0.93, 0.94, 0.96, 0.95, 
    0.95, 0.95, 0.95, 0.93, 0.91, 0.81, 0.86, 0.84, 0.8, 0.88, 0.77, 0.62, 
    0.76, 0.76, 0.79, 0.76, 0.75, 0.7, 0.77, 0.91, 0.96, 0.96, 0.95, 0.96, 
    0.98, 0.97, 0.96, 0.98, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.96, 0.93, 
    0.96, 0.95, 0.94, 0.95, 0.91, 0.93, 0.96, 0.93, 0.9, 0.92, 0.89, 0.93, 
    0.93, 0.92, 0.96, 0.96, 0.98, 0.98, 0.98, 0.95, 0.95, 0.98, 0.93, 0.94, 
    0.93, 0.92, 0.92, 0.91, 0.9, 0.9, 0.89, 0.89, 0.9, 0.86, 0.89, 0.96, 
    0.97, 0.96, 0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.88, 
    0.88, 0.97, 0.97, 0.95, 0.93, 0.95, 0.95, 0.95, 0.93, 0.96, 0.98, 0.99, 
    0.99, 0.99, 0.97, 0.96, 0.98, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 
    0.96, 0.97, 0.96, 0.96, 0.96, 0.94, 0.92, 0.9, 0.89, 0.86, 0.84, 0.79, 
    0.77, 0.83, 0.75, 0.75, 0.7, 0.9, 0.87, 0.87, 0.9, 0.9, 0.91, 0.91, 0.86, 
    0.89, 0.86, 0.82, 0.85, 0.85, 0.89, 0.79, 0.77, 0.83, 0.89, 0.9, 0.9, 
    0.9, 0.88, 0.86, 0.86, 0.88, 0.9, 0.84, 0.82, 0.8, 0.77, 0.81, 0.8, 0.77, 
    0.85, 0.88, 0.89, 0.9, 0.93, 0.89, 0.85, 0.91, 0.94, 0.94, 0.93, 0.87, 
    0.91, 0.92, 0.92, 0.94, 0.97, 0.98, 0.99, 0.99, 0.99, 0.97, 0.97, 0.95, 
    0.96, 0.98, 0.96, 0.93, 0.92, 0.93, 0.93, 0.82, 0.79, 0.81, 0.9, 0.86, 
    0.85, 0.89, 0.84, 0.86, 0.8, 0.79, 0.8, 0.8, 0.8, 0.83, 0.87, 0.8, 0.78, 
    0.78, 0.87, 0.85, 0.82, 0.85, 0.89, 0.91, 0.91, 0.91, 0.93, 0.94, 0.97, 
    0.98, 0.98, 0.92, 0.95, 0.91, 0.92, 0.94, 0.96, 0.97, 0.97, 0.98, 0.99, 
    0.98, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.96, 0.92, 
    0.94, 0.95, 0.94, 0.94, 0.91, 0.91, 0.93, 0.98, 0.99, 0.98, 0.96, 0.94, 
    0.94, 0.98, 0.98, 0.99, 0.99, 0.99, 0.97, 0.95, 0.92, 0.92, 0.88, 0.83, 
    0.81, 0.8, 0.78, 0.76, 0.79, 0.75, 0.8, 0.86, 0.82, 0.79, 0.81, 0.88, 
    0.83, 0.81, 0.92, 0.92, 0.87, 0.86, 0.89, 0.87, 0.86, 0.91, 0.91, 0.91, 
    0.89, 0.86, 0.86, 0.84, 0.84, 0.82, 0.8, 0.84, 0.87, 0.88, 0.93, 0.94, 
    0.96, 0.96, 0.98, 0.99, 0.99, 1, 1, 0.99, 0.99, 0.9, 0.92, 0.9, 0.95, 
    0.9, 0.94, 0.94, 0.92, 0.92, 0.93, 0.97, 0.97, 0.97, 0.98, 0.99, 0.99, 
    0.98, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 
    0.95, 0.91, 0.89, 0.89, 0.88, 0.95, 0.93, 0.94, 0.94, 0.93, 0.92, 0.85, 
    0.96, 0.9, 0.95, 0.96, 0.96, 0.95, 0.85, 0.79, 0.94, 0.96, 0.93, 0.94, 
    0.79, 0.83, 0.78, 0.75, 0.81, 0.9, 0.84, 0.94, 0.94, 0.93, 0.92, 0.92, 
    0.9, 0.91, 0.91, 0.88, 0.92, 0.89, 0.91, 0.91, 0.9, 0.89, 0.93, 0.92, 
    0.9, 0.88, 0.92, 0.93, 0.96, 0.97, 0.98, 0.96, 0.96, 0.96, 0.95, 0.97, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.98, 0.97, 0.98, 0.95, 
    0.93, 0.96, 0.96, 0.97, 0.98, 0.93, 0.95, 0.96, 0.88, 0.84, 0.87, 0.91, 
    0.82, 0.88, 0.93, 0.96, 0.92, 0.88, 0.86, 0.9, 0.95, 0.95, 0.99, 0.97, 
    0.88, 0.95, 0.91, 0.9, 0.83, 0.83, 0.89, 0.95, 0.98, 0.98, 0.97, 0.93, 
    0.82, 0.82, 0.82, 0.85, 0.9, 0.96, 0.98, 0.99, 0.96, 0.96, 0.98, 0.97, 
    0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 0.95, 1, 0.95, 0.99, 1, 
    0.99, 0.99, 0.98, 0.99, 0.98, 0.99, 0.99, 0.98, 0.96, 0.97, 0.99, 0.99, 
    0.98, 0.97, 0.96, 0.96, 0.95, 0.95, 0.96, 0.95, 0.98, 0.98, 0.99, 1, 
    0.95, 0.94, 1, 0.99, 0.96, 0.95, 0.94, 0.91, 0.84, 0.89, 0.89, 0.87, 
    0.84, 0.86, 0.87, 0.88, 0.88, 0.88, 0.89, 0.9, 0.9, 0.91, 0.94, 0.97, 
    0.97, 0.94, 0.95, 0.96, 0.97, 0.98, 0.87, 0.91, 0.92, 0.93, 0.93, 0.86, 
    0.88, 0.84, 0.87, 0.84, 0.87, 0.87, 0.87, 0.89, 0.91, 0.9, 0.91, 0.91, 
    0.94, 0.98, 0.96, 0.91, 0.91, 0.89, 0.87, 0.85, 0.84, 0.89, 0.88, 0.91, 
    0.87, 0.88, 0.9, 0.89, 0.9, 0.91, 0.89, 0.9, 0.9, 0.88, 0.87, 0.88, 0.93, 
    0.92, 0.89, 0.81, 0.91, 0.98, 0.99, 0.99, 1, 0.99, 0.95, 0.97, 0.96, 
    0.98, 0.97, 0.96, 0.95, 0.95, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 1, 
    1, 1, 0.95, 0.88, 0.98, 0.97, 0.96, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 1, 0.99, 0.99, 0.98, 0.98, 0.92, 0.9, 0.91, 0.93, 0.95, 0.98, 
    0.99, 0.99, 1, 0.99, 0.98, 0.89, 0.9, 0.91, 0.92, 0.9, 0.93, 0.93, 0.88, 
    0.9, 0.92, 0.89, 0.91, 0.92, 0.94, 0.92, 0.86, 0.82, 0.92, 0.92, 0.94, 
    0.95, 0.96, 0.94, 0.98, 0.93, 0.89, 0.9, 0.92, 0.88, 0.86, 0.87, 0.88, 
    0.9, 0.91, 0.92, 0.97, 0.98, 0.99, 1, 1, 1, 1, 0.99, 0.99, 0.92, 0.9, 
    0.87, 0.86, 0.88, 0.86, 0.87, 0.97, 0.86, 0.86, 0.82, 0.87, 0.87, 0.9, 
    0.89, 0.86, 0.86, 0.87, 0.89, 0.9, 0.85, 0.9, 0.85, 0.88, 0.9, 0.88, 0.9, 
    0.81, 0.82, 0.81, 0.83, 0.85, 0.86, 0.82, 0.84, 0.8, 0.84, 0.9, 0.91, 
    0.75, 0.71, 0.68, 0.67, 0.85, 0.84, 0.79, 0.81, 0.91, 0.67, 0.71, 0.7, 
    0.72, 0.9, 0.73, 0.86, 0.81, 0.92, 0.85, 0.91, 0.91, 0.9, 0.97, 0.98, 
    0.95, 0.92, 0.95, 0.95, 0.94, 0.95, 0.95, 0.95, 0.95, 0.97, 0.99, 1, 
    0.99, 0.99, 1, 1, 0.99, 0.96, 0.96, 0.94, 0.93, 0.94, 0.94, 0.94, 0.96, 
    0.99, 0.99, 1, 1, 1, 0.98, 0.99, 0.99, 0.99, 1, 1, 1, 0.97, 0.95, 0.91, 
    0.9, 0.91, 0.95, 0.97, 0.97, 0.98, 0.98, 0.99, 1, 1, 1, 1, 0.99, 0.99, 1, 
    0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.91, 0.86, 0.85, 0.88, 0.94, 
    0.92, 0.91, 1, 0.89, 0.9, 0.91, 0.88, 0.87, 1, 1, 0.88, 0.9, 1, 0.9, 
    0.92, 0.92, 1, 1, 0.94, 0.93, 0.96, 0.95, 0.94, 0.95, 0.97, 0.95, 0.97, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.99, 0.98, 0.96, 0.95, 0.96, 
    0.96, 0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.95, 0.96, 0.97, 0.89, 
    0.92, 0.97, 0.98, 0.99, 0.99, 0.99, 1, 0.98, 1, 1, 1, 0.99, 1, 0.99, 
    0.99, 0.99, 0.97, 0.93, 0.9, 0.91, 0.95, 0.96, 0.89, 0.92, 0.96, 0.97, 
    0.99, 1, 1, 0.97, 0.95, 0.99, 1, 0.99, 0.96, 0.93, 0.89, 0.88, 0.86, 
    0.83, 0.78, 0.87, 0.97, 0.97, 0.98, 0.99, 0.98, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.95, 0.95, 0.95, 0.93, 0.89, 0.86, 0.83, 0.87, 0.92, 0.97, 0.99, 
    0.95, 0.9, 0.89, 0.88, 0.9, 0.9, 0.85, 0.88, 0.85, 0.9, 0.93, 0.95, 0.88, 
    0.88, 0.92, 0.92, 0.91, 0.94, 0.89, 0.91, 0.92, 0.84, 0.89, 0.89, 0.89, 
    0.91, 0.92, 0.91, 0.9, 0.87, 0.86, 0.92, 0.88, 0.87, 0.87, 0.84, 0.85, 
    0.85, 0.85, 0.83, 0.82, 0.78, 0.75, 0.76, 0.71, 0.62, 0.66, 0.75, 0.65, 
    0.66, 0.7, 0.74, 0.72, 0.75, 0.73, 0.71, 0.71, 0.71, 0.72, 0.73, 0.73, 
    0.76, 0.74, 0.72, 0.72, 0.72, 0.7, 0.68, 0.66, 0.64, 0.61, 0.6, 0.61, 
    0.61, 0.93, 0.92, 0.92, 0.92, 0.62, 0.62, 0.73, 0.56, 0.59, 0.63, 0.69, 
    0.68, 0.69, 0.69, 0.68, 0.66, 0.64, 0.62, 0.6, 0.58, 0.57, 0.63, 0.61, 
    0.56, 0.53, 0.53, 0.54, 0.59, 0.55, 0.57, 0.68, 0.62, 0.6, 0.59, 0.57, 
    0.55, 0.73, 0.75, 0.72, 0.7, 0.69, 0.69, 0.91, 0.68, 0.68, 0.67, 0.86, 
    0.86, 0.85, 0.6, 0.59, 0.57, 0.61, 0.67, 0.63, 0.63, 0.55, 0.5, 0.52, 
    0.54, 0.5, 0.5, 0.52, 0.53, 0.59, 0.68, 0.81, 0.77, 0.8, 0.82, 0.81, 
    0.81, 0.71, 0.81, 0.79, 0.77, 0.79, 0.79, 0.88, 0.79, 0.8, 0.81, 0.82, 
    0.83, 0.83, 0.84, 0.85, 0.85, 0.83, 0.84, 0.84, 0.83, 0.83, 0.82, 0.81, 
    0.79, 0.82, 0.86, 0.88, 0.86, 0.86, 0.87, 0.87, 0.87, 0.87, 0.83, 0.82, 
    0.87, 0.93, 0.95, 0.94, 0.92, 0.91, 0.88, 0.86, 0.88, 0.89, 0.9, 0.88, 
    0.85, 0.81, 0.79, 0.77, 0.77, 0.82, 0.88, 0.85, 0.77, 0.81, 0.81, 0.82, 
    0.85, 0.9, 0.96, 0.9, 0.93, 0.93, 0.99, 0.99, 1, 1, 0.99, 0.99, 0.99, 
    0.98, 0.99, 0.96, 0.97, 0.96, 0.94, 0.95, 0.95, 0.97, 0.98, 0.94, 0.96, 
    0.97, 0.95, 0.97, 0.99, 1, 1, 1, 1, 1, 1, 0.98, 0.96, 0.91, 0.92, 0.93, 
    0.9, 0.9, 0.94, 0.92, 0.92, 0.92, 0.96, 0.88, 0.88, 0.87, 0.9, 0.91, 0.9, 
    0.9, 0.91, 0.91, 0.9, 0.91, 0.86, 0.88, 0.86, 0.89, 0.89, 0.92, 0.93, 
    0.86, 0.9, 0.91, 0.88, 0.87, 0.87, 0.87, 0.87, 0.89, 0.88, 0.88, 0.91, 
    0.9, 0.89, 0.89, 0.87, 0.85, 0.87, 0.87, 0.86, 0.86, 0.87, 0.85, 0.78, 
    0.8, 0.79, 0.79, 0.8, 0.9, 0.92, 0.84, 0.88, 0.97, 0.99, 0.94, 0.91, 
    0.91, 0.91, 0.92, 0.91, 0.9, 0.9, 0.9, 0.91, 0.93, 0.94, 0.94, 0.92, 
    0.99, 0.99, 1, 1, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.97, 
    0.97, 0.98, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.97, 0.98, 0.97, 0.96, 0.96, 0.93, 
    0.93, 0.98, 0.98, 0.98, 0.99, 0.98, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 
    0.98, 1, 1, 1, 1, 0.95, 1, 0.94, 0.99, 0.97, 0.99, 1, 1, 0.97, 1, 1, 
    0.99, 0.89, 1, 1, 1, 1, 0.98, 1, 1, 1, 0.99, 0.99, 0.98, 0.88, 0.9, 0.97, 
    0.92, 0.95, 0.94, 0.96, 0.96, 0.98, 0.98, 0.98, 0.99, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.99, 1, 1, 0.99, 0.86, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0.98, 0.96, 0.95, 0.94, 0.93, 0.89, 0.92, 0.9, 0.87, 0.96, 0.88, 0.87, 
    0.89, 0.89, 0.91, 0.96, 0.95, 0.95, 0.98, 0.95, 0.93, 0.92, 0.9, 0.93, 
    0.96, 0.99, 1, 1, 1, 1, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 0.99, 1, 1, 1, 1, 
    1, 1, 1, 1, 0.99, 0.99, 0.97, 0.99, 0.97, 0.99, 0.99, 0.97, 0.97, 0.93, 
    0.91, 0.93, 0.93, 0.87, 0.93, 0.96, 0.88, 0.93, 0.91, 0.95, 0.85, 0.97, 
    0.81, 0.85, 0.84, 0.83, 0.84, 0.86, 0.87, 0.86, 0.89, 0.9, 0.9, 0.89, 
    0.87, 0.89, 0.9, 0.91, 0.94, 0.98, 0.97, 0.97, 0.98, 0.99, 1, 1, 1, 1, 1, 
    0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.97, 0.98, 0.97, 1, 0.96, 0.96, 
    0.96, 0.96, 0.93, 0.94, 0.9, 0.94, 0.93, 0.95, 0.95, 0.96, 0.93, 0.96, 
    0.95, 0.93, 0.93, 0.91, 0.9, 0.91, 0.95, 0.95, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.99, 1, 0.97, 0.99, 1, 1, 0.98, 0.99, 0.98, 0.92, 0.87, 0.88, 
    0.92, 0.82, 0.89, 0.9, 0.84, 0.87, 0.89, 0.92, 0.96, 0.97, 0.99, 0.99, 
    0.97, 0.98, 0.98, 0.99, 0.9, 0.88, 0.85, 0.86, 0.95, 0.98, 0.98, 0.99, 
    0.98, 0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.93, 0.96, 0.92, 
    0.92, 0.87, 0.86, 0.91, 0.86, 0.85, 0.85, 0.86, 0.84, 0.86, 0.85, 0.85, 
    0.84, 0.88, 0.89, 0.98, 0.98, 0.98, 0.96, 0.94, 0.98, 0.9, 0.94, 0.99, 
    0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.94, 0.79, 0.92, 0.88, 
    0.89, 0.89, 0.92, 0.95, 0.97, 0.96, 0.93, 0.92, 0.93, 0.9, 0.96, 0.96, 
    0.95, 0.9, 0.94, 0.9, 0.94, 0.93, 0.94, 0.91, 0.95, 0.95, 0.94, 0.92, 
    0.88, 0.86, 0.88, 0.9, 0.87, 0.92, 0.95, 0.93, 0.94, 0.94, 0.94, 0.94, 
    0.97, 0.96, 0.96, 0.97, 0.95, 0.98, 0.98, 0.97, 0.98, 0.97, 0.98, 0.97, 
    0.96, 0.95, 0.93, 0.91, 0.92, 0.9, 0.9, 0.93, 0.92, 0.9, 0.9, 0.88, 0.89, 
    0.9, 0.95, 0.91, 0.88, 0.86, 0.83, 0.8, 0.77, 0.74, 0.86, 0.83, 0.79, 
    0.79, 0.83, 0.83, 0.84, 0.84, 0.83, 0.83, 0.83, 0.83, 0.84, 0.85, 0.92, 
    0.93, 0.89, 0.88, 0.88, 0.88, 0.91, 0.94, 0.9, 0.91, 0.92, 0.92, 0.97, 
    0.97, 0.96, 0.96, 0.95, 0.96, 0.97, 0.96, 0.97, 0.92, 0.95, 0.97, 0.94, 
    0.89, 0.89, 0.91, 0.9, 0.87, 0.84, 0.83, 0.82, 0.86, 0.83, 0.84, 0.83, 
    0.82, 0.77, 0.72, 0.75, 0.79, 0.8, 0.81, 0.83, 0.85, 0.87, 0.82, 0.86, 
    0.84, 0.81, 0.85, 0.83, 0.82, 0.78, 0.76, 0.78, 0.79, 0.79, 0.81, 0.83, 
    0.8, 0.82, 0.81, 0.78, 0.8, 0.82, 0.82, 0.83, 0.82, 0.83, 0.81, 0.83, 
    0.86, 0.85, 0.87, 0.84, 0.89, 0.85, 0.9, 0.88, 0.84, 0.86, 0.89, 0.89, 
    0.86, 0.87, 0.84, 0.9, 0.89, 0.89, 0.89, 0.92, 0.89, 0.92, 0.89, 0.88, 
    0.9, 0.9, 0.9, 0.89, 0.92, 0.88, 0.88, 0.89, 0.91, 0.88, 0.91, 0.89, 
    0.91, 0.89, 0.9, 0.92, 0.89, 0.9, 0.89, 0.89, 0.91, 0.92, 0.88, 0.93, 
    0.94, 0.95, 0.95, 0.94, 0.94, 0.96, 0.95, 0.95, 0.96, 0.96, 0.96, 0.94, 
    0.95, 0.94, 0.95, 0.95, 0.94, 0.88, 0.9, 0.93, 0.96, 0.94, 0.93, 0.92, 
    0.92, 0.93, 0.94, 0.94, 0.93, 0.89, 0.91, 0.9, 0.85, 0.93, 0.89, 0.91, 
    0.89, 0.87, 0.91, 0.9, 0.85, 0.88, 0.87, 0.9, 0.9, 0.91, 0.92, 0.89, 
    0.92, 0.9, 0.92, 0.93, 0.89, 0.91, 0.92, 0.93, 0.9, 0.93, 0.92, 0.91, 
    0.86, 0.86, 0.88, 0.89, 0.92, 0.92, 0.92, 0.94, 0.94, 0.93, 0.93, 0.93, 
    0.95, 0.95, 0.97, 0.97, 0.96, 0.95, 0.94, 0.93, 0.94, 0.94, 0.93, 0.93, 
    0.93, 0.94, 0.94, 0.92, 0.93, 0.95, 0.97, 0.97, 0.98, 0.94, 0.94, 0.93, 
    0.93, 0.93, 0.94, 0.95, 0.98, 0.99, 0.98, 0.92, 0.91, 0.89, 0.89, 0.9, 
    0.97, 0.98, 0.97, 0.95, 0.95, 0.95, 0.95, 0.97, 0.98, 0.97, 0.95, 0.94, 
    0.95, 0.95, 0.96, 0.97, 0.97, 0.98, 0.99, 0.98, 0.94, 0.92, 0.9, 0.89, 
    0.97, 0.97, 0.98, 0.97, 0.98, 0.96, 0.96, 0.98, 0.95, 0.94, 0.95, 0.93, 
    0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.94, 0.95, 0.94, 0.93, 0.94, 0.93, 
    0.87, 0.88, 0.88, 0.89, 0.87, 0.86, 0.87, 0.91, 0.9, 0.91, 0.92, 0.93, 
    0.89, 0.82, 0.78, 0.76, 0.78, 0.78, 0.73, 0.78, 0.77, 0.74, 0.71, 0.73, 
    0.76, 0.74, 0.84, 0.93, 0.96, 0.94, 0.93, 0.94, 0.93, 0.86, 0.77, 0.8, 
    0.85, 0.83, 0.83, 0.83, 0.82, 0.78, 0.81, 0.8, 0.79, 0.78, 0.76, 0.76, 
    0.76, 0.8, 0.81, 0.82, 0.85, 0.92, 0.93, 0.9, 0.89, 0.88, 0.88, 0.88, 
    0.9, 0.9, 0.91, 0.91, 0.94, 0.96, 0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 
    0.93, 0.88, 0.85, 0.8, 0.83, 0.85, 0.91, 0.96, 0.97, 0.98, 0.98, 0.97, 
    0.94, 0.91, 0.93, 0.92, 0.93, 0.93, 0.95, 0.92, 0.92, 0.91, 0.91, 0.93, 
    0.89, 0.98, 0.98, 0.98, 0.98, 0.97, 0.94, 0.95, 0.97, 0.95, 0.91, 0.9, 
    0.91, 0.9, 0.88, 0.82, 0.83, 0.9, 0.91, 0.9, 0.88, 0.87, 0.89, 0.85, 
    0.88, 0.92, 0.95, 0.97, 0.98, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.93, 0.93, 0.89, 0.9, 
    0.91, 0.89, 0.88, 0.85, 0.86, 0.87, 0.91, 0.92, 0.89, 0.92, 0.92, 0.92, 
    0.94, 0.89, 0.87, 0.94, 0.94, 0.95, 0.95, 0.92, 0.95, 0.91, 0.89, 0.89, 
    0.89, 0.9, 0.89, 0.89, 0.89, 0.89, 0.92, 0.9, 0.91, 0.93, 0.93, 0.94, 
    0.94, 0.96, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 
    0.95, 0.88, 0.88, 0.88, 0.89, 0.93, 0.96, 0.98, 0.98, 0.97, 0.96, 0.95, 
    0.95, 0.95, 0.92, 0.92, 0.81, 0.89, 0.93, 0.92, 0.89, 0.88, 0.9, 0.88, 
    0.88, 0.92, 0.97, 0.98, 0.98, 0.9, 0.78, 0.83, 0.93, 0.9, 0.79, 0.72, 
    0.73, 0.75, 0.71, 0.83, 0.87, 0.88, 0.88, 0.9, 0.86, 0.87, 0.9, 0.95, 
    0.89, 0.93, 0.93, 0.95, 0.91, 0.92, 0.96, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.93, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.98, 0.97, 0.98, 0.99, 0.98, 0.97, 0.96, 0.96, 0.97, 0.96, 0.97, 
    0.95, 0.86, 0.83, 0.85, 0.83, 0.78, 0.81, 0.88, 0.84, 0.79, 0.91, 0.88, 
    0.86, 0.87, 0.91, 0.93, 0.86, 0.86, 0.85, 0.87, 0.88, 0.87, 0.87, 0.88, 
    0.92, 0.95, 0.93, 0.94, 0.97, 0.97, 0.97, 0.98, 0.98, 0.95, 0.93, 0.95, 
    0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.96, 0.96, 0.97, 0.96, 0.96, 0.97, 
    0.98, 0.96, 0.98, 0.96, 0.97, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.96, 
    0.94, 0.94, 0.96, 0.96, 0.95, 0.92, 0.88, 0.89, 0.87, 0.85, 0.83, 0.84, 
    0.82, 0.83, 0.83, 0.85, 0.73, 0.77, 0.8, 0.82, 0.83, 0.83, 0.82, 0.77, 
    0.8, 0.84, 0.81, 0.86, 0.89, 0.84, 0.81, 0.82, 0.86, 0.86, 0.86, 0.86, 
    0.87, 0.89, 0.89, 0.87, 0.91, 0.89, 0.9, 0.89, 0.96, 0.98, 0.94, 0.91, 
    0.92, 0.91, 0.89, 0.89, 0.86, 0.89, 0.93, 0.95, 0.95, 0.97, 0.96, 0.96, 
    0.96, 0.96, 0.92, 0.92, 0.93, 0.93, 0.92, 0.92, 0.91, 0.88, 0.84, 0.83, 
    0.83, 0.88, 0.82, 0.79, 0.79, 0.82, 0.8, 0.78, 0.74, 0.74, 0.76, 0.78, 
    0.76, 0.79, 0.75, 0.75, 0.73, 0.77, 0.78, 0.78, 0.8, 0.82, 0.81, 0.8, 
    0.79, 0.76, 0.77, 0.77, 0.78, 0.85, 0.92, 0.89, 0.93, 0.93, 0.93, 0.93, 
    0.95, 0.97, 0.98, 0.99, 0.98, 0.97, 0.98, 0.96, 0.98, 0.97, 0.98, 0.97, 
    0.97, 0.96, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.96, 0.94, 0.93, 0.92, 0.97, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.95, 0.98, 0.96, 0.95, 0.98, 0.98, 0.97, 0.97, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.96, 0.98, 0.99, 0.99, 
    0.98, 0.95, 0.94, 0.9, 0.86, 0.85, 0.86, 0.87, 0.88, 0.87, 0.87, 0.88, 
    0.84, 0.85, 0.86, 0.85, 0.86, 0.87, 0.85, 0.83, 0.85, 0.83, 0.83, 0.83, 
    0.77, 0.83, 0.79, 0.86, 0.92, 0.85, 0.84, 0.78, 0.78, 0.78, 0.77, 0.76, 
    0.76, 0.75, 0.73, 0.71, 0.71, 0.7, 0.68, 0.7, 0.69, 0.68, 0.68, 0.67, 
    0.66, 0.65, 0.65, 0.65, 0.65, 0.65, 0.62, 0.62, 0.65, 0.68, 0.68, 0.66, 
    0.66, 0.67, 0.65, 0.6, 0.58, 0.58, 0.58, 0.66, 0.67, 0.67, 0.68, 0.68, 
    0.68, 0.68, 0.69, 0.7, 0.71, 0.72, 0.74, 0.68, 0.71, 0.72, 0.73, 0.75, 
    0.78, 0.81, 0.82, 0.83, 0.8, 0.8, 0.81, 0.95, 0.95, 0.94, 0.93, 0.93, 
    0.92, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.92, 0.92, 0.92, 0.92, 0.92, 
    0.92, 0.93, 0.93, 0.93, 0.94, 0.94, 0.9, 0.78, 0.81, 0.86, 0.9, 0.94, 
    0.95, 0.93, 0.9, 0.88, 0.89, 0.87, 0.84, 0.83, 0.82, 0.83, 0.84, 0.84, 
    0.87, 0.84, 0.82, 0.83, 0.87, 0.89, 0.88, 0.86, 0.83, 0.87, 0.74, 0.75, 
    0.79, 0.83, 0.89, 0.91, 0.92, 0.9, 0.87, 0.89, 0.85, 0.89, 0.91, 0.93, 
    0.9, 0.94, 0.95, 0.94, 0.96, 0.97, 0.98, 0.98, 0.99, 0.98, 0.92, 0.92, 
    0.91, 0.92, 0.92, 0.92, 0.89, 0.89, 0.94, 0.92, 0.89, 0.89, 0.88, 0.92, 
    0.91, 0.92, 0.9, 0.92, 0.91, 0.92, 0.92, 0.94, 0.93, 0.93, 0.94, 0.91, 
    0.9, 0.9, 0.92, 0.91, 0.92, 0.93, 0.94, 0.95, 0.96, 0.98, 0.99, 0.99, 
    0.99, 0.95, 0.93, 0.91, 0.89, 0.86, 0.82, 0.89, 0.9, 0.93, 0.93, 0.94, 
    0.94, 0.94, 0.93, 0.92, 0.93, 0.93, 0.94, 0.94, 0.93, 0.92, 0.91, 0.9, 
    0.87, 0.87, 0.88, 0.89, 0.9, 0.92, 0.93, 0.95, 0.95, 0.97, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.96, 0.94, 0.94, 
    0.94, 0.95, 0.95, 0.96, 0.98, 0.99, 0.98, 0.98, 0.99, 0.99, 0.99, 0.95, 
    0.9, 0.86, 0.83, 0.82, 0.88, 0.94, 0.95, 0.95, 0.94, 0.9, 0.91, 0.93, 
    0.93, 0.95, 0.89, 0.94, 0.92, 0.91, 0.92, 0.89, 0.94, 0.93, 0.91, 0.9, 
    0.9, 0.91, 0.94, 0.93, 0.91, 0.94, 0.94, 0.89, 0.89, 0.92, 0.91, 0.9, 
    0.89, 0.88, 0.9, 0.9, 0.89, 0.93, 0.95, 0.93, 0.95, 0.93, 0.92, 0.95, 
    0.92, 0.93, 0.89, 0.93, 0.92, 0.94, 0.92, 0.94, 0.91, 0.91, 0.92, 0.94, 
    0.92, 0.93, 0.91, 0.92, 0.93, 0.93, 0.97, 0.98, 0.98, 0.98, 0.95, 0.91, 
    0.93, 0.93, 0.97, 0.97, 0.97, 0.96, 0.95, 0.89, 0.91, 0.92, 0.89, 0.93, 
    0.92, 0.92, 0.92, 0.95, 0.94, 0.93, 0.96, 0.96, 0.96, 0.97, 0.97, 0.95, 
    0.95, 0.94, 0.94, 0.94, 0.95, 0.95, 0.94, 0.93, 0.93, 0.94, 0.94, 0.94, 
    0.89, 0.92, 0.91, 0.86, 0.86, 0.87, 0.89, 0.91, 0.93, 0.93, 0.94, 0.95, 
    0.96, 0.95, 0.95, 0.96, 0.97, 0.98, 0.98, 0.95, 0.95, 0.96, 0.96, 0.98, 
    0.98, 0.98, 0.97, 0.95, 0.97, 0.97, 0.97, 0.97, 0.95, 0.94, 0.92, 0.93, 
    0.95, 0.94, 0.95, 0.95, 0.94, 0.93, 0.94, 0.93, 0.93, 0.95, 0.96, 0.97, 
    0.98, 0.97, 0.95, 0.96, 0.94, 0.9, 0.9, 0.83, 0.82, 0.81, 0.86, 0.84, 
    0.88, 0.92, 0.93, 0.88, 0.89, 0.89, 0.89, 0.9, 0.93, 0.96, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.96, 0.94, 0.93, 0.91, 0.88, 
    0.87, 0.85, 0.84, 0.84, 0.82, 0.79, 0.76, 0.74, 0.78, 0.82, 0.81, 0.86, 
    0.85, 0.8, 0.75, 0.73, 0.81, 0.7, 0.69, 0.72, 0.71, 0.64, 0.61, 0.61, 
    0.74, 0.81, 0.76, 0.76, 0.79, 0.76, 0.76, 0.75, 0.71, 0.71, 0.77, 0.71, 
    0.82, 0.79, 0.81, 0.77, 0.79, 0.78, 0.77, 0.79, 0.78, 0.8, 0.84, 0.83, 
    0.72, 0.74, 0.67, 0.74, 0.71, 0.85, 0.85, 0.69, 0.67, 0.77, 0.78, 0.85, 
    0.87, 0.77, 0.78, 0.73, 0.72, 0.71, 0.73, 0.7, 0.67, 0.83, 0.81, 0.78, 
    0.73, 0.82, 0.75, 0.71, 0.74, 0.7, 0.72, 0.73, 0.74, 0.72, 0.74, 0.71, 
    0.67, 0.7, 0.68, 0.73, 0.76, 0.76, 0.75, 0.74, 0.75, 0.73, 0.78, 0.78, 
    0.8, 0.77, 0.8, 0.87, 0.86, 0.91, 0.93, 0.93, 0.94, 0.93, 0.94, 0.93, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 
    0.94, 0.95, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.94, 0.95, 0.96, 
    0.94, 0.93, 0.9, 0.9, 0.89, 0.88, 0.87, 0.89, 0.92, 0.93, 0.94, 0.93, 
    0.9, 0.88, 0.91, 0.9, 0.86, 0.87, 0.89, 0.88, 0.86, 0.85, 0.82, 0.76, 
    0.76, 0.75, 0.79, 0.8, 0.78, 0.8, 0.82, 0.76, 0.72, 0.79, 0.72, 0.76, 
    0.8, 0.78, 0.8, 0.66, 0.64, 0.7, 0.67, 0.72, 0.76, 0.8, 0.81, 0.81, 0.83, 
    0.87, 0.8, 0.79, 0.88, 0.89, 0.89, 0.68, 0.77, 0.64, 0.66, 0.64, 0.74, 
    0.63, 0.7, 0.81, 0.71, 0.69, 0.7, 0.8, 0.75, 0.74, 0.69, 0.77, 0.83, 
    0.82, 0.77, 0.76, 0.82, 0.77, 0.79, 0.69, 0.81, 0.79, 0.72, 0.76, 0.76, 
    0.79, 0.8, 0.75, 0.78, 0.76, 0.74, 0.73, 0.69, 0.76, 0.82, 0.72, 0.73, 
    0.71, 0.68, 0.73, 0.71, 0.73, 0.73, 0.7, 0.7, 0.7, 0.72, 0.69, 0.7, 0.71, 
    0.72, 0.72, 0.76, 0.79, 0.81, 0.81, 0.82, 0.87, 0.9, 0.89, 0.89, 0.89, 
    0.89, 0.88, 0.9, 0.9, 0.91, 0.91, 0.91, 0.91, 0.92, 0.93, 0.93, 0.94, 
    0.95, 0.93, 0.95, 0.94, 0.95, 0.96, 0.96, 0.96, 0.98, 0.98, 0.99, 0.99, 
    0.98, 0.98, 0.98, 0.97, 0.98, 0.98, 0.97, 0.96, 0.95, 0.94, 0.92, 0.94, 
    0.93, 0.97, 0.98, 0.99, 0.98, 0.96, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.94, 0.93, 0.89, 0.93, 0.96, 0.93, 0.91, 0.93, 0.91, 0.89, 
    0.89, 0.88, 0.92, 0.94, 0.97, 0.98, 0.98, 0.97, 0.91, 0.95, 0.94, 0.92, 
    0.9, 0.89, 0.88, 0.87, 0.88, 0.88, 0.88, 0.9, 0.89, 0.87, 0.86, 0.87, 
    0.87, 0.86, 0.88, 0.85, 0.86, 0.87, 0.88, 0.88, 0.91, 0.89, 0.89, 0.88, 
    0.84, 0.83, 0.84, 0.83, 0.8, 0.83, 0.84, 0.83, 0.8, 0.81, 0.8, 0.82, 
    0.82, 0.87, 0.84, 0.76, 0.8, 0.76, 0.73, 0.8, 0.78, 0.74, 0.71, 0.68, 
    0.75, 0.69, 0.64, 0.72, 0.74, 0.69, 0.66, 0.59, 0.67, 0.73, 0.64, 0.65, 
    0.66, 0.75, 0.83, 0.87, 0.83, 0.88, 0.74, 0.72, 0.79, 0.74, 0.71, 0.83, 
    0.8, 0.79, 0.87, 0.79, 0.77, 0.77, 0.84, 0.83, 0.7, 0.8, 0.63, 0.59, 
    0.62, 0.65, 0.64, 0.63, 0.84, 0.83, 0.83, 0.8, 0.76, 0.65, 0.63, 0.67, 
    0.69, 0.62, 0.6, 0.53, 0.52, 0.53, 0.64, 0.5, 0.57, 0.54, 0.61, 0.64, 
    0.66, 0.71, 0.74, 0.76, 0.77, 0.82, 0.78, 0.76, 0.82, 0.82, 0.73, 0.76, 
    0.76, 0.77, 0.83, 0.89, 0.85, 0.85, 0.83, 0.88, 0.88, 0.83, 0.86, 0.89, 
    0.92, 0.94, 0.96, 0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.98, 0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.96, 
    0.96, 0.95, 0.96, 0.93, 0.93, 0.92, 0.93, 0.93, 0.93, 0.91, 0.96, 0.9, 
    0.91, 0.92, 0.92, 0.92, 0.95, 0.96, 0.96, 0.95, 0.93, 0.88, 0.86, 0.85, 
    0.82, 0.82, 0.83, 0.85, 0.87, 0.86, 0.86, 0.85, 0.86, 0.85, 0.87, 0.84, 
    0.88, 0.86, 0.84, 0.83, 0.82, 0.85, 0.85, 0.85, 0.84, 0.81, 0.83, 0.82, 
    0.81, 0.81, 0.79, 0.83, 0.87, 0.88, 0.85, 0.83, 0.88, 0.85, 0.82, 0.82, 
    0.82, 0.78, 0.72, 0.68, 0.7, 0.71, 0.86, 0.89, 0.92, 0.9, 0.88, 0.88, 
    0.88, 0.85, 0.86, 0.82, 0.7, 0.66, 0.65, 0.74, 0.76, 0.73, 0.83, 0.68, 
    0.66, 0.78, 0.8, 0.82, 0.82, 0.88, 0.87, 0.85, 0.9, 0.82, 0.8, 0.83, 
    0.92, 0.86, 0.86, 0.86, 0.86, 0.83, 0.81, 0.82, 0.79, 0.81, 0.87, 0.85, 
    0.85, 0.82, 0.86, 0.88, 0.91, 0.91, 0.92, 0.94, 0.95, 0.96, 0.95, 0.95, 
    0.96, 0.96, 0.96, 0.97, 0.98, 0.98, 0.96, 0.98, 0.98, 0.98, 0.99, 0.99, 
    0.95, 0.92, 0.92, 0.93, 0.91, 0.93, 0.96, 0.96, 0.98, 0.99, 0.98, 0.95, 
    0.92, 0.92, 0.92, 0.92, 0.9, 0.9, 0.9, 0.92, 0.94, 0.9, 0.91, 0.91, 0.91, 
    0.95, 0.98, 0.98, 0.98, 0.97, 0.96, 0.95, 0.93, 0.92, 0.91, 0.87, 0.87, 
    0.89, 0.91, 0.92, 0.93, 0.94, 0.87, 0.88, 0.87, 0.84, 0.86, 0.88, 0.88, 
    0.9, 0.86, 0.9, 0.87, 0.88, 0.87, 0.86, 0.83, 0.84, 0.81, 0.81, 0.73, 
    0.78, 0.78, 0.76, 0.79, 0.77, 0.78, 0.75, 0.76, 0.76, 0.76, 0.76, 0.77, 
    0.8, 0.78, 0.7, 0.8, 0.69, 0.69, 0.74, 0.69, 0.69, 0.73, 0.76, 0.78, 
    0.74, 0.81, 0.86, 0.88, 0.91, 0.9, 0.94, 0.94, 0.91, 0.92, 0.93, 0.95, 
    0.95, 0.86, 0.83, 0.75, 0.89, 0.86, 0.94, 0.93, 0.89, 0.89, 0.93, 0.92, 
    0.92, 0.88, 0.88, 0.88, 0.85, 0.85, 0.86, 0.85, 0.84, 0.78, 0.82, 0.79, 
    0.86, 0.83, 0.84, 0.92, 0.92, 0.91, 0.89, 0.83, 0.85, 0.8, 0.81, 0.84, 
    0.79, 0.78, 0.8, 0.81, 0.76, 0.73, 0.74, 0.73, 0.71, 0.74, 0.74, 0.73, 
    0.72, 0.74, 0.79, 0.86, 0.9, 0.89, 0.89, 0.86, 0.9, 0.84, 0.76, 0.76, 
    0.76, 0.78, 0.82, 0.84, 0.92, 0.93, 0.95, 0.93, 0.88, 0.88, 0.86, 0.78, 
    0.8, 0.73, 0.67, 0.81, 0.65, 0.64, 0.61, 0.62, 0.67, 0.69, 0.7, 0.72, 
    0.8, 0.82, 0.88, 0.81, 0.77, 0.62, 0.75, 0.69, 0.58, 0.6, 0.66, 0.64, 
    0.66, 0.85, 0.86, 0.84, 0.88, 0.87, 0.91, 0.93, 0.9, 0.89, 0.92, 0.91, 
    0.86, 0.8, 0.79, 0.76, 0.76, 0.73, 0.77, 0.75, 0.78, 0.79, 0.77, 0.79, 
    0.72, 0.73, 0.71, 0.71, 0.8, 0.78, 0.75, 0.83, 0.84, 0.78, 0.79, 0.83, 
    0.86, 0.84, 0.87, 0.85, 0.89, 0.85, 0.8, 0.81, 0.8, 0.8, 0.8, 0.78, 0.77, 
    0.77, 0.85, 0.85, 0.83, 0.84, 0.84, 0.76, 0.82, 0.88, 0.92, 0.77, 0.74, 
    0.79, 0.78, 0.77, 0.79, 0.88, 0.8, 0.85, 0.78, 0.79, 0.8, 0.78, 0.8, 
    0.79, 0.76, 0.76, 0.83, 0.81, 0.77, 0.73, 0.89, 0.76, 0.78, 0.76, 0.75, 
    0.76, 0.67, 0.68, 0.81, 0.79, 0.8, 0.83, 0.79, 0.79, 0.79, 0.79, 0.78, 
    0.79, 0.77, 0.79, 0.77, 0.74, 0.76, 0.75, 0.77, 0.83, 0.82, 0.77, 0.77, 
    0.84, 0.74, 0.84, 0.74, 0.79, 0.76, 0.82, 0.85, 0.83, 0.79, 0.78, 0.75, 
    0.75, 0.78, 0.79, 0.82, 0.78, 0.81, 0.82, 0.83, 0.84, 0.85, 0.87, 0.88, 
    0.87, 0.88, 0.87, 0.88, 0.88, 0.89, 0.88, 0.88, 0.89, 0.9, 0.92, 0.91, 
    0.92, 0.93, 0.92, 0.92, 0.93, 0.91, 0.92, 0.91, 0.9, 0.9, 0.89, 0.88, 
    0.88, 0.88, 0.88, 0.87, 0.88, 0.9, 0.89, 0.87, 0.87, 0.81, 0.82, 0.84, 
    0.85, 0.85, 0.85, 0.86, 0.86, 0.87, 0.88, 0.89, 0.88, 0.89, 0.88, 0.88, 
    0.9, 0.91, 0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 0.94, 0.92, 0.91, 0.91, 
    0.91, 0.91, 0.92, 0.92, 0.91, 0.9, 0.92, 0.94, 0.95, 0.96, 0.95, 0.91, 
    0.88, 0.9, 0.92, 0.94, 0.95, 0.96, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.94, 0.92, 0.94, 0.94, 0.95, 0.95, 0.95, 0.94, 0.95, 
    0.96, 0.97, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 
    0.96, 0.95, 0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 0.98, 0.98, 
    0.98, 0.97, 0.96, 0.94, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.94, 0.95, 0.97, 0.98, 0.95, 0.91, 0.87, 0.91, 0.91, 0.91, 0.91, 0.91, 
    0.91, 0.91, 0.9, 0.89, 0.88, 0.88, 0.91, 0.83, 0.93, 0.85, 0.85, 0.87, 
    0.85, 0.87, 0.86, 0.87, 0.87, 0.87, 0.87, 0.85, 0.85, 0.84, 0.84, 0.83, 
    0.87, 0.86, 0.93, 0.93, 0.91, 0.89, 0.86, 0.82, 0.85, 0.85, 0.84, 0.83, 
    0.85, 0.85, 0.83, 0.79, 0.82, 0.79, 0.83, 0.82, 0.83, 0.8, 0.86, 0.85, 
    0.83, 0.83, 0.83, 0.82, 0.82, 0.83, 0.82, 0.78, 0.75, 0.83, 0.84, 0.81, 
    0.73, 0.74, 0.78, 0.75, 0.7, 0.72, 0.76, 0.68, 0.72, 0.77, 0.76, 0.79, 
    0.77, 0.76, 0.75, 0.75, 0.73, 0.7, 0.72, 0.68, 0.67, 0.68, 0.75, 0.65, 
    0.72, 0.8, 0.63, 0.74, 0.72, 0.73, 0.66, 0.67, 0.59, 0.66, 0.72, 0.57, 
    0.69, 0.62, 0.75, 0.61, 0.69, 0.6, 0.66, 0.67, 0.64, 0.67, 0.7, 0.67, 
    0.67, 0.65, 0.68, 0.69, 0.7, 0.69, 0.74, 0.76, 0.77, 0.79, 0.79, 0.81, 
    0.82, 0.85, 0.85, 0.85, 0.83, 0.83, 0.85, 0.86, 0.85, 0.87, 0.87, 0.84, 
    0.84, 0.83, 0.83, 0.8, 0.78, 0.79, 0.78, 0.8, 0.76, 0.78, 0.67, 0.78, 
    0.75, 0.8, 0.77, 0.77, 0.69, 0.72, 0.76, 0.65, 0.66, 0.67, 0.61, 0.71, 
    0.64, 0.66, 0.66, 0.75, 0.69, 0.76, 0.74, 0.62, 0.79, 0.8, 0.79, 0.74, 
    0.75, 0.74, 0.71, 0.77, 0.75, 0.74, 0.74, 0.72, 0.73, 0.77, 0.73, 0.71, 
    0.68, 0.71, 0.76, 0.78, 0.82, 0.82, 0.8, 0.73, 0.75, 0.84, 0.74, 0.85, 
    0.8, 0.73, 0.82, 0.69, 0.79, 0.72, 0.68, 0.63, 0.62, 0.6, 0.59, 0.62, 
    0.65, 0.61, 0.59, 0.57, 0.72, 0.61, 0.59, 0.74, 0.78, 0.82, 0.84, 0.83, 
    0.83, 0.82, 0.8, 0.82, 0.8, 0.8, 0.79, 0.8, 0.79, 0.82, 0.81, 0.83, 0.82, 
    0.85, 0.85, 0.86, 0.86, 0.85, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.86, 0.84, 0.85, 0.85, 0.85, 0.84, 0.83, 0.84, 
    0.83, 0.82, 0.82, 0.81, 0.81, 0.82, 0.83, 0.81, 0.82, 0.82, 0.82, 0.82, 
    0.82, 0.8, 0.8, 0.79, 0.77, 0.77, 0.75, 0.79, 0.73, 0.75, 0.76, 0.75, 
    0.69, 0.64, 0.67, 0.64, 0.71, 0.67, 0.72, 0.77, 0.73, 0.73, 0.75, 0.77, 
    0.77, 0.78, 0.83, 0.84, 0.83, 0.82, 0.84, 0.84, 0.83, 0.84, 0.84, 0.84, 
    0.84, 0.84, 0.84, 0.84, 0.83, 0.84, 0.84, 0.84, 0.85, 0.86, 0.84, 0.83, 
    0.84, 0.85, 0.86, 0.84, 0.85, 0.87, 0.88, 0.88, 0.88, 0.89, 0.89, 0.89, 
    0.89, 0.89, 0.89, 0.9, 0.89, 0.89, 0.89, 0.9, 0.89, 0.87, 0.87, 0.9, 
    0.92, 0.93, 0.92, 0.93, 0.93, 0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.92, 
    0.93, 0.92, 0.91, 0.92, 0.93, 0.94, 0.94, 0.93, 0.94, 0.93, 0.95, 0.93, 
    0.94, 0.95, 0.94, 0.96, 0.95, 0.95, 0.95, 0.95, 0.94, 0.91, 0.92, 0.93, 
    0.92, 0.92, 0.92, 0.92, 0.92, 0.9, 0.92, 0.91, 0.9, 0.9, 0.9, 0.9, 0.89, 
    0.89, 0.89, 0.9, 0.89, 0.8, 0.85, 0.84, 0.86, 0.9, 0.92, 0.92, 0.91, 
    0.88, 0.89, 0.88, 0.88, 0.87, 0.86, 0.84, 0.82, 0.82, 0.8, 0.8, 0.79, 
    0.76, 0.75, 0.8, 0.79, 0.78, 0.77, 0.77, 0.72, 0.77, 0.77, 0.67, 0.71, 
    0.7, 0.69, 0.72, 0.74, 0.67, 0.68, 0.69, 0.67, 0.66, 0.7, 0.71, 0.71, 
    0.74, 0.78, 0.82, 0.84, 0.85, 0.86, 0.87, 0.88, 0.9, 0.91, 0.93, 0.94, 
    0.94, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 0.94, 0.91, 0.87, 
    0.85, 0.86, 0.86, 0.86, 0.85, 0.83, 0.83, 0.83, 0.83, 0.82, 0.81, 0.81, 
    0.79, 0.79, 0.79, 0.78, 0.78, 0.79, 0.79, 0.78, 0.79, 0.79, 0.77, 0.8, 
    0.81, 0.81, 0.85, 0.79, 0.81, 0.82, 0.8, 0.74, 0.72, 0.73, 0.72, 0.72, 
    0.78, 0.75, 0.68, 0.71, 0.73, 0.76, 0.75, 0.74, 0.73, 0.8, 0.79, 0.74, 
    0.71, 0.77, 0.78, 0.79, 0.77, 0.74, 0.76, 0.75, 0.73, 0.71, 0.7, 0.71, 
    0.73, 0.76, 0.75, 0.82, 0.78, 0.74, 0.72, 0.72, 0.72, 0.68, 0.72, 0.72, 
    0.73, 0.75, 0.76, 0.76, 0.77, 0.8, 0.78, 0.76, 0.74, 0.75, 0.75, 0.72, 
    0.7, 0.73, 0.79, 0.84, 0.86, 0.87, 0.88, 0.88, 0.87, 0.89, 0.87, 0.78, 
    0.8, 0.82, 0.79, 0.83, 0.85, 0.79, 0.84, 0.89, 0.84, 0.89, 0.9, 0.9, 
    0.89, 0.89, 0.9, 0.89, 0.9, 0.93, 0.95, 0.95, 0.94, 0.94, 0.92, 0.92, 
    0.91, 0.93, 0.93, 0.93, 0.95, 0.95, 0.94, 0.93, 0.92, 0.91, 0.91, 0.92, 
    0.93, 0.94, 0.95, 0.94, 0.93, 0.94, 0.94, 0.94, 0.95, 0.96, 0.97, 0.98, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.93, 0.99, 0.99, 0.99, 
    0.97, 0.98, 0.96, 0.94, 0.94, 0.95, 0.98, 0.99, 0.99, 0.94, 0.89, 0.87, 
    0.85, 0.83, 0.8, 0.85, 0.83, 0.84, 0.84, 0.87, 0.88, 0.98, 0.88, 0.89, 
    0.91, 0.93, 0.96, 0.98, 0.99, 0.98, 0.96, 0.95, 0.94, 0.95, 0.95, 0.94, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 0.96, 0.94, 0.92, 0.92, 0.92, 0.91, 
    0.92, 0.93, 0.94, 0.97, 0.98, 0.98, 0.97, 0.96, 0.95, 0.94, 0.91, 0.93, 
    0.9, 0.9, 0.87, 0.92, 0.94, 0.94, 0.95, 0.96, 0.94, 0.95, 0.95, 0.94, 
    0.93, 0.9, 0.9, 0.9, 0.91, 0.93, 0.94, 0.95, 0.95, 0.96, 0.97, 0.97, 
    0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.93, 0.89, 0.83, 
    0.85, 0.85, 0.75, 0.79, 0.86, 0.84, 0.83, 0.82, 0.81, 0.81, 0.81, 0.82, 
    0.83, 0.83, 0.83, 0.84, 0.9, 0.9, 0.9, 0.9, 0.87, 0.89, 0.89, 0.87, 0.77, 
    0.73, 0.77, 0.77, 0.87, 0.85, 0.83, 0.81, 0.82, 0.83, 0.84, 0.85, 0.87, 
    0.89, 0.93, 0.8, 0.76, 0.75, 0.77, 0.81, 0.84, 0.87, 0.84, 0.82, 0.81, 
    0.81, 0.79, 0.85, 0.69, 0.64, 0.76, 0.79, 0.77, 0.78, 0.77, 0.78, 0.74, 
    0.77, 0.77, 0.76, 0.81, 0.73, 0.77, 0.73, 0.7, 0.73, 0.74, 0.73, 0.76, 
    0.75, 0.74, 0.73, 0.73, 0.72, 0.73, 0.75, 0.72, 0.72, 0.7, 0.72, 0.71, 
    0.73, 0.73, 0.74, 0.75, 0.76, 0.8, 0.83, 0.81, 0.79, 0.79, 0.78, 0.77, 
    0.79, 0.79, 0.78, 0.77, 0.76, 0.76, 0.77, 0.77, 0.86, 0.75, 0.75, 0.78, 
    0.83, 0.78, 0.8, 0.8, 0.79, 0.78, 0.78, 0.79, 0.8, 0.8, 0.79, 0.76, 0.76, 
    0.76, 0.76, 0.76, 0.77, 0.78, 0.79, 0.77, 0.77, 0.77, 0.74, 0.72, 0.72, 
    0.73, 0.72, 0.76, 0.73, 0.72, 0.72, 0.71, 0.71, 0.67, 0.7, 0.68, 0.7, 
    0.71, 0.68, 0.7, 0.68, 0.68, 0.69, 0.67, 0.67, 0.67, 0.67, 0.68, 0.65, 
    0.7, 0.65, 0.69, 0.7, 0.71, 0.71, 0.72, 0.75, 0.78, 0.76, 0.76, 0.77, 
    0.78, 0.75, 0.74, 0.76, 0.77, 0.78, 0.78, 0.77, 0.78, 0.73, 0.73, 0.72, 
    0.69, 0.71, 0.71, 0.74, 0.77, 0.69, 0.69, 0.77, 0.75, 0.73, 0.81, 0.86, 
    0.71, 0.73, 0.73, 0.73, 0.69, 0.7, 0.7, 0.7, 0.66, 0.8, 0.73, 0.8, 0.8, 
    0.78, 0.83, 0.82, 0.79, 0.8, 0.81, 0.82, 0.83, 0.82, 0.79, 0.85, 0.82, 
    0.84, 0.8, 0.83, 0.83, 0.8, 0.75, 0.75, 0.81, 0.74, 0.78, 0.73, 0.81, 
    0.65, 0.65, 0.7, 0.78, 0.85, 0.83, 0.85, 0.81, 0.78, 0.77, 0.74, 0.75, 
    0.69, 0.7, 0.71, 0.81, 0.82, 0.88, 0.89, 0.88, 0.81, 0.84, 0.83, 0.85, 
    0.85, 0.79, 0.74, 0.73, 0.67, 0.8, 0.63, 0.61, 0.62, 0.66, 0.65, 0.76, 
    0.85, 0.75, 0.75, 0.8, 0.85, 0.89, 0.9, 0.91, 0.89, 0.92, 0.94, 0.94, 
    0.93, 0.87, 0.88, 0.89, 0.88, 0.89, 0.89, 0.91, 0.91, 0.91, 0.89, 0.88, 
    0.91, 0.94, 0.94, 0.91, 0.92, 0.94, 0.94, 0.93, 0.93, 0.93, 0.93, 0.94, 
    0.94, 0.95, 0.94, 0.94, 0.95, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.95, 
    0.96, 0.95, 0.95, 0.9, 0.9, 0.91, 0.93, 0.93, 0.93, 0.9, 0.91, 0.91, 
    0.92, 0.94, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.95, 0.95, 
    0.95, 0.95, 0.91, 0.92, 0.93, 0.92, 0.91, 0.91, 0.92, 0.91, 0.91, 0.91, 
    0.92, 0.92, 0.93, 0.93, 0.9, 0.88, 0.9, 0.9, 0.92, 0.92, 0.93, 0.92, 
    0.88, 0.8, 0.81, 0.79, 0.84, 0.84, 0.85, 0.85, 0.82, 0.81, 0.81, 0.8, 
    0.79, 0.8, 0.81, 0.82, 0.87, 0.91, 0.89, 0.91, 0.92, 0.92, 0.92, 0.92, 
    0.88, 0.88, 0.87, 0.84, 0.8, 0.82, 0.84, 0.88, 0.88, 0.89, 0.9, 0.9, 
    0.86, 0.81, 0.85, 0.87, 0.9, 0.9, 0.9, 0.93, 0.87, 0.81, 0.9, 0.88, 0.89, 
    0.81, 0.87, 0.83, 0.82, 0.78, 0.83, 0.8, 0.78, 0.77, 0.77, 0.79, 0.88, 
    0.89, 0.9, 0.87, 0.89, 0.93, 0.94, 0.91, 0.83, 0.82, 0.87, 0.87, 0.88, 
    0.89, 0.88, 0.9, 0.9, 0.91, 0.93, 0.94, 0.92, 0.91, 0.93, 0.92, 0.88, 
    0.91, 0.95, 0.96, 0.97, 0.97, 0.96, 0.95, 0.94, 0.94, 0.96, 0.95, 0.94, 
    0.96, 0.96, 0.95, 0.96, 0.96, 0.96, 0.95, 0.96, 0.96, 0.96, 0.96, 0.97, 
    0.96, 0.96, 0.95, 0.93, 0.92, 0.98, 0.98, 0.98, 0.96, 0.95, 0.92, 0.88, 
    0.84, 0.81, 0.8, 0.81, 0.8, 0.83, 0.85, 0.85, 0.79, 0.79, 0.8, 0.82, 
    0.85, 0.89, 0.89, 0.87, 0.86, 0.88, 0.87, 0.89, 0.87, 0.86, 0.85, 0.85, 
    0.88, 0.85, 0.84, 0.83, 0.72, 0.83, 0.87, 0.87, 0.87, 0.87, 0.86, 0.84, 
    0.85, 0.84, 0.82, 0.81, 0.87, 0.87, 0.88, 0.9, 0.9, 0.89, 0.9, 0.89, 
    0.89, 0.89, 0.88, 0.86, 0.84, 0.82, 0.82, 0.87, 0.86, 0.9, 0.89, 0.88, 
    0.89, 0.89, 0.89, 0.87, 0.87, 0.88, 0.88, 0.9, 0.86, 0.91, 0.89, 0.88, 
    0.9, 0.92, 0.91, 0.91, 0.91, 0.91, 0.89, 0.9, 0.86, 0.83, 0.77, 0.89, 
    0.86, 0.85, 0.85, 0.83, 0.82, 0.81, 0.79, 0.78, 0.83, 0.82, 0.78, 0.85, 
    0.88, 0.86, 0.89, 0.88, 0.9, 0.9, 0.9, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 
    0.9, 0.92, 0.91, 0.93, 0.95, 0.97, 0.98, 0.98, 0.97, 0.95, 0.96, 0.93, 
    0.92, 0.93, 0.93, 0.94, 0.94, 0.93, 0.94, 0.96, 0.96, 0.95, 0.94, 0.92, 
    0.92, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.92, 0.91, 0.9, 0.9, 0.9, 
    0.89, 0.89, 0.92, 0.93, 0.92, 0.9, 0.91, 0.89, 0.87, 0.87, 0.88, 0.91, 
    0.9, 0.9, 0.86, 0.88, 0.88, 0.86, 0.88, 0.88, 0.88, 0.89, 0.89, 0.89, 
    0.91, 0.92, 0.93, 0.9, 0.89, 0.88, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 
    0.89, 0.88, 0.88, 0.9, 0.88, 0.86, 0.85, 0.84, 0.83, 0.85, 0.84, 0.85, 
    0.87, 0.85, 0.85, 0.87, 0.85, 0.86, 0.87, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.87, 0.85, 0.87, 0.86, 0.86, 0.87, 0.86, 0.87, 0.86, 0.86, 0.85, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.85, 0.85, 0.86, 0.87, 0.87, 0.86, 
    0.87, 0.86, 0.87, 0.86, 0.86, 0.86, 0.87, 0.87, 0.87, 0.87, 0.87, 0.88, 
    0.86, 0.84, 0.84, 0.82, 0.82, 0.83, 0.82, 0.83, 0.75, 0.8, 0.81, 0.83, 
    0.82, 0.83, 0.87, 0.85, 0.85, 0.84, 0.84, 0.85, 0.84, 0.84, 0.85, 0.86, 
    0.84, 0.86, 0.85, 0.85, 0.86, 0.84, 0.84, 0.91, 0.89, 0.9, 0.87, 0.85, 
    0.84, 0.84, 0.78, 0.81, 0.73, 0.77, 0.8, 0.79, 0.8, 0.76, 0.8, 0.77, 
    0.79, 0.76, 0.74, 0.77, 0.76, 0.75, 0.79, 0.78, 0.76, 0.8, 0.78, 0.79, 
    0.72, 0.64, 0.67, 0.72, 0.75, 0.71, 0.73, 0.75, 0.81, 0.8, 0.78, 0.77, 
    0.79, 0.74, 0.77, 0.76, 0.76, 0.78, 0.81, 0.74, 0.81, 0.84, 0.84, 0.82, 
    0.74, 0.79, 0.76, 0.78, 0.72, 0.68, 0.68, 0.68, 0.7, 0.69, 0.69, 0.69, 
    0.68, 0.67, 0.63, 0.58, 0.58, 0.58, 0.58, 0.51, 0.44, 0.5, 0.47, 0.59, 
    0.55, 0.43, 0.48, 0.68, 0.78, 0.77, 0.76, 0.76, 0.76, 0.77, 0.8, 0.82, 
    0.83, 0.84, 0.87, 0.86, 0.88, 0.88, 0.88, 0.87, 0.86, 0.85, 0.84, 0.84, 
    0.86, 0.86, 0.87, 0.87, 0.89, 0.89, 0.89, 0.88, 0.89, 0.89, 0.89, 0.89, 
    0.89, 0.91, 0.9, 0.9, 0.92, 0.93, 0.92, 0.94, 0.93, 0.92, 0.94, 0.96, 
    0.96, 0.96, 0.95, 0.96, 0.94, 0.92, 0.89, 0.88, 0.87, 0.86, 0.81, 0.83, 
    0.89, 0.86, 0.85, 0.86, 0.84, 0.84, 0.83, 0.84, 0.82, 0.81, 0.82, 0.78, 
    0.81, 0.86, 0.8, 0.78, 0.81, 0.78, 0.81, 0.82, 0.81, 0.78, 0.83, 0.83, 
    0.83, 0.89, 0.86, 0.81, 0.75, 0.81, 0.83, 0.76, 0.78, 0.79, 0.77, 0.76, 
    0.75, 0.7, 0.75, 0.7, 0.69, 0.71, 0.65, 0.71, 0.68, 0.63, 0.62, 0.63, 
    0.66, 0.69, 0.73, 0.71, 0.72, 0.7, 0.86, 0.79, 0.77, 0.76, 0.75, 0.73, 
    0.76, 0.79, 0.8, 0.86, 0.82, 0.84, 0.84, 0.83, 0.78, 0.85, 0.83, 0.85, 
    0.69, 0.76, 0.74, 0.71, 0.73, 0.73, 0.75, 0.77, 0.79, 0.83, 0.88, 0.9, 
    0.92, 0.9, 0.9, 0.89, 0.89, 0.86, 0.79, 0.78, 0.83, 0.84, 0.85, 0.85, 
    0.85, 0.79, 0.84, 0.85, 0.88, 0.93, 0.91, 0.89, 0.89, 0.87, 0.89, 0.89, 
    0.9, 0.89, 0.88, 0.87, 0.87, 0.87, 0.87, 0.89, 0.9, 0.9, 0.91, 0.92, 
    0.91, 0.91, 0.9, 0.89, 0.88, 0.89, 0.89, 0.89, 0.88, 0.87, 0.87, 0.87, 
    0.88, 0.92, 0.92, 0.92, 0.9, 0.9, 0.9, 0.86, 0.88, 0.83, 0.82, 0.83, 
    0.85, 0.9, 0.9, 0.91, 0.9, 0.89, 0.89, 0.88, 0.89, 0.89, 0.88, 0.86, 
    0.89, 0.89, 0.89, 0.9, 0.88, 0.91, 0.9, 0.9, 0.88, 0.89, 0.87, 0.86, 
    0.87, 0.91, 0.94, 0.93, 0.95, 0.94, 0.95, 0.96, 0.95, 0.97, 0.94, 0.93, 
    0.8, 0.85, 0.85, 0.86, 0.87, 0.9, 0.93, 0.93, 0.94, 0.94, 0.92, 0.95, 
    0.94, 0.95, 0.94, 0.91, 0.84, 0.87, 0.87, 0.85, 0.83, 0.83, 0.89, 0.95, 
    0.94, 0.93, 0.92, 0.93, 0.92, 0.92, 0.92, 0.96, 0.97, 0.95, 0.96, 0.96, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 
    0.97, 0.96, 0.96, 0.95, 0.97, 0.96, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 0.97, 0.95, 
    0.95, 0.95, 0.93, 0.92, 0.87, 0.84, 0.79, 0.84, 0.92, 0.94, 0.94, 0.93, 
    0.92, 0.92, 0.92, 0.92, 0.91, 0.9, 0.92, 0.92, 0.92, 0.94, 0.96, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.98, 0.96, 0.96, 0.97, 
    0.96, 0.94, 0.92, 0.88, 0.85, 0.85, 0.88, 0.92, 0.93, 0.95, 0.96, 0.94, 
    0.95, 0.92, 0.89, 0.89, 0.9, 0.91, 0.91, 0.92, 0.93, 0.93, 0.88, 0.9, 
    0.9, 0.9, 0.86, 0.84, 0.82, 0.77, 0.65, 0.72, 0.67, 0.65, 0.67, 0.66, 
    0.69, 0.63, 0.69, 0.65, 0.67, 0.75, 0.78, 0.84, 0.87, 0.86, 0.85, 0.84, 
    0.86, 0.88, 0.87, 0.89, 0.85, 0.86, 0.85, 0.83, 0.81, 0.81, 0.78, 0.79, 
    0.79, 0.79, 0.8, 0.81, 0.81, 0.85, 0.82, 0.81, 0.81, 0.79, 0.78, 0.74, 
    0.79, 0.79, 0.8, 0.79, 0.8, 0.79, 0.8, 0.81, 0.82, 0.81, 0.81, 0.79, 0.8, 
    0.8, 0.8, 0.79, 0.79, 0.79, 0.81, 0.81, 0.81, 0.82, 0.8, 0.73, 0.71, 
    0.74, 0.7, 0.69, 0.74, 0.75, 0.76, 0.78, 0.8, 0.77, 0.75, 0.71, 0.76, 
    0.74, 0.72, 0.76, 0.78, 0.77, 0.8, 0.8, 0.83, 0.84, 0.82, 0.78, 0.81, 
    0.82, 0.78, 0.8, 0.8, 0.8, 0.8, 0.79, 0.83, 0.83, 0.83, 0.81, 0.8, 0.74, 
    0.78, 0.82, 0.77, 0.79, 0.69, 0.8, 0.8, 0.81, 0.78, 0.76, 0.78, 0.77, 
    0.76, 0.77, 0.81, 0.82, 0.82, 0.79, 0.79, 0.81, 0.8, 0.81, 0.78, 0.8, 
    0.82, 0.82, 0.82, 0.83, 0.81, 0.86, 0.86, 0.84, 0.83, 0.81, 0.84, 0.84, 
    0.84, 0.85, 0.85, 0.86, 0.88, 0.89, 0.88, 0.87, 0.86, 0.89, 0.86, 0.87, 
    0.84, 0.87, 0.89, 0.91, 0.91, 0.91, 0.91, 0.92, 0.93, 0.93, 0.92, 0.91, 
    0.93, 0.95, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.94, 0.95, 0.95, 0.96, 
    0.96, 0.96, 0.97, 0.96, 0.96, 0.95, 0.94, 0.92, 0.9, 0.89, 0.89, 0.89, 
    0.88, 0.89, 0.89, 0.89, 0.89, 0.9, 0.9, 0.89, 0.89, 0.89, 0.9, 0.9, 0.89, 
    0.88, 0.89, 0.89, 0.88, 0.88, 0.88, 0.87, 0.88, 0.89, 0.9, 0.92, 0.93, 
    0.91, 0.9, 0.91, 0.91, 0.89, 0.88, 0.89, 0.89, 0.91, 0.91, 0.91, 0.91, 
    0.91, 0.91, 0.92, 0.93, 0.96, 0.97, 0.96, 0.96, 0.96, 0.95, 0.96, 0.97, 
    0.93, 0.96, 0.96, 0.95, 0.97, 0.98, 0.99, 0.99, 0.98, 0.97, 0.95, 0.96, 
    0.95, 0.94, 0.96, 0.98, 0.98, 0.97, 0.97, 0.96, 0.97, 0.96, 0.97, 0.95, 
    0.96, 0.96, 0.96, 0.96, 0.95, 0.91, 0.91, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.94, 0.95, 0.95, 0.94, 0.94, 0.91, 0.91, 0.85, 0.84, 0.9, 0.87, 0.93, 
    0.92, 0.87, 0.85, 0.83, 0.82, 0.86, 0.92, 0.9, 0.87, 0.85, 0.84, 0.83, 
    0.82, 0.92, 0.89, 0.84, 0.82, 0.85, 0.9, 0.97, 0.97, 0.95, 0.9, 0.9, 
    0.92, 0.9, 0.88, 0.89, 0.86, 0.79, 0.79, 0.78, 0.79, 0.78, 0.82, 0.88, 
    0.83, 0.82, 0.88, 0.89, 0.86, 0.88, 0.92, 0.88, 0.88, 0.87, 0.88, 0.89, 
    0.89, 0.86, 0.89, 0.88, 0.86, 0.95, 0.93, 0.92, 0.91, 0.87, 0.83, 0.81, 
    0.81, 0.81, 0.88, 0.86, 0.89, 0.91, 0.92, 0.91, 0.89, 0.87, 0.88, 0.89, 
    0.91, 0.89, 0.86, 0.88, 0.89, 0.9, 0.86, 0.85, 0.82, 0.85, 0.86, 0.87, 
    0.93, 0.92, 0.91, 0.93, 0.87, 0.94, 0.97, 0.95, 0.96, 0.94, 0.92, 0.89, 
    0.84, 0.85, 0.81, 0.86, 0.87, 0.85, 0.88, 0.85, 0.89, 0.92, 0.92, 0.9, 
    0.9, 0.91, 0.92, 0.94, 0.95, 0.96, 0.96, 0.96, 0.91, 0.92, 0.93, 0.95, 
    0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 0.99, 0.98, 
    0.98, 0.98, 0.97, 0.95, 0.89, 0.87, 0.86, 0.87, 0.86, 0.87, 0.9, 0.91, 
    0.92, 0.9, 0.91, 0.93, 0.94, 0.95, 0.95, 0.95, 0.95, 0.98, 0.98, 0.99, 
    0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.98, 0.89, 0.87, 0.9, 0.9, 0.93, 
    0.91, 0.92, 0.89, 0.88, 0.86, 0.84, 0.83, 0.85, 0.84, 0.73, 0.71, 0.73, 
    0.75, 0.74, 0.73, 0.74, 0.72, 0.72, 0.75, 0.77, 0.79, 0.78, 0.85, 0.9, 
    0.89, 0.9, 0.89, 0.88, 0.88, 0.85, 0.85, 0.86, 0.86, 0.88, 0.83, 0.84, 
    0.81, 0.78, 0.81, 0.76, 0.75, 0.78, 0.78, 0.76, 0.79, 0.76, 0.74, 0.74, 
    0.75, 0.72, 0.78, 0.65, 0.68, 0.73, 0.78, 0.82, 0.73, 0.69, 0.79, 0.8, 
    0.82, 0.77, 0.69, 0.76, 0.7, 0.72, 0.76, 0.8, 0.83, 0.73, 0.76, 0.79, 
    0.68, 0.69, 0.71, 0.7, 0.75, 0.73, 0.69, 0.75, 0.72, 0.78, 0.82, 0.8, 
    0.74, 0.76, 0.78, 0.77, 0.78, 0.73, 0.77, 0.84, 0.74, 0.83, 0.71, 0.79, 
    0.82, 0.76, 0.78, 0.75, 0.77, 0.79, 0.78, 0.84, 0.83, 0.8, 0.86, 0.83, 
    0.79, 0.77, 0.79, 0.77, 0.79, 0.82, 0.84, 0.85, 0.87, 0.84, 0.81, 0.83, 
    0.81, 0.72, 0.74, 0.78, 0.72, 0.81, 0.85, 0.82, 0.8, 0.78, 0.83, 0.85, 
    0.84, 0.85, 0.76, 0.78, 0.79, 0.78, 0.78, 0.77, 0.76, 0.77, 0.76, 0.74, 
    0.78, 0.78, 0.79, 0.78, 0.77, 0.77, 0.79, 0.8, 0.78, 0.77, 0.79, 0.8, 
    0.79, 0.79, 0.79, 0.72, 0.85, 0.76, 0.77, 0.81, 0.75, 0.75, 0.81, 0.84, 
    0.81, 0.79, 0.81, 0.79, 0.79, 0.79, 0.81, 0.76, 0.79, 0.73, 0.84, 0.83, 
    0.75, 0.79, 0.8, 0.75, 0.8, 0.79, 0.8, 0.77, 0.78, 0.77, 0.75, 0.78, 
    0.81, 0.74, 0.8, 0.76, 0.8, 0.75, 0.78, 0.82, 0.78, 0.82, 0.8, 0.84, 
    0.83, 0.8, 0.77, 0.78, 0.77, 0.79, 0.83, 0.78, 0.78, 0.78, 0.79, 0.79, 
    0.8, 0.81, 0.8, 0.82, 0.8, 0.81, 0.83, 0.84, 0.85, 0.82, 0.84, 0.85, 
    0.84, 0.8, 0.8, 0.79, 0.8, 0.8, 0.83, 0.74, 0.75, 0.71, 0.72, 0.74, 0.73, 
    0.68, 0.69, 0.76, 0.75, 0.73, 0.72, 0.71, 0.79, 0.67, 0.74, 0.74, 0.72, 
    0.7, 0.7, 0.69, 0.7, 0.69, 0.72, 0.74, 0.69, 0.67, 0.67, 0.67, 0.73, 
    0.65, 0.77, 0.82, 0.84, 0.86, 0.87, 0.88, 0.88, 0.87, 0.87, 0.88, 0.88, 
    0.9, 0.88, 0.89, 0.89, 0.89, 0.89, 0.89, 0.9, 0.89, 0.92, 0.92, 0.92, 
    0.93, 0.95, 0.95, 0.93, 0.94, 0.93, 0.93, 0.92, 0.9, 0.9, 0.9, 0.88, 0.9, 
    0.9, 0.89, 0.87, 0.91, 0.91, 0.93, 0.9, 0.88, 0.91, 0.92, 0.94, 0.91, 
    0.91, 0.93, 0.94, 0.93, 0.91, 0.91, 0.9, 0.91, 0.92, 0.9, 0.9, 0.91, 
    0.91, 0.92, 0.92, 0.92, 0.92, 0.91, 0.92, 0.91, 0.93, 0.93, 0.93, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 
    0.93, 0.94, 0.93, 0.93, 0.93, 0.92, 0.93, 0.92, 0.92, 0.91, 0.89, 0.9, 
    0.91, 0.92, 0.9, 0.88, 0.89, 0.89, 0.9, 0.9, 0.9, 0.91, 0.91, 0.92, 0.81, 
    0.76, 0.77, 0.8, 0.86, 0.86, 0.86, 0.89, 0.89, 0.86, 0.86, 0.9, 0.89, 
    0.84, 0.87, 0.84, 0.8, 0.81, 0.81, 0.8, 0.77, 0.8, 0.8, 0.84, 0.85, 0.85, 
    0.83, 0.86, 0.84, 0.84, 0.84, 0.83, 0.86, 0.85, 0.85, 0.86, 0.84, 0.85, 
    0.84, 0.84, 0.83, 0.83, 0.84, 0.82, 0.82, 0.86, 0.86, 0.83, 0.8, 0.79, 
    0.81, 0.78, 0.78, 0.8, 0.81, 0.76, 0.77, 0.78, 0.77, 0.75, 0.71, 0.7, 
    0.69, 0.74, 0.77, 0.69, 0.7, 0.72, 0.71, 0.71, 0.77, 0.76, 0.76, 0.74, 
    0.72, 0.72, 0.72, 0.72, 0.73, 0.75, 0.77, 0.78, 0.78, 0.79, 0.82, 0.87, 
    0.85, 0.83, 0.82, 0.81, 0.81, 0.8, 0.83, 0.82, 0.82, 0.81, 0.79, 0.81, 
    0.83, 0.84, 0.84, 0.87, 0.88, 0.68, 0.78, 0.82, 0.68, 0.68, 0.71, 0.7, 
    0.75, 0.87, 0.85, 0.88, 0.87, 0.86, 0.81, 0.83, 0.84, 0.8, 0.85, 0.81, 
    0.79, 0.83, 0.85, 0.89, 0.87, 0.9, 0.94, 0.85, 0.82, 0.86, 0.89, 0.9, 
    0.88, 0.87, 0.79, 0.76, 0.83, 0.79, 0.83, 0.88, 0.88, 0.89, 0.88, 0.87, 
    0.89, 0.88, 0.9, 0.9, 0.9, 0.89, 0.92, 0.9, 0.92, 0.92, 0.91, 0.9, 0.87, 
    0.85, 0.85, 0.85, 0.9, 0.92, 0.83, 0.83, 0.78, 0.82, 0.84, 0.75, 0.69, 
    0.79, 0.87, 0.87, 0.86, 0.86, 0.81, 0.82, 0.83, 0.87, 0.91, 0.88, 0.85, 
    0.85, 0.8, 0.82, 0.8, 0.79, 0.86, 0.86, 0.89, 0.76, 0.75, 0.76, 0.75, 
    0.74, 0.76, 0.8, 0.75, 0.8, 0.86, 0.87, 0.89, 0.86, 0.93, 0.95, 0.94, 
    0.94, 0.92, 0.9, 0.89, 0.89, 0.9, 0.87, 0.91, 0.93, 0.94, 0.93, 0.94, 
    0.91, 0.89, 0.89, 0.89, 0.88, 0.85, 0.86, 0.87, 0.87, 0.88, 0.86, 0.82, 
    0.81, 0.85, 0.81, 0.82, 0.85, 0.82, 0.84, 0.83, 0.83, 0.82, 0.83, 0.86, 
    0.87, 0.85, 0.86, 0.86, 0.91, 0.92, 0.93, 0.87, 0.87, 0.89, 0.92, 0.92, 
    0.88, 0.89, 0.82, 0.88, 0.83, 0.83, 0.83, 0.82, 0.84, 0.84, 0.88, 0.84, 
    0.86, 0.91, 0.93, 0.86, 0.85, 0.81, 0.8, 0.81, 0.81, 0.82, 0.79, 0.74, 
    0.76, 0.77, 0.73, 0.76, 0.71, 0.76, 0.72, 0.73, 0.78, 0.78, 0.72, 0.76, 
    0.77, 0.78, 0.78, 0.74, 0.67, 0.74, 0.73, 0.73, 0.71, 0.72, 0.71, 0.77, 
    0.73, 0.78, 0.82, 0.83, 0.83, 0.83, 0.82, 0.81, 0.83, 0.81, 0.81, 0.88, 
    0.9, 0.89, 0.87, 0.87, 0.87, 0.86, 0.86, 0.85, 0.86, 0.86, 0.85, 0.85, 
    0.85, 0.82, 0.82, 0.82, 0.81, 0.82, 0.82, 0.83, 0.82, 0.83, 0.84, 0.85, 
    0.84, 0.84, 0.84, 0.85, 0.85, 0.85, 0.84, 0.85, 0.86, 0.86, 0.86, 0.86, 
    0.86, 0.86, 0.85, 0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.84, 0.85, 0.85, 
    0.85, 0.86, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 0.84, 0.85, 0.81, 0.79, 
    0.83, 0.81, 0.8, 0.79, 0.79, 0.83, 0.81, 0.82, 0.83, 0.82, 0.84, 0.85, 
    0.84, 0.86, 0.85, 0.83, 0.85, 0.82, 0.82, 0.82, 0.85, 0.86, 0.87, 0.86, 
    0.85, 0.85, 0.85, 0.84, 0.86, 0.84, 0.84, 0.83, 0.81, 0.81, 0.81, 0.84, 
    0.84, 0.84, 0.85, 0.84, 0.85, 0.86, 0.87, 0.87, 0.88, 0.87, 0.85, 0.87, 
    0.86, 0.86, 0.86, 0.85, 0.84, 0.83, 0.81, 0.84, 0.83, 0.84, 0.84, 0.87, 
    0.85, 0.86, 0.84, 0.81, 0.8, 0.8, 0.81, 0.82, 0.81, 0.81, 0.8, 0.8, 0.79, 
    0.81, 0.8, 0.79, 0.78, 0.8, 0.74, 0.74, 0.76, 0.76, 0.8, 0.74, 0.75, 
    0.79, 0.8, 0.85, 0.85, 0.81, 0.82, 0.81, 0.83, 0.78, 0.78, 0.78, 0.81, 
    0.77, 0.78, 0.76, 0.74, 0.81, 0.84, 0.83, 0.85, 0.87, 0.88, 0.88, 0.9, 
    0.9, 0.83, 0.82, 0.81, 0.83, 0.85, 0.89, 0.9, 0.93, 0.93, 0.93, 0.94, 
    0.94, 0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.96, 0.97, 0.91, 0.92, 0.93, 
    0.92, 0.95, 0.96, 0.94, 0.91, 0.9, 0.93, 0.92, 0.93, 0.9, 0.92, 0.92, 
    0.93, 0.92, 0.92, 0.92, 0.91, 0.88, 0.86, 0.87, 0.86, 0.86, 0.84, 0.87, 
    0.88, 0.85, 0.87, 0.87, 0.86, 0.86, 0.85, 0.82, 0.83, 0.83, 0.82, 0.84, 
    0.83, 0.81, 0.82, 0.8, 0.8, 0.81, 0.8, 0.81, 0.8, 0.8, 0.79, 0.78, 0.79, 
    0.79, 0.79, 0.79, 0.78, 0.77, 0.78, 0.76, 0.75, 0.76, 0.75, 0.78, 0.78, 
    0.81, 0.8, 0.8, 0.82, 0.84, 0.84, 0.83, 0.85, 0.84, 0.85, 0.87, 0.86, 
    0.83, 0.88, 0.88, 0.89, 0.89, 0.88, 0.89, 0.9, 0.87, 0.86, 0.89, 0.89, 
    0.85, 0.81, 0.82, 0.83, 0.8, 0.73, 0.78, 0.78, 0.78, 0.81, 0.82, 0.81, 
    0.83, 0.87, 0.87, 0.86, 0.83, 0.82, 0.82, 0.82, 0.87, 0.87, 0.85, 0.87, 
    0.87, 0.87, 0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 0.84, 0.8, 0.83, 0.82, 
    0.81, 0.85, 0.88, 0.87, 0.86, 0.85, 0.85, 0.84, 0.85, 0.87, 0.86, 0.85, 
    0.85, 0.83, 0.82, 0.83, 0.78, 0.81, 0.76, 0.79, 0.79, 0.78, 0.8, 0.79, 
    0.79, 0.79, 0.81, 0.83, 0.84, 0.84, 0.82, 0.82, 0.81, 0.8, 0.79, 0.77, 
    0.75, 0.76, 0.78, 0.81, 0.78, 0.79, 0.81, 0.8, 0.8, 0.82, 0.82, 0.81, 
    0.83, 0.8, 0.81, 0.8, 0.81, 0.8, 0.82, 0.85, 0.84, 0.8, 0.8, 0.8, 0.8, 
    0.76, 0.76, 0.75, 0.79, 0.77, 0.58, 0.53, 0.46, 0.42, 0.46, 0.43, 0.4, 
    0.45, 0.5, 0.63, 0.71, 0.65, 0.54, 0.54, 0.58, 0.46, 0.5, 0.6, 0.66, 
    0.64, 0.63, 0.61, 0.68, 0.53, 0.48, 0.72, 0.85, 0.89, 0.94, 0.96, 0.93, 
    0.91, 0.84, 0.78, 0.88, 0.85, 0.86, 0.65, 0.66, 0.64, 0.65, 0.7, 0.67, 
    0.74, 0.76, 0.78, 0.79, 0.7, 0.71, 0.71, 0.74, 0.64, 0.78, 0.87, 0.91, 
    0.91, 0.9, 0.89, 0.88, 0.88, 0.82, 0.79, 0.76, 0.77, 0.78, 0.84, 0.89, 
    0.86, 0.86, 0.89, 0.83, 0.83, 0.74, 0.73, 0.75, 0.87, 0.96, 0.95, 0.95, 
    0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.97, 0.97, 0.96, 0.97, 0.96, 0.96, 
    0.95, 0.93, 0.93, 0.9, 0.96, 0.93, 0.92, 0.9, 0.89, 0.86, 0.87, 0.87, 
    0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 0.91, 0.92, 0.89, 0.86, 0.83, 
    0.79, 0.77, 0.8, 0.79, 0.79, 0.81, 0.82, 0.81, 0.81, 0.81, 0.81, 0.78, 
    0.8, 0.8, 0.8, 0.82, 0.81, 0.83, 0.83, 0.81, 0.79, 0.77, 0.73, 0.71, 0.7, 
    0.69, 0.7, 0.67, 0.65, 0.71, 0.74, 0.77, 0.77, 0.8, 0.82, 0.83, 0.84, 
    0.85, 0.85, 0.85, 0.86, 0.86, 0.85, 0.83, 0.81, 0.79, 0.77, 0.75, 0.77, 
    0.77, 0.78, 0.75, 0.76, 0.74, 0.77, 0.77, 0.76, 0.76, 0.82, 0.83, 0.84, 
    0.81, 0.81, 0.8, 0.77, 0.79, 0.79, 0.79, 0.78, 0.76, 0.75, 0.74, 0.73, 
    0.75, 0.77, 0.76, 0.77, 0.78, 0.78, 0.8, 0.81, 0.82, 0.81, 0.81, 0.8, 
    0.8, 0.8, 0.8, 0.76, 0.82, 0.83, 0.85, 0.86, 0.85, 0.86, 0.85, 0.85, 
    0.84, 0.82, 0.84, 0.84, 0.83, 0.85, 0.84, 0.87, 0.88, 0.91, 0.9, 0.89, 
    0.88, 0.84, 0.81, 0.8, 0.83, 0.83, 0.83, 0.82, 0.82, 0.84, 0.87, 0.88, 
    0.84, 0.8, 0.75, 0.77, 0.81, 0.83, 0.88, 0.87, 0.88, 0.89, 0.9, 0.92, 
    0.93, 0.92, 0.91, 0.91, 0.92, 0.91, 0.92, 0.91, 0.91, 0.91, 0.89, 0.88, 
    0.87, 0.86, 0.85, 0.84, 0.83, 0.85, 0.83, 0.8, 0.8, 0.82, 0.82, 0.84, 
    0.84, 0.82, 0.78, 0.86, 0.86, 0.85, 0.84, 0.76, 0.82, 0.84, 0.84, 0.8, 
    0.82, 0.84, 0.82, 0.8, 0.88, 0.89, 0.89, 0.88, 0.86, 0.87, 0.9, 0.89, 
    0.89, 0.87, 0.87, 0.86, 0.87, 0.88, 0.9, 0.9, 0.89, 0.87, 0.86, 0.86, 
    0.83, 0.8, 0.81, 0.81, 0.86, 0.84, 0.82, 0.83, 0.82, 0.84, 0.85, 0.87, 
    0.88, 0.88, 0.89, 0.9, 0.88, 0.89, 0.93, 0.93, 0.9, 0.87, 0.85, 0.84, 
    0.87, 0.87, 0.87, 0.86, 0.88, 0.87, 0.86, 0.87, 0.87, 0.87, 0.87, 0.88, 
    0.89, 0.88, 0.89, 0.88, 0.88, 0.9, 0.91, 0.9, 0.9, 0.91, 0.91, 0.92, 
    0.92, 0.93, 0.92, 0.92, 0.91, 0.88, 0.88, 0.89, 0.89, 0.88, 0.88, 0.9, 
    0.9, 0.91, 0.9, 0.91, 0.91, 0.92, 0.92, 0.92, 0.88, 0.83, 0.83, 0.84, 
    0.84, 0.86, 0.85, 0.87, 0.89, 0.9, 0.9, 0.9, 0.9, 0.9, 0.89, 0.88, 0.89, 
    0.86, 0.85, 0.84, 0.86, 0.86, 0.89, 0.89, 0.88, 0.88, 0.86, 0.86, 0.86, 
    0.85, 0.85, 0.84, 0.84, 0.84, 0.83, 0.83, 0.83, 0.86, 0.86, 0.87, 0.88, 
    0.9, 0.93, 0.94, 0.94, 0.94, 0.93, 0.93, 0.94, 0.94, 0.95, 0.95, 0.94, 
    0.95, 0.94, 0.93, 0.91, 0.94, 0.93, 0.94, 0.92, 0.94, 0.96, 0.94, 0.96, 
    0.96, 0.97, 0.97, 0.95, 0.93, 0.95, 0.87, 0.91, 0.91, 0.87, 0.89, 0.89, 
    0.89, 0.89, 0.9, 0.9, 0.86, 0.86, 0.85, 0.82, 0.84, 0.83, 0.81, 0.81, 
    0.66, 0.67, 0.67, 0.65, 0.66, 0.64, 0.64, 0.68, 0.76, 0.73, 0.72, 0.63, 
    0.79, 0.79, 0.78, 0.77, 0.79, 0.78, 0.79, 0.8, 0.81, 0.83, 0.84, 0.83, 
    0.79, 0.8, 0.82, 0.8, 0.77, 0.78, 0.78, 0.78, 0.79, 0.8, 0.8, 0.8, 0.8, 
    0.84, 0.83, 0.83, 0.8, 0.78, 0.81, 0.81, 0.8, 0.84, 0.82, 0.82, 0.85, 
    0.84, 0.76, 0.79, 0.8, 0.82, 0.84, 0.84, 0.83, 0.78, 0.8, 0.81, 0.79, 
    0.79, 0.84, 0.81, 0.79, 0.79, 0.84, 0.84, 0.86, 0.84, 0.84, 0.86, 0.86, 
    0.77, 0.74, 0.7, 0.74, 0.82, 0.87, 0.77, 0.82, 0.82, 0.85, 0.86, 0.78, 
    0.72, 0.83, 0.87, 0.83, 0.87, 0.8, 0.76, 0.82, 0.81, 0.88, 0.87, 0.87, 
    0.86, 0.84, 0.83, 0.84, 0.8, 0.84, 0.81, 0.82, 0.84, 0.83, 0.83, 0.83, 
    0.84, 0.81, 0.77, 0.74, 0.8, 0.82, 0.84, 0.86, 0.87, 0.89, 0.9, 0.9, 0.9, 
    0.88, 0.91, 0.84, 0.83, 0.73, 0.86, 0.89, 0.85, 0.87, 0.88, 0.88, 0.87, 
    0.86, 0.85, 0.84, 0.82, 0.83, 0.83, 0.85, 0.86, 0.83, 0.84, 0.79, 0.75, 
    0.67, 0.63, 0.68, 0.72, 0.8, 0.86, 0.88, 0.88, 0.86, 0.86, 0.89, 0.89, 
    0.9, 0.96, 0.96, 0.95, 0.93, 0.94, 0.93, 0.94, 0.93, 0.94, 0.96, 0.93, 
    0.95, 0.91, 0.88, 0.89, 0.91, 0.88, 0.86, 0.87, 0.87, 0.86, 0.84, 0.87, 
    0.86, 0.9, 0.92, 0.93, 0.93, 0.92, 0.92, 0.93, 0.93, 0.92, 0.89, 0.89, 
    0.87, 0.87, 0.9, 0.84, 0.81, 0.8, 0.84, 0.83, 0.83, 0.87, 0.85, 0.82, 
    0.77, 0.84, 0.84, 0.88, 0.91, 0.92, 0.94, 0.92, 0.93, 0.95, 0.91, 0.88, 
    0.85, 0.81, 0.82, 0.84, 0.87, 0.86, 0.8, 0.81, 0.84, 0.76, 0.72, 0.72, 
    0.76, 0.82, 0.81, 0.81, 0.83, 0.83, 0.85, 0.86, 0.87, 0.86, 0.87, 0.88, 
    0.88, 0.89, 0.89, 0.89, 0.89, 0.89, 0.87, 0.87, 0.88, 0.88, 0.9, 0.92, 
    0.94, 0.95, 0.95, 0.96, 0.97, 0.95, 0.96, 0.97, 0.97, 0.98, 0.98, 0.99, 
    0.99, 0.99, 0.98, 0.98, 0.97, 0.94, 0.91, 0.9, 0.91, 0.9, 0.92, 0.95, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 0.96, 
    0.95, 0.94, 0.92, 0.91, 0.88, 0.92, 0.91, 0.89, 0.91, 0.9, 0.89, 0.89, 
    0.89, 0.88, 0.89, 0.88, 0.89, 0.9, 0.92, 0.9, 0.89, 0.87, 0.89, 0.92, 
    0.91, 0.91, 0.93, 0.93, 0.93, 0.94, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 0.97, 0.97, 
    0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.9, 
    0.87, 0.86, 0.83, 0.84, 0.84, 0.79, 0.79, 0.8, 0.81, 0.83, 0.84, 0.85, 
    0.86, 0.84, 0.73, 0.84, 0.86, 0.88, 0.85, 0.82, 0.75, 0.83, 0.77, 0.8, 
    0.81, 0.83, 0.85, 0.87, 0.87, 0.88, 0.89, 0.86, 0.87, 0.87, 0.88, 0.9, 
    0.9, 0.9, 0.87, 0.87, 0.89, 0.87, 0.87, 0.9, 0.92, 0.91, 0.9, 0.92, 0.91, 
    0.89, 0.92, 0.9, 0.9, 0.89, 0.91, 0.89, 0.9, 0.88, 0.91, 0.9, 0.91, 0.91, 
    0.9, 0.86, 0.87, 0.89, 0.92, 0.92, 0.91, 0.91, 0.9, 0.91, 0.91, 0.9, 
    0.91, 0.91, 0.89, 0.87, 0.86, 0.88, 0.86, 0.86, 0.87, 0.87, 0.85, 0.87, 
    0.89, 0.89, 0.88, 0.89, 0.86, 0.87, 0.87, 0.89, 0.9, 0.9, 0.9, 0.88, 
    0.89, 0.89, 0.88, 0.9, 0.87, 0.89, 0.88, 0.88, 0.89, 0.88, 0.88, 0.88, 
    0.83, 0.88, 0.91, 0.9, 0.9, 0.88, 0.9, 0.93, 0.93, 0.88, 0.86, 0.87, 
    0.88, 0.88, 0.87, 0.89, 0.87, 0.87, 0.84, 0.87, 0.89, 0.88, 0.88, 0.89, 
    0.82, 0.82, 0.86, 0.86, 0.86, 0.93, 0.94, 0.95, 0.95, 0.97, 0.98, 0.96, 
    0.96, 0.96, 0.94, 0.93, 0.93, 0.83, 0.88, 0.82, 0.79, 0.83, 0.84, 0.87, 
    0.81, 0.79, 0.86, 0.88, 0.88, 0.93, 0.94, 0.9, 0.89, 0.88, 0.88, 0.91, 
    0.92, 0.91, 0.91, 0.93, 0.92, 0.9, 0.92, 0.92, 0.95, 0.92, 0.92, 0.92, 
    0.94, 0.91, 0.91, 0.92, 0.9, 0.93, 0.95, 0.94, 0.98, 0.96, 0.97, 0.97, 
    0.96, 0.95, 0.96, 0.97, 0.97, 0.97, 0.96, 0.97, 0.96, 0.95, 0.95, 0.97, 
    0.94, 0.94, 0.95, 0.96, 0.94, 0.96, 0.96, 0.97, 0.95, 0.97, 0.97, 0.98, 
    0.96, 0.95, 0.95, 0.97, 0.97, 0.98, 0.96, 0.95, 0.95, 0.95, 0.95, 0.96, 
    0.96, 0.96, 0.96, 0.95, 0.9, 0.88, 0.96, 0.97, 0.95, 0.95, 0.95, 1, 0.96, 
    0.96, 0.95, 0.96, 0.92, 0.88, 0.86, 0.93, 0.9, 0.87, 0.91, 0.86, 0.9, 
    0.88, 0.87, 0.86, 0.86, 0.86, 0.87, 0.93, 0.91, 0.88, 0.87, 0.88, 0.89, 
    0.89, 0.9, 0.9, 0.88, 0.87, 0.83, 0.79, 0.85, 0.86, 0.84, 0.9, 0.89, 
    0.91, 0.91, 0.93, 0.95, 0.9, 0.92, 0.93, 0.94, 0.96, 0.95, 0.96, 0.97, 
    0.96, 0.95, 0.94, 0.91, 0.92, 0.91, 0.93, 0.94, 0.94, 0.91, 0.89, 0.91, 
    0.92, 0.92, 0.94, 0.94, 0.94, 0.93, 0.94, 0.88, 0.92, 0.93, 0.94, 0.93, 
    0.91, 0.92, 0.9, 0.92, 0.89, 0.9, 0.89, 0.9, 0.9, 0.86, 0.86, 0.9, 0.88, 
    0.87, 0.85, 0.83, 0.86, 0.82, 0.79, 0.82, 0.82, 0.83, 0.8, 0.76, 0.73, 
    0.83, 0.83, 0.84, 0.8, 0.78, 0.84, 0.86, 0.89, 0.89, 0.89, 0.9, 0.9, 0.9, 
    0.91, 0.87, 0.93, 0.94, 0.95, 0.95, 0.95, 0.97, 0.98, 0.98, 0.97, 0.91, 
    0.94, 0.94, 0.95, 0.96, 0.93, 0.94, 0.94, 0.94, 0.95, 0.9, 0.89, 0.91, 
    0.9, 0.93, 0.91, 0.95, 0.96, 0.97, 0.99, 0.99, 0.98, 0.98, 0.99, 0.99, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 0.98, 
    0.95, 0.93, 0.95, 0.95, 0.95, 0.94, 0.92, 0.92, 0.93, 0.93, 0.9, 0.88, 
    0.87, 0.92, 0.97, 0.97, 0.97, 0.98, 1, 0.99, 0.99, 0.99, 0.99, 0.96, 
    0.97, 0.96, 0.96, 0.98, 0.91, 0.97, 0.97, 0.98, 0.98, 0.96, 0.93, 0.94, 
    0.94, 0.94, 0.92, 0.95, 0.92, 0.93, 0.97, 0.98, 0.98, 0.91, 0.98, 0.98, 
    0.97, 0.94, 0.93, 0.91, 0.9, 0.9, 0.89, 0.88, 0.86, 0.81, 0.83, 0.83, 
    0.79, 0.76, 0.79, 0.75, 0.81, 0.78, 0.81, 0.82, 0.83, 0.82, 0.73, 0.82, 
    0.85, 0.81, 0.79, 0.77, 0.86, 0.92, 0.94, 0.95, 0.86, 0.95, 0.91, 0.91, 
    0.89, 0.8, 0.93, 0.93, 0.95, 0.97, 0.86, 0.95, 0.95, 0.92, 0.91, 0.95, 
    0.92, 0.91, 0.91, 0.89, 0.88, 0.89, 0.89, 0.87, 0.87, 0.88, 0.9, 0.91, 
    0.9, 0.93, 0.95, 0.97, 0.98, 0.98, 0.99, 0.98, 0.91, 0.9, 0.95, 0.93, 
    0.94, 0.97, 0.97, 0.97, 0.98, 0.94, 0.96, 0.94, 0.93, 0.93, 0.91, 0.89, 
    0.91, 0.93, 0.91, 0.94, 0.96, 0.91, 0.92, 0.89, 0.84, 0.92, 0.92, 0.92, 
    0.89, 0.87, 0.79, 0.86, 0.85, 0.79, 0.83, 0.86, 0.84, 0.91, 0.91, 0.89, 
    0.9, 0.82, 0.85, 0.86, 0.89, 0.85, 0.9, 0.88, 0.89, 0.81, 0.87, 0.85, 
    0.9, 0.85, 0.87, 0.91, 0.95, 0.93, 0.91, 0.92, 0.89, 0.88, 0.95, 0.94, 
    0.92, 0.89, 0.91, 0.9, 0.87, 0.93, 0.91, 0.9, 0.89, 0.89, 0.92, 0.92, 
    0.91, 0.91, 0.93, 0.92, 0.93, 0.93, 0.94, 0.97, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.98, 0.96, 0.94, 0.93, 0.91, 0.88, 0.9, 0.92, 0.92, 0.9, 
    0.92, 0.95, 0.96, 0.95, 0.94, 0.97, 0.95, 0.94, 0.95, 0.96, 0.97, 0.98, 
    0.97, 0.96, 0.96, 0.95, 0.96, 0.95, 0.94, 0.94, 0.93, 0.94, 0.89, 0.93, 
    0.95, 0.96, 0.94, 0.96, 0.95, 0.94, 0.93, 0.93, 0.9, 0.92, 0.94, 0.94, 
    0.92, 0.92, 0.94, 0.93, 0.9, 0.94, 0.94, 0.92, 0.9, 0.92, 0.92, 0.87, 
    0.9, 0.93, 0.95, 0.93, 0.95, 0.95, 0.96, 0.95, 0.97, 0.97, 0.96, 0.97, 
    0.92, 0.89, 0.89, 0.88, 0.9, 0.93, 0.91, 0.93, 0.94, 0.93, 0.95, 0.95, 
    0.96, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.98, 0.98, 0.98, 0.95, 0.92, 
    0.94, 0.95, 0.9, 0.83, 0.83, 0.75, 0.93, 0.94, 0.93, 0.97, 0.97, 0.9, 
    0.93, 0.92, 0.92, 0.92, 0.95, 0.96, 0.95, 0.93, 0.92, 0.94, 0.92, 0.9, 
    0.93, 0.93, 0.95, 0.94, 0.95, 0.94, 0.92, 0.9, 0.91, 0.92, 0.92, 0.82, 
    0.84, 0.89, 0.98, 0.96, 0.92, 0.93, 0.96, 0.94, 0.93, 0.89, 0.9, 0.92, 
    0.93, 0.93, 0.93, 0.9, 0.9, 0.89, 0.92, 0.92, 0.87, 0.9, 0.97, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.98, 1, 0.98, 0.9, 0.98, 0.98, 0.98, 0.91, 0.93, 
    0.92, 0.92, 0.92, 0.97, 0.98, 0.97, 0.9, 0.91, 0.94, 0.96, 0.97, 0.98, 
    0.98, 0.98, 0.99, 0.97, 0.97, 0.98, 0.98, 0.95, 0.98, 0.93, 0.92, 0.91, 
    0.91, 0.92, 0.94, 0.96, 0.96, 0.95, 0.94, 0.92, 0.96, 0.95, 0.93, 0.89, 
    0.89, 0.92, 0.97, 0.94, 0.93, 0.96, 0.98, 0.97, 0.97, 0.93, 0.92, 0.89, 
    0.85, 0.83, 0.81, 0.81, 0.79, 0.78, 0.8, 0.84, 0.86, 0.84, 0.83, 0.85, 
    0.85, 0.83, 0.8, 0.8, 0.86, 0.85, 0.8, 0.73, 0.78, 0.78, 0.77, 0.73, 
    0.76, 0.7, 0.64, 0.64, 0.8, 0.66, 0.62, 0.62, 0.63, 0.71, 0.74, 0.81, 
    0.85, 0.8, 0.89, 0.93, 0.94, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 0.93, 
    0.9, 0.88, 0.89, 0.87, 0.88, 0.82, 0.82, 0.82, 0.79, 0.78, 0.79, 0.79, 
    0.83, 0.64, 0.75, 0.81, 0.75, 0.69, 0.7, 0.69, 0.7, 0.81, 0.85, 0.89, 
    0.73, 0.81, 0.85, 0.75, 0.85, 0.81, 0.81, 0.83, 0.85, 0.86, 0.9, 0.88, 
    0.87, 0.89, 0.85, 0.75, 0.87, 0.9, 0.96, 0.96, 0.97, 0.96, 0.93, 0.92, 
    0.93, 0.93, 0.89, 0.86, 0.84, 0.83, 0.87, 0.75, 0.89, 0.87, 0.79, 0.75, 
    0.71, 0.7, 0.75, 0.72, 0.76, 0.75, 0.84, 0.8, 0.88, 0.86, 0.92, 0.88, 
    0.82, 0.84, 0.87, 0.93, 0.9, 0.9, 0.9, 0.92, 0.92, 0.91, 0.91, 0.92, 
    0.92, 0.91, 0.92, 0.91, 0.92, 0.91, 0.92, 0.91, 0.91, 0.91, 0.87, 0.86, 
    0.76, 0.82, 0.71, 0.78, 0.83, 0.82, 0.82, 0.84, 0.79, 0.87, 0.78, 0.83, 
    0.84, 0.88, 0.89, 0.9, 0.88, 0.9, 0.89, 0.87, 0.88, 0.86, 0.86, 0.84, 
    0.87, 0.91, 0.8, 0.88, 0.88, 0.85, 0.76, 0.79, 0.79, 0.79, 0.82, 0.84, 
    0.84, 0.83, 0.87, 0.88, 0.89, 0.89, 0.89, 0.89, 0.87, 0.87, 0.89, 0.9, 
    0.9, 0.92, 0.9, 0.89, 0.88, 0.86, 0.86, 0.8, 0.84, 0.77, 0.77, 0.9, 0.79, 
    0.69, 0.82, 0.84, 0.85, 0.82, 0.88, 0.91, 0.9, 0.89, 0.79, 0.9, 0.93, 
    0.88, 0.91, 0.92, 0.94, 0.95, 0.97, 0.93, 0.95, 0.92, 0.9, 0.92, 0.9, 
    0.91, 0.89, 0.9, 0.91, 0.9, 0.94, 0.92, 0.93, 0.88, 0.94, 0.94, 0.94, 
    0.94, 0.95, 0.94, 0.97, 0.98, 0.98, 0.98, 0.98, 0.95, 0.98, 0.99, 0.97, 
    0.98, 0.98, 0.99, 0.97, 0.99, 0.99, 0.99, 0.99, 0.98, 0.91, 0.97, 0.98, 
    0.97, 0.96, 0.97, 0.97, 0.95, 0.97, 0.96, 0.98, 0.95, 0.97, 0.97, 0.96, 
    0.95, 0.96, 0.97, 0.97, 0.98, 0.95, 0.99, 0.96, 0.92, 0.93, 0.94, 0.95, 
    0.92, 0.87, 0.92, 0.88, 0.93, 0.89, 0.86, 0.93, 0.94, 0.94, 0.95, 0.96, 
    0.94, 0.93, 0.95, 0.96, 0.97, 0.93, 0.92, 0.94, 0.95, 0.92, 0.91, 0.92, 
    0.93, 0.94, 0.93, 0.91, 0.92, 0.93, 1, 0.92, 0.92, 0.86, 0.91, 0.89, 
    0.91, 0.93, 0.97, 0.95, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.93, 0.91, 0.89, 
    0.9, 0.91, 0.9, 0.91, 0.95, 0.91, 0.91, 0.97, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.98, 0.96, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.94, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.94, 0.99, 0.99, 0.93, 
    0.88, 0.85, 0.85, 0.86, 0.85, 0.87, 0.88, 0.9, 0.89, 0.88, 0.89, 0.88, 
    0.91, 0.91, 0.87, 0.87, 0.91, 0.91, 0.91, 0.93, 0.92, 0.89, 0.89, 0.9, 
    0.92, 0.95, 0.92, 0.87, 0.89, 0.9, 0.86, 0.91, 0.87, 0.94, 0.93, 0.96, 
    0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.98, 0.99, 
    0.99, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.99, 0.97, 0.94, 0.92, 0.95, 
    0.95, 0.98, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.96, 0.97, 0.96, 0.97, 0.97, 0.97, 0.97, 0.95, 0.97, 0.96, 
    0.97, 0.96, 0.97, 0.98, 0.95, 0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.94, 0.96, 0.95, 0.95, 0.94, 0.95, 0.97, 0.97, 0.96, 0.97, 0.97, 
    0.97, 0.96, 0.95, 0.94, 0.94, 0.96, 0.96, 0.96, 0.93, 0.92, 0.93, 0.9, 
    0.88, 0.92, 0.87, 0.9, 0.93, 0.93, 0.92, 0.91, 0.9, 0.89, 0.9, 0.91, 
    0.92, 0.92, 0.92, 0.93, 0.95, 0.96, 0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.95, 0.96, 0.98, 0.98, 0.96, 
    0.95, 0.94, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.95, 0.92, 0.92, 0.93, 
    0.96, 0.87, 0.94, 0.87, 0.92, 0.89, 0.89, 0.94, 0.96, 0.98, 0.96, 0.94, 
    0.95, 0.98, 0.98, 0.98, 0.94, 0.95, 0.95, 0.94, 0.97, 0.97, 0.97, 0.94, 
    0.94, 0.92, 0.89, 0.91, 0.89, 0.94, 0.9, 0.97, 0.96, 0.92, 0.92, 0.86, 
    0.85, 0.88, 0.97, 0.95, 0.97, 0.97, 0.99, 0.98, 0.98, 0.95, 0.93, 0.96, 
    0.95, 0.92, 0.91, 0.89, 0.91, 0.9, 0.86, 0.83, 0.86, 0.87, 0.88, 0.87, 
    0.88, 0.9, 0.95, 0.98, 0.99, 0.95, 0.97, 0.98, 0.95, 0.94, 0.94, 0.96, 
    0.98, 0.98, 0.98, 0.98, 0.99, 0.96, 0.91, 0.87, 0.89, 0.82, 0.92, 0.8, 
    0.87, 0.87, 0.9, 0.91, 0.87, 0.83, 0.86, 0.91, 0.98, 0.94, 0.91, 0.86, 
    0.86, 0.85, 0.86, 0.87, 0.9, 0.89, 0.92, 0.94, 0.95, 0.93, 0.95, 0.96, 
    0.96, 0.96, 0.96, 0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.98, 0.95, 0.92, 
    0.91, 0.9, 0.9, 0.85, 0.86, 0.84, 0.85, 0.89, 0.87, 0.78, 0.83, 0.79, 
    0.77, 0.77, 0.92, 0.88, 0.96, 0.96, 0.94, 0.96, 0.97, 0.98, 0.92, 0.93, 
    0.93, 0.91, 0.89, 0.91, 0.85, 0.9, 0.85, 0.84, 0.86, 0.84, 0.86, 0.87, 
    0.88, 0.88, 0.92, 0.96, 0.9, 0.95, 0.95, 0.94, 0.93, 0.97, 0.96, 0.88, 
    0.96, 0.9, 0.91, 0.89, 0.88, 0.89, 0.89, 0.87, 0.88, 0.9, 0.92, 0.91, 
    0.89, 0.89, 0.9, 0.9, 0.89, 0.89, 0.89, 0.92, 0.91, 0.9, 0.92, 0.92, 
    0.89, 0.89, 0.91, 0.94, 0.93, 0.95, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.98, 0.97, 0.95, 0.94, 0.93, 0.94, 0.97, 0.96, 0.97, 0.99, 0.99, 
    0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.97, 0.95, 0.92, 0.92, 0.97, 0.98, 0.96, 0.96, 0.94, 0.96, 0.98, 
    0.98, 0.97, 0.93, 0.92, 0.91, 0.91, 0.92, 0.93, 0.92, 0.94, 0.9, 0.88, 
    0.86, 0.83, 0.9, 0.9, 0.88, 0.9, 0.87, 0.85, 0.87, 0.93, 0.95, 0.92, 
    0.87, 0.88, 0.93, 0.93, 0.92, 0.87, 0.94, 0.97, 0.91, 0.89, 0.91, 0.9, 
    0.92, 0.9, 0.88, 0.89, 0.87, 0.79, 0.91, 0.93, 0.76, 0.7, 0.72, 0.81, 
    0.87, 0.71, 0.8, 0.79, 0.78, 0.78, 0.8, 0.78, 0.79, 0.75, 0.71, 0.71, 
    0.74, 0.69, 0.77, 0.76, 0.75, 0.76, 0.85, 0.94, 0.89, 0.87, 0.86, 0.88, 
    0.87, 0.89, 0.9, 0.9, 0.89, 0.92, 0.94, 0.97, 0.89, 0.9, 0.89, 0.85, 
    0.84, 0.85, 0.9, 0.84, 0.8, 0.83, 0.81, 0.83, 0.88, 0.89, 0.96, 0.96, 
    0.94, 0.97, 0.98, 0.99, 0.99, 0.99, 0.97, 0.93, 0.89, 0.9, 0.91, 0.89, 
    0.9, 0.89, 0.9, 0.9, 0.91, 0.91, 0.93, 0.94, 0.94, 0.95, 0.91, 0.9, 0.91, 
    0.94, 0.96, 0.94, 0.92, 0.9, 0.87, 0.85, 0.88, 0.89, 0.92, 0.92, 0.88, 
    0.86, 1, 0.85, 0.83, 0.81, 0.84, 0.85, 1, 0.88, 0.9, 0.89, 0.91, 0.95, 
    0.91, 0.9, 0.94, 0.96, 0.97, 0.96, 0.95, 0.87, 0.86, 0.88, 0.86, 0.87, 
    0.77, 0.72, 0.82, 0.76, 0.78, 0.77, 0.78, 0.79, 0.76, 0.8, 0.76, 0.75, 
    0.86, 0.94, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.97, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.94, 0.95, 0.94, 0.95, 0.95, 0.98, 
    0.99, 0.99, 0.98, 0.95, 0.98, 0.84, 0.89, 0.86, 0.86, 0.85, 0.87, 0.88, 
    0.91, 0.96, 0.99, 0.99, 0.99, 0.99, 0.96, 0.95, 0.9, 0.91, 0.97, 0.95, 
    0.96, 0.9, 0.97, 0.88, 0.83, 0.79, 0.77, 0.76, 0.87, 0.84, 0.9, 0.92, 
    0.93, 0.95, 0.97, 0.95, 0.99, 0.99, 0.99, 0.96, 0.95, 0.98, 0.89, 0.86, 
    0.85, 0.87, 0.86, 0.82, 0.86, 0.91, 0.9, 0.9, 0.91, 0.88, 0.86, 0.88, 
    0.91, 0.93, 0.96, 0.93, 0.93, 0.96, 0.96, 0.98, 0.99, 0.99, 0.97, 0.96, 
    0.95, 0.94, 0.91, 0.91, 0.9, 0.87, 0.87, 0.86, 0.9, 0.92, 0.92, 0.89, 
    0.89, 0.9, 0.9, 0.85, 0.85, 0.88, 0.92, 0.91, 0.91, 0.85, 0.86, 0.86, 
    0.85, 0.84, 0.84, 0.82, 0.84, 0.86, 0.89, 0.91, 0.93, 0.89, 0.93, 0.86, 
    0.94, 0.91, 0.91, 0.84, 0.82, 0.77, 0.79, 0.8, 0.78, 0.78, 0.82, 0.76, 
    0.87, 0.8, 0.78, 0.71, 0.76, 0.75, 0.78, 0.79, 0.81, 0.84, 0.85, 0.87, 
    0.85, 0.84, 0.83, 0.83, 0.78, 0.77, 0.69, 0.72, 0.79, 0.83, 0.82, 0.81, 
    0.76, 0.79, 0.8, 0.83, 0.82, 0.91, 0.89, 0.88, 0.95, 0.97, 0.95, 0.95, 
    0.96, 0.95, 0.92, 0.92, 0.91, 0.88, 0.83, 0.84, 0.85, 0.85, 0.86, 0.84, 
    0.85, 0.83, 0.83, 0.84, 0.83, 0.82, 0.84, 0.9, 0.86, 0.8, 0.85, 0.8, 
    0.81, 0.92, 0.87, 0.9, 0.92, 0.89, 0.94, 0.92, 0.91, 0.89, 0.85, 0.85, 
    0.8, 0.89, 0.91, 0.85, 0.84, 0.88, 0.89, 0.91, 0.9, 0.91, 0.9, 0.91, 0.9, 
    0.88, 0.83, 0.87, 0.89, 0.9, 0.94, 0.95, 0.93, 0.95, 0.96, 0.95, 0.95, 
    0.95, 0.96, 0.97, 0.97, 0.97, 0.93, 0.89, 0.95, 0.96, 0.96, 0.95, 0.96, 
    0.96, 0.96, 0.9, 0.94, 0.96, 0.94, 0.96, 0.96, 0.95, 0.94, 0.95, 0.94, 
    0.93, 0.94, 0.95, 0.93, 0.87, 0.89, 0.9, 0.91, 0.95, 0.97, 0.97, 0.97, 
    0.98, 0.98, 0.97, 0.97, 0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 
    0.95, 0.96, 0.96, 0.97, 0.98, 0.93, 0.96, 0.98, 0.98, 0.98, 0.96, 0.94, 
    0.96, 0.96, 0.88, 0.86, 0.87, 0.87, 0.89, 0.86, 0.88, 0.85, 0.84, 0.84, 
    0.84, 0.82, 0.81, 0.83, 0.83, 0.85, 0.83, 0.78, 0.83, 0.85, 0.81, 0.81, 
    0.8, 0.79, 0.75, 0.73, 0.78, 0.78, 0.8, 0.93, 0.97, 0.9, 0.84, 0.84, 
    0.85, 0.85, 0.89, 0.93, 0.91, 0.99, 0.89, 0.89, 0.9, 0.93, 0.95, 0.96, 
    0.98, 0.98, 0.98, 0.99, 0.99, 0.96, 0.98, 0.99, 0.96, 0.95, 0.95, 0.93, 
    0.91, 0.89, 0.92, 0.96, 0.97, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 0.98, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.96, 0.94, 
    0.89, 0.92, 0.87, 0.86, 0.81, 0.77, 0.79, 0.72, 0.73, 0.77, 0.8, 0.82, 
    0.88, 0.9, 0.94, 0.94, 0.94, 0.92, 0.87, 0.9, 0.91, 0.89, 0.84, 0.82, 
    0.76, 0.66, 0.84, 0.61, 0.62, 0.62, 0.64, 0.62, 0.62, 0.72, 0.77, 0.82, 
    0.83, 0.87, 0.88, 0.83, 0.82, 0.93, 0.94, 0.84, 0.79, 0.75, 0.71, 0.68, 
    0.68, 0.71, 0.79, 0.95, 0.84, 0.84, 0.83, 0.85, 0.85, 0.87, 0.88, 0.85, 
    0.88, 0.92, 0.95, 0.97, 0.98, 0.98, 0.9, 0.91, 0.95, 0.97, 0.97, 0.93, 
    0.91, 0.9, 0.91, 0.91, 0.94, 0.95, 0.96, 0.98, 0.98, 0.98, 0.98, 0.89, 
    0.93, 0.95, 0.91, 0.92, 0.95, 0.95, 0.87, 0.95, 0.88, 0.88, 0.87, 0.87, 
    0.86, 0.84, 0.86, 0.85, 0.92, 0.97, 0.9, 0.94, 0.96, 0.91, 0.96, 0.98, 
    0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 0.98, 0.99, 0.99, 0.99, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.97, 0.89, 0.89, 0.97, 
    0.98, 0.95, 0.93, 0.92, 0.93, 0.93, 0.93, 0.93, 0.91, 0.86, 0.85, 0.87, 
    0.89, 0.87, 0.88, 0.86, 0.87, 0.87, 0.88, 0.9, 0.92, 0.95, 0.96, 0.98, 
    0.98, 0.97, 0.96, 0.97, 0.98, 0.98, 0.99, 0.98, 0.98, 0.98, 0.94, 0.86, 
    0.84, 0.85, 0.85, 0.89, 0.92, 0.94, 0.94, 0.92, 0.91, 0.93, 0.91, 0.89, 
    0.93, 0.92, 0.91, 0.92, 0.95, 0.9, 0.92, 0.91, 0.84, 0.89, 0.85, 0.86, 
    0.84, 0.81, 0.86, 0.83, 0.84, 0.83, 0.75, 0.84, 0.96, 0.82, 0.71, 0.8, 
    0.83, 0.95, 0.97, 0.98, 0.98, 0.97, 0.96, 0.96, 0.95, 0.95, 0.94, 0.95, 
    0.95, 0.95, 0.98, 0.97, 0.96, 0.94, 0.96, 0.94, 0.93, 0.94, 0.94, 0.92, 
    0.97, 0.96, 0.98, 0.99, 0.99, 0.99, 0.95, 0.92, 0.92, 0.97, 0.98, 0.98, 
    0.98, 0.96, 0.96, 0.91, 0.98, 0.97, 0.98, 0.99, 0.97, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 1, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 
    0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.96, 0.96, 0.98, 0.99, 
    0.99, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.94, 0.94, 0.95, 0.94, 0.95, 
    0.92, 0.88, 0.77, 0.79, 0.79, 0.79, 0.78, 0.77, 0.78, 0.75, 0.75, 0.71, 
    0.68, 0.72, 0.7, 0.7, 0.74, 0.77, 0.83, 0.84, 0.88, 0.89, 0.92, 0.92, 
    0.94, 0.96, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 
    0.98, 0.96, 0.95, 0.93, 0.92, 0.93, 0.94, 0.96, 0.96, 0.97, 0.98, 0.96, 
    0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.94, 0.9, 0.87, 0.9, 0.89, 0.9, 0.84, 0.82, 0.92, 
    0.92, 0.92, 0.91, 0.92, 0.9, 0.89, 0.9, 0.92, 0.94, 0.95, 0.94, 0.97, 
    0.95, 0.93, 0.86, 0.85, 0.84, 0.91, 0.83, 0.83, 0.83, 0.91, 0.88, 0.84, 
    0.86, 0.84, 0.85, 0.85, 0.83, 0.85, 0.87, 0.88, 0.89, 0.92, 0.93, 0.94, 
    0.94, 0.93, 0.93, 0.94, 0.95, 0.98, 0.99, 0.99, 0.99, 0.97, 0.97, 0.97, 
    0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.91, 0.89, 0.89, 0.9, 0.93, 0.96, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.92, 0.86, 0.91, 
    0.91, 0.9, 0.94, 0.95, 0.98, 0.97, 0.94, 0.91, 0.87, 0.85, 0.84, 0.83, 
    0.84, 0.83, 0.84, 0.82, 0.81, 0.84, 0.93, 0.92, 0.97, 0.98, 0.97, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.97, 0.94, 0.93, 0.94, 0.9, 
    0.85, 0.77, 0.85, 0.83, 0.84, 0.89, 0.7, 0.71, 0.73, 0.82, 0.83, 0.84, 
    0.84, 0.86, 0.89, 0.91, 0.92, 0.91, 0.91, 0.9, 0.9, 0.89, 0.92, 0.97, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.95, 0.94, 0.94, 0.96, 0.96, 0.93, 0.96, 
    0.96, 0.96, 0.9, 0.91, 0.95, 0.87, 0.87, 0.92, 0.92, 0.98, 0.98, 0.99, 
    0.99, 0.97, 0.95, 0.95, 0.97, 0.97, 0.96, 0.95, 0.94, 0.94, 0.95, 0.94, 
    0.94, 0.95, 0.95, 0.95, 0.96, 0.97, 0.97, 0.99, 0.99, 0.99, 0.98, 0.95, 
    0.93, 0.93, 0.94, 0.95, 0.96, 0.97, 0.95, 0.98, 0.97, 0.97, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 
    0.99, 0.99, 1, 1, 0.98, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 
    0.99, 0.99, 0.97, 0.95, 0.93, 0.9, 0.9, 0.87, 0.85, 0.83, 0.83, 0.85, 
    0.86, 0.85, 0.86, 0.86, 0.9, 0.89, 0.91, 0.91, 0.91, 0.91, 0.92, 0.94, 
    0.94, 0.93, 0.92, 0.94, 0.95, 0.95, 0.94, 0.95, 0.95, 0.96, 0.95, 0.97, 
    0.98, 0.98, 0.95, 0.98, 0.97, 0.97, 0.98, 0.96, 0.96, 0.98, 0.98, 0.99, 
    0.99, 0.98, 0.97, 0.98, 0.95, 0.98, 0.98, 0.96, 0.98, 0.98, 0.97, 0.96, 
    0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 
    0.97, 0.97, 0.98, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 
    0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.96, 0.98, 0.95, 0.98, 0.96, 
    0.94, 0.97, 0.96, 0.95, 0.97, 0.95, 0.91, 0.89, 0.85, 0.85, 0.84, 0.83, 
    0.83, 0.86, 0.82, 0.79, 0.78, 0.76, 0.71, 0.72, 0.71, 0.73, 0.73, 0.7, 
    0.69, 0.67, 0.69, 0.64, 0.66, 0.64, 0.7, 0.7, 0.72, 0.71, 0.76, 0.75, 
    0.8, 0.8, 0.81, 0.93, 0.95, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.93, 0.97, 0.99, 0.97, 0.97, 
    0.86, 0.76, 0.8, 0.76, 0.76, 0.75, 0.75, 0.77, 0.76, 0.77, 0.77, 0.82, 
    0.82, 0.84, 0.84, 0.84, 0.85, 0.81, 0.83, 0.86, 0.89, 0.9, 0.93, 0.94, 
    0.93, 0.9, 0.89, 0.91, 0.96, 0.96, 0.96, 0.96, 0.95, 0.92, 0.92, 0.93, 
    0.93, 0.92, 0.92, 0.92, 0.89, 0.84, 0.93, 0.83, 0.83, 0.85, 0.87, 0.82, 
    0.87, 0.87, 0.83, 0.82, 0.82, 0.83, 0.86, 0.84, 0.86, 0.82, 0.73, 0.72, 
    0.77, 0.79, 0.77, 0.78, 0.79, 0.76, 0.8, 0.82, 0.83, 0.86, 0.82, 0.84, 
    0.83, 0.86, 0.85, 0.88, 0.83, 0.86, 0.86, 0.88, 0.88, 0.88, 0.93, 0.89, 
    0.88, 0.87, 0.87, 0.91, 0.95, 0.96, 0.98, 0.99, 0.99, 0.99, 0.98, 0.97, 
    0.83, 0.86, 0.9, 0.92, 0.92, 0.94, 0.93, 0.92, 0.87, 0.88, 0.85, 0.88, 
    0.9, 0.9, 0.89, 0.86, 0.9, 0.91, 0.89, 0.91, 0.84, 0.87, 0.88, 0.84, 
    0.82, 0.81, 0.83, 0.84, 0.83, 0.85, 0.86, 0.86, 0.89, 0.87, 0.89, 0.91, 
    0.9, 0.91, 0.89, 0.86, 0.87, 0.9, 0.93, 0.94, 0.96, 0.95, 0.94, 0.93, 
    0.91, 0.93, 0.89, 0.89, 0.89, 0.94, 0.93, 0.89, 0.87, 0.87, 0.86, 0.89, 
    0.93, 0.95, 0.94, 0.93, 0.91, 0.9, 0.9, 0.94, 0.92, 0.92, 0.92, 0.92, 
    0.93, 0.92, 0.92, 0.91, 0.95, 0.95, 0.93, 0.93, 0.91, 0.89, 0.94, 0.97, 
    0.97, 0.98, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.96, 0.94, 0.93, 0.94, 0.94, 0.95, 0.98, 0.99, 0.98, 0.98, 0.96, 
    0.94, 0.95, 0.97, 0.99, 0.98, 0.96, 0.96, 0.97, 0.96, 0.95, 0.94, 0.91, 
    0.94, 0.97, 0.98, 0.94, 0.94, 0.94, 0.98, 0.94, 0.93, 0.98, 0.99, 0.96, 
    0.83, 0.72, 0.82, 0.8, 0.8, 0.79, 0.87, 0.89, 0.87, 0.84, 0.81, 0.88, 
    0.9, 0.91, 0.89, 0.9, 0.9, 0.87, 0.88, 0.86, 0.86, 0.89, 0.87, 0.82, 
    0.82, 0.82, 0.79, 0.81, 0.76, 0.71, 0.72, 0.74, 0.79, 0.8, 0.81, 0.84, 
    0.85, 0.87, 0.85, 0.78, 0.77, 0.77, 0.78, 0.77, 0.78, 0.77, 0.74, 0.8, 
    0.78, 0.73, 0.8, 0.82, 0.82, 0.83, 0.84, 0.88, 0.94, 0.96, 0.98, 0.99, 1, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.95, 
    0.93, 0.89, 0.83, 0.84, 0.77, 0.81, 0.83, 0.86, 0.86, 0.88, 0.88, 0.91, 
    0.93, 0.94, 0.94, 0.94, 0.94, 0.96, 0.93, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.96, 0.94, 0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 0.96, 0.96, 0.96, 0.97, 
    0.91, 0.9, 0.89, 0.89, 0.88, 0.86, 0.91, 0.9, 0.9, 0.91, 0.92, 0.92, 
    0.92, 0.91, 0.93, 0.93, 0.95, 0.96, 0.93, 0.93, 0.92, 0.96, 0.93, 0.9, 
    0.91, 0.91, 0.93, 0.93, 0.93, 0.93, 0.91, 0.91, 0.92, 0.91, 0.93, 0.92, 
    0.93, 0.9, 0.93, 0.92, 0.93, 0.93, 0.96, 0.92, 0.89, 0.89, 0.87, 0.86, 
    0.88, 0.9, 0.87, 0.85, 0.87, 0.86, 0.82, 0.81, 0.79, 0.83, 0.81, 0.78, 
    0.7, 0.75, 0.69, 0.68, 0.67, 0.71, 0.71, 0.7, 0.69, 0.75, 0.74, 0.73, 
    0.75, 0.76, 0.78, 0.77, 0.8, 0.8, 0.83, 0.86, 0.9, 0.94, 0.92, 0.92, 
    0.93, 0.96, 0.98, 0.99, 0.95, 0.95, 0.95, 0.94, 0.96, 0.95, 0.95, 0.92, 
    0.95, 0.9, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.97, 0.94, 0.91, 
    0.95, 0.96, 0.97, 0.94, 0.85, 0.83, 0.79, 0.78, 0.88, 0.9, 0.92, 0.97, 
    0.98, 0.99, 0.99, 0.97, 0.94, 0.88, 0.88, 0.94, 0.95, 0.96, 0.94, 0.92, 
    0.94, 0.96, 0.92, 0.92, 0.91, 0.9, 0.86, 0.9, 0.89, 0.85, 0.83, 0.89, 
    0.92, 0.91, 0.92, 0.93, 0.95, 0.95, 0.96, 0.95, 0.96, 0.94, 0.89, 0.9, 
    0.97, 0.94, 0.94, 0.94, 0.91, 0.94, 0.93, 0.94, 0.92, 0.95, 0.94, 0.94, 
    0.96, 0.98, 0.98, 0.99, 0.97, 0.94, 0.94, 0.95, 0.96, 0.98, 0.97, 0.98, 
    0.98, 0.98, 0.97, 0.97, 0.94, 0.93, 0.92, 0.92, 0.88, 0.85, 0.89, 0.87, 
    0.84, 0.85, 0.86, 0.86, 0.85, 0.86, 0.88, 0.91, 0.92, 0.87, 0.85, 0.89, 
    0.88, 0.89, 0.88, 0.87, 0.89, 0.89, 0.88, 0.91, 0.91, 0.92, 0.91, 0.9, 
    0.88, 0.86, 0.85, 0.84, 0.84, 0.84, 0.83, 0.79, 0.78, 0.73, 0.71, 0.79, 
    0.85, 0.79, 0.73, 0.73, 0.84, 0.88, 0.82, 0.85, 0.85, 0.89, 0.88, 0.84, 
    0.86, 0.85, 0.85, 0.8, 0.81, 0.82, 0.84, 0.83, 0.82, 0.81, 0.82, 0.82, 
    0.82, 0.82, 0.8, 0.84, 0.86, 0.83, 0.83, 0.85, 0.85, 0.87, 0.86, 0.87, 
    0.9, 0.9, 0.86, 0.86, 0.86, 0.81, 0.8, 0.8, 0.82, 0.77, 0.77, 0.79, 0.8, 
    0.77, 0.74, 0.78, 0.78, 0.71, 0.69, 0.69, 0.78, 0.7, 0.7, 0.69, 0.77, 
    0.74, 0.76, 0.72, 0.77, 0.76, 0.77, 0.76, 0.8, 0.81, 0.79, 0.82, 0.8, 
    0.83, 0.83, 0.85, 0.86, 0.85, 0.85, 0.86, 0.85, 0.84, 0.83, 0.83, 0.8, 
    0.81, 0.82, 0.82, 0.83, 0.83, 0.89, 0.9, 0.92, 0.91, 0.87, 0.87, 0.8, 
    0.81, 0.81, 0.78, 0.69, 0.7, 0.72, 0.82, 0.93, 0.91, 0.92, 0.91, 0.86, 
    0.84, 0.83, 0.85, 0.88, 0.82, 0.84, 0.83, 0.87, 0.89, 0.92, 0.9, 0.65, 
    0.66, 0.73, 0.68, 0.71, 0.73, 0.71, 0.72, 0.71, 0.73, 0.74, 0.78, 0.82, 
    0.87, 0.88, 0.86, 0.86, 0.85, 0.86, 0.88, 0.87, 0.9, 0.9, 0.91, 0.89, 
    0.91, 0.94, 0.92, 0.94, 0.93, 0.96, 0.96, 0.96, 0.92, 0.91, 0.96, 0.97, 
    0.97, 0.94, 0.93, 0.88, 0.87, 0.89, 0.9, 0.89, 0.87, 0.87, 0.86, 0.84, 
    0.83, 0.83, 0.81, 0.8, 0.81, 0.82, 0.8, 0.79, 0.8, 0.82, 0.83, 0.78, 
    0.77, 0.79, 0.72, 0.73, 0.76, 0.82, 0.82, 0.86, 0.88, 0.89, 0.9, 0.93, 
    0.92, 0.89, 0.89, 0.89, 0.89, 0.91, 0.91, 0.91, 0.92, 0.93, 0.93, 0.94, 
    0.93, 0.94, 0.94, 0.93, 0.92, 0.91, 0.93, 0.92, 0.93, 0.93, 0.92, 0.9, 
    0.9, 0.91, 0.91, 0.95, 0.93, 0.91, 0.91, 0.9, 0.9, 0.91, 0.9, 0.91, 0.91, 
    0.86, 0.87, 0.91, 0.93, 0.78, 0.78, 0.77, 0.7, 0.72, 0.74, 0.77, 0.79, 
    0.82, 0.79, 0.79, 0.76, 0.77, 0.77, 0.79, 0.8, 0.78, 0.8, 0.78, 0.78, 
    0.77, 0.79, 0.84, 0.84, 0.86, 0.88, 0.88, 0.87, 0.86, 0.88, 0.88, 0.91, 
    0.93, 0.92, 0.89, 0.9, 0.87, 0.82, 0.81, 0.83, 0.82, 0.87, 0.88, 0.89, 
    0.9, 0.93, 0.94, 0.95, 0.95, 0.94, 0.88, 0.88, 0.84, 0.84, 0.84, 0.78, 
    0.79, 0.77, 0.83, 0.9, 0.85, 0.76, 0.79, 0.74, 0.8, 0.91, 0.87, 0.88, 
    0.91, 0.86, 0.95, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.96, 0.98, 0.98, 0.99, 0.99, 0.98, 0.97, 0.97, 0.98, 0.99, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 
    0.95, 0.9, 0.94, 0.96, 0.98, 0.98, 0.99, 0.98, 0.97, 0.98, 0.98, 0.96, 
    0.94, 0.94, 0.95, 0.96, 0.96, 0.96, 0.97, 0.98, 0.98, 0.97, 0.92, 0.9, 
    0.89, 0.87, 0.85, 0.86, 0.89, 0.91, 0.91, 0.91, 0.91, 0.91, 0.92, 0.92, 
    0.9, 0.91, 0.93, 0.94, 0.94, 0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.96, 0.97, 0.97, 0.96, 0.96, 0.96, 0.97, 0.97, 0.98, 0.98, 0.97, 
    0.97, 0.97, 0.97, 0.95, 0.94, 0.89, 0.89, 0.91, 0.94, 0.94, 0.97, 0.95, 
    0.92, 0.9, 0.9, 0.9, 0.94, 0.98, 0.99, 0.93, 0.91, 0.97, 0.99, 0.99, 
    0.99, 0.98, 0.98, 0.99, 0.99, 0.92, 0.97, 0.97, 0.95, 0.95, 0.97, 0.97, 
    0.96, 0.97, 0.96, 0.95, 0.94, 0.93, 0.93, 0.9, 0.94, 0.94, 0.95, 0.96, 
    0.96, 0.95, 0.93, 0.92, 0.9, 0.89, 0.88, 0.9, 0.89, 0.91, 0.88, 0.8, 
    0.83, 0.82, 0.81, 0.79, 0.86, 0.89, 0.91, 0.9, 0.89, 0.89, 0.87, 0.88, 
    0.89, 0.87, 0.88, 0.91, 0.9, 0.85, 0.88, 0.84, 0.86, 0.9, 0.87, 0.91, 
    0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.91, 0.88, 0.86, 0.87, 
    0.84, 0.83, 0.84, 0.84, 0.88, 0.87, 0.87, 0.87, 0.87, 0.81, 0.84, 0.82, 
    0.78, 0.79, 0.83, 0.81, 0.8, 0.81, 0.83, 0.77, 0.85, 0.84, 0.81, 0.79, 
    0.92, 0.91, 0.84, 0.81, 0.78, 0.83, 0.85, 0.69, 0.7, 0.72, 0.73, 0.78, 
    0.8, 0.69, 0.71, 0.81, 0.75, 0.7, 0.76, 0.69, 0.76, 0.77, 0.73, 0.82, 
    0.81, 0.79, 0.83, 0.81, 0.81, 0.83, 0.77, 0.69, 0.7, 0.77, 0.79, 0.82, 
    0.75, 0.72, 0.66, 0.64, 0.62, 0.7, 0.67, 0.71, 0.67, 0.71, 0.7, 0.73, 
    0.7, 0.69, 0.71, 0.72, 0.7, 0.69, 0.69, 0.73, 0.92, 0.92, 0.96, 0.79, 
    0.84, 0.89, 0.86, 0.85, 0.76, 0.75, 0.7, 0.71, 0.72, 0.71, 0.72, 0.72, 
    0.73, 0.75, 0.78, 0.81, 0.8, 0.78, 0.74, 0.7, 0.67, 0.71, 0.71, 0.67, 
    0.83, 0.82, 0.67, 0.71, 0.66, 0.68, 0.75, 0.74, 0.68, 0.82, 0.75, 0.83, 
    0.85, 0.75, 0.72, 0.81, 0.8, 0.76, 0.76, 0.77, 0.83, 0.77, 0.7, 0.84, 
    0.84, 0.76, 0.75, 0.86, 0.8, 0.9, 0.85, 0.8, 0.83, 0.78, 0.59, 0.71, 
    0.78, 0.72, 0.78, 0.66, 0.7, 0.8, 0.89, 0.92, 0.94, 0.82, 0.78, 0.76, 
    0.73, 0.72, 0.74, 0.8, 0.79, 0.76, 0.7, 0.68, 0.77, 0.7, 0.68, 0.77, 0.8, 
    0.74, 0.74, 0.76, 0.72, 0.71, 0.73, 0.81, 0.78, 0.78, 0.79, 0.62, 0.69, 
    0.65, 0.65, 0.63, 0.61, 0.62, 0.59, 0.59, 0.6, 0.69, 0.83, 0.86, 0.88, 
    0.7, 0.67, 0.69, 0.91, 0.74, 0.69, 0.74, 0.68, 0.83, 0.86, 0.74, 0.74, 
    0.69, 0.83, 0.84, 0.82, 0.69, 0.71, 0.69, 0.85, 0.88, 0.7, 0.72, 0.73, 
    0.68, 0.68, 0.79, 0.9, 0.83, 0.83, 0.9, 0.8, 0.8, 0.72, 0.74, 0.74, 0.79, 
    0.88, 0.78, 0.73, 0.76, 0.79, 0.78, 0.78, 0.78, 0.7, 0.78, 0.71, 0.68, 
    0.78, 0.79, 0.75, 0.79, 0.79, 0.75, 0.77, 0.67, 0.76, 0.78, 0.69, 0.7, 
    0.72, 0.69, 0.61, 0.62, 0.65, 0.66, 0.69, 0.7, 0.72, 0.7, 0.65, 0.65, 
    0.64, 0.61, 0.58, 0.56, 0.57, 0.6, 0.61, 0.62, 0.62, 0.61, 0.52, 0.54, 
    0.61, 0.58, 0.61, 0.6, 0.57, 0.69, 0.61, 0.77, 0.67, 0.64, 0.66, 0.67, 
    0.66, 0.67, 0.8, 0.62, 0.66, 0.56, 0.52, 0.65, 0.54, 0.57, 0.56, 0.54, 
    0.61, 0.74, 0.68, 0.53, 0.59, 0.6, 0.73, 0.61, 0.69, 0.68, 0.76, 0.74, 
    0.76, 0.78, 0.79, 0.86, 0.86, 0.83, 0.82, 0.85, 0.86, 0.86, 0.82, 0.83, 
    0.82, 0.78, 0.78, 0.79, 0.81, 0.81, 0.82, 0.83, 0.84, 0.84, 0.86, 0.88, 
    0.88, 0.87, 0.88, 0.89, 0.91, 0.91, 0.88, 0.85, 0.79, 0.72, 0.73, 0.65, 
    0.77, 0.73, 0.75, 0.84, 0.65, 0.79, 0.84, 0.78, 0.65, 0.61, 0.63, 0.66, 
    0.64, 0.66, 0.64, 0.6, 0.63, 0.62, 0.6, 0.63, 0.65, 0.63, 0.62, 0.64, 
    0.62, 0.6, 0.63, 0.63, 0.6, 0.6, 0.61, 0.6, 0.6, 0.62, 0.62, 0.64, 0.63, 
    0.62, 0.62, 0.65, 0.66, 0.65, 0.67, 0.65, 0.65, 0.68, 0.66, 0.72, 0.73, 
    0.74, 0.74, 0.74, 0.74, 0.73, 0.72, 0.72, 0.73, 0.74, 0.75, 0.74, 0.74, 
    0.74, 0.75, 0.71, 0.68, 0.73, 0.74, 0.63, 0.58, 0.59, 0.62, 0.69, 0.57, 
    0.55, 0.65, 0.77, 0.8, 0.81, 0.8, 0.8, 0.82, 0.83, 0.82, 0.81, 0.79, 
    0.76, 0.75, 0.74, 0.73, 0.74, 0.77, 0.79, 0.81, 0.82, 0.83, 0.81, 0.81, 
    0.8, 0.8, 0.79, 0.78, 0.77, 0.77, 0.75, 0.74, 0.74, 0.73, 0.72, 0.73, 
    0.74, 0.78, 0.8, 0.82, 0.84, 0.84, 0.8, 0.77, 0.74, 0.76, 0.76, 0.75, 
    0.74, 0.74, 0.74, 0.73, 0.74, 0.74, 0.74, 0.73, 0.72, 0.7, 0.74, 0.73, 
    0.72, 0.71, 0.71, 0.72, 0.73, 0.73, 0.73, 0.73, 0.74, 0.75, 0.75, 0.76, 
    0.77, 0.77, 0.76, 0.76, 0.76, 0.76, 0.75, 0.75, 0.73, 0.72, 0.71, 0.7, 
    0.7, 0.7, 0.69, 0.69, 0.7, 0.69, 0.68, 0.69, 0.68, 0.68, 0.71, 0.71, 
    0.71, 0.71, 0.71, 0.72, _, 0.73, 0.72, 0.71, 0.72, 0.75, 0.74, 0.76, 
    0.77, 0.79, 0.81, 0.82, 0.84, 0.86, 0.88, 0.89, 0.9, 0.92, 0.96, 0.96, 
    0.96, 0.97, 0.96, 0.97, 0.96, 0.91, 0.87, 0.84, 0.88, 0.9, 0.83, 0.83, 
    0.84, 0.83, 0.81, 0.79, 0.77, 0.78, 0.79, 0.78, 0.79, 0.8, 0.76, 0.76, 
    0.76, 0.77, 0.78, 0.79, 0.8, 0.74, 0.77, 0.76, 0.84, 0.82, 0.82, 0.88, 
    0.88, 0.89, 0.93, 0.94, 0.95, 0.94, 0.95, 0.94, 0.96, 0.97, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.86, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.92, 0.92, 0.92, 0.96, 0.96, 0.93, 0.93, 0.89, 0.86, 0.86, 0.89, 0.88, 
    0.88, 0.89, 0.89, 0.87, 0.87, 0.87, 0.87, 0.88, 0.87, 0.89, 0.87, 0.87, 
    0.88, 0.87, 0.86, 0.88, 0.87, 0.86, 0.91, 0.9, 0.93, 0.96, 0.97, 0.97, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 
    0.96, 0.96, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.96, 0.94, 0.94, 0.92, 0.93, 
    0.95, 0.96, 0.94, 0.95, 0.96, 0.98, 0.98, 0.96, 0.96, 0.93, 0.93, 0.89, 
    0.95, 0.96, 0.97, 0.97, 0.96, 0.97, 0.98, 0.98, 0.99, 0.98, 0.88, 0.8, 
    0.8, 0.77, 0.79, 0.83, 0.81, 0.73, 0.76, 0.76, 0.8, 0.76, 0.8, 0.88, 
    0.83, 0.83, 0.8, 0.79, 0.86, 0.87, 0.9, 0.91, 0.94, 0.95, 0.95, 0.93, 
    0.95, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.95, 0.94, 0.93, 
    0.97, 0.98, 0.99, 0.99, 0.97, 0.95, 0.94, 0.95, 0.95, 0.93, 0.91, 0.95, 
    0.95, 0.94, 0.93, 0.89, 0.85, 0.84, 0.83, 0.89, 0.92, 0.91, 0.88, 0.9, 
    0.91, 0.96, 0.91, 0.92, 0.91, 0.92, 0.93, 0.93, 0.93, 0.94, 0.93, 0.94, 
    0.93, 0.93, 0.92, 0.92, 0.93, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.91, 
    0.97, 0.97, 0.98, 0.98, 0.97, 0.95, 0.97, 0.97, 0.96, 0.94, 0.92, 0.88, 
    0.84, 0.92, 0.94, 0.94, 0.92, 0.91, 0.96, 0.93, 0.89, 0.94, 0.93, 0.94, 
    0.92, 0.9, 0.94, 0.93, 0.92, 0.91, 0.96, 0.91, 0.86, 0.9, 0.9, 0.89, 
    0.89, 0.91, 0.92, 0.9, 1, 0.9, 0.89, 0.9, 0.89, 0.88, 0.95, 0.94, 0.93, 
    0.93, 0.9, 0.92, 0.92, 0.94, 0.94, 0.93, 0.94, 0.91, 0.91, 0.91, 0.93, 
    0.93, 0.93, 0.93, 0.91, 0.89, 0.89, 0.87, 0.89, 0.86, 0.89, 0.88, 0.87, 
    0.89, 0.89, 0.87, 0.89, 0.88, 0.8, 0.79, 0.83, 0.83, 0.8, 0.76, 0.81, 
    0.77, 0.67, 0.67, 0.69, 0.69, 0.65, 0.65, 0.62, 0.63, 0.64, 0.64, 0.74, 
    0.88, 0.86, 0.81, 0.77, 0.79, 0.75, 0.68, 0.66, 0.7, 0.69, 0.61, 0.67, 
    0.72, 0.69, 0.7, 0.73, 0.82, 0.75, 0.84, 0.8, 0.84, 0.83, 0.89, 0.84, 
    0.83, 0.83, 0.9, 0.91, 0.87, 0.86, 0.85, 0.84, 0.83, 0.91, 0.86, 0.79, 
    0.82, 0.71, 0.87, 0.88, 0.89, 0.88, 0.83, 0.82, 0.86, 0.85, 0.88, 0.73, 
    0.85, 0.79, 0.81, 0.77, 0.73, 0.69, 0.7, 0.73, 0.66, 0.8, 0.86, 0.8, 
    0.73, 0.75, 0.84, 0.83, 0.87, 0.85, 0.86, 0.78, 0.77, 0.86, 0.83, 0.72, 
    0.84, 0.83, 0.82, 0.84, 0.85, 0.76, 0.79, 0.76, 0.75, 0.76, 0.77, 0.82, 
    0.82, 0.78, 0.8, 0.77, 0.74, 0.79, 0.8, 0.78, 0.73, 0.78, 0.76, 0.76, 
    0.79, 0.74, 0.75, 0.76, 0.77, 0.79, 0.77, 0.77, 0.75, 0.75, 0.76, 0.74, 
    0.81, 0.76, 0.78, 0.82, 0.84, 0.81, 0.74, 0.74, 0.72, 0.73, 0.71, 0.7, 
    0.71, 0.67, 0.78, 0.67, 0.77, 0.79, 0.78, 0.8, 0.76, 0.75, 0.77, 0.72, 
    0.74, 0.76, 0.81, 0.82, 0.7, 0.76, 0.65, 0.74, 0.73, 0.69, 0.73, 0.7, 
    0.62, 0.61, 0.66, 0.64, 0.6, 0.62, 0.66, 0.64, 0.63, 0.68, 0.64, 0.63, 
    0.62, 0.64, 0.63, 0.63, 0.61, 0.63, 0.65, 0.6, 0.61, 0.62, 0.61, 0.63, 
    0.64, 0.63, 0.65, 0.64, 0.65, 0.65, 0.69, 0.72, 0.76, 0.76, 0.76, 0.74, 
    0.74, 0.74, 0.71, 0.71, 0.7, 0.73, 0.73, 0.76, 0.72, 0.69, 0.74, 0.93, 
    0.88, 0.81, 0.77, 0.77, 0.8, 0.84, 0.81, 0.77, 0.78, 0.84, 0.86, 0.85, 
    0.77, 0.92, 0.93, 0.83, 0.81, 0.83, 0.88, 0.96, 0.96, 0.93, 0.95, 0.97, 
    0.97, 0.97, 0.96, 0.95, 0.95, 0.9, 0.88, 0.91, 0.9, 0.92, 0.88, 0.85, 
    0.87, 0.86, 0.83, 0.84, 0.81, 0.79, 0.86, 0.75, 0.8, 0.7, 0.82, 0.82, 
    0.78, 0.8, 0.77, 0.84, 0.77, 0.78, 0.81, 0.79, 0.75, 0.75, 0.84, 0.74, 
    0.72, 0.65, 0.69, 0.6, 0.63, 0.62, 0.59, 0.63, 0.67, 0.77, 0.72, 0.67, 
    0.6, 0.63, 0.71, 0.63, 0.56, 0.63, 0.58, 0.75, 0.77, 0.67, 0.59, 0.61, 
    0.72, 0.85, 0.66, 0.62, 0.52, 0.69, 0.66, 0.7, 0.75, 0.73, 0.57, 0.58, 
    0.62, 0.62, 0.69, 0.7, 0.71, 0.7, 0.68, 0.74, 0.74, 0.75, 0.75, 0.72, 
    0.69, 0.71, 0.85, 0.74, 0.82, 0.75, 0.79, 0.81, 0.78, 0.87, 0.85, 0.83, 
    0.85, 0.75, 0.8, 0.85, 0.86, 0.83, 0.86, 0.88, 0.88, 0.83, 0.84, 0.87, 
    0.81, 0.87, 0.87, 0.87, 0.8, 0.81, 0.8, 0.82, 0.83, 0.79, 0.8, 0.77, 
    0.76, 0.79, 0.74, 0.77, 0.68, 0.77, 0.73, 0.71, 0.69, 0.6, 0.63, 0.75, 
    0.74, 0.72, 0.72, 0.73, 0.72, 0.72, 0.74, 0.74, 0.71, 0.71, 0.71, 0.77, 
    0.77, 0.8, 0.81, 0.8, 0.7, 0.72, 0.79, 0.78, 0.78, 0.69, 0.69, 0.71, 
    0.72, 0.75, 0.63, 0.77, 0.67, 0.7, 0.67, 0.75, 0.71, 0.66, 0.75, 0.68, 
    0.59, 0.52, 0.53, 0.62, 0.69, 0.76, 0.7, 0.78, 0.88, 0.81, 0.73, 0.73, 
    0.72, 0.71, 0.65, 0.66, 0.64, 0.63, 0.69, 0.66, 0.66, 0.69, 0.69, 0.72, 
    0.68, 0.68, 0.67, 0.7, 0.61, 0.73, 0.69, 0.56, 0.61, 0.76, 0.81, 0.83, 
    0.8, 0.81, 0.82, 0.76, 0.78, 0.82, 0.82, 0.84, 0.86, 0.85, 0.86, 0.86, 
    0.87, 0.85, 0.84, 0.83, 0.83, 0.84, 0.86, 0.88, 0.92, 0.9, 0.89, 0.87, 
    0.86, 0.85, 0.83, 0.84, 0.81, 0.76, 0.74, 0.72, 0.72, 0.68, 0.78, 0.91, 
    0.72, 0.72, 0.67, 0.69, 0.66, 0.63, 0.64, 0.72, 0.69, 0.77, 0.73, 0.76, 
    0.77, 0.89, 0.89, 0.87, 0.92, 0.91, 0.88, 0.85, 0.94, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.98, 0.99, 0.99, 0.98, 0.92, 0.83, 0.88, 0.88, 0.86, 0.9, 
    0.89, 0.87, 0.85, 0.81, 0.76, 0.8, 0.81, 0.83, 0.88, 0.85, 0.65, 0.69, 
    0.83, 0.81, 0.81, 0.78, 0.77, 0.75, 0.79, 0.71, 0.83, 0.78, 0.78, 0.74, 
    0.83, 0.79, 0.7, 0.67, 0.6, 0.62, 0.67, 0.77, 0.66, 0.82, 0.81, 0.82, 
    0.67, 0.73, 0.79, 0.71, 0.69, 0.69, 0.78, 0.67, 0.52, 0.47, 0.57, 0.57, 
    0.6, 0.64, 0.69, 0.57, 0.53, 0.51, 0.45, 0.81, 0.67, 0.66, 0.72, 0.63, 
    0.61, 0.55, 0.66, 0.71, 0.71, 0.69, 0.83, 0.8, 0.79, 0.86, 0.79, 0.73, 
    0.76, 0.66, 0.64, 0.72, 0.73, 0.59, 0.8, 0.63, 0.56, 0.72, 0.71, 0.64, 
    0.55, 0.57, 0.56, 0.64, 0.76, 0.82, 0.83, 0.89, 0.91, 0.89, 0.85, 0.79, 
    0.74, 0.83, 0.82, 0.79, 0.78, 0.8, 0.8, 0.75, 0.8, 0.84, 0.84, 0.82, 
    0.79, 0.8, 0.78, 0.74, 0.71, 0.7, 0.65, 0.81, 0.87, 0.8, 0.77, 0.71, 
    0.81, 0.88, 0.84, 0.78, 0.77, 0.81, 0.89, 0.8, 0.81, 0.8, 0.75, 0.76, 
    0.77, 0.74, 0.7, 0.67, 0.69, 0.64, 0.65, 0.68, 0.69, 0.72, 0.73, 0.75, 
    0.78, 0.83, 0.84, 0.78, 0.76, 0.76, 0.74, 0.87, 0.85, 0.69, 0.68, 0.66, 
    0.69, 0.73, 0.77, 0.8, 0.8, 0.81, 0.82, 0.85, 0.89, 0.91, 0.81, 0.82, 
    0.82, 0.83, 0.83, 0.87, 0.87, 0.89, 0.9, 0.95, 0.96, 0.93, 0.87, 0.89, 
    0.83, 0.83, 0.85, 0.82, 0.8, 0.84, 0.81, 0.84, 0.82, 0.86, 0.8, 0.82, 
    0.7, 0.73, 0.68, 0.7, 0.83, 0.8, 0.78, 0.85, 0.81, 0.89, 0.85, 0.82, 
    0.88, 0.85, 0.87, 0.81, 0.74, 0.78, 0.68, 0.82, 0.68, 0.62, 0.62, 0.65, 
    0.72, 0.71, 0.85, 0.75, 0.75, 0.82, 0.83, 0.78, 0.73, 0.82, 0.86, 0.81, 
    0.69, 0.81, 0.74, 0.83, 0.73, 0.69, 0.78, 0.83, 0.83, 0.68, 0.66, 0.74, 
    0.63, 0.65, 0.83, 0.69, 0.68, 0.82, 0.78, 0.74, 0.83, 0.79, 0.68, 0.68, 
    0.75, 0.73, 0.76, 0.79, 0.78, 0.85, 0.84, 0.81, 0.8, 0.72, 0.67, 0.69, 
    0.79, 0.84, 0.66, 0.7, 0.7, 0.79, 0.76, 0.68, 0.8, 0.73, 0.76, 0.8, 0.74, 
    0.86, 0.86, 0.82, 0.83, 0.77, 0.8, 0.73, 0.78, 0.65, 0.69, 0.68, 0.66, 
    0.64, 0.67, 0.59, 0.6, 0.67, 0.82, 0.79, 0.69, 0.79, 0.68, 0.66, 0.67, 
    0.81, 0.72, 0.71, 0.73, 0.77, 0.71, 0.68, 0.69, 0.77, 0.71, 0.68, 0.71, 
    0.69, 0.74, 0.76, 0.73, 0.87, 0.86, 0.8, 0.73, 0.76, 0.78, 0.81, 0.87, 
    0.85, 0.79, 0.87, 0.86, 0.89, 0.83, 0.85, 0.81, 0.88, 0.85, 0.76, 0.79, 
    0.83, 0.77, 0.87, 0.85, 0.84, 0.81, 0.79, 0.77, 0.74, 0.79, 0.79, 0.75, 
    0.73, 0.71, 0.8, 0.85, 0.83, 0.83, 0.82, 0.83, 0.8, 0.76, 0.77, 0.78, 
    0.74, 0.76, 0.8, 0.72, 0.7, 0.74, 0.73, 0.76, 0.79, 0.74, 0.72, 0.74, 
    0.72, 0.75, 0.74, 0.8, 0.68, 0.7, 0.73, 0.72, 0.7, 0.69, 0.7, 0.74, 0.73, 
    0.72, 0.72, 0.7, 0.81, 0.67, 0.67, 0.68, 0.7, 0.79, 0.83, 0.87, 0.83, 
    0.9, 0.9, 0.9, 0.9, 0.86, 0.86, 0.87, 0.86, 0.86, 0.86, 0.85, 0.83, 0.84, 
    0.82, 0.85, 0.81, 0.83, 0.82, 0.84, 0.95, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.95, 0.95, 0.94, 0.94, 0.95, 0.97, 0.97, 0.97, 0.99, 0.97, 0.97, 0.95, 
    0.92, 0.92, 0.93, 0.94, 0.92, 0.9, 0.88, 0.84, 0.81, 0.87, 0.9, 0.92, 
    0.93, 0.93, 0.95, 0.95, 0.94, 0.94, 0.99, 0.97, 0.96, 0.97, 0.98, 0.98, 
    0.99, 0.98, 0.94, 0.92, 0.92, 0.9, 0.91, 0.92, 0.94, 0.89, 0.88, 0.89, 
    0.93, 0.95, 0.95, 0.9, 0.93, 0.93, 0.94, 0.91, 0.96, 0.95, 0.95, 0.95, 
    0.85, 0.83, 0.87, 0.87, 0.91, 0.94, 0.95, 0.83, 0.84, 0.86, 0.82, 0.85, 
    0.83, 0.85, 0.85, 0.88, 0.89, 0.89, 0.9, 0.84, 0.85, 0.84, 0.86, 0.9, 
    0.88, 0.9, 0.89, 0.9, 0.89, 0.89, 0.9, 0.97, 0.93, 0.94, 0.91, 0.9, 0.91, 
    0.89, 0.88, 0.92, 0.85, 0.82, 0.83, 0.86, 0.87, 0.91, 0.93, 0.95, 0.95, 
    0.94, 0.93, 0.92, 0.92, 0.88, 0.8, 0.82, 0.87, 0.9, 0.91, 0.89, 0.9, 
    0.89, 0.87, 0.79, 0.75, 0.73, 0.72, 0.72, 0.69, 0.79, 0.85, 0.82, 0.84, 
    0.74, 0.8, 0.77, 0.75, 0.77, 0.73, 0.72, 0.78, 0.81, 0.81, 0.84, 0.79, 
    0.82, 0.8, 0.78, 0.8, 0.8, 0.81, 0.84, 0.8, 0.83, 0.82, 0.81, 0.79, 0.83, 
    0.86, 0.87, 0.87, 0.88, 0.89, 0.84, 0.88, 0.89, 0.9, 0.92, 0.91, 0.91, 
    0.89, 0.9, 0.87, 0.87, 0.87, 0.86, 0.89, 0.74, 0.8, 0.8, 0.82, 0.82, 
    0.82, 0.81, 0.85, 0.84, 0.82, 0.84, 0.87, 0.88, 0.93, 0.96, 0.94, 0.94, 
    0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 0.98, 0.97, 0.89, 0.87, 0.93, 0.89, 
    0.92, 0.9, 0.86, 0.84, 0.8, 0.82, 0.82, 0.85, 0.76, 0.76, 0.73, 0.76, 
    0.78, 0.78, 0.75, 0.76, 0.77, 0.76, 0.78, 0.75, 0.72, 0.74, 0.75, 0.77, 
    0.77, 0.82, 0.8, 0.81, 0.83, 0.75, 0.82, 0.78, 0.81, 0.8, 0.83, 0.85, 
    0.85, 0.78, 0.83, 0.8, 0.76, 0.72, 0.7, 0.76, 0.8, 0.7, 0.76, 0.68, 0.71, 
    0.78, 0.72, 0.75, 0.76, 0.84, 0.77, 0.74, 0.8, 0.78, 0.75, 0.79, 0.77, 
    0.78, 0.79, 0.81, 0.82, 0.82, 0.82, 0.82, 0.81, 0.83, 0.84, 0.84, 0.83, 
    0.83, 0.83, 0.7, 0.72, 0.8, 0.71, 0.78, 0.79, 0.79, 0.76, 0.77, 0.77, 
    0.77, 0.79, 0.83, 0.81, 0.79, 0.79, 0.79, 0.77, 0.79, 0.8, 0.8, 0.78, 
    0.8, 0.79, 0.79, 0.79, 0.73, 0.75, 0.75, 0.77, 0.77, 0.77, 0.77, 0.77, 
    0.8, 0.74, 0.76, 0.81, 0.81, 0.81, 0.81, 0.82, 0.81, 0.79, 0.81, 0.77, 
    0.79, 0.8, 0.79, 0.83, 0.76, 0.73, 0.66, 0.71, 0.72, 0.66, 0.71, 0.67, 
    0.72, 0.68, 0.65, 0.77, 0.63, 0.69, 0.7, 0.72, 0.71, 0.68, 0.68, 0.7, 
    0.69, 0.69, 0.74, 0.72, 0.69, 0.71, 0.74, 0.75, 0.75, 0.76, 0.77, 0.78, 
    0.77, 0.75, 0.75, 0.77, 0.73, 0.79, 0.74, 0.81, 0.87, 0.87, 0.87, 0.87, 
    0.87, 0.87, 0.86, 0.86, 0.87, 0.87, 0.87, 0.86, 0.87, 0.87, 0.88, 0.88, 
    0.88, 0.89, 0.89, 0.9, 0.9, 0.89, 0.88, 0.89, 0.9, 0.9, 0.9, 0.9, 0.9, 
    0.89, 0.89, 0.89, 0.88, 0.89, 0.87, 0.85, 0.84, 0.84, 0.84, 0.84, 0.83, 
    0.82, 0.84, 0.85, 0.83, 0.84, 0.79, 0.8, 0.79, 0.78, 0.78, 0.77, 0.82, 
    0.79, 0.78, 0.78, 0.78, 0.79, 0.81, 0.79, 0.82, 0.82, 0.85, 0.82, 0.82, 
    0.84, 0.83, 0.82, 0.84, 0.84, 0.84, 0.85, 0.85, 0.8, 0.77, 0.75, 0.76, 
    0.77, 0.76, 0.75, 0.76, 0.78, 0.77, 0.75, 0.76, 0.75, 0.77, 0.77, 0.78, 
    0.82, 0.86, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.85, 0.85, 0.84, 0.84, 
    0.85, 0.87, 0.85, 0.82, 0.82, 0.83, 0.83, 0.85, 0.87, 0.86, 0.87, 0.89, 
    0.89, 0.88, 0.87, 0.87, 0.91, 0.9, 0.87, 0.86, 0.84, 0.82, 0.83, 0.84, 
    0.83, 0.85, 0.86, 0.89, 0.89, 0.88, 0.9, 0.86, 0.82, 0.81, 0.83, 0.85, 
    0.83, 0.87, 0.9, 0.87, 0.88, 0.86, 0.86, 0.84, 0.83, 0.83, 0.82, 0.81, 
    0.78, 0.78, 0.79, 0.81, 0.77, 0.81, 0.79, 0.76, 0.79, 0.8, 0.76, 0.77, 
    0.78, 0.78, 0.78, 0.82, 0.85, 0.82, 0.82, 0.84, 0.73, 0.69, 0.72, 0.79, 
    0.8, 0.8, 0.83, 0.83, 0.83, 0.8, 0.82, 0.84, 0.85, 0.8, 0.79, 0.79, 0.82, 
    0.83, 0.83, 0.83, 0.82, 0.84, 0.81, 0.82, 0.84, 0.84, 0.84, 0.83, 0.83, 
    0.82, 0.84, 0.81, 0.8, 0.8, 0.8, 0.8, 0.79, 0.79, 0.79, 0.79, 0.79, 0.81, 
    0.81, 0.82, 0.8, 0.79, 0.8, 0.81, 0.8, 0.79, 0.8, 0.79, 0.79, 0.8, 0.82, 
    0.82, 0.83, 0.84, 0.87, 0.89, 0.87, 0.84, 0.84, 0.83, 0.84, 0.86, 0.87, 
    0.85, 0.83, 0.82, 0.82, 0.82, 0.81, 0.81, 0.79, 0.8, 0.81, 0.81, 0.82, 
    0.83, 0.82, 0.83, 0.84, 0.85, 0.82, 0.83, 0.85, 0.86, 0.84, 0.89, 0.9, 
    0.86, 0.86, 0.87, 0.86, 0.88, 0.88, 0.88, 0.89, 0.88, 0.88, 0.88, 0.85, 
    0.87, 0.82, 0.89, 0.88, 0.85, 0.84, 0.85, 0.86, 0.86, 0.83, 0.87, 0.87, 
    0.91, 0.84, 0.83, 0.78, 0.78, 0.81, 0.77, 0.73, 0.77, 0.83, 0.75, 0.79, 
    0.89, 0.91, 0.89, 0.84, 0.81, 0.85, 0.88, 0.89, 0.76, 0.89, 0.86, 0.83, 
    0.83, 0.84, 0.88, 0.87, 0.87, 0.89, 0.88, 0.88, 0.88, 0.9, 0.9, 0.89, 
    0.89, 0.89, 0.89, 0.88, 0.87, 0.85, 0.85, 0.85, 0.87, 0.88, 0.89, 0.9, 
    0.9, 0.92, 0.92, 0.93, 0.91, 0.87, 0.84, 0.85, 0.82, 0.86, 0.86, 0.84, 
    0.83, 0.84, 0.84, 0.82, 0.83, 0.82, 0.75, 0.79, 0.75, 0.74, 0.72, 0.79, 
    0.75, 0.73, 0.75, 0.74, 0.72, 0.74, 0.73, 0.74, 0.67, 0.67, 0.7, 0.66, 
    0.66, 0.67, 0.7, 0.68, 0.72, 0.75, 0.7, 0.69, 0.71, 0.68, 0.7, 0.71, 0.7, 
    0.69, 0.7, 0.7, 0.71, 0.76, 0.75, 0.76, 0.74, 0.75, 0.79, 0.79, 0.83, 
    0.82, 0.82, 0.85, 0.85, 0.85, 0.84, 0.84, 0.85, 0.83, 0.85, 0.85, 0.84, 
    0.85, 0.83, 0.81, 0.79, 0.77, 0.75, 0.78, 0.78, 0.79, 0.78, 0.77, 0.79, 
    0.81, 0.8, 0.79, 0.8, 0.78, 0.77, 0.78, 0.79, 0.77, 0.79, 0.78, 0.79, 
    0.79, 0.78, 0.77, 0.76, 0.76, 0.74, 0.73, 0.74, 0.73, 0.72, 0.72, 0.75, 
    0.78, 0.81, 0.83, 0.82, 0.83, 0.8, 0.82, 0.83, 0.81, 0.79, 0.81, 0.83, 
    0.83, 0.83, 0.84, 0.84, 0.85, 0.85, 0.84, 0.84, 0.83, 0.83, 0.87, 0.86, 
    0.89, 0.79, 0.89, 0.87, 0.85, 0.86, 0.85, 0.84, 0.82, 0.83, 0.83, 0.83, 
    0.84, 0.86, 0.89, 0.72, 0.74, 0.76, 0.74, 0.8, 0.8, 0.79, 0.76, 0.74, 
    0.76, 0.73, 0.74, 0.72, 0.72, 0.74, 0.75, 0.78, 0.84, 0.86, 0.84, 0.82, 
    0.83, 0.81, 0.83, 0.78, 0.82, 0.83, 0.82, 0.84, 0.82, 0.83, 0.83, 0.84, 
    0.83, 0.83, 0.83, 0.84, 0.85, 0.86, 0.76, 0.76, 0.81, 0.81, 0.79, 0.82, 
    0.82, 0.84, 0.85, 0.84, 0.87, 0.89, 0.81, 0.77, 0.8, 0.81, 0.69, 0.72, 
    0.77, 0.79, 0.81, 0.85, 0.86, 0.85, 0.86, 0.83, 0.8, 0.85, 0.86, 0.88, 
    0.87, 0.87, 0.86, 0.87, 0.91, 0.88, 0.91, 0.9, 0.89, 0.91, 0.92, 0.91, 
    0.92, 0.92, 0.96, 0.97, 0.96, 0.97, 0.96, 0.94, 0.93, 0.9, 0.91, 0.94, 
    0.94, 0.96, 0.95, 0.95, 0.94, 0.93, 0.91, 0.91, 0.9, 0.9, 0.9, 0.89, 0.9, 
    0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 0.87, 0.87, 0.85, 0.85, 0.83, 0.84, 
    0.82, 0.82, 0.83, 0.82, 0.84, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.84, 
    0.84, 0.84, 0.83, 0.84, 0.84, 0.83, 0.81, 0.82, 0.8, 0.83, 0.83, 0.82, 
    0.81, 0.81, 0.79, 0.78, 0.76, 0.77, 0.82, 0.8, 0.8, 0.79, 0.78, 0.77, 
    0.77, 0.76, 0.75, 0.77, 0.77, 0.77, 0.75, 0.75, 0.74, 0.77, 0.77, 0.76, 
    0.77, 0.77, 0.77, 0.76, 0.76, 0.76, 0.78, 0.76, 0.78, 0.77, 0.78, 0.79, 
    0.8, 0.79, 0.79, 0.78, 0.79, 0.78, 0.78, 0.77, 0.79, 0.77, 0.77, 0.75, 
    0.75, 0.78, 0.77, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.79, 0.79, 0.79, 
    0.78, 0.78, 0.78, 0.76, 0.79, 0.78, 0.77, 0.77, 0.77, 0.77, 0.76, 0.75, 
    0.75, 0.76, 0.75, 0.77, 0.78, 0.78, 0.79, 0.77, 0.77, 0.75, 0.78, 0.77, 
    0.76, 0.72, 0.74, 0.73, 0.75, 0.75, 0.74, 0.76, 0.77, 0.78, 0.76, 0.77, 
    0.77, 0.79, 0.8, 0.8, 0.82, 0.83, 0.81, 0.8, 0.79, 0.77, 0.8, 0.81, 0.79, 
    0.78, 0.79, 0.82, 0.81, 0.78, 0.79, 0.79, 0.8, 0.8, 0.76, 0.77, 0.76, 
    0.76, 0.76, 0.72, 0.77, 0.78, 0.83, 0.84, 0.85, 0.84, 0.84, 0.85, 0.85, 
    0.87, 0.86, 0.86, 0.87, 0.87, 0.86, 0.86, 0.87, 0.87, 0.84, 0.85, 0.84, 
    0.86, 0.86, 0.9, 0.92, 0.92, 0.92, 0.91, 0.87, 0.89, 0.86, 0.82, 0.82, 
    0.78, 0.77, 0.79, 0.79, 0.79, 0.79, 0.78, 0.8, 0.81, 0.83, 0.83, 0.81, 
    0.81, 0.8, 0.82, 0.83, 0.83, 0.83, 0.83, 0.82, 0.82, 0.81, 0.8, 0.78, 
    0.79, 0.78, 0.79, 0.8, 0.81, 0.8, 0.8, 0.79, 0.8, 0.79, 0.76, 0.77, 0.78, 
    0.78, 0.78, 0.78, 0.77, 0.81, 0.82, 0.83, 0.84, 0.85, 0.83, 0.82, 0.81, 
    0.83, 0.83, 0.83, 0.82, 0.81, 0.81, 0.81, 0.81, 0.79, 0.79, 0.77, 0.77, 
    0.77, 0.79, 0.78, 0.79, 0.78, 0.78, 0.78, 0.78, 0.78, 0.77, 0.77, 0.77, 
    0.77, 0.75, 0.75, 0.75, 0.76, 0.77, 0.77, 0.77, 0.78, 0.79, 0.78, 0.79, 
    0.79, 0.78, 0.79, 0.81, 0.8, 0.81, 0.81, 0.79, 0.79, 0.8, 0.79, 0.8, 
    0.79, 0.79, 0.78, 0.78, 0.77, 0.75, 0.75, 0.73, 0.75, 0.75, 0.75, 0.75, 
    0.75, 0.74, 0.75, 0.75, 0.76, 0.77, 0.78, 0.78, 0.77, 0.77, 0.77, 0.74, 
    0.75, 0.76, 0.75, 0.74, 0.74, 0.75, 0.74, 0.74, 0.75, 0.76, 0.76, 0.75, 
    0.74, 0.75, 0.77, 0.76, 0.77, 0.73, 0.77, 0.75, 0.76, 0.77, 0.77, 0.77, 
    0.77, 0.76, 0.78, 0.77, 0.76, 0.77, 0.78, 0.73, 0.75, 0.74, 0.74, 0.75, 
    0.75, 0.77, 0.79, 0.79, 0.77, 0.75, 0.79, 0.79, 0.79, 0.81, 0.79, 0.8, 
    0.8, 0.8, 0.78, 0.78, 0.77, 0.77, 0.78, 0.79, 0.77, 0.75, 0.77, 0.78, 
    0.8, 0.79, 0.79, 0.78, 0.79, 0.81, 0.81, 0.8, 0.81, 0.79, 0.79, 0.78, 
    0.79, 0.8, 0.79, 0.78, 0.79, 0.8, 0.79, 0.79, 0.78, 0.77, 0.78, 0.78, 
    0.78, 0.78, 0.78, 0.78, 0.79, 0.79, 0.78, 0.79, 0.79, 0.79, 0.8, 0.8, 
    0.81, 0.8, 0.78, 0.82, 0.81, 0.81, 0.81, 0.8, 0.81, 0.78, 0.8, 0.81, 
    0.81, 0.81, 0.82, 0.82, 0.84, 0.84, 0.84, 0.85, 0.83, 0.82, 0.8, 0.79, 
    0.83, 0.87, 0.89, 0.86, 0.88, 0.85, 0.84, 0.79, 0.78, 0.71, 0.63, 0.69, 
    0.75, 0.7, 0.75, 0.69, 0.68, 0.7, 0.75, 0.76, 0.8, 0.77, 0.74, 0.8, 0.79, 
    0.79, 0.78, 0.79, 0.79, 0.8, 0.79, 0.79, 0.78, 0.77, 0.77, 0.73, 0.76, 
    0.76, 0.78, 0.78, 0.81, 0.82, 0.83, 0.81, 0.84, 0.85, 0.84, 0.83, 0.84, 
    0.81, 0.78, 0.79, 0.8, 0.8, 0.77, 0.76, 0.69, 0.71, 0.79, 0.78, 0.78, 
    0.79, 0.8, 0.83, 0.77, 0.7, 0.65, 0.61, 0.61, 0.67, 0.69, 0.71, 0.77, 
    0.8, 0.81, 0.78, 0.8, 0.8, 0.8, 0.77, 0.79, 0.79, 0.82, 0.83, 0.84, 0.84, 
    0.85, 0.87, 0.85, 0.86, 0.86, 0.85, 0.84, 0.86, 0.85, 0.86, 0.83, 0.81, 
    0.81, 0.82, 0.83, 0.8, 0.81, 0.78, 0.78, 0.81, 0.84, 0.82, 0.84, 0.84, 
    0.85, 0.85, 0.85, 0.85, 0.86, 0.86, 0.85, 0.86, 0.85, 0.84, 0.84, 0.84, 
    0.84, 0.89, 0.89, 0.86, 0.85, 0.85, 0.86, 0.89, 0.88, 0.88, 0.87, 0.87, 
    0.87, 0.88, 0.87, 0.85, 0.87, 0.87, 0.9, 0.91, 0.91, 0.89, 0.89, 0.91, 
    0.9, 0.89, 0.91, 0.88, 0.9, 0.91, 0.88, 0.87, 0.84, 0.84, 0.84, 0.83, 
    0.87, 0.88, 0.9, 0.86, 0.87, 0.89, 0.87, 0.84, 0.88, 0.86, 0.89, 0.89, 
    0.91, 0.89, 0.89, 0.86, 0.87, 0.85, 0.81, 0.84, 0.84, 0.79, 0.81, 0.76, 
    0.8, 0.82, 0.77, 0.85, 0.82, 0.88, 0.89, 0.86, 0.89, 0.88, 0.88, 0.82, 
    0.84, 0.71, 0.69, 0.68, 0.72, 0.74, 0.77, 0.87, 0.87, 0.76, 0.76, 0.84, 
    0.87, 0.87, 0.88, 0.85, 0.86, 0.87, 0.9, 0.91, 0.84, 0.79, 0.82, 0.86, 
    0.89, 0.91, 0.9, 0.89, 0.87, 0.87, 0.87, 0.88, 0.84, 0.81, 0.86, 0.88, 
    0.87, 0.85, 0.88, 0.92, 0.94, 0.92, 0.92, 0.93, 0.9, 0.88, 0.86, 0.86, 
    0.86, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.83, 0.81, 0.82, 0.82, 
    0.82, 0.88, 0.83, 0.85, 0.88, 0.9, 0.91, 0.9, 0.87, 0.86, 0.85, 0.84, 
    0.83, 0.82, 0.81, 0.8, 0.8, 0.81, 0.79, 0.79, 0.79, 0.78, 0.79, 0.78, 
    0.79, 0.79, 0.79, 0.81, 0.81, 0.8, 0.79, 0.79, 0.79, 0.8, 0.81, 0.81, 
    0.8, 0.79, 0.78, 0.77, 0.79, 0.79, 0.79, 0.81, 0.81, 0.82, 0.82, 0.81, 
    0.81, 0.82, 0.82, 0.83, 0.83, 0.84, 0.83, 0.83, 0.83, 0.82, 0.83, 0.84, 
    0.85, 0.85, 0.84, 0.84, 0.83, 0.82, 0.81, 0.81, 0.8, 0.8, 0.8, 0.8, 0.81, 
    0.81, 0.82, 0.83, 0.84, 0.85, 0.85, 0.86, 0.86, 0.86, 0.85, 0.85, 0.86, 
    0.86, 0.84, 0.84, 0.84, 0.85, 0.81, 0.81, 0.85, 0.85, 0.85, 0.83, 0.83, 
    0.82, 0.8, 0.79, 0.78, 0.77, 0.79, 0.81, 0.82, 0.8, 0.8, 0.78, 0.78, 
    0.78, 0.78, 0.85, 0.78, 0.79, 0.84, 0.84, 0.84, 0.83, 0.84, 0.77, 0.78, 
    0.77, 0.8, 0.81, 0.83, 0.8, 0.81, 0.82, 0.86, 0.86, 0.84, 0.87, 0.87, 
    0.88, 0.89, 0.87, 0.83, 0.79, 0.74, 0.84, 0.86, 0.86, 0.86, 0.86, 0.87, 
    0.89, 0.9, 0.9, 0.9, 0.92, 0.92, 0.92, 0.92, 0.9, 0.9, 0.91, 0.9, 0.9, 
    0.89, 0.86, 0.87, 0.87, 0.85, 0.85, 0.84, 0.82, 0.81, 0.79, 0.8, 0.82, 
    0.75, 0.83, 0.84, 0.83, 0.83, 0.86, 0.86, 0.84, 0.83, 0.83, 0.83, 0.83, 
    0.81, 0.76, 0.73, 0.8, 0.72, 0.81, 0.8, 0.81, 0.82, 0.82, 0.81, 0.8, 0.8, 
    0.78, 0.69, 0.7, 0.76, 0.8, 0.83, 0.86, 0.86, 0.87, 0.78, 0.86, 0.86, 
    0.88, 0.88, 0.89, 0.87, 0.8, 0.81, 0.81, 0.81, 0.8, 0.8, 0.83, 0.82, 
    0.81, 0.82, 0.84, 0.82, 0.83, 0.83, 0.82, 0.82, 0.82, 0.83, 0.83, 0.82, 
    0.82, 0.85, 0.84, 0.85, 0.81, 0.81, 0.8, 0.82, 0.81, 0.83, 0.83, 0.82, 
    0.84, 0.85, 0.84, 0.83, 0.84, 0.83, 0.84, 0.85, 0.85, 0.85, 0.84, 0.83, 
    0.85, 0.85, 0.84, 0.82, 0.82, 0.82, 0.81, 0.82, 0.82, 0.82, 0.82, 0.83, 
    0.84, 0.85, 0.84, 0.85, 0.86, 0.86, 0.86, 0.85, 0.84, 0.83, 0.85, 0.83, 
    0.82, 0.84, 0.83, 0.84, 0.84, 0.83, 0.82, 0.82, 0.82, 0.83, 0.84, 0.84, 
    0.85, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.84, 
    0.81, 0.82, 0.81, 0.81, 0.82, 0.82, 0.79, 0.81, 0.78, 0.79, 0.76, 0.77, 
    0.77, 0.78, 0.79, 0.81, 0.82, 0.84, 0.85, 0.87, 0.88, 0.88, 0.87, 0.88, 
    0.88, 0.81, 0.78, 0.79, 0.79, 0.8, 0.81, 0.79, 0.78, 0.81, 0.81, 0.81, 
    0.82, 0.82, 0.85, 0.84, 0.84, 0.85, 0.82, 0.81, 0.82, 0.82, 0.82, 0.83, 
    0.83, 0.85, 0.85, 0.84, 0.86, 0.85, 0.87, 0.85, 0.85, 0.86, 0.86, 0.88, 
    0.9, 0.89, 0.91, 0.92, 0.93, 0.93, 0.94, 0.93, 0.93, 0.93, 0.88, 0.88, 
    0.87, 0.86, 0.85, 0.84, 0.83, 0.83, 0.83, 0.81, 0.79, 0.8, 0.82, 0.79, 
    0.78, 0.8, 0.8, 0.81, 0.82, 0.82, 0.84, 0.85, 0.83, 0.72, 0.74, 0.81, 
    0.79, 0.82, 0.8, 0.75, 0.66, 0.68, 0.7, 0.68, 0.68, 0.74, 0.78, 0.77, 
    0.8, 0.8, 0.82, 0.82, 0.85, 0.87, 0.86, 0.85, 0.85, 0.85, 0.86, 0.87, 
    0.88, 0.88, 0.87, 0.87, 0.87, 0.87, 0.86, 0.85, 0.85, 0.86, 0.87, 0.87, 
    0.86, 0.87, 0.88, 0.88, 0.85, 0.86, 0.89, 0.91, 0.89, 0.85, 0.84, 0.85, 
    0.83, 0.82, 0.81, 0.81, 0.77, 0.79, 0.78, 0.78, 0.77, 0.77, 0.77, 0.76, 
    0.78, 0.8, 0.79, 0.8, 0.81, 0.82, 0.83, 0.83, 0.83, 0.82, 0.83, 0.84, 
    0.82, 0.82, 0.8, 0.8, 0.72, 0.69, 0.82, 0.83, 0.87, 0.86, 0.87, 0.87, 
    0.88, 0.89, 0.91, 0.93, 0.92, 0.93, 0.94, 0.95, 0.95, 0.93, 0.9, 0.87, 
    0.88, 0.88, 0.87, 0.8, 0.8, 0.79, 0.77, 0.76, 0.75, 0.77, 0.8, 0.81, 
    0.82, 0.81, 0.83, 0.82, 0.81, 0.81, 0.84, 0.84, 0.84, 0.85, 0.85, 0.84, 
    0.84, 0.82, 0.82, 0.84, 0.84, 0.82, 0.79, 0.81, 0.79, 0.76, 0.74, 0.79, 
    0.78, 0.77, 0.81, 0.82, 0.82, 0.76, 0.81, 0.78, 0.81, 0.81, 0.84, 0.84, 
    0.81, 0.82, 0.81, 0.81, 0.77, 0.76, 0.79, 0.82, 0.84, 0.8, 0.83, 0.81, 
    0.84, 0.83, 0.82, 0.83, 0.83, 0.84, 0.85, 0.85, 0.82, 0.82, 0.8, 0.79, 
    0.79, 0.81, 0.81, 0.82, 0.82, 0.82, 0.81, 0.81, 0.82, 0.81, 0.85, 0.84, 
    0.83, 0.83, 0.81, 0.81, 0.81, 0.82, 0.8, 0.82, 0.82, 0.81, 0.79, 0.8, 
    0.78, 0.79, 0.76, 0.77, 0.78, 0.79, 0.77, 0.76, 0.77, 0.78, 0.79, 0.8, 
    0.82, 0.83, 0.83, 0.85, 0.85, 0.84, 0.83, 0.84, 0.85, 0.84, 0.85, 0.85, 
    0.85, 0.85, 0.85, 0.85, 0.83, 0.83, 0.81, 0.8, 0.8, 0.8, 0.79, 0.81, 
    0.82, 0.82, 0.83, 0.84, 0.84, 0.84, 0.85, 0.85, 0.85, 0.85, 0.84, 0.85, 
    0.84, 0.83, 0.83, 0.82, 0.82, 0.82, 0.83, 0.81, 0.81, 0.82, 0.81, 0.81, 
    0.8, 0.81, 0.75, 0.72, 0.76, 0.76, 0.74, 0.74, 0.8, 0.76, 0.79, 0.75, 
    0.78, 0.77, 0.77, 0.75, 0.73, 0.76, 0.79, 0.78, 0.8, 0.79, 0.78, 0.8, 
    0.8, 0.84, 0.84, 0.85, 0.86, 0.85, 0.84, 0.82, 0.82, 0.76, 0.78, 0.73, 
    0.74, 0.78, 0.8, 0.82, 0.79, 0.8, 0.83, 0.84, 0.83, 0.84, 0.84, 0.85, 
    0.84, 0.82, 0.82, 0.82, 0.81, 0.81, 0.81, 0.79, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.8, 0.79, 0.79, 0.78, 0.8, 0.79, 0.81, 0.81, 0.82, 0.83, 0.84, 0.84, 
    0.86, 0.87, 0.89, 0.9, 0.89, 0.88, 0.88, 0.85, 0.84, 0.81, 0.82, 0.8, 
    0.78, 0.79, 0.83, 0.87, 0.87, 0.85, 0.84, 0.86, 0.86, 0.83, 0.8, 0.83, 
    0.83, 0.81, 0.81, 0.81, 0.84, 0.85, 0.86, 0.88, 0.88, 0.89, 0.89, 0.91, 
    0.92, 0.93, 0.93, 0.92, 0.92, 0.91, 0.92, 0.86, 0.87, 0.85, 0.85, 0.86, 
    0.85, 0.83, 0.82, 0.83, 0.8, 0.8, 0.78, 0.83, 0.83, 0.81, 0.82, 0.81, 
    0.81, 0.8, 0.83, 0.8, 0.81, 0.8, 0.81, 0.79, 0.82, 0.82, 0.83, 0.83, 
    0.85, 0.86, 0.87, 0.87, 0.87, 0.87, 0.88, 0.89, 0.89, 0.88, 0.89, 0.85, 
    0.85, 0.83, 0.83, 0.82, 0.81, 0.82, 0.81, 0.82, 0.84, 0.84, 0.84, 0.85, 
    0.87, 0.87, 0.87, 0.87, 0.87, 0.88, 0.87, 0.87, 0.87, 0.85, 0.85, 0.83, 
    0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.84, 0.83, 0.83, 0.84, 0.86, 
    0.86, 0.87, 0.86, 0.86, 0.87, 0.87, 0.87, 0.87, 0.86, 0.86, 0.85, 0.85, 
    0.83, 0.83, 0.81, 0.8, 0.82, 0.82, 0.82, 0.83, 0.84, 0.83, 0.85, 0.85, 
    0.85, 0.86, 0.87, 0.87, 0.87, 0.88, 0.88, 0.89, 0.88, 0.88, 0.85, 0.9, 
    0.89, 0.89, 0.86, 0.86, 0.82, 0.82, 0.83, 0.83, 0.83, 0.83, 0.85, 0.88, 
    0.92, 0.91, 0.92, 0.92, 0.92, 0.91, 0.93, 0.94, 0.94, 0.93, 0.93, 0.92, 
    0.93, 0.93, 0.94, 0.92, 0.89, 0.88, 0.89, 0.88, 0.87, 0.88, 0.88, 0.9, 
    0.92, 0.95, 0.96, 0.97, 0.97, 0.97, 0.94, 0.92, 0.91, 0.91, 0.9, 0.89, 
    0.89, 0.87, 0.88, 0.85, 0.85, 0.86, 0.84, 0.85, 0.85, 0.85, 0.87, 0.87, 
    0.85, 0.85, 0.84, 0.85, 0.85, 0.88, 0.88, 0.88, 0.88, 0.88, 0.87, 0.88, 
    0.87, 0.88, 0.88, 0.88, 0.88, 0.89, 0.89, 0.89, 0.88, 0.89, 0.89, 0.9, 
    0.91, 0.92, 0.81, 0.85, 0.86, 0.86, 0.86, 0.89, 0.81, 0.83, 0.82, 0.84, 
    0.85, 0.85, 0.86, 0.86, 0.87, 0.85, 0.82, 0.82, 0.87, 0.79, 0.83, 0.81, 
    0.8, 0.81, 0.82, 0.83, 0.78, 0.79, 0.85, 0.88, 0.87, 0.86, 0.86, 0.88, 
    0.89, 0.88, 0.86, 0.85, 0.85, 0.85, 0.84, 0.84, 0.84, 0.82, 0.85, 0.83, 
    0.83, 0.81, 0.85, 0.82, 0.82, 0.85, 0.86, 0.87, 0.87, 0.87, 0.86, 0.86, 
    0.83, 0.84, 0.81, 0.81, 0.8, 0.75, 0.72, 0.74, 0.72, 0.78, 0.81, 0.79, 
    0.86, 0.86, 0.88, 0.87, 0.86, 0.88, 0.87, 0.85, 0.82, 0.76, 0.65, 0.74, 
    0.72, 0.7, 0.72, 0.65, 0.64, 0.66, 0.7, 0.74, 0.72, 0.75, 0.76, 0.79, 
    0.8, 0.82, 0.79, 0.78, 0.74, 0.7, 0.73, 0.77, 0.76, 0.75, 0.76, 0.76, 
    0.76, 0.74, 0.79, 0.76, 0.76, 0.78, 0.76, 0.73, 0.78, 0.78, 0.82, 0.87, 
    0.87, 0.83, 0.87, 0.91, 0.93, 0.93, 0.94, 0.95, 0.94, 0.89, 0.9, 0.9, 
    0.87, 0.89, 0.92, 0.93, 0.91, 0.92, 0.9, 0.91, 0.91, 0.9, 0.9, 0.89, 
    0.87, 0.87, 0.87, 0.87, 0.87, 0.86, 0.86, 0.84, 0.84, 0.83, 0.81, 0.78, 
    0.8, 0.75, 0.76, 0.73, 0.73, 0.74, 0.73, 0.72, 0.73, 0.73, 0.69, 0.67, 
    0.65, 0.6, 0.6, 0.61, 0.8, 0.79, 0.6, 0.65, 0.79, 0.79, 0.83, 0.81, 0.87, 
    0.77, 0.73, 0.81, 0.77, 0.75, 0.75, 0.82, 0.82, 0.82, 0.82, 0.82, 0.81, 
    0.82, 0.81, 0.8, 0.83, 0.8, 0.79, 0.77, 0.77, 0.77, 0.76, 0.75, 0.77, 
    0.71, 0.69, 0.68, 0.7, 0.71, 0.69, 0.76, 0.71, 0.76, 0.79, 0.81, 0.82, 
    0.83, 0.84, 0.86, 0.84, 0.87, 0.84, 0.79, 0.8, 0.79, 0.71, 0.82, 0.87, 
    0.87, 0.86, 0.85, 0.81, 0.8, 0.83, 0.85, 0.86, 0.87, 0.9, 0.9, 0.9, 0.9, 
    0.91, 0.91, 0.92, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 0.94, 0.93, 
    0.94, 0.94, 0.93, 0.93, 0.92, 0.93, 0.92, 0.93, 0.94, 0.95, 0.94, 0.95, 
    0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.94, 0.94, 0.92, 0.88, 0.87, 
    0.87, 0.88, 0.87, 0.87, 0.91, 0.91, 0.89, 0.94, 0.95, 0.94, 0.96, 0.96, 
    0.95, 0.94, 0.94, 0.94, 0.95, 0.94, 0.94, 0.93, 0.93, 0.92, 0.91, 0.92, 
    0.9, 0.87, 0.89, 0.87, 0.86, 0.87, 0.87, 0.89, 0.93, 0.94, 0.93, 0.93, 
    0.93, 0.92, 0.88, 0.85, 0.87, 0.89, 0.86, 0.85, 0.82, 0.79, 0.83, 0.82, 
    0.82, 0.82, 0.82, 0.82, 0.79, 0.8, 0.82, 0.84, 0.86, 0.86, 0.87, 0.9, 
    0.92, 0.89, 0.89, 0.88, 0.88, 0.89, 0.89, 0.88, 0.88, 0.89, 0.87, 0.88, 
    0.86, 0.95, 0.95, 0.95, 0.96, 0.96, 0.94, 0.96, 0.96, 0.96, 0.95, 0.95, 
    0.97, 0.98, 0.98, 0.98, 0.97, 0.98, 0.95, 0.96, 0.86, 0.86, 0.85, 0.88, 
    0.86, 0.84, 0.87, 0.87, 0.87, 0.88, 0.88, 0.88, 0.88, 0.87, 0.88, 0.89, 
    0.91, 0.92, 0.93, 0.94, 0.96, 0.96, 0.96, 0.95, 0.95, 0.94, 0.93, 0.93, 
    0.92, 0.92, 0.85, 0.9, 0.91, 0.9, 0.91, 0.89, 0.92, 0.88, 0.9, 0.9, 0.91, 
    0.92, 0.95, 0.95, 0.93, 0.91, 0.93, 0.93, 0.93, 0.91, 0.9, 0.89, 0.88, 
    0.86, 0.84, 0.86, 0.85, 0.83, 0.85, 0.87, 0.87, 0.92, 0.93, 0.93, 0.97, 
    0.98, 0.96, 0.88, 0.86, 0.87, 0.91, 0.93, 0.97, 0.97, 0.96, 0.97, 0.95, 
    0.94, 0.93, 0.91, 0.91, 0.9, 0.9, 0.9, 0.94, 0.9, 0.92, 0.92, 0.94, 0.95, 
    0.95, 0.94, 0.95, 0.93, 0.96, 0.95, 0.95, 0.97, 0.95, 0.92, 0.9, 0.94, 
    0.91, 0.87, 0.89, 0.92, 0.88, 0.88, 0.92, 0.91, 0.9, 0.92, 0.92, 0.92, 
    0.91, 0.9, 0.9, 0.93, 0.93, 0.92, 0.92, 0.93, 0.91, 0.94, 0.94, 0.93, 
    0.95, 0.92, 0.92, 0.94, 0.93, 0.93, 0.92, 0.93, 0.94, 0.92, 0.94, 0.93, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.94, 0.95, 0.96, 0.96, 
    0.94, 0.89, 0.86, 0.84, 0.74, 0.84, 0.84, 0.87, 0.84, 0.85, 0.85, 0.88, 
    0.86, 0.84, 0.84, 0.86, 0.84, 0.91, 0.86, 0.87, 0.84, 0.84, 0.85, 0.81, 
    0.8, 0.84, 0.84, 0.84, 0.87, 0.83, 0.84, 0.83, 0.83, 0.84, 0.85, 0.85, 
    0.84, 0.89, 0.86, 0.87, 0.84, 0.84, 0.84, 0.82, 0.8, 0.78, 0.78, 0.8, 
    0.8, 0.8, 0.79, 0.81, 0.82, 0.84, 0.83, 0.84, 0.87, 0.87, 0.86, 0.85, 
    0.87, 0.87, 0.89, 0.9, 0.89, 0.91, 0.9, 0.91, 0.88, 0.9, 0.86, 0.89, 
    0.87, 0.89, 0.84, 0.87, 0.85, 0.88, 0.88, 0.87, 0.87, 0.92, 0.91, 0.92, 
    0.92, 0.92, 0.91, 0.91, 0.92, 0.93, 0.91, 0.9, 0.9, 0.89, 0.87, 0.88, 
    0.87, 0.91, 0.88, 0.91, 0.91, 0.91, 0.9, 0.92, 0.92, 0.9, 0.91, 0.92, 
    0.93, 0.94, 0.92, 0.93, 0.94, 0.92, 0.91, 0.89, 0.87, 0.86, 0.86, 0.83, 
    0.83, 0.82, 0.77, 0.77, 0.78, 0.78, 0.84, 0.88, 0.94, 0.94, 0.93, 0.93, 
    0.96, 0.97, 0.98, 0.98, 0.98, 0.97, 0.96, 0.95, 0.94, 0.93, 0.91, 0.88, 
    0.9, 0.91, 0.91, 0.87, 0.74, 0.78, 0.83, 0.84, 0.84, 0.82, 0.8, 0.92, 
    0.81, 0.84, 0.89, 0.92, 0.84, 0.85, 0.87, 0.8, 0.85, 0.89, 0.91, 0.85, 
    0.84, 0.85, 0.86, 0.87, 0.86, 0.86, 0.86, 0.88, 0.9, 0.94, 0.91, 0.91, 
    0.92, 0.92, 0.93, 0.92, 0.93, 0.91, 0.89, 0.89, 0.91, 0.91, 0.9, 0.93, 
    0.91, 0.91, 0.9, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.93, 0.93, 0.94, 
    0.94, 0.95, 0.95, 0.96, 0.92, 0.92, 0.92, 0.92, 0.91, 0.86, 0.82, 0.83, 
    0.86, 0.86, 0.89, 0.93, 0.95, 0.94, 0.96, 0.97, 0.96, 0.96, 0.97, 0.98, 
    0.98, 0.97, 0.98, 0.97, 0.97, 0.97, 0.97, 0.93, 0.89, 0.91, 0.92, 0.94, 
    0.93, 0.9, 0.93, 0.85, 0.9, 0.93, 0.92, 0.93, 0.94, 0.95, 0.95, 0.96, 
    0.97, 0.96, 0.97, 0.95, 0.95, 0.93, 0.92, 0.93, 0.93, 0.94, 0.94, 0.91, 
    0.91, 0.87, 0.84, 0.85, 0.83, 0.89, 0.96, 0.95, 0.96, 0.95, 0.95, 0.94, 
    0.95, 0.93, 0.89, 0.85, 0.87, 0.89, 0.89, 0.88, 0.89, 0.88, 0.88, 0.87, 
    0.79, 0.85, 0.84, 0.87, 0.91, 0.89, 0.89, 0.92, 0.94, 0.93, 0.9, 0.88, 
    0.9, 0.87, 0.87, 0.95, 0.95, 0.91, 0.89, 0.89, 0.88, 0.87, 0.88, 0.89, 
    0.91, 0.92, 0.95, 0.97, 0.94, 0.93, 0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 
    0.92, 0.91, 0.91, 0.92, 0.92, 0.91, 0.88, 0.87, 0.85, 0.92, 0.92, 0.96, 
    0.95, 0.96, 0.97, 0.96, 0.94, 0.92, 0.91, 0.94, 0.97, 0.98, 0.97, 0.96, 
    0.95, 0.96, 0.95, 0.95, 0.96, 0.96, 0.94, 0.92, 0.94, 0.91, 0.95, 0.95, 
    0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.95, 0.93, 0.93, 0.91, 0.93, 0.95, 
    0.95, 0.96, 0.91, 0.88, 0.86, 0.9, 0.93, 0.92, 0.93, 0.93, 0.91, 0.92, 
    0.93, 0.94, 0.92, 0.91, 0.91, 0.91, 0.93, 0.96, 0.98, 0.98, 0.98, 0.98, 
    0.96, 0.97, 0.99, 0.96, 0.95, 0.96, 0.96, 0.96, 0.97, 0.96, 0.95, 0.95, 
    0.93, 0.91, 0.92, 0.93, 0.93, 0.94, 0.95, 0.95, 0.94, 0.94, 0.95, 0.96, 
    0.95, 0.96, 0.92, 0.94, 0.95, 0.91, 0.88, 0.9, 0.89, 0.87, 0.83, 0.79, 
    0.82, 0.84, 0.85, 0.88, 0.89, 0.91, 0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 
    0.91, 0.92, 0.9, 0.88, 0.87, 0.93, 0.88, 0.89, 0.89, 0.88, 0.8, 0.83, 
    0.87, 0.84, 0.9, 0.91, 0.91, 0.9, 0.89, 0.75, 0.8, 0.76, 0.73, 0.8, 0.77, 
    0.78, 0.81, 0.8, 0.83, 0.84, 0.88, 0.9, 0.86, 0.81, 0.85, 0.92, 0.89, 
    0.9, 0.91, 0.92, 0.93, 0.95, 0.93, 0.9, 0.96, 0.98, 0.96, 0.93, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 
    0.95, 0.92, 0.97, 0.98, 0.98, 0.97, 0.96, 0.92, 0.91, 0.9, 0.87, 0.89, 
    0.83, 0.8, 0.77, 0.78, 0.87, 0.9, 0.92, 0.91, 0.93, 0.87, 0.89, 0.85, 
    0.77, 0.76, 0.75, 0.88, 0.85, 0.82, 0.79, 0.87, 0.81, 0.78, 0.85, 0.79, 
    0.78, 0.78, 0.85, 0.84, 0.75, 0.79, 0.77, 0.84, 0.89, 0.85, 0.86, 0.87, 
    0.87, 0.86, 0.83, 0.78, 0.75, 0.74, 0.75, 0.78, 0.82, 0.84, 0.85, 0.87, 
    0.89, 0.9, 0.91, 0.96, 0.97, 0.97, 0.94, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.96, 0.95, 0.95, 0.94, 0.96, 
    0.96, 0.95, 0.95, 0.95, 0.97, 0.95, 0.93, 0.91, 0.91, 0.87, 0.83, 0.83, 
    0.88, 0.89, 0.87, 0.88, 0.88, 0.91, 0.93, 0.95, 0.96, 0.97, 0.98, 0.98, 
    0.97, 0.92, 0.92, 0.83, 0.83, 0.79, 0.77, 0.76, 0.76, 0.75, 0.77, 0.74, 
    0.81, 0.81, 0.82, 0.85, 0.85, 0.85, 0.85, 0.82, 0.77, 0.78, 0.76, 0.74, 
    0.78, 0.81, 0.86, 0.85, 0.77, 0.77, 0.78, 0.73, 0.78, 0.79, 0.79, 0.78, 
    0.8, 0.8, 0.85, 0.96, 0.97, 0.96, 0.97, 0.95, 0.94, 0.96, 0.98, 0.99, 
    0.99, 0.93, 0.93, 0.93, 0.94, 0.93, 0.94, 0.95, 0.96, 0.95, 0.93, 0.93, 
    0.94, 0.93, 0.93, 0.94, 0.94, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.98, 0.96, 0.95, 0.93, 0.9, 0.89, 0.85, 0.94, 
    0.82, 0.88, 0.88, 0.89, 0.91, 0.93, 0.95, 0.93, 0.93, 0.93, 0.92, 0.91, 
    0.94, 0.95, 0.98, 0.98, 0.97, 0.95, 0.95, 0.93, 0.88, 0.89, 0.87, 0.89, 
    0.92, 0.94, 0.94, 0.94, 0.94, 0.93, 0.89, 0.89, 0.89, 0.91, 0.91, 0.91, 
    0.88, 0.83, 0.81, 0.79, 0.78, 0.78, 0.69, 0.77, 0.72, 0.67, 0.7, 0.79, 
    0.7, 0.75, 0.68, 0.67, 0.7, 0.76, 0.79, 0.79, 0.82, 0.76, 0.89, 0.93, 
    0.92, 0.88, 0.86, 0.88, 0.92, 0.93, 0.93, 0.81, 0.77, 0.75, 0.84, 0.8, 
    0.8, 0.84, 0.86, 0.82, 0.87, 0.91, 0.96, 0.93, 0.95, 0.98, 0.99, 0.96, 
    0.95, 0.94, 0.97, 0.96, 0.97, 0.99, 0.98, 0.98, 0.98, 0.97, 0.97, 0.98, 
    0.95, 0.86, 0.84, 0.89, 0.92, 0.94, 0.96, 0.98, 0.95, 0.94, 0.97, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.88, 0.88, 0.89, 0.91, 0.95, 
    0.93, 0.93, 0.81, 0.87, 0.86, 0.93, 0.87, 0.88, 0.91, 0.94, 0.92, 0.91, 
    0.89, 0.89, 0.84, 0.88, 0.91, 0.88, 0.89, 0.89, 0.9, 0.92, 0.94, 0.94, 
    0.91, 0.91, 0.9, 0.88, 0.94, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.97, 0.96, 0.97, 
    0.98, 0.96, 0.97, 0.96, 0.97, 0.99, 0.98, 0.97, 0.94, 0.92, 0.93, 0.96, 
    0.97, 0.98, 0.98, 0.97, 0.96, 0.95, 0.95, 0.94, 0.9, 0.92, 0.94, 0.93, 
    0.9, 0.9, 0.9, 0.89, 0.88, 0.88, 0.85, 0.93, 0.9, 0.92, 0.97, 0.98, 0.98, 
    0.98, 0.98, 0.97, 0.98, 0.98, 0.96, 0.94, 0.93, 0.95, 0.97, 0.96, 0.97, 
    0.99, 0.98, 0.91, 0.91, 0.93, 0.93, 0.84, 0.83, 0.84, 0.85, 0.83, 0.8, 
    0.83, 0.83, 0.83, 0.81, 0.83, 0.83, 0.99, 0.84, 0.84, 0.85, 0.89, 0.89, 
    0.88, 0.84, 0.8, 0.8, 0.82, 0.82, 0.82, 0.81, 0.8, 0.8, 0.79, 0.77, 0.87, 
    0.78, 0.81, 0.82, 0.83, 0.82, 0.85, 0.84, 0.81, 0.82, 0.81, 0.85, 0.8, 1, 
    1, 1, 0.72, 0.72, 0.8, 0.83, 0.85, 0.88, 0.88, 0.89, 0.9, 0.88, 0.89, 
    0.84, 0.86, 0.85, 0.93, 0.96, 0.97, 0.95, 0.9, 0.92, 0.94, 0.95, 0.94, 
    0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.96, 0.92, 0.9, 0.87, 0.87, 0.85, 0.82, 0.82, 0.72, 0.84, 0.84, 0.85, 
    0.9, 0.91, 0.9, 0.92, 0.87, 0.87, 0.9, 0.88, 0.95, 0.96, 0.96, 0.97, 
    0.96, 0.97, 0.96, 0.96, 0.88, 0.85, 0.85, 0.86, 0.86, 0.86, 0.87, 0.94, 
    0.94, 0.95, 0.92, 0.94, 0.92, 0.93, 0.93, 0.94, 0.92, 0.96, 0.97, 0.98, 
    0.98, 0.98, 0.98, 0.95, 0.96, 0.96, 0.97, 0.98, 0.97, 0.97, 0.98, 0.96, 
    0.96, 0.97, 0.97, 0.95, 0.97, 0.98, 0.98, 0.98, 0.99, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.94, 0.95, 0.95, 0.93, 0.93, 
    0.93, 0.94, 0.95, 0.95, 0.97, 0.97, 0.97, 0.97, 0.95, 0.93, 0.95, 0.96, 
    0.96, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.97, 0.97, 0.97, 0.96, 0.96, 
    0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 0.96, 
    0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.96, 0.95, 0.86, 0.82, 0.91, 0.89, 0.89, 0.91, 0.89, 0.93, 
    0.92, 0.94, 0.95, 0.9, 0.92, 0.91, 0.92, 0.93, 0.92, 0.9, 0.93, 0.95, 
    0.95, 0.95, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.93, 0.97, 0.98, 0.97, 0.91, 0.9, 
    0.97, 0.94, 0.92, 0.91, 0.92, 0.89, 0.81, 0.83, 0.79, 0.84, 0.78, 0.8, 
    0.82, 0.86, 0.86, 0.89, 0.82, 0.87, 0.83, 0.81, 0.81, 0.85, 0.86, 0.86, 
    0.84, 0.83, 0.87, 0.89, 0.88, 0.93, 0.96, 0.96, 0.95, 0.95, 0.96, 0.95, 
    0.95, 0.95, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    1, 0.99, 0.98, 0.94, 0.95, 0.93, 0.93, 0.93, 0.91, 0.84, 0.82, 0.88, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.95, 0.96, 0.98, 0.98, 0.95, 
    0.95, 0.96, 0.91, 0.92, 0.92, 0.88, 0.92, 0.93, 0.94, 0.91, 0.91, 0.93, 
    0.92, 0.88, 0.89, 0.91, 0.9, 0.9, 0.94, 0.92, 0.95, 0.97, 0.96, 0.98, 
    0.98, 0.99, 0.96, 0.96, 0.93, 0.94, 0.93, 0.94, 0.95, 0.92, 0.91, 0.95, 
    0.94, 0.96, 0.97, 0.97, 0.93, 0.94, 0.94, 0.94, 0.93, 0.92, 0.93, 0.93, 
    0.93, 0.95, 0.97, 0.93, 0.93, 0.94, 0.94, 0.96, 0.93, 0.92, 0.96, 0.96, 
    0.96, 0.96, 0.96, 0.98, 0.98, 0.96, 0.92, 0.97, 0.98, 0.98, 0.97, 0.97, 
    0.98, 0.97, 0.95, 0.91, 0.91, 0.89, 0.9, 0.85, 0.83, 0.85, 0.86, 0.86, 
    0.85, 0.87, 0.92, 0.85, 0.82, 0.91, 0.96, 0.97, 0.98, 0.98, 0.96, 0.98, 
    0.97, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.96, 0.96, 0.96, 0.95, 0.94, 0.96, 
    0.96, 0.95, 0.97, 0.94, 0.94, 0.96, 0.94, 0.96, 0.97, 0.96, 0.97, 0.96, 
    0.97, 0.96, 0.95, 0.96, 0.97, 0.96, 0.96, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.97, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.96, 0.97, 0.98, 0.97, 0.94, 
    0.93, 0.93, 0.93, 0.93, 0.91, 0.9, 0.95, 0.92, 0.91, 0.93, 0.93, 0.95, 
    0.97, 0.97, 0.98, 0.97, 0.95, 0.95, 0.95, 0.93, 0.89, 0.92, 0.9, 0.9, 
    0.9, 0.92, 0.92, 0.91, 0.89, 0.92, 0.93, 0.95, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.96, 0.93, 0.89, 0.86, 0.95, 0.93, 0.96, 0.96, 0.94, 0.92, 0.95, 
    0.93, 0.94, 0.95, 0.97, 0.97, 0.98, 0.97, 0.96, 0.97, 0.97, 0.97, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.97, 0.96, 0.95, 0.93, 0.91, 0.89, 0.91, 0.92, 0.93, 0.93, 
    0.94, 0.97, 0.98, 0.98, 0.97, 0.98, 0.97, 0.94, 0.92, 0.93, 0.91, 0.88, 
    0.9, 0.89, 0.88, 0.88, 0.87, 0.84, 0.87, 0.87, 0.94, 0.96, 0.94, 0.96, 
    0.94, 0.94, 0.93, 0.92, 0.93, 0.93, 0.92, 0.9, 0.91, 0.89, 0.91, 0.91, 
    0.91, 0.91, 0.92, 0.92, 0.93, 0.94, 0.95, 0.95, 0.96, 0.95, 0.97, 0.96, 
    0.96, 0.96, 0.95, 0.96, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.93, 
    0.94, 0.94, 0.93, 0.94, 0.95, 0.95, 0.96, 0.97, 0.97, 0.93, 0.96, 0.96, 
    0.95, 0.96, 0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.98, 0.98, 0.98, 0.96, 
    0.95, 0.92, 0.88, 0.89, 0.89, 0.88, 0.89, 0.87, 0.89, 0.87, 0.89, 0.92, 
    0.91, 0.91, 0.91, 0.93, 0.92, 0.93, 0.95, 0.94, 0.95, 0.95, 0.96, 0.96, 
    0.94, 0.94, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.96, 
    0.96, 0.96, 0.96, 0.96, 0.97, 0.98, 0.97, 0.97, 0.97, 0.98, 1, 0.99, 
    0.98, 0.96, 0.97, 0.97, 0.94, 0.92, 0.92, 0.91, 0.91, 0.93, 0.93, 0.91, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.94, 0.95, 0.94, 0.94, 0.94, 0.9, 0.89, 0.9, 0.93, 0.97, 0.97, 
    0.96, 0.93, 0.89, 0.93, 0.87, 0.81, 0.87, 0.92, 0.94, 0.94, 0.96, 0.95, 
    0.97, 0.97, 0.98, 0.98, 0.97, 0.97, 0.94, 0.93, 0.88, 0.84, 0.87, 0.94, 
    0.94, 0.93, 0.95, 0.94, 0.89, 0.9, 0.91, 0.89, 0.88, 0.89, 0.94, 0.94, 
    0.95, 0.93, 0.94, 0.94, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 
    0.93, 0.93, 0.94, 0.95, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.95, 
    0.97, 0.95, 0.96, 0.93, 0.95, 0.97, 0.97, 0.96, 0.94, 0.94, 0.92, 0.83, 
    0.91, 0.95, 0.97, 0.98, 0.98, 0.99, 0.97, 0.98, 0.95, 0.94, 0.94, 0.93, 
    0.92, 0.92, 0.89, 0.85, 0.81, 0.83, 0.85, 0.85, 0.88, 0.87, 0.83, 0.96, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.95, 0.97, 0.98, 0.98, 0.98, 0.97, 
    0.97, 0.95, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.96, 0.97, 0.98, 0.97, 0.95, 0.92, 0.92, 0.95, 0.97, 0.98, 
    0.98, 0.96, 0.93, 0.96, 0.98, 0.97, 0.98, 0.99, 0.99, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.95, 0.91, 0.93, 0.85, 0.89, 0.91, 
    0.92, 0.94, 0.96, 0.95, 0.97, 0.96, 0.93, 0.94, 0.93, 0.94, 0.95, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.96, 0.96, 
    0.96, 0.96, 0.95, 0.95, 0.94, 0.94, 0.93, 0.94, 0.94, 0.93, 0.91, 0.91, 
    0.91, 0.92, 0.9, 0.89, 0.89, 0.89, 0.9, 0.93, 0.94, 0.92, 0.93, 0.93, 
    0.93, 0.94, 0.95, 0.96, 0.96, 0.95, 0.95, 0.95, 0.94, 0.93, 0.92, 0.92, 
    0.78, 0.87, 0.87, 0.61, 0.72, 0.73, 0.73, 0.72, 0.78, 0.79, 0.77, 0.77, 
    0.77, 0.79, 0.83, 0.85, 0.88, 0.9, 0.89, 0.88, 0.92, 0.9, 0.9, 0.87, 
    0.87, 0.9, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.95, 0.93, 0.93, 
    0.91, 0.91, 0.89, 0.92, 0.94, 0.94, 0.96, 0.98, 0.97, 0.97, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.91, 0.92, 0.91, 0.9, 1, 0.92, 0.91, 0.93, 0.97, 0.88, 0.94, 0.91, 
    0.93, 0.9, 0.9, 0.92, 0.9, 0.9, 0.9, 0.92, 0.94, 0.89, 0.92, 0.89, 0.91, 
    0.91, 0.9, 0.88, 0.89, 0.89, 0.9, 0.91, 0.89, 0.9, 0.9, 0.93, 0.93, 0.91, 
    0.9, 0.91, 0.87, 0.9, 0.93, 0.96, 0.96, 0.95, 0.91, 0.93, 0.9, 0.88, 
    0.85, 0.85, 0.89, 0.87, 0.89, 0.91, 0.92, 0.91, 0.94, 0.9, 0.91, 0.92, 
    0.91, 0.95, 0.97, 0.97, 0.97, 0.97, 0.98, 0.96, 0.96, 0.96, 0.95, 0.96, 
    0.95, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.95, 0.95, 0.96, 0.96, 0.95, 
    0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 
    0.97, 0.98, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.95, 0.96, 0.97, 0.96, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 
    0.91, 0.91, 0.93, 0.95, 0.97, 0.97, 0.94, 0.98, 0.98, 0.98, 0.98, 0.96, 
    0.9, 0.94, 0.93, 0.92, 0.9, 0.91, 0.95, 0.96, 0.94, 0.93, 0.91, 0.9, 0.9, 
    0.86, 0.92, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.97, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.96, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.94, 0.94, 0.97, 0.96, 0.95, 0.96, 0.97, 0.96, 0.95, 0.93, 0.96, 0.94, 
    0.94, 0.94, 0.95, 0.94, 0.95, 0.92, 0.9, 0.9, 0.9, 0.91, 0.94, 0.96, 
    0.97, 0.97, 0.93, 0.95, 0.95, 0.96, 0.96, 0.93, 0.94, 0.94, 0.95, 0.95, 
    0.92, 0.92, 0.94, 0.93, 0.92, 0.94, 0.95, 0.91, 0.95, 0.89, 0.95, 0.96, 
    0.95, 0.96, 0.98, 0.98, 0.98, 0.94, 0.94, 0.84, 0.87, 0.91, 0.91, 0.93, 
    0.96, 0.93, 0.94, 0.97, 0.97, 0.97, 0.96, 0.97, 0.97, 0.95, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.95, 0.96, 0.96, 0.94, 0.95, 0.94, 0.93, 0.95, 0.93, 0.96, 0.95, 0.92, 
    0.92, 0.91, 0.93, 0.94, 0.95, 0.95, 0.93, 0.97, 0.97, 0.91, 0.96, 0.96, 
    0.97, 0.97, 0.96, 0.95, 0.92, 0.94, 0.95, 0.94, 0.95, 0.95, 0.94, 0.91, 
    0.95, 0.92, 0.93, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 0.98, 0.98, 0.99, 
    0.99, 0.98, 0.96, 0.96, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.94, 0.92, 
    0.94, 0.96, 0.96, 0.96, 0.95, 0.93, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.94, 0.94, 0.94, 0.88, 0.87, 0.88, 0.88, 0.9, 0.91, 0.92, 0.93, 
    0.95, 0.96, 0.95, 0.95, 0.94, 0.94, 0.95, 0.94, 0.96, 0.96, 0.96, 0.91, 
    0.86, 0.93, 0.89, 0.8, 0.75, 0.78, 0.73, 0.74, 0.69, 0.72, 0.71, 0.7, 
    0.75, 0.73, 0.77, 0.78, 0.8, 0.8, 0.78, 0.77, 0.74, 0.75, 0.73, 0.74, 
    0.72, 0.74, 0.74, 0.73, 0.71, 0.74, 0.72, 0.71, 0.71, 0.72, 0.71, 0.74, 
    0.74, 0.77, 0.82, 0.8, 0.82, 0.86, 0.84, 0.86, 0.84, 0.81, 0.8, 0.79, 
    0.82, 0.81, 0.81, 0.76, 0.79, 0.79, 0.78, 0.82, 0.84, 0.87, 0.89, 0.84, 
    0.83, 0.86, 0.87, 0.89, 0.86, 0.89, 0.88, 0.89, 0.9, 0.92, 0.93, 0.94, 
    0.95, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.98, 0.97, 0.98, 0.98, 0.97, 0.97, 0.86, 0.85, 0.93, 0.95, 0.9, 
    0.88, 0.86, 0.93, 0.9, 0.92, 0.94, 0.96, 0.94, 0.96, 0.98, 0.98, 0.99, 
    0.98, 0.95, 0.96, 0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.94, 
    0.93, 0.91, 0.9, 0.91, 0.92, 0.86, 0.9, 0.92, 0.81, 0.92, 0.93, 0.91, 
    0.9, 0.85, 0.82, 0.87, 0.91, 0.95, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.97, 0.97, 0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 0.97, 0.94, 0.94, 
    0.94, 0.94, 0.94, 0.91, 0.93, 0.95, 0.98, 0.98, 0.98, 0.93, 0.92, 0.92, 
    0.89, 0.89, 0.95, 0.95, 0.88, 0.86, 0.98, 0.98, 0.94, 0.92, 0.92, 0.92, 
    0.93, 0.95, 0.89, 0.86, 0.79, 0.85, 0.85, 0.86, 0.88, 0.9, 0.89, 0.94, 
    0.94, 0.93, 0.93, 0.94, 0.91, 0.9, 0.93, 0.95, 0.95, 0.97, 0.98, 0.98, 
    0.98, 0.97, 0.97, 0.99, 0.96, 0.95, 0.93, 0.91, 0.88, 0.85, 0.87, 0.89, 
    0.91, 0.89, 0.89, 0.85, 0.82, 0.8, 0.87, 0.9, 0.94, 0.93, 0.87, 0.84, 
    0.85, 0.81, 0.82, 0.81, 0.83, 0.82, 0.83, 0.82, 0.81, 0.8, 0.68, 0.82, 
    0.81, 0.85, 0.85, 0.86, 0.87, 0.88, 0.9, 0.89, 0.86, 0.89, 0.93, 0.87, 
    0.91, 0.91, 0.95, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.94, 
    0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.97, 0.97, 0.94, 0.93, 0.94, 0.92, 0.87, 0.88, 0.82, 0.88, 0.93, 
    0.86, 0.86, 0.84, 0.88, 0.96, 0.98, 0.98, 0.96, 0.99, 0.99, 0.99, 0.97, 
    0.89, 0.92, 0.86, 0.92, 0.91, 0.94, 0.94, 0.95, 0.95, 0.96, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 
    0.97, 0.98, 0.98, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.96, 0.97, 0.96, 0.91, 0.96, 0.96, 0.97, 0.97, 0.98, 0.98, 0.99, 
    0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.9, 0.95, 0.87, 
    0.86, 0.89, 0.91, 0.91, 0.92, 0.88, 0.95, 0.93, 0.91, 0.88, 0.88, 0.87, 
    0.88, 0.9, 0.93, 0.94, 0.95, 0.94, 0.92, 0.92, 0.9, 0.92, 0.92, 0.92, 
    0.97, 0.94, 0.95, 0.93, 0.94, 0.93, 0.93, 0.92, 0.92, 0.93, 0.94, 0.94, 
    0.95, 0.94, 0.93, 0.94, 0.95, 0.96, 0.94, 0.92, 0.94, 0.87, 0.9, 0.87, 
    0.88, 0.8, 0.91, 0.86, 0.79, 0.82, 0.82, 0.82, 0.85, 0.86, 0.86, 0.86, 
    0.85, 0.87, 0.91, 0.94, 0.93, 0.9, 0.92, 0.92, 0.91, 0.92, 0.89, 0.87, 
    0.91, 0.88, 0.89, 0.89, 0.86, 0.87, 0.88, 0.85, 0.84, 0.85, 0.8, 0.77, 
    0.83, 0.81, 0.79, 0.8, 0.77, 0.78, 0.81, 0.72, 0.75, 0.73, 0.74, 0.73, 
    0.75, 0.76, 0.76, 0.75, 0.75, 0.73, 0.71, 0.71, 0.74, 0.75, 0.77, 0.8, 
    0.83, 0.91, 0.94, 0.95, 0.92, 0.88, 0.87, 0.88, 0.9, 0.91, 0.96, 0.98, 
    0.98, 0.99, 0.99, 0.98, 0.92, 0.9, 0.92, 0.96, 0.97, 0.98, 0.97, 0.97, 
    0.97, 0.93, 0.94, 0.95, 0.95, 0.94, 0.93, 0.92, 0.94, 0.94, 0.93, 0.91, 
    0.9, 0.9, 0.88, 0.89, 0.94, 0.96, 0.97, 0.88, 0.92, 0.94, 0.91, 0.96, 
    0.93, 0.95, 0.93, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.97, 0.97, 0.95, 0.94, 0.95, 0.95, 0.96, 0.96, 0.95, 0.94, 0.96, 0.93, 
    0.93, 0.95, 0.97, 0.95, 0.96, 0.97, 0.94, 0.94, 0.97, 0.94, 0.85, 0.93, 
    0.9, 0.93, 0.88, 0.84, 0.85, 0.85, 0.84, 0.86, 0.91, 0.88, 0.89, 0.86, 
    0.84, 0.83, 0.92, 0.93, 0.91, 0.91, 0.94, 0.93, 0.97, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.96, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.94, 0.95, 0.96, 0.96, 0.96, 0.95, 0.92, 0.93, 0.94, 0.95, 
    0.94, 0.92, 0.93, 0.92, 0.9, 0.9, 0.9, 0.9, 0.93, 0.94, 0.95, 0.95, 0.96, 
    0.96, 0.96, 0.95, 0.95, 0.93, 0.94, 0.94, 0.94, 0.92, 0.92, 0.91, 0.93, 
    0.95, 0.94, 0.94, 0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.93, 0.94, 
    0.95, 0.95, 0.95, 0.95, 0.93, 0.93, 0.92, 0.91, 0.93, 0.93, 0.93, 0.91, 
    0.91, 0.92, 0.93, 0.91, 0.9, 0.9, 0.91, 0.92, 0.93, 0.93, 0.92, 0.92, 
    0.93, 0.93, 0.92, 0.9, 0.87, 0.87, 0.85, 0.84, 0.9, 0.89, 0.84, 0.84, 
    0.86, 0.87, 0.88, 0.88, 0.88, 0.83, 0.85, 0.84, 0.84, 0.82, 0.83, 0.82, 
    0.79, 0.76, 0.77, 0.75, 0.7, 0.71, 0.73, 0.76, 0.71, 0.72, 0.73, 0.82, 
    0.81, 0.79, 0.66, 0.75, 0.74, 0.74, 0.74, 0.77, 0.79, 0.82, 0.84, 0.85, 
    0.8, 0.81, 0.79, 0.77, 0.72, 0.75, 0.72, 0.77, 0.78, 0.78, 0.77, 0.77, 
    0.79, 0.8, 0.78, 0.76, 0.74, 0.75, 0.73, 0.73, 0.74, 0.75, 0.77, 0.8, 
    0.79, 0.81, 0.79, 0.81, 0.82, 0.81, 0.82, 0.82, 0.81, 0.81, 0.8, 0.79, 
    0.8, 0.82, 0.83, 0.83, 0.84, 0.83, 0.85, 0.86, 0.88, 0.88, 0.88, 0.88, 
    0.89, 0.89, 0.89, 0.88, 0.88, 0.88, 0.88, 0.89, 0.9, 0.9, 0.9, 0.91, 
    0.89, 0.89, 0.88, 0.9, 0.93, 0.95, 0.93, 0.95, 0.95, 0.95, 0.96, 0.96, 
    0.97, 0.97, 0.97, 0.98, 0.98, 0.99, 0.98, 0.95, 0.94, 0.91, 0.81, 0.88, 
    0.93, 0.9, 0.9, 0.89, 0.86, 0.88, 0.89, 0.86, 0.86, 0.92, 0.95, 0.98, 
    0.98, 0.95, 0.94, 0.94, 0.93, 0.94, 0.86, 0.87, 0.87, 0.85, 0.82, 0.82, 
    0.8, 0.8, 0.83, 0.85, 0.77, 0.78, 0.81, 0.81, 0.81, 0.84, 0.8, 0.85, 
    0.76, 0.77, 0.75, 0.76, 0.72, 0.81, 0.79, 0.79, 0.76, 0.76, 0.8, 0.76, 
    0.78, 0.8, 0.79, 0.79, 0.78, 0.74, 0.71, 0.74, 0.75, 0.73, 0.75, 0.76, 
    0.75, 0.76, 0.73, 0.77, 0.72, 0.75, 0.71, 0.74, 0.72, 0.72, 0.71, 0.71, 
    0.7, 0.72, 0.75, 0.75, 0.75, 0.76, 0.78, 0.78, 0.79, 0.84, 0.84, 0.86, 
    0.88, 0.9, 0.85, 0.76, 0.81, 0.79, 0.8, 0.78, 0.8, 0.79, 0.83, 0.86, 
    0.86, 0.85, 0.85, 0.88, 0.88, 0.89, 0.88, 0.89, 0.86, 0.87, 0.88, 0.86, 
    0.86, 0.86, 0.85, 0.87, 0.88, 0.89, 0.87, 0.89, 0.9, 0.9, 0.89, 0.89, 
    0.9, 0.9, 0.92, 0.92, 0.92, 0.91, 0.91, 0.91, 0.91, 0.91, 0.91, 0.9, 0.9, 
    0.91, 0.91, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 0.92, 
    0.92, 0.91, 0.92, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.94, 0.93, 0.94, 
    0.9, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.9, 
    0.91, 0.91, 0.91, 0.9, 0.89, 0.9, 0.92, 0.91, 0.91, 0.93, 0.94, 0.95, 
    0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.92, 0.91, 0.93, 0.91, 0.92, 0.88, 
    0.83, 0.82, 0.8, 0.87, 0.75, 0.86, 0.88, 0.89, 0.94, 0.97, 0.94, 0.97, 
    0.95, 0.97, 0.97, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.96, 0.96, 
    0.95, 0.96, 0.97, 0.97, 0.96, 0.96, 0.93, 0.92, 0.89, 0.85, 0.88, 0.87, 
    0.87, 0.85, 0.82, 0.83, 0.82, 0.77, 0.78, 0.77, 0.79, 0.82, 0.78, 0.73, 
    0.73, 0.76, 0.74, 0.75, 0.76, 0.77, 0.77, 0.76, 0.76, 0.76, 0.8, 0.81, 
    0.82, 0.81, 0.79, 0.78, 0.82, 0.88, 0.86, 0.88, 0.89, 0.9, 0.91, 0.92, 
    0.91, 0.9, 0.89, 0.89, 0.88, 0.89, 0.89, 0.88, 0.88, 0.87, 0.87, 0.88, 
    0.88, 0.9, 0.89, 0.88, 0.88, 0.89, 0.9, 0.9, 0.9, 0.91, 0.9, 0.9, 0.91, 
    0.91, 0.89, 0.88, 0.89, 0.86, 0.84, 0.84, 0.81, 0.82, 0.81, 0.83, 0.82, 
    0.82, 0.8, 0.83, 0.85, 0.85, 0.86, 0.86, 0.85, 0.86, 0.89, 0.87, 0.93, 
    0.89, 0.89, 0.92, 0.89, 0.87, 0.84, 0.85, 0.84, 0.85, 0.86, 0.87, 0.86, 
    0.85, 0.85, 0.84, 0.82, 0.84, 0.83, 0.82, 0.83, 0.8, 0.83, 0.81, 0.82, 
    0.85, 0.83, 0.8, 0.81, 0.82, 0.83, 0.85, 0.85, 0.85, 0.86, 0.85, 0.86, 
    0.86, 0.86, 0.84, 0.8, 0.77, 0.7, 0.74, 0.75, 0.78, 0.74, 0.78, 0.76, 
    0.76, 0.79, 0.75, 0.8, 0.75, 0.78, 0.76, 0.79, 0.81, 0.79, 0.73, 0.76, 
    0.81, 0.76, 0.74, 0.77, 0.83, 0.83, 0.84, 0.81, 0.77, 0.73, 0.7, 0.72, 
    0.74, 0.78, 0.79, 0.79, 0.82, 0.83, 0.85, 0.86, 0.86, 0.86, 0.84, 0.86, 
    0.85, 0.86, 0.85, 0.82, 0.86, 0.83, 0.85, 0.8, 0.79, 0.77, 0.81, 0.86, 
    0.87, 0.84, 0.78, 0.8, 0.82, 0.81, 0.84, 0.87, 0.86, 0.88, 0.88, 0.83, 
    0.83, 0.79, 0.8, 0.88, 0.89, 0.87, 0.86, 0.88, 0.89, 0.93, 0.91, 0.87, 
    0.86, 0.88, 0.85, 0.81, 0.83, 0.77, 0.79, 0.9, 0.92, 0.9, 0.91, 0.9, 
    0.86, 0.84, 0.82, 0.87, 0.86, 0.86, 0.87, 0.86, 0.84, 0.86, 0.84, 0.82, 
    0.82, 0.82, 0.82, 0.82, 0.83, 0.8, 0.85, 0.84, 0.81, 0.82, 0.84, 0.84, 
    0.85, 0.89, 0.91, 0.91, 0.9, 0.91, 0.91, 0.92, 0.91, 0.91, 0.91, 0.91, 
    0.91, 0.91, 0.91, 0.91, 0.92, 0.92, 0.93, 0.96, 0.98, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.97, 0.98, 0.98, 0.97, 0.93, 0.94, 0.96, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.98, 0.97, 0.98, 0.99, 0.97, 0.97, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.97, 0.96, 0.89, 0.9, 0.94, 0.94, 0.92, 0.92, 0.93, 0.92, 
    0.93, 0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.97, 0.95, 0.92, 0.95, 
    0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.94, 0.92, 0.91, 0.92, 0.95, 0.94, 
    0.97, 0.97, 0.91, 0.92, 0.96, 0.95, 0.93, 0.88, 0.9, 0.93, 0.94, 0.95, 
    0.94, 0.89, 0.85, 0.84, 0.81, 0.85, 0.83, 0.78, 0.75, 0.73, 0.75, 0.79, 
    0.75, 0.76, 0.75, 0.75, 0.74, 0.77, 0.79, 0.81, 0.8, 0.8, 0.8, 0.81, 
    0.81, 0.75, 0.76, 0.74, 0.75, 0.74, 0.77, 0.73, 0.79, 0.75, 0.7, 0.68, 
    0.78, 0.78, 0.8, 0.83, 0.84, 0.85, 0.88, 0.85, 0.87, 0.9, 0.88, 0.86, 
    0.84, 0.86, 0.79, 0.79, 0.79, 0.8, 0.81, 0.76, 0.81, 0.8, 0.83, 0.85, 
    0.81, 0.8, 0.83, 0.81, 0.79, 0.84, 0.85, 0.8, 0.77, 0.75, 0.84, 0.82, 
    0.78, 0.75, 0.72, 0.8, 0.77, 0.76, 0.77, 0.79, 0.79, 0.79, 0.74, 0.77, 
    0.76, 0.78, 0.77, 0.76, 0.75, 0.75, 0.76, 0.77, 0.79, 0.78, 0.78, 0.78, 
    0.77, 0.83, 0.81, 0.83, 0.79, 0.77, 0.81, 0.84, 0.86, 0.84, 0.83, 0.82, 
    0.79, 0.77, 0.67, 0.79, 0.79, 0.8, 0.83, 0.86, 0.78, 0.76, 0.77, 0.8, 
    0.82, 0.83, 0.88, 0.81, 0.79, 0.78, 0.78, 0.8, 0.79, 0.78, 0.75, 0.77, 
    0.77, 0.77, 0.78, 0.77, 0.75, 0.78, 0.76, 0.78, 0.79, 0.78, 0.78, 0.8, 
    0.83, 0.83, 0.82, 0.82, 0.84, 0.83, 0.82, 0.79, 0.79, 0.82, 0.8, 0.79, 
    0.77, 0.73, 0.81, 0.81, 0.81, 0.82, 0.8, 0.78, 0.8, 0.78, 0.79, 0.8, 
    0.81, 0.82, 0.83, 0.83, 0.83, 0.83, 0.83, 0.85, 0.84, 0.8, 0.81, 0.77, 
    0.75, 0.7, 0.71, 0.76, 0.79, 0.78, 0.73, 0.75, 0.82, 0.74, 0.7, 0.71, 
    0.84, 0.76, 0.79, 0.73, 0.74, 0.76, 0.76, 0.79, 0.73, 0.71, 0.75, 0.74, 
    0.81, 0.74, 0.77, 0.72, 0.77, 0.8, 0.7, 0.75, 0.74, 0.74, 0.75, 0.75, 
    0.77, 0.78, 0.74, 0.74, 0.74, 0.76, 0.78, 0.74, 0.74, 0.74, 0.74, 0.77, 
    0.71, 0.74, 0.71, 0.71, 0.71, 0.69, 0.69, 0.72, 0.7, 0.7, 0.73, 0.73, 
    0.74, 0.77, 0.75, 0.77, 0.77, 0.77, 0.76, 0.73, 0.74, 0.75, 0.76, 0.78, 
    0.75, 0.75, 0.77, 0.77, 0.78, 0.81, 0.83, 0.87, 0.88, 0.78, 0.78, 0.82, 
    0.83, 0.87, 0.86, 0.86, 0.77, 0.82, 0.8, 0.83, 0.81, 0.82, 0.89, 0.82, 
    0.8, 0.81, 0.81, 0.81, 0.81, 0.81, 0.79, 0.79, 0.79, 0.78, 0.79, 0.77, 
    0.75, 0.75, 0.78, 0.82, 0.82, 0.81, 0.82, 0.83, 0.83, 0.8, 0.79, 0.81, 
    0.81, 0.81, 0.86, 0.86, 0.88, 0.89, 0.87, 0.84, 0.78, 0.8, 0.78, 0.79, 
    0.79, 0.8, 0.77, 0.77, 0.77, 0.8, 0.81, 0.81, 0.79, 0.78, 0.81, 0.82, 
    0.84, 0.81, 0.83, 0.84, 0.82, 0.77, 0.71, 0.65, 0.73, 0.7, 0.67, 0.73, 
    0.7, 0.72, 0.73, 0.71, 0.68, 0.66, 0.64, 0.64, 0.67, 0.66, 0.76, 0.81, 
    0.79, 0.81, 0.83, 0.83, 0.84, 0.82, 0.83, 0.81, 0.82, 0.81, 0.79, 0.81, 
    0.82, 0.8, 0.81, 0.79, 0.79, 0.8, 0.8, 0.79, 0.79, 0.8, 0.79, 0.84, 0.82, 
    0.84, 0.84, 0.86, 0.87, 0.87, 0.88, 0.88, 0.88, 0.88, 0.89, 0.9, 0.91, 
    0.94, 0.94, 0.94, 0.94, 0.96, 0.97, 0.96, 0.94, 0.91, 0.89, 0.92, 0.89, 
    0.9, 0.88, 0.87, 0.88, 0.89, 0.9, 0.89, 0.91, 0.91, 0.92, 0.93, 0.93, 
    0.93, 0.92, 0.92, 0.91, 0.91, 0.9, 0.9, 0.93, 0.92, 0.92, 0.92, 0.91, 
    0.91, 0.9, 0.89, 0.88, 0.87, 0.88, 0.89, 0.9, 0.89, 0.88, 0.88, 0.9, 
    0.91, 0.9, 0.91, 0.9, 0.9, 0.91, 0.88, 0.88, 0.84, 0.89, 0.86, 0.86, 
    0.87, 0.87, 0.86, 0.87, 0.88, 0.88, 0.88, 0.86, 0.87, 0.87, 0.87, 0.84, 
    0.82, 0.83, 0.82, 0.81, 0.81, 0.82, 0.8, 0.81, 0.8, 0.79, 0.81, 0.81, 
    0.82, 0.83, 0.86, 0.84, 0.86, 0.85, 0.84, 0.84, 0.82, 0.81, 0.83, 0.84, 
    0.83, 0.84, 0.85, 0.85, 0.85, 0.86, 0.87, 0.9, 0.9, 0.89, 0.9, 0.9, 0.88, 
    0.88, 0.88, 0.89, 0.88, 0.87, 0.87, 0.86, 0.87, 0.88, 0.89, 0.88, 0.87, 
    0.87, 0.88, 0.88, 0.88, 0.85, 0.85, 0.85, 0.85, 0.85, 0.84, 0.84, 0.83, 
    0.82, 0.81, 0.77, 0.81, 0.82, 0.85, 0.89, 0.9, 0.87, 0.87, 0.87, 0.78, 
    0.78, 0.75, 0.84, 0.88, 0.86, 0.87, 0.87, 0.87, 0.88, 0.88, 0.87, 0.88, 
    0.88, 0.88, 0.88, 0.9, 0.88, 0.87, 0.87, 0.78, 0.74, 0.78, 0.81, 0.87, 
    0.86, 0.84, 0.83, 0.86, 0.87, 0.87, 0.86, 0.86, 0.85, 0.85, 0.83, 0.82, 
    0.82, 0.82, 0.85, 0.84, 0.84, 0.84, 0.83, 0.84, 0.85, 0.83, 0.83, 0.83, 
    0.85, 0.82, 0.81, 0.81, 0.8, 0.77, 0.83, 0.82, 0.82, 0.85, 0.84, 0.84, 
    0.82, 0.8, 0.8, 0.85, 0.83, 0.85, 0.86, 0.85, 0.86, 0.88, 0.88, 0.87, 
    0.85, 0.84, 0.84, 0.84, 0.84, 0.85, 0.85, 0.85, 0.86, 0.86, 0.84, 0.86, 
    0.87, 0.86, 0.86, 0.88, 0.87, 0.88, 0.87, 0.89, 0.88, 0.88, 0.88, 0.86, 
    0.87, 0.89, 0.89, 0.88, 0.87, 0.84, 0.89, 0.89, 0.9, 0.91, 0.92, 0.92, 
    0.92, 0.9, 0.9, 0.89, 0.86, 0.85, 0.87, 0.89, 0.89, 0.87, 0.88, 0.85, 
    0.83, 0.85, 0.83, 0.84, 0.87, 0.88, 0.86, 0.85, 0.85, 0.89, 0.91, 0.87, 
    0.9, 0.88, 0.88, 0.88, 0.91, 0.89, 0.95, 0.95, 0.87, 0.8, 0.75, 0.82, 
    0.92, 0.89, 0.94, 0.89, 0.87, 0.85, 0.89, 0.91, 0.9, 0.86, 0.85, 0.85, 
    0.85, 0.84, 0.86, 0.86, 0.85, 0.86, 0.85, 0.83, 0.83, 0.82, 0.82, 0.81, 
    0.81, 0.82, 0.84, 0.82, 0.8, 0.8, 0.79, 0.8, 0.8, 0.78, 0.78, 0.77, 0.78, 
    0.79, 0.78, 0.78, 0.8, 0.77, 0.8, 0.81, 0.77, 0.74, 0.72, 0.73, 0.75, 
    0.8, 0.81, 0.82, 0.81, 0.81, 0.82, 0.81, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 
    0.81, 0.79, 0.8, 0.8, 0.79, 0.77, 0.76, 0.79, 0.8, 0.78, 0.8, 0.81, 0.81, 
    0.8, 0.79, 0.8, 0.82, 0.81, 0.8, 0.82, 0.83, 0.86, 0.86, 0.86, 0.86, 
    0.87, 0.88, 0.86, 0.85, 0.89, 0.88, 0.88, 0.9, 0.93, 0.94, 0.93, 0.89, 
    0.9, 0.94, 0.95, 0.94, 0.83, 0.83, 0.83, 0.85, 0.85, 0.87, 0.9, 0.91, 
    0.93, 0.93, 0.94, 0.96, 0.95, 0.95, 0.95, 0.95, 0.93, 0.9, 0.85, 0.86, 
    0.87, 0.89, 0.87, 0.85, 0.83, 0.84, 0.84, 0.89, 0.87, 0.91, 0.88, 0.9, 
    0.92, 0.91, 0.94, 0.91, 0.9, 0.87, 0.84, 0.87, 0.88, 0.86, 0.93, 0.95, 
    0.92, 0.92, 0.93, 0.92, 0.91, 0.91, 0.93, 0.93, 0.93, 0.93, 0.93, 0.93, 
    0.94, 0.96, 0.95, 0.93, 0.92, 0.94, 0.95, 0.94, 0.94, 0.95, 0.95, 0.96, 
    0.96, 0.96, 0.94, 0.93, 0.94, 0.94, 0.96, 0.95, 0.95, 0.94, 0.93, 0.93, 
    0.92, 0.94, 0.95, 0.95, 0.94, 0.94, 0.94, 0.95, 0.94, 0.93, 0.94, 0.94, 
    0.93, 0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 0.96, 0.96, 0.96, 0.96, 0.88, 
    0.93, 0.9, 0.87, 0.9, 0.92, 0.92, 0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 
    0.98, 0.96, 0.96, 0.95, 0.97, 0.97, 0.95, 0.96, 0.97, 0.97, 0.95, 0.95, 
    0.96, 0.95, 0.93, 0.91, 0.94, 0.93, 0.91, 0.91, 0.89, 0.9, 0.91, 0.85, 
    0.89, 0.88, 0.88, 0.88, 0.88, 0.88, 0.87, 0.88, 0.88, 0.89, 0.89, 0.87, 
    0.87, 0.88, 0.87, 0.87, 0.87, 0.88, 0.87, 0.87, 0.88, 0.88, 0.88, 0.88, 
    0.88, 0.88, 0.86, 0.86, 0.85, 0.84, 0.87, 0.89, 0.89, 0.9, 0.88, 0.87, 
    0.87, 0.85, 0.83, 0.84, 0.83, 0.82, 0.83, 0.83, 0.83, 0.84, 0.85, 0.84, 
    0.84, 0.84, 0.84, 0.85, 0.85, 0.85, 0.83, 0.86, 0.84, 0.82, 0.76, 0.7, 
    0.73, 0.81, 0.85, 0.88, 0.87, 0.87, 0.88, 0.85, 0.85, 0.85, 0.87, 0.85, 
    0.84, 0.84, 0.8, 0.82, 0.82, 0.79, 0.78, 0.77, 0.77, 0.76, 0.78, 0.77, 
    0.78, 0.78, 0.77, 0.75, 0.76, 0.78, 0.75, 0.74, 0.77, 0.76, 0.77, 0.78, 
    0.77, 0.75, 0.81, 0.84, 0.85, 0.87, 0.89, 0.9, 0.88, 0.86, 0.86, 0.83, 
    0.87, 0.86, 0.82, 0.8, 0.79, 0.82, 0.8, 0.82, 0.84, 0.86, 0.88, 0.84, 
    0.8, 0.78, 0.78, 0.74, 0.79, 0.79, 0.78, 0.75, 0.57, 0.76, 0.78, 0.85, 
    0.84, 0.83, 0.83, 0.83, 0.82, 0.83, 0.82, 0.82, 0.82, 0.82, 0.81, 0.78, 
    0.79, 0.77, 0.76, 0.76, 0.79, 0.8, 0.78, 0.77, 0.81, 0.83, 0.81, 0.82, 
    0.81, 0.79, 0.79, 0.79, 0.81, 0.82, 0.83, 0.83, 0.82, 0.8, 0.78, 0.77, 
    0.77, 0.77, 0.78, 0.76, 0.77, 0.78, 0.78, 0.77, 0.77, 0.78, 0.79, 0.81, 
    0.81, 0.81, 0.81, 0.81, 0.82, 0.82, 0.82, 0.81, 0.8, 0.78, 0.79, 0.81, 
    0.82, 0.82, 0.81, 0.8, 0.76, 0.74, 0.74, 0.79, 0.82, 0.79, 0.83, 0.87, 
    0.86, 0.88, 0.84, 0.76, 0.66, 0.72, 0.72, 0.76, 0.83, 0.81, 0.8, 0.76, 
    0.76, 0.76, 0.77, 0.79, 0.76, 0.78, 0.77, 0.79, 0.85, 0.81, 0.81, 0.78, 
    0.79, 0.72, 0.65, 0.62, 0.62, 0.72, 0.83, 0.84, 0.83, 0.83, 0.84, 0.84, 
    0.83, 0.83, 0.83, 0.79, 0.83, 0.84, 0.83, 0.81, 0.81, 0.8, 0.83, 0.83, 
    0.83, 0.82, 0.81, 0.81, 0.82, 0.81, 0.8, 0.83, 0.84, 0.85, 0.83, 0.84, 
    0.85, 0.84, 0.83, 0.84, 0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.83, 
    0.83, 0.82, 0.82, 0.81, 0.81, 0.81, 0.81, 0.82, 0.81, 0.81, 0.81, 0.81, 
    0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.81, 0.82, 0.83, 0.83, 0.83, 0.84, 
    0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 0.83, 0.82, 0.83, 0.83, 0.84, 
    0.84, 0.83, 0.84, 0.83, 0.83, 0.84, 0.85, 0.86, 0.85, 0.85, 0.86, 0.85, 
    0.84, 0.83, 0.84, 0.83, 0.86, 0.87, 0.87, 0.87, 0.89, 0.83, 0.81, 0.83, 
    0.81, 0.81, 0.82, 0.81, 0.82, 0.83, 0.82, 0.81, 0.81, 0.82, 0.87, 0.76, 
    0.73, 0.69, 0.75, 0.85, 0.87, 0.89, 0.86, 0.84, 0.84, 0.85, 0.88, 0.9, 
    0.9, 0.88, 0.9, 0.9, 0.9, 0.9, 0.89, 0.91, 0.91, 0.92, 0.91, 0.92, 0.9, 
    0.9, 0.87, 0.9, 0.9, 0.89, 0.87, 0.82, 0.85, 0.82, 0.85, 0.76, 0.71, 
    0.71, 0.7, 0.7, 0.68, 0.73, 0.77, 0.78, 0.79, 0.79, 0.78, 0.8, 0.84, 
    0.84, 0.85, 0.86, 0.87, 0.88, 0.88, 0.88, 0.89, 0.89, 0.86, 0.87, 0.87, 
    0.88, 0.87, 0.89, 0.88, 0.87, 0.88, 0.87, 0.89, 0.89, 0.88, 0.88, 0.88, 
    0.91, 0.95, 0.94, 0.92, 0.92, 0.92, 0.94, 0.94, 0.94, 0.94, 0.94, 0.94, 
    0.95, 0.96, 0.98, 0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.96, 0.96, 0.96, 
    0.96, 0.96, 0.96, 0.96, 0.95, 0.89, 0.89, 0.9, 0.94, 0.94, 0.96, 0.97, 
    0.97, 0.97, 0.96, 0.96, 0.85, 0.81, 0.84, 0.87, 0.88, 0.88, 0.89, 0.93, 
    0.94, 0.95, 0.95, 0.86, 0.79, 0.85, 0.85, 0.88, 0.89, 0.88, 0.87, 0.87, 
    0.92, 0.92, 0.89, 0.88, 0.88, 0.93, 0.91, 0.81, 0.84, 0.83, 0.83, 0.87, 
    0.85, 0.93, 0.96, 0.95, 0.96, 0.98, 0.97, 0.98, 0.98, 0.96, 0.94, 0.93, 
    0.92, 0.91, 0.91, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.91, 0.91, 0.89, 0.88, 
    0.88, 0.85, 0.83, 0.84, 0.84, 0.78, 0.84, 0.79, 0.79, 0.83, 0.83, 0.82, 
    0.82, 0.84, 0.83, 0.83, 0.84, 0.83, 0.84, 0.84, 0.83, 0.85, 0.86, 0.87, 
    0.84, 0.85, 0.84, 0.84, 0.86, 0.86, 0.86, 0.88, 0.89, 0.88, 0.89, 0.87, 
    0.86, 0.85, 0.86, 0.87, 0.87, 0.86, 0.86, 0.88, 0.88, 0.89, 0.91, 0.93, 
    0.96, 0.95, 0.97, 0.96, 0.88, 0.88, 0.88, 0.92, 0.95, 0.94, 0.92, 0.93, 
    0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.91, 0.91, 0.89, 0.9, 0.91, 
    0.9, 0.89, 0.91, 0.91, 0.91, 0.89, 0.88, 0.88, 0.87, 0.87, 0.88, 0.87, 
    0.87, 0.87, 0.87, 0.87, 0.86, 0.87, 0.87, 0.87, 0.87, 0.89, 0.9, 0.91, 
    0.89, 0.88, 0.88, 0.89, 0.86, 0.89, 0.92, 0.92, 0.92, 0.9, 0.94, 0.93, 
    0.93, 0.94, 0.92, 0.9, 0.89, 0.89, 0.89, 0.86, 0.89, 0.92, 0.91, 0.9, 
    0.84, 0.83, 0.91, 0.93, 0.91, 0.92, 0.91, 0.91, 0.89, 0.9, 0.91, 0.92, 
    0.91, 0.9, 0.86, 0.82, 0.83, 0.86, 0.89, 0.87, 0.88, 0.89, 0.9, 0.9, 
    0.91, 0.9, 0.91, 0.9, 0.9, 0.92, 0.92, 0.91, 0.87, 0.88, 0.9, 0.92, 0.92, 
    0.93, 0.91, 0.93, 0.95, 0.96, 0.94, 0.89, 0.83, 0.82, 0.87, 0.91, 0.91, 
    0.89, 0.9, 0.91, 0.91, 0.91, 0.93, 0.94, 0.96, 0.97, 0.98, 0.98, 0.97, 
    0.89, 0.89, 0.95, 0.95, 0.94, 0.91, 0.92, 0.93, 0.94, 0.94, 0.94, 0.92, 
    0.91, 0.91, 0.91, 0.91, 0.98, 0.92, 0.9, 0.89, 0.89, 0.9, 0.89, 0.91, 
    0.89, 0.88, 0.88, 0.9, 0.9, 0.91, 0.88, 0.89, 0.9, 0.93, 0.91, 0.92, 
    0.92, 0.92, 0.93, 0.92, 0.92, 0.88, 0.89, 0.9, 0.9, 0.93, 0.92, 0.93, 
    0.92, 0.92, 0.92, 0.89, 0.89, 0.9, 0.91, 0.89, 0.89, 0.88, 0.89, 0.88, 
    0.86, 0.85, 0.86, 0.9, 0.87, 0.86, 0.85, 0.85, 0.87, 0.86, 0.83, 0.84, 
    0.86, 0.86, 0.83, 0.83, 0.84, 0.83, 0.91, 0.87, 0.89, 0.89, 0.9, 0.87, 
    0.85, 0.82, 0.88, 0.84, 0.74, 0.68, 0.68, 0.65, 0.67, 0.7, 0.64, 0.65, 
    0.66, 0.76, 0.65, 0.66, 0.79, 0.75, 0.79, 0.8, 0.82, 0.83, 0.82, 0.82, 
    0.82, 0.82, 0.83, 0.84, 0.83, 0.83, 0.84, 0.83, 0.84, 0.84, 0.83, 0.83, 
    0.83, 0.83, 0.84, 0.83, 0.83, 0.82, 0.82, 0.82, 0.81, 0.81, 0.81, 0.82, 
    0.83, 0.8, 0.78, 0.8, 0.78, 0.78, 0.79, 0.8, 0.8, 0.79, 0.78, 0.81, 0.85, 
    0.87, 0.85, 0.84, 0.84, 0.86, 0.85, 0.83, 0.82, 0.82, 0.7, 0.73, 0.71, 
    0.65, 0.66, 0.67, 0.65, 0.64, 0.64, 0.68, 0.65, 0.71, 0.74, 0.78, 0.83, 
    0.86, 0.79, 0.76, 0.77, 0.7, 0.71, 0.8, 0.76, 0.7, 0.69, 0.71, 0.77, 
    0.64, 0.65, 0.69, 0.82, 0.81, 0.79, 0.79, 0.74, 0.77, 0.83, 0.85, 0.85, 
    0.84, 0.84, 0.84, 0.83, 0.84, 0.83, 0.84, 0.84, 0.83, 0.83, 0.83, 0.83, 
    0.83, 0.82, 0.82, 0.8, 0.83, 0.82, 0.82, 0.81, 0.81, 0.81, 0.81, 0.81, 
    0.8, 0.8, 0.8, 0.8, 0.81, 0.8, 0.8, 0.78, 0.77, 0.78, 0.78, 0.76, 0.8, 
    0.77, 0.74, 0.74, 0.74, 0.74, 0.75, 0.74, 0.72, 0.74, 0.78, 0.8, 0.82, 
    0.83, 0.84, 0.75, 0.81, 0.73, 0.69, 0.7, 0.7, 0.72, 0.83, 0.86, 0.84, 
    0.84, 0.83, 0.84, 0.83, 0.83, 0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.83, 
    0.83, 0.83, 0.83, 0.83, 0.83, 0.82, 0.8, 0.79, 0.79, 0.77, 0.76, 0.81, 
    0.76, 0.78, 0.84, 0.84, 0.84, 0.85, 0.85, 0.84, 0.84, 0.84, 0.85, 0.84, 
    0.83, 0.82, 0.8, 0.8, 0.76, 0.82, 0.8, 0.78, 0.79, 0.82, 0.83, 0.82, 
    0.82, 0.82, 0.83, 0.86, 0.89, 0.92, 0.91, 0.9, 0.88, 0.89, 0.89, 0.89, 
    0.88, 0.89, 0.91, 0.9, 0.9, 0.87, 0.89, 0.94, 0.94, 0.94, 0.94, 0.93, 
    0.92, 0.92, 0.92, 0.93, 0.95, 0.96, 0.97, 0.96, 0.89, 0.92, 0.93, 0.9, 
    0.93, 0.92, 0.95, 0.96, 0.96, 0.97, 0.98, 0.97, 0.95, 0.92, 0.88, 0.85, 
    0.84, 0.84, 0.83, 0.85, 0.85, 0.82, 0.82, 0.75, 0.64, 0.7, 0.72, 0.76, 
    0.73, 0.76, 0.79, 0.75, 0.76, 0.77, 0.83, 0.84, 0.75, 0.75, 0.74, 0.71, 
    0.69, 0.7, 0.74, 0.73, 0.78, 0.83, 0.83, 0.8, 0.74, 0.77, 0.83, 0.83, 
    0.78, 0.83, 0.81, 0.8, 0.81, 0.82, 0.8, 0.85, 0.82, 0.83, 0.83, 0.85, 
    0.87, 0.9, 0.92, 0.92, 0.91, 0.85, 0.86, 0.91, 0.95, 0.97, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.97, 0.97, 0.97, 0.97, 0.97, 0.96, 0.96, 0.97, 0.96, 
    0.96, 0.96, 0.95, 0.95, 0.94, 0.95, 0.93, 0.95, 0.95, 0.91, 0.91, 0.95, 
    0.96, 0.97, 0.97, 0.97, 0.96, 0.96, 0.95, 0.93, 0.93, 0.93, 0.94, 0.88, 
    0.94, 0.89, 0.86, 0.88, 0.88, 0.85, 0.9, 0.87, 0.91, 0.95, 0.97, 0.97, 
    0.96, 0.93, 0.9, 0.91, 0.9, 0.92, 0.89, 0.93, 0.95, 0.95, 0.93, 0.93, 
    0.94, 0.95, 0.94, 0.95, 0.93, 0.94, 0.94, 0.95, 0.96, 0.95, 0.91, 0.93, 
    0.94, 0.95, 0.97, 0.96, 0.89, 0.88, 0.85, 0.83, 0.84, 0.86, 0.87, 0.89, 
    0.9, 0.91, 0.91, 0.89, 0.9, 0.9, 0.9, 0.86, 0.92, 0.94, 0.95, 0.89, 0.9, 
    0.84, 0.9, 0.84, 0.81, 0.8, 0.82, 0.84, 0.81, 0.81, 0.86, 0.83, 0.84, 
    0.81, 0.71, 0.69, 0.72, 0.75, 0.76, 0.79, 0.87, 0.87, 0.85, 0.84, 0.87, 
    0.87, 0.84, 0.85, 0.84, 0.85, 0.9, 0.9, 0.93, 0.94, 0.83, 0.9, 0.88, 
    0.94, 0.94, 0.95, 0.9, 0.86, 0.84, 0.87, 0.83, 0.87, 0.84, 0.85, 0.83, 
    0.8, 0.81, 0.79, 0.79, 0.83, 0.86, 0.81, 0.76, 0.79, 0.78, 0.79, 0.82, 
    0.83, 0.91, 0.83, 0.87, 0.9, 0.89, 0.89, 0.92, 0.92, 0.88, 0.84, 0.8, 
    0.8, 0.73, 0.79, 0.8, 0.83, 0.86, 0.88, 0.89, 0.93, 0.92, 0.89, 0.87, 
    0.88, 0.88, 0.92, 0.81, 0.89, 0.9, 0.82, 0.83, 0.84, 0.85, 0.87, 0.9, 
    0.88, 0.89, 0.89, 0.93, 0.92, 0.92, 0.92, 0.92, 0.91, 0.92, 0.91, 0.9, 
    0.91, 0.91, 0.88, 0.87, 0.86, 0.85, 0.85, 0.83, 0.84, 0.84, 0.83, 0.83, 
    0.83, 0.84, 0.84, 0.82, 0.79, 0.71, 0.82, 0.84, 0.8, 0.79, 0.78, 0.79, 
    0.78, 0.77, 0.73, 0.7, 0.67, 0.67, 0.64, 0.62, 0.59, 0.6, 0.61, 0.62, 
    0.6, 0.61, 0.73, 0.8, 0.82, 0.82, 0.79, 0.79, 0.81, 0.83, 0.87, 0.88, 
    0.89, 0.89, 0.85, 0.89, 0.89, 0.89, 0.88, 0.88, 0.88, 0.88, 0.86, 0.87, 
    0.87, 0.86, 0.85, 0.84, 0.85, 0.87, 0.82, 0.78, 0.73, 0.65, 0.66, 0.73, 
    0.76, 0.78, 0.76, 0.76, 0.73, 0.73, 0.73, 0.89, 0.77, 0.81, 0.81, 0.81, 
    0.8, 0.82, 0.84, 0.85, 0.85, 0.84, 0.82, 0.8, 0.77, 0.77, 0.76, 0.77, 
    0.74, 0.7, 0.68, 0.66, 0.64, 0.65, 0.64, 0.65, 0.67, 0.72, 0.76, 0.75, 
    0.76, 0.76, 0.74, 0.72, 0.69, 0.68, 0.71, 0.72, 0.7, 0.68, 0.66, 0.67, 
    0.67, 0.73, 0.77, 0.75, 0.75, 0.75, 0.76, 0.77, 0.79, 0.81, 0.85, 0.87, 
    0.87, 0.87, 0.88, 0.88, 0.88, 0.84, 0.81, 0.81, 0.79, 0.76, 0.73, 0.75, 
    0.72, 0.72, 0.73, 0.78, 0.81, 0.84, 0.86, 0.82, 0.8, 0.82, 0.8, 0.71, 
    0.7, 0.74, 0.83, 0.83, 0.83, 0.84, 0.82, 0.84, 0.83, 0.85, 0.84, 0.83, 
    0.83, 0.84, 0.84, 0.82, 0.83, 0.84, 0.83, 0.82, 0.81, 0.83, 0.85, 0.87, 
    0.88, 0.87, 0.87, 0.87, 0.86, 0.86, 0.86, 0.87, 0.86, 0.85, 0.87, 0.84, 
    0.84, 0.84, 0.83, 0.83, 0.83, 0.84, 0.83, 0.84, 0.84, 0.85, 0.86, 0.86, 
    0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.84, 0.83, 0.82, 0.82, 0.84, 0.87, 
    0.86, 0.85, 0.84, 0.83, 0.83, 0.83, 0.84, 0.85, 0.86, 0.87, 0.87, 0.88, 
    0.87, 0.88, 0.88, 0.89, 0.89, 0.9, 0.89, 0.89, 0.87, 0.89, 0.91, 0.91, 
    0.86, 0.81, 0.76, 0.87, 0.89, 0.89, 0.86, 0.93, 0.93, 0.91, 0.9, 0.87, 
    0.86, 0.89, 0.9, 0.9, 0.9, 0.9, 0.91, 0.93, 0.95, 0.94, 0.92, 0.89, 0.87, 
    0.89, 0.88, 0.87, 0.89, 0.86, 0.83, 0.8, 0.75, 0.78, 0.72, 0.7, 0.72, 
    0.72, 0.7, 0.8, 0.72, 0.64, 0.61, 0.61, 0.64, 0.61, 0.63, 0.66, 0.7, 
    0.76, 0.8, 0.83, 0.72, 0.65, 0.62, 0.65, 0.65, 0.56, 0.83, 0.79, 0.81, 
    0.74, 0.66, 0.58, 0.66, 0.68, 0.74, 0.62, 0.7, 0.61, 0.75, 0.72, 0.68, 
    0.6, 0.76, 0.67, 0.77, 0.71, 0.69, 0.72, 0.74, 0.76, 0.76, 0.78, 0.74, 
    0.7, 0.71, 0.72, 0.71, 0.79, 0.73, 0.74, 0.75, 0.72, 0.8, 0.72, 0.79, 
    0.66, 0.73, 0.79, 0.82, 0.82, 0.75, 0.75, 0.76, 0.82, 0.75, 0.8, 0.74, 
    0.75, 0.75, 0.81, 0.78, 0.75, 0.78, 0.77, 0.76, 0.73, 0.71, 0.79, 0.77, 
    0.79, 0.78, 0.76, 0.72, 0.72, 0.73, 0.74, 0.74, 0.75, 0.75, 0.73, 0.78, 
    0.78, 0.74, 0.79, 0.82, 0.76, 0.71, 0.68, 0.72, 0.73, 0.72, 0.75, 0.74, 
    0.77, 0.79, 0.78, 0.77, 0.74, 0.76, 0.74, 0.73, 0.71, 0.72, 0.73, 0.73, 
    0.71, 0.7, 0.71, 0.71, 0.7, 0.72, 0.74, 0.75, 0.75, 0.74, 0.73, 0.73, 
    0.73, 0.73, 0.75, 0.75, 0.76, 0.73, 0.66, 0.71, 0.73, 0.7, 0.75, 0.77, 
    0.8, 0.82, 0.81, 0.81, 0.81, 0.81, 0.78, 0.79, 0.79, 0.8, 0.8, 0.79, 
    0.78, 0.79, 0.77, 0.77, 0.77, 0.77, 0.76, 0.74, 0.75, 0.75, 0.75, 0.75, 
    0.74, 0.74, 0.75, 0.76, 0.76, 0.77, 0.78, 0.78, 0.78, 0.79, 0.77, 0.77, 
    0.78, 0.79, 0.8, 0.81, 0.79, 0.81, 0.81, 0.8, 0.79, 0.79, 0.8, 0.8, 0.79, 
    0.78, 0.79, 0.79, 0.79, 0.78, 0.78, 0.78, 0.78, 0.78, 0.79, 0.79, 0.8, 
    0.81, 0.81, 0.82, 0.82, 0.82, 0.82, 0.82, 0.82, 0.83, 0.83, 0.83, 0.82, 
    0.83, 0.83, 0.83, 0.84, 0.84, 0.83, 0.83, 0.83, 0.83, 0.82, 0.82, 0.83, 
    0.83, 0.83, 0.83, 0.83, 0.83, 0.83, 0.82, 0.82, 0.82, 0.83, 0.82, 0.82, 
    0.82, 0.81, 0.82, 0.83, 0.82, 0.84, 0.84, 0.84, 0.86, 0.87, 0.86, 0.84, 
    0.79, 0.83, 0.82, 0.81, 0.84, 0.83, 0.83, 0.83, 0.76, 0.76, 0.79, 0.82, 
    0.84, 0.83, 0.82, 0.84, 0.82, 0.81, 0.81, 0.82, 0.82, 0.79, 0.79, 0.78, 
    0.8, 0.8, 0.8, 0.77, 0.75, 0.72, 0.7, 0.76, 0.82, 0.79, 0.77, 0.79, 0.78, 
    0.8, 0.82, 0.8, 0.8, 0.81, 0.84, 0.83, 0.83, 0.72, 0.75, 0.78, 0.81, 
    0.79, 0.79, 0.78, 0.77, 0.76, 0.78, 0.73, 0.76, 0.75, 0.73, 0.76, 0.76, 
    0.78, 0.8, 0.78, 0.78, 0.79, 0.83, 0.84, 0.83, 0.84, 0.85, 0.85, 0.84, 
    0.85, 0.86, 0.85, 0.83, 0.84, 0.83, 0.83, 0.82, 0.82, 0.85, 0.83, 0.82, 
    0.81, 0.73, 0.79, 0.74, 0.76, 0.78, 0.77, 0.79, 0.82, 0.8, 0.81, 0.82, 
    0.82, 0.83, 0.81, 0.82, 0.83, 0.82, 0.83, 0.85, 0.86, 0.86, 0.87, 0.87, 
    0.87, 0.87, 0.86, 0.85, 0.86, 0.86, 0.85, 0.87, 0.87, 0.87, 0.89, 0.88, 
    0.9, 0.85, 0.82, 0.88, 0.89, 0.87, 0.87, 0.87, 0.87, 0.86, 0.83, 0.83, 
    0.82, 0.81, 0.86, 0.81, 0.84, 0.83, 0.83, 0.84, 0.85, 0.85, 0.85, 0.84, 
    0.84, 0.85, 0.86, 0.86, 0.86, 0.87, 0.87, 0.87, 0.87, 0.88, 0.89, 0.9, 
    0.86, 0.91, 0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.89, 0.89, 0.88, 0.89, 0.88, 
    0.88, 0.87, 0.85, 0.86, 0.86, 0.85, 0.85, 0.84, 0.82, 0.81, 0.84, 0.83, 
    0.82, 0.83, 0.82, 0.84, 0.83, 0.83, 0.81, 0.82, 0.81, 0.79, 0.79, 0.79, 
    0.79, 0.8, 0.8, 0.8, 0.79, 0.8, 0.8, 0.82, 0.78, 0.79, 0.78, 0.77, 0.76, 
    0.73, 0.75, 0.77, 0.73, 0.71, 0.74, 0.75, 0.76, 0.73, 0.76, 0.76, 0.65, 
    0.76, 0.77, 0.78, 0.8, 0.76, 0.65, 0.74, 0.78, 0.75, 0.73, 0.73, 0.73, 
    0.73, 0.72, 0.72, 0.7, 0.71, 0.71, 0.7, 0.69, 0.7, 0.71, 0.7, 0.71, 0.7, 
    0.72, 0.7, 0.71, 0.72, 0.73, 0.74, 0.74, 0.73, 0.72, 0.73, 0.75, 0.75, 
    0.77, 0.77, 0.76, 0.76, 0.75, 0.75, 0.76, 0.77, 0.77, 0.8, 0.74, 0.78, 
    0.73, 0.71, 0.74, 0.76, 0.79, 0.78, 0.79, 0.79, 0.77, 0.77, 0.77, 0.74, 
    0.73, 0.74, 0.74, 0.77, 0.79, 0.8, 0.8, 0.8, 0.77, 0.77, 0.8, 0.76, 0.79, 
    0.8, 0.78, 0.75, 0.78, 0.79, 0.78, 0.82, 0.83, 0.81, 0.78, 0.76, 0.73, 
    0.73, 0.76, 0.72, 0.73, 0.75, 0.76, 0.76, 0.79, 0.8, 0.78, 0.79, 0.8, 
    0.79, 0.79, 0.78, 0.8, 0.82, 0.83, 0.82, 0.81, 0.8, 0.79, 0.81, 0.8, 
    0.79, 0.79, 0.77, 0.79, 0.8, 0.81, 0.8, 0.81, 0.8, 0.79, 0.8, 0.77, 0.76, 
    0.76, 0.77, 0.78, 0.78, 0.79, 0.78, 0.8, 0.79, 0.79, 0.8, 0.79, 0.78, 
    0.79, 0.8, 0.81, 0.78, 0.8, 0.8, 0.81, 0.82, 0.83, 0.85, 0.86, 0.85, 
    0.82, 0.83, 0.82, 0.78, 0.78, 0.78, 0.76, 0.77, 0.79, 0.8, 0.81, 0.78, 
    0.79, 0.8, 0.81, 0.81, 0.83, 0.84, 0.82, 0.83, 0.8, 0.78, 0.8, 0.78, 
    0.76, 0.75, 0.76, 0.77, 0.79, 0.79, 0.81, 0.82, 0.83, 0.82, 0.82, 0.8, 
    0.81, 0.8, 0.81, 0.81, 0.78, 0.79, 0.81, 0.81, 0.83, 0.83, 0.83, 0.85, 
    0.84, 0.83, 0.83, 0.82, 0.8, 0.82, 0.76, 0.75, 0.76, 0.73, 0.76, 0.71, 
    0.72, 0.74, 0.72, 0.7, 0.69, 0.7, 0.7, 0.72, 0.78, 0.84, 0.85, 0.85, 
    0.86, 0.86, 0.81, 0.74, 0.73, 0.75, 0.79, 0.77, 0.81, 0.78, 0.76, 0.76, 
    0.78, 0.78, 0.78, 0.77, 0.77, 0.79, 0.8, 0.81, 0.79, 0.75, 0.78, 0.83, 
    0.84, 0.85, 0.85, 0.81, 0.8, 0.8, 0.82, 0.86, 0.85, 0.83, 0.8, 0.8, 0.77, 
    0.78, 0.79, 0.78, 0.78, 0.78, 0.79, 0.79, 0.73, 0.75, 0.22, 0.77, 0.78, 
    0.84, 0.81, 0.78, 0.77, 0.79, 0.76, 0.8, 0.73, 0.66, 0.66, 0.64, 0.61, 
    0.58, 0.55, 0.53, 0.58, 0.61, 0.59, 0.65, 0.61, 0.6, 0.65, 0.64, 0.64, 
    0.71, 0.71, 0.71, 0.69, 0.71, 0.71, 0.76, 0.75, 0.75, 0.74, 0.7, 0.67, 
    0.68, 0.75, 0.81, 0.82, 0.78, 0.81, 0.77, 0.76, 0.78, 0.8, 0.83, 0.77, 
    0.79, 0.81, 0.8, 0.74, 0.78, 0.82, 0.8, 0.77, 0.76, 0.74, 0.74, 0.74, 
    0.74, 0.74, 0.74, 0.73, 0.72, 0.72, 0.75, 0.79, 0.8, 0.81, 0.82, 0.85, 
    0.85, 0.83, 0.82, 0.81, 0.8, 0.81, 0.78, 0.79, 0.76, 0.72, 0.74, 0.73, 
    0.72, 0.72, 0.72, 0.72, 0.74, 0.76, 0.77, 0.77, 0.76, 0.78, 0.74, 0.8, 
    0.76, 0.77, 0.78, 0.78, 0.78, 0.77, 0.73, 0.62, 0.67, 0.74, 0.72, 0.72, 
    0.73, 0.68, 0.72, 0.7, 0.69, 0.65, 0.68, 0.71, 0.73, 0.75, 0.84, 0.84, 
    0.86, 0.88, 0.85, 0.83, 0.84, 0.83, 0.82, 0.82, 0.81, 0.8, 0.8, 0.79, 
    0.81, 0.75, 0.75, 0.74, 0.78, 0.81, 0.82, 0.8, 0.83, 0.83, 0.83, 0.83, 
    0.82, 0.81, 0.82, 0.82, 0.84, 0.83, 0.83, 0.82, 0.81, 0.8, 0.79, 0.77, 
    0.77, 0.77, 0.75, 0.75, 0.69, 0.7, 0.74, 0.76, 0.75, 0.72, 0.75, 0.78, 
    0.79, 0.76, 0.71, 0.74, 0.73, 0.79, 0.81, 0.8, 0.78, 0.75, 0.79, 0.78, 
    0.79, 0.78, 0.78, 0.79, 0.79, 0.78, 0.78, 0.79, 0.81, 0.81, 0.82, 0.84, 
    0.84, 0.83, 0.82, 0.83, 0.84, 0.84, 0.85, 0.85, 0.85, 0.85, 0.86, 0.87, 
    0.87, 0.9, 0.88, 0.86, 0.87, 0.81, 0.79, 0.82, 0.83, 0.84, 0.85, 0.84, 
    0.82, 0.81, 0.82, 0.81, 0.82, 0.82, 0.85, 0.87, 0.86, 0.84, 0.83, 0.62, 
    0.64, 0.65, 0.65, 0.66, 0.74, 0.73, 0.74, 0.69, 0.74, 0.82, 0.86, 0.88, 
    0.91, 0.9, 0.9, 0.9, 0.9, 0.9, 0.89, 0.87, 0.81, 0.8, 0.87, 0.9, 0.9, 
    0.89, 0.9, 0.87, 0.83, 0.8, 0.76, 0.77, 0.8, 0.8, 0.83, 0.81, 0.81, 0.82, 
    0.8, 0.83, 0.85, 0.88, 0.87, 0.79, 0.85, 0.82, 0.79, 0.77, 0.74, 0.74, 
    0.71, 0.68, 0.7, 0.75, 0.78, 0.8, 0.81, 0.77, 0.79, 0.74, 0.76, 0.76, 
    0.8, 0.83, 0.85, 0.89, 0.86, 0.88, 0.87, 0.84, 0.85, 0.89, 0.88, 0.87, 
    0.89, 0.89, 0.9, 0.92, 0.91, 0.93, 0.93, 0.93, 0.92, 0.91, 0.92, 0.92, 
    0.93, 0.95, 0.95, 0.93, 0.81, 0.82, 0.8, 0.77, 0.79, 0.73, 0.8, 0.81, 
    0.8, 0.83, 0.82, 0.87, 0.87, 0.87, 0.85, 0.84, 0.84, 0.82, 0.8, 0.8, 
    0.74, 0.76, 0.77, 0.79, 0.78, 0.77, 0.78, 0.77, 0.77, 0.76, 0.75, 0.76, 
    0.74, 0.76, 0.75, 0.74, 0.74, 0.76, 0.79, 0.82, 0.83, 0.75, 0.72, 0.75, 
    0.73, 0.7, 0.74, 0.78, 0.73, 0.67, 0.64, 0.51, 0.54, 0.5, 0.56, 0.7, 
    0.76, 0.76, 0.73, 0.81, 0.81, 0.79, 0.73, 0.66, 0.73, 0.82, 0.83, 0.78, 
    0.75, 0.74, 0.74, 0.76, 0.77, 0.78, 0.78, 0.85, 0.89, 0.88, 0.9, 0.9, 
    0.9, 0.89, 0.89, 0.92, 0.93, 0.92, 0.93, 0.93, 0.92, 0.92, 0.92, 0.94, 
    0.88, 0.86, 0.91, 0.92, 0.93, 0.87, 0.87, 0.89, 0.88, 0.86, 0.85, 0.84, 
    0.84, 0.85, 0.85, 0.86, 0.87, 0.87, 0.85, 0.83, 0.82, 0.82, 0.85, 0.82, 
    0.83, 0.83, 0.83, 0.82, 0.81, 0.79, 0.81, 0.81, 0.85, 0.84, 0.82, 0.82, 
    0.82, 0.82, 0.82, 0.82, 0.83, 0.85, 0.85, 0.88, 0.88, 0.88, 0.86, 0.87, 
    0.88, 0.88, 0.87, 0.86, 0.84, 0.85, 0.85, 0.86, 0.84, 0.84, 0.83, 0.84, 
    0.84, 0.83, 0.82, 0.81, 0.81, 0.84, 0.84, 0.85, 0.85, 0.85, 0.86, 0.84, 
    0.84, 0.87, 0.87, 0.88, 0.87, 0.88, 0.88, 0.87, 0.84, 0.83, 0.81, 0.79, 
    0.79, 0.78, 0.77, 0.78, 0.81, 0.8, 0.8, 0.81, 0.81, 0.79, 0.81, 0.81, 
    0.81, 0.81, 0.79, 0.76, 0.79, 0.82, 0.8, 0.77, 0.81, 0.83, 0.8, 0.77, 
    0.8, 0.81, 0.82, 0.8, 0.8, 0.8, 0.8, 0.8, 0.81, 0.8, 0.79, 0.81, 0.81, 
    0.8, 0.8, 0.79, 0.77, 0.74, 0.74, 0.73, 0.73, 0.67, 0.66, 0.67, 0.69, 
    0.73, 0.77, 0.77, 0.76, 0.81, 0.83, 0.84, 0.83, 0.82, 0.84, 0.85, 0.83, 
    0.8, 0.8, 0.79, 0.76, 0.76, 0.74, 0.73, 0.73, 0.74, 0.72, 0.73, 0.71, 
    0.66, 0.68, 0.7, 0.71, 0.76, 0.75, 0.77, 0.75, 0.76, 0.76, 0.77, 0.76, 
    0.76, 0.73, 0.76, 0.75, 0.75, 0.73, 0.7, 0.73, 0.7, 0.73, 0.69, 0.66, 
    0.67, 0.66, 0.63, 0.63, 0.64, 0.69, 0.71, 0.75, 0.72, 0.79, 0.78, 0.78, 
    0.81, 0.81, 0.81, 0.81, 0.78, 0.74, 0.72, 0.74, 0.74, 0.74, 0.76, 0.73, 
    0.75, 0.77, 0.75, 0.76, 0.76, 0.76, 0.77, 0.79, 0.81, 0.8, 0.82, 0.86, 
    0.84, 0.84, 0.84, 0.83, 0.78, 0.77, 0.75, 0.77, 0.75, 0.75, 0.75, 0.75, 
    0.75, 0.77, 0.79, 0.82, 0.79, 0.77, 0.79, 0.82, 0.82, 0.86, 0.84, 0.84, 
    0.84, 0.82, 0.83, 0.75, 0.75, 0.75, 0.7, 0.73, 0.68, 0.65, 0.68, 0.62, 
    0.62, 0.66, 0.68, 0.71, 0.72, 0.72, 0.78, 0.8, 0.82, 0.83, 0.83, 0.84, 
    0.86, 0.85, 0.84, 0.85, 0.85, 0.85, 0.82, 0.81, 0.79, 0.78, 0.79, 0.79, 
    0.8, 0.8, 0.83, 0.84, 0.86, 0.86, 0.86, 0.86, 0.87, 0.87, 0.86, 0.86, 
    0.88, 0.88, 0.87, 0.87, 0.86, 0.85, 0.84, 0.76, 0.79, 0.8, 0.76, 0.73, 
    0.69, 0.74, 0.81, 0.8, 0.81, 0.78, 0.81, 0.82, 0.87, 0.85, 0.85, 0.87, 
    0.83, 0.85, 0.78, 0.88, 0.89, 0.84, 0.84, 0.83, 0.82, 0.83, 0.84, 0.81, 
    0.8, 0.81, 0.81, 0.81, 0.82, 0.81, 0.82, 0.84, 0.84, 0.85, 0.84, 0.86, 
    0.85, 0.86, 0.86, 0.85, 0.85, 0.86, 0.85, 0.84, 0.84, 0.84, 0.83, 0.82, 
    0.81, 0.81, 0.82, 0.81, 0.82, 0.81, 0.79, 0.8, 0.8, 0.79, 0.75, 0.83, 
    0.83, 0.88, 0.86, 0.88, 0.87, 0.88, 0.88, 0.88, 0.89, 0.89, 0.9, 0.91, 
    0.91, 0.91, 0.91, 0.92, 0.92, 0.93, 0.93, 0.93, 0.92, 0.92, 0.92, 0.92, 
    0.92, 0.93, 0.94, 0.94, 0.93, 0.92, 0.92, 0.9, 0.89, 0.87, 0.84, 0.81, 
    0.82, 0.82, 0.84, 0.9, 0.95, 0.95, 0.94, 0.93, 0.93, 0.94, 0.95, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 
    0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.95, 0.97, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.96, 0.97, 0.97, 0.97, 
    0.97, 0.99, 0.97, 0.98, 0.98, 0.98, 0.99, 0.97, 0.96, 0.95, 0.95, 0.94, 
    0.95, 0.95, 0.96, 0.97, 0.97, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.97, 
    0.96, 0.96, 0.92, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.95, 0.94, 0.93, 0.93, 0.92, 0.93, 0.94, 0.9, 0.95, 0.96, 0.96, 
    0.95, 0.92, 0.91, 0.9, 0.87, 0.83, 0.81, 0.79, 0.84, 0.76, 0.77, 0.71, 
    0.84, 0.83, 0.8, 0.81, 0.86, 0.89, 0.92, 0.92, 0.94, 0.94, 0.96, 0.96, 
    0.97, 0.95, 0.96, 0.94, 0.96, 0.95, 0.95, 0.94, 0.93, 0.95, 0.93, 0.93, 
    0.89, 0.88, 0.89, 0.94, 0.93, 0.92, 0.88, 0.87, 0.89, 0.88, 0.87, 0.81, 
    0.77, 0.82, 0.86, 0.84, 0.89, 0.95, 0.96, 0.96, 0.97, 0.91, 0.92, 0.94, 
    0.95, 0.94, 0.93, 0.93, 0.93, 0.93, 0.92, 0.92, 0.91, 0.92, 0.93, 0.92, 
    0.93, 0.93, 0.92, 0.91, 0.91, 0.91, 0.9, 0.89, 0.89, 0.93, 0.95, 0.94, 
    0.95, 0.94, 0.91, 0.92, 0.91, 0.9, 0.91, 0.91, 0.89, 0.87, 0.86, 0.82, 
    0.79, 0.9, 0.87, 0.84, 0.86, 0.9, 0.88, 0.9, 0.89, 0.89, 0.88, 0.91, 
    0.92, 0.9, 0.91, 0.9, 0.89, 0.89, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 
    0.93, 0.92, 0.9, 0.89, 0.88, 0.91, 0.87, 0.88, 0.89, 0.91, 0.84, 0.87, 
    0.87, 0.88, 0.86, 0.89, 0.89, 0.89, 0.88, 0.85, 0.88, 0.89, 0.9, 0.89, 
    0.89, 0.89, 0.89, 0.89, 0.9, 0.9, 0.91, 0.91, 0.9, 0.9, 0.87, 0.85, 0.84, 
    0.84, 0.81, 0.77, 0.77, 0.78, 0.8, 0.8, 0.78, 0.76, 0.75, 0.74, 0.7, 
    0.69, 0.73, 0.76, 0.79, 0.81, 0.83, 0.87, 0.87, 0.88, 0.89, 0.88, 0.88, 
    0.88, 0.88, 0.87, 0.91, 0.92, 0.93, 0.91, 0.91, 0.91, 0.9, 0.9, 0.88, 
    0.89, 0.89, 0.9, 0.9, 0.85, 0.86, 0.81, 0.82, 0.83, 0.84, 0.84, 0.86, 
    0.85, 0.84, 0.8, 0.79, 0.84, 0.84, 0.83, 0.84, 0.8, 0.82, 0.77, 0.82, 
    0.84, 0.85, 0.9, 0.85, 0.87, 0.85, 0.87, 0.9, 0.91, 0.91, 0.93, 0.93, 
    0.93, 0.92, 0.91, 0.89, 0.91, 0.92, 0.91, 0.91, 0.91, 0.9, 0.9, 0.9, 0.9, 
    0.91, 0.9, 0.92, 0.92, 0.92, 0.93, 0.93, 0.94, 0.94, 0.94, 0.96, 0.96, 
    0.96, 0.97, 0.96, 0.96, 0.9, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.93, 
    0.94, 0.96, 0.96, 0.95, 0.96, 0.95, 0.96, 0.96, 0.95, 0.94, 0.96, 0.97, 
    0.94, 0.95, 0.95, 0.92, 0.91, 0.93, 0.93, 0.91, 0.92, 0.91, 0.92, 0.92, 
    0.94, 0.9, 0.94, 0.94, 0.93, 0.93, 0.95, 0.95, 0.94, 0.94, 0.94, 0.93, 
    0.91, 0.92, 0.92, 0.92, 0.9, 0.91, 0.9, 0.89, 0.88, 0.86, 0.87, 0.84, 
    0.86, 0.82, 0.85, 0.87, 0.87, 0.88, 0.88, 0.88, 0.88, 0.89, 0.88, 0.87, 
    0.88, 0.83, 0.86, 0.84, 0.84, 0.83, 0.83, 0.84, 0.83, 0.75, 0.82, 0.83, 
    0.81, 0.81, 0.8, 0.83, 0.83, 0.8, 0.84, 0.82, 0.85, 0.87, 0.88, 0.86, 
    0.88, 0.83, 0.88, 0.86, 0.87, 0.86, 0.85, 0.86, 0.83, 0.85, 0.88, 0.89, 
    0.87, 0.87, 0.88, 0.88, 0.9, 0.88, 0.91, 0.92, 0.93, 0.94, 0.93, 0.93, 
    0.93, 0.94, 0.9, 0.91, 0.86, 0.84, 0.84, 0.83, 0.79, 0.77, 0.82, 0.83, 
    0.85, 0.85, 0.85, 0.8, 0.85, 0.87, 0.87, 0.88, 0.89, 0.87, 0.86, 0.87, 
    0.82, 0.82, 0.81, 0.76, 0.74, 0.74, 0.75, 0.77, 0.81, 0.88, 0.93, 0.93, 
    0.92, 0.91, 0.93, 0.94, 0.95, 0.97, 0.94, 0.97, 0.97, 0.97, 0.96, 0.95, 
    0.94, 0.93, 0.91, 0.89, 0.94, 0.93, 0.91, 0.9, 0.86, 0.81, 0.78, 0.79, 
    0.81, 0.8, 0.79, 0.79, 0.82, 0.85, 0.85, 0.87, 0.89, 0.89, 0.91, 0.92, 
    0.9, 0.89, 0.88, 0.88, 0.85, 0.88, 0.86, 0.84, 0.82, 0.82, 0.8, 0.78, 
    0.84, 0.82, 0.88, 0.88, 0.86, 0.88, 0.93, 0.9, 0.93, 0.91, 0.93, 0.9, 
    0.9, 0.9, 0.86, 0.86, 0.86, 0.84, 0.87, 0.76, 0.78, 0.75, 0.75, 0.75, 
    0.79, 0.81, 0.82, 0.82, 0.83, 0.85, 0.87, 0.89, 0.91, 0.84, 0.86, 0.79, 
    0.77, 0.8, 0.78, 0.8, 0.81, 0.83, 0.8, 0.81, 0.81, 0.8, 0.81, 0.79, 0.77, 
    0.79, 0.82, 0.83, 0.83, 0.83, 0.85, 0.86, 0.88, 0.85, 0.87, 0.87, 0.86, 
    0.86, 0.86, 0.85, 0.81, 0.82, 0.82, 0.82, 0.8, 0.8, 0.81, 0.79, 0.84, 
    0.84, 0.8, 0.85, 0.85, 0.87, 0.84, 0.87, 0.87, 0.88, 0.86, 0.86, 0.85, 
    0.86, 0.82, 0.79, 0.74, 0.8, 0.78, 0.77, 0.73, 0.76, 0.83, 0.85, 0.84, 
    0.83, 0.86, 0.8, 0.83, 0.84, 0.84, 0.83, 0.82, 0.8, 0.83, 0.8, 0.82, 
    0.83, 0.81, 0.81, 0.8, 0.81, 0.81, 0.81, 0.81, 0.88, 0.87, 0.88, 0.88, 
    0.89, 0.91, 0.92, 0.92, 0.92, 0.92, 0.91, 0.92, 0.92, 0.93, 0.95, 0.92, 
    0.87, 0.89, 0.9, 0.91, 0.9, 0.88, 0.87, 0.89, 0.89, 0.88, 0.88, 0.88, 
    0.89, 0.92, 0.96, 0.97, 0.97, 0.96, 0.95, 0.95, 0.95, 0.94, 0.94, 0.95, 
    0.94, 0.94, 0.96, 0.96, 0.93, 0.93, 0.93, 0.91, 0.91, 0.9, 0.91, 0.92, 
    0.92, 0.91, 0.87, 0.86, 0.88, 0.89, 0.92, 0.94, 0.95, 0.93, 0.93, 0.95, 
    0.96, 0.96, 0.95, 0.95, 0.94, 0.93, 0.87, 0.88, 0.89, 0.89, 0.91, 0.88, 
    0.9, 0.9, 0.91, 0.92, 0.95, 0.94, 0.93, 0.93, 0.91, 0.9, 0.88, 0.87, 
    0.88, 0.84, 0.87, 0.76, 0.8, 0.81, 0.77, 0.76, 0.76, 0.81, 0.82, 0.79, 
    0.78, 0.77, 0.76, 0.84, 0.88, 0.84, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 
    0.85, 0.82, 0.86, 0.85, 0.81, 0.86, 0.87, 0.88, 0.88, 0.86, 0.89, 0.88, 
    0.86, 0.85, 0.89, 0.9, 0.91, 0.93, 0.92, 0.92, 0.93, 0.94, 0.94, 0.95, 
    0.96, 0.95, 0.95, 0.95, 0.95, 0.93, 0.94, 0.94, 0.95, 0.95, 0.95, 0.94, 
    0.92, 0.93, 0.96, 0.93, 0.93, 0.94, 0.94, 0.93, 0.94, 0.93, 0.93, 0.93, 
    0.93, 0.93, 0.91, 0.92, 0.93, 0.94, 0.93, 0.93, 0.92, 0.89, 0.93, 0.92, 
    0.92, 0.92, 0.92, 0.94, 0.95, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 
    0.94, 0.95, 0.94, 0.93, 0.92, 0.91, 0.91, 0.91, 0.9, 0.91, 0.92, 0.92, 
    0.89, 0.89, 0.9, 0.89, 0.85, 0.87, 0.85, 0.86, 0.88, 0.9, 0.92, 0.93, 
    0.94, 0.9, 0.93, 0.82, 0.9, 0.84, 0.89, 0.92, 0.86, 0.84, 0.81, 0.83, 
    0.84, 0.89, 0.85, 0.83, 0.89, 0.87, 0.87, 0.89, 0.85, 0.82, 0.81, 0.76, 
    0.83, 0.82, 0.83, 0.89, 0.82, 0.83, 0.8, 0.8, 0.86, 0.84, 0.8, 0.84, 
    0.83, 0.79, 0.86, 0.87, 0.8, 0.89, 0.81, 0.8, 0.91, 0.82, 0.81, 0.84, 
    0.85, 0.84, 0.86, 0.87, 0.9, 0.92, 0.92, 0.93, 0.92, 0.93, 0.92, 0.91, 
    0.88, 0.89, 0.91, 0.93, 0.92, 0.95, 0.94, 0.95, 0.95, 0.93, 0.87, 0.86, 
    0.81, 0.78, 0.85, 0.82, 0.77, 0.81, 0.86, 0.9, 0.91, 0.94, 0.95, 0.95, 
    0.95, 0.96, 0.96, 0.96, 0.97, 0.97, 0.95, 0.93, 0.91, 0.89, 0.89, 0.95, 
    0.93, 0.91, 0.91, 0.85, 0.83, 0.86, 0.87, 0.83, 0.83, 0.82, 0.86, 0.86, 
    0.87, 0.89, 0.9, 0.91, 0.85, 0.9, 0.89, 0.88, 0.95, 0.97, 0.96, 0.96, 
    0.96, 0.95, 0.95, 0.95, 0.94, 0.92, 0.93, 0.91, 0.91, 0.9, 0.9, 0.95, 
    0.96, 0.96, 0.95, 0.9, 0.91, 0.92, 0.96, 0.97, 0.98, 0.98, 0.98, 0.97, 
    0.96, 0.97, 0.95, 0.94, 0.89, 0.85, 0.8, 0.77, 0.79, 0.74, 0.74, 0.82, 
    0.86, 0.93, 0.81, 0.78, 0.76, 0.74, 0.72, 0.67, 0.69, 0.74, 0.72, 0.75, 
    0.76, 0.81, 0.88, 0.89, 0.84, 0.83, 0.84, 0.87, 0.82, 0.8, 0.83, 0.85, 
    0.86, 0.9, 0.92, 0.94, 0.95, 0.97, 0.97, 0.96, 0.95, 0.94, 0.91, 0.93, 
    0.94, 0.94, 0.9, 0.95, 0.97, 0.97, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 
    0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.98, 0.98, 
    0.98, 0.97, 0.9, 0.95, 0.91, 0.81, 0.82, 0.88, 0.9, 0.88, 0.87, 0.83, 
    0.8, 0.83, 0.91, 0.89, 0.9, 0.86, 0.85, 0.85, 0.85, 0.84, 0.8, 0.8, 0.74, 
    0.75, 0.79, 0.87, 0.89, 0.89, 0.89, 0.87, 0.89, 0.87, 0.85, 0.84, 0.86, 
    0.87, 0.88, 0.89, 0.91, 0.92, 0.93, 0.93, 0.94, 0.93, 0.93, 0.95, 0.94, 
    0.93, 0.94, 0.95, 0.95, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.98, 0.96, 0.93, 0.94, 0.96, 0.96, 0.97, 0.94, 0.95, 
    0.95, 0.94, 0.95, 0.92, 0.89, 0.93, 0.91, 0.91, 0.92, 0.93, 0.93, 0.91, 
    0.95, 0.96, 0.96, 0.95, 0.94, 0.94, 0.94, 0.94, 0.95, 0.95, 0.96, 0.96, 
    0.96, 0.94, 0.91, 0.94, 0.92, 0.9, 0.89, 0.94, 0.91, 0.89, 0.85, 0.89, 
    0.93, 0.92, 0.93, 0.92, 0.93, 0.94, 0.96, 0.97, 0.94, 0.85, 0.92, 0.93, 
    0.93, 0.89, 0.92, 0.95, 0.95, 0.92, 0.96, 0.95, 0.95, 0.91, 0.7, 0.84, 
    0.6, 0.57, 0.84, 0.76, 0.89, 0.84, 0.9, 0.86, 0.9, 0.73, 0.87, 0.83, 
    0.82, 0.93, 0.49, 0.69, 0.84, 0.89, 0.94, 0.93, 0.88, 0.91, 0.92, 0.94, 
    0.95, 0.89, 0.9, 0.9, 0.9, 0.92, 0.91, 0.93, 0.91, 0.93, 0.94, 0.95, 
    0.94, 0.93, 0.93, 0.93, 0.93, 0.93, 0.95, 0.96, 0.96, 0.96, 0.94, 0.97, 
    0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.96, 0.96, 0.98, 0.98, 0.98, 0.98, 
    0.97, 0.94, 0.91, 0.93, 0.95, 0.92, 0.92, 0.96, 0.96, 0.97, 0.97, 0.97, 
    0.98, 0.98, 0.97, 0.97, 0.93, 0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.99, 0.98, 0.96, 0.95, 0.94, 0.91, 0.87, 0.91, 
    0.93, 0.91, 0.87, 0.86, 0.88, 0.89, 0.9, 0.9, 0.92, 0.95, 0.97, 0.94, 
    0.94, 0.96, 0.98, 0.98, 0.97, 0.89, 0.94, 0.93, 0.96, 0.96, 0.98, 0.99, 
    0.99, 0.98, 0.98, 0.97, 0.98, 0.97, 0.96, 0.96, 0.98, 0.96, 0.96, 0.95, 
    0.96, 0.95, 0.96, 0.95, 0.94, 0.97, 0.94, 0.91, 0.94, 0.96, 0.96, 0.97, 
    0.97, 0.96, 0.95, 0.95, 0.94, 0.93, 0.94, 0.94, 0.94, 0.95, 0.96, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.94, 0.91, 0.87, 0.87, 0.88, 0.9, 0.92, 0.94, 0.95, 0.97, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.95, 0.94, 0.95, 0.97, 0.96, 0.96, 0.97, 0.98, 
    0.98, 0.98, 0.9, 0.92, 0.94, 0.91, 0.89, 0.91, 0.9, 0.91, 0.91, 0.88, 
    0.88, 0.89, 0.91, 0.88, 0.84, 0.86, 0.85, 0.87, 0.81, 0.82, 0.79, 0.78, 
    0.88, 0.89, 0.78, 0.84, 0.85, 0.85, 0.82, 0.82, 0.85, 0.72, 0.72, 0.75, 
    0.84, 0.74, 0.8, 0.86, 0.84, 0.89, 0.9, 0.93, 0.87, 0.89, 0.89, 0.88, 
    0.88, 0.9, 0.92, 0.94, 0.96, 0.96, 0.91, 0.94, 0.93, 0.96, 0.96, 0.97, 
    0.98, 0.96, 0.97, 0.98, 0.98, 0.96, 0.98, 0.97, 0.95, 0.94, 0.95, 0.95, 
    0.98, 0.98, 0.98, 0.98, 0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 
    0.99, 0.99, 0.97, 0.97, 0.97, 0.96, 0.94, 0.86, 0.86, 0.88, 0.91, 0.91, 
    0.88, 0.79, 0.8, 0.84, 0.86, 0.92, 0.94, 0.94, 0.94, 0.92, 0.93, 0.93, 
    0.9, 0.88, 0.86, 0.9, 0.91, 0.91, 0.93, 0.95, 0.92, 0.9, 0.89, 0.89, 
    0.92, 0.9, 0.85, 0.86, 0.88, 0.88, 0.91, 0.91, 0.89, 0.88, 0.84, 0.84, 
    0.79, 0.86, 0.83, 0.94, 0.86, 0.86, 0.84, 0.86, 0.85, 0.76, 0.74, 0.74, 
    0.84, 0.83, 0.82, 0.79, 0.81, 0.82, 0.8, 0.73, 0.79, 0.76, 0.8, 0.79, 
    0.79, 0.79, 0.79, 0.8, 0.82, 0.82, 0.87, 0.88, 0.85, 0.84, 0.86, 0.94, 
    0.97, 0.98, 0.98, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.94, 0.89, 
    0.85, 0.86, 0.9, 0.9, 0.85, 0.85, 0.9, 0.9, 0.91, 0.9, 0.85, 0.85, 0.82, 
    0.85, 0.83, 0.82, 0.81, 0.86, 0.87, 0.83, 0.79, 0.79, 0.77, 0.81, 0.85, 
    0.87, 0.88, 0.88, 0.9, 0.91, 0.91, 0.94, 0.94, 0.91, 0.92, 0.89, 0.9, 
    0.9, 0.93, 0.91, 0.9, 0.9, 0.93, 0.97, 0.98, 0.99, 0.98, 0.98, 0.97, 
    0.94, 0.9, 0.87, 0.87, 0.83, 0.8, 0.84, 0.86, 0.89, 0.83, 0.86, 0.85, 
    0.85, 0.86, 0.87, 0.92, 0.96, 0.91, 0.92, 0.92, 0.92, 0.92, 0.91, 0.9, 
    0.96, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.98, 
    0.95, 0.97, 0.98, 0.95, 0.95, 0.93, 0.92, 0.93, 0.92, 0.95, 0.97, 0.98, 
    0.97, 0.92, 0.9, 0.9, 0.88, 0.91, 0.91, 0.85, 0.79, 0.76, 0.82, 0.86, 
    0.88, 0.95, 0.97, 0.98, 0.96, 0.86, 0.88, 0.87, 0.97, 0.98, 0.84, 0.81, 
    0.83, 0.83, 0.78, 0.83, 0.84, 0.88, 0.86, 0.94, 0.96, 0.9, 0.96, 0.94, 
    0.97, 0.92, 0.95, 0.95, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.97, 0.96, 0.88, 0.86, 0.86, 0.86, 0.88, 0.9, 
    0.95, 0.94, 0.96, 0.96, 0.97, 0.96, 0.97, 0.97, 0.96, 0.98, 0.98, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.97, 0.97, 0.97, 0.98, 0.97, 
    0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.94, 0.92, 
    0.93, 0.93, 0.91, 0.93, 0.92, 0.94, 0.94, 0.88, 0.91, 0.9, 0.91, 0.93, 
    0.94, 0.94, 0.93, 0.91, 0.91, 0.95, 0.98, 0.98, 0.99, 0.98, 0.98, 0.97, 
    0.98, 0.96, 0.95, 0.94, 0.86, 0.92, 0.87, 0.91, 0.87, 0.87, 0.85, 0.89, 
    0.89, 0.88, 0.92, 0.9, 0.92, 0.9, 0.91, 0.87, 0.91, 0.91, 0.91, 0.91, 
    0.92, 0.92, 0.93, 0.94, 0.91, 0.95, 0.9, 0.93, 0.88, 0.88, 0.88, 0.82, 
    0.79, 0.88, 0.86, 0.9, 0.91, 0.76, 0.9, 0.89, 0.89, 0.86, 0.87, 0.87, 
    0.86, 0.9, 0.94, 0.96, 0.97, 0.92, 0.95, 0.93, 0.94, 0.95, 0.92, 0.95, 
    0.95, 0.97, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.94, 0.89, 0.85, 0.89, 0.91, 0.83, 0.87, 
    0.81, 0.83, 0.91, 0.92, 0.96, 0.94, 0.97, 0.94, 0.93, 0.92, 0.96, 0.98, 
    0.99, 0.99, 0.98, 0.97, 0.95, 0.97, 0.98, 0.99, 0.98, 0.99, 0.99, 0.99, 
    0.97, 0.99, 0.95, 0.99, 0.91, 0.82, 0.83, 0.87, 0.96, 0.92, 0.9, 0.97, 
    0.97, 0.98, 0.98, 0.98, 0.97, 0.96, 0.91, 0.9, 0.9, 0.91, 0.9, 0.93, 
    0.87, 0.87, 0.87, 0.81, 0.83, 0.87, 0.84, 0.87, 0.86, 0.88, 0.89, 0.89, 
    0.89, 0.87, 0.8, 0.82, 0.89, 0.97, 0.96, 0.95, 0.95, 0.94, 0.85, 0.73, 
    0.81, 0.87, 0.91, 0.93, 0.9, 0.91, 0.89, 0.9, 0.92, 0.95, 0.98, 0.97, 
    0.98, 0.98, 0.94, 0.94, 0.96, 0.97, 0.97, 0.97, 0.87, 0.98, 0.91, 0.93, 
    0.96, 0.95, 0.94, 0.96, 0.96, 0.97, 0.97, 0.95, 0.93, 0.91, 0.93, 0.97, 
    0.95, 0.96, 0.97, 0.98, 0.98, 0.9, 0.84, 0.87, 0.78, 0.88, 0.93, 0.96, 
    0.97, 0.95, 0.93, 0.97, 0.98, 0.99, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.96, 0.94, 
    1, 0.93, 0.92, 0.92, 0.92, 0.95, 0.96, 0.95, 0.95, 0.8, 0.8, 0.92, 0.88, 
    0.89, 0.86, 0.78, 0.82, 0.84, 0.87, 0.83, 0.86, 0.86, 0.87, 0.89, 0.91, 
    0.92, 0.9, 0.93, 0.93, 0.92, 0.95, 0.97, 0.94, 0.91, 0.91, 0.93, 0.94, 
    0.89, 0.83, 0.85, 0.85, 0.9, 0.92, 0.91, 0.92, 0.91, 0.94, 0.95, 0.95, 
    0.95, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.96, 
    0.96, 0.94, 0.96, 0.97, 0.97, 0.96, 0.96, 0.94, 0.95, 0.96, 0.97, 0.93, 
    0.98, 0.98, 0.98, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.95, 0.91, 0.89, 
    0.86, 0.84, 0.84, 0.83, 0.83, 0.81, 0.81, 0.82, 0.82, 0.85, 0.87, 0.89, 
    0.89, 0.91, 0.86, 0.7, 0.71, 0.87, 0.89, 0.91, 0.89, 0.88, 0.88, 0.88, 
    0.88, 0.9, 0.86, 0.9, 0.9, 0.94, 0.93, 0.93, 0.87, 0.87, 0.79, 0.84, 
    0.89, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.95, 0.9, 0.9, 0.88, 0.91, 1, 0.98, 0.98, 0.95, 0.96, 0.97, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 1, 0.99, 0.98, 
    0.95, 0.91, 0.92, 0.89, 0.88, 0.88, 0.9, 0.89, 0.9, 0.92, 0.91, 0.9, 
    0.91, 0.93, 0.94, 0.89, 0.91, 0.95, 0.93, 0.96, 0.97, 0.97, 0.97, 0.97, 
    0.98, 0.98, 0.99, 0.99, 0.93, 0.96, 0.98, 0.99, 0.99, 0.98, 0.97, 0.97, 
    0.95, 0.96, 0.97, 0.98, 0.97, 0.92, 0.93, 0.96, 0.96, 0.94, 0.96, 0.97, 
    0.98, 0.98, 0.98, 0.97, 0.98, 0.98, 0.96, 0.96, 0.97, 0.94, 0.87, 0.83, 
    0.89, 0.93, 0.94, 0.95, 0.95, 0.95, 0.95, 0.97, 0.98, 0.98, 0.97, 0.98, 
    0.99, 0.99, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 
    1, 1, 1, 1, 1, 1, 1, 1, 0.99, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 
    0.99, 1, 1, 0.99, 1, 1, 0.99, 1, 0.99, 1, 1, 1, 0.99, 1, 1, 0.99, 0.99, 
    0.97, 0.96, 0.95, 0.94, 0.93, 0.93, 0.94, 0.95, 0.97, 0.95, 0.91, 0.93, 
    0.92, 0.95, 0.98, 0.87, 0.94, 0.92, 0.92, 0.94, 0.94, 0.95, 0.96, 0.97, 
    0.88, 0.8, 0.82, 0.83, 0.85, 0.83, 0.85, 0.94, 0.91, 0.92, 0.92, 0.97, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.91, 0.94, 0.88, 0.93, 0.95, 0.93, 
    0.95, 0.96, 0.87, 0.94, 0.9, 0.97, 0.98, 0.91, 0.93, 0.92, 0.93, 0.9, 
    0.92, 0.87, 0.85, 0.82, 0.83, 0.9, 0.89, 0.93, 0.93, 0.93, 0.96, 0.95, 
    0.94, 0.95, 0.96, 0.95, 0.95, 0.96, 0.97, 0.97, 0.95, 0.95, 0.95, 0.95, 
    0.92, 0.96, 0.97, 0.96, 0.92, 0.92, 0.93, 0.91, 0.92, 0.95, 0.96, 0.98, 
    0.99, 0.98, 0.9, 0.91, 0.93, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.96, 
    0.97, 0.99, 0.99, 0.98, 0.98, 0.98, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.97, 0.98, 0.94, 0.93, 
    0.94, 0.93, 0.94, 0.94, 0.96, 0.96, 0.94, 0.94, 0.93, 0.93, 0.92, 0.92, 
    0.92, 0.89, 0.82, 0.83, 0.8, 0.81, 0.9, 0.92, 0.97, 0.98, 0.97, 0.96, 
    0.96, 0.97, 0.96, 0.96, 0.97, 0.98, 1, 0.98, 1, 0.98, 0.98, 0.98, 0.98, 
    0.97, 0.96, 0.97, 0.97, 0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.98, 0.96, 
    0.96, 0.95, 0.96, 0.94, 0.97, 0.98, 0.98, 0.98, 0.96, 0.98, 0.98, 0.99, 
    0.99, 0.98, 0.99, 0.98, 0.96, 0.97, 0.98, 0.99, 0.99, 0.98, 0.97, 0.97, 
    0.96, 0.93, 0.92, 0.93, 0.91, 0.94, 0.94, 0.93, 0.97, 0.94, 0.94, 0.97, 
    0.98, 0.98, 0.99, 0.96, 0.97, 0.99, 0.99, 0.96, 0.98, 0.99, 0.99, 0.99, 
    0.96, 0.98, 0.97, 0.98, 0.98, 0.97, 0.96, 0.94, 0.93, 0.97, 0.97, 0.97, 
    0.96, 0.96, 0.95, 0.93, 0.94, 0.94, 0.95, 0.95, 0.97, 0.97, 0.97, 0.92, 
    0.91, 0.9, 0.91, 0.9, 0.88, 0.89, 0.89, 0.89, 0.88, 0.88, 0.86, 0.82, 
    0.82, 0.85, 0.86, 0.88, 0.87, 0.93, 0.86, 0.87, 0.92, 0.93, 0.92, 0.94, 
    0.94, 0.93, 0.93, 0.95, 0.96, 0.97, 0.95, 0.94, 0.97, 0.96, 0.92, 0.93, 
    0.91, 0.93, 0.93, 0.91, 0.93, 0.92, 0.91, 0.89, 0.9, 0.9, 0.89, 0.9, 0.9, 
    0.91, 0.92, 0.94, 0.94, 0.94, 0.94, 0.92, 0.93, 0.92, 0.81, 0.88, 0.89, 
    0.91, 0.89, 0.88, 0.86, 0.83, 0.85, 0.79, 0.76, 0.76, 0.74, 0.82, 0.85, 
    0.87, 0.87, 0.84, 0.77, 0.8, 0.85, 0.89, 0.95, 0.94, 0.96, 0.97, 0.97, 
    0.92, 0.93, 0.96, 0.95, 0.94, 0.94, 0.95, 0.95, 0.97, 0.97, 0.89, 0.85, 
    0.92, 0.93, 0.94, 0.89, 0.92, 0.93, 0.93, 0.93, 0.92, 0.93, 0.93, 0.93, 
    0.94, 0.94, 0.96, 0.96, 0.96, 0.94, 0.94, 0.96, 0.97, 0.97, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.98, 0.96, 0.98, 0.99, 0.98, 0.98, 0.96, 0.97, 1, 
    0.99, 0.98, 0.98, 0.99, 0.99, 0.99, 0.93, 0.89, 0.87, 0.87, 0.83, 0.87, 
    0.92, 0.94, 0.98, 0.98, 0.98, 0.88, 0.86, 0.77, 0.9, 0.9, 0.93, 0.91, 
    0.91, 0.9, 0.91, 0.84, 0.81, 0.81, 0.81, 0.83, 0.81, 0.84, 0.84, 0.89, 
    0.89, 0.86, 0.89, 0.88, 0.86, 0.87, 0.89, 0.88, 0.85, 0.82, 0.83, 0.83, 
    0.84, 0.86, 0.85, 0.85, 0.89, 0.9, 0.93, 0.92, 0.94, 0.94, 0.96, 0.96, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.87, 0.95, 0.97, 0.98, 0.97, 0.96, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 0.99, 0.99, 0.97, 0.97, 
    0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.9, 
    0.95, 0.93, 0.95, 0.97, 0.98, 0.98, 0.97, 0.95, 0.89, 0.87, 0.96, 0.96, 
    0.92, 0.93, 0.91, 0.93, 0.9, 0.89, 0.87, 0.88, 0.88, 0.88, 0.88, 0.9, 
    0.9, 0.9, 0.85, 0.92, 0.86, 0.86, 0.91, 0.93, 0.95, 0.94, 0.94, 0.91, 
    0.94, 0.92, 0.89, 0.87, 0.86, 0.87, 0.88, 0.85, 0.88, 0.9, 0.9, 0.91, 
    0.93, 0.9, 0.94, 0.94, 0.92, 0.93, 0.94, 0.96, 0.97, 0.97, 0.97, 0.96, 
    0.97, 0.98, 0.98, 0.97, 0.97, 0.98, 0.98, 0.99, 0.99, 0.91, 0.9, 0.87, 
    0.89, 0.93, 0.94, 0.91, 0.86, 0.87, 0.91, 0.87, 0.81, 0.94, 0.83, 0.85, 
    0.85, 0.84, 0.84, 0.87, 0.91, 0.94, 0.85, 0.82, 0.79, 0.84, 0.83, 0.85, 
    0.88, 0.88, 0.88, 0.88, 0.83, 0.77, 0.77, 0.82, 0.85, 0.91, 0.94, 0.91, 
    0.92, 0.91, 0.91, 0.89, 0.91, 0.89, 0.87, 0.86, 0.77, 0.89, 0.95, 0.93, 
    0.95, 0.95, 0.96, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.96, 0.86, 0.85, 0.89, 0.88, 0.82, 0.78, 0.85, 0.86, 0.89, 0.96, 0.98, 
    0.97, 0.97, 0.88, 0.85, 0.83, 0.83, 0.84, 0.87, 0.87, 0.89, 0.9, 0.94, 
    0.95, 0.96, 0.94, 0.95, 0.91, 0.91, 0.87, 0.85, 0.87, 0.86, 0.81, 0.87, 
    0.89, 0.87, 0.89, 0.89, 0.83, 0.81, 0.72, 0.79, 0.79, 0.85, 0.77, 0.84, 
    0.92, 0.9, 0.9, 0.87, 0.88, 0.86, 0.87, 0.88, 0.87, 0.93, 0.94, 0.93, 
    0.92, 0.9, 0.91, 0.93, 0.9, 0.91, 0.93, 0.91, 0.93, 0.93, 0.9, 0.89, 
    0.91, 0.83, 0.85, 0.86, 0.81, 0.82, 0.8, 0.78, 0.78, 0.79, 0.79, 0.8, 
    0.84, 0.8, 0.81, 0.85, 0.91, 0.89, 0.87, 0.87, 0.86, 0.86, 0.84, 0.83, 
    0.84, 0.81, 0.82, 0.79, 0.77, 0.77, 0.77, 0.79, 0.76, 0.77, 0.77, 0.93, 
    0.89, 0.9, 0.89, 0.85, 0.82, 0.83, 0.9, 0.87, 0.81, 0.85, 0.82, 0.84, 
    0.82, 0.94, 0.87, 0.85, 0.85, 0.81, 0.92, 0.87, 0.86, 0.82, 0.85, 0.9, 
    0.79, 0.85, 0.82, 0.85, 0.81, 0.82, 0.78, 0.8, 0.81, 0.81, 0.81, 0.84, 
    0.83, 0.86, 0.87, 0.87, 0.87, 0.88, 0.84, 0.86, 0.92, 0.91, 0.95, 0.96, 
    0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.95, 0.96, 0.96, 0.95, 0.95, 0.95, 
    0.94, 0.94, 0.93, 0.91, 0.9, 0.9, 0.92, 0.94, 0.93, 0.87, 0.87, 0.86, 
    0.87, 0.88, 0.86, 0.85, 0.86, 0.87, 0.87, 0.86, 0.87, 0.86, 0.87, 0.87, 
    0.87, 0.84, 0.86, 0.86, 0.85, 0.8, 0.79, 0.8, 0.82, 0.82, 0.81, 0.82, 
    0.83, 0.82, 0.83, 0.83, 0.83, 0.85, 0.83, 0.82, 0.82, 0.82, 0.83, 0.85, 
    0.86, 0.82, 0.81, 0.83, 0.82, 0.79, 0.83, 0.85, 0.83, 0.83, 0.87, 0.84, 
    0.85, 0.84, 0.85, 0.85, 0.86, 0.89, 0.83, 0.86, 0.84, 0.87, 0.83, 0.84, 
    0.84, 0.79, 0.8, 0.8, 0.84, 0.8, 0.81, 0.83, 0.85, 0.87, 0.87, 0.86, 
    0.85, 0.85, 0.83, 0.83, 0.85, 0.81, 0.82, 0.83, 0.77, 0.77, 0.78, 0.76, 
    0.82, 0.82, 0.84, 0.89, 0.89, 0.88, 0.84, 0.86, 0.89, 0.87, 0.91, 0.82, 
    0.78, 0.8, 0.88, 0.91, 0.89, 0.86, 0.87, 0.88, 0.89, 0.86, 0.83, 0.83, 
    0.85, 0.85, 0.86, 0.82, 0.84, 0.79, 0.81, 0.81, 0.79, 0.8, 0.81, 0.86, 
    0.81, 0.79, 0.81, 0.85, 0.85, 0.84, 0.85, 0.85, 0.85, 0.85, 0.87, 0.88, 
    0.88, 0.88, 0.86, 0.83, 0.81, 0.81, 0.82, 0.81, 0.83, 0.84, 0.83, 0.85, 
    0.83, 0.84, 0.82, 0.81, 0.82, 0.87, 0.84, 0.84, 0.86, 0.87, 0.88, 0.88, 
    0.88, 0.88, 0.89, 0.91, 0.91, 0.92, 0.92, 0.91, 0.92, 0.92, 0.91, 0.92, 
    0.92, 0.93, 0.92, 0.93, 0.93, 0.94, 0.94, 0.97, 0.98, 0.99, 0.99, 0.96, 
    0.98, 0.97, 0.96, 0.98, 0.97, 0.96, 0.94, 0.95, 0.96, 0.93, 0.94, 0.96, 
    0.96, 0.98, 0.98, 0.98, 0.99, 0.95, 0.94, 0.97, 0.98, 0.97, 0.96, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.96, 0.95, 
    0.95, 0.9, 0.93, 0.98, 0.99, 0.99, 0.97, 0.96, 0.95, 0.91, 0.9, 0.9, 
    0.91, 0.9, 0.87, 0.87, 0.93, 0.89, 0.87, 0.86, 0.92, 0.89, 0.85, 0.86, 
    0.87, 0.87, 0.84, 0.83, 0.83, 0.84, 0.88, 0.91, 0.9, 0.86, 0.87, 0.85, 
    0.87, 0.86, 0.85, 0.82, 0.78, 0.82, 0.81, 0.77, 0.74, 0.69, 0.66, 0.66, 
    0.63, 0.63, 0.6, 0.61, 0.61, 0.63, 0.61, 0.64, 0.66, 0.66, 0.65, 0.65, 
    0.67, 0.62, 0.6, 0.6, 0.6, 0.64, 0.83, 0.79, 0.9, 0.86, 0.83, 0.86, 0.69, 
    0.74, 0.72, 0.74, 0.63, 0.73, 0.74, 0.63, 0.59, 0.57, 0.65, 0.83, 0.76, 
    0.77, 0.66, 0.65, 0.62, 0.63, 0.68, 0.71, 0.79, 0.8, 0.81, 0.85, 0.85, 
    0.74, 0.85, 0.81, 0.84, 0.85, 0.86, 0.87, 0.88, 0.84, 0.69, 0.68, 0.69, 
    0.64, 0.61, 0.66, 0.69, 0.73, 0.87, 0.72, 0.7, 0.73, 0.7, 0.69, 0.71, 
    0.72, 0.76, 0.81, 0.85, 0.84, _, 0.83, 0.83, 0.83, 0.95, 0.94, 0.92, 
    0.92, 0.91, 0.94, 0.94, 0.95, 0.94, 0.96, 0.98, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.97, 0.93, 0.92, 0.93, 0.97, 0.98, 0.98, 0.98, 0.99, 
    0.99, 0.97, 0.96, 0.96, 0.94, 0.95, 0.94, 0.96, 0.95, 0.92, 0.95, 0.94, 
    0.95, 0.92, 0.85, 0.86, 0.82, 0.82, 0.86, 0.79, 0.81, 0.81, 0.8, 0.82, 
    0.8, 0.79, 0.78, 0.91, 0.94, 0.93, 0.97, 0.97, 0.97, 0.94, 0.93, 0.9, 
    0.92, 0.92, 0.92, 0.94, 0.9, 0.81, 0.79, 0.81, 0.89, 0.88, 0.95, 0.91, 
    0.85, 0.83, 0.84, 0.87, 0.84, 0.91, 0.94, 0.95, 0.95, 0.94, 0.93, 0.93, 
    0.95, 0.97, 0.96, 0.93, 0.88, 0.91, 0.93, 0.93, 0.94, 0.93, 0.93, 0.91, 
    0.93, 0.95, 0.91, 0.85, 0.87, 0.9, 0.87, 0.89, 0.89, 0.84, 0.89, 0.94, 
    0.92, 0.91, 0.87, 0.85, 0.86, 0.8, 0.8, 0.82, 0.86, 0.87, 0.88, 0.86, 
    0.85, 0.83, 0.84, 0.84, 0.85, 0.87, 0.91, 0.91, 0.93, 0.94, 0.95, 0.96, 
    0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.95, 0.94, 0.91, 0.89, 
    0.88, 0.86, 0.85, 0.84, 0.84, 0.83, 0.79, 0.78, 0.79, 0.83, 0.81, 0.81, 
    0.77, 0.75, 0.81, 0.78, 0.75, 0.71, 0.7, 0.72, 0.7, 0.7, 0.74, 0.73, 
    0.72, 0.73, 0.77, 0.86, 0.86, 0.67, 0.67, 0.68, 0.65, 0.66, 0.66, 0.69, 
    0.68, 0.68, 0.67, 0.67, 0.7, 0.67, 0.77, 0.76, 0.72, 0.66, 0.64, 0.64, 
    0.7, 0.68, 0.69, 0.66, 0.81, 0.84, 0.77, 0.62, 0.83, 0.79, 0.78, 0.82, 
    0.89, 0.91, 0.92, 0.91, 0.9, 0.87, 0.84, 0.8, 0.82, 0.83, 0.83, 0.79, 
    0.81, 0.82, 0.85, 0.81, 0.81, 0.8, 0.8, 0.78, 0.8, 0.82, 0.78, 0.8, 0.82, 
    0.79, 0.83, 0.83, 0.8, 0.83, 0.77, 0.74, 0.73, 0.73, 0.7, 0.73, 0.72, 
    0.73, 0.73, 0.8, 0.79, 0.8, 0.81, 0.7, 0.74, 0.79, 0.83, 0.87, 0.9, 0.87, 
    0.85, 0.85, 0.85, 0.89, 0.91, 0.88, 0.89, 0.87, 0.93, 0.95, 0.93, 0.92, 
    0.89, 0.86, 0.71, 0.77, 0.85, 0.9, 0.86, 0.88, 0.89, 0.9, 0.9, 0.94, 
    0.97, 0.98, 0.98, 0.96, 0.97, 0.98, 0.98, 0.93, 0.94, 0.94, 0.92, 0.93, 
    0.93, 0.93, 0.92, 0.91, 0.89, 0.87, 0.87, 0.82, 0.84, 0.84, 0.88, 0.89, 
    0.89, 0.9, 0.91, 0.92, 0.93, 0.95, 0.95, 0.96, 0.95, 0.96, 0.96, 0.96, 
    0.95, 0.96, 0.96, 0.97, 0.96, 0.93, 0.96, 0.97, 0.97, 0.98, 0.97, 0.94, 
    0.95, 0.94, 0.95, 0.95, 0.93, 0.97, 0.97, 0.96, 0.95, 0.96, 0.93, 0.95, 
    0.93, 0.94, 0.95, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 0.92, 0.91, 
    0.91, 0.87, 0.85, 0.86, 0.85, 0.85, 0.83, 0.82, 0.83, 0.81, 0.87, 0.9, 
    0.9, 0.88, 0.87, 0.85, 0.81, 0.82, 0.81, 0.78, 0.79, 0.75, 0.79, 0.8, 
    0.81, 0.82, 0.88, 0.89, 0.89, 0.93, 0.93, 0.91, 0.93, 0.93, 0.93, 0.91, 
    0.92, 0.9, 0.92, 0.92, 0.97, 0.97, 0.97, 0.96, 0.92, 0.89, 0.89, 0.9, 
    0.89, 0.9, 0.93, 0.96, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.94, 0.92, 
    0.92, 0.91, 0.91, 0.92, 0.94, 0.97, 0.96, 0.96, 0.96, 0.92, 0.9, 0.9, 
    0.91, 0.94, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.97, 0.92, 
    0.91, 0.92, 0.94, 0.95, 0.92, 0.91, 0.92, 0.92, 0.92, 0.95, 0.95, 0.94, 
    0.93, 0.95, 0.95, 0.93, 0.9, 0.95, 0.92, 0.96, 0.91, 0.89, 0.9, 0.93, 
    0.94, 0.95, 0.95, 0.95, 0.94, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.93, 
    0.92, 0.9, 0.9, 0.9, 0.92, 0.92, 0.93, 0.93, 0.93, 0.9, 0.9, 0.89, 0.87, 
    0.86, 0.85, 0.87, 0.86, 0.86, 0.85, 0.89, 0.83, 0.78, 0.72, 0.76, 0.83, 
    0.81, 0.82, 0.82, 0.84, 0.84, 0.83, 0.79, 0.81, 0.85, 0.78, 0.81, 0.86, 
    0.75, 0.79, 0.81, 0.82, 0.8, 0.85, 0.81, 0.78, 0.74, 0.72, 0.7, 0.77, 
    0.78, 0.82, 0.76, 0.73, 0.71, 0.74, 0.78, 0.76, 0.73, 0.73, 0.74, 0.71, 
    0.82, 0.81, 0.82, 0.84, 0.84, 0.83, 0.81, 0.82, 0.81, 0.81, 0.84, 0.8, 
    0.78, 0.83, 0.77, 0.77, 0.83, 0.84, 0.84, 0.8, 0.8, 0.81, 0.8, 0.78, 
    0.76, 0.74, 0.7, 0.61, 0.76, 0.72, 0.76, 0.75, 0.71, 0.67, 0.67, 0.81, 
    0.78, 0.75, 0.73, 0.75, 0.71, 0.74, 0.69, 0.75, 0.74, 0.77, 0.8, 0.86, 
    0.78, 0.77, 0.76, 0.79, 0.76, 0.81, 0.73, 0.8, 0.8, 0.73, 0.72, 0.72, 
    0.74, 0.76, 0.79, 0.76, 0.73, 0.72, 0.72, 0.73, 0.73, 0.74, 0.72, 0.74, 
    0.73, 0.75, 0.73, 0.74, 0.73, 0.73, 0.73, 0.74, 0.73, 0.72, 0.72, 0.73, 
    0.72, 0.72, 0.75, 0.74, 0.75, 0.77, 0.78, 0.8, 0.79, 0.8, 0.83, 0.86, 
    0.63, 0.67, 0.79, 0.7, 0.72, 0.76, 0.8, 0.8, 0.82, 0.91, 0.95, 0.95, 
    0.95, 0.97, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    1, 1, 1, 1, 0.99, 1, 0.99, 0.88, 0.87, 0.93, 0.96, 0.92, 0.88, 0.87, 
    0.84, 0.81, 0.81, 0.79, 0.79, 0.82, 0.82, 0.81, 0.8, 0.79, 0.8, 0.79, 
    0.81, 0.82, 0.82, 0.85, 0.86, 0.89, 0.88, 0.9, 0.91, 0.91, 0.93, 0.94, 
    0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.98, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.97, 0.93, 0.91, 0.92, 0.86, 0.85, 0.79, 0.76, 
    0.78, 0.75, 0.72, 0.71, 0.73, 0.69, 0.66, 0.73, 0.68, 0.64, 0.67, 0.67, 
    0.65, 0.66, 0.67, 0.68, 0.76, 0.89, 0.78, 0.76, 0.74, 0.72, 0.71, 0.77, 
    0.75, 0.77, 0.71, 0.74, 0.74, 0.75, 0.71, 0.76, 0.71, 0.72, 0.71, 0.68, 
    0.74, 0.73, 0.7, 0.75, 0.77, 0.76, 0.78, 0.79, 0.76, 0.82, 0.8, 0.82, 
    0.8, 0.79, 0.78, 0.72, 0.72, 0.75, 0.74, 0.71, 0.78, 0.72, 0.75, 0.86, 
    0.79, 0.77, 0.82, 0.82, 0.71, 0.69, 0.74, 0.73, 0.76, 0.7, 0.81, 0.83, 
    0.69, 0.72, 0.7, 0.72, 0.72, 0.74, 0.73, 0.74, 0.76, 0.76, 0.75, 0.76, 
    0.74, 0.74, 0.77, 0.77, 0.74, 0.78, 0.82, 0.87, 0.87, 0.87, 0.86, 0.8, 
    0.77, 0.74, 0.74, 0.76, 0.74, 0.77, 0.78, 0.72, 0.7, 0.72, 0.79, 0.74, 
    0.73, 0.72, 0.85, 0.75, 0.77, 0.78, 0.78, 0.77, 0.73, 0.76, 0.79, 0.72, 
    0.73, 0.74, 0.68, 0.68, 0.71, 0.7, 0.73, 0.73, 0.7, 0.73, 0.7, 0.75, 
    0.67, 0.71, 0.71, 0.7, 0.7, 0.7, 0.7, 0.75, 0.74, 0.65, 0.64, 0.75, 0.72, 
    0.69, 0.68, 0.71, 0.72, 0.7, 0.71, 0.75, 0.75, 0.75, 0.78, 0.72, 0.73, 
    0.73, 0.73, 0.71, 0.72, 0.75, 0.76, 0.74, 0.71, 0.68, 0.7, 0.69, 0.68, 
    0.67, 0.7, 0.7, 0.74, 0.78, 0.8, 0.81, 0.82, 0.84, 0.84, 0.88, 0.89, 
    0.86, 0.85, 0.86, 0.86, 0.85, 0.83, 0.82, 0.81, 0.82, 0.84, 0.85, 0.86, 
    0.87, 0.88, 0.88, 0.9, 0.9, 0.9, 0.89, 0.89, 0.9, 0.94, 0.93, 0.95, 0.92, 
    0.92, 0.93, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.95, 0.96, 0.96, 0.97, 
    0.98, 0.99, 0.97, 0.92, 0.94, 0.96, 0.97, 0.98, 0.93, 0.92, 0.91, 0.92, 
    0.94, 0.96, 0.93, 0.93, 0.91, 0.93, 0.94, 0.93, 0.88, 0.91, 0.91, 0.91, 
    0.94, 0.96, 0.95, 0.91, 0.91, 0.99, 0.98, 0.96, 0.91, 0.86, 0.89, 0.85, 
    0.8, 0.79, 0.78, 0.77, 0.76, 0.75, 0.81, 0.72, 0.84, 0.82, 0.74, 0.77, 
    0.78, 0.75, 0.84, 0.76, 0.75, 0.81, 0.83, 0.9, 0.77, 0.78, 0.9, 0.79, 
    0.75, 0.8, 0.83, 0.79, 0.75, 0.73, 0.68, 0.72, 0.71, 0.74, 0.73, 0.72, 
    0.74, 0.75, 0.75, 0.77, 0.74, 0.72, 0.7, 0.72, 0.76, 0.72, 0.73, 0.66, 
    0.67, 0.63, 0.64, 0.65, 0.67, 0.64, 0.68, 0.71, 0.7, 0.68, 0.68, 0.73, 
    0.72, 0.83, 0.69, 0.75, 0.78, 0.72, 0.77, 0.9, 0.89, 0.87, 0.87, 0.91, 
    0.8, 0.75, 0.81, 0.73, 0.88, 0.87, 0.85, 0.91, 0.81, 0.83, 0.8, 0.74, 
    0.72, 0.7, 0.77, 0.75, 0.76, 0.75, 0.74, 0.74, 0.78, 0.7, 0.7, 0.76, 
    0.73, 0.69, 0.71, 0.68, 0.68, 0.67, 0.68, 0.67, 0.66, 0.67, 0.67, 0.65, 
    0.69, 0.68, 0.73, 0.79, 0.81, 0.79, 0.77, 0.75, 0.74, 0.75, 0.74, 0.77, 
    0.84, 0.84, 0.78, 0.67, 0.75, 0.93, 0.7, 0.61, 0.7, 0.72, 0.67, 0.6, 
    0.58, 0.66, 0.72, 0.8, 0.78, 0.77, 0.73, 0.66, 0.73, 0.73, 0.77, 0.78, 
    0.77, 0.79, 0.83, 0.89, 0.96, 0.97, 0.96, 0.95, 0.94, 0.95, 0.96, 0.96, 
    0.96, 0.96, 0.95, 0.94, 0.95, 0.96, 0.97, 0.98, 0.97, 0.98, 0.98, 0.93, 
    0.91, 0.91, 0.89, 0.89, 0.87, 0.86, 0.88, 0.9, 0.89, 0.94, 0.94, 0.89, 
    0.92, 0.91, 0.96, 0.9, 0.9, 0.89, 0.86, 0.87, 0.8, 0.76, 0.78, 0.81, 
    0.81, 0.8, 0.76, 0.75, 0.68, 0.77, 0.8, 0.77, 0.73, 0.72, 0.8, 0.77, 
    0.79, 0.73, 0.77, 0.8, 0.74, 0.74, 0.74, 0.75, 0.75, 0.73, 0.73, 0.71, 
    0.68, 0.71, 0.73, 0.75, 0.74, 0.72, 0.74, 0.76, 0.72, 0.76, 0.76, 0.77, 
    0.77, 0.79, 0.76, 0.82, 0.8, 0.8, 0.77, 0.71, 0.77, 0.78, 0.79, 0.76, 
    0.73, 0.77, 0.73, 0.68, 0.81, 0.84, 0.81, 0.79, 0.79, 0.76, 0.74, 0.79, 
    0.78, 0.76, 0.74, 0.76, 0.75, 0.77, 0.77, 0.8, 0.77, 0.75, 0.75, 0.76, 
    0.73, 0.74, 0.75, 0.74, 0.72, 0.72, 0.75, 0.76, 0.73, 0.77, 0.76, 0.73, 
    0.72, 0.78, 0.73, 0.74, 0.72, 0.71, 0.7, 0.7, 0.71, 0.75, 0.76, 0.72, 
    0.73, 0.72, 0.79, 0.76, 0.81, 0.82, 0.78, 0.77, 0.71, 0.71, 0.69, 0.72, 
    0.72, 0.72, 0.73, 0.79, 0.81, 0.81, 0.81, 0.81, 0.77, 0.8, 0.73, 0.69, 
    0.73, 0.72, 0.75, 0.82, 0.79, 0.8, 0.77, 0.73, 0.7, 0.74, 0.68, 0.76, 
    0.72, 0.71, 0.7, 0.78, 0.79, 0.77, 0.76, 0.76, 0.81, 0.79, 0.78, 0.77, 
    0.74, 0.68, 0.67, 0.77, 0.73, 0.7, 0.64, 0.69, 0.66, 0.72, 0.72, 0.7, 
    0.69, 0.69, 0.83, 0.84, 0.81, 0.78, 0.75, 0.77, 0.77, 0.76, 0.76, 0.77, 
    0.82, 0.72, 0.76, 0.76, 0.79, 0.79, 0.77, 0.72, 0.71, 0.72, 0.77, 0.8, 
    0.89, 0.91, 0.87, 0.91, 0.88, 0.85, 0.94, 0.91, 0.94, 0.94, 0.94, 0.95, 
    0.93, 0.91, 0.91, 0.88, 0.87, 0.87, 0.85, 0.85, 0.82, 0.83, 0.82, 0.86, 
    0.79, 0.87, 0.87, 0.88, 0.89, 0.86, 0.82, 0.81, 0.76, 0.74, 0.78, 0.8, 
    0.81, 0.86, 0.83, 0.9, 0.8, 0.8, 0.9, 0.82, 0.79, 0.78, 0.75, 0.85, 0.87, 
    0.88, 0.85, 0.84, 0.89, 0.89, 0.88, 0.84, 0.87, 0.87, 0.87, 0.87, 0.91, 
    0.91, 0.92, 0.89, 0.89, 0.88, 0.89, 0.88, 0.83, 0.82, 0.79, 0.82, 0.83, 
    0.78, 0.83, 0.83, 0.84, 0.81, 0.8, 0.83, 0.83, 0.86, 0.84, 0.87, 0.88, 
    0.89, 0.9, 0.9, 0.87, 0.87, 0.84, 0.84, 0.81, 0.78, 0.82, 0.82, 0.79, 
    0.84, 0.82, 0.82, 0.82, 0.86, 0.81, 0.85, 0.87, 0.87, 0.9, 0.91, 0.91, 
    0.92, 0.92, 0.92, 0.91, 0.92, 0.9, 0.91, 0.9, 0.88, 0.86, 0.85, 0.86, 
    0.86, 0.87, 0.88, 0.89, 0.86, 0.88, 0.87, 0.86, 0.85, 0.85, 0.86, 0.85, 
    0.85, 0.84, 0.86, 0.85, 0.86, 0.85, 0.84, 0.85, 0.84, 0.86, 0.85, 0.86, 
    0.85, 0.85, 0.86, 0.85, 0.89, 0.93, 0.91, 0.94, 0.93, 0.94, 0.94, 0.97, 
    0.93, 0.88, 0.91, 0.94, 0.94, 0.97, 0.98, 0.93, 0.96, 0.95, 0.96, 0.96, 
    0.96, 0.95, 0.92, 0.92, 0.95, 0.97, 0.92, 0.95, 0.96, 0.93, 0.91, 0.92, 
    0.94, 0.96, 0.97, 0.97, 0.98, 0.98, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 
    0.99, 0.99, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.94, 0.95, 
    0.92, 0.96, 0.97, 0.97, 0.97, 0.96, 0.94, 0.96, 0.97, 0.96, 0.94, 0.93, 
    0.93, 0.93, 0.93, 0.92, 0.94, 0.93, 0.92, 0.92, 0.92, 0.92, 0.91, 0.93, 
    0.94, 0.92, 0.91, 0.91, 0.9, 0.9, 0.9, 0.89, 0.88, 0.88, 0.86, 0.85, 
    0.85, 0.84, 0.85, 0.86, 0.87, 0.85, 0.84, 0.8, 0.78, 0.82, 0.78, 0.75, 
    0.76, 0.74, 0.7, 0.72, 0.76, 0.78, 0.85, 0.88, 0.9, 0.94, 0.92, 0.89, 
    0.9, 0.9, 0.85, 0.86, 0.82, 0.89, 0.85, 0.87, 0.9, 0.84, 0.82, 0.86, 
    0.82, 0.81, 0.83, 0.82, 0.83, 0.83, 0.83, 0.82, 0.8, 0.79, 0.87, 0.8, 
    0.74, 0.75, 0.73, 0.72, 0.71, 0.82, 0.71, 0.62, 0.74, 0.63, 0.56, 0.7, 
    0.77, 0.75, 0.63, 0.59, 0.62, 0.64, 0.65, 0.62, 0.6, 0.71, 0.64, 0.79, 
    0.72, 0.68, 0.66, 0.69, 0.84, 0.59, 0.51, 0.47, 0.51, 0.52, 0.48, 0.5, 
    0.51, 0.58, 0.88, 0.71, 0.69, 0.64, 0.69, 0.64, 0.83, 0.72, 0.68, 0.7, 
    0.7, 0.63, 0.63, 0.81, 0.66, 0.63, 0.65, 0.65, 0.62, 0.64, 0.65, 0.62, 
    0.62, 0.65, 0.69, 0.79, 0.61, 0.55, 0.6, 0.69, 0.78, 0.83, 0.83, 0.86, 
    0.86, 0.83, 0.82, 0.81, 0.81, 0.77, 0.76, 0.72, 0.75, 0.75, 0.77, 0.82, 
    0.83, 0.83, 0.84, 0.87, 0.86, 0.85, 0.84, 0.86, 0.86, 0.85, 0.86, 0.85, 
    0.87, 0.88, 0.88, 0.84, 0.85, 0.83, 0.79, 0.83, 0.81, 0.85, 0.88, 0.94, 
    0.95, 0.91, 0.95, 0.94, 0.91, 0.91, 0.87, 0.85, 0.85, 0.87, 0.83, 0.89, 
    0.89, 0.87, 0.88, 0.91, 0.91, 0.92, 0.93, 0.93, 0.93, 0.89, 0.89, 0.9, 
    0.87, 0.88, 0.91, 0.97, 0.96, 0.95, 0.91, 0.91, 0.93, 0.95, 0.85, 0.86, 
    0.79, 0.73, 0.68, 0.67, 0.68, 0.7, 0.77, 0.76, 0.66, 0.69, 0.72, 0.79, 
    0.69, 0.88, 0.85, 0.83, 0.85, 0.86, 0.87, 0.86, 0.77, 0.81, 0.82, 0.87, 
    0.77, 0.86, 0.81, 0.84, 0.82, 0.83, 0.83, 0.84, 0.84, 0.85, 0.84, 0.82, 
    0.81, 0.84, 0.77, 0.78, 0.73, 0.75, 0.8, 0.71, 0.7, 0.68, 0.7, 0.66, 
    0.67, 0.71, 0.79, 0.64, 0.62, 0.65, 0.66, 0.67, 0.69, 0.7, 0.66, 0.69, 
    0.69, 0.72, 0.78, 0.77, 0.77, 0.84, 0.91, 0.93, 0.91, 0.94, 0.96, 0.97, 
    0.98, 0.98, 0.95, 0.94, 0.96, 0.96, 0.92, 0.92, 0.91, 0.97, 0.96, 0.95, 
    0.92, 0.87, 0.81, 0.79, 0.8, 0.78, 0.81, 0.84, 0.83, 0.84, 0.81, 0.82, 
    0.83, 0.8, 0.81, 0.8, 0.81, 0.8, 0.79, 0.8, 0.77, 0.78, 0.79, 0.78, 0.83, 
    0.85, 0.84, 0.81, 0.79, 0.85, 0.86, 0.84, 0.86, 0.84, 0.89, 0.9, 0.93, 
    0.94, 0.96, 0.97, 0.96, 0.96, 0.97, 0.97, 0.96, 0.97, 0.96, 0.95, 0.94, 
    0.95, 0.94, 0.94, 0.93, 0.92, 0.93, 0.93, 0.93, 0.93, 0.95, 0.95, 0.96, 
    0.92, 0.91, 0.88, 0.86, 0.86, 0.84, 0.84, 0.86, 0.86, 0.86, 0.86, 0.88, 
    0.9, 0.92, 0.91, 0.89, 0.94, 0.97, 0.98, 0.98, 0.98, 0.96, 0.94, 0.93, 
    0.92, 0.9, 0.88, 0.88, 0.83, 0.82, 0.82, 0.81, 0.78, 0.8, 0.81, 0.78, 
    0.8, 0.78, 0.71, 0.71, 0.76, 0.73, 0.67, 0.75, 0.74, 0.76, 0.69, 0.64, 
    0.68, 0.64, 0.7, 0.78, 0.63, 0.5, 0.82, 0.75, 0.69, 0.82, 0.59, 0.81, 
    0.76, 0.78, 0.78, 0.78, 0.79, 0.8, 0.82, 0.81, 0.81, 0.81, 0.8, 0.8, 0.8, 
    0.8, 0.77, 0.76, 0.78, 0.78, 0.78, 0.78, 0.78, 0.8, 0.79, 0.79, 0.78, 
    0.77, 0.76, 0.79, 0.76, 0.77, 0.79, 0.78, 0.79, 0.8, 0.8, 0.79, 0.81, 
    0.81, 0.81, 0.82, 0.81, 0.85, 0.82, 0.85, 0.88, 0.85, 0.83, 0.81, 0.86, 
    0.85, 0.83, 0.82, 0.81, 0.78, 0.82, 0.77, 0.8, 0.76, 0.76, 0.81, 0.73, 
    0.72, 0.72, 0.77, 0.74, 0.78, 0.71, 0.72, 0.74, 0.75, 0.75, 0.77, 0.71, 
    0.75, 0.73, 0.74, 0.66, 0.68, 0.74, 0.7, 0.75, 0.65, 0.66, 0.69, 0.71, 
    0.73, 0.66, 0.72, 0.7, 0.72, 0.73, 0.74, 0.68, 0.77, 0.79, 0.8, 0.8, 0.8, 
    0.79, 0.79, 0.76, 0.71, 0.6, 0.67, 0.67, 0.74, 0.75, 0.72, 0.74, 0.73, 
    0.72, 0.71, 0.75, 0.74, 0.71, 0.72, 0.75, 0.73, 0.72, 0.74, 0.69, 0.76, 
    0.77, 0.78, 0.77, 0.81, 0.84, 0.84, 0.84, 0.83, 0.81, 0.82, 0.81, 0.81, 
    0.81, 0.82, 0.81, 0.77, 0.83, 0.8, 0.83, 0.82, 0.8, 0.78, 0.77, 0.76, 
    0.76, 0.74, 0.8, 0.78, 0.78, 0.82, 0.8, 0.76, 0.78, 0.73, 0.68, 0.67, 
    0.68, 0.74, 0.72, 0.67, 0.67, 0.72, 0.67, 0.71, 0.77, 0.78, 0.75, 0.7, 
    0.74, 0.74, 0.63, 0.64, 0.67, 0.68, 0.66, 0.72, 0.75, 0.74, 0.76, 0.77, 
    0.78, 0.79, 0.8, 0.75, 0.81, 0.78, 0.8, 0.81, 0.8, 0.79, 0.74, 0.72, 
    0.73, 0.79, 0.78, 0.74, 0.76, 0.79, 0.77, 0.8, 0.81, 0.82, 0.81, 0.8, 
    0.77, 0.79, 0.79, 0.8, 0.72, 0.76, 0.75, 0.76, 0.78, 0.79, 0.8, 0.81, 
    0.83, 0.82, 0.8, 0.82, 0.81, 0.82, 0.8, 0.81, 0.82, 0.81, 0.75, 0.77, 
    0.77, 0.74, 0.74, 0.75, 0.73, 0.75, 0.75, 0.73, 0.75, 0.77, 0.79, 0.76, 
    0.79, 0.81, 0.79, 0.8, 0.8, 0.8, 0.81, 0.8, 0.74, 0.82, 0.81, 0.8, 0.81, 
    0.89, 0.79, 0.8, 0.85, 0.87, 0.81, 0.86, 0.85, 0.85, 0.85, 0.85, 0.83, 
    0.88, 0.87, 0.87, 0.87, 0.87, 0.87, 0.86, 0.82, 0.8, 0.83, 0.82, 0.82, 
    0.79, 0.77, 0.78, 0.77, 0.76, 0.79, 0.77, 0.76, 0.76, 0.75, 0.76, 0.76, 
    0.73, 0.75, 0.71, 0.72, 0.7, 0.68, 0.74, 0.72, 0.71, 0.73, 0.72, 0.71, 
    0.73, 0.74, 0.7, 0.71, 0.75, 0.73, 0.76, 0.79, 0.81, 0.83, 0.83, 0.81, 
    0.82, 0.79, 0.75, 0.73, 0.73, 0.72, 0.72, 0.73, 0.83, 0.86, 0.8, 0.84, 
    0.87, 0.87, 0.86, 0.86, 0.85, 0.84, 0.85, 0.84, 0.85, 0.85, 0.84, 0.81, 
    0.81, 0.8, 0.78, 0.81, 0.81, 0.81, 0.82, 0.78, 0.76, 0.76, 0.76, 0.77, 
    0.77, 0.77, 0.77, 0.77, 0.77, 0.77, 0.75, 0.75, 0.77, 0.76, 0.77, 0.77, 
    0.77, 0.75, 0.75, 0.74, 0.79, 0.85, 0.81, 0.74, 0.85, 0.87, 0.9, 0.91, 
    0.91, 0.91, 0.9, 0.9, 0.91, 0.9, 0.9, 0.89, 0.91, 0.91, 0.9, 0.89, 0.89, 
    0.89, 0.9, 0.9, 0.9, 0.9, 0.9, 0.89, 0.89, 0.88, 0.88, 0.87, 0.87, 0.87, 
    0.87, 0.86, 0.86, 0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 0.86, 0.86, 0.85, 
    0.84, 0.83, 0.83, 0.83, 0.82, 0.83, 0.83, 0.82, 0.82, 0.83, 0.83, 0.83, 
    0.83, 0.83, 0.84, 0.84, 0.82, 0.83, 0.84, 0.84, 0.84, 0.85, 0.84, 0.83, 
    0.83, 0.83, 0.82, 0.82, 0.82, 0.81, 0.82, 0.83, 0.82, 0.82, 0.82, 0.8, 
    0.8, 0.8, 0.8, 0.82, 0.81, 0.8, 0.8, 0.8, 0.79, 0.8, 0.81, 0.8, 0.79, 
    0.83, 0.83, 0.81, 0.83, 0.84, 0.82, 0.83, 0.84, 0.82, 0.81, 0.82, 0.81, 
    0.81, 0.81, 0.83, 0.83, 0.83, 0.82, 0.8, 0.8, 0.78, 0.76, 0.78, 0.81, 
    0.84, 0.84, 0.8, 0.79, 0.79, 0.8, 0.8, 0.78, 0.78, 0.77, 0.76, 0.77, 
    0.78, 0.77, 0.76, 0.77, 0.79, 0.78, 0.78, 0.79, 0.78, 0.77, 0.76, 0.76, 
    0.75, 0.76, 0.82, 0.79, 0.79, 0.78, 0.77, 0.77, 0.76, 0.76, 0.78, 0.77, 
    0.8, 0.79, 0.84, 0.77, 0.76, 0.75, 0.76, 0.75, 0.78, 0.8, 0.75, 0.76, 
    0.78, 0.82, 0.73, 0.72, 0.74, 0.76, 0.78, 0.78, 0.77, 0.78, 0.79, 0.77, 
    0.77, 0.77, 0.77, 0.78, 0.79, 0.8, 0.81, 0.8, 0.8, 0.73, 0.75, 0.74, 
    0.73, 0.73, 0.74, 0.75, 0.75, 0.75, 0.77, 0.76, 0.77, 0.72, 0.71, 0.72, 
    0.74, 0.74, 0.75, 0.75, 0.74, 0.76, 0.73, 0.77, 0.76, 0.75, 0.74, 0.76, 
    0.74, 0.75, 0.75, 0.71, 0.69, 0.78, 0.72, 0.74, 0.73, 0.73, 0.75, 0.75, 
    0.74, 0.71, 0.71, 0.73, 0.72, 0.69, 0.86, 0.73, 0.74, 0.76, 0.75, 0.75, 
    0.75, 0.74, 0.77, 0.76, 0.77, 0.75, 0.78, 0.74, 0.75, 0.76, 0.76, 0.77, 
    0.78, 0.77, 0.77, 0.75, 0.75, 0.75, 0.76, 0.79, 0.76, 0.76, 0.77, 0.78, 
    0.79, 0.8, 0.79, 0.78, 0.77, 0.77, 0.79, 0.79, 0.79, 0.78, 0.79, 0.79, 
    0.79, 0.78, 0.8, 0.79, 0.78, 0.78, 0.77, 0.78, 0.78, 0.78, 0.78, 0.77, 
    0.77, 0.76, 0.77, 0.77, 0.77, 0.75, 0.77, 0.76, 0.76, 0.77, 0.78, 0.79, 
    0.79, 0.79, 0.81, 0.83, 0.83, 0.82, 0.79, 0.76, 0.79, 0.77, 0.76, 0.76, 
    0.78, 0.77, 0.77, 0.74, 0.74, 0.74, 0.75, 0.75, 0.75, 0.74, 0.77, 0.75, 
    0.75, 0.75, 0.72, 0.73, 0.75, 0.71, 0.71, 0.72, 0.72, 0.69, 0.74, 0.72, 
    0.71, 0.75, 0.77, 0.78, 0.76, 0.78, 0.74, 0.78, 0.8, 0.85, 0.85, 0.86, 
    0.85, 0.69, 0.67, 0.76, 0.82, 0.83, 0.83, 0.85, 0.88, 0.84, 0.86, 0.84, 
    0.85, 0.86, 0.71, 0.78, 0.75, 0.73, 0.79, 0.8, 0.83, 0.84, 0.87, 0.88, 
    0.91, 0.91, 0.88, 0.88, 0.84, 0.82, 0.82, 0.86, 0.85, 0.81, 0.8, 0.82, 
    0.79, 0.7, 0.71, 0.78, 0.79, 0.74, 0.74, 0.71, 0.72, 0.71, 0.74, 0.75, 
    0.8, 0.83, 0.84, 0.84, 0.82, 0.8, 0.79, 0.8, 0.81, 0.8, 0.79, 0.79, 0.87, 
    0.88, 0.79, 0.85, 0.88, 0.89, 0.85, 0.83, 0.85, 0.89, 0.9, 0.88, 0.89, 
    0.83, 0.76, 0.78, 0.86, 0.87, 0.9, 0.89, 0.9, 0.92, 0.89, 0.84, 0.81, 
    0.79, 0.78, 0.81, 0.79, 0.77, 0.79, 0.81, 0.83, 0.85, 0.86, 0.82, 0.86, 
    0.9, 0.91, 0.92, 0.93, 0.94, 0.96, 0.94, 0.92, 0.91, 0.9, 0.91, 0.9, 
    0.84, 0.81, 0.75, 0.81, 0.84, 0.85, 0.81, 0.81, 0.69, 0.67, 0.74, 0.71, 
    0.84, 0.83, 0.81, 0.78, 0.7, 0.86, 0.85, 0.82, 0.82, 0.73, 0.76, 0.82, 
    0.8, 0.79, 0.78, 0.78, 0.77, 0.76, 0.81, 0.83, 0.83, 0.78, 0.78, 0.83, 
    0.87, 0.85, 0.86, 0.87, 0.88, 0.91, 0.89, 0.87, 0.85, 0.87, 0.85, 0.84, 
    0.84, 0.85, 0.85, 0.85, 0.84, 0.83, 0.84, 0.84, 0.86, 0.87, 0.86, 0.88, 
    0.89, 0.88, 0.85, 0.85, 0.82, 0.84, 0.83, 0.82, 0.83, 0.84, 0.82, 0.84, 
    0.84, 0.9, 0.94, 0.93, 0.93, 0.92, 0.92, 0.93, 0.93, 0.93, 0.91, 0.91, 
    0.9, 0.92, 0.94, 0.93, 0.91, 0.9, 0.91, 0.92, 0.92, 0.91, 0.91, 0.89, 
    0.89, 0.9, 0.9, 0.9, 0.89, 0.9, 0.91, 0.92, 0.92, 0.92, 0.91, 0.92, 0.91, 
    0.91, 0.88, 0.89, 0.87, 0.9, 0.9, 0.9, 0.88, 0.89, 0.9, 0.9, 0.88, 0.9, 
    0.93, 0.92, 0.89, 0.89, 0.9, 0.87, 0.9, 0.91, 0.89, 0.88, 0.9, 0.87, 
    0.87, 0.89, 0.9, 0.9, 0.9, 0.85, 0.86, 0.86, 0.86, 0.87, 0.91, 0.83, 
    0.87, 0.87, 0.89, 0.88, 0.89, 0.85, 0.86, 0.84, 0.81, 0.79, 0.8, 0.83, 
    0.81, 0.84, 0.82, 0.83, 0.85, 0.85, 0.83, 0.87, 0.85, 0.83, 0.85, 0.85, 
    0.79, 0.8, 0.85, 0.86, 0.87, 0.85, 0.9, 0.9, 0.84, 0.83, 0.85, 0.87, 
    0.79, 0.85, 0.85, 0.84, 0.84, 0.86, 0.85, 0.86, 0.82, 0.83, 0.83, 0.85, 
    0.85, 0.85, 0.85, 0.86, 0.85, 0.85, 0.85, 0.86, 0.86, 0.86, 0.85, 0.84, 
    0.86, 0.87, 0.87, 0.9, 0.91, 0.9, 0.89, 0.87, 0.86, 0.85, 0.88, 0.85, 
    0.85, 0.84, 0.86, 0.87, 0.94, 0.82, 0.8, 0.82, 0.84, 0.79, 0.8, 0.88, 
    0.8, 0.82, 0.84, 0.85, 0.81, 0.75, 0.72, 0.75, 0.78, 0.83, 0.79, 0.74, 
    0.73, 0.73, 0.8, 0.84, 0.8, 0.69, 0.71, 0.62, 0.72, 0.85, 0.87, 0.75, 
    0.75, 0.8, 0.83, 0.83, 0.83, 0.8, 0.75, 0.78, 0.82, 0.82, 0.82, 0.83, 
    0.84, 0.83, 0.84, 0.82, 0.81, 0.82, 0.79, 0.8, 0.8, 0.76, 0.78, 0.79, 
    0.8, 0.78, 0.78, 0.8, 0.8, 0.79, 0.8, 0.8, 0.8, 0.81, 0.85, 0.85, 0.85, 
    0.83, 0.85, 0.86, 0.86, 0.84, 0.83, 0.83, 0.81, 0.82, 0.82, 0.82, 0.81, 
    0.83, 0.82, 0.82, 0.82, 0.82, 0.83, 0.82, 0.83, 0.82, 0.8, 0.81, 0.82, 
    0.82, 0.83, 0.83, 0.84, 0.83, 0.84, 0.84, 0.88, 0.89, 0.9, 0.9, 0.9, 
    0.92, 0.94, 0.91, 0.9, 0.92, 0.92, 0.92, 0.91, 0.88, 0.89, 0.88, 0.92, 
    0.95, 0.93, 0.92, 0.91, 0.89, 0.88, 0.86, 0.86, 0.84, 0.83, 0.85, 0.82, 
    0.83, 0.82, 0.8, 0.8, 0.79, 0.79, 0.79, 0.79, 0.79, 0.75, 0.74, 0.74, 
    0.75, 0.74, 0.76, 0.77, 0.8, 0.82, 0.81, 0.81, 0.8, 0.8, 0.72, 0.8, 0.79, 
    0.78, 0.75, 0.76, 0.79, 0.72, 0.77, 0.79, 0.79, 0.81, 0.73, 0.75, 0.78, 
    0.74, 0.73, 0.7, 0.69, 0.66, 0.65, 0.75, 0.78, 0.79, 0.8, 0.74, 0.71, 
    0.7, 0.74, 0.73, 0.77, 0.78, 0.78, 0.81, 0.79, 0.81, 0.83, 0.81, 0.84, 
    0.83, 0.85, 0.9, 0.8, 0.81, 0.8, 0.82, 0.8, 0.75, 0.71, 0.7, 0.68, 0.68, 
    0.67, 0.68, 0.69, 0.69, 0.69, 0.74, 0.74, 0.75, 0.76, 0.77, 0.75, 0.72, 
    0.74, 0.73, 0.77, 0.76, 0.77, 0.77, 0.76, 0.76, 0.77, 0.74, 0.75, 0.77, 
    0.76, 0.77, 0.78, 0.8, 0.79, 0.8, 0.78, 0.79, 0.75, 0.74, 0.75, 0.74, 
    0.74, 0.72, 0.7, 0.69, 0.69, 0.71, 0.68, 0.66, 0.68, 0.71, 0.7, 0.69, 
    0.66, 0.67, 0.66, 0.67, 0.68, 0.67, 0.67, 0.67, 0.67, 0.67, 0.67, 0.68, 
    0.69, 0.69, 0.69, 0.68, 0.69, 0.69, 0.69, 0.7, 0.72, 0.7, 0.7, 0.71, 
    0.71, 0.71, 0.7, 0.7, 0.71, 0.73, 0.73, 0.73, 0.71, 0.7, 0.73, 0.73, 
    0.73, 0.72, 0.72, 0.72, 0.73, 0.73, 0.72, 0.73, 0.73, 0.74, 0.74, 0.75, 
    0.75, 0.75, 0.75, 0.75, 0.74, 0.76, 0.77, 0.77, 0.74, 0.74, 0.76, 0.76, 
    0.76, 0.75, 0.74, 0.75, 0.75, 0.76, 0.75, 0.74, 0.75, 0.75, 0.75, 0.74, 
    0.77, 0.78, 0.79, 0.79, 0.78, 0.8, 0.79, 0.77, 0.79, 0.8, 0.8, 0.79, 
    0.78, 0.78, 0.78, 0.77, 0.78, 0.79, 0.81, 0.83, 0.83, 0.8, 0.76, 0.75, 
    0.72, 0.79, 0.78, 0.83, 0.83, 0.82, 0.81, 0.81, 0.81, 0.81, 0.82, 0.82, 
    0.83, 0.82, 0.82, 0.83, 0.82, 0.84, 0.83, 0.84, 0.83, 0.77, 0.81, 0.78, 
    0.77, 0.8, 0.8, 0.8, 0.85, 0.84, 0.86, 0.88, 0.9, 0.9, 0.89, 0.91, 0.91, 
    0.91, 0.91, 0.94, 0.86, 0.87, 0.85, 0.85, 0.85, 0.82, 0.79, 0.85, 0.89, 
    0.9, 0.85, 0.83, 0.84, 0.83, 0.88, 0.87, 0.89, 0.9, 0.91, 0.9, 0.91, 
    0.88, 0.86, 0.84, 0.86, 0.82, 0.8, 0.79, 0.79, 0.77, 0.77, 0.8, 0.79, 
    0.78, 0.84, 0.76, 0.73, 0.74, 0.73, 0.72, 0.74, 0.73, 0.71, 0.7, 0.66, 
    0.64, 0.6, 0.63, 0.65, 0.67, 0.72, 0.81, 0.8, 0.79, 0.8, 0.82, 0.81, 
    0.78, 0.76, 0.76, 0.74, 0.74, 0.74, 0.73, 0.73, 0.71, 0.71, 0.71, 0.71, 
    0.71, 0.72, 0.69, 0.72, 0.72, 0.72, 0.7, 0.71, 0.71, 0.73, 0.72, 0.72, 
    0.74, 0.74, 0.75, 0.77, 0.78, 0.76, 0.76, 0.75, 0.77, 0.76, 0.74, 0.76, 
    0.76, 0.76, 0.78, 0.79, 0.78, 0.78, 0.78, 0.77, 0.76, 0.77, 0.76, 0.77, 
    0.76, 0.76, 0.76, 0.76, 0.78, 0.77, 0.78, 0.78, 0.78, 0.78, 0.79, 0.79, 
    0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.8, 0.79, 
    0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.79, 0.78, 0.77, 
    0.77, 0.77, 0.77, 0.76, 0.75, 0.74, 0.74, 0.75, 0.76, 0.75, 0.75, 0.74, 
    0.74, 0.75, 0.77, 0.78, 0.77, 0.78, 0.77, 0.77, 0.78, 0.79, 0.78, 0.75, 
    0.76, 0.79, 0.79, 0.79, 0.79, 0.77, 0.8, 0.8, 0.8, 0.8, 0.81, 0.79, 0.8, 
    0.77, 0.78, 0.78, 0.77, 0.75, 0.73, 0.74, 0.73, 0.74, 0.74, 0.74, 0.74, 
    0.76, 0.76, 0.76 ;
}
