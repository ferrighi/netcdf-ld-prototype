netcdf SN99880 {
dimensions:
	time = UNLIMITED ; // (59360 currently)
	station_id = 7 ;
variables:
	double time(time) ;
		time:standard_name = "time" ;
		time:long_name = "Time of measurement" ;
		time:calendar = "standard" ;
		time:units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:axis = "T" ;
	double latitude ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:units = "degree_north" ;
	double longitude ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:units = "degree_east" ;
	char station_id(station_id) ;
		station_id:cf_role = "timeseries_id" ;
	float air_temperature_2m(time) ;
		air_temperature_2m:long_name = "Air temperature" ;
		air_temperature_2m:coverage_content_type = "coordinate" ;
		air_temperature_2m:standard_name = "air_temperature" ;
		air_temperature_2m:units = "K" ;
	float air_pressure_at_sea_level(time) ;
		air_pressure_at_sea_level:long_name = "Air pressure at sea level" ;
		air_pressure_at_sea_level:coverage_content_type = "coordinate" ;
		air_pressure_at_sea_level:standard_name = "air_pressure_at_sea_level" ;
		air_pressure_at_sea_level:units = "Pa" ;
	float air_pressure_at_sea_level_qnh(time) ;
		air_pressure_at_sea_level_qnh:long_name = "Air pressure (QNH)" ;
		air_pressure_at_sea_level_qnh:coverage_content_type = "coordinate" ;
		air_pressure_at_sea_level_qnh:standard_name = "air_pressure_at_sea_level_qnh" ;
		air_pressure_at_sea_level_qnh:units = "hPa" ;
	float wind_speed_10m(time) ;
		wind_speed_10m:long_name = "Mean wind speed" ;
		wind_speed_10m:coverage_content_type = "coordinate" ;
		wind_speed_10m:standard_name = "wind_speed" ;
		wind_speed_10m:units = "m s-1" ;
	float relative_humidity(time) ;
		relative_humidity:long_name = "Relative air humidity" ;
		relative_humidity:coverage_content_type = "coordinate" ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:units = "1" ;
	float surface_air_pressure_2m(time) ;
		surface_air_pressure_2m:long_name = "Air pressure at station level" ;
		surface_air_pressure_2m:coverage_content_type = "coordinate" ;
		surface_air_pressure_2m:standard_name = "surface_air_pressure" ;
		surface_air_pressure_2m:units = "Pa" ;
	float wind_from_direction_10m(time) ;
		wind_from_direction_10m:long_name = "Wind direction" ;
		wind_from_direction_10m:coverage_content_type = "coordinate" ;
		wind_from_direction_10m:standard_name = "wind_from_direction" ;
		wind_from_direction_10m:units = "degree" ;

// global attributes:
		:station_name = "PYRAMIDEN" ;
		:wigos_identifier = "0-20000-0-01024" ;
		:wmo_identifier = "01024" ;
		:date_created = "2019-09-03T09:58:12.415858+00:00" ;
		:Conventions = "ACDD-1.3 CF-1.6" ;
		:title = "Observations from station PYRAMIDEN SN99880" ;
		:institution = "Norwegian Meteorological Institute" ;
		:source = "Meterological surface observation via frost.met.no" ;
		//:history = "2019-09-03T09:58:12.415858+00:00: frost write netcdf" ;
		:history = "https://github.com/ferrighi/netcdf-ld-prototype/blob/master/files/data-provenance-sios.ttl" ; 
		:references = "" ;
		:acknowledgment = "frost.met.no" ;
		:comment = "Observations based on data from frost.met.no" ;
		:creator_email = "observasjon@met.no" ;
		:creator_name = "Norwegian Meteorological Institute" ;
		:creator_url = "https://met.no" ;
		:geospatial_bounds = "POINT(16.360300 78.655700)" ;
		:geospatial_bounds_crs = "latlon" ;
		:geospatial_lat_max = "78.655700" ;
		:geospatial_lat_min = "78.655700" ;
		:geospatial_lon_max = "16.360300" ;
		:geospatial_lon_min = "16.360300" ;
		:id = "metno_obs_SN99880" ;
		:keywords = "observations" ;
		:metadata_link = "https://oaipmh.met.no/oai/?verb=GetRecord&metadataPrefix=iso&identifier=SN99880" ;
		:summary = "Surface meteorological observations from the observation network operated by the Norwegian Meteorological Institute. Data are received and quality controlled using the local KVALOBS system. Observation stations are normally operated according to WMO requirements, although specifications are not followed on some remote stations for practical matters. Stations may have more parameters than reported in this dataset." ;
		:time_coverage_start = "2012-11-16T10:00:00" ;
		:time_coverage_end = "2019-09-03T10:00:00" ;
		:featureType = "timeSeries" ;
data:

 time = 1353060000, 1353063600, 1353067200, 1353070800, 1353074400, 
    1353078000, 1353081600, 1353085200, 1353088800, 1353092400, 1353096000, 
    1353099600, 1353103200, 1353106800, 1353110400, 1353114000, 1353117600, 
    1353121200, 1353124800, 1353128400, 1353132000, 1353135600, 1353139200, 
    1353142800, 1353146400, 1353150000, 1353153600, 1353157200, 1353160800, 
    1353164400, 1353168000, 1353171600, 1353175200, 1353178800, 1353182400, 
    1353186000, 1353189600, 1353193200, 1353196800, 1353200400, 1353204000, 
    1353207600, 1353211200, 1353214800, 1353218400, 1353222000, 1353225600, 
    1353229200, 1353232800, 1353236400, 1353240000, 1353243600, 1353247200, 
    1353250800, 1353254400, 1353258000, 1353261600, 1353265200, 1353268800, 
    1353272400, 1353276000, 1353279600, 1353283200, 1353286800, 1353290400, 
    1353294000, 1353297600, 1353301200, 1353304800, 1353308400, 1353312000, 
    1353315600, 1353319200, 1353322800, 1353326400, 1353330000, 1353333600, 
    1353337200, 1353340800, 1353344400, 1353348000, 1353351600, 1353355200, 
    1353358800, 1353362400, 1353366000, 1353369600, 1353373200, 1353376800, 
    1353380400, 1353384000, 1353387600, 1353391200, 1353394800, 1353398400, 
    1353402000, 1353405600, 1353409200, 1353412800, 1353416400, 1353420000, 
    1353423600, 1353427200, 1353430800, 1353434400, 1353438000, 1353441600, 
    1353445200, 1353448800, 1353452400, 1353456000, 1353459600, 1353463200, 
    1353466800, 1353470400, 1353474000, 1353477600, 1353481200, 1353484800, 
    1353488400, 1353492000, 1353495600, 1353499200, 1353502800, 1353506400, 
    1353510000, 1353513600, 1353517200, 1353520800, 1353524400, 1353528000, 
    1353531600, 1353535200, 1353538800, 1353542400, 1353546000, 1353549600, 
    1353553200, 1353556800, 1353560400, 1353564000, 1353567600, 1353571200, 
    1353574800, 1353578400, 1353582000, 1353585600, 1353589200, 1353592800, 
    1353596400, 1353600000, 1353603600, 1353607200, 1353610800, 1353614400, 
    1353618000, 1353621600, 1353625200, 1353628800, 1353632400, 1353636000, 
    1353639600, 1353643200, 1353646800, 1353650400, 1353654000, 1353657600, 
    1353661200, 1353664800, 1353668400, 1353672000, 1353675600, 1353679200, 
    1353682800, 1353686400, 1353690000, 1353693600, 1353697200, 1353700800, 
    1353704400, 1353708000, 1353711600, 1353715200, 1353718800, 1353722400, 
    1353726000, 1353729600, 1353733200, 1353736800, 1353740400, 1353744000, 
    1353747600, 1353751200, 1353754800, 1353758400, 1353762000, 1353765600, 
    1353769200, 1353772800, 1353776400, 1353780000, 1353783600, 1353787200, 
    1353790800, 1353794400, 1353798000, 1353801600, 1353805200, 1353808800, 
    1353812400, 1353816000, 1353819600, 1353823200, 1353826800, 1353830400, 
    1353834000, 1353837600, 1353841200, 1353844800, 1353848400, 1353852000, 
    1353855600, 1353859200, 1353862800, 1353866400, 1353870000, 1353873600, 
    1353877200, 1353880800, 1353884400, 1353888000, 1353891600, 1353895200, 
    1353898800, 1353902400, 1353906000, 1353909600, 1353913200, 1353916800, 
    1353920400, 1353924000, 1353927600, 1353931200, 1353934800, 1353938400, 
    1353942000, 1353945600, 1353949200, 1353952800, 1353956400, 1353960000, 
    1353963600, 1353967200, 1353970800, 1353974400, 1353978000, 1353981600, 
    1353985200, 1353988800, 1353992400, 1353996000, 1353999600, 1354003200, 
    1354006800, 1354010400, 1354014000, 1354017600, 1354021200, 1354024800, 
    1354028400, 1354032000, 1354035600, 1354039200, 1354042800, 1354046400, 
    1354050000, 1354053600, 1354057200, 1354060800, 1354064400, 1354068000, 
    1354071600, 1354075200, 1354078800, 1354082400, 1354086000, 1354089600, 
    1354093200, 1354096800, 1354100400, 1354104000, 1354107600, 1354111200, 
    1354114800, 1354118400, 1354122000, 1354125600, 1354129200, 1354132800, 
    1354136400, 1354140000, 1354143600, 1354147200, 1354150800, 1354154400, 
    1354158000, 1354161600, 1354165200, 1354168800, 1354172400, 1354176000, 
    1354179600, 1354183200, 1354186800, 1354190400, 1354194000, 1354197600, 
    1354201200, 1354204800, 1354208400, 1354212000, 1354215600, 1354219200, 
    1354222800, 1354226400, 1354230000, 1354233600, 1354237200, 1354240800, 
    1354244400, 1354248000, 1354251600, 1354255200, 1354258800, 1354262400, 
    1354266000, 1354269600, 1354273200, 1354276800, 1354280400, 1354284000, 
    1354287600, 1354291200, 1354294800, 1354298400, 1354302000, 1354305600, 
    1354309200, 1354312800, 1354316400, 1354320000, 1354323600, 1354327200, 
    1354330800, 1354334400, 1354338000, 1354341600, 1354345200, 1354348800, 
    1354352400, 1354356000, 1354359600, 1354363200, 1354366800, 1354370400, 
    1354374000, 1354377600, 1354381200, 1354384800, 1354388400, 1354392000, 
    1354395600, 1354399200, 1354402800, 1354406400, 1354410000, 1354413600, 
    1354417200, 1354420800, 1354424400, 1354428000, 1354431600, 1354435200, 
    1354438800, 1354442400, 1354446000, 1354449600, 1354453200, 1354456800, 
    1354460400, 1354464000, 1354467600, 1354471200, 1354474800, 1354478400, 
    1354482000, 1354485600, 1354489200, 1354492800, 1354496400, 1354500000, 
    1354503600, 1354507200, 1354510800, 1354514400, 1354518000, 1354521600, 
    1354525200, 1354528800, 1354532400, 1354536000, 1354539600, 1354543200, 
    1354546800, 1354550400, 1354554000, 1354557600, 1354561200, 1354564800, 
    1354568400, 1354572000, 1354575600, 1354579200, 1354582800, 1354586400, 
    1354590000, 1354593600, 1354597200, 1354600800, 1354604400, 1354608000, 
    1354611600, 1354615200, 1354618800, 1354622400, 1354626000, 1354629600, 
    1354633200, 1354636800, 1354640400, 1354644000, 1354647600, 1354651200, 
    1354654800, 1354658400, 1354662000, 1354665600, 1354669200, 1354672800, 
    1354676400, 1354680000, 1354683600, 1354687200, 1354690800, 1354694400, 
    1354698000, 1354701600, 1354705200, 1354708800, 1354712400, 1354716000, 
    1354719600, 1354723200, 1354726800, 1354730400, 1354734000, 1354737600, 
    1354741200, 1354744800, 1354748400, 1354752000, 1354755600, 1354759200, 
    1354762800, 1354766400, 1354770000, 1354773600, 1354777200, 1354780800, 
    1354784400, 1354788000, 1354791600, 1354795200, 1354798800, 1354802400, 
    1354806000, 1354809600, 1354813200, 1354816800, 1354820400, 1354824000, 
    1354827600, 1354831200, 1354834800, 1354838400, 1354842000, 1354845600, 
    1354849200, 1354852800, 1354856400, 1354860000, 1354863600, 1354867200, 
    1354870800, 1354874400, 1354878000, 1354881600, 1354885200, 1354888800, 
    1354892400, 1354896000, 1354899600, 1354903200, 1354906800, 1354910400, 
    1354914000, 1354917600, 1354921200, 1354924800, 1354928400, 1354932000, 
    1354935600, 1354939200, 1354942800, 1354946400, 1354950000, 1354953600, 
    1354957200, 1354960800, 1354964400, 1354968000, 1354971600, 1354975200, 
    1354978800, 1354982400, 1354986000, 1354989600, 1354993200, 1354996800, 
    1355000400, 1355004000, 1355007600, 1355011200, 1355014800, 1355018400, 
    1355022000, 1355025600, 1355029200, 1355032800, 1355036400, 1355040000, 
    1355043600, 1355047200, 1355050800, 1355054400, 1355058000, 1355061600, 
    1355065200, 1355068800, 1355072400, 1355076000, 1355079600, 1355083200, 
    1355086800, 1355090400, 1355094000, 1355097600, 1355101200, 1355104800, 
    1355108400, 1355112000, 1355115600, 1355119200, 1355122800, 1355126400, 
    1355130000, 1355133600, 1355137200, 1355140800, 1355144400, 1355148000, 
    1355151600, 1355155200, 1355158800, 1355162400, 1355166000, 1355169600, 
    1355173200, 1355176800, 1355180400, 1355184000, 1355187600, 1355191200, 
    1355194800, 1355198400, 1355202000, 1355205600, 1355209200, 1355212800, 
    1355216400, 1355220000, 1355223600, 1355227200, 1355230800, 1355234400, 
    1355238000, 1355241600, 1355245200, 1355248800, 1355252400, 1355256000, 
    1355259600, 1355263200, 1355266800, 1355270400, 1355274000, 1355277600, 
    1355281200, 1355284800, 1355288400, 1355292000, 1355295600, 1355299200, 
    1355302800, 1355306400, 1355310000, 1355313600, 1355317200, 1355320800, 
    1355324400, 1355328000, 1355331600, 1355335200, 1355338800, 1355342400, 
    1355346000, 1355349600, 1355353200, 1355356800, 1355360400, 1355364000, 
    1355367600, 1355371200, 1355374800, 1355378400, 1355382000, 1355385600, 
    1355389200, 1355392800, 1355396400, 1355400000, 1355403600, 1355407200, 
    1355410800, 1355414400, 1355418000, 1355421600, 1355425200, 1355428800, 
    1355432400, 1355436000, 1355439600, 1355443200, 1355446800, 1355450400, 
    1355454000, 1355457600, 1355461200, 1355464800, 1355468400, 1355472000, 
    1355475600, 1355479200, 1355482800, 1355486400, 1355490000, 1355493600, 
    1355497200, 1355500800, 1355504400, 1355508000, 1355511600, 1355515200, 
    1355518800, 1355522400, 1355526000, 1355529600, 1355533200, 1355536800, 
    1355540400, 1355544000, 1355547600, 1355551200, 1355554800, 1355558400, 
    1355562000, 1355565600, 1355569200, 1355572800, 1355576400, 1355580000, 
    1355583600, 1355587200, 1355590800, 1355594400, 1355598000, 1355601600, 
    1355605200, 1355608800, 1355612400, 1355616000, 1355619600, 1355623200, 
    1355626800, 1355630400, 1355634000, 1355637600, 1355641200, 1355644800, 
    1355648400, 1355652000, 1355655600, 1355659200, 1355662800, 1355666400, 
    1355670000, 1355673600, 1355677200, 1355680800, 1355684400, 1355688000, 
    1355691600, 1355695200, 1355698800, 1355702400, 1355706000, 1355709600, 
    1355713200, 1355716800, 1355720400, 1355724000, 1355727600, 1355731200, 
    1355734800, 1355738400, 1355742000, 1355745600, 1355749200, 1355752800, 
    1355756400, 1355760000, 1355763600, 1355767200, 1355770800, 1355774400, 
    1355778000, 1355781600, 1355785200, 1355788800, 1355792400, 1355796000, 
    1355799600, 1355803200, 1355806800, 1355810400, 1355814000, 1355817600, 
    1355821200, 1355824800, 1355828400, 1355832000, 1355835600, 1355839200, 
    1355842800, 1355846400, 1355850000, 1355853600, 1355857200, 1355860800, 
    1355864400, 1355868000, 1355871600, 1355875200, 1355878800, 1355882400, 
    1355886000, 1355889600, 1355893200, 1355896800, 1355900400, 1355904000, 
    1355907600, 1355911200, 1355914800, 1355918400, 1355922000, 1355925600, 
    1355929200, 1355932800, 1355936400, 1355940000, 1355943600, 1355947200, 
    1355950800, 1355954400, 1355958000, 1355961600, 1355965200, 1355968800, 
    1355972400, 1355976000, 1355979600, 1355983200, 1355986800, 1355990400, 
    1355994000, 1355997600, 1356001200, 1356004800, 1356008400, 1356012000, 
    1356015600, 1356019200, 1356022800, 1356026400, 1356030000, 1356033600, 
    1356037200, 1356040800, 1356044400, 1356048000, 1356051600, 1356055200, 
    1356058800, 1356062400, 1356066000, 1356069600, 1356073200, 1356076800, 
    1356080400, 1356084000, 1356087600, 1356091200, 1356094800, 1356098400, 
    1356102000, 1356105600, 1356109200, 1356112800, 1356116400, 1356120000, 
    1356123600, 1356127200, 1356130800, 1356134400, 1356138000, 1356141600, 
    1356145200, 1356148800, 1356152400, 1356156000, 1356159600, 1356163200, 
    1356166800, 1356170400, 1356174000, 1356177600, 1356181200, 1356184800, 
    1356188400, 1356192000, 1356195600, 1356199200, 1356202800, 1356206400, 
    1356210000, 1356213600, 1356217200, 1356220800, 1356224400, 1356228000, 
    1356231600, 1356235200, 1356238800, 1356242400, 1356246000, 1356249600, 
    1356253200, 1356256800, 1356260400, 1356264000, 1356267600, 1356271200, 
    1356274800, 1356278400, 1356282000, 1356285600, 1356289200, 1356292800, 
    1356296400, 1356300000, 1356303600, 1356307200, 1356310800, 1356314400, 
    1356318000, 1356321600, 1356325200, 1356328800, 1356332400, 1356336000, 
    1356339600, 1356343200, 1356346800, 1356350400, 1356354000, 1356357600, 
    1356361200, 1356364800, 1356368400, 1356372000, 1356375600, 1356379200, 
    1356382800, 1356386400, 1356390000, 1356393600, 1356397200, 1356400800, 
    1356404400, 1356408000, 1356411600, 1356415200, 1356418800, 1356422400, 
    1356426000, 1356429600, 1356433200, 1356436800, 1356440400, 1356444000, 
    1356447600, 1356451200, 1356454800, 1356458400, 1356462000, 1356465600, 
    1356469200, 1356472800, 1356476400, 1356480000, 1356483600, 1356487200, 
    1356490800, 1356494400, 1356498000, 1356501600, 1356505200, 1356508800, 
    1356512400, 1356516000, 1356519600, 1356523200, 1356526800, 1356530400, 
    1356534000, 1356537600, 1356541200, 1356544800, 1356548400, 1356552000, 
    1356555600, 1356559200, 1356562800, 1356566400, 1356570000, 1356573600, 
    1356577200, 1356580800, 1356584400, 1356588000, 1356591600, 1356595200, 
    1356598800, 1356602400, 1356606000, 1356609600, 1356613200, 1356616800, 
    1356620400, 1356624000, 1356627600, 1356631200, 1356634800, 1356638400, 
    1356642000, 1356645600, 1356649200, 1356652800, 1356656400, 1356660000, 
    1356663600, 1356667200, 1356670800, 1356674400, 1356678000, 1356681600, 
    1356685200, 1356688800, 1356692400, 1356696000, 1356699600, 1356703200, 
    1356706800, 1356710400, 1356714000, 1356717600, 1356721200, 1356724800, 
    1356728400, 1356732000, 1356735600, 1356739200, 1356742800, 1356746400, 
    1356750000, 1356753600, 1356757200, 1356760800, 1356764400, 1356768000, 
    1356771600, 1356775200, 1356778800, 1356782400, 1356786000, 1356789600, 
    1356793200, 1356796800, 1356800400, 1356804000, 1356807600, 1356811200, 
    1356814800, 1356818400, 1356822000, 1356825600, 1356829200, 1356832800, 
    1356836400, 1356840000, 1356843600, 1356847200, 1356850800, 1356854400, 
    1356858000, 1356861600, 1356865200, 1356868800, 1356872400, 1356876000, 
    1356879600, 1356883200, 1356886800, 1356890400, 1356894000, 1356897600, 
    1356901200, 1356904800, 1356908400, 1356912000, 1356915600, 1356919200, 
    1356922800, 1356926400, 1356930000, 1356933600, 1356937200, 1356940800, 
    1356944400, 1356948000, 1356951600, 1356955200, 1356958800, 1356962400, 
    1356966000, 1356969600, 1356973200, 1356976800, 1356980400, 1356984000, 
    1356987600, 1356991200, 1356994800, 1356998400, 1357002000, 1357005600, 
    1357009200, 1357012800, 1357016400, 1357020000, 1357023600, 1357027200, 
    1357030800, 1357034400, 1357038000, 1357041600, 1357045200, 1357048800, 
    1357052400, 1357056000, 1357059600, 1357063200, 1357066800, 1357070400, 
    1357074000, 1357077600, 1357081200, 1357084800, 1357088400, 1357092000, 
    1357095600, 1357099200, 1357102800, 1357106400, 1357110000, 1357113600, 
    1357117200, 1357120800, 1357124400, 1357128000, 1357131600, 1357135200, 
    1357138800, 1357142400, 1357146000, 1357149600, 1357153200, 1357156800, 
    1357160400, 1357164000, 1357167600, 1357171200, 1357174800, 1357178400, 
    1357182000, 1357185600, 1357189200, 1357192800, 1357196400, 1357200000, 
    1357203600, 1357207200, 1357210800, 1357214400, 1357218000, 1357221600, 
    1357225200, 1357228800, 1357232400, 1357236000, 1357239600, 1357243200, 
    1357246800, 1357250400, 1357254000, 1357257600, 1357261200, 1357264800, 
    1357268400, 1357272000, 1357275600, 1357279200, 1357282800, 1357286400, 
    1357290000, 1357293600, 1357297200, 1357300800, 1357304400, 1357308000, 
    1357311600, 1357315200, 1357318800, 1357322400, 1357326000, 1357329600, 
    1357333200, 1357336800, 1357340400, 1357344000, 1357347600, 1357351200, 
    1357354800, 1357358400, 1357362000, 1357365600, 1357369200, 1357372800, 
    1357376400, 1357380000, 1357383600, 1357387200, 1357390800, 1357394400, 
    1357398000, 1357401600, 1357405200, 1357408800, 1357412400, 1357416000, 
    1357419600, 1357423200, 1357426800, 1357430400, 1357434000, 1357437600, 
    1357441200, 1357444800, 1357448400, 1357452000, 1357455600, 1357459200, 
    1357462800, 1357466400, 1357470000, 1357473600, 1357477200, 1357480800, 
    1357484400, 1357488000, 1357491600, 1357495200, 1357498800, 1357502400, 
    1357506000, 1357509600, 1357513200, 1357516800, 1357520400, 1357524000, 
    1357527600, 1357531200, 1357534800, 1357538400, 1357542000, 1357545600, 
    1357549200, 1357552800, 1357556400, 1357560000, 1357563600, 1357567200, 
    1357570800, 1357574400, 1357578000, 1357581600, 1357585200, 1357588800, 
    1357592400, 1357596000, 1357599600, 1357603200, 1357606800, 1357610400, 
    1357614000, 1357617600, 1357621200, 1357624800, 1357628400, 1357632000, 
    1357635600, 1357639200, 1357642800, 1357646400, 1357650000, 1357653600, 
    1357657200, 1357660800, 1357664400, 1357668000, 1357671600, 1357675200, 
    1357678800, 1357682400, 1357686000, 1357689600, 1357693200, 1357696800, 
    1357700400, 1357704000, 1357707600, 1357711200, 1357714800, 1357718400, 
    1357722000, 1357725600, 1357729200, 1357732800, 1357736400, 1357740000, 
    1357743600, 1357747200, 1357750800, 1357754400, 1357758000, 1357761600, 
    1357765200, 1357768800, 1357772400, 1357776000, 1357779600, 1357783200, 
    1357786800, 1357790400, 1357794000, 1357797600, 1357801200, 1357804800, 
    1357808400, 1357812000, 1357815600, 1357819200, 1357822800, 1357826400, 
    1357830000, 1357833600, 1357837200, 1357840800, 1357844400, 1357848000, 
    1357851600, 1357855200, 1357858800, 1357862400, 1357866000, 1357869600, 
    1357873200, 1357876800, 1357880400, 1357884000, 1357887600, 1357891200, 
    1357894800, 1357898400, 1357902000, 1357905600, 1357909200, 1357912800, 
    1357916400, 1357920000, 1357923600, 1357927200, 1357930800, 1357934400, 
    1357938000, 1357941600, 1357945200, 1357948800, 1357952400, 1357956000, 
    1357959600, 1357963200, 1357966800, 1357970400, 1357974000, 1357977600, 
    1357981200, 1357984800, 1357988400, 1357992000, 1357995600, 1357999200, 
    1358002800, 1358006400, 1358010000, 1358013600, 1358017200, 1358020800, 
    1358024400, 1358028000, 1358031600, 1358035200, 1358038800, 1358042400, 
    1358046000, 1358049600, 1358053200, 1358056800, 1358060400, 1358064000, 
    1358067600, 1358071200, 1358074800, 1358078400, 1358082000, 1358085600, 
    1358089200, 1358092800, 1358096400, 1358100000, 1358103600, 1358107200, 
    1358110800, 1358114400, 1358118000, 1358121600, 1358125200, 1358128800, 
    1358132400, 1358136000, 1358139600, 1358143200, 1358146800, 1358150400, 
    1358154000, 1358157600, 1358161200, 1358164800, 1358168400, 1358172000, 
    1358175600, 1358179200, 1358182800, 1358186400, 1358190000, 1358193600, 
    1358197200, 1358200800, 1358204400, 1358208000, 1358211600, 1358215200, 
    1358218800, 1358222400, 1358226000, 1358229600, 1358233200, 1358236800, 
    1358240400, 1358244000, 1358247600, 1358251200, 1358254800, 1358258400, 
    1358262000, 1358265600, 1358269200, 1358272800, 1358276400, 1358280000, 
    1358283600, 1358287200, 1358290800, 1358294400, 1358298000, 1358301600, 
    1358305200, 1358308800, 1358312400, 1358316000, 1358319600, 1358323200, 
    1358326800, 1358330400, 1358334000, 1358337600, 1358341200, 1358344800, 
    1358348400, 1358352000, 1358355600, 1358359200, 1358362800, 1358366400, 
    1358370000, 1358373600, 1358377200, 1358380800, 1358384400, 1358388000, 
    1358391600, 1358395200, 1358398800, 1358402400, 1358406000, 1358409600, 
    1358413200, 1358416800, 1358420400, 1358424000, 1358427600, 1358431200, 
    1358434800, 1358438400, 1358442000, 1358445600, 1358449200, 1358452800, 
    1358456400, 1358460000, 1358463600, 1358467200, 1358470800, 1358474400, 
    1358478000, 1358481600, 1358485200, 1358488800, 1358492400, 1358496000, 
    1358499600, 1358503200, 1358506800, 1358510400, 1358514000, 1358517600, 
    1358521200, 1358524800, 1358528400, 1358532000, 1358535600, 1358539200, 
    1358542800, 1358546400, 1358550000, 1358553600, 1358557200, 1358560800, 
    1358564400, 1358568000, 1358571600, 1358575200, 1358578800, 1358582400, 
    1358586000, 1358589600, 1358593200, 1358596800, 1358600400, 1358604000, 
    1358607600, 1358611200, 1358614800, 1358618400, 1358622000, 1358625600, 
    1358629200, 1358632800, 1358636400, 1358640000, 1358643600, 1358647200, 
    1358650800, 1358654400, 1358658000, 1358661600, 1358665200, 1358668800, 
    1358672400, 1358676000, 1358679600, 1358683200, 1358686800, 1358690400, 
    1358694000, 1358697600, 1358701200, 1358704800, 1358708400, 1358712000, 
    1358715600, 1358719200, 1358722800, 1358726400, 1358730000, 1358733600, 
    1358737200, 1358740800, 1358744400, 1358748000, 1358751600, 1358755200, 
    1358758800, 1358762400, 1358766000, 1358769600, 1358773200, 1358776800, 
    1358780400, 1358784000, 1358787600, 1358791200, 1358794800, 1358798400, 
    1358802000, 1358805600, 1358809200, 1358812800, 1358816400, 1358820000, 
    1358823600, 1358827200, 1358830800, 1358834400, 1358838000, 1358841600, 
    1358845200, 1358848800, 1358852400, 1358856000, 1358859600, 1358863200, 
    1358866800, 1358870400, 1358874000, 1358877600, 1358881200, 1358884800, 
    1358888400, 1358892000, 1358895600, 1358899200, 1358902800, 1358906400, 
    1358910000, 1358913600, 1358917200, 1358920800, 1358924400, 1358928000, 
    1358931600, 1358935200, 1358938800, 1358942400, 1358946000, 1358949600, 
    1358953200, 1358956800, 1358960400, 1358964000, 1358967600, 1358971200, 
    1358974800, 1358978400, 1358982000, 1358985600, 1358989200, 1358992800, 
    1358996400, 1359000000, 1359003600, 1359007200, 1359010800, 1359014400, 
    1359018000, 1359021600, 1359025200, 1359028800, 1359032400, 1359036000, 
    1359039600, 1359043200, 1359046800, 1359050400, 1359054000, 1359057600, 
    1359061200, 1359064800, 1359068400, 1359072000, 1359075600, 1359079200, 
    1359082800, 1359086400, 1359090000, 1359093600, 1359097200, 1359100800, 
    1359104400, 1359108000, 1359111600, 1359115200, 1359118800, 1359122400, 
    1359126000, 1359129600, 1359133200, 1359136800, 1359140400, 1359144000, 
    1359147600, 1359151200, 1359154800, 1359158400, 1359162000, 1359165600, 
    1359169200, 1359172800, 1359176400, 1359180000, 1359183600, 1359187200, 
    1359190800, 1359194400, 1359198000, 1359201600, 1359205200, 1359208800, 
    1359212400, 1359216000, 1359219600, 1359223200, 1359226800, 1359230400, 
    1359234000, 1359237600, 1359241200, 1359244800, 1359248400, 1359252000, 
    1359255600, 1359259200, 1359262800, 1359266400, 1359270000, 1359273600, 
    1359277200, 1359280800, 1359284400, 1359288000, 1359291600, 1359295200, 
    1359298800, 1359302400, 1359306000, 1359309600, 1359313200, 1359316800, 
    1359320400, 1359324000, 1359327600, 1359331200, 1359334800, 1359338400, 
    1359342000, 1359345600, 1359349200, 1359352800, 1359356400, 1359360000, 
    1359363600, 1359367200, 1359370800, 1359374400, 1359378000, 1359381600, 
    1359385200, 1359388800, 1359392400, 1359396000, 1359399600, 1359403200, 
    1359406800, 1359410400, 1359414000, 1359417600, 1359421200, 1359424800, 
    1359428400, 1359432000, 1359435600, 1359439200, 1359442800, 1359446400, 
    1359450000, 1359453600, 1359457200, 1359460800, 1359464400, 1359468000, 
    1359471600, 1359475200, 1359478800, 1359482400, 1359486000, 1359489600, 
    1359493200, 1359496800, 1359500400, 1359504000, 1359507600, 1359511200, 
    1359514800, 1359518400, 1359522000, 1359525600, 1359529200, 1359532800, 
    1359536400, 1359540000, 1359543600, 1359547200, 1359550800, 1359554400, 
    1359558000, 1359561600, 1359565200, 1359568800, 1359572400, 1359576000, 
    1359579600, 1359583200, 1359586800, 1359590400, 1359594000, 1359597600, 
    1359601200, 1359604800, 1359608400, 1359612000, 1359615600, 1359619200, 
    1359622800, 1359626400, 1359630000, 1359633600, 1359637200, 1359640800, 
    1359644400, 1359648000, 1359651600, 1359655200, 1359658800, 1359662400, 
    1359666000, 1359669600, 1359673200, 1359676800, 1359680400, 1359684000, 
    1359687600, 1359691200, 1359694800, 1359698400, 1359702000, 1359705600, 
    1359709200, 1359712800, 1359716400, 1359720000, 1359723600, 1359727200, 
    1359730800, 1359734400, 1359738000, 1359741600, 1359745200, 1359748800, 
    1359752400, 1359756000, 1359759600, 1359763200, 1359766800, 1359770400, 
    1359774000, 1359777600, 1359781200, 1359784800, 1359788400, 1359792000, 
    1359795600, 1359799200, 1359802800, 1359806400, 1359810000, 1359813600, 
    1359817200, 1359820800, 1359824400, 1359828000, 1359831600, 1359835200, 
    1359838800, 1359842400, 1359846000, 1359849600, 1359853200, 1359856800, 
    1359860400, 1359864000, 1359867600, 1359871200, 1359874800, 1359878400, 
    1359882000, 1359885600, 1359889200, 1359892800, 1359896400, 1359900000, 
    1359903600, 1359907200, 1359910800, 1359914400, 1359918000, 1359921600, 
    1359925200, 1359928800, 1359932400, 1359936000, 1359939600, 1359943200, 
    1359946800, 1359950400, 1359954000, 1359957600, 1359961200, 1359964800, 
    1359968400, 1359972000, 1359975600, 1359979200, 1359982800, 1359986400, 
    1359990000, 1359993600, 1359997200, 1360000800, 1360004400, 1360008000, 
    1360011600, 1360015200, 1360018800, 1360022400, 1360026000, 1360029600, 
    1360033200, 1360036800, 1360040400, 1360044000, 1360047600, 1360051200, 
    1360054800, 1360058400, 1360062000, 1360065600, 1360069200, 1360072800, 
    1360076400, 1360080000, 1360083600, 1360087200, 1360090800, 1360094400, 
    1360098000, 1360101600, 1360105200, 1360108800, 1360112400, 1360116000, 
    1360119600, 1360123200, 1360126800, 1360130400, 1360134000, 1360137600, 
    1360141200, 1360144800, 1360148400, 1360152000, 1360155600, 1360159200, 
    1360162800, 1360166400, 1360170000, 1360173600, 1360177200, 1360180800, 
    1360184400, 1360188000, 1360191600, 1360195200, 1360198800, 1360202400, 
    1360206000, 1360209600, 1360213200, 1360216800, 1360220400, 1360224000, 
    1360227600, 1360231200, 1360234800, 1360238400, 1360242000, 1360245600, 
    1360249200, 1360252800, 1360256400, 1360260000, 1360263600, 1360267200, 
    1360270800, 1360274400, 1360278000, 1360281600, 1360285200, 1360288800, 
    1360292400, 1360296000, 1360299600, 1360303200, 1360306800, 1360310400, 
    1360314000, 1360317600, 1360321200, 1360324800, 1360328400, 1360332000, 
    1360335600, 1360339200, 1360342800, 1360346400, 1360350000, 1360353600, 
    1360357200, 1360360800, 1360364400, 1360368000, 1360371600, 1360375200, 
    1360378800, 1360382400, 1360386000, 1360389600, 1360393200, 1360396800, 
    1360400400, 1360404000, 1360407600, 1360411200, 1360414800, 1360418400, 
    1360422000, 1360425600, 1360429200, 1360432800, 1360436400, 1360440000, 
    1360443600, 1360447200, 1360450800, 1360454400, 1360458000, 1360461600, 
    1360465200, 1360468800, 1360472400, 1360476000, 1360479600, 1360483200, 
    1360486800, 1360490400, 1360494000, 1360497600, 1360501200, 1360504800, 
    1360508400, 1360512000, 1360515600, 1360519200, 1360522800, 1360526400, 
    1360530000, 1360533600, 1360537200, 1360540800, 1360544400, 1360548000, 
    1360551600, 1360555200, 1360558800, 1360562400, 1360566000, 1360569600, 
    1360573200, 1360576800, 1360580400, 1360584000, 1360587600, 1360591200, 
    1360594800, 1360598400, 1360602000, 1360605600, 1360609200, 1360612800, 
    1360616400, 1360620000, 1360623600, 1360627200, 1360630800, 1360634400, 
    1360638000, 1360641600, 1360645200, 1360648800, 1360652400, 1360656000, 
    1360659600, 1360663200, 1360666800, 1360670400, 1360674000, 1360677600, 
    1360681200, 1360684800, 1360688400, 1360692000, 1360695600, 1360699200, 
    1360702800, 1360706400, 1360710000, 1360713600, 1360717200, 1360720800, 
    1360724400, 1360728000, 1360731600, 1360735200, 1360738800, 1360742400, 
    1360746000, 1360749600, 1360753200, 1360756800, 1360760400, 1360764000, 
    1360767600, 1360771200, 1360774800, 1360778400, 1360782000, 1360785600, 
    1360789200, 1360792800, 1360796400, 1360800000, 1360803600, 1360807200, 
    1360810800, 1360814400, 1360818000, 1360821600, 1360825200, 1360828800, 
    1360832400, 1360836000, 1360839600, 1360843200, 1360846800, 1360850400, 
    1360854000, 1360857600, 1360861200, 1360864800, 1360868400, 1360872000, 
    1360875600, 1360879200, 1360882800, 1360886400, 1360890000, 1360893600, 
    1360897200, 1360900800, 1360904400, 1360908000, 1360911600, 1360915200, 
    1360918800, 1360922400, 1360926000, 1360929600, 1360933200, 1360936800, 
    1360940400, 1360944000, 1360947600, 1360951200, 1360954800, 1360958400, 
    1360962000, 1360965600, 1360969200, 1360972800, 1360976400, 1360980000, 
    1360983600, 1360987200, 1360990800, 1360994400, 1360998000, 1361001600, 
    1361005200, 1361008800, 1361012400, 1361016000, 1361019600, 1361023200, 
    1361026800, 1361030400, 1361034000, 1361037600, 1361041200, 1361044800, 
    1361048400, 1361052000, 1361055600, 1361059200, 1361062800, 1361066400, 
    1361070000, 1361073600, 1361077200, 1361080800, 1361084400, 1361088000, 
    1361091600, 1361095200, 1361098800, 1361102400, 1361106000, 1361109600, 
    1361113200, 1361116800, 1361120400, 1361124000, 1361127600, 1361131200, 
    1361134800, 1361138400, 1361142000, 1361145600, 1361149200, 1361152800, 
    1361156400, 1361160000, 1361163600, 1361167200, 1361170800, 1361174400, 
    1361178000, 1361181600, 1361185200, 1361188800, 1361192400, 1361196000, 
    1361199600, 1361203200, 1361206800, 1361210400, 1361214000, 1361217600, 
    1361221200, 1361224800, 1361228400, 1361232000, 1361235600, 1361239200, 
    1361242800, 1361246400, 1361250000, 1361253600, 1361257200, 1361260800, 
    1361264400, 1361268000, 1361271600, 1361275200, 1361278800, 1361282400, 
    1361286000, 1361289600, 1361293200, 1361296800, 1361300400, 1361304000, 
    1361307600, 1361311200, 1361314800, 1361318400, 1361322000, 1361325600, 
    1361329200, 1361332800, 1361336400, 1361340000, 1361343600, 1361347200, 
    1361350800, 1361354400, 1361358000, 1361361600, 1361365200, 1361368800, 
    1361372400, 1361376000, 1361379600, 1361383200, 1361386800, 1361390400, 
    1361394000, 1361397600, 1361401200, 1361404800, 1361408400, 1361412000, 
    1361415600, 1361419200, 1361422800, 1361426400, 1361430000, 1361433600, 
    1361437200, 1361440800, 1361444400, 1361448000, 1361451600, 1361455200, 
    1361458800, 1361462400, 1361466000, 1361469600, 1361473200, 1361476800, 
    1361480400, 1361484000, 1361487600, 1361491200, 1361494800, 1361498400, 
    1361502000, 1361505600, 1361509200, 1361512800, 1361516400, 1361520000, 
    1361523600, 1361527200, 1361530800, 1361534400, 1361538000, 1361541600, 
    1361545200, 1361548800, 1361552400, 1361556000, 1361559600, 1361563200, 
    1361566800, 1361570400, 1361574000, 1361577600, 1361581200, 1361584800, 
    1361588400, 1361592000, 1361595600, 1361599200, 1361602800, 1361606400, 
    1361610000, 1361613600, 1361617200, 1361620800, 1361624400, 1361628000, 
    1361631600, 1361635200, 1361638800, 1361642400, 1361646000, 1361649600, 
    1361653200, 1361656800, 1361660400, 1361664000, 1361667600, 1361671200, 
    1361674800, 1361678400, 1361682000, 1361685600, 1361689200, 1361692800, 
    1361696400, 1361700000, 1361703600, 1361707200, 1361710800, 1361714400, 
    1361718000, 1361721600, 1361725200, 1361728800, 1361732400, 1361736000, 
    1361739600, 1361743200, 1361746800, 1361750400, 1361754000, 1361757600, 
    1361761200, 1361764800, 1361768400, 1361772000, 1361775600, 1361779200, 
    1361782800, 1361786400, 1361790000, 1361793600, 1361797200, 1361800800, 
    1361804400, 1361808000, 1361811600, 1361815200, 1361818800, 1361822400, 
    1361826000, 1361829600, 1361833200, 1361836800, 1361840400, 1361844000, 
    1361847600, 1361851200, 1361854800, 1361858400, 1361862000, 1361865600, 
    1361869200, 1361872800, 1361876400, 1361880000, 1361883600, 1361887200, 
    1361890800, 1361894400, 1361898000, 1361901600, 1361905200, 1361908800, 
    1361912400, 1361916000, 1361919600, 1361923200, 1361926800, 1361930400, 
    1361934000, 1361937600, 1361941200, 1361944800, 1361948400, 1361952000, 
    1361955600, 1361959200, 1361962800, 1361966400, 1361970000, 1361973600, 
    1361977200, 1361980800, 1361984400, 1361988000, 1361991600, 1361995200, 
    1361998800, 1362002400, 1362006000, 1362009600, 1362013200, 1362016800, 
    1362020400, 1362024000, 1362027600, 1362031200, 1362034800, 1362038400, 
    1362042000, 1362045600, 1362049200, 1362052800, 1362056400, 1362060000, 
    1362063600, 1362067200, 1362070800, 1362074400, 1362078000, 1362081600, 
    1362085200, 1362088800, 1362092400, 1362096000, 1362099600, 1362103200, 
    1362106800, 1362110400, 1362114000, 1362117600, 1362121200, 1362124800, 
    1362128400, 1362132000, 1362135600, 1362139200, 1362142800, 1362146400, 
    1362150000, 1362153600, 1362157200, 1362160800, 1362164400, 1362168000, 
    1362171600, 1362175200, 1362178800, 1362182400, 1362186000, 1362189600, 
    1362193200, 1362196800, 1362200400, 1362204000, 1362207600, 1362211200, 
    1362214800, 1362218400, 1362222000, 1362225600, 1362229200, 1362232800, 
    1362236400, 1362240000, 1362243600, 1362247200, 1362250800, 1362254400, 
    1362258000, 1362261600, 1362265200, 1362268800, 1362272400, 1362276000, 
    1362279600, 1362283200, 1362286800, 1362290400, 1362294000, 1362297600, 
    1362301200, 1362304800, 1362308400, 1362312000, 1362315600, 1362319200, 
    1362322800, 1362326400, 1362330000, 1362333600, 1362337200, 1362340800, 
    1362344400, 1362348000, 1362351600, 1362355200, 1362358800, 1362362400, 
    1362366000, 1362369600, 1362373200, 1362376800, 1362380400, 1362384000, 
    1362387600, 1362391200, 1362394800, 1362398400, 1362402000, 1362405600, 
    1362409200, 1362412800, 1362416400, 1362420000, 1362423600, 1362427200, 
    1362430800, 1362434400, 1362438000, 1362441600, 1362445200, 1362448800, 
    1362452400, 1362456000, 1362459600, 1362463200, 1362466800, 1362470400, 
    1362474000, 1362477600, 1362481200, 1362484800, 1362488400, 1362492000, 
    1362495600, 1362499200, 1362502800, 1362506400, 1362510000, 1362513600, 
    1362517200, 1362520800, 1362524400, 1362528000, 1362531600, 1362535200, 
    1362538800, 1362542400, 1362546000, 1362549600, 1362553200, 1362556800, 
    1362560400, 1362564000, 1362567600, 1362571200, 1362574800, 1362578400, 
    1362582000, 1362585600, 1362589200, 1362592800, 1362596400, 1362600000, 
    1362603600, 1362607200, 1362610800, 1362614400, 1362618000, 1362621600, 
    1362625200, 1362628800, 1362632400, 1362636000, 1362639600, 1362643200, 
    1362646800, 1362650400, 1362654000, 1362657600, 1362661200, 1362664800, 
    1362668400, 1362672000, 1362675600, 1362679200, 1362682800, 1362686400, 
    1362690000, 1362693600, 1362697200, 1362700800, 1362704400, 1362708000, 
    1362711600, 1362715200, 1362718800, 1362722400, 1362726000, 1362729600, 
    1362733200, 1362736800, 1362740400, 1362744000, 1362747600, 1362751200, 
    1362754800, 1362758400, 1362762000, 1362765600, 1362769200, 1362772800, 
    1362776400, 1362780000, 1362783600, 1362787200, 1362790800, 1362794400, 
    1362798000, 1362801600, 1362805200, 1362808800, 1362812400, 1362816000, 
    1362819600, 1362823200, 1362826800, 1362830400, 1362834000, 1362837600, 
    1362841200, 1362844800, 1362848400, 1362852000, 1362855600, 1362859200, 
    1362862800, 1362866400, 1362870000, 1362873600, 1362877200, 1362880800, 
    1362884400, 1362888000, 1362891600, 1362895200, 1362898800, 1362902400, 
    1362906000, 1362909600, 1362913200, 1362916800, 1362920400, 1362924000, 
    1362927600, 1362931200, 1362934800, 1362938400, 1362942000, 1362945600, 
    1362949200, 1362952800, 1362956400, 1362960000, 1362963600, 1362967200, 
    1362970800, 1362974400, 1362978000, 1362981600, 1362985200, 1362988800, 
    1362992400, 1362996000, 1362999600, 1363003200, 1363006800, 1363010400, 
    1363014000, 1363017600, 1363021200, 1363024800, 1363028400, 1363032000, 
    1363035600, 1363039200, 1363042800, 1363046400, 1363050000, 1363053600, 
    1363057200, 1363060800, 1363064400, 1363068000, 1363071600, 1363075200, 
    1363078800, 1363082400, 1363086000, 1363089600, 1363093200, 1363096800, 
    1363100400, 1363104000, 1363107600, 1363111200, 1363114800, 1363118400, 
    1363122000, 1363125600, 1363129200, 1363132800, 1363136400, 1363140000, 
    1363143600, 1363147200, 1363150800, 1363154400, 1363158000, 1363161600, 
    1363165200, 1363168800, 1363172400, 1363176000, 1363179600, 1363183200, 
    1363186800, 1363190400, 1363194000, 1363197600, 1363201200, 1363204800, 
    1363208400, 1363212000, 1363215600, 1363219200, 1363222800, 1363226400, 
    1363230000, 1363233600, 1363237200, 1363240800, 1363244400, 1363248000, 
    1363251600, 1363255200, 1363258800, 1363262400, 1363266000, 1363269600, 
    1363273200, 1363276800, 1363280400, 1363284000, 1363287600, 1363291200, 
    1363294800, 1363298400, 1363302000, 1363305600, 1363309200, 1363312800, 
    1363316400, 1363320000, 1363323600, 1363327200, 1363330800, 1363334400, 
    1363338000, 1363341600, 1363345200, 1363348800, 1363352400, 1363356000, 
    1363359600, 1363363200, 1363366800, 1363370400, 1363374000, 1363377600, 
    1363381200, 1363384800, 1363388400, 1363392000, 1363395600, 1363399200, 
    1363402800, 1363406400, 1363410000, 1363413600, 1363417200, 1363420800, 
    1363424400, 1363428000, 1363431600, 1363435200, 1363438800, 1363442400, 
    1363446000, 1363449600, 1363453200, 1363456800, 1363460400, 1363464000, 
    1363467600, 1363471200, 1363474800, 1363478400, 1363482000, 1363485600, 
    1363489200, 1363492800, 1363496400, 1363500000, 1363503600, 1363507200, 
    1363510800, 1363514400, 1363518000, 1363521600, 1363525200, 1363528800, 
    1363532400, 1363536000, 1363539600, 1363543200, 1363546800, 1363550400, 
    1363554000, 1363557600, 1363561200, 1363564800, 1363568400, 1363572000, 
    1363575600, 1363579200, 1363582800, 1363586400, 1363590000, 1363593600, 
    1363597200, 1363600800, 1363604400, 1363608000, 1363611600, 1363615200, 
    1363618800, 1363622400, 1363626000, 1363629600, 1363633200, 1363636800, 
    1363640400, 1363644000, 1363647600, 1363651200, 1363654800, 1363658400, 
    1363662000, 1363665600, 1363669200, 1363672800, 1363676400, 1363680000, 
    1363683600, 1363687200, 1363690800, 1363694400, 1363698000, 1363701600, 
    1363705200, 1363708800, 1363712400, 1363716000, 1363719600, 1363723200, 
    1363726800, 1363730400, 1363734000, 1363737600, 1363741200, 1363744800, 
    1363748400, 1363752000, 1363755600, 1363759200, 1363762800, 1363766400, 
    1363770000, 1363773600, 1363777200, 1363780800, 1363784400, 1363788000, 
    1363791600, 1363795200, 1363798800, 1363802400, 1363806000, 1363809600, 
    1363813200, 1363816800, 1363820400, 1363824000, 1363827600, 1363831200, 
    1363834800, 1363838400, 1363842000, 1363845600, 1363849200, 1363852800, 
    1363856400, 1363860000, 1363863600, 1363867200, 1363870800, 1363874400, 
    1363878000, 1363881600, 1363885200, 1363888800, 1363892400, 1363896000, 
    1363899600, 1363903200, 1363906800, 1363910400, 1363914000, 1363917600, 
    1363921200, 1363924800, 1363928400, 1363932000, 1363935600, 1363939200, 
    1363942800, 1363946400, 1363950000, 1363953600, 1363957200, 1363960800, 
    1363964400, 1363968000, 1363971600, 1363975200, 1363978800, 1363982400, 
    1363986000, 1363989600, 1363993200, 1363996800, 1364000400, 1364004000, 
    1364007600, 1364011200, 1364014800, 1364018400, 1364022000, 1364025600, 
    1364029200, 1364032800, 1364036400, 1364040000, 1364043600, 1364047200, 
    1364050800, 1364054400, 1364058000, 1364061600, 1364065200, 1364068800, 
    1364072400, 1364076000, 1364079600, 1364083200, 1364086800, 1364090400, 
    1364094000, 1364097600, 1364101200, 1364104800, 1364108400, 1364112000, 
    1364115600, 1364119200, 1364122800, 1364126400, 1364130000, 1364133600, 
    1364137200, 1364140800, 1364144400, 1364148000, 1364151600, 1364155200, 
    1364158800, 1364162400, 1364166000, 1364169600, 1364173200, 1364176800, 
    1364180400, 1364184000, 1364187600, 1364191200, 1364194800, 1364198400, 
    1364202000, 1364205600, 1364209200, 1364212800, 1364216400, 1364220000, 
    1364223600, 1364227200, 1364230800, 1364234400, 1364238000, 1364241600, 
    1364245200, 1364248800, 1364252400, 1364256000, 1364259600, 1364263200, 
    1364266800, 1364270400, 1364274000, 1364277600, 1364281200, 1364284800, 
    1364288400, 1364292000, 1364295600, 1364299200, 1364302800, 1364306400, 
    1364310000, 1364313600, 1364317200, 1364320800, 1364324400, 1364328000, 
    1364331600, 1364335200, 1364338800, 1364342400, 1364346000, 1364349600, 
    1364353200, 1364356800, 1364360400, 1364364000, 1364367600, 1364371200, 
    1364374800, 1364378400, 1364382000, 1364385600, 1364389200, 1364392800, 
    1364396400, 1364400000, 1364403600, 1364407200, 1364410800, 1364414400, 
    1364418000, 1364421600, 1364425200, 1364428800, 1364432400, 1364436000, 
    1364439600, 1364443200, 1364446800, 1364450400, 1364454000, 1364457600, 
    1364461200, 1364464800, 1364468400, 1364472000, 1364475600, 1364479200, 
    1364482800, 1364486400, 1364490000, 1364493600, 1364497200, 1364500800, 
    1364504400, 1364508000, 1364511600, 1364515200, 1364518800, 1364522400, 
    1364526000, 1364529600, 1364533200, 1364536800, 1364540400, 1364544000, 
    1364547600, 1364551200, 1364554800, 1364558400, 1364562000, 1364565600, 
    1364569200, 1364572800, 1364576400, 1364580000, 1364583600, 1364587200, 
    1364590800, 1364594400, 1364598000, 1364601600, 1364605200, 1364608800, 
    1364612400, 1364616000, 1364619600, 1364623200, 1364626800, 1364630400, 
    1364634000, 1364637600, 1364641200, 1364644800, 1364648400, 1364652000, 
    1364655600, 1364659200, 1364662800, 1364666400, 1364670000, 1364673600, 
    1364677200, 1364680800, 1364684400, 1364688000, 1364691600, 1364695200, 
    1364698800, 1364702400, 1364706000, 1364709600, 1364713200, 1364716800, 
    1364720400, 1364724000, 1364727600, 1364731200, 1364734800, 1364738400, 
    1364742000, 1364745600, 1364749200, 1364752800, 1364756400, 1364760000, 
    1364763600, 1364767200, 1364770800, 1364774400, 1364778000, 1364781600, 
    1364785200, 1364788800, 1364792400, 1364796000, 1364799600, 1364803200, 
    1364806800, 1364810400, 1364814000, 1364817600, 1364821200, 1364824800, 
    1364828400, 1364832000, 1364835600, 1364839200, 1364842800, 1364846400, 
    1364850000, 1364853600, 1364857200, 1364860800, 1364864400, 1364868000, 
    1364871600, 1364875200, 1364878800, 1364882400, 1364886000, 1364889600, 
    1364893200, 1364896800, 1364900400, 1364904000, 1364907600, 1364911200, 
    1364914800, 1364918400, 1364922000, 1364925600, 1364929200, 1364932800, 
    1364936400, 1364940000, 1364943600, 1364947200, 1364950800, 1364954400, 
    1364958000, 1364961600, 1364965200, 1364968800, 1364972400, 1364976000, 
    1364979600, 1364983200, 1364986800, 1364990400, 1364994000, 1364997600, 
    1365001200, 1365004800, 1365008400, 1365012000, 1365015600, 1365019200, 
    1365022800, 1365026400, 1365030000, 1365033600, 1365037200, 1365040800, 
    1365044400, 1365048000, 1365051600, 1365055200, 1365058800, 1365062400, 
    1365066000, 1365069600, 1365073200, 1365076800, 1365080400, 1365084000, 
    1365087600, 1365091200, 1365094800, 1365098400, 1365102000, 1365105600, 
    1365109200, 1365112800, 1365116400, 1365120000, 1365123600, 1365127200, 
    1365130800, 1365134400, 1365138000, 1365141600, 1365145200, 1365148800, 
    1365152400, 1365156000, 1365159600, 1365163200, 1365166800, 1365170400, 
    1365174000, 1365177600, 1365181200, 1365184800, 1365188400, 1365192000, 
    1365195600, 1365199200, 1365202800, 1365206400, 1365210000, 1365213600, 
    1365217200, 1365220800, 1365224400, 1365228000, 1365231600, 1365235200, 
    1365238800, 1365242400, 1365246000, 1365249600, 1365253200, 1365256800, 
    1365260400, 1365264000, 1365267600, 1365271200, 1365274800, 1365278400, 
    1365282000, 1365285600, 1365289200, 1365292800, 1365296400, 1365300000, 
    1365303600, 1365307200, 1365310800, 1365314400, 1365318000, 1365321600, 
    1365325200, 1365328800, 1365332400, 1365336000, 1365339600, 1365343200, 
    1365346800, 1365350400, 1365354000, 1365357600, 1365361200, 1365364800, 
    1365368400, 1365372000, 1365375600, 1365379200, 1365382800, 1365386400, 
    1365390000, 1365393600, 1365397200, 1365400800, 1365404400, 1365408000, 
    1365411600, 1365415200, 1365418800, 1365422400, 1365426000, 1365429600, 
    1365433200, 1365436800, 1365440400, 1365444000, 1365447600, 1365451200, 
    1365454800, 1365458400, 1365462000, 1365465600, 1365469200, 1365472800, 
    1365476400, 1365480000, 1365483600, 1365487200, 1365490800, 1365494400, 
    1365498000, 1365501600, 1365505200, 1365508800, 1365512400, 1365516000, 
    1365519600, 1365523200, 1365526800, 1365530400, 1365534000, 1365537600, 
    1365541200, 1365544800, 1365548400, 1365552000, 1365555600, 1365559200, 
    1365562800, 1365566400, 1365570000, 1365573600, 1365577200, 1365580800, 
    1365584400, 1365588000, 1365591600, 1365595200, 1365598800, 1365602400, 
    1365606000, 1365609600, 1365613200, 1365616800, 1365620400, 1365624000, 
    1365627600, 1365631200, 1365634800, 1365638400, 1365642000, 1365645600, 
    1365649200, 1365652800, 1365656400, 1365660000, 1365663600, 1365667200, 
    1365670800, 1365674400, 1365678000, 1365681600, 1365685200, 1365688800, 
    1365692400, 1365696000, 1365699600, 1365703200, 1365706800, 1365710400, 
    1365714000, 1365717600, 1365721200, 1365724800, 1365728400, 1365732000, 
    1365735600, 1365739200, 1365742800, 1365746400, 1365750000, 1365753600, 
    1365757200, 1365760800, 1365764400, 1365768000, 1365771600, 1365775200, 
    1365778800, 1365782400, 1365786000, 1365789600, 1365793200, 1365796800, 
    1365800400, 1365804000, 1365807600, 1365811200, 1365814800, 1365818400, 
    1365822000, 1365825600, 1365829200, 1365832800, 1365836400, 1365840000, 
    1365843600, 1365847200, 1365850800, 1365854400, 1365858000, 1365861600, 
    1365865200, 1365868800, 1365872400, 1365876000, 1365879600, 1365883200, 
    1365886800, 1365890400, 1365894000, 1365897600, 1365901200, 1365904800, 
    1365908400, 1365912000, 1365915600, 1365919200, 1365922800, 1365926400, 
    1365930000, 1365933600, 1365937200, 1365940800, 1365944400, 1365948000, 
    1365951600, 1365955200, 1365958800, 1365962400, 1365966000, 1365969600, 
    1365973200, 1365976800, 1365980400, 1365984000, 1365987600, 1365991200, 
    1365994800, 1365998400, 1366002000, 1366005600, 1366009200, 1366012800, 
    1366016400, 1366020000, 1366023600, 1366027200, 1366030800, 1366034400, 
    1366038000, 1366041600, 1366045200, 1366048800, 1366052400, 1366056000, 
    1366059600, 1366063200, 1366066800, 1366070400, 1366074000, 1366077600, 
    1366081200, 1366084800, 1366088400, 1366092000, 1366095600, 1366099200, 
    1366102800, 1366106400, 1366110000, 1366113600, 1366117200, 1366120800, 
    1366124400, 1366128000, 1366131600, 1366135200, 1366138800, 1366142400, 
    1366146000, 1366149600, 1366153200, 1366156800, 1366160400, 1366164000, 
    1366167600, 1366171200, 1366174800, 1366178400, 1366182000, 1366185600, 
    1366189200, 1366192800, 1366196400, 1366200000, 1366203600, 1366207200, 
    1366210800, 1366214400, 1366218000, 1366221600, 1366225200, 1366228800, 
    1366232400, 1366236000, 1366239600, 1366243200, 1366246800, 1366250400, 
    1366254000, 1366257600, 1366261200, 1366264800, 1366268400, 1366272000, 
    1366275600, 1366279200, 1366282800, 1366286400, 1366290000, 1366293600, 
    1366297200, 1366300800, 1366304400, 1366308000, 1366311600, 1366315200, 
    1366318800, 1366322400, 1366326000, 1366329600, 1366333200, 1366336800, 
    1366340400, 1366344000, 1366347600, 1366351200, 1366354800, 1366358400, 
    1366362000, 1366365600, 1366369200, 1366372800, 1366376400, 1366380000, 
    1366383600, 1366387200, 1366390800, 1366394400, 1366398000, 1366401600, 
    1366405200, 1366408800, 1366412400, 1366416000, 1366419600, 1366423200, 
    1366426800, 1366430400, 1366434000, 1366437600, 1366441200, 1366444800, 
    1366448400, 1366452000, 1366455600, 1366459200, 1366462800, 1366466400, 
    1366470000, 1366473600, 1366477200, 1366480800, 1366484400, 1366488000, 
    1366491600, 1366495200, 1366498800, 1366502400, 1366506000, 1366509600, 
    1366513200, 1366516800, 1366520400, 1366524000, 1366527600, 1366531200, 
    1366534800, 1366538400, 1366542000, 1366545600, 1366549200, 1366552800, 
    1366556400, 1366560000, 1366563600, 1366567200, 1366570800, 1366574400, 
    1366578000, 1366581600, 1366585200, 1366588800, 1366592400, 1366596000, 
    1366599600, 1366603200, 1366606800, 1366610400, 1366614000, 1366617600, 
    1366621200, 1366624800, 1366628400, 1366632000, 1366635600, 1366639200, 
    1366642800, 1366646400, 1366650000, 1366653600, 1366657200, 1366660800, 
    1366664400, 1366668000, 1366671600, 1366675200, 1366678800, 1366682400, 
    1366686000, 1366689600, 1366693200, 1366696800, 1366700400, 1366704000, 
    1366707600, 1366711200, 1366714800, 1366718400, 1366722000, 1366725600, 
    1366729200, 1366732800, 1366736400, 1366740000, 1366743600, 1366747200, 
    1366750800, 1366754400, 1366758000, 1366761600, 1366765200, 1366768800, 
    1366772400, 1366776000, 1366779600, 1366783200, 1366786800, 1366790400, 
    1366794000, 1366797600, 1366801200, 1366804800, 1366808400, 1366812000, 
    1366815600, 1366819200, 1366822800, 1366826400, 1366830000, 1366833600, 
    1366837200, 1366840800, 1366844400, 1366848000, 1366851600, 1366855200, 
    1366858800, 1366862400, 1366866000, 1366869600, 1366873200, 1366876800, 
    1366880400, 1366884000, 1366887600, 1366891200, 1366894800, 1366898400, 
    1366902000, 1366905600, 1366909200, 1366912800, 1366916400, 1366920000, 
    1366923600, 1366927200, 1366930800, 1366934400, 1366938000, 1366941600, 
    1366945200, 1366948800, 1366952400, 1366956000, 1366959600, 1366963200, 
    1366966800, 1366970400, 1366974000, 1366977600, 1366981200, 1366984800, 
    1366988400, 1366992000, 1366995600, 1366999200, 1367002800, 1367006400, 
    1367010000, 1367013600, 1367017200, 1367020800, 1367024400, 1367028000, 
    1367031600, 1367035200, 1367038800, 1367042400, 1367046000, 1367049600, 
    1367053200, 1367056800, 1367060400, 1367064000, 1367067600, 1367071200, 
    1367074800, 1367078400, 1367082000, 1367085600, 1367089200, 1367092800, 
    1367096400, 1367100000, 1367103600, 1367107200, 1367110800, 1367114400, 
    1367118000, 1367121600, 1367125200, 1367128800, 1367132400, 1367136000, 
    1367139600, 1367143200, 1367146800, 1367150400, 1367154000, 1367157600, 
    1367161200, 1367164800, 1367168400, 1367172000, 1367175600, 1367179200, 
    1367182800, 1367186400, 1367190000, 1367193600, 1367197200, 1367200800, 
    1367204400, 1367208000, 1367211600, 1367215200, 1367218800, 1367222400, 
    1367226000, 1367229600, 1367233200, 1367236800, 1367240400, 1367244000, 
    1367247600, 1367251200, 1367254800, 1367258400, 1367262000, 1367265600, 
    1367269200, 1367272800, 1367276400, 1367280000, 1367283600, 1367287200, 
    1367290800, 1367294400, 1367298000, 1367301600, 1367305200, 1367308800, 
    1367312400, 1367316000, 1367319600, 1367323200, 1367326800, 1367330400, 
    1367334000, 1367337600, 1367341200, 1367344800, 1367348400, 1367352000, 
    1367355600, 1367359200, 1367362800, 1367366400, 1367370000, 1367373600, 
    1367377200, 1367380800, 1367384400, 1367388000, 1367391600, 1367395200, 
    1367398800, 1367402400, 1367406000, 1367409600, 1367413200, 1367416800, 
    1367420400, 1367424000, 1367427600, 1367431200, 1367434800, 1367438400, 
    1367442000, 1367445600, 1367449200, 1367452800, 1367456400, 1367460000, 
    1367463600, 1367467200, 1367470800, 1367474400, 1367478000, 1367481600, 
    1367485200, 1367488800, 1367492400, 1367496000, 1367499600, 1367503200, 
    1367506800, 1367510400, 1367514000, 1367517600, 1367521200, 1367524800, 
    1367528400, 1367532000, 1367535600, 1367539200, 1367542800, 1367546400, 
    1367550000, 1367553600, 1367557200, 1367560800, 1367564400, 1367568000, 
    1367571600, 1367575200, 1367578800, 1367582400, 1367586000, 1367589600, 
    1367593200, 1367596800, 1367600400, 1367604000, 1367607600, 1367611200, 
    1367614800, 1367618400, 1367622000, 1367625600, 1367629200, 1367632800, 
    1367636400, 1367640000, 1367643600, 1367647200, 1367650800, 1367654400, 
    1367658000, 1367661600, 1367665200, 1367668800, 1367672400, 1367676000, 
    1367679600, 1367683200, 1367686800, 1367690400, 1367694000, 1367697600, 
    1367701200, 1367704800, 1367708400, 1367712000, 1367715600, 1367719200, 
    1367722800, 1367726400, 1367730000, 1367733600, 1367737200, 1367740800, 
    1367744400, 1367748000, 1367751600, 1367755200, 1367758800, 1367762400, 
    1367766000, 1367769600, 1367773200, 1367776800, 1367780400, 1367784000, 
    1367787600, 1367791200, 1367794800, 1367798400, 1367802000, 1367805600, 
    1367809200, 1367812800, 1367816400, 1367820000, 1367823600, 1367827200, 
    1367830800, 1367834400, 1367838000, 1367841600, 1367845200, 1367848800, 
    1367852400, 1367856000, 1367859600, 1367863200, 1367866800, 1367870400, 
    1367874000, 1367877600, 1367881200, 1367884800, 1367888400, 1367892000, 
    1367895600, 1367899200, 1367902800, 1367906400, 1367910000, 1367913600, 
    1367917200, 1367920800, 1367924400, 1367928000, 1367931600, 1367935200, 
    1367938800, 1367942400, 1367946000, 1367949600, 1367953200, 1367956800, 
    1367960400, 1367964000, 1367967600, 1367971200, 1367974800, 1367978400, 
    1367982000, 1367985600, 1367989200, 1367992800, 1367996400, 1368000000, 
    1368003600, 1368007200, 1368010800, 1368014400, 1368018000, 1368021600, 
    1368025200, 1368028800, 1368032400, 1368036000, 1368039600, 1368043200, 
    1368046800, 1368050400, 1368054000, 1368057600, 1368061200, 1368064800, 
    1368068400, 1368072000, 1368075600, 1368079200, 1368082800, 1368086400, 
    1368090000, 1368093600, 1368097200, 1368100800, 1368104400, 1368108000, 
    1368111600, 1368115200, 1368118800, 1368122400, 1368126000, 1368129600, 
    1368133200, 1368136800, 1368140400, 1368144000, 1368147600, 1368151200, 
    1368154800, 1368158400, 1368162000, 1368165600, 1368169200, 1368172800, 
    1368176400, 1368180000, 1368183600, 1368187200, 1368190800, 1368194400, 
    1368198000, 1368201600, 1368205200, 1368208800, 1368212400, 1368216000, 
    1368219600, 1368223200, 1368226800, 1368230400, 1368234000, 1368237600, 
    1368241200, 1368244800, 1368248400, 1368252000, 1368255600, 1368259200, 
    1368262800, 1368266400, 1368270000, 1368273600, 1368277200, 1368280800, 
    1368284400, 1368288000, 1368291600, 1368295200, 1368298800, 1368302400, 
    1368306000, 1368309600, 1368313200, 1368316800, 1368320400, 1368324000, 
    1368327600, 1368331200, 1368334800, 1368338400, 1368342000, 1368345600, 
    1368349200, 1368352800, 1368356400, 1368360000, 1368363600, 1368367200, 
    1368370800, 1368374400, 1368378000, 1368381600, 1368385200, 1368388800, 
    1368392400, 1368396000, 1368399600, 1368403200, 1368406800, 1368410400, 
    1368414000, 1368417600, 1368421200, 1368424800, 1368428400, 1368432000, 
    1368435600, 1368439200, 1368442800, 1368446400, 1368450000, 1368453600, 
    1368457200, 1368460800, 1368464400, 1368468000, 1368471600, 1368475200, 
    1368478800, 1368482400, 1368486000, 1368489600, 1368493200, 1368496800, 
    1368500400, 1368504000, 1368507600, 1368511200, 1368514800, 1368518400, 
    1368522000, 1368525600, 1368529200, 1368532800, 1368536400, 1368540000, 
    1368543600, 1368547200, 1368550800, 1368554400, 1368558000, 1368561600, 
    1368565200, 1368568800, 1368572400, 1368576000, 1368579600, 1368583200, 
    1368586800, 1368590400, 1368594000, 1368597600, 1368601200, 1368604800, 
    1368608400, 1368612000, 1368615600, 1368619200, 1368622800, 1368626400, 
    1368630000, 1368633600, 1368637200, 1368640800, 1368644400, 1368648000, 
    1368651600, 1368655200, 1368658800, 1368662400, 1368666000, 1368669600, 
    1368673200, 1368676800, 1368680400, 1368684000, 1368687600, 1368691200, 
    1368694800, 1368698400, 1368702000, 1368705600, 1368709200, 1368712800, 
    1368716400, 1368720000, 1368723600, 1368727200, 1368730800, 1368734400, 
    1368738000, 1368741600, 1368745200, 1368748800, 1368752400, 1368756000, 
    1368759600, 1368763200, 1368766800, 1368770400, 1368774000, 1368777600, 
    1368781200, 1368784800, 1368788400, 1368792000, 1368795600, 1368799200, 
    1368802800, 1368806400, 1368810000, 1368813600, 1368817200, 1368820800, 
    1368824400, 1368828000, 1368831600, 1368835200, 1368838800, 1368842400, 
    1368846000, 1368849600, 1368853200, 1368856800, 1368860400, 1368864000, 
    1368867600, 1368871200, 1368874800, 1368878400, 1368882000, 1368885600, 
    1368889200, 1368892800, 1368896400, 1368900000, 1368903600, 1368907200, 
    1368910800, 1368914400, 1368918000, 1368921600, 1368925200, 1368928800, 
    1368932400, 1368936000, 1368939600, 1368943200, 1368946800, 1368950400, 
    1368954000, 1368957600, 1368961200, 1368964800, 1368968400, 1368972000, 
    1368975600, 1368979200, 1368982800, 1368986400, 1368990000, 1368993600, 
    1368997200, 1369000800, 1369004400, 1369008000, 1369011600, 1369015200, 
    1369018800, 1369022400, 1369026000, 1369029600, 1369033200, 1369036800, 
    1369040400, 1369044000, 1369047600, 1369051200, 1369054800, 1369058400, 
    1369062000, 1369065600, 1369069200, 1369072800, 1369076400, 1369080000, 
    1369083600, 1369087200, 1369090800, 1369094400, 1369098000, 1369101600, 
    1369105200, 1369108800, 1369112400, 1369116000, 1369119600, 1369123200, 
    1369126800, 1369130400, 1369134000, 1369137600, 1369141200, 1369144800, 
    1369148400, 1369152000, 1369155600, 1369159200, 1369162800, 1369166400, 
    1369170000, 1369173600, 1369177200, 1369180800, 1369184400, 1369188000, 
    1369191600, 1369195200, 1369198800, 1369202400, 1369206000, 1369209600, 
    1369213200, 1369216800, 1369220400, 1369224000, 1369227600, 1369231200, 
    1369234800, 1369238400, 1369242000, 1369245600, 1369249200, 1369252800, 
    1369256400, 1369260000, 1369263600, 1369267200, 1369270800, 1369274400, 
    1369278000, 1369281600, 1369285200, 1369288800, 1369292400, 1369296000, 
    1369299600, 1369303200, 1369306800, 1369310400, 1369314000, 1369317600, 
    1369321200, 1369324800, 1369328400, 1369332000, 1369335600, 1369339200, 
    1369342800, 1369346400, 1369350000, 1369353600, 1369357200, 1369360800, 
    1369364400, 1369368000, 1369371600, 1369375200, 1369378800, 1369382400, 
    1369386000, 1369389600, 1369393200, 1369396800, 1369400400, 1369404000, 
    1369407600, 1369411200, 1369414800, 1369418400, 1369422000, 1369425600, 
    1369429200, 1369432800, 1369436400, 1369440000, 1369443600, 1369447200, 
    1369450800, 1369454400, 1369458000, 1369461600, 1369465200, 1369468800, 
    1369472400, 1369476000, 1369479600, 1369483200, 1369486800, 1369490400, 
    1369494000, 1369497600, 1369501200, 1369504800, 1369508400, 1369512000, 
    1369515600, 1369519200, 1369522800, 1369526400, 1369530000, 1369533600, 
    1369537200, 1369540800, 1369544400, 1369548000, 1369551600, 1369555200, 
    1369558800, 1369562400, 1369566000, 1369569600, 1369573200, 1369576800, 
    1369580400, 1369584000, 1369587600, 1369591200, 1369594800, 1369598400, 
    1369602000, 1369605600, 1369609200, 1369612800, 1369616400, 1369620000, 
    1369623600, 1369627200, 1369630800, 1369634400, 1369638000, 1369641600, 
    1369645200, 1369648800, 1369652400, 1369656000, 1369659600, 1369663200, 
    1369666800, 1369670400, 1369674000, 1369677600, 1369681200, 1369684800, 
    1369688400, 1369692000, 1369695600, 1369699200, 1369702800, 1369706400, 
    1369710000, 1369713600, 1369717200, 1369720800, 1369724400, 1369728000, 
    1369731600, 1369735200, 1369738800, 1369742400, 1369746000, 1369749600, 
    1369753200, 1369756800, 1369760400, 1369764000, 1369767600, 1369771200, 
    1369774800, 1369778400, 1369782000, 1369785600, 1369789200, 1369792800, 
    1369796400, 1369800000, 1369803600, 1369807200, 1369810800, 1369814400, 
    1369818000, 1369821600, 1369825200, 1369828800, 1369832400, 1369836000, 
    1369839600, 1369843200, 1369846800, 1369850400, 1369854000, 1369857600, 
    1369861200, 1369864800, 1369868400, 1369872000, 1369875600, 1369879200, 
    1369882800, 1369886400, 1369890000, 1369893600, 1369897200, 1369900800, 
    1369904400, 1369908000, 1369911600, 1369915200, 1369918800, 1369922400, 
    1369926000, 1369929600, 1369933200, 1369936800, 1369940400, 1369944000, 
    1369947600, 1369951200, 1369954800, 1369958400, 1369962000, 1369965600, 
    1369969200, 1369972800, 1369976400, 1369980000, 1369983600, 1369987200, 
    1369990800, 1369994400, 1369998000, 1370001600, 1370005200, 1370008800, 
    1370012400, 1370016000, 1370019600, 1370023200, 1370026800, 1370030400, 
    1370034000, 1370037600, 1370041200, 1370044800, 1370048400, 1370052000, 
    1370055600, 1370059200, 1370062800, 1370066400, 1370070000, 1370073600, 
    1370077200, 1370080800, 1370084400, 1370088000, 1370091600, 1370095200, 
    1370098800, 1370102400, 1370106000, 1370109600, 1370113200, 1370116800, 
    1370120400, 1370124000, 1370127600, 1370131200, 1370134800, 1370138400, 
    1370142000, 1370145600, 1370149200, 1370152800, 1370156400, 1370160000, 
    1370163600, 1370167200, 1370170800, 1370174400, 1370178000, 1370181600, 
    1370185200, 1370188800, 1370192400, 1370196000, 1370199600, 1370203200, 
    1370206800, 1370210400, 1370214000, 1370217600, 1370221200, 1370224800, 
    1370228400, 1370232000, 1370235600, 1370239200, 1370242800, 1370246400, 
    1370250000, 1370253600, 1370257200, 1370260800, 1370264400, 1370268000, 
    1370271600, 1370275200, 1370278800, 1370282400, 1370286000, 1370289600, 
    1370293200, 1370296800, 1370300400, 1370304000, 1370307600, 1370311200, 
    1370314800, 1370318400, 1370322000, 1370325600, 1370329200, 1370332800, 
    1370336400, 1370340000, 1370343600, 1370347200, 1370350800, 1370354400, 
    1370358000, 1370361600, 1370365200, 1370368800, 1370372400, 1370376000, 
    1370379600, 1370383200, 1370386800, 1370390400, 1370394000, 1370397600, 
    1370401200, 1370404800, 1370408400, 1370412000, 1370415600, 1370419200, 
    1370422800, 1370426400, 1370430000, 1370433600, 1370437200, 1370440800, 
    1370444400, 1370448000, 1370451600, 1370455200, 1370458800, 1370462400, 
    1370466000, 1370469600, 1370473200, 1370476800, 1370480400, 1370484000, 
    1370487600, 1370491200, 1370494800, 1370498400, 1370502000, 1370505600, 
    1370509200, 1370512800, 1370516400, 1370520000, 1370523600, 1370527200, 
    1370530800, 1370534400, 1370538000, 1370541600, 1370545200, 1370548800, 
    1370552400, 1370556000, 1370559600, 1370563200, 1370566800, 1370570400, 
    1370574000, 1370577600, 1370581200, 1370584800, 1370588400, 1370592000, 
    1370595600, 1370599200, 1370602800, 1370606400, 1370610000, 1370613600, 
    1370617200, 1370620800, 1370624400, 1370628000, 1370631600, 1370635200, 
    1370638800, 1370642400, 1370646000, 1370649600, 1370653200, 1370656800, 
    1370660400, 1370664000, 1370667600, 1370671200, 1370674800, 1370678400, 
    1370682000, 1370685600, 1370689200, 1370692800, 1370696400, 1370700000, 
    1370703600, 1370707200, 1370710800, 1370714400, 1370718000, 1370721600, 
    1370725200, 1370728800, 1370732400, 1370736000, 1370739600, 1370743200, 
    1370746800, 1370750400, 1370754000, 1370757600, 1370761200, 1370764800, 
    1370768400, 1370772000, 1370775600, 1370779200, 1370782800, 1370786400, 
    1370790000, 1370793600, 1370797200, 1370800800, 1370804400, 1370808000, 
    1370811600, 1370815200, 1370818800, 1370822400, 1370826000, 1370829600, 
    1370833200, 1370836800, 1370840400, 1370844000, 1370847600, 1370851200, 
    1370854800, 1370858400, 1370862000, 1370865600, 1370869200, 1370872800, 
    1370876400, 1370880000, 1370883600, 1370887200, 1370890800, 1370894400, 
    1370898000, 1370901600, 1370905200, 1370908800, 1370912400, 1370916000, 
    1370919600, 1370923200, 1370926800, 1370930400, 1370934000, 1370937600, 
    1370941200, 1370944800, 1370948400, 1370952000, 1370955600, 1370959200, 
    1370962800, 1370966400, 1370970000, 1370973600, 1370977200, 1370980800, 
    1370984400, 1370988000, 1370991600, 1370995200, 1370998800, 1371002400, 
    1371006000, 1371009600, 1371013200, 1371016800, 1371020400, 1371024000, 
    1371027600, 1371031200, 1371034800, 1371038400, 1371042000, 1371045600, 
    1371049200, 1371052800, 1371056400, 1371060000, 1371063600, 1371067200, 
    1371070800, 1371074400, 1371078000, 1371081600, 1371085200, 1371088800, 
    1371092400, 1371096000, 1371099600, 1371103200, 1371106800, 1371110400, 
    1371114000, 1371117600, 1371121200, 1371124800, 1371128400, 1371132000, 
    1371135600, 1371139200, 1371142800, 1371146400, 1371150000, 1371153600, 
    1371157200, 1371160800, 1371164400, 1371168000, 1371171600, 1371175200, 
    1371178800, 1371182400, 1371186000, 1371189600, 1371193200, 1371196800, 
    1371200400, 1371204000, 1371207600, 1371211200, 1371214800, 1371218400, 
    1371222000, 1371225600, 1371229200, 1371232800, 1371236400, 1371240000, 
    1371243600, 1371247200, 1371250800, 1371254400, 1371258000, 1371261600, 
    1371265200, 1371268800, 1371272400, 1371276000, 1371279600, 1371283200, 
    1371286800, 1371290400, 1371294000, 1371297600, 1371301200, 1371304800, 
    1371308400, 1371312000, 1371315600, 1371319200, 1371322800, 1371326400, 
    1371330000, 1371333600, 1371337200, 1371340800, 1371344400, 1371348000, 
    1371351600, 1371355200, 1371358800, 1371362400, 1371366000, 1371369600, 
    1371373200, 1371376800, 1371380400, 1371384000, 1371387600, 1371391200, 
    1371394800, 1371398400, 1371402000, 1371405600, 1371409200, 1371412800, 
    1371416400, 1371420000, 1371423600, 1371427200, 1371430800, 1371434400, 
    1371438000, 1371441600, 1371445200, 1371448800, 1371452400, 1371456000, 
    1371459600, 1371463200, 1371466800, 1371470400, 1371474000, 1371477600, 
    1371481200, 1371484800, 1371488400, 1371492000, 1371495600, 1371499200, 
    1371502800, 1371506400, 1371510000, 1371513600, 1371517200, 1371520800, 
    1371524400, 1371528000, 1371531600, 1371535200, 1371538800, 1371542400, 
    1371546000, 1371549600, 1371553200, 1371556800, 1371560400, 1371564000, 
    1371567600, 1371571200, 1371574800, 1371578400, 1371582000, 1371585600, 
    1371589200, 1371592800, 1371596400, 1371600000, 1371603600, 1371607200, 
    1371610800, 1371614400, 1371618000, 1371621600, 1371625200, 1371628800, 
    1371632400, 1371636000, 1371639600, 1371643200, 1371646800, 1371650400, 
    1371654000, 1371657600, 1371661200, 1371664800, 1371668400, 1371672000, 
    1371675600, 1371679200, 1371682800, 1371686400, 1371690000, 1371693600, 
    1371697200, 1371700800, 1371704400, 1371708000, 1371711600, 1371715200, 
    1371718800, 1371722400, 1371726000, 1371729600, 1371733200, 1371736800, 
    1371740400, 1371744000, 1371747600, 1371751200, 1371754800, 1371758400, 
    1371762000, 1371765600, 1371769200, 1371772800, 1371776400, 1371780000, 
    1371783600, 1371787200, 1371790800, 1371794400, 1371798000, 1371801600, 
    1371805200, 1371808800, 1371812400, 1371816000, 1371819600, 1371823200, 
    1371826800, 1371830400, 1371834000, 1371837600, 1371841200, 1371844800, 
    1371848400, 1371852000, 1371855600, 1371859200, 1371862800, 1371866400, 
    1371870000, 1371873600, 1371877200, 1371880800, 1371884400, 1371888000, 
    1371891600, 1371895200, 1371898800, 1371902400, 1371906000, 1371909600, 
    1371913200, 1371916800, 1371920400, 1371924000, 1371927600, 1371931200, 
    1371934800, 1371938400, 1371942000, 1371945600, 1371949200, 1371952800, 
    1371956400, 1371960000, 1371963600, 1371967200, 1371970800, 1371974400, 
    1371978000, 1371981600, 1371985200, 1371988800, 1371992400, 1371996000, 
    1371999600, 1372003200, 1372006800, 1372010400, 1372014000, 1372017600, 
    1372021200, 1372024800, 1372028400, 1372032000, 1372035600, 1372039200, 
    1372042800, 1372046400, 1372050000, 1372053600, 1372057200, 1372060800, 
    1372064400, 1372068000, 1372071600, 1372075200, 1372078800, 1372082400, 
    1372086000, 1372089600, 1372093200, 1372096800, 1372100400, 1372104000, 
    1372107600, 1372111200, 1372114800, 1372118400, 1372122000, 1372125600, 
    1372129200, 1372132800, 1372136400, 1372140000, 1372143600, 1372147200, 
    1372150800, 1372154400, 1372158000, 1372161600, 1372165200, 1372168800, 
    1372172400, 1372176000, 1372179600, 1372183200, 1372186800, 1372190400, 
    1372194000, 1372197600, 1372201200, 1372204800, 1372208400, 1372212000, 
    1372215600, 1372219200, 1372222800, 1372226400, 1372230000, 1372233600, 
    1372237200, 1372240800, 1372244400, 1372248000, 1372251600, 1372255200, 
    1372258800, 1372262400, 1372266000, 1372269600, 1372273200, 1372276800, 
    1372280400, 1372284000, 1372287600, 1372291200, 1372294800, 1372298400, 
    1372302000, 1372305600, 1372309200, 1372312800, 1372316400, 1372320000, 
    1372323600, 1372327200, 1372330800, 1372334400, 1372338000, 1372341600, 
    1372345200, 1372348800, 1372352400, 1372356000, 1372359600, 1372363200, 
    1372366800, 1372370400, 1372374000, 1372377600, 1372381200, 1372384800, 
    1372388400, 1372392000, 1372395600, 1372399200, 1372402800, 1372406400, 
    1372410000, 1372413600, 1372417200, 1372420800, 1372424400, 1372428000, 
    1372431600, 1372435200, 1372438800, 1372442400, 1372446000, 1372449600, 
    1372453200, 1372456800, 1372460400, 1372464000, 1372467600, 1372471200, 
    1372474800, 1372478400, 1372482000, 1372485600, 1372489200, 1372492800, 
    1372496400, 1372500000, 1372503600, 1372507200, 1372510800, 1372514400, 
    1372518000, 1372521600, 1372525200, 1372528800, 1372532400, 1372536000, 
    1372539600, 1372543200, 1372546800, 1372550400, 1372554000, 1372557600, 
    1372561200, 1372564800, 1372568400, 1372572000, 1372575600, 1372579200, 
    1372582800, 1372586400, 1372590000, 1372593600, 1372597200, 1372600800, 
    1372604400, 1372608000, 1372611600, 1372615200, 1372618800, 1372622400, 
    1372626000, 1372629600, 1372633200, 1372636800, 1372640400, 1372644000, 
    1372647600, 1372651200, 1372654800, 1372658400, 1372662000, 1372665600, 
    1372669200, 1372672800, 1372676400, 1372680000, 1372683600, 1372687200, 
    1372690800, 1372694400, 1372698000, 1372701600, 1372705200, 1372708800, 
    1372712400, 1372716000, 1372719600, 1372723200, 1372726800, 1372730400, 
    1372734000, 1372737600, 1372741200, 1372744800, 1372748400, 1372752000, 
    1372755600, 1372759200, 1372762800, 1372766400, 1372770000, 1372773600, 
    1372777200, 1372780800, 1372784400, 1372788000, 1372791600, 1372795200, 
    1372798800, 1372802400, 1372806000, 1372809600, 1372813200, 1372816800, 
    1372820400, 1372824000, 1372827600, 1372831200, 1372834800, 1372838400, 
    1372842000, 1372845600, 1372849200, 1372852800, 1372856400, 1372860000, 
    1372863600, 1372867200, 1372870800, 1372874400, 1372878000, 1372881600, 
    1372885200, 1372888800, 1372892400, 1372896000, 1372899600, 1372903200, 
    1372906800, 1372910400, 1372914000, 1372917600, 1372921200, 1372924800, 
    1372928400, 1372932000, 1372935600, 1372939200, 1372942800, 1372946400, 
    1372950000, 1372953600, 1372957200, 1372960800, 1372964400, 1372968000, 
    1372971600, 1372975200, 1372978800, 1372982400, 1372986000, 1372989600, 
    1372993200, 1372996800, 1373000400, 1373004000, 1373007600, 1373011200, 
    1373014800, 1373018400, 1373022000, 1373025600, 1373029200, 1373032800, 
    1373036400, 1373040000, 1373043600, 1373047200, 1373050800, 1373054400, 
    1373058000, 1373061600, 1373065200, 1373068800, 1373072400, 1373076000, 
    1373079600, 1373083200, 1373086800, 1373090400, 1373094000, 1373097600, 
    1373101200, 1373104800, 1373108400, 1373112000, 1373115600, 1373119200, 
    1373122800, 1373126400, 1373130000, 1373133600, 1373137200, 1373140800, 
    1373144400, 1373148000, 1373151600, 1373155200, 1373158800, 1373162400, 
    1373166000, 1373169600, 1373173200, 1373176800, 1373180400, 1373184000, 
    1373187600, 1373191200, 1373194800, 1373198400, 1373202000, 1373205600, 
    1373209200, 1373212800, 1373216400, 1373220000, 1373223600, 1373227200, 
    1373230800, 1373234400, 1373238000, 1373241600, 1373245200, 1373248800, 
    1373252400, 1373256000, 1373259600, 1373263200, 1373266800, 1373270400, 
    1373274000, 1373277600, 1373281200, 1373284800, 1373288400, 1373292000, 
    1373295600, 1373299200, 1373302800, 1373306400, 1373310000, 1373313600, 
    1373317200, 1373320800, 1373324400, 1373328000, 1373331600, 1373335200, 
    1373338800, 1373342400, 1373346000, 1373349600, 1373353200, 1373356800, 
    1373360400, 1373364000, 1373367600, 1373371200, 1373374800, 1373378400, 
    1373382000, 1373385600, 1373389200, 1373392800, 1373396400, 1373400000, 
    1373403600, 1373407200, 1373410800, 1373414400, 1373418000, 1373421600, 
    1373425200, 1373428800, 1373432400, 1373436000, 1373439600, 1373443200, 
    1373446800, 1373450400, 1373454000, 1373457600, 1373461200, 1373464800, 
    1373468400, 1373472000, 1373475600, 1373479200, 1373482800, 1373486400, 
    1373490000, 1373493600, 1373497200, 1373500800, 1373504400, 1373508000, 
    1373511600, 1373515200, 1373518800, 1373522400, 1373526000, 1373529600, 
    1373533200, 1373536800, 1373540400, 1373544000, 1373547600, 1373551200, 
    1373554800, 1373558400, 1373562000, 1373565600, 1373569200, 1373572800, 
    1373576400, 1373580000, 1373583600, 1373587200, 1373590800, 1373594400, 
    1373598000, 1373601600, 1373605200, 1373608800, 1373612400, 1373616000, 
    1373619600, 1373623200, 1373626800, 1373630400, 1373634000, 1373637600, 
    1373641200, 1373644800, 1373648400, 1373652000, 1373655600, 1373659200, 
    1373662800, 1373666400, 1373670000, 1373673600, 1373677200, 1373680800, 
    1373684400, 1373688000, 1373691600, 1373695200, 1373698800, 1373702400, 
    1373706000, 1373709600, 1373713200, 1373716800, 1373720400, 1373724000, 
    1373727600, 1373731200, 1373734800, 1373738400, 1373742000, 1373745600, 
    1373749200, 1373752800, 1373756400, 1373760000, 1373763600, 1373767200, 
    1373770800, 1373774400, 1373778000, 1373781600, 1373785200, 1373788800, 
    1373792400, 1373796000, 1373799600, 1373803200, 1373806800, 1373810400, 
    1373814000, 1373817600, 1373821200, 1373824800, 1373828400, 1373832000, 
    1373835600, 1373839200, 1373842800, 1373846400, 1373850000, 1373853600, 
    1373857200, 1373860800, 1373864400, 1373868000, 1373871600, 1373875200, 
    1373878800, 1373882400, 1373886000, 1373889600, 1373893200, 1373896800, 
    1373900400, 1373904000, 1373907600, 1373911200, 1373914800, 1373918400, 
    1373922000, 1373925600, 1373929200, 1373932800, 1373936400, 1373940000, 
    1373943600, 1373947200, 1373950800, 1373954400, 1373958000, 1373961600, 
    1373965200, 1373968800, 1373972400, 1373976000, 1373979600, 1373983200, 
    1373986800, 1373990400, 1373994000, 1373997600, 1374001200, 1374004800, 
    1374008400, 1374012000, 1374015600, 1374019200, 1374022800, 1374026400, 
    1374030000, 1374033600, 1374037200, 1374040800, 1374044400, 1374048000, 
    1374051600, 1374055200, 1374058800, 1374062400, 1374066000, 1374069600, 
    1374073200, 1374076800, 1374080400, 1374084000, 1374087600, 1374091200, 
    1374094800, 1374098400, 1374102000, 1374105600, 1374109200, 1374112800, 
    1374116400, 1374120000, 1374123600, 1374127200, 1374130800, 1374134400, 
    1374138000, 1374141600, 1374145200, 1374148800, 1374152400, 1374156000, 
    1374159600, 1374163200, 1374166800, 1374170400, 1374174000, 1374177600, 
    1374181200, 1374184800, 1374188400, 1374192000, 1374195600, 1374199200, 
    1374202800, 1374206400, 1374210000, 1374213600, 1374217200, 1374220800, 
    1374224400, 1374228000, 1374231600, 1374235200, 1374238800, 1374242400, 
    1374246000, 1374249600, 1374253200, 1374256800, 1374260400, 1374264000, 
    1374267600, 1374271200, 1374274800, 1374278400, 1374282000, 1374285600, 
    1374289200, 1374292800, 1374296400, 1374300000, 1374303600, 1374307200, 
    1374310800, 1374314400, 1374318000, 1374321600, 1374325200, 1374328800, 
    1374332400, 1374336000, 1374339600, 1374343200, 1374346800, 1374350400, 
    1374354000, 1374357600, 1374361200, 1374364800, 1374368400, 1374372000, 
    1374375600, 1374379200, 1374382800, 1374386400, 1374390000, 1374393600, 
    1374397200, 1374400800, 1374404400, 1374408000, 1374411600, 1374415200, 
    1374418800, 1374422400, 1374426000, 1374429600, 1374433200, 1374436800, 
    1374440400, 1374444000, 1374447600, 1374451200, 1374454800, 1374458400, 
    1374462000, 1374465600, 1374469200, 1374472800, 1374476400, 1374480000, 
    1374483600, 1374487200, 1374490800, 1374494400, 1374498000, 1374501600, 
    1374505200, 1374508800, 1374512400, 1374516000, 1374519600, 1374523200, 
    1374526800, 1374530400, 1374534000, 1374537600, 1374541200, 1374544800, 
    1374548400, 1374552000, 1374555600, 1374559200, 1374562800, 1374566400, 
    1374570000, 1374573600, 1374577200, 1374580800, 1374584400, 1374588000, 
    1374591600, 1374595200, 1374598800, 1374602400, 1374606000, 1374609600, 
    1374613200, 1374616800, 1374620400, 1374624000, 1374627600, 1374631200, 
    1374634800, 1374638400, 1374642000, 1374645600, 1374649200, 1374652800, 
    1374656400, 1374660000, 1374663600, 1374667200, 1374670800, 1374674400, 
    1374678000, 1374681600, 1374685200, 1374688800, 1374692400, 1374696000, 
    1374699600, 1374703200, 1374706800, 1374710400, 1374714000, 1374717600, 
    1374721200, 1374724800, 1374728400, 1374732000, 1374735600, 1374739200, 
    1374742800, 1374746400, 1374750000, 1374753600, 1374757200, 1374760800, 
    1374764400, 1374768000, 1374771600, 1374775200, 1374778800, 1374782400, 
    1374786000, 1374789600, 1374793200, 1374796800, 1374800400, 1374804000, 
    1374807600, 1374811200, 1374814800, 1374818400, 1374822000, 1374825600, 
    1374829200, 1374832800, 1374836400, 1374840000, 1374843600, 1374847200, 
    1374850800, 1374854400, 1374858000, 1374861600, 1374865200, 1374868800, 
    1374872400, 1374876000, 1374879600, 1374883200, 1374886800, 1374890400, 
    1374894000, 1374897600, 1374901200, 1374904800, 1374908400, 1374912000, 
    1374915600, 1374919200, 1374922800, 1374926400, 1374930000, 1374933600, 
    1374937200, 1374940800, 1374944400, 1374948000, 1374951600, 1374955200, 
    1374958800, 1374962400, 1374966000, 1374969600, 1374973200, 1374976800, 
    1374980400, 1374984000, 1374987600, 1374991200, 1374994800, 1374998400, 
    1375002000, 1375005600, 1375009200, 1375012800, 1375016400, 1375020000, 
    1375023600, 1375027200, 1375030800, 1375034400, 1375038000, 1375041600, 
    1375045200, 1375048800, 1375052400, 1375056000, 1375059600, 1375063200, 
    1375066800, 1375070400, 1375074000, 1375077600, 1375081200, 1375084800, 
    1375088400, 1375092000, 1375095600, 1375099200, 1375102800, 1375106400, 
    1375110000, 1375113600, 1375117200, 1375120800, 1375124400, 1375128000, 
    1375131600, 1375135200, 1375138800, 1375142400, 1375146000, 1375149600, 
    1375153200, 1375156800, 1375160400, 1375164000, 1375167600, 1375171200, 
    1375174800, 1375178400, 1375182000, 1375185600, 1375189200, 1375192800, 
    1375196400, 1375200000, 1375203600, 1375207200, 1375210800, 1375214400, 
    1375218000, 1375221600, 1375225200, 1375228800, 1375232400, 1375236000, 
    1375239600, 1375243200, 1375246800, 1375250400, 1375254000, 1375257600, 
    1375261200, 1375264800, 1375268400, 1375272000, 1375275600, 1375279200, 
    1375282800, 1375286400, 1375290000, 1375293600, 1375297200, 1375300800, 
    1375304400, 1375308000, 1375311600, 1375315200, 1375318800, 1375322400, 
    1375326000, 1375329600, 1375333200, 1375336800, 1375340400, 1375344000, 
    1375347600, 1375351200, 1375354800, 1375358400, 1375362000, 1375365600, 
    1375369200, 1375372800, 1375376400, 1375380000, 1375383600, 1375387200, 
    1375390800, 1375394400, 1375398000, 1375401600, 1375405200, 1375408800, 
    1375412400, 1375416000, 1375419600, 1375423200, 1375426800, 1375430400, 
    1375434000, 1375437600, 1375441200, 1375444800, 1375448400, 1375452000, 
    1375455600, 1375459200, 1375462800, 1375466400, 1375470000, 1375473600, 
    1375477200, 1375480800, 1375484400, 1375488000, 1375491600, 1375495200, 
    1375498800, 1375502400, 1375506000, 1375509600, 1375513200, 1375516800, 
    1375520400, 1375524000, 1375527600, 1375531200, 1375534800, 1375538400, 
    1375542000, 1375545600, 1375549200, 1375552800, 1375556400, 1375560000, 
    1375563600, 1375567200, 1375570800, 1375574400, 1375578000, 1375581600, 
    1375585200, 1375588800, 1375592400, 1375596000, 1375599600, 1375603200, 
    1375606800, 1375610400, 1375614000, 1375617600, 1375621200, 1375624800, 
    1375628400, 1375632000, 1375635600, 1375639200, 1375642800, 1375646400, 
    1375650000, 1375653600, 1375657200, 1375660800, 1375664400, 1375668000, 
    1375671600, 1375675200, 1375678800, 1375682400, 1375686000, 1375689600, 
    1375693200, 1375696800, 1375700400, 1375704000, 1375707600, 1375711200, 
    1375714800, 1375718400, 1375722000, 1375725600, 1375729200, 1375732800, 
    1375736400, 1375740000, 1375743600, 1375747200, 1375750800, 1375754400, 
    1375758000, 1375761600, 1375765200, 1375768800, 1375772400, 1375776000, 
    1375779600, 1375783200, 1375786800, 1375790400, 1375794000, 1375797600, 
    1375801200, 1375804800, 1375808400, 1375812000, 1375815600, 1375819200, 
    1375822800, 1375826400, 1375830000, 1375833600, 1375837200, 1375840800, 
    1375844400, 1375848000, 1375851600, 1375855200, 1375858800, 1375862400, 
    1375866000, 1375869600, 1375873200, 1375876800, 1375880400, 1375884000, 
    1375887600, 1375891200, 1375894800, 1375898400, 1375902000, 1375905600, 
    1375909200, 1375912800, 1375916400, 1375920000, 1375923600, 1375927200, 
    1375930800, 1375934400, 1375938000, 1375941600, 1375945200, 1375948800, 
    1375952400, 1375956000, 1375959600, 1375963200, 1375966800, 1375970400, 
    1375974000, 1375977600, 1375981200, 1375984800, 1375988400, 1375992000, 
    1375995600, 1375999200, 1376002800, 1376006400, 1376010000, 1376013600, 
    1376017200, 1376020800, 1376024400, 1376028000, 1376031600, 1376035200, 
    1376038800, 1376042400, 1376046000, 1376049600, 1376053200, 1376056800, 
    1376060400, 1376064000, 1376067600, 1376071200, 1376074800, 1376078400, 
    1376082000, 1376085600, 1376089200, 1376092800, 1376096400, 1376100000, 
    1376103600, 1376107200, 1376110800, 1376114400, 1376118000, 1376121600, 
    1376125200, 1376128800, 1376132400, 1376136000, 1376139600, 1376143200, 
    1376146800, 1376150400, 1376154000, 1376157600, 1376161200, 1376164800, 
    1376168400, 1376172000, 1376175600, 1376179200, 1376182800, 1376186400, 
    1376190000, 1376193600, 1376197200, 1376200800, 1376204400, 1376208000, 
    1376211600, 1376215200, 1376218800, 1376222400, 1376226000, 1376229600, 
    1376233200, 1376236800, 1376240400, 1376244000, 1376247600, 1376251200, 
    1376254800, 1376258400, 1376262000, 1376265600, 1376269200, 1376272800, 
    1376276400, 1376280000, 1376283600, 1376287200, 1376290800, 1376294400, 
    1376298000, 1376301600, 1376305200, 1376308800, 1376312400, 1376316000, 
    1376319600, 1376323200, 1376326800, 1376330400, 1376334000, 1376337600, 
    1376341200, 1376344800, 1376348400, 1376352000, 1376355600, 1376359200, 
    1376362800, 1376366400, 1376370000, 1376373600, 1376377200, 1376380800, 
    1376384400, 1376388000, 1376391600, 1376395200, 1376398800, 1376402400, 
    1376406000, 1376409600, 1376413200, 1376416800, 1376420400, 1376424000, 
    1376427600, 1376431200, 1376434800, 1376438400, 1376442000, 1376445600, 
    1376449200, 1376452800, 1376456400, 1376460000, 1376463600, 1376467200, 
    1376470800, 1376474400, 1376478000, 1376481600, 1376485200, 1376488800, 
    1376492400, 1376496000, 1376499600, 1376503200, 1376506800, 1376510400, 
    1376514000, 1376517600, 1376521200, 1376524800, 1376528400, 1376532000, 
    1376535600, 1376539200, 1376542800, 1376546400, 1376550000, 1376553600, 
    1376557200, 1376560800, 1376564400, 1376568000, 1376571600, 1376575200, 
    1376578800, 1376582400, 1376586000, 1376589600, 1376593200, 1376596800, 
    1376600400, 1376604000, 1376607600, 1376611200, 1376614800, 1376618400, 
    1376622000, 1376625600, 1376629200, 1376632800, 1376636400, 1376640000, 
    1376643600, 1376647200, 1376650800, 1376654400, 1376658000, 1376661600, 
    1376665200, 1376668800, 1376672400, 1376676000, 1376679600, 1376683200, 
    1376686800, 1376690400, 1376694000, 1376697600, 1376701200, 1376704800, 
    1376708400, 1376712000, 1376715600, 1376719200, 1376722800, 1376726400, 
    1376730000, 1376733600, 1376737200, 1376740800, 1376744400, 1376748000, 
    1376751600, 1376755200, 1376758800, 1376762400, 1376766000, 1376769600, 
    1376773200, 1376776800, 1376780400, 1376784000, 1376787600, 1376791200, 
    1376794800, 1376798400, 1376802000, 1376805600, 1376809200, 1376812800, 
    1376816400, 1376820000, 1376823600, 1376827200, 1376830800, 1376834400, 
    1376838000, 1376841600, 1376845200, 1376848800, 1376852400, 1376856000, 
    1376859600, 1376863200, 1376866800, 1376870400, 1376874000, 1376877600, 
    1376881200, 1376884800, 1376888400, 1376892000, 1376895600, 1376899200, 
    1376902800, 1376906400, 1376910000, 1376913600, 1376917200, 1376920800, 
    1376924400, 1376928000, 1376931600, 1376935200, 1376938800, 1376942400, 
    1376946000, 1376949600, 1376953200, 1376956800, 1376960400, 1376964000, 
    1376967600, 1376971200, 1376974800, 1376978400, 1376982000, 1376985600, 
    1376989200, 1376992800, 1376996400, 1377000000, 1377003600, 1377007200, 
    1377010800, 1377014400, 1377018000, 1377021600, 1377025200, 1377028800, 
    1377032400, 1377036000, 1377039600, 1377043200, 1377046800, 1377050400, 
    1377054000, 1377057600, 1377061200, 1377064800, 1377068400, 1377072000, 
    1377075600, 1377079200, 1377082800, 1377086400, 1377090000, 1377093600, 
    1377097200, 1377100800, 1377104400, 1377108000, 1377111600, 1377115200, 
    1377118800, 1377122400, 1377126000, 1377129600, 1377133200, 1377136800, 
    1377140400, 1377144000, 1377147600, 1377151200, 1377154800, 1377158400, 
    1377162000, 1377165600, 1377169200, 1377172800, 1377176400, 1377180000, 
    1377183600, 1377187200, 1377190800, 1377194400, 1377198000, 1377201600, 
    1377205200, 1377208800, 1377212400, 1377216000, 1377219600, 1377223200, 
    1377226800, 1377230400, 1377234000, 1377237600, 1377241200, 1377244800, 
    1377248400, 1377252000, 1377255600, 1377259200, 1377262800, 1377266400, 
    1377270000, 1377273600, 1377277200, 1377280800, 1377284400, 1377288000, 
    1377291600, 1377295200, 1377298800, 1377302400, 1377306000, 1377309600, 
    1377313200, 1377316800, 1377320400, 1377324000, 1377327600, 1377331200, 
    1377334800, 1377338400, 1377342000, 1377345600, 1377349200, 1377352800, 
    1377356400, 1377360000, 1377363600, 1377367200, 1377370800, 1377374400, 
    1377378000, 1377381600, 1377385200, 1377388800, 1377392400, 1377396000, 
    1377399600, 1377403200, 1377406800, 1377410400, 1377414000, 1377417600, 
    1377421200, 1377424800, 1377428400, 1377432000, 1377435600, 1377439200, 
    1377442800, 1377446400, 1377450000, 1377453600, 1377457200, 1377460800, 
    1377464400, 1377468000, 1377471600, 1377475200, 1377478800, 1377482400, 
    1377486000, 1377489600, 1377493200, 1377496800, 1377500400, 1377504000, 
    1377507600, 1377511200, 1377514800, 1377518400, 1377522000, 1377525600, 
    1377529200, 1377532800, 1377536400, 1377540000, 1377543600, 1377547200, 
    1377550800, 1377554400, 1377558000, 1377561600, 1377565200, 1377568800, 
    1377572400, 1377576000, 1377579600, 1377583200, 1377586800, 1377590400, 
    1377594000, 1377597600, 1377601200, 1377604800, 1377608400, 1377612000, 
    1377615600, 1377619200, 1377622800, 1377626400, 1377630000, 1377633600, 
    1377637200, 1377640800, 1377644400, 1377648000, 1377651600, 1377655200, 
    1377658800, 1377662400, 1377666000, 1377669600, 1377673200, 1377676800, 
    1377680400, 1377684000, 1377687600, 1377691200, 1377694800, 1377698400, 
    1377702000, 1377705600, 1377709200, 1377712800, 1377716400, 1377720000, 
    1377723600, 1377727200, 1377730800, 1377734400, 1377738000, 1377741600, 
    1377745200, 1377748800, 1377752400, 1377756000, 1377759600, 1377763200, 
    1377766800, 1377770400, 1377774000, 1377777600, 1377781200, 1377784800, 
    1377788400, 1377792000, 1377795600, 1377799200, 1377802800, 1377806400, 
    1377810000, 1377813600, 1377817200, 1377820800, 1377824400, 1377828000, 
    1377831600, 1377835200, 1377838800, 1377842400, 1377846000, 1377849600, 
    1377853200, 1377856800, 1377860400, 1377864000, 1377867600, 1377871200, 
    1377874800, 1377878400, 1377882000, 1377885600, 1377889200, 1377892800, 
    1377896400, 1377900000, 1377903600, 1377907200, 1377910800, 1377914400, 
    1377918000, 1377921600, 1377925200, 1377928800, 1377932400, 1377936000, 
    1377939600, 1377943200, 1377946800, 1377950400, 1377954000, 1377957600, 
    1377961200, 1377964800, 1377968400, 1377972000, 1377975600, 1377979200, 
    1377982800, 1377986400, 1377990000, 1377993600, 1377997200, 1378000800, 
    1378004400, 1378008000, 1378011600, 1378015200, 1378018800, 1378022400, 
    1378026000, 1378029600, 1378033200, 1378036800, 1378040400, 1378044000, 
    1378047600, 1378051200, 1378054800, 1378058400, 1378062000, 1378065600, 
    1378069200, 1378072800, 1378076400, 1378080000, 1378083600, 1378087200, 
    1378090800, 1378094400, 1378098000, 1378101600, 1378105200, 1378108800, 
    1378112400, 1378116000, 1378119600, 1378123200, 1378126800, 1378130400, 
    1378134000, 1378137600, 1378141200, 1378144800, 1378148400, 1378152000, 
    1378155600, 1378159200, 1378162800, 1378166400, 1378170000, 1378173600, 
    1378177200, 1378180800, 1378184400, 1378188000, 1378191600, 1378195200, 
    1378198800, 1378202400, 1378206000, 1378209600, 1378213200, 1378216800, 
    1378220400, 1378224000, 1378227600, 1378231200, 1378234800, 1378238400, 
    1378242000, 1378245600, 1378249200, 1378252800, 1378256400, 1378260000, 
    1378263600, 1378267200, 1378270800, 1378274400, 1378278000, 1378281600, 
    1378285200, 1378288800, 1378292400, 1378296000, 1378299600, 1378303200, 
    1378306800, 1378310400, 1378314000, 1378317600, 1378321200, 1378324800, 
    1378328400, 1378332000, 1378335600, 1378339200, 1378342800, 1378346400, 
    1378350000, 1378353600, 1378357200, 1378360800, 1378364400, 1378368000, 
    1378371600, 1378375200, 1378378800, 1378382400, 1378386000, 1378389600, 
    1378393200, 1378396800, 1378400400, 1378404000, 1378407600, 1378411200, 
    1378414800, 1378418400, 1378422000, 1378425600, 1378429200, 1378432800, 
    1378436400, 1378440000, 1378443600, 1378447200, 1378450800, 1378454400, 
    1378458000, 1378461600, 1378465200, 1378468800, 1378472400, 1378476000, 
    1378479600, 1378483200, 1378486800, 1378490400, 1378494000, 1378497600, 
    1378501200, 1378504800, 1378508400, 1378512000, 1378515600, 1378519200, 
    1378522800, 1378526400, 1378530000, 1378533600, 1378537200, 1378540800, 
    1378544400, 1378548000, 1378551600, 1378555200, 1378558800, 1378562400, 
    1378566000, 1378569600, 1378573200, 1378576800, 1378580400, 1378584000, 
    1378587600, 1378591200, 1378594800, 1378598400, 1378602000, 1378605600, 
    1378609200, 1378612800, 1378616400, 1378620000, 1378623600, 1378627200, 
    1378630800, 1378634400, 1378638000, 1378641600, 1378645200, 1378648800, 
    1378652400, 1378656000, 1378659600, 1378663200, 1378666800, 1378670400, 
    1378674000, 1378677600, 1378681200, 1378684800, 1378688400, 1378692000, 
    1378695600, 1378699200, 1378702800, 1378706400, 1378710000, 1378713600, 
    1378717200, 1378720800, 1378724400, 1378728000, 1378731600, 1378735200, 
    1378738800, 1378742400, 1378746000, 1378749600, 1378753200, 1378756800, 
    1378760400, 1378764000, 1378767600, 1378771200, 1378774800, 1378778400, 
    1378782000, 1378785600, 1378789200, 1378792800, 1378796400, 1378800000, 
    1378803600, 1378807200, 1378810800, 1378814400, 1378818000, 1378821600, 
    1378825200, 1378828800, 1378832400, 1378836000, 1378839600, 1378843200, 
    1378846800, 1378850400, 1378854000, 1378857600, 1378861200, 1378864800, 
    1378868400, 1378872000, 1378875600, 1378879200, 1378882800, 1378886400, 
    1378890000, 1378893600, 1378897200, 1378900800, 1378904400, 1378908000, 
    1378911600, 1378915200, 1378918800, 1378922400, 1378926000, 1378929600, 
    1378933200, 1378936800, 1378940400, 1378944000, 1378947600, 1378951200, 
    1378954800, 1378958400, 1378962000, 1378965600, 1378969200, 1378972800, 
    1378976400, 1378980000, 1378983600, 1378987200, 1378990800, 1378994400, 
    1378998000, 1379001600, 1379005200, 1379008800, 1379012400, 1379016000, 
    1379019600, 1379023200, 1379026800, 1379030400, 1379034000, 1379037600, 
    1379041200, 1379044800, 1379048400, 1379052000, 1379055600, 1379059200, 
    1379062800, 1379066400, 1379070000, 1379073600, 1379077200, 1379080800, 
    1379084400, 1379088000, 1379091600, 1379095200, 1379098800, 1379102400, 
    1379106000, 1379109600, 1379113200, 1379116800, 1379120400, 1379124000, 
    1379127600, 1379131200, 1379134800, 1379138400, 1379142000, 1379145600, 
    1379149200, 1379152800, 1379156400, 1379160000, 1379163600, 1379167200, 
    1379170800, 1379174400, 1379178000, 1379181600, 1379185200, 1379188800, 
    1379192400, 1379196000, 1379199600, 1379203200, 1379206800, 1379210400, 
    1379214000, 1379217600, 1379221200, 1379224800, 1379228400, 1379232000, 
    1379235600, 1379239200, 1379242800, 1379246400, 1379250000, 1379253600, 
    1379257200, 1379260800, 1379264400, 1379268000, 1379271600, 1379275200, 
    1379278800, 1379282400, 1379286000, 1379289600, 1379293200, 1379296800, 
    1379300400, 1379304000, 1379307600, 1379311200, 1379314800, 1379318400, 
    1379322000, 1379325600, 1379329200, 1379332800, 1379336400, 1379340000, 
    1379343600, 1379347200, 1379350800, 1379354400, 1379358000, 1379361600, 
    1379365200, 1379368800, 1379372400, 1379376000, 1379379600, 1379383200, 
    1379386800, 1379390400, 1379394000, 1379397600, 1379401200, 1379404800, 
    1379408400, 1379412000, 1379415600, 1379419200, 1379422800, 1379426400, 
    1379430000, 1379433600, 1379437200, 1379440800, 1379444400, 1379448000, 
    1379451600, 1379455200, 1379458800, 1379462400, 1379466000, 1379469600, 
    1379473200, 1379476800, 1379480400, 1379484000, 1379487600, 1379491200, 
    1379494800, 1379498400, 1379502000, 1379505600, 1379509200, 1379512800, 
    1379516400, 1379520000, 1379523600, 1379527200, 1379530800, 1379534400, 
    1379538000, 1379541600, 1379545200, 1379548800, 1379552400, 1379556000, 
    1379559600, 1379563200, 1379566800, 1379570400, 1379574000, 1379577600, 
    1379581200, 1379584800, 1379588400, 1379592000, 1379595600, 1379599200, 
    1379602800, 1379606400, 1379610000, 1379613600, 1379617200, 1379620800, 
    1379624400, 1379628000, 1379631600, 1379635200, 1379638800, 1379642400, 
    1379646000, 1379649600, 1379653200, 1379656800, 1379660400, 1379664000, 
    1379667600, 1379671200, 1379674800, 1379678400, 1379682000, 1379685600, 
    1379689200, 1379692800, 1379696400, 1379700000, 1379703600, 1379707200, 
    1379710800, 1379714400, 1379718000, 1379721600, 1379725200, 1379728800, 
    1379732400, 1379736000, 1379739600, 1379743200, 1379746800, 1379750400, 
    1379754000, 1379757600, 1379761200, 1379764800, 1379768400, 1379772000, 
    1379775600, 1379779200, 1379782800, 1379786400, 1379790000, 1379793600, 
    1379797200, 1379800800, 1379804400, 1379808000, 1379811600, 1379815200, 
    1379818800, 1379822400, 1379826000, 1379829600, 1379833200, 1379836800, 
    1379840400, 1379844000, 1379847600, 1379851200, 1379854800, 1379858400, 
    1379862000, 1379865600, 1379869200, 1379872800, 1379876400, 1379880000, 
    1379883600, 1379887200, 1379890800, 1379894400, 1379898000, 1379901600, 
    1379905200, 1379908800, 1379912400, 1379916000, 1379919600, 1379923200, 
    1379926800, 1379930400, 1379934000, 1379937600, 1379941200, 1379944800, 
    1379948400, 1379952000, 1379955600, 1379959200, 1379962800, 1379966400, 
    1379970000, 1379973600, 1379977200, 1379980800, 1379984400, 1379988000, 
    1379991600, 1379995200, 1379998800, 1380002400, 1380006000, 1380009600, 
    1380013200, 1380016800, 1380020400, 1380024000, 1380027600, 1380031200, 
    1380034800, 1380038400, 1380042000, 1380045600, 1380049200, 1380052800, 
    1380056400, 1380060000, 1380063600, 1380067200, 1380070800, 1380074400, 
    1380078000, 1380081600, 1380085200, 1380088800, 1380092400, 1380096000, 
    1380099600, 1380103200, 1380106800, 1380110400, 1380114000, 1380117600, 
    1380121200, 1380124800, 1380128400, 1380132000, 1380135600, 1380139200, 
    1380142800, 1380146400, 1380150000, 1380153600, 1380157200, 1380160800, 
    1380164400, 1380168000, 1380171600, 1380175200, 1380178800, 1380182400, 
    1380186000, 1380189600, 1380193200, 1380196800, 1380200400, 1380204000, 
    1380207600, 1380211200, 1380214800, 1380218400, 1380222000, 1380225600, 
    1380229200, 1380232800, 1380236400, 1380240000, 1380243600, 1380247200, 
    1380250800, 1380254400, 1380258000, 1380261600, 1380265200, 1380268800, 
    1380272400, 1380276000, 1380279600, 1380283200, 1380286800, 1380290400, 
    1380294000, 1380297600, 1380301200, 1380304800, 1380308400, 1380312000, 
    1380315600, 1380319200, 1380322800, 1380326400, 1380330000, 1380333600, 
    1380337200, 1380340800, 1380344400, 1380348000, 1380351600, 1380355200, 
    1380358800, 1380362400, 1380366000, 1380369600, 1380373200, 1380376800, 
    1380380400, 1380384000, 1380387600, 1380391200, 1380394800, 1380398400, 
    1380402000, 1380405600, 1380409200, 1380412800, 1380416400, 1380420000, 
    1380423600, 1380427200, 1380430800, 1380434400, 1380438000, 1380441600, 
    1380445200, 1380448800, 1380452400, 1380456000, 1380459600, 1380463200, 
    1380466800, 1380470400, 1380474000, 1380477600, 1380481200, 1380484800, 
    1380488400, 1380492000, 1380495600, 1380499200, 1380502800, 1380506400, 
    1380510000, 1380513600, 1380517200, 1380520800, 1380524400, 1380528000, 
    1380531600, 1380535200, 1380538800, 1380542400, 1380546000, 1380549600, 
    1380553200, 1380556800, 1380560400, 1380564000, 1380567600, 1380571200, 
    1380574800, 1380578400, 1380582000, 1380585600, 1380589200, 1380592800, 
    1380596400, 1380600000, 1380603600, 1380607200, 1380610800, 1380614400, 
    1380618000, 1380621600, 1380625200, 1380628800, 1380632400, 1380636000, 
    1380639600, 1380643200, 1380646800, 1380650400, 1380654000, 1380657600, 
    1380661200, 1380664800, 1380668400, 1380672000, 1380675600, 1380679200, 
    1380682800, 1380686400, 1380690000, 1380693600, 1380697200, 1380700800, 
    1380704400, 1380708000, 1380711600, 1380715200, 1380718800, 1380722400, 
    1380726000, 1380729600, 1380733200, 1380736800, 1380740400, 1380744000, 
    1380747600, 1380751200, 1380754800, 1380758400, 1380762000, 1380765600, 
    1380769200, 1380772800, 1380776400, 1380780000, 1380783600, 1380787200, 
    1380790800, 1380794400, 1380798000, 1380801600, 1380805200, 1380808800, 
    1380812400, 1380816000, 1380819600, 1380823200, 1380826800, 1380830400, 
    1380834000, 1380837600, 1380841200, 1380844800, 1380848400, 1380852000, 
    1380855600, 1380859200, 1380862800, 1380866400, 1380870000, 1380873600, 
    1380877200, 1380880800, 1380884400, 1380888000, 1380891600, 1380895200, 
    1380898800, 1380902400, 1380906000, 1380909600, 1380913200, 1380916800, 
    1380920400, 1380924000, 1380927600, 1380931200, 1380934800, 1380938400, 
    1380942000, 1380945600, 1380949200, 1380952800, 1380956400, 1380960000, 
    1380963600, 1380967200, 1380970800, 1380974400, 1380978000, 1380981600, 
    1380985200, 1380988800, 1380992400, 1380996000, 1380999600, 1381003200, 
    1381006800, 1381010400, 1381014000, 1381017600, 1381021200, 1381024800, 
    1381028400, 1381032000, 1381035600, 1381039200, 1381042800, 1381046400, 
    1381050000, 1381053600, 1381057200, 1381060800, 1381064400, 1381068000, 
    1381071600, 1381075200, 1381078800, 1381082400, 1381086000, 1381089600, 
    1381093200, 1381096800, 1381100400, 1381104000, 1381107600, 1381111200, 
    1381114800, 1381118400, 1381122000, 1381125600, 1381129200, 1381132800, 
    1381136400, 1381140000, 1381143600, 1381147200, 1381150800, 1381154400, 
    1381158000, 1381161600, 1381165200, 1381168800, 1381172400, 1381176000, 
    1381179600, 1381183200, 1381186800, 1381190400, 1381194000, 1381197600, 
    1381201200, 1381204800, 1381208400, 1381212000, 1381215600, 1381219200, 
    1381222800, 1381226400, 1381230000, 1381233600, 1381237200, 1381240800, 
    1381244400, 1381248000, 1381251600, 1381255200, 1381258800, 1381262400, 
    1381266000, 1381269600, 1381273200, 1381276800, 1381280400, 1381284000, 
    1381287600, 1381291200, 1381294800, 1381298400, 1381302000, 1381305600, 
    1381309200, 1381312800, 1381316400, 1381320000, 1381323600, 1381327200, 
    1381330800, 1381334400, 1381338000, 1381341600, 1381345200, 1381348800, 
    1381352400, 1381356000, 1381359600, 1381363200, 1381366800, 1381370400, 
    1381374000, 1381377600, 1381381200, 1381384800, 1381388400, 1381392000, 
    1381395600, 1381399200, 1381402800, 1381406400, 1381410000, 1381413600, 
    1381417200, 1381420800, 1381424400, 1381428000, 1381431600, 1381435200, 
    1381438800, 1381442400, 1381446000, 1381449600, 1381453200, 1381456800, 
    1381460400, 1381464000, 1381467600, 1381471200, 1381474800, 1381478400, 
    1381482000, 1381485600, 1381489200, 1381492800, 1381496400, 1381500000, 
    1381503600, 1381507200, 1381510800, 1381514400, 1381518000, 1381521600, 
    1381525200, 1381528800, 1381532400, 1381536000, 1381539600, 1381543200, 
    1381546800, 1381550400, 1381554000, 1381557600, 1381561200, 1381564800, 
    1381568400, 1381572000, 1381575600, 1381579200, 1381582800, 1381586400, 
    1381590000, 1381593600, 1381597200, 1381600800, 1381604400, 1381608000, 
    1381611600, 1381615200, 1381618800, 1381622400, 1381626000, 1381629600, 
    1381633200, 1381636800, 1381640400, 1381644000, 1381647600, 1381651200, 
    1381654800, 1381658400, 1381662000, 1381665600, 1381669200, 1381672800, 
    1381676400, 1381680000, 1381683600, 1381687200, 1381690800, 1381694400, 
    1381698000, 1381701600, 1381705200, 1381708800, 1381712400, 1381716000, 
    1381719600, 1381723200, 1381726800, 1381730400, 1381734000, 1381737600, 
    1381741200, 1381744800, 1381748400, 1381752000, 1381755600, 1381759200, 
    1381762800, 1381766400, 1381770000, 1381773600, 1381777200, 1381780800, 
    1381784400, 1381788000, 1381791600, 1381795200, 1381798800, 1381802400, 
    1381806000, 1381809600, 1381813200, 1381816800, 1381820400, 1381824000, 
    1381827600, 1381831200, 1381834800, 1381838400, 1381842000, 1381845600, 
    1381849200, 1381852800, 1381856400, 1381860000, 1381863600, 1381867200, 
    1381870800, 1381874400, 1381878000, 1381881600, 1381885200, 1381888800, 
    1381892400, 1381896000, 1381899600, 1381903200, 1381906800, 1381910400, 
    1381914000, 1381917600, 1381921200, 1381924800, 1381928400, 1381932000, 
    1381935600, 1381939200, 1381942800, 1381946400, 1381950000, 1381953600, 
    1381957200, 1381960800, 1381964400, 1381968000, 1381971600, 1381975200, 
    1381978800, 1381982400, 1381986000, 1381989600, 1381993200, 1381996800, 
    1382000400, 1382004000, 1382007600, 1382011200, 1382014800, 1382018400, 
    1382022000, 1382025600, 1382029200, 1382032800, 1382036400, 1382040000, 
    1382043600, 1382047200, 1382050800, 1382054400, 1382058000, 1382061600, 
    1382065200, 1382068800, 1382072400, 1382076000, 1382079600, 1382083200, 
    1382086800, 1382090400, 1382094000, 1382097600, 1382101200, 1382104800, 
    1382108400, 1382112000, 1382115600, 1382119200, 1382122800, 1382126400, 
    1382130000, 1382133600, 1382137200, 1382140800, 1382144400, 1382148000, 
    1382151600, 1382155200, 1382158800, 1382162400, 1382166000, 1382169600, 
    1382173200, 1382176800, 1382180400, 1382184000, 1382187600, 1382191200, 
    1382194800, 1382198400, 1382202000, 1382205600, 1382209200, 1382212800, 
    1382216400, 1382220000, 1382223600, 1382227200, 1382230800, 1382234400, 
    1382238000, 1382241600, 1382245200, 1382248800, 1382252400, 1382256000, 
    1382259600, 1382263200, 1382266800, 1382270400, 1382274000, 1382277600, 
    1382281200, 1382284800, 1382288400, 1382292000, 1382295600, 1382299200, 
    1382302800, 1382306400, 1382310000, 1382313600, 1382317200, 1382320800, 
    1382324400, 1382328000, 1382331600, 1382335200, 1382338800, 1382342400, 
    1382346000, 1382349600, 1382353200, 1382356800, 1382360400, 1382364000, 
    1382367600, 1382371200, 1382374800, 1382378400, 1382382000, 1382385600, 
    1382389200, 1382392800, 1382396400, 1382400000, 1382403600, 1382407200, 
    1382410800, 1382414400, 1382418000, 1382421600, 1382425200, 1382428800, 
    1382432400, 1382436000, 1382439600, 1382443200, 1382446800, 1382450400, 
    1382454000, 1382457600, 1382461200, 1382464800, 1382468400, 1382472000, 
    1382475600, 1382479200, 1382482800, 1382486400, 1382490000, 1382493600, 
    1382497200, 1382500800, 1382504400, 1382508000, 1382511600, 1382515200, 
    1382518800, 1382522400, 1382526000, 1382529600, 1382533200, 1382536800, 
    1382540400, 1382544000, 1382547600, 1382551200, 1382554800, 1382558400, 
    1382562000, 1382565600, 1382569200, 1382572800, 1382576400, 1382580000, 
    1382583600, 1382587200, 1382590800, 1382594400, 1382598000, 1382601600, 
    1382605200, 1382608800, 1382612400, 1382616000, 1382619600, 1382623200, 
    1382626800, 1382630400, 1382634000, 1382637600, 1382641200, 1382644800, 
    1382648400, 1382652000, 1382655600, 1382659200, 1382662800, 1382666400, 
    1382670000, 1382673600, 1382677200, 1382680800, 1382684400, 1382688000, 
    1382691600, 1382695200, 1382698800, 1382702400, 1382706000, 1382709600, 
    1382713200, 1382716800, 1382720400, 1382724000, 1382727600, 1382731200, 
    1382734800, 1382738400, 1382742000, 1382745600, 1382749200, 1382752800, 
    1382756400, 1382760000, 1382763600, 1382767200, 1382770800, 1382774400, 
    1382778000, 1382781600, 1382785200, 1382788800, 1382792400, 1382796000, 
    1382799600, 1382803200, 1382806800, 1382810400, 1382814000, 1382817600, 
    1382821200, 1382824800, 1382828400, 1382832000, 1382835600, 1382839200, 
    1382842800, 1382846400, 1382850000, 1382853600, 1382857200, 1382860800, 
    1382864400, 1382868000, 1382871600, 1382875200, 1382878800, 1382882400, 
    1382886000, 1382889600, 1382893200, 1382896800, 1382900400, 1382904000, 
    1382907600, 1382911200, 1382914800, 1382918400, 1382922000, 1382925600, 
    1382929200, 1382932800, 1382936400, 1382940000, 1382943600, 1382947200, 
    1382950800, 1382954400, 1382958000, 1382961600, 1382965200, 1382968800, 
    1382972400, 1382976000, 1382979600, 1382983200, 1382986800, 1382990400, 
    1382994000, 1382997600, 1383001200, 1383004800, 1383008400, 1383012000, 
    1383015600, 1383019200, 1383022800, 1383026400, 1383030000, 1383033600, 
    1383037200, 1383040800, 1383044400, 1383048000, 1383051600, 1383055200, 
    1383058800, 1383062400, 1383066000, 1383069600, 1383073200, 1383076800, 
    1383080400, 1383084000, 1383087600, 1383091200, 1383094800, 1383098400, 
    1383102000, 1383105600, 1383109200, 1383112800, 1383116400, 1383120000, 
    1383123600, 1383127200, 1383130800, 1383134400, 1383138000, 1383141600, 
    1383145200, 1383148800, 1383152400, 1383156000, 1383159600, 1383163200, 
    1383166800, 1383170400, 1383174000, 1383177600, 1383181200, 1383184800, 
    1383188400, 1383192000, 1383195600, 1383199200, 1383202800, 1383206400, 
    1383210000, 1383213600, 1383217200, 1383220800, 1383224400, 1383228000, 
    1383231600, 1383235200, 1383238800, 1383242400, 1383246000, 1383249600, 
    1383253200, 1383256800, 1383260400, 1383264000, 1383267600, 1383271200, 
    1383274800, 1383278400, 1383282000, 1383285600, 1383289200, 1383292800, 
    1383296400, 1383300000, 1383303600, 1383307200, 1383310800, 1383314400, 
    1383318000, 1383321600, 1383325200, 1383328800, 1383332400, 1383336000, 
    1383339600, 1383343200, 1383346800, 1383350400, 1383354000, 1383357600, 
    1383361200, 1383364800, 1383368400, 1383372000, 1383375600, 1383379200, 
    1383382800, 1383386400, 1383390000, 1383393600, 1383397200, 1383400800, 
    1383404400, 1383408000, 1383411600, 1383415200, 1383418800, 1383422400, 
    1383426000, 1383429600, 1383433200, 1383436800, 1383440400, 1383444000, 
    1383447600, 1383451200, 1383454800, 1383458400, 1383462000, 1383465600, 
    1383469200, 1383472800, 1383476400, 1383480000, 1383483600, 1383487200, 
    1383490800, 1383494400, 1383498000, 1383501600, 1383505200, 1383508800, 
    1383512400, 1383516000, 1383519600, 1383523200, 1383526800, 1383530400, 
    1383534000, 1383537600, 1383541200, 1383544800, 1383548400, 1383552000, 
    1383555600, 1383559200, 1383562800, 1383566400, 1383570000, 1383573600, 
    1383577200, 1383580800, 1383584400, 1383588000, 1383591600, 1383595200, 
    1383598800, 1383602400, 1383606000, 1383609600, 1383613200, 1383616800, 
    1383620400, 1383624000, 1383627600, 1383631200, 1383634800, 1383638400, 
    1383642000, 1383645600, 1383649200, 1383652800, 1383656400, 1383660000, 
    1383663600, 1383667200, 1383670800, 1383674400, 1383678000, 1383681600, 
    1383685200, 1383688800, 1383692400, 1383696000, 1383699600, 1383703200, 
    1383706800, 1383710400, 1383714000, 1383717600, 1383721200, 1383724800, 
    1383728400, 1383732000, 1383735600, 1383739200, 1383742800, 1383746400, 
    1383750000, 1383753600, 1383757200, 1383760800, 1383764400, 1383768000, 
    1383771600, 1383775200, 1383778800, 1383782400, 1383786000, 1383789600, 
    1383793200, 1383796800, 1383800400, 1383804000, 1383807600, 1383811200, 
    1383814800, 1383818400, 1383822000, 1383825600, 1383829200, 1383832800, 
    1383836400, 1383840000, 1383843600, 1383847200, 1383850800, 1383854400, 
    1383858000, 1383861600, 1383865200, 1383868800, 1383872400, 1383876000, 
    1383879600, 1383883200, 1383886800, 1383890400, 1383894000, 1383897600, 
    1383901200, 1383904800, 1383908400, 1383912000, 1383915600, 1383919200, 
    1383922800, 1383926400, 1383930000, 1383933600, 1383937200, 1383940800, 
    1383944400, 1383948000, 1383951600, 1383955200, 1383958800, 1383962400, 
    1383966000, 1383969600, 1383973200, 1383976800, 1383980400, 1383984000, 
    1383987600, 1383991200, 1383994800, 1383998400, 1384002000, 1384005600, 
    1384009200, 1384012800, 1384016400, 1384020000, 1384023600, 1384027200, 
    1384030800, 1384034400, 1384038000, 1384041600, 1384045200, 1384048800, 
    1384052400, 1384056000, 1384059600, 1384063200, 1384066800, 1384070400, 
    1384074000, 1384077600, 1384081200, 1384084800, 1384088400, 1384092000, 
    1384095600, 1384099200, 1384102800, 1384106400, 1384110000, 1384113600, 
    1384117200, 1384120800, 1384124400, 1384128000, 1384131600, 1384135200, 
    1384138800, 1384142400, 1384146000, 1384149600, 1384153200, 1384156800, 
    1384160400, 1384164000, 1384167600, 1384171200, 1384174800, 1384178400, 
    1384182000, 1384185600, 1384189200, 1384192800, 1384196400, 1384200000, 
    1384203600, 1384207200, 1384210800, 1384214400, 1384218000, 1384221600, 
    1384225200, 1384228800, 1384232400, 1384236000, 1384239600, 1384243200, 
    1384246800, 1384250400, 1384254000, 1384257600, 1384261200, 1384264800, 
    1384268400, 1384272000, 1384275600, 1384279200, 1384282800, 1384286400, 
    1384290000, 1384293600, 1384297200, 1384300800, 1384304400, 1384308000, 
    1384311600, 1384315200, 1384318800, 1384322400, 1384326000, 1384329600, 
    1384333200, 1384336800, 1384340400, 1384344000, 1384347600, 1384351200, 
    1384354800, 1384358400, 1384362000, 1384365600, 1384369200, 1384372800, 
    1384376400, 1384380000, 1384383600, 1384387200, 1384390800, 1384394400, 
    1384398000, 1384401600, 1384405200, 1384408800, 1384412400, 1384416000, 
    1384419600, 1384423200, 1384426800, 1384430400, 1384434000, 1384437600, 
    1384441200, 1384444800, 1384448400, 1384452000, 1384455600, 1384459200, 
    1384462800, 1384466400, 1384470000, 1384473600, 1384477200, 1384480800, 
    1384484400, 1384488000, 1384491600, 1384495200, 1384498800, 1384502400, 
    1384506000, 1384509600, 1384513200, 1384516800, 1384520400, 1384524000, 
    1384527600, 1384531200, 1384534800, 1384538400, 1384542000, 1384545600, 
    1384549200, 1384552800, 1384556400, 1384560000, 1384563600, 1384567200, 
    1384570800, 1384574400, 1384578000, 1384581600, 1384585200, 1384588800, 
    1384592400, 1384596000, 1384599600, 1384603200, 1384606800, 1384610400, 
    1384614000, 1384617600, 1384621200, 1384624800, 1384628400, 1384632000, 
    1384635600, 1384639200, 1384642800, 1384646400, 1384650000, 1384653600, 
    1384657200, 1384660800, 1384664400, 1384668000, 1384671600, 1384675200, 
    1384678800, 1384682400, 1384686000, 1384689600, 1384693200, 1384696800, 
    1384700400, 1384704000, 1384707600, 1384711200, 1384714800, 1384718400, 
    1384722000, 1384725600, 1384729200, 1384732800, 1384736400, 1384740000, 
    1384743600, 1384747200, 1384750800, 1384754400, 1384758000, 1384761600, 
    1384765200, 1384768800, 1384772400, 1384776000, 1384779600, 1384783200, 
    1384786800, 1384790400, 1384794000, 1384797600, 1384801200, 1384804800, 
    1384808400, 1384812000, 1384815600, 1384819200, 1384822800, 1384826400, 
    1384830000, 1384833600, 1384837200, 1384840800, 1384844400, 1384848000, 
    1384851600, 1384855200, 1384858800, 1384862400, 1384866000, 1384869600, 
    1384873200, 1384876800, 1384880400, 1384884000, 1384887600, 1384891200, 
    1384894800, 1384898400, 1384902000, 1384905600, 1384909200, 1384912800, 
    1384916400, 1384920000, 1384923600, 1384927200, 1384930800, 1384934400, 
    1384938000, 1384941600, 1384945200, 1384948800, 1384952400, 1384956000, 
    1384959600, 1384963200, 1384966800, 1384970400, 1384974000, 1384977600, 
    1384981200, 1384984800, 1384988400, 1384992000, 1384995600, 1384999200, 
    1385002800, 1385006400, 1385010000, 1385013600, 1385017200, 1385020800, 
    1385024400, 1385028000, 1385031600, 1385035200, 1385038800, 1385042400, 
    1385046000, 1385049600, 1385053200, 1385056800, 1385060400, 1385064000, 
    1385067600, 1385071200, 1385074800, 1385078400, 1385082000, 1385085600, 
    1385089200, 1385092800, 1385096400, 1385100000, 1385103600, 1385107200, 
    1385110800, 1385114400, 1385118000, 1385121600, 1385125200, 1385128800, 
    1385132400, 1385136000, 1385139600, 1385143200, 1385146800, 1385150400, 
    1385154000, 1385157600, 1385161200, 1385164800, 1385168400, 1385172000, 
    1385175600, 1385179200, 1385182800, 1385186400, 1385190000, 1385193600, 
    1385197200, 1385200800, 1385204400, 1385208000, 1385211600, 1385215200, 
    1385218800, 1385222400, 1385226000, 1385229600, 1385233200, 1385236800, 
    1385240400, 1385244000, 1385247600, 1385251200, 1385254800, 1385258400, 
    1385262000, 1385265600, 1385269200, 1385272800, 1385276400, 1385280000, 
    1385283600, 1385287200, 1385290800, 1385294400, 1385298000, 1385301600, 
    1385305200, 1385308800, 1385312400, 1385316000, 1385319600, 1385323200, 
    1385326800, 1385330400, 1385334000, 1385337600, 1385341200, 1385344800, 
    1385348400, 1385352000, 1385355600, 1385359200, 1385362800, 1385366400, 
    1385370000, 1385373600, 1385377200, 1385380800, 1385384400, 1385388000, 
    1385391600, 1385395200, 1385398800, 1385402400, 1385406000, 1385409600, 
    1385413200, 1385416800, 1385420400, 1385424000, 1385427600, 1385431200, 
    1385434800, 1385438400, 1385442000, 1385445600, 1385449200, 1385452800, 
    1385456400, 1385460000, 1385463600, 1385467200, 1385470800, 1385474400, 
    1385478000, 1385481600, 1385485200, 1385488800, 1385492400, 1385496000, 
    1385499600, 1385503200, 1385506800, 1385510400, 1385514000, 1385517600, 
    1385521200, 1385524800, 1385528400, 1385532000, 1385535600, 1385539200, 
    1385542800, 1385546400, 1385550000, 1385553600, 1385557200, 1385560800, 
    1385564400, 1385568000, 1385571600, 1385575200, 1385578800, 1385582400, 
    1385586000, 1385589600, 1385593200, 1385596800, 1385600400, 1385604000, 
    1385607600, 1385611200, 1385614800, 1385618400, 1385622000, 1385625600, 
    1385629200, 1385632800, 1385636400, 1385640000, 1385643600, 1385647200, 
    1385650800, 1385654400, 1385658000, 1385661600, 1385665200, 1385668800, 
    1385672400, 1385676000, 1385679600, 1385683200, 1385686800, 1385690400, 
    1385694000, 1385697600, 1385701200, 1385704800, 1385708400, 1385712000, 
    1385715600, 1385719200, 1385722800, 1385726400, 1385730000, 1385733600, 
    1385737200, 1385740800, 1385744400, 1385748000, 1385751600, 1385755200, 
    1385758800, 1385762400, 1385766000, 1385769600, 1385773200, 1385776800, 
    1385780400, 1385784000, 1385787600, 1385791200, 1385794800, 1385798400, 
    1385802000, 1385805600, 1385809200, 1385812800, 1385816400, 1385820000, 
    1385823600, 1385827200, 1385830800, 1385834400, 1385838000, 1385841600, 
    1385845200, 1385848800, 1385852400, 1385856000, 1385859600, 1385863200, 
    1385866800, 1385870400, 1385874000, 1385877600, 1385881200, 1385884800, 
    1385888400, 1385892000, 1385895600, 1385899200, 1385902800, 1385906400, 
    1385910000, 1385913600, 1385917200, 1385920800, 1385924400, 1385928000, 
    1385931600, 1385935200, 1385938800, 1385942400, 1385946000, 1385949600, 
    1385953200, 1385956800, 1385960400, 1385964000, 1385967600, 1385971200, 
    1385974800, 1385978400, 1385982000, 1385985600, 1385989200, 1385992800, 
    1385996400, 1386000000, 1386003600, 1386007200, 1386010800, 1386014400, 
    1386018000, 1386021600, 1386025200, 1386028800, 1386032400, 1386036000, 
    1386039600, 1386043200, 1386046800, 1386050400, 1386054000, 1386057600, 
    1386061200, 1386064800, 1386068400, 1386072000, 1386075600, 1386079200, 
    1386082800, 1386086400, 1386090000, 1386093600, 1386097200, 1386100800, 
    1386104400, 1386108000, 1386111600, 1386115200, 1386118800, 1386122400, 
    1386126000, 1386129600, 1386133200, 1386136800, 1386140400, 1386144000, 
    1386147600, 1386151200, 1386154800, 1386158400, 1386162000, 1386165600, 
    1386169200, 1386172800, 1386176400, 1386180000, 1386183600, 1386187200, 
    1386190800, 1386194400, 1386198000, 1386201600, 1386205200, 1386208800, 
    1386212400, 1386216000, 1386219600, 1386223200, 1386226800, 1386230400, 
    1386234000, 1386237600, 1386241200, 1386244800, 1386248400, 1386252000, 
    1386255600, 1386259200, 1386262800, 1386266400, 1386270000, 1386273600, 
    1386277200, 1386280800, 1386284400, 1386288000, 1386291600, 1386295200, 
    1386298800, 1386302400, 1386306000, 1386309600, 1386313200, 1386316800, 
    1386320400, 1386324000, 1386327600, 1386331200, 1386334800, 1386338400, 
    1386342000, 1386345600, 1386349200, 1386352800, 1386356400, 1386360000, 
    1386363600, 1386367200, 1386370800, 1386374400, 1386378000, 1386381600, 
    1386385200, 1386388800, 1386392400, 1386396000, 1386399600, 1386403200, 
    1386406800, 1386410400, 1386414000, 1386417600, 1386421200, 1386424800, 
    1386428400, 1386432000, 1386435600, 1386439200, 1386442800, 1386446400, 
    1386450000, 1386453600, 1386457200, 1386460800, 1386464400, 1386468000, 
    1386471600, 1386475200, 1386478800, 1386482400, 1386486000, 1386489600, 
    1386493200, 1386496800, 1386500400, 1386504000, 1386507600, 1386511200, 
    1386514800, 1386518400, 1386522000, 1386525600, 1386529200, 1386532800, 
    1386536400, 1386540000, 1386543600, 1386547200, 1386550800, 1386554400, 
    1386558000, 1386561600, 1386565200, 1386568800, 1386572400, 1386576000, 
    1386579600, 1386583200, 1386586800, 1386590400, 1386594000, 1386597600, 
    1386601200, 1386604800, 1386608400, 1386612000, 1386615600, 1386619200, 
    1386622800, 1386626400, 1386630000, 1386633600, 1386637200, 1386640800, 
    1386644400, 1386648000, 1386651600, 1386655200, 1386658800, 1386662400, 
    1386666000, 1386669600, 1386673200, 1386676800, 1386680400, 1386684000, 
    1386687600, 1386691200, 1386694800, 1386698400, 1386702000, 1386705600, 
    1386709200, 1386712800, 1386716400, 1386720000, 1386723600, 1386727200, 
    1386730800, 1386734400, 1386738000, 1386741600, 1386745200, 1386748800, 
    1386752400, 1386756000, 1386759600, 1386763200, 1386766800, 1386770400, 
    1386774000, 1386777600, 1386781200, 1386784800, 1386788400, 1386792000, 
    1386795600, 1386799200, 1386802800, 1386806400, 1386810000, 1386813600, 
    1386817200, 1386820800, 1386824400, 1386828000, 1386831600, 1386835200, 
    1386838800, 1386842400, 1386846000, 1386849600, 1386853200, 1386856800, 
    1386860400, 1386864000, 1386867600, 1386871200, 1386874800, 1386878400, 
    1386882000, 1386885600, 1386889200, 1386892800, 1386896400, 1386900000, 
    1386903600, 1386907200, 1386910800, 1386914400, 1386918000, 1386921600, 
    1386925200, 1386928800, 1386932400, 1386936000, 1386939600, 1386943200, 
    1386946800, 1386950400, 1386954000, 1386957600, 1386961200, 1386964800, 
    1386968400, 1386972000, 1386975600, 1386979200, 1386982800, 1386986400, 
    1386990000, 1386993600, 1386997200, 1387000800, 1387004400, 1387008000, 
    1387011600, 1387015200, 1387018800, 1387022400, 1387026000, 1387029600, 
    1387033200, 1387036800, 1387040400, 1387044000, 1387047600, 1387051200, 
    1387054800, 1387058400, 1387062000, 1387065600, 1387069200, 1387072800, 
    1387076400, 1387080000, 1387083600, 1387087200, 1387090800, 1387094400, 
    1387098000, 1387101600, 1387105200, 1387108800, 1387112400, 1387116000, 
    1387119600, 1387123200, 1387126800, 1387130400, 1387134000, 1387137600, 
    1387141200, 1387144800, 1387148400, 1387152000, 1387155600, 1387159200, 
    1387162800, 1387166400, 1387170000, 1387173600, 1387177200, 1387180800, 
    1387184400, 1387188000, 1387191600, 1387195200, 1387198800, 1387202400, 
    1387206000, 1387209600, 1387213200, 1387216800, 1387220400, 1387224000, 
    1387227600, 1387231200, 1387234800, 1387238400, 1387242000, 1387245600, 
    1387249200, 1387252800, 1387256400, 1387260000, 1387263600, 1387267200, 
    1387270800, 1387274400, 1387278000, 1387281600, 1387285200, 1387288800, 
    1387292400, 1387296000, 1387299600, 1387303200, 1387306800, 1387310400, 
    1387314000, 1387317600, 1387321200, 1387324800, 1387328400, 1387332000, 
    1387335600, 1387339200, 1387342800, 1387346400, 1387350000, 1387353600, 
    1387357200, 1387360800, 1387364400, 1387368000, 1387371600, 1387375200, 
    1387378800, 1387382400, 1387386000, 1387389600, 1387393200, 1387396800, 
    1387400400, 1387404000, 1387407600, 1387411200, 1387414800, 1387418400, 
    1387422000, 1387425600, 1387429200, 1387432800, 1387436400, 1387440000, 
    1387443600, 1387447200, 1387450800, 1387454400, 1387458000, 1387461600, 
    1387465200, 1387468800, 1387472400, 1387476000, 1387479600, 1387483200, 
    1387486800, 1387490400, 1387494000, 1387497600, 1387501200, 1387504800, 
    1387508400, 1387512000, 1387515600, 1387519200, 1387522800, 1387526400, 
    1387530000, 1387533600, 1387537200, 1387540800, 1387544400, 1387548000, 
    1387551600, 1387555200, 1387558800, 1387562400, 1387566000, 1387569600, 
    1387573200, 1387576800, 1387580400, 1387584000, 1387587600, 1387591200, 
    1387594800, 1387598400, 1387602000, 1387605600, 1387609200, 1387612800, 
    1387616400, 1387620000, 1387623600, 1387627200, 1387630800, 1387634400, 
    1387638000, 1387641600, 1387645200, 1387648800, 1387652400, 1387656000, 
    1387659600, 1387663200, 1387666800, 1387670400, 1387674000, 1387677600, 
    1387681200, 1387684800, 1387688400, 1387692000, 1387695600, 1387699200, 
    1387702800, 1387706400, 1387710000, 1387713600, 1387717200, 1387720800, 
    1387724400, 1387728000, 1387731600, 1387735200, 1387738800, 1387742400, 
    1387746000, 1387749600, 1387753200, 1387756800, 1387760400, 1387764000, 
    1387767600, 1387771200, 1387774800, 1387778400, 1387782000, 1387785600, 
    1387789200, 1387792800, 1387796400, 1387800000, 1387803600, 1387807200, 
    1387810800, 1387814400, 1387818000, 1387821600, 1387825200, 1387828800, 
    1387832400, 1387836000, 1387839600, 1387843200, 1387846800, 1387850400, 
    1387854000, 1387857600, 1387861200, 1387864800, 1387868400, 1387872000, 
    1387875600, 1387879200, 1387882800, 1387886400, 1387890000, 1387893600, 
    1387897200, 1387900800, 1387904400, 1387908000, 1387911600, 1387915200, 
    1387918800, 1387922400, 1387926000, 1387929600, 1387933200, 1387936800, 
    1387940400, 1387944000, 1387947600, 1387951200, 1387954800, 1387958400, 
    1387962000, 1387965600, 1387969200, 1387972800, 1387976400, 1387980000, 
    1387983600, 1387987200, 1387990800, 1387994400, 1387998000, 1388001600, 
    1388005200, 1388008800, 1388012400, 1388016000, 1388019600, 1388023200, 
    1388026800, 1388030400, 1388034000, 1388037600, 1388041200, 1388044800, 
    1388048400, 1388052000, 1388055600, 1388059200, 1388062800, 1388066400, 
    1388070000, 1388073600, 1388077200, 1388080800, 1388084400, 1388088000, 
    1388091600, 1388095200, 1388098800, 1388102400, 1388106000, 1388109600, 
    1388113200, 1388116800, 1388120400, 1388124000, 1388127600, 1388131200, 
    1388134800, 1388138400, 1388142000, 1388145600, 1388149200, 1388152800, 
    1388156400, 1388160000, 1388163600, 1388167200, 1388170800, 1388174400, 
    1388178000, 1388181600, 1388185200, 1388188800, 1388192400, 1388196000, 
    1388199600, 1388203200, 1388206800, 1388210400, 1388214000, 1388217600, 
    1388221200, 1388224800, 1388228400, 1388232000, 1388235600, 1388239200, 
    1388242800, 1388246400, 1388250000, 1388253600, 1388257200, 1388260800, 
    1388264400, 1388268000, 1388271600, 1388275200, 1388278800, 1388282400, 
    1388286000, 1388289600, 1388293200, 1388296800, 1388300400, 1388304000, 
    1388307600, 1388311200, 1388314800, 1388318400, 1388322000, 1388325600, 
    1388329200, 1388332800, 1388336400, 1388340000, 1388343600, 1388347200, 
    1388350800, 1388354400, 1388358000, 1388361600, 1388365200, 1388368800, 
    1388372400, 1388376000, 1388379600, 1388383200, 1388386800, 1388390400, 
    1388394000, 1388397600, 1388401200, 1388404800, 1388408400, 1388412000, 
    1388415600, 1388419200, 1388422800, 1388426400, 1388430000, 1388433600, 
    1388437200, 1388440800, 1388444400, 1388448000, 1388451600, 1388455200, 
    1388458800, 1388462400, 1388466000, 1388469600, 1388473200, 1388476800, 
    1388480400, 1388484000, 1388487600, 1388491200, 1388494800, 1388498400, 
    1388502000, 1388505600, 1388509200, 1388512800, 1388516400, 1388520000, 
    1388523600, 1388527200, 1388530800, 1388534400, 1388538000, 1388541600, 
    1388545200, 1388548800, 1388552400, 1388556000, 1388559600, 1388563200, 
    1388566800, 1388570400, 1388574000, 1388577600, 1388581200, 1388584800, 
    1388588400, 1388592000, 1388595600, 1388599200, 1388602800, 1388606400, 
    1388610000, 1388613600, 1388617200, 1388620800, 1388624400, 1388628000, 
    1388631600, 1388635200, 1388638800, 1388642400, 1388646000, 1388649600, 
    1388653200, 1388656800, 1388660400, 1388664000, 1388667600, 1388671200, 
    1388674800, 1388678400, 1388682000, 1388685600, 1388689200, 1388692800, 
    1388696400, 1388700000, 1388703600, 1388707200, 1388710800, 1388714400, 
    1388718000, 1388721600, 1388725200, 1388728800, 1388732400, 1388736000, 
    1388739600, 1388743200, 1388746800, 1388750400, 1388754000, 1388757600, 
    1388761200, 1388764800, 1388768400, 1388772000, 1388775600, 1388779200, 
    1388782800, 1388786400, 1388790000, 1388793600, 1388797200, 1388800800, 
    1388804400, 1388808000, 1388811600, 1388815200, 1388818800, 1388822400, 
    1388826000, 1388829600, 1388833200, 1388836800, 1388840400, 1388844000, 
    1388847600, 1388851200, 1388854800, 1388858400, 1388862000, 1388865600, 
    1388869200, 1388872800, 1388876400, 1388880000, 1388883600, 1388887200, 
    1388890800, 1388894400, 1388898000, 1388901600, 1388905200, 1388908800, 
    1388912400, 1388916000, 1388919600, 1388923200, 1388926800, 1388930400, 
    1388934000, 1388937600, 1388941200, 1388944800, 1388948400, 1388952000, 
    1388955600, 1388959200, 1388962800, 1388966400, 1388970000, 1388973600, 
    1388977200, 1388980800, 1388984400, 1388988000, 1388991600, 1388995200, 
    1388998800, 1389002400, 1389006000, 1389009600, 1389013200, 1389016800, 
    1389020400, 1389024000, 1389027600, 1389031200, 1389034800, 1389038400, 
    1389042000, 1389045600, 1389049200, 1389052800, 1389056400, 1389060000, 
    1389063600, 1389067200, 1389070800, 1389074400, 1389078000, 1389081600, 
    1389085200, 1389088800, 1389092400, 1389096000, 1389099600, 1389103200, 
    1389106800, 1389110400, 1389114000, 1389117600, 1389121200, 1389124800, 
    1389128400, 1389132000, 1389135600, 1389139200, 1389142800, 1389146400, 
    1389150000, 1389153600, 1389157200, 1389160800, 1389164400, 1389168000, 
    1389171600, 1389175200, 1389178800, 1389182400, 1389186000, 1389189600, 
    1389193200, 1389196800, 1389200400, 1389204000, 1389207600, 1389211200, 
    1389214800, 1389218400, 1389222000, 1389225600, 1389229200, 1389232800, 
    1389236400, 1389240000, 1389243600, 1389247200, 1389250800, 1389254400, 
    1389258000, 1389261600, 1389265200, 1389268800, 1389272400, 1389276000, 
    1389279600, 1389283200, 1389286800, 1389290400, 1389294000, 1389297600, 
    1389301200, 1389304800, 1389308400, 1389312000, 1389315600, 1389319200, 
    1389322800, 1389326400, 1389330000, 1389333600, 1389337200, 1389340800, 
    1389344400, 1389348000, 1389351600, 1389355200, 1389358800, 1389362400, 
    1389366000, 1389369600, 1389373200, 1389376800, 1389380400, 1389384000, 
    1389387600, 1389391200, 1389394800, 1389398400, 1389402000, 1389405600, 
    1389409200, 1389412800, 1389416400, 1389420000, 1389423600, 1389427200, 
    1389430800, 1389434400, 1389438000, 1389441600, 1389445200, 1389448800, 
    1389452400, 1389456000, 1389459600, 1389463200, 1389466800, 1389470400, 
    1389474000, 1389477600, 1389481200, 1389484800, 1389488400, 1389492000, 
    1389495600, 1389499200, 1389502800, 1389506400, 1389510000, 1389513600, 
    1389517200, 1389520800, 1389524400, 1389528000, 1389531600, 1389535200, 
    1389538800, 1389542400, 1389546000, 1389549600, 1389553200, 1389556800, 
    1389560400, 1389564000, 1389567600, 1389571200, 1389574800, 1389578400, 
    1389582000, 1389585600, 1389589200, 1389592800, 1389596400, 1389600000, 
    1389603600, 1389607200, 1389610800, 1389614400, 1389618000, 1389621600, 
    1389625200, 1389628800, 1389632400, 1389636000, 1389639600, 1389643200, 
    1389646800, 1389650400, 1389654000, 1389657600, 1389661200, 1389664800, 
    1389668400, 1389672000, 1389675600, 1389679200, 1389682800, 1389686400, 
    1389690000, 1389693600, 1389697200, 1389700800, 1389704400, 1389708000, 
    1389711600, 1389715200, 1389718800, 1389722400, 1389726000, 1389729600, 
    1389733200, 1389736800, 1389740400, 1389744000, 1389747600, 1389751200, 
    1389754800, 1389758400, 1389762000, 1389765600, 1389769200, 1389772800, 
    1389776400, 1389780000, 1389783600, 1389787200, 1389790800, 1389794400, 
    1389798000, 1389801600, 1389805200, 1389808800, 1389812400, 1389816000, 
    1389819600, 1389823200, 1389826800, 1389830400, 1389834000, 1389837600, 
    1389841200, 1389844800, 1389848400, 1389852000, 1389855600, 1389859200, 
    1389862800, 1389866400, 1389870000, 1389873600, 1389877200, 1389880800, 
    1389884400, 1389888000, 1389891600, 1389895200, 1389898800, 1389902400, 
    1389906000, 1389909600, 1389913200, 1389916800, 1389920400, 1389924000, 
    1389927600, 1389931200, 1389934800, 1389938400, 1389942000, 1389945600, 
    1389949200, 1389952800, 1389956400, 1389960000, 1389963600, 1389967200, 
    1389970800, 1389974400, 1389978000, 1389981600, 1389985200, 1389988800, 
    1389992400, 1389996000, 1389999600, 1390003200, 1390006800, 1390010400, 
    1390014000, 1390017600, 1390021200, 1390024800, 1390028400, 1390032000, 
    1390035600, 1390039200, 1390042800, 1390046400, 1390050000, 1390053600, 
    1390057200, 1390060800, 1390064400, 1390068000, 1390071600, 1390075200, 
    1390078800, 1390082400, 1390086000, 1390089600, 1390093200, 1390096800, 
    1390100400, 1390104000, 1390107600, 1390111200, 1390114800, 1390118400, 
    1390122000, 1390125600, 1390129200, 1390132800, 1390136400, 1390140000, 
    1390143600, 1390147200, 1390150800, 1390154400, 1390158000, 1390161600, 
    1390165200, 1390168800, 1390172400, 1390176000, 1390179600, 1390183200, 
    1390186800, 1390190400, 1390194000, 1390197600, 1390201200, 1390204800, 
    1390208400, 1390212000, 1390215600, 1390219200, 1390222800, 1390226400, 
    1390230000, 1390233600, 1390237200, 1390240800, 1390244400, 1390248000, 
    1390251600, 1390255200, 1390258800, 1390262400, 1390266000, 1390269600, 
    1390273200, 1390276800, 1390280400, 1390284000, 1390287600, 1390291200, 
    1390294800, 1390298400, 1390302000, 1390305600, 1390309200, 1390312800, 
    1390316400, 1390320000, 1390323600, 1390327200, 1390330800, 1390334400, 
    1390338000, 1390341600, 1390345200, 1390348800, 1390352400, 1390356000, 
    1390359600, 1390363200, 1390366800, 1390370400, 1390374000, 1390377600, 
    1390381200, 1390384800, 1390388400, 1390392000, 1390395600, 1390399200, 
    1390402800, 1390406400, 1390410000, 1390413600, 1390417200, 1390420800, 
    1390424400, 1390428000, 1390431600, 1390435200, 1390438800, 1390442400, 
    1390446000, 1390449600, 1390453200, 1390456800, 1390460400, 1390464000, 
    1390467600, 1390471200, 1390474800, 1390478400, 1390482000, 1390485600, 
    1390489200, 1390492800, 1390496400, 1390500000, 1390503600, 1390507200, 
    1390510800, 1390514400, 1390518000, 1390521600, 1390525200, 1390528800, 
    1390532400, 1390536000, 1390539600, 1390543200, 1390546800, 1390550400, 
    1390554000, 1390557600, 1390561200, 1390564800, 1390568400, 1390572000, 
    1390575600, 1390579200, 1390582800, 1390586400, 1390590000, 1390593600, 
    1390597200, 1390600800, 1390604400, 1390608000, 1390611600, 1390615200, 
    1390618800, 1390622400, 1390626000, 1390629600, 1390633200, 1390636800, 
    1390640400, 1390644000, 1390647600, 1390651200, 1390654800, 1390658400, 
    1390662000, 1390665600, 1390669200, 1390672800, 1390676400, 1390680000, 
    1390683600, 1390687200, 1390690800, 1390694400, 1390698000, 1390701600, 
    1390705200, 1390708800, 1390712400, 1390716000, 1390719600, 1390723200, 
    1390726800, 1390730400, 1390734000, 1390737600, 1390741200, 1390744800, 
    1390748400, 1390752000, 1390755600, 1390759200, 1390762800, 1390766400, 
    1390770000, 1390773600, 1390777200, 1390780800, 1390784400, 1390788000, 
    1390791600, 1390795200, 1390798800, 1390802400, 1390806000, 1390809600, 
    1390813200, 1390816800, 1390820400, 1390824000, 1390827600, 1390831200, 
    1390834800, 1390838400, 1390842000, 1390845600, 1390849200, 1390852800, 
    1390856400, 1390860000, 1390863600, 1390867200, 1390870800, 1390874400, 
    1390878000, 1390881600, 1390885200, 1390888800, 1390892400, 1390896000, 
    1390899600, 1390903200, 1390906800, 1390910400, 1390914000, 1390917600, 
    1390921200, 1390924800, 1390928400, 1390932000, 1390935600, 1390939200, 
    1390942800, 1390946400, 1390950000, 1390953600, 1390957200, 1390960800, 
    1390964400, 1390968000, 1390971600, 1390975200, 1390978800, 1390982400, 
    1390986000, 1390989600, 1390993200, 1390996800, 1391000400, 1391004000, 
    1391007600, 1391011200, 1391014800, 1391018400, 1391022000, 1391025600, 
    1391029200, 1391032800, 1391036400, 1391040000, 1391043600, 1391047200, 
    1391050800, 1391054400, 1391058000, 1391061600, 1391065200, 1391068800, 
    1391072400, 1391076000, 1391079600, 1391083200, 1391086800, 1391090400, 
    1391094000, 1391097600, 1391101200, 1391104800, 1391108400, 1391112000, 
    1391115600, 1391119200, 1391122800, 1391126400, 1391130000, 1391133600, 
    1391137200, 1391140800, 1391144400, 1391148000, 1391151600, 1391155200, 
    1391158800, 1391162400, 1391166000, 1391169600, 1391173200, 1391176800, 
    1391180400, 1391184000, 1391187600, 1391191200, 1391194800, 1391198400, 
    1391202000, 1391205600, 1391209200, 1391212800, 1391216400, 1391220000, 
    1391223600, 1391227200, 1391230800, 1391234400, 1391238000, 1391241600, 
    1391245200, 1391248800, 1391252400, 1391256000, 1391259600, 1391263200, 
    1391266800, 1391270400, 1391274000, 1391277600, 1391281200, 1391284800, 
    1391288400, 1391292000, 1391295600, 1391299200, 1391302800, 1391306400, 
    1391310000, 1391313600, 1391317200, 1391320800, 1391324400, 1391328000, 
    1391331600, 1391335200, 1391338800, 1391342400, 1391346000, 1391349600, 
    1391353200, 1391356800, 1391360400, 1391364000, 1391367600, 1391371200, 
    1391374800, 1391378400, 1391382000, 1391385600, 1391389200, 1391392800, 
    1391396400, 1391400000, 1391403600, 1391407200, 1391410800, 1391414400, 
    1391418000, 1391421600, 1391425200, 1391428800, 1391432400, 1391436000, 
    1391439600, 1391443200, 1391446800, 1391450400, 1391454000, 1391457600, 
    1391461200, 1391464800, 1391468400, 1391472000, 1391475600, 1391479200, 
    1391482800, 1391486400, 1391490000, 1391493600, 1391497200, 1391500800, 
    1391504400, 1391508000, 1391511600, 1391515200, 1391518800, 1391522400, 
    1391526000, 1391529600, 1391533200, 1391536800, 1391540400, 1391544000, 
    1391547600, 1391551200, 1391554800, 1391558400, 1391562000, 1391565600, 
    1391569200, 1391572800, 1391576400, 1391580000, 1391583600, 1391587200, 
    1391590800, 1391594400, 1391598000, 1391601600, 1391605200, 1391608800, 
    1391612400, 1391616000, 1391619600, 1391623200, 1391626800, 1391630400, 
    1391634000, 1391637600, 1391641200, 1391644800, 1391648400, 1391652000, 
    1391655600, 1391659200, 1391662800, 1391666400, 1391670000, 1391673600, 
    1391677200, 1391680800, 1391684400, 1391688000, 1391691600, 1391695200, 
    1391698800, 1391702400, 1391706000, 1391709600, 1391713200, 1391716800, 
    1391720400, 1391724000, 1391727600, 1391731200, 1391734800, 1391738400, 
    1391742000, 1391745600, 1391749200, 1391752800, 1391756400, 1391760000, 
    1391763600, 1391767200, 1391770800, 1391774400, 1391778000, 1391781600, 
    1391785200, 1391788800, 1391792400, 1391796000, 1391799600, 1391803200, 
    1391806800, 1391810400, 1391814000, 1391817600, 1391821200, 1391824800, 
    1391828400, 1391832000, 1391835600, 1391839200, 1391842800, 1391846400, 
    1391850000, 1391853600, 1391857200, 1391860800, 1391864400, 1391868000, 
    1391871600, 1391875200, 1391878800, 1391882400, 1391886000, 1391889600, 
    1391893200, 1391896800, 1391900400, 1391904000, 1391907600, 1391911200, 
    1391914800, 1391918400, 1391922000, 1391925600, 1391929200, 1391932800, 
    1391936400, 1391940000, 1391943600, 1391947200, 1391950800, 1391954400, 
    1391958000, 1391961600, 1391965200, 1391968800, 1391972400, 1391976000, 
    1391979600, 1391983200, 1391986800, 1391990400, 1391994000, 1391997600, 
    1392001200, 1392004800, 1392008400, 1392012000, 1392015600, 1392019200, 
    1392022800, 1392026400, 1392030000, 1392033600, 1392037200, 1392040800, 
    1392044400, 1392048000, 1392051600, 1392055200, 1392058800, 1392062400, 
    1392066000, 1392069600, 1392073200, 1392076800, 1392080400, 1392084000, 
    1392087600, 1392091200, 1392094800, 1392098400, 1392102000, 1392105600, 
    1392109200, 1392112800, 1392116400, 1392120000, 1392123600, 1392127200, 
    1392130800, 1392134400, 1392138000, 1392141600, 1392145200, 1392148800, 
    1392152400, 1392156000, 1392159600, 1392163200, 1392166800, 1392170400, 
    1392174000, 1392177600, 1392181200, 1392184800, 1392188400, 1392192000, 
    1392195600, 1392199200, 1392202800, 1392206400, 1392210000, 1392213600, 
    1392217200, 1392220800, 1392224400, 1392228000, 1392231600, 1392235200, 
    1392238800, 1392242400, 1392246000, 1392249600, 1392253200, 1392256800, 
    1392260400, 1392264000, 1392267600, 1392271200, 1392274800, 1392278400, 
    1392282000, 1392285600, 1392289200, 1392292800, 1392296400, 1392300000, 
    1392303600, 1392307200, 1392310800, 1392314400, 1392318000, 1392321600, 
    1392325200, 1392328800, 1392332400, 1392336000, 1392339600, 1392343200, 
    1392346800, 1392350400, 1392354000, 1392357600, 1392361200, 1392364800, 
    1392368400, 1392372000, 1392375600, 1392379200, 1392382800, 1392386400, 
    1392390000, 1392393600, 1392397200, 1392400800, 1392404400, 1392408000, 
    1392411600, 1392415200, 1392418800, 1392422400, 1392426000, 1392429600, 
    1392433200, 1392436800, 1392440400, 1392444000, 1392447600, 1392451200, 
    1392454800, 1392458400, 1392462000, 1392465600, 1392469200, 1392472800, 
    1392476400, 1392480000, 1392483600, 1392487200, 1392490800, 1392494400, 
    1392498000, 1392501600, 1392505200, 1392508800, 1392512400, 1392516000, 
    1392519600, 1392523200, 1392526800, 1392530400, 1392534000, 1392537600, 
    1392541200, 1392544800, 1392548400, 1392552000, 1392555600, 1392559200, 
    1392562800, 1392566400, 1392570000, 1392573600, 1392577200, 1392580800, 
    1392584400, 1392588000, 1392591600, 1392595200, 1392598800, 1392602400, 
    1392606000, 1392609600, 1392613200, 1392616800, 1392620400, 1392624000, 
    1392627600, 1392631200, 1392634800, 1392638400, 1392642000, 1392645600, 
    1392649200, 1392652800, 1392656400, 1392660000, 1392663600, 1392667200, 
    1392670800, 1392674400, 1392678000, 1392681600, 1392685200, 1392688800, 
    1392692400, 1392696000, 1392699600, 1392703200, 1392706800, 1392710400, 
    1392714000, 1392717600, 1392721200, 1392724800, 1392728400, 1392732000, 
    1392735600, 1392739200, 1392742800, 1392746400, 1392750000, 1392753600, 
    1392757200, 1392760800, 1392764400, 1392768000, 1392771600, 1392775200, 
    1392778800, 1392782400, 1392786000, 1392789600, 1392793200, 1392796800, 
    1392800400, 1392804000, 1392807600, 1392811200, 1392814800, 1392818400, 
    1392822000, 1392825600, 1392829200, 1392832800, 1392836400, 1392840000, 
    1392843600, 1392847200, 1392850800, 1392854400, 1392858000, 1392861600, 
    1392865200, 1392868800, 1392872400, 1392876000, 1392879600, 1392883200, 
    1392886800, 1392890400, 1392894000, 1392897600, 1392901200, 1392904800, 
    1392908400, 1392912000, 1392915600, 1392919200, 1392922800, 1392926400, 
    1392930000, 1392933600, 1392937200, 1392940800, 1392944400, 1392948000, 
    1392951600, 1392955200, 1392958800, 1392962400, 1392966000, 1392969600, 
    1392973200, 1392976800, 1392980400, 1392984000, 1392987600, 1392991200, 
    1392994800, 1392998400, 1393002000, 1393005600, 1393009200, 1393012800, 
    1393016400, 1393020000, 1393023600, 1393027200, 1393030800, 1393034400, 
    1393038000, 1393041600, 1393045200, 1393048800, 1393052400, 1393056000, 
    1393059600, 1393063200, 1393066800, 1393070400, 1393074000, 1393077600, 
    1393081200, 1393084800, 1393088400, 1393092000, 1393095600, 1393099200, 
    1393102800, 1393106400, 1393110000, 1393113600, 1393117200, 1393120800, 
    1393124400, 1393128000, 1393131600, 1393135200, 1393138800, 1393142400, 
    1393146000, 1393149600, 1393153200, 1393156800, 1393160400, 1393164000, 
    1393167600, 1393171200, 1393174800, 1393178400, 1393182000, 1393185600, 
    1393189200, 1393192800, 1393196400, 1393200000, 1393203600, 1393207200, 
    1393210800, 1393214400, 1393218000, 1393221600, 1393225200, 1393228800, 
    1393232400, 1393236000, 1393239600, 1393243200, 1393246800, 1393250400, 
    1393254000, 1393257600, 1393261200, 1393264800, 1393268400, 1393272000, 
    1393275600, 1393279200, 1393282800, 1393286400, 1393290000, 1393293600, 
    1393297200, 1393300800, 1393304400, 1393308000, 1393311600, 1393315200, 
    1393318800, 1393322400, 1393326000, 1393329600, 1393333200, 1393336800, 
    1393340400, 1393344000, 1393347600, 1393351200, 1393354800, 1393358400, 
    1393362000, 1393365600, 1393369200, 1393372800, 1393376400, 1393380000, 
    1393383600, 1393387200, 1393390800, 1393394400, 1393398000, 1393401600, 
    1393405200, 1393408800, 1393412400, 1393416000, 1393419600, 1393423200, 
    1393426800, 1393430400, 1393434000, 1393437600, 1393441200, 1393444800, 
    1393448400, 1393452000, 1393455600, 1393459200, 1393462800, 1393466400, 
    1393470000, 1393473600, 1393477200, 1393480800, 1393484400, 1393488000, 
    1393491600, 1393495200, 1393498800, 1393502400, 1393506000, 1393509600, 
    1393513200, 1393516800, 1393520400, 1393524000, 1393527600, 1393531200, 
    1393534800, 1393538400, 1393542000, 1393545600, 1393549200, 1393552800, 
    1393556400, 1393560000, 1393563600, 1393567200, 1393570800, 1393574400, 
    1393578000, 1393581600, 1393585200, 1393588800, 1393592400, 1393596000, 
    1393599600, 1393603200, 1393606800, 1393610400, 1393614000, 1393617600, 
    1393621200, 1393624800, 1393628400, 1393632000, 1393635600, 1393639200, 
    1393642800, 1393646400, 1393650000, 1393653600, 1393657200, 1393660800, 
    1393664400, 1393668000, 1393671600, 1393675200, 1393678800, 1393682400, 
    1393686000, 1393689600, 1393693200, 1393696800, 1393700400, 1393704000, 
    1393707600, 1393711200, 1393714800, 1393718400, 1393722000, 1393725600, 
    1393729200, 1393732800, 1393736400, 1393740000, 1393743600, 1393747200, 
    1393750800, 1393754400, 1393758000, 1393761600, 1393765200, 1393768800, 
    1393772400, 1393776000, 1393779600, 1393783200, 1393786800, 1393790400, 
    1393794000, 1393797600, 1393801200, 1393804800, 1393808400, 1393812000, 
    1393815600, 1393819200, 1393822800, 1393826400, 1393830000, 1393833600, 
    1393837200, 1393840800, 1393844400, 1393848000, 1393851600, 1393855200, 
    1393858800, 1393862400, 1393866000, 1393869600, 1393873200, 1393876800, 
    1393880400, 1393884000, 1393887600, 1393891200, 1393894800, 1393898400, 
    1393902000, 1393905600, 1393909200, 1393912800, 1393916400, 1393920000, 
    1393923600, 1393927200, 1393930800, 1393934400, 1393938000, 1393941600, 
    1393945200, 1393948800, 1393952400, 1393956000, 1393959600, 1393963200, 
    1393966800, 1393970400, 1393974000, 1393977600, 1393981200, 1393984800, 
    1393988400, 1393992000, 1393995600, 1393999200, 1394002800, 1394006400, 
    1394010000, 1394013600, 1394017200, 1394020800, 1394024400, 1394028000, 
    1394031600, 1394035200, 1394038800, 1394042400, 1394046000, 1394049600, 
    1394053200, 1394056800, 1394060400, 1394064000, 1394067600, 1394071200, 
    1394074800, 1394078400, 1394082000, 1394085600, 1394089200, 1394092800, 
    1394096400, 1394100000, 1394103600, 1394107200, 1394110800, 1394114400, 
    1394118000, 1394121600, 1394125200, 1394128800, 1394132400, 1394136000, 
    1394139600, 1394143200, 1394146800, 1394150400, 1394154000, 1394157600, 
    1394161200, 1394164800, 1394168400, 1394172000, 1394175600, 1394179200, 
    1394182800, 1394186400, 1394190000, 1394193600, 1394197200, 1394200800, 
    1394204400, 1394208000, 1394211600, 1394215200, 1394218800, 1394222400, 
    1394226000, 1394229600, 1394233200, 1394236800, 1394240400, 1394244000, 
    1394247600, 1394251200, 1394254800, 1394258400, 1394262000, 1394265600, 
    1394269200, 1394272800, 1394276400, 1394280000, 1394283600, 1394287200, 
    1394290800, 1394294400, 1394298000, 1394301600, 1394305200, 1394308800, 
    1394312400, 1394316000, 1394319600, 1394323200, 1394326800, 1394330400, 
    1394334000, 1394337600, 1394341200, 1394344800, 1394348400, 1394352000, 
    1394355600, 1394359200, 1394362800, 1394366400, 1394370000, 1394373600, 
    1394377200, 1394380800, 1394384400, 1394388000, 1394391600, 1394395200, 
    1394398800, 1394402400, 1394406000, 1394409600, 1394413200, 1394416800, 
    1394420400, 1394424000, 1394427600, 1394431200, 1394434800, 1394438400, 
    1394442000, 1394445600, 1394449200, 1394452800, 1394456400, 1394460000, 
    1394463600, 1394467200, 1394470800, 1394474400, 1394478000, 1394481600, 
    1394485200, 1394488800, 1394492400, 1394496000, 1394499600, 1394503200, 
    1394506800, 1394510400, 1394514000, 1394517600, 1394521200, 1394524800, 
    1394528400, 1394532000, 1394535600, 1394539200, 1394542800, 1394546400, 
    1394550000, 1394553600, 1394557200, 1394560800, 1394564400, 1394568000, 
    1394571600, 1394575200, 1394578800, 1394582400, 1394586000, 1394589600, 
    1394593200, 1394596800, 1394600400, 1394604000, 1394607600, 1394611200, 
    1394614800, 1394618400, 1394622000, 1394625600, 1394629200, 1394632800, 
    1394636400, 1394640000, 1394643600, 1394647200, 1394650800, 1394654400, 
    1394658000, 1394661600, 1394665200, 1394668800, 1394672400, 1394676000, 
    1394679600, 1394683200, 1394686800, 1394690400, 1394694000, 1394697600, 
    1394701200, 1394704800, 1394708400, 1394712000, 1394715600, 1394719200, 
    1394722800, 1394726400, 1394730000, 1394733600, 1394737200, 1394740800, 
    1394744400, 1394748000, 1394751600, 1394755200, 1394758800, 1394762400, 
    1394766000, 1394769600, 1394773200, 1394776800, 1394780400, 1394784000, 
    1394787600, 1394791200, 1394794800, 1394798400, 1394802000, 1394805600, 
    1394809200, 1394812800, 1394816400, 1394820000, 1394823600, 1394827200, 
    1394830800, 1394834400, 1394838000, 1394841600, 1394845200, 1394848800, 
    1394852400, 1394856000, 1394859600, 1394863200, 1394866800, 1394870400, 
    1394874000, 1394877600, 1394881200, 1394884800, 1394888400, 1394892000, 
    1394895600, 1394899200, 1394902800, 1394906400, 1394910000, 1394913600, 
    1394917200, 1394920800, 1394924400, 1394928000, 1394931600, 1394935200, 
    1394938800, 1394942400, 1394946000, 1394949600, 1394953200, 1394956800, 
    1394960400, 1394964000, 1394967600, 1394971200, 1394974800, 1394978400, 
    1394982000, 1394985600, 1394989200, 1394992800, 1394996400, 1395000000, 
    1395003600, 1395007200, 1395010800, 1395014400, 1395018000, 1395021600, 
    1395025200, 1395028800, 1395032400, 1395036000, 1395039600, 1395043200, 
    1395046800, 1395050400, 1395054000, 1395057600, 1395061200, 1395064800, 
    1395068400, 1395072000, 1395075600, 1395079200, 1395082800, 1395086400, 
    1395090000, 1395093600, 1395097200, 1395100800, 1395104400, 1395108000, 
    1395111600, 1395115200, 1395118800, 1395122400, 1395126000, 1395129600, 
    1395133200, 1395136800, 1395140400, 1395144000, 1395147600, 1395151200, 
    1395154800, 1395158400, 1395162000, 1395165600, 1395169200, 1395172800, 
    1395176400, 1395180000, 1395183600, 1395187200, 1395190800, 1395194400, 
    1395198000, 1395201600, 1395205200, 1395208800, 1395212400, 1395216000, 
    1395219600, 1395223200, 1395226800, 1395230400, 1395234000, 1395237600, 
    1395241200, 1395244800, 1395248400, 1395252000, 1395255600, 1395259200, 
    1395262800, 1395266400, 1395270000, 1395273600, 1395277200, 1395280800, 
    1395284400, 1395288000, 1395291600, 1395295200, 1395298800, 1395302400, 
    1395306000, 1395309600, 1395313200, 1395316800, 1395320400, 1395324000, 
    1395327600, 1395331200, 1395334800, 1395338400, 1395342000, 1395345600, 
    1395349200, 1395352800, 1395356400, 1395360000, 1395363600, 1395367200, 
    1395370800, 1395374400, 1395378000, 1395381600, 1395385200, 1395388800, 
    1395392400, 1395396000, 1395399600, 1395403200, 1395406800, 1395410400, 
    1395414000, 1395417600, 1395421200, 1395424800, 1395428400, 1395432000, 
    1395435600, 1395439200, 1395442800, 1395446400, 1395450000, 1395453600, 
    1395457200, 1395460800, 1395464400, 1395468000, 1395471600, 1395475200, 
    1395478800, 1395482400, 1395486000, 1395489600, 1395493200, 1395496800, 
    1395500400, 1395504000, 1395507600, 1395511200, 1395514800, 1395518400, 
    1395522000, 1395525600, 1395529200, 1395532800, 1395536400, 1395540000, 
    1395543600, 1395547200, 1395550800, 1395554400, 1395558000, 1395561600, 
    1395565200, 1395568800, 1395572400, 1395576000, 1395579600, 1395583200, 
    1395586800, 1395590400, 1395594000, 1395597600, 1395601200, 1395604800, 
    1395608400, 1395612000, 1395615600, 1395619200, 1395622800, 1395626400, 
    1395630000, 1395633600, 1395637200, 1395640800, 1395644400, 1395648000, 
    1395651600, 1395655200, 1395658800, 1395662400, 1395666000, 1395669600, 
    1395673200, 1395676800, 1395680400, 1395684000, 1395687600, 1395691200, 
    1395694800, 1395698400, 1395702000, 1395705600, 1395709200, 1395712800, 
    1395716400, 1395720000, 1395723600, 1395727200, 1395730800, 1395734400, 
    1395738000, 1395741600, 1395745200, 1395748800, 1395752400, 1395756000, 
    1395759600, 1395763200, 1395766800, 1395770400, 1395774000, 1395777600, 
    1395781200, 1395784800, 1395788400, 1395792000, 1395795600, 1395799200, 
    1395802800, 1395806400, 1395810000, 1395813600, 1395817200, 1395820800, 
    1395824400, 1395828000, 1395831600, 1395835200, 1395838800, 1395842400, 
    1395846000, 1395849600, 1395853200, 1395856800, 1395860400, 1395864000, 
    1395867600, 1395871200, 1395874800, 1395878400, 1395882000, 1395885600, 
    1395889200, 1395892800, 1395896400, 1395900000, 1395903600, 1395907200, 
    1395910800, 1395914400, 1395918000, 1395921600, 1395925200, 1395928800, 
    1395932400, 1395936000, 1395939600, 1395943200, 1395946800, 1395950400, 
    1395954000, 1395957600, 1395961200, 1395964800, 1395968400, 1395972000, 
    1395975600, 1395979200, 1395982800, 1395986400, 1395990000, 1395993600, 
    1395997200, 1396000800, 1396004400, 1396008000, 1396011600, 1396015200, 
    1396018800, 1396022400, 1396026000, 1396029600, 1396033200, 1396036800, 
    1396040400, 1396044000, 1396047600, 1396051200, 1396054800, 1396058400, 
    1396062000, 1396065600, 1396069200, 1396072800, 1396076400, 1396080000, 
    1396083600, 1396087200, 1396090800, 1396094400, 1396098000, 1396101600, 
    1396105200, 1396108800, 1396112400, 1396116000, 1396119600, 1396123200, 
    1396126800, 1396130400, 1396134000, 1396137600, 1396141200, 1396144800, 
    1396148400, 1396152000, 1396155600, 1396159200, 1396162800, 1396166400, 
    1396170000, 1396173600, 1396177200, 1396180800, 1396184400, 1396188000, 
    1396191600, 1396195200, 1396198800, 1396202400, 1396206000, 1396209600, 
    1396213200, 1396216800, 1396220400, 1396224000, 1396227600, 1396231200, 
    1396234800, 1396238400, 1396242000, 1396245600, 1396249200, 1396252800, 
    1396256400, 1396260000, 1396263600, 1396267200, 1396270800, 1396274400, 
    1396278000, 1396281600, 1396285200, 1396288800, 1396292400, 1396296000, 
    1396299600, 1396303200, 1396306800, 1396310400, 1396314000, 1396317600, 
    1396321200, 1396324800, 1396328400, 1396332000, 1396335600, 1396339200, 
    1396342800, 1396346400, 1396350000, 1396353600, 1396357200, 1396360800, 
    1396364400, 1396368000, 1396371600, 1396375200, 1396378800, 1396382400, 
    1396386000, 1396389600, 1396393200, 1396396800, 1396400400, 1396404000, 
    1396407600, 1396411200, 1396414800, 1396418400, 1396422000, 1396425600, 
    1396429200, 1396432800, 1396436400, 1396440000, 1396443600, 1396447200, 
    1396450800, 1396454400, 1396458000, 1396461600, 1396465200, 1396468800, 
    1396472400, 1396476000, 1396479600, 1396483200, 1396486800, 1396490400, 
    1396494000, 1396497600, 1396501200, 1396504800, 1396508400, 1396512000, 
    1396515600, 1396519200, 1396522800, 1396526400, 1396530000, 1396533600, 
    1396537200, 1396540800, 1396544400, 1396548000, 1396551600, 1396555200, 
    1396558800, 1396562400, 1396566000, 1396569600, 1396573200, 1396576800, 
    1396580400, 1396584000, 1396587600, 1396591200, 1396594800, 1396598400, 
    1396602000, 1396605600, 1396609200, 1396612800, 1396616400, 1396620000, 
    1396623600, 1396627200, 1396630800, 1396634400, 1396638000, 1396641600, 
    1396645200, 1396648800, 1396652400, 1396656000, 1396659600, 1396663200, 
    1396666800, 1396670400, 1396674000, 1396677600, 1396681200, 1396684800, 
    1396688400, 1396692000, 1396695600, 1396699200, 1396702800, 1396706400, 
    1396710000, 1396713600, 1396717200, 1396720800, 1396724400, 1396728000, 
    1396731600, 1396735200, 1396738800, 1396742400, 1396746000, 1396749600, 
    1396753200, 1396756800, 1396760400, 1396764000, 1396767600, 1396771200, 
    1396774800, 1396778400, 1396782000, 1396785600, 1396789200, 1396792800, 
    1396796400, 1396800000, 1396803600, 1396807200, 1396810800, 1396814400, 
    1396818000, 1396821600, 1396825200, 1396828800, 1396832400, 1396836000, 
    1396839600, 1396843200, 1396846800, 1396850400, 1396854000, 1396857600, 
    1396861200, 1396864800, 1396868400, 1396872000, 1396875600, 1396879200, 
    1396882800, 1396886400, 1396890000, 1396893600, 1396897200, 1396900800, 
    1396904400, 1396908000, 1396911600, 1396915200, 1396918800, 1396922400, 
    1396926000, 1396929600, 1396933200, 1396936800, 1396940400, 1396944000, 
    1396947600, 1396951200, 1396954800, 1396958400, 1396962000, 1396965600, 
    1396969200, 1396972800, 1396976400, 1396980000, 1396983600, 1396987200, 
    1396990800, 1396994400, 1396998000, 1397001600, 1397005200, 1397008800, 
    1397012400, 1397016000, 1397019600, 1397023200, 1397026800, 1397030400, 
    1397034000, 1397037600, 1397041200, 1397044800, 1397048400, 1397052000, 
    1397055600, 1397059200, 1397062800, 1397066400, 1397070000, 1397073600, 
    1397077200, 1397080800, 1397084400, 1397088000, 1397091600, 1397095200, 
    1397098800, 1397102400, 1397106000, 1397109600, 1397113200, 1397116800, 
    1397120400, 1397124000, 1397127600, 1397131200, 1397134800, 1397138400, 
    1397142000, 1397145600, 1397149200, 1397152800, 1397156400, 1397160000, 
    1397163600, 1397167200, 1397170800, 1397174400, 1397178000, 1397181600, 
    1397185200, 1397188800, 1397192400, 1397196000, 1397199600, 1397203200, 
    1397206800, 1397210400, 1397214000, 1397217600, 1397221200, 1397224800, 
    1397228400, 1397232000, 1397235600, 1397239200, 1397242800, 1397246400, 
    1397250000, 1397253600, 1397257200, 1397260800, 1397264400, 1397268000, 
    1397271600, 1397275200, 1397278800, 1397282400, 1397286000, 1397289600, 
    1397293200, 1397296800, 1397300400, 1397304000, 1397307600, 1397311200, 
    1397314800, 1397318400, 1397322000, 1397325600, 1397329200, 1397332800, 
    1397336400, 1397340000, 1397343600, 1397347200, 1397350800, 1397354400, 
    1397358000, 1397361600, 1397365200, 1397368800, 1397372400, 1397376000, 
    1397379600, 1397383200, 1397386800, 1397390400, 1397394000, 1397397600, 
    1397401200, 1397404800, 1397408400, 1397412000, 1397415600, 1397419200, 
    1397422800, 1397426400, 1397430000, 1397433600, 1397437200, 1397440800, 
    1397444400, 1397448000, 1397451600, 1397455200, 1397458800, 1397462400, 
    1397466000, 1397469600, 1397473200, 1397476800, 1397480400, 1397484000, 
    1397487600, 1397491200, 1397494800, 1397498400, 1397502000, 1397505600, 
    1397509200, 1397512800, 1397516400, 1397520000, 1397523600, 1397527200, 
    1397530800, 1397534400, 1397538000, 1397541600, 1397545200, 1397548800, 
    1397552400, 1397556000, 1397559600, 1397563200, 1397566800, 1397570400, 
    1397574000, 1397577600, 1397581200, 1397584800, 1397588400, 1397592000, 
    1397595600, 1397599200, 1397602800, 1397606400, 1397610000, 1397613600, 
    1397617200, 1397620800, 1397624400, 1397628000, 1397631600, 1397635200, 
    1397638800, 1397642400, 1397646000, 1397649600, 1397653200, 1397656800, 
    1397660400, 1397664000, 1397667600, 1397671200, 1397674800, 1397678400, 
    1397682000, 1397685600, 1397689200, 1397692800, 1397696400, 1397700000, 
    1397703600, 1397707200, 1397710800, 1397714400, 1397718000, 1397721600, 
    1397725200, 1397728800, 1397732400, 1397736000, 1397739600, 1397743200, 
    1397746800, 1397750400, 1397754000, 1397757600, 1397761200, 1397764800, 
    1397768400, 1397772000, 1397775600, 1397779200, 1397782800, 1397786400, 
    1397790000, 1397793600, 1397797200, 1397800800, 1397804400, 1397808000, 
    1397811600, 1397815200, 1397818800, 1397822400, 1397826000, 1397829600, 
    1397833200, 1397836800, 1397840400, 1397844000, 1397847600, 1397851200, 
    1397854800, 1397858400, 1397862000, 1397865600, 1397869200, 1397872800, 
    1397876400, 1397880000, 1397883600, 1397887200, 1397890800, 1397894400, 
    1397898000, 1397901600, 1397905200, 1397908800, 1397912400, 1397916000, 
    1397919600, 1397923200, 1397926800, 1397930400, 1397934000, 1397937600, 
    1397941200, 1397944800, 1397948400, 1397952000, 1397955600, 1397959200, 
    1397962800, 1397966400, 1397970000, 1397973600, 1397977200, 1397980800, 
    1397984400, 1397988000, 1397991600, 1397995200, 1397998800, 1398002400, 
    1398006000, 1398009600, 1398013200, 1398016800, 1398020400, 1398024000, 
    1398027600, 1398031200, 1398034800, 1398038400, 1398042000, 1398045600, 
    1398049200, 1398052800, 1398056400, 1398060000, 1398063600, 1398067200, 
    1398070800, 1398074400, 1398078000, 1398081600, 1398085200, 1398088800, 
    1398092400, 1398096000, 1398099600, 1398103200, 1398106800, 1398110400, 
    1398114000, 1398117600, 1398121200, 1398124800, 1398128400, 1398132000, 
    1398135600, 1398139200, 1398142800, 1398146400, 1398150000, 1398153600, 
    1398157200, 1398160800, 1398164400, 1398168000, 1398171600, 1398175200, 
    1398178800, 1398182400, 1398186000, 1398189600, 1398193200, 1398196800, 
    1398200400, 1398204000, 1398207600, 1398211200, 1398214800, 1398218400, 
    1398222000, 1398225600, 1398229200, 1398232800, 1398236400, 1398240000, 
    1398243600, 1398247200, 1398250800, 1398254400, 1398258000, 1398261600, 
    1398265200, 1398268800, 1398272400, 1398276000, 1398279600, 1398283200, 
    1398286800, 1398290400, 1398294000, 1398297600, 1398301200, 1398304800, 
    1398308400, 1398312000, 1398315600, 1398319200, 1398322800, 1398326400, 
    1398330000, 1398333600, 1398337200, 1398340800, 1398344400, 1398348000, 
    1398351600, 1398355200, 1398358800, 1398362400, 1398366000, 1398369600, 
    1398373200, 1398376800, 1398380400, 1398384000, 1398387600, 1398391200, 
    1398394800, 1398398400, 1398402000, 1398405600, 1398409200, 1398412800, 
    1398416400, 1398420000, 1398423600, 1398427200, 1398430800, 1398434400, 
    1398438000, 1398441600, 1398445200, 1398448800, 1398452400, 1398456000, 
    1398459600, 1398463200, 1398466800, 1398470400, 1398474000, 1398477600, 
    1398481200, 1398484800, 1398488400, 1398492000, 1398495600, 1398499200, 
    1398502800, 1398506400, 1398510000, 1398513600, 1398517200, 1398520800, 
    1398524400, 1398528000, 1398531600, 1398535200, 1398538800, 1398542400, 
    1398546000, 1398549600, 1398553200, 1398556800, 1398560400, 1398564000, 
    1398567600, 1398571200, 1398574800, 1398578400, 1398582000, 1398585600, 
    1398589200, 1398592800, 1398596400, 1398600000, 1398603600, 1398607200, 
    1398610800, 1398614400, 1398618000, 1398621600, 1398625200, 1398628800, 
    1398632400, 1398636000, 1398639600, 1398643200, 1398646800, 1398650400, 
    1398654000, 1398657600, 1398661200, 1398664800, 1398668400, 1398672000, 
    1398675600, 1398679200, 1398682800, 1398686400, 1398690000, 1398693600, 
    1398697200, 1398700800, 1398704400, 1398708000, 1398711600, 1398715200, 
    1398718800, 1398722400, 1398726000, 1398729600, 1398733200, 1398736800, 
    1398740400, 1398744000, 1398747600, 1398751200, 1398754800, 1398758400, 
    1398762000, 1398765600, 1398769200, 1398772800, 1398776400, 1398780000, 
    1398783600, 1398787200, 1398790800, 1398794400, 1398798000, 1398801600, 
    1398805200, 1398808800, 1398812400, 1398816000, 1398819600, 1398823200, 
    1398826800, 1398830400, 1398834000, 1398837600, 1398841200, 1398844800, 
    1398848400, 1398852000, 1398855600, 1398859200, 1398862800, 1398866400, 
    1398870000, 1398873600, 1398877200, 1398880800, 1398884400, 1398888000, 
    1398891600, 1398895200, 1398898800, 1398902400, 1398906000, 1398909600, 
    1398913200, 1398916800, 1398920400, 1398924000, 1398927600, 1398931200, 
    1398934800, 1398938400, 1398942000, 1398945600, 1398949200, 1398952800, 
    1398956400, 1398960000, 1398963600, 1398967200, 1398970800, 1398974400, 
    1398978000, 1398981600, 1398985200, 1398988800, 1398992400, 1398996000, 
    1398999600, 1399003200, 1399006800, 1399010400, 1399014000, 1399017600, 
    1399021200, 1399024800, 1399028400, 1399032000, 1399035600, 1399039200, 
    1399042800, 1399046400, 1399050000, 1399053600, 1399057200, 1399060800, 
    1399064400, 1399068000, 1399071600, 1399075200, 1399078800, 1399082400, 
    1399086000, 1399089600, 1399093200, 1399096800, 1399100400, 1399104000, 
    1399107600, 1399111200, 1399114800, 1399118400, 1399122000, 1399125600, 
    1399129200, 1399132800, 1399136400, 1399140000, 1399143600, 1399147200, 
    1399150800, 1399154400, 1399158000, 1399161600, 1399165200, 1399168800, 
    1399172400, 1399176000, 1399179600, 1399183200, 1399186800, 1399190400, 
    1399194000, 1399197600, 1399201200, 1399204800, 1399208400, 1399212000, 
    1399215600, 1399219200, 1399222800, 1399226400, 1399230000, 1399233600, 
    1399237200, 1399240800, 1399244400, 1399248000, 1399251600, 1399255200, 
    1399258800, 1399262400, 1399266000, 1399269600, 1399273200, 1399276800, 
    1399280400, 1399284000, 1399287600, 1399291200, 1399294800, 1399298400, 
    1399302000, 1399305600, 1399309200, 1399312800, 1399316400, 1399320000, 
    1399323600, 1399327200, 1399330800, 1399334400, 1399338000, 1399341600, 
    1399345200, 1399348800, 1399352400, 1399356000, 1399359600, 1399363200, 
    1399366800, 1399370400, 1399374000, 1399377600, 1399381200, 1399384800, 
    1399388400, 1399392000, 1399395600, 1399399200, 1399402800, 1399406400, 
    1399410000, 1399413600, 1399417200, 1399420800, 1399424400, 1399428000, 
    1399431600, 1399435200, 1399438800, 1399442400, 1399446000, 1399449600, 
    1399453200, 1399456800, 1399460400, 1399464000, 1399467600, 1399471200, 
    1399474800, 1399478400, 1399482000, 1399485600, 1399489200, 1399492800, 
    1399496400, 1399500000, 1399503600, 1399507200, 1399510800, 1399514400, 
    1399518000, 1399521600, 1399525200, 1399528800, 1399532400, 1399536000, 
    1399539600, 1399543200, 1399546800, 1399550400, 1399554000, 1399557600, 
    1399561200, 1399564800, 1399568400, 1399572000, 1399575600, 1399579200, 
    1399582800, 1399586400, 1399590000, 1399593600, 1399597200, 1399600800, 
    1399604400, 1399608000, 1399611600, 1399615200, 1399618800, 1399622400, 
    1399626000, 1399629600, 1399633200, 1399636800, 1399640400, 1399644000, 
    1399647600, 1399651200, 1399654800, 1399658400, 1399662000, 1399665600, 
    1399669200, 1399672800, 1399676400, 1399680000, 1399683600, 1399687200, 
    1399690800, 1399694400, 1399698000, 1399701600, 1399705200, 1399708800, 
    1399712400, 1399716000, 1399719600, 1399723200, 1399726800, 1399730400, 
    1399734000, 1399737600, 1399741200, 1399744800, 1399748400, 1399752000, 
    1399755600, 1399759200, 1399762800, 1399766400, 1399770000, 1399773600, 
    1399777200, 1399780800, 1399784400, 1399788000, 1399791600, 1399795200, 
    1399798800, 1399802400, 1399806000, 1399809600, 1399813200, 1399816800, 
    1399820400, 1399824000, 1399827600, 1399831200, 1399834800, 1399838400, 
    1399842000, 1399845600, 1399849200, 1399852800, 1399856400, 1399860000, 
    1399863600, 1399867200, 1399870800, 1399874400, 1399878000, 1399881600, 
    1399885200, 1399888800, 1399892400, 1399896000, 1399899600, 1399903200, 
    1399906800, 1399910400, 1399914000, 1399917600, 1399921200, 1399924800, 
    1399928400, 1399932000, 1399935600, 1399939200, 1399942800, 1399946400, 
    1399950000, 1399953600, 1399957200, 1399960800, 1399964400, 1399968000, 
    1399971600, 1399975200, 1399978800, 1399982400, 1399986000, 1399989600, 
    1399993200, 1399996800, 1400000400, 1400004000, 1400007600, 1400011200, 
    1400014800, 1400018400, 1400022000, 1400025600, 1400029200, 1400032800, 
    1400036400, 1400040000, 1400043600, 1400047200, 1400050800, 1400054400, 
    1400058000, 1400061600, 1400065200, 1400068800, 1400072400, 1400076000, 
    1400079600, 1400083200, 1400086800, 1400090400, 1400094000, 1400097600, 
    1400101200, 1400104800, 1400108400, 1400112000, 1400115600, 1400119200, 
    1400122800, 1400126400, 1400130000, 1400133600, 1400137200, 1400140800, 
    1400144400, 1400148000, 1400151600, 1400155200, 1400158800, 1400162400, 
    1400166000, 1400169600, 1400173200, 1400176800, 1400180400, 1400184000, 
    1400187600, 1400191200, 1400194800, 1400198400, 1400202000, 1400205600, 
    1400209200, 1400212800, 1400216400, 1400220000, 1400223600, 1400227200, 
    1400230800, 1400234400, 1400238000, 1400241600, 1400245200, 1400248800, 
    1400252400, 1400256000, 1400259600, 1400263200, 1400266800, 1400270400, 
    1400274000, 1400277600, 1400281200, 1400284800, 1400288400, 1400292000, 
    1400295600, 1400299200, 1400302800, 1400306400, 1400310000, 1400313600, 
    1400317200, 1400320800, 1400324400, 1400328000, 1400331600, 1400335200, 
    1400338800, 1400342400, 1400346000, 1400349600, 1400353200, 1400356800, 
    1400360400, 1400364000, 1400367600, 1400371200, 1400374800, 1400378400, 
    1400382000, 1400385600, 1400389200, 1400392800, 1400396400, 1400400000, 
    1400403600, 1400407200, 1400410800, 1400414400, 1400418000, 1400421600, 
    1400425200, 1400428800, 1400432400, 1400436000, 1400439600, 1400443200, 
    1400446800, 1400450400, 1400454000, 1400457600, 1400461200, 1400464800, 
    1400468400, 1400472000, 1400475600, 1400479200, 1400482800, 1400486400, 
    1400490000, 1400493600, 1400497200, 1400500800, 1400504400, 1400508000, 
    1400511600, 1400515200, 1400518800, 1400522400, 1400526000, 1400529600, 
    1400533200, 1400536800, 1400540400, 1400544000, 1400547600, 1400551200, 
    1400554800, 1400558400, 1400562000, 1400565600, 1400569200, 1400572800, 
    1400576400, 1400580000, 1400583600, 1400587200, 1400590800, 1400594400, 
    1400598000, 1400601600, 1400605200, 1400608800, 1400612400, 1400616000, 
    1400619600, 1400623200, 1400626800, 1400630400, 1400634000, 1400637600, 
    1400641200, 1400644800, 1400648400, 1400652000, 1400655600, 1400659200, 
    1400662800, 1400666400, 1400670000, 1400673600, 1400677200, 1400680800, 
    1400684400, 1400688000, 1400691600, 1400695200, 1400698800, 1400702400, 
    1400706000, 1400709600, 1400713200, 1400716800, 1400720400, 1400724000, 
    1400727600, 1400731200, 1400734800, 1400738400, 1400742000, 1400745600, 
    1400749200, 1400752800, 1400756400, 1400760000, 1400763600, 1400767200, 
    1400770800, 1400774400, 1400778000, 1400781600, 1400785200, 1400788800, 
    1400792400, 1400796000, 1400799600, 1400803200, 1400806800, 1400810400, 
    1400814000, 1400817600, 1400821200, 1400824800, 1400828400, 1400832000, 
    1400835600, 1400839200, 1400842800, 1400846400, 1400850000, 1400853600, 
    1400857200, 1400860800, 1400864400, 1400868000, 1400871600, 1400875200, 
    1400878800, 1400882400, 1400886000, 1400889600, 1400893200, 1400896800, 
    1400900400, 1400904000, 1400907600, 1400911200, 1400914800, 1400918400, 
    1400922000, 1400925600, 1400929200, 1400932800, 1400936400, 1400940000, 
    1400943600, 1400947200, 1400950800, 1400954400, 1400958000, 1400961600, 
    1400965200, 1400968800, 1400972400, 1400976000, 1400979600, 1400983200, 
    1400986800, 1400990400, 1400994000, 1400997600, 1401001200, 1401004800, 
    1401008400, 1401012000, 1401015600, 1401019200, 1401022800, 1401026400, 
    1401030000, 1401033600, 1401037200, 1401040800, 1401044400, 1401048000, 
    1401051600, 1401055200, 1401058800, 1401062400, 1401066000, 1401069600, 
    1401073200, 1401076800, 1401080400, 1401084000, 1401087600, 1401091200, 
    1401094800, 1401098400, 1401102000, 1401105600, 1401109200, 1401112800, 
    1401116400, 1401120000, 1401123600, 1401127200, 1401130800, 1401134400, 
    1401138000, 1401141600, 1401145200, 1401148800, 1401152400, 1401156000, 
    1401159600, 1401163200, 1401166800, 1401170400, 1401174000, 1401177600, 
    1401181200, 1401184800, 1401188400, 1401192000, 1401195600, 1401199200, 
    1401202800, 1401206400, 1401210000, 1401213600, 1401217200, 1401220800, 
    1401224400, 1401228000, 1401231600, 1401235200, 1401238800, 1401242400, 
    1401246000, 1401249600, 1401253200, 1401256800, 1401260400, 1401264000, 
    1401267600, 1401271200, 1401274800, 1401278400, 1401282000, 1401285600, 
    1401289200, 1401292800, 1401296400, 1401300000, 1401303600, 1401307200, 
    1401310800, 1401314400, 1401318000, 1401321600, 1401325200, 1401328800, 
    1401332400, 1401336000, 1401339600, 1401343200, 1401346800, 1401350400, 
    1401354000, 1401357600, 1401361200, 1401364800, 1401368400, 1401372000, 
    1401375600, 1401379200, 1401382800, 1401386400, 1401390000, 1401393600, 
    1401397200, 1401400800, 1401404400, 1401408000, 1401411600, 1401415200, 
    1401418800, 1401422400, 1401426000, 1401429600, 1401433200, 1401436800, 
    1401440400, 1401444000, 1401447600, 1401451200, 1401454800, 1401458400, 
    1401462000, 1401465600, 1401469200, 1401472800, 1401476400, 1401480000, 
    1401483600, 1401487200, 1401490800, 1401494400, 1401498000, 1401501600, 
    1401505200, 1401508800, 1401512400, 1401516000, 1401519600, 1401523200, 
    1401526800, 1401530400, 1401534000, 1401537600, 1401541200, 1401544800, 
    1401548400, 1401552000, 1401555600, 1401559200, 1401562800, 1401566400, 
    1401570000, 1401573600, 1401577200, 1401580800, 1401584400, 1401588000, 
    1401591600, 1401595200, 1401598800, 1401602400, 1401606000, 1401609600, 
    1401613200, 1401616800, 1401620400, 1401624000, 1401627600, 1401631200, 
    1401634800, 1401638400, 1401642000, 1401645600, 1401649200, 1401652800, 
    1401656400, 1401660000, 1401663600, 1401667200, 1401670800, 1401674400, 
    1401678000, 1401681600, 1401685200, 1401688800, 1401692400, 1401696000, 
    1401699600, 1401703200, 1401706800, 1401710400, 1401714000, 1401717600, 
    1401721200, 1401724800, 1401728400, 1401732000, 1401735600, 1401739200, 
    1401742800, 1401746400, 1401750000, 1401753600, 1401757200, 1401760800, 
    1401764400, 1401768000, 1401771600, 1401775200, 1401778800, 1401782400, 
    1401786000, 1401789600, 1401793200, 1401796800, 1401800400, 1401804000, 
    1401807600, 1401811200, 1401814800, 1401818400, 1401822000, 1401825600, 
    1401829200, 1401832800, 1401836400, 1401840000, 1401843600, 1401847200, 
    1401850800, 1401854400, 1401858000, 1401861600, 1401865200, 1401868800, 
    1401872400, 1401876000, 1401879600, 1401883200, 1401886800, 1401890400, 
    1401894000, 1401897600, 1401901200, 1401904800, 1401908400, 1401912000, 
    1401915600, 1401919200, 1401922800, 1401926400, 1401930000, 1401933600, 
    1401937200, 1401940800, 1401944400, 1401948000, 1401951600, 1401955200, 
    1401958800, 1401962400, 1401966000, 1401969600, 1401973200, 1401976800, 
    1401980400, 1401984000, 1401987600, 1401991200, 1401994800, 1401998400, 
    1402002000, 1402005600, 1402009200, 1402012800, 1402016400, 1402020000, 
    1402023600, 1402027200, 1402030800, 1402034400, 1402038000, 1402041600, 
    1402045200, 1402048800, 1402052400, 1402056000, 1402059600, 1402063200, 
    1402066800, 1402070400, 1402074000, 1402077600, 1402081200, 1402084800, 
    1402088400, 1402092000, 1402095600, 1402099200, 1402102800, 1402106400, 
    1402110000, 1402113600, 1402117200, 1402120800, 1402124400, 1402128000, 
    1402131600, 1402135200, 1402138800, 1402142400, 1402146000, 1402149600, 
    1402153200, 1402156800, 1402160400, 1402164000, 1402167600, 1402171200, 
    1402174800, 1402178400, 1402182000, 1402185600, 1402189200, 1402192800, 
    1402196400, 1402200000, 1402203600, 1402207200, 1402210800, 1402214400, 
    1402218000, 1402221600, 1402225200, 1402228800, 1402232400, 1402236000, 
    1402239600, 1402243200, 1402246800, 1402250400, 1402254000, 1402257600, 
    1402261200, 1402264800, 1402268400, 1402272000, 1402275600, 1402279200, 
    1402282800, 1402286400, 1402290000, 1402293600, 1402297200, 1402300800, 
    1402304400, 1402308000, 1402311600, 1402315200, 1402318800, 1402322400, 
    1402326000, 1402329600, 1402333200, 1402336800, 1402340400, 1402344000, 
    1402347600, 1402351200, 1402354800, 1402358400, 1402362000, 1402365600, 
    1402369200, 1402372800, 1402376400, 1402380000, 1402383600, 1402387200, 
    1402390800, 1402394400, 1402398000, 1402401600, 1402405200, 1402408800, 
    1402412400, 1402416000, 1402419600, 1402423200, 1402426800, 1402430400, 
    1402434000, 1402437600, 1402441200, 1402444800, 1402448400, 1402452000, 
    1402455600, 1402459200, 1402462800, 1402466400, 1402470000, 1402473600, 
    1402477200, 1402480800, 1402484400, 1402488000, 1402491600, 1402495200, 
    1402498800, 1402502400, 1402506000, 1402509600, 1402513200, 1402516800, 
    1402520400, 1402524000, 1402527600, 1402531200, 1402534800, 1402538400, 
    1402542000, 1402545600, 1402549200, 1402552800, 1402556400, 1402560000, 
    1402563600, 1402567200, 1402570800, 1402574400, 1402578000, 1402581600, 
    1402585200, 1402588800, 1402592400, 1402596000, 1402599600, 1402603200, 
    1402606800, 1402610400, 1402614000, 1402617600, 1402621200, 1402624800, 
    1402628400, 1402632000, 1402635600, 1402639200, 1402642800, 1402646400, 
    1402650000, 1402653600, 1402657200, 1402660800, 1402664400, 1402668000, 
    1402671600, 1402675200, 1402678800, 1402682400, 1402686000, 1402689600, 
    1402693200, 1402696800, 1402700400, 1402704000, 1402707600, 1402711200, 
    1402714800, 1402718400, 1402722000, 1402725600, 1402729200, 1402732800, 
    1402736400, 1402740000, 1402743600, 1402747200, 1402750800, 1402754400, 
    1402758000, 1402761600, 1402765200, 1402768800, 1402772400, 1402776000, 
    1402779600, 1402783200, 1402786800, 1402790400, 1402794000, 1402797600, 
    1402801200, 1402804800, 1402808400, 1402812000, 1402815600, 1402819200, 
    1402822800, 1402826400, 1402830000, 1402833600, 1402837200, 1402840800, 
    1402844400, 1402848000, 1402851600, 1402855200, 1402858800, 1402862400, 
    1402866000, 1402869600, 1402873200, 1402876800, 1402880400, 1402884000, 
    1402887600, 1402891200, 1402894800, 1402898400, 1402902000, 1402905600, 
    1402909200, 1402912800, 1402916400, 1402920000, 1402923600, 1402927200, 
    1402930800, 1402934400, 1402938000, 1402941600, 1402945200, 1402948800, 
    1402952400, 1402956000, 1402959600, 1402963200, 1402966800, 1402970400, 
    1402974000, 1402977600, 1402981200, 1402984800, 1402988400, 1402992000, 
    1402995600, 1402999200, 1403002800, 1403006400, 1403010000, 1403013600, 
    1403017200, 1403020800, 1403024400, 1403028000, 1403031600, 1403035200, 
    1403038800, 1403042400, 1403046000, 1403049600, 1403053200, 1403056800, 
    1403060400, 1403064000, 1403067600, 1403071200, 1403074800, 1403078400, 
    1403082000, 1403085600, 1403089200, 1403092800, 1403096400, 1403100000, 
    1403103600, 1403107200, 1403110800, 1403114400, 1403118000, 1403121600, 
    1403125200, 1403128800, 1403132400, 1403136000, 1403139600, 1403143200, 
    1403146800, 1403150400, 1403154000, 1403157600, 1403161200, 1403164800, 
    1403168400, 1403172000, 1403175600, 1403179200, 1403182800, 1403186400, 
    1403190000, 1403193600, 1403197200, 1403200800, 1403204400, 1403208000, 
    1403211600, 1403215200, 1403218800, 1403222400, 1403226000, 1403229600, 
    1403233200, 1403236800, 1403240400, 1403244000, 1403247600, 1403251200, 
    1403254800, 1403258400, 1403262000, 1403265600, 1403269200, 1403272800, 
    1403276400, 1403280000, 1403283600, 1403287200, 1403290800, 1403294400, 
    1403298000, 1403301600, 1403305200, 1403308800, 1403312400, 1403316000, 
    1403319600, 1403323200, 1403326800, 1403330400, 1403334000, 1403337600, 
    1403341200, 1403344800, 1403348400, 1403352000, 1403355600, 1403359200, 
    1403362800, 1403366400, 1403370000, 1403373600, 1403377200, 1403380800, 
    1403384400, 1403388000, 1403391600, 1403395200, 1403398800, 1403402400, 
    1403406000, 1403409600, 1403413200, 1403416800, 1403420400, 1403424000, 
    1403427600, 1403431200, 1403434800, 1403438400, 1403442000, 1403445600, 
    1403449200, 1403452800, 1403456400, 1403460000, 1403463600, 1403467200, 
    1403470800, 1403474400, 1403478000, 1403481600, 1403485200, 1403488800, 
    1403492400, 1403496000, 1403499600, 1403503200, 1403506800, 1403510400, 
    1403514000, 1403517600, 1403521200, 1403524800, 1403528400, 1403532000, 
    1403535600, 1403539200, 1403542800, 1403546400, 1403550000, 1403553600, 
    1403557200, 1403560800, 1403564400, 1403568000, 1403571600, 1403575200, 
    1403578800, 1403582400, 1403586000, 1403589600, 1403593200, 1403596800, 
    1403600400, 1403604000, 1403607600, 1403611200, 1403614800, 1403618400, 
    1403622000, 1403625600, 1403629200, 1403632800, 1403636400, 1403640000, 
    1403643600, 1403647200, 1403650800, 1403654400, 1403658000, 1403661600, 
    1403665200, 1403668800, 1403672400, 1403676000, 1403679600, 1403683200, 
    1403686800, 1403690400, 1403694000, 1403697600, 1403701200, 1403704800, 
    1403708400, 1403712000, 1403715600, 1403719200, 1403722800, 1403726400, 
    1403730000, 1403733600, 1403737200, 1403740800, 1403744400, 1403748000, 
    1403751600, 1403755200, 1403758800, 1403762400, 1403766000, 1403769600, 
    1403773200, 1403776800, 1403780400, 1403784000, 1403787600, 1403791200, 
    1403794800, 1403798400, 1403802000, 1403805600, 1403809200, 1403812800, 
    1403816400, 1403820000, 1403823600, 1403827200, 1403830800, 1403834400, 
    1403838000, 1403841600, 1403845200, 1403848800, 1403852400, 1403856000, 
    1403859600, 1403863200, 1403866800, 1403870400, 1403874000, 1403877600, 
    1403881200, 1403884800, 1403888400, 1403892000, 1403895600, 1403899200, 
    1403902800, 1403906400, 1403910000, 1403913600, 1403917200, 1403920800, 
    1403924400, 1403928000, 1403931600, 1403935200, 1403938800, 1403942400, 
    1403946000, 1403949600, 1403953200, 1403956800, 1403960400, 1403964000, 
    1403967600, 1403971200, 1403974800, 1403978400, 1403982000, 1403985600, 
    1403989200, 1403992800, 1403996400, 1404000000, 1404003600, 1404007200, 
    1404010800, 1404014400, 1404018000, 1404021600, 1404025200, 1404028800, 
    1404032400, 1404036000, 1404039600, 1404043200, 1404046800, 1404050400, 
    1404054000, 1404057600, 1404061200, 1404064800, 1404068400, 1404072000, 
    1404075600, 1404079200, 1404082800, 1404086400, 1404090000, 1404093600, 
    1404097200, 1404100800, 1404104400, 1404108000, 1404111600, 1404115200, 
    1404118800, 1404122400, 1404126000, 1404129600, 1404133200, 1404136800, 
    1404140400, 1404144000, 1404147600, 1404151200, 1404154800, 1404158400, 
    1404162000, 1404165600, 1404169200, 1404172800, 1404176400, 1404180000, 
    1404183600, 1404187200, 1404190800, 1404194400, 1404198000, 1404201600, 
    1404205200, 1404208800, 1404212400, 1404216000, 1404219600, 1404223200, 
    1404226800, 1404230400, 1404234000, 1404237600, 1404241200, 1404244800, 
    1404248400, 1404252000, 1404255600, 1404259200, 1404262800, 1404266400, 
    1404270000, 1404273600, 1404277200, 1404280800, 1404284400, 1404288000, 
    1404291600, 1404295200, 1404298800, 1404302400, 1404306000, 1404309600, 
    1404313200, 1404316800, 1404320400, 1404324000, 1404327600, 1404331200, 
    1404334800, 1404338400, 1404342000, 1404345600, 1404349200, 1404352800, 
    1404356400, 1404360000, 1404363600, 1404367200, 1404370800, 1404374400, 
    1404378000, 1404381600, 1404385200, 1404388800, 1404392400, 1404396000, 
    1404399600, 1404403200, 1404406800, 1404410400, 1404414000, 1404417600, 
    1404421200, 1404424800, 1404428400, 1404432000, 1404435600, 1404439200, 
    1404442800, 1404446400, 1404450000, 1404453600, 1404457200, 1404460800, 
    1404464400, 1404468000, 1404471600, 1404475200, 1404478800, 1404482400, 
    1404486000, 1404489600, 1404493200, 1404496800, 1404500400, 1404504000, 
    1404507600, 1404511200, 1404514800, 1404518400, 1404522000, 1404525600, 
    1404529200, 1404532800, 1404536400, 1404540000, 1404543600, 1404547200, 
    1404550800, 1404554400, 1404558000, 1404561600, 1404565200, 1404568800, 
    1404572400, 1404576000, 1404579600, 1404583200, 1404586800, 1404590400, 
    1404594000, 1404597600, 1404601200, 1404604800, 1404608400, 1404612000, 
    1404615600, 1404619200, 1404622800, 1404626400, 1404630000, 1404633600, 
    1404637200, 1404640800, 1404644400, 1404648000, 1404651600, 1404655200, 
    1404658800, 1404662400, 1404666000, 1404669600, 1404673200, 1404676800, 
    1404680400, 1404684000, 1404687600, 1404691200, 1404694800, 1404698400, 
    1404702000, 1404705600, 1404709200, 1404712800, 1404716400, 1404720000, 
    1404723600, 1404727200, 1404730800, 1404734400, 1404738000, 1404741600, 
    1404745200, 1404748800, 1404752400, 1404756000, 1404759600, 1404763200, 
    1404766800, 1404770400, 1404774000, 1404777600, 1404781200, 1404784800, 
    1404788400, 1404792000, 1404795600, 1404799200, 1404802800, 1404806400, 
    1404810000, 1404813600, 1404817200, 1404820800, 1404824400, 1404828000, 
    1404831600, 1404835200, 1404838800, 1404842400, 1404846000, 1404849600, 
    1404853200, 1404856800, 1404860400, 1404864000, 1404867600, 1404871200, 
    1404874800, 1404878400, 1404882000, 1404885600, 1404889200, 1404892800, 
    1404896400, 1404900000, 1404903600, 1404907200, 1404910800, 1404914400, 
    1404918000, 1404921600, 1404925200, 1404928800, 1404932400, 1404936000, 
    1404939600, 1404943200, 1404946800, 1404950400, 1404954000, 1404957600, 
    1404961200, 1404964800, 1404968400, 1404972000, 1404975600, 1404979200, 
    1404982800, 1404986400, 1404990000, 1404993600, 1404997200, 1405000800, 
    1405004400, 1405008000, 1405011600, 1405015200, 1405018800, 1405022400, 
    1405026000, 1405029600, 1405033200, 1405036800, 1405040400, 1405044000, 
    1405047600, 1405051200, 1405054800, 1405058400, 1405062000, 1405065600, 
    1405069200, 1405072800, 1405076400, 1405080000, 1405083600, 1405087200, 
    1405090800, 1405094400, 1405098000, 1405101600, 1405105200, 1405108800, 
    1405112400, 1405116000, 1405119600, 1405123200, 1405126800, 1405130400, 
    1405134000, 1405137600, 1405141200, 1405144800, 1405148400, 1405152000, 
    1405155600, 1405159200, 1405162800, 1405166400, 1405170000, 1405173600, 
    1405177200, 1405180800, 1405184400, 1405188000, 1405191600, 1405195200, 
    1405198800, 1405202400, 1405206000, 1405209600, 1405213200, 1405216800, 
    1405220400, 1405224000, 1405227600, 1405231200, 1405234800, 1405238400, 
    1405242000, 1405245600, 1405249200, 1405252800, 1405256400, 1405260000, 
    1405263600, 1405267200, 1405270800, 1405274400, 1405278000, 1405281600, 
    1405285200, 1405288800, 1405292400, 1405296000, 1405299600, 1405303200, 
    1405306800, 1405310400, 1405314000, 1405317600, 1405321200, 1405324800, 
    1405328400, 1405332000, 1405335600, 1405339200, 1405342800, 1405346400, 
    1405350000, 1405353600, 1405357200, 1405360800, 1405364400, 1405368000, 
    1405371600, 1405375200, 1405378800, 1405382400, 1405386000, 1405389600, 
    1405393200, 1405396800, 1405400400, 1405404000, 1405407600, 1405411200, 
    1405414800, 1405418400, 1405422000, 1405425600, 1405429200, 1405432800, 
    1405436400, 1405440000, 1405443600, 1405447200, 1405450800, 1405454400, 
    1405458000, 1405461600, 1405465200, 1405468800, 1405472400, 1405476000, 
    1405479600, 1405483200, 1405486800, 1405490400, 1405494000, 1405497600, 
    1405501200, 1405504800, 1405508400, 1405512000, 1405515600, 1405519200, 
    1405522800, 1405526400, 1405530000, 1405533600, 1405537200, 1405540800, 
    1405544400, 1405548000, 1405551600, 1405555200, 1405558800, 1405562400, 
    1405566000, 1405569600, 1405573200, 1405576800, 1405580400, 1405584000, 
    1405587600, 1405591200, 1405594800, 1405598400, 1405602000, 1405605600, 
    1405609200, 1405612800, 1405616400, 1405620000, 1405623600, 1405627200, 
    1405630800, 1405634400, 1405638000, 1405641600, 1405645200, 1405648800, 
    1405652400, 1405656000, 1405659600, 1405663200, 1405666800, 1405670400, 
    1405674000, 1405677600, 1405681200, 1405684800, 1405688400, 1405692000, 
    1405695600, 1405699200, 1405702800, 1405706400, 1405710000, 1405713600, 
    1405717200, 1405720800, 1405724400, 1405728000, 1405731600, 1405735200, 
    1405738800, 1405742400, 1405746000, 1405749600, 1405753200, 1405756800, 
    1405760400, 1405764000, 1405767600, 1405771200, 1405774800, 1405778400, 
    1405782000, 1405785600, 1405789200, 1405792800, 1405796400, 1405800000, 
    1405803600, 1405807200, 1405810800, 1405814400, 1405818000, 1405821600, 
    1405825200, 1405828800, 1405832400, 1405836000, 1405839600, 1405843200, 
    1405846800, 1405850400, 1405854000, 1405857600, 1405861200, 1405864800, 
    1405868400, 1405872000, 1405875600, 1405879200, 1405882800, 1405886400, 
    1405890000, 1405893600, 1405897200, 1405900800, 1405904400, 1405908000, 
    1405911600, 1405915200, 1405918800, 1405922400, 1405926000, 1405929600, 
    1405933200, 1405936800, 1405940400, 1405944000, 1405947600, 1405951200, 
    1405954800, 1405958400, 1405962000, 1405965600, 1405969200, 1405972800, 
    1405976400, 1405980000, 1405983600, 1405987200, 1405990800, 1405994400, 
    1405998000, 1406001600, 1406005200, 1406008800, 1406012400, 1406016000, 
    1406019600, 1406023200, 1406026800, 1406030400, 1406034000, 1406037600, 
    1406041200, 1406044800, 1406048400, 1406052000, 1406055600, 1406059200, 
    1406062800, 1406066400, 1406070000, 1406073600, 1406077200, 1406080800, 
    1406084400, 1406088000, 1406091600, 1406095200, 1406098800, 1406102400, 
    1406106000, 1406109600, 1406113200, 1406116800, 1406120400, 1406124000, 
    1406127600, 1406131200, 1406134800, 1406138400, 1406142000, 1406145600, 
    1406149200, 1406152800, 1406156400, 1406160000, 1406163600, 1406167200, 
    1406170800, 1406174400, 1406178000, 1406181600, 1406185200, 1406188800, 
    1406192400, 1406196000, 1406199600, 1406203200, 1406206800, 1406210400, 
    1406214000, 1406217600, 1406221200, 1406224800, 1406228400, 1406232000, 
    1406235600, 1406239200, 1406242800, 1406246400, 1406250000, 1406253600, 
    1406257200, 1406260800, 1406264400, 1406268000, 1406271600, 1406275200, 
    1406278800, 1406282400, 1406286000, 1406289600, 1406293200, 1406296800, 
    1406300400, 1406304000, 1406307600, 1406311200, 1406314800, 1406318400, 
    1406322000, 1406325600, 1406329200, 1406332800, 1406336400, 1406340000, 
    1406343600, 1406347200, 1406350800, 1406354400, 1406358000, 1406361600, 
    1406365200, 1406368800, 1406372400, 1406376000, 1406379600, 1406383200, 
    1406386800, 1406390400, 1406394000, 1406397600, 1406401200, 1406404800, 
    1406408400, 1406412000, 1406415600, 1406419200, 1406422800, 1406426400, 
    1406430000, 1406433600, 1406437200, 1406440800, 1406444400, 1406448000, 
    1406451600, 1406455200, 1406458800, 1406462400, 1406466000, 1406469600, 
    1406473200, 1406476800, 1406480400, 1406484000, 1406487600, 1406491200, 
    1406494800, 1406498400, 1406502000, 1406505600, 1406509200, 1406512800, 
    1406516400, 1406520000, 1406523600, 1406527200, 1406530800, 1406534400, 
    1406538000, 1406541600, 1406545200, 1406548800, 1406552400, 1406556000, 
    1406559600, 1406563200, 1406566800, 1406570400, 1406574000, 1406577600, 
    1406581200, 1406584800, 1406588400, 1406592000, 1406595600, 1406599200, 
    1406602800, 1406606400, 1406610000, 1406613600, 1406617200, 1406620800, 
    1406624400, 1406628000, 1406631600, 1406635200, 1406638800, 1406642400, 
    1406646000, 1406649600, 1406653200, 1406656800, 1406660400, 1406664000, 
    1406667600, 1406671200, 1406674800, 1406678400, 1406682000, 1406685600, 
    1406689200, 1406692800, 1406696400, 1406700000, 1406703600, 1406707200, 
    1406710800, 1406714400, 1406718000, 1406721600, 1406725200, 1406728800, 
    1406732400, 1406736000, 1406739600, 1406743200, 1406746800, 1406750400, 
    1406754000, 1406757600, 1406761200, 1406764800, 1406768400, 1406772000, 
    1406775600, 1406779200, 1406782800, 1406786400, 1406790000, 1406793600, 
    1406797200, 1406800800, 1406804400, 1406808000, 1406811600, 1406815200, 
    1406818800, 1406822400, 1406826000, 1406829600, 1406833200, 1406836800, 
    1406840400, 1406844000, 1406847600, 1406851200, 1406854800, 1406858400, 
    1406862000, 1406865600, 1406869200, 1406872800, 1406876400, 1406880000, 
    1406883600, 1406887200, 1406890800, 1406894400, 1406898000, 1406901600, 
    1406905200, 1406908800, 1406912400, 1406916000, 1406919600, 1406923200, 
    1406926800, 1406930400, 1406934000, 1406937600, 1406941200, 1406944800, 
    1406948400, 1406952000, 1406955600, 1406959200, 1406962800, 1406966400, 
    1406970000, 1406973600, 1406977200, 1406980800, 1406984400, 1406988000, 
    1406991600, 1406995200, 1406998800, 1407002400, 1407006000, 1407009600, 
    1407013200, 1407016800, 1407020400, 1407024000, 1407027600, 1407031200, 
    1407034800, 1407038400, 1407042000, 1407045600, 1407049200, 1407052800, 
    1407056400, 1407060000, 1407063600, 1407067200, 1407070800, 1407074400, 
    1407078000, 1407081600, 1407085200, 1407088800, 1407092400, 1407096000, 
    1407099600, 1407103200, 1407106800, 1407110400, 1407114000, 1407117600, 
    1407121200, 1407124800, 1407128400, 1407132000, 1407135600, 1407139200, 
    1407142800, 1407146400, 1407150000, 1407153600, 1407157200, 1407160800, 
    1407164400, 1407168000, 1407171600, 1407175200, 1407178800, 1407182400, 
    1407186000, 1407189600, 1407193200, 1407196800, 1407200400, 1407204000, 
    1407207600, 1407211200, 1407214800, 1407218400, 1407222000, 1407225600, 
    1407229200, 1407232800, 1407236400, 1407240000, 1407243600, 1407247200, 
    1407250800, 1407254400, 1407258000, 1407261600, 1407265200, 1407268800, 
    1407272400, 1407276000, 1407279600, 1407283200, 1407286800, 1407290400, 
    1407294000, 1407297600, 1407301200, 1407304800, 1407308400, 1407312000, 
    1407315600, 1407319200, 1407322800, 1407326400, 1407330000, 1407333600, 
    1407337200, 1407340800, 1407344400, 1407348000, 1407351600, 1407355200, 
    1407358800, 1407362400, 1407366000, 1407369600, 1407373200, 1407376800, 
    1407380400, 1407384000, 1407387600, 1407391200, 1407394800, 1407398400, 
    1407402000, 1407405600, 1407409200, 1407412800, 1407416400, 1407420000, 
    1407423600, 1407427200, 1407430800, 1407434400, 1407438000, 1407441600, 
    1407445200, 1407448800, 1407452400, 1407456000, 1407459600, 1407463200, 
    1407466800, 1407470400, 1407474000, 1407477600, 1407481200, 1407484800, 
    1407488400, 1407492000, 1407495600, 1407499200, 1407502800, 1407506400, 
    1407510000, 1407513600, 1407517200, 1407520800, 1407524400, 1407528000, 
    1407531600, 1407535200, 1407538800, 1407542400, 1407546000, 1407549600, 
    1407553200, 1407556800, 1407560400, 1407564000, 1407567600, 1407571200, 
    1407574800, 1407578400, 1407582000, 1407585600, 1407589200, 1407592800, 
    1407596400, 1407600000, 1407603600, 1407607200, 1407610800, 1407614400, 
    1407618000, 1407621600, 1407625200, 1407628800, 1407632400, 1407636000, 
    1407639600, 1407643200, 1407646800, 1407650400, 1407654000, 1407657600, 
    1407661200, 1407664800, 1407668400, 1407672000, 1407675600, 1407679200, 
    1407682800, 1407686400, 1407690000, 1407693600, 1407697200, 1407700800, 
    1407704400, 1407708000, 1407711600, 1407715200, 1407718800, 1407722400, 
    1407726000, 1407729600, 1407733200, 1407736800, 1407740400, 1407744000, 
    1407747600, 1407751200, 1407754800, 1407758400, 1407762000, 1407765600, 
    1407769200, 1407772800, 1407776400, 1407780000, 1407783600, 1407787200, 
    1407790800, 1407794400, 1407798000, 1407801600, 1407805200, 1407808800, 
    1407812400, 1407816000, 1407819600, 1407823200, 1407826800, 1407830400, 
    1407834000, 1407837600, 1407841200, 1407844800, 1407848400, 1407852000, 
    1407855600, 1407859200, 1407862800, 1407866400, 1407870000, 1407873600, 
    1407877200, 1407880800, 1407884400, 1407888000, 1407891600, 1407895200, 
    1407898800, 1407902400, 1407906000, 1407909600, 1407913200, 1407916800, 
    1407920400, 1407924000, 1407927600, 1407931200, 1407934800, 1407938400, 
    1407942000, 1407945600, 1407949200, 1407952800, 1407956400, 1407960000, 
    1407963600, 1407967200, 1407970800, 1407974400, 1407978000, 1407981600, 
    1407985200, 1407988800, 1407992400, 1407996000, 1407999600, 1408003200, 
    1408006800, 1408010400, 1408014000, 1408017600, 1408021200, 1408024800, 
    1408028400, 1408032000, 1408035600, 1408039200, 1408042800, 1408046400, 
    1408050000, 1408053600, 1408057200, 1408060800, 1408064400, 1408068000, 
    1408071600, 1408075200, 1408078800, 1408082400, 1408086000, 1408089600, 
    1408093200, 1408096800, 1408100400, 1408104000, 1408107600, 1408111200, 
    1408114800, 1408118400, 1408122000, 1408125600, 1408129200, 1408132800, 
    1408136400, 1408140000, 1408143600, 1408147200, 1408150800, 1408154400, 
    1408158000, 1408161600, 1408165200, 1408168800, 1408172400, 1408176000, 
    1408179600, 1408183200, 1408186800, 1408190400, 1408194000, 1408197600, 
    1408201200, 1408204800, 1408208400, 1408212000, 1408215600, 1408219200, 
    1408222800, 1408226400, 1408230000, 1408233600, 1408237200, 1408240800, 
    1408244400, 1408248000, 1408251600, 1408255200, 1408258800, 1408262400, 
    1408266000, 1408269600, 1408273200, 1408276800, 1408280400, 1408284000, 
    1408287600, 1408291200, 1408294800, 1408298400, 1408302000, 1408305600, 
    1408309200, 1408312800, 1408316400, 1408320000, 1408323600, 1408327200, 
    1408330800, 1408334400, 1408338000, 1408341600, 1408345200, 1408348800, 
    1408352400, 1408356000, 1408359600, 1408363200, 1408366800, 1408370400, 
    1408374000, 1408377600, 1408381200, 1408384800, 1408388400, 1408392000, 
    1408395600, 1408399200, 1408402800, 1408406400, 1408410000, 1408413600, 
    1408417200, 1408420800, 1408424400, 1408428000, 1408431600, 1408435200, 
    1408438800, 1408442400, 1408446000, 1408449600, 1408453200, 1408456800, 
    1408460400, 1408464000, 1408467600, 1408471200, 1408474800, 1408478400, 
    1408482000, 1408485600, 1408489200, 1408492800, 1408496400, 1408500000, 
    1408503600, 1408507200, 1408510800, 1408514400, 1408518000, 1408521600, 
    1408525200, 1408528800, 1408532400, 1408536000, 1408539600, 1408543200, 
    1408546800, 1408550400, 1408554000, 1408557600, 1408561200, 1408564800, 
    1408568400, 1408572000, 1408575600, 1408579200, 1408582800, 1408586400, 
    1408590000, 1408593600, 1408597200, 1408600800, 1408604400, 1408608000, 
    1408611600, 1408615200, 1408618800, 1408622400, 1408626000, 1408629600, 
    1408633200, 1408636800, 1408640400, 1408644000, 1408647600, 1408651200, 
    1408654800, 1408658400, 1408662000, 1408665600, 1408669200, 1408672800, 
    1408676400, 1408680000, 1408683600, 1408687200, 1408690800, 1408694400, 
    1408698000, 1408701600, 1408705200, 1408708800, 1408712400, 1408716000, 
    1408719600, 1408723200, 1408726800, 1408730400, 1408734000, 1408737600, 
    1408741200, 1408744800, 1408748400, 1408752000, 1408755600, 1408759200, 
    1408762800, 1408766400, 1408770000, 1408773600, 1408777200, 1408780800, 
    1408784400, 1408788000, 1408791600, 1408795200, 1408798800, 1408802400, 
    1408806000, 1408809600, 1408813200, 1408816800, 1408820400, 1408824000, 
    1408827600, 1408831200, 1408834800, 1408838400, 1408842000, 1408845600, 
    1408849200, 1408852800, 1408856400, 1408860000, 1408863600, 1408867200, 
    1408870800, 1408874400, 1408878000, 1408881600, 1408885200, 1408888800, 
    1408892400, 1408896000, 1408899600, 1408903200, 1408906800, 1408910400, 
    1408914000, 1408917600, 1408921200, 1408924800, 1408928400, 1408932000, 
    1408935600, 1408939200, 1408942800, 1408946400, 1408950000, 1408953600, 
    1408957200, 1408960800, 1408964400, 1408968000, 1408971600, 1408975200, 
    1408978800, 1408982400, 1408986000, 1408989600, 1408993200, 1408996800, 
    1409000400, 1409004000, 1409007600, 1409011200, 1409014800, 1409018400, 
    1409022000, 1409025600, 1409029200, 1409032800, 1409036400, 1409040000, 
    1409043600, 1409047200, 1409050800, 1409054400, 1409058000, 1409061600, 
    1409065200, 1409068800, 1409072400, 1409076000, 1409079600, 1409083200, 
    1409086800, 1409090400, 1409094000, 1409097600, 1409101200, 1409104800, 
    1409108400, 1409112000, 1409115600, 1409119200, 1409122800, 1409126400, 
    1409130000, 1409133600, 1409137200, 1409140800, 1409144400, 1409148000, 
    1409151600, 1409155200, 1409158800, 1409162400, 1409166000, 1409169600, 
    1409173200, 1409176800, 1409180400, 1409184000, 1409187600, 1409191200, 
    1409194800, 1409198400, 1409202000, 1409205600, 1409209200, 1409212800, 
    1409216400, 1409220000, 1409223600, 1409227200, 1409230800, 1409234400, 
    1409238000, 1409241600, 1409245200, 1409248800, 1409252400, 1409256000, 
    1409259600, 1409263200, 1409266800, 1409270400, 1409274000, 1409277600, 
    1409281200, 1409284800, 1409288400, 1409292000, 1409295600, 1409299200, 
    1409302800, 1409306400, 1409310000, 1409313600, 1409317200, 1409320800, 
    1409324400, 1409328000, 1409331600, 1409335200, 1409338800, 1409342400, 
    1409346000, 1409349600, 1409353200, 1409356800, 1409360400, 1409364000, 
    1409367600, 1409371200, 1409374800, 1409378400, 1409382000, 1409385600, 
    1409389200, 1409392800, 1409396400, 1409400000, 1409403600, 1409407200, 
    1409410800, 1409414400, 1409418000, 1409421600, 1409425200, 1409428800, 
    1409432400, 1409436000, 1409439600, 1409443200, 1409446800, 1409450400, 
    1409454000, 1409457600, 1409461200, 1409464800, 1409468400, 1409472000, 
    1409475600, 1409479200, 1409482800, 1409486400, 1409490000, 1409493600, 
    1409497200, 1409500800, 1409504400, 1409508000, 1409511600, 1409515200, 
    1409518800, 1409522400, 1409526000, 1409529600, 1409533200, 1409536800, 
    1409540400, 1409544000, 1409547600, 1409551200, 1409554800, 1409558400, 
    1409562000, 1409565600, 1409569200, 1409572800, 1409576400, 1409580000, 
    1409583600, 1409587200, 1409590800, 1409594400, 1409598000, 1409601600, 
    1409605200, 1409608800, 1409612400, 1409616000, 1409619600, 1409623200, 
    1409626800, 1409630400, 1409634000, 1409637600, 1409641200, 1409644800, 
    1409648400, 1409652000, 1409655600, 1409659200, 1409662800, 1409666400, 
    1409670000, 1409673600, 1409677200, 1409680800, 1409684400, 1409688000, 
    1409691600, 1409695200, 1409698800, 1409702400, 1409706000, 1409709600, 
    1409713200, 1409716800, 1409720400, 1409724000, 1409727600, 1409731200, 
    1409734800, 1409738400, 1409742000, 1409745600, 1409749200, 1409752800, 
    1409756400, 1409760000, 1409763600, 1409767200, 1409770800, 1409774400, 
    1409778000, 1409781600, 1409785200, 1409788800, 1409792400, 1409796000, 
    1409799600, 1409803200, 1409806800, 1409810400, 1409814000, 1409817600, 
    1409821200, 1409824800, 1409828400, 1409832000, 1409835600, 1409839200, 
    1409842800, 1409846400, 1409850000, 1409853600, 1409857200, 1409860800, 
    1409864400, 1409868000, 1409871600, 1409875200, 1409878800, 1409882400, 
    1409886000, 1409889600, 1409893200, 1409896800, 1409900400, 1409904000, 
    1409907600, 1409911200, 1409914800, 1409918400, 1409922000, 1409925600, 
    1409929200, 1409932800, 1409936400, 1409940000, 1409943600, 1409947200, 
    1409950800, 1409954400, 1409958000, 1409961600, 1409965200, 1409968800, 
    1409972400, 1409976000, 1409979600, 1409983200, 1409986800, 1409990400, 
    1409994000, 1409997600, 1410001200, 1410004800, 1410008400, 1410012000, 
    1410015600, 1410019200, 1410022800, 1410026400, 1410030000, 1410033600, 
    1410037200, 1410040800, 1410044400, 1410048000, 1410051600, 1410055200, 
    1410058800, 1410062400, 1410066000, 1410069600, 1410073200, 1410076800, 
    1410080400, 1410084000, 1410087600, 1410091200, 1410094800, 1410098400, 
    1410102000, 1410105600, 1410109200, 1410112800, 1410116400, 1410120000, 
    1410123600, 1410127200, 1410130800, 1410134400, 1410138000, 1410141600, 
    1410145200, 1410148800, 1410152400, 1410156000, 1410159600, 1410163200, 
    1410166800, 1410170400, 1410174000, 1410177600, 1410181200, 1410184800, 
    1410188400, 1410192000, 1410195600, 1410199200, 1410202800, 1410206400, 
    1410210000, 1410213600, 1410217200, 1410220800, 1410224400, 1410228000, 
    1410231600, 1410235200, 1410238800, 1410242400, 1410246000, 1410249600, 
    1410253200, 1410256800, 1410260400, 1410264000, 1410267600, 1410271200, 
    1410274800, 1410278400, 1410282000, 1410285600, 1410289200, 1410292800, 
    1410296400, 1410300000, 1410303600, 1410307200, 1410310800, 1410314400, 
    1410318000, 1410321600, 1410325200, 1410328800, 1410332400, 1410336000, 
    1410339600, 1410343200, 1410346800, 1410350400, 1410354000, 1410357600, 
    1410361200, 1410364800, 1410368400, 1410372000, 1410375600, 1410379200, 
    1410382800, 1410386400, 1410390000, 1410393600, 1410397200, 1410400800, 
    1410404400, 1410408000, 1410411600, 1410415200, 1410418800, 1410422400, 
    1410426000, 1410429600, 1410433200, 1410436800, 1410440400, 1410444000, 
    1410447600, 1410451200, 1410454800, 1410458400, 1410462000, 1410465600, 
    1410469200, 1410472800, 1410476400, 1410480000, 1410483600, 1410487200, 
    1410490800, 1410494400, 1410498000, 1410501600, 1410505200, 1410508800, 
    1410512400, 1410516000, 1410519600, 1410523200, 1410526800, 1410530400, 
    1410534000, 1410537600, 1410541200, 1410544800, 1410548400, 1410552000, 
    1410555600, 1410559200, 1410562800, 1410566400, 1410570000, 1410573600, 
    1410577200, 1410580800, 1410584400, 1410588000, 1410591600, 1410595200, 
    1410598800, 1410602400, 1410606000, 1410609600, 1410613200, 1410616800, 
    1410620400, 1410624000, 1410627600, 1410631200, 1410634800, 1410638400, 
    1410642000, 1410645600, 1410649200, 1410652800, 1410656400, 1410660000, 
    1410663600, 1410667200, 1410670800, 1410674400, 1410678000, 1410681600, 
    1410685200, 1410688800, 1410692400, 1410696000, 1410699600, 1410703200, 
    1410706800, 1410710400, 1410714000, 1410717600, 1410721200, 1410724800, 
    1410728400, 1410732000, 1410735600, 1410739200, 1410742800, 1410746400, 
    1410750000, 1410753600, 1410757200, 1410760800, 1410764400, 1410768000, 
    1410771600, 1410775200, 1410778800, 1410782400, 1410786000, 1410789600, 
    1410793200, 1410796800, 1410800400, 1410804000, 1410807600, 1410811200, 
    1410814800, 1410818400, 1410822000, 1410825600, 1410829200, 1410832800, 
    1410836400, 1410840000, 1410843600, 1410847200, 1410850800, 1410854400, 
    1410858000, 1410861600, 1410865200, 1410868800, 1410872400, 1410876000, 
    1410879600, 1410883200, 1410886800, 1410890400, 1410894000, 1410897600, 
    1410901200, 1410904800, 1410908400, 1410912000, 1410915600, 1410919200, 
    1410922800, 1410926400, 1410930000, 1410933600, 1410937200, 1410940800, 
    1410944400, 1410948000, 1410951600, 1410955200, 1410958800, 1410962400, 
    1410966000, 1410969600, 1410973200, 1410976800, 1410980400, 1410984000, 
    1410987600, 1410991200, 1410994800, 1410998400, 1411002000, 1411005600, 
    1411009200, 1411012800, 1411016400, 1411020000, 1411023600, 1411027200, 
    1411030800, 1411034400, 1411038000, 1411041600, 1411045200, 1411048800, 
    1411052400, 1411056000, 1411059600, 1411063200, 1411066800, 1411070400, 
    1411074000, 1411077600, 1411081200, 1411084800, 1411088400, 1411092000, 
    1411095600, 1411099200, 1411102800, 1411106400, 1411110000, 1411113600, 
    1411117200, 1411120800, 1411124400, 1411128000, 1411131600, 1411135200, 
    1411138800, 1411142400, 1411146000, 1411149600, 1411153200, 1411156800, 
    1411160400, 1411164000, 1411167600, 1411171200, 1411174800, 1411178400, 
    1411182000, 1411185600, 1411189200, 1411192800, 1411196400, 1411200000, 
    1411203600, 1411207200, 1411210800, 1411214400, 1411218000, 1411221600, 
    1411225200, 1411228800, 1411232400, 1411236000, 1411239600, 1411243200, 
    1411246800, 1411250400, 1411254000, 1411257600, 1411261200, 1411264800, 
    1411268400, 1411272000, 1411275600, 1411279200, 1411282800, 1411286400, 
    1411290000, 1411293600, 1411297200, 1411300800, 1411304400, 1411308000, 
    1411311600, 1411315200, 1411318800, 1411322400, 1411326000, 1411329600, 
    1411333200, 1411336800, 1411340400, 1411344000, 1411347600, 1411351200, 
    1411354800, 1411358400, 1411362000, 1411365600, 1411369200, 1411372800, 
    1411376400, 1411380000, 1411383600, 1411387200, 1411390800, 1411394400, 
    1411398000, 1411401600, 1411405200, 1411408800, 1411412400, 1411416000, 
    1411419600, 1411423200, 1411426800, 1411430400, 1411434000, 1411437600, 
    1411441200, 1411444800, 1411448400, 1411452000, 1411455600, 1411459200, 
    1411462800, 1411466400, 1411470000, 1411473600, 1411477200, 1411480800, 
    1411484400, 1411488000, 1411491600, 1411495200, 1411498800, 1411502400, 
    1411506000, 1411509600, 1411513200, 1411516800, 1411520400, 1411524000, 
    1411527600, 1411531200, 1411534800, 1411538400, 1411542000, 1411545600, 
    1411549200, 1411552800, 1411556400, 1411560000, 1411563600, 1411567200, 
    1411570800, 1411574400, 1411578000, 1411581600, 1411585200, 1411588800, 
    1411592400, 1411596000, 1411599600, 1411603200, 1411606800, 1411610400, 
    1411614000, 1411617600, 1411621200, 1411624800, 1411628400, 1411632000, 
    1411635600, 1411639200, 1411642800, 1411646400, 1411650000, 1411653600, 
    1411657200, 1411660800, 1411664400, 1411668000, 1411671600, 1411675200, 
    1411678800, 1411682400, 1411686000, 1411689600, 1411693200, 1411696800, 
    1411700400, 1411704000, 1411707600, 1411711200, 1411714800, 1411718400, 
    1411722000, 1411725600, 1411729200, 1411732800, 1411736400, 1411740000, 
    1411743600, 1411747200, 1411750800, 1411754400, 1411758000, 1411761600, 
    1411765200, 1411768800, 1411772400, 1411776000, 1411779600, 1411783200, 
    1411786800, 1411790400, 1411794000, 1411797600, 1411801200, 1411804800, 
    1411808400, 1411812000, 1411815600, 1411819200, 1411822800, 1411826400, 
    1411830000, 1411833600, 1411837200, 1411840800, 1411844400, 1411848000, 
    1411851600, 1411855200, 1411858800, 1411862400, 1411866000, 1411869600, 
    1411873200, 1411876800, 1411880400, 1411884000, 1411887600, 1411891200, 
    1411894800, 1411898400, 1411902000, 1411905600, 1411909200, 1411912800, 
    1411916400, 1411920000, 1411923600, 1411927200, 1411930800, 1411934400, 
    1411938000, 1411941600, 1411945200, 1411948800, 1411952400, 1411956000, 
    1411959600, 1411963200, 1411966800, 1411970400, 1411974000, 1411977600, 
    1411981200, 1411984800, 1411988400, 1411992000, 1411995600, 1411999200, 
    1412002800, 1412006400, 1412010000, 1412013600, 1412017200, 1412020800, 
    1412024400, 1412028000, 1412031600, 1412035200, 1412038800, 1412042400, 
    1412046000, 1412049600, 1412053200, 1412056800, 1412060400, 1412064000, 
    1412067600, 1412071200, 1412074800, 1412078400, 1412082000, 1412085600, 
    1412089200, 1412092800, 1412096400, 1412100000, 1412103600, 1412107200, 
    1412110800, 1412114400, 1412118000, 1412121600, 1412125200, 1412128800, 
    1412132400, 1412136000, 1412139600, 1412143200, 1412146800, 1412150400, 
    1412154000, 1412157600, 1412161200, 1412164800, 1412168400, 1412172000, 
    1412175600, 1412179200, 1412182800, 1412186400, 1412190000, 1412193600, 
    1412197200, 1412200800, 1412204400, 1412208000, 1412211600, 1412215200, 
    1412218800, 1412222400, 1412226000, 1412229600, 1412233200, 1412236800, 
    1412240400, 1412244000, 1412247600, 1412251200, 1412254800, 1412258400, 
    1412262000, 1412265600, 1412269200, 1412272800, 1412276400, 1412280000, 
    1412283600, 1412287200, 1412290800, 1412294400, 1412298000, 1412301600, 
    1412305200, 1412308800, 1412312400, 1412316000, 1412319600, 1412323200, 
    1412326800, 1412330400, 1412334000, 1412337600, 1412341200, 1412344800, 
    1412348400, 1412352000, 1412355600, 1412359200, 1412362800, 1412366400, 
    1412370000, 1412373600, 1412377200, 1412380800, 1412384400, 1412388000, 
    1412391600, 1412395200, 1412398800, 1412402400, 1412406000, 1412409600, 
    1412413200, 1412416800, 1412420400, 1412424000, 1412427600, 1412431200, 
    1412434800, 1412438400, 1412442000, 1412445600, 1412449200, 1412452800, 
    1412456400, 1412460000, 1412463600, 1412467200, 1412470800, 1412474400, 
    1412478000, 1412481600, 1412485200, 1412488800, 1412492400, 1412496000, 
    1412499600, 1412503200, 1412506800, 1412510400, 1412514000, 1412517600, 
    1412521200, 1412524800, 1412528400, 1412532000, 1412535600, 1412539200, 
    1412542800, 1412546400, 1412550000, 1412553600, 1412557200, 1412560800, 
    1412564400, 1412568000, 1412571600, 1412575200, 1412578800, 1412582400, 
    1412586000, 1412589600, 1412593200, 1412596800, 1412600400, 1412604000, 
    1412607600, 1412611200, 1412614800, 1412618400, 1412622000, 1412625600, 
    1412629200, 1412632800, 1412636400, 1412640000, 1412643600, 1412647200, 
    1412650800, 1412654400, 1412658000, 1412661600, 1412665200, 1412668800, 
    1412672400, 1412676000, 1412679600, 1412683200, 1412686800, 1412690400, 
    1412694000, 1412697600, 1412701200, 1412704800, 1412708400, 1412712000, 
    1412715600, 1412719200, 1412722800, 1412726400, 1412730000, 1412733600, 
    1412737200, 1412740800, 1412744400, 1412748000, 1412751600, 1412755200, 
    1412758800, 1412762400, 1412766000, 1412769600, 1412773200, 1412776800, 
    1412780400, 1412784000, 1412787600, 1412791200, 1412794800, 1412798400, 
    1412802000, 1412805600, 1412809200, 1412812800, 1412816400, 1412820000, 
    1412823600, 1412827200, 1412830800, 1412834400, 1412838000, 1412841600, 
    1412845200, 1412848800, 1412852400, 1412856000, 1412859600, 1412863200, 
    1412866800, 1412870400, 1412874000, 1412877600, 1412881200, 1412884800, 
    1412888400, 1412892000, 1412895600, 1412899200, 1412902800, 1412906400, 
    1412910000, 1412913600, 1412917200, 1412920800, 1412924400, 1412928000, 
    1412931600, 1412935200, 1412938800, 1412942400, 1412946000, 1412949600, 
    1412953200, 1412956800, 1412960400, 1412964000, 1412967600, 1412971200, 
    1412974800, 1412978400, 1412982000, 1412985600, 1412989200, 1412992800, 
    1412996400, 1413000000, 1413003600, 1413007200, 1413010800, 1413014400, 
    1413018000, 1413021600, 1413025200, 1413028800, 1413032400, 1413036000, 
    1413039600, 1413043200, 1413046800, 1413050400, 1413054000, 1413057600, 
    1413061200, 1413064800, 1413068400, 1413072000, 1413075600, 1413079200, 
    1413082800, 1413086400, 1413090000, 1413093600, 1413097200, 1413100800, 
    1413104400, 1413108000, 1413111600, 1413115200, 1413118800, 1413122400, 
    1413126000, 1413129600, 1413133200, 1413136800, 1413140400, 1413144000, 
    1413147600, 1413151200, 1413154800, 1413158400, 1413162000, 1413165600, 
    1413169200, 1413172800, 1413176400, 1413180000, 1413183600, 1413187200, 
    1413190800, 1413194400, 1413198000, 1413201600, 1413205200, 1413208800, 
    1413212400, 1413216000, 1413219600, 1413223200, 1413226800, 1413230400, 
    1413234000, 1413237600, 1413241200, 1413244800, 1413248400, 1413252000, 
    1413255600, 1413259200, 1413262800, 1413266400, 1413270000, 1413273600, 
    1413277200, 1413280800, 1413284400, 1413288000, 1413291600, 1413295200, 
    1413298800, 1413302400, 1413306000, 1413309600, 1413313200, 1413316800, 
    1413320400, 1413324000, 1413327600, 1413331200, 1413334800, 1413338400, 
    1413342000, 1413345600, 1413349200, 1413352800, 1413356400, 1413360000, 
    1413363600, 1413367200, 1413370800, 1413374400, 1413378000, 1413381600, 
    1413385200, 1413388800, 1413392400, 1413396000, 1413399600, 1413403200, 
    1413406800, 1413410400, 1413414000, 1413417600, 1413421200, 1413424800, 
    1413428400, 1413432000, 1413435600, 1413439200, 1413442800, 1413446400, 
    1413450000, 1413453600, 1413457200, 1413460800, 1413464400, 1413468000, 
    1413471600, 1413475200, 1413478800, 1413482400, 1413486000, 1413489600, 
    1413493200, 1413496800, 1413500400, 1413504000, 1413507600, 1413511200, 
    1413514800, 1413518400, 1413522000, 1413525600, 1413529200, 1413532800, 
    1413536400, 1413540000, 1413543600, 1413547200, 1413550800, 1413554400, 
    1413558000, 1413561600, 1413565200, 1413568800, 1413572400, 1413576000, 
    1413579600, 1413583200, 1413586800, 1413590400, 1413594000, 1413597600, 
    1413601200, 1413604800, 1413608400, 1413612000, 1413615600, 1413619200, 
    1413622800, 1413626400, 1413630000, 1413633600, 1413637200, 1413640800, 
    1413644400, 1413648000, 1413651600, 1413655200, 1413658800, 1413662400, 
    1413666000, 1413669600, 1413673200, 1413676800, 1413680400, 1413684000, 
    1413687600, 1413691200, 1413694800, 1413698400, 1413702000, 1413705600, 
    1413709200, 1413712800, 1413716400, 1413720000, 1413723600, 1413727200, 
    1413730800, 1413734400, 1413738000, 1413741600, 1413745200, 1413748800, 
    1413752400, 1413756000, 1413759600, 1413763200, 1413766800, 1413770400, 
    1413774000, 1413777600, 1413781200, 1413784800, 1413788400, 1413792000, 
    1413795600, 1413799200, 1413802800, 1413806400, 1413810000, 1413813600, 
    1413817200, 1413820800, 1413824400, 1413828000, 1413831600, 1413835200, 
    1413838800, 1413842400, 1413846000, 1413849600, 1413853200, 1413856800, 
    1413860400, 1413864000, 1413867600, 1413871200, 1413874800, 1413878400, 
    1413882000, 1413885600, 1413889200, 1413892800, 1413896400, 1413900000, 
    1413903600, 1413907200, 1413910800, 1413914400, 1413918000, 1413921600, 
    1413925200, 1413928800, 1413932400, 1413936000, 1413939600, 1413943200, 
    1413946800, 1413950400, 1413954000, 1413957600, 1413961200, 1413964800, 
    1413968400, 1413972000, 1413975600, 1413979200, 1413982800, 1413986400, 
    1413990000, 1413993600, 1413997200, 1414000800, 1414004400, 1414008000, 
    1414011600, 1414015200, 1414018800, 1414022400, 1414026000, 1414029600, 
    1414033200, 1414036800, 1414040400, 1414044000, 1414047600, 1414051200, 
    1414054800, 1414058400, 1414062000, 1414065600, 1414069200, 1414072800, 
    1414076400, 1414080000, 1414083600, 1414087200, 1414090800, 1414094400, 
    1414098000, 1414101600, 1414105200, 1414108800, 1414112400, 1414116000, 
    1414119600, 1414123200, 1414126800, 1414130400, 1414134000, 1414137600, 
    1414141200, 1414144800, 1414148400, 1414152000, 1414155600, 1414159200, 
    1414162800, 1414166400, 1414170000, 1414173600, 1414177200, 1414180800, 
    1414184400, 1414188000, 1414191600, 1414195200, 1414198800, 1414202400, 
    1414206000, 1414209600, 1414213200, 1414216800, 1414220400, 1414224000, 
    1414227600, 1414231200, 1414234800, 1414238400, 1414242000, 1414245600, 
    1414249200, 1414252800, 1414256400, 1414260000, 1414263600, 1414267200, 
    1414270800, 1414274400, 1414278000, 1414281600, 1414285200, 1414288800, 
    1414292400, 1414296000, 1414299600, 1414303200, 1414306800, 1414310400, 
    1414314000, 1414317600, 1414321200, 1414324800, 1414328400, 1414332000, 
    1414335600, 1414339200, 1414342800, 1414346400, 1414350000, 1414353600, 
    1414357200, 1414360800, 1414364400, 1414368000, 1414371600, 1414375200, 
    1414378800, 1414382400, 1414386000, 1414389600, 1414393200, 1414396800, 
    1414400400, 1414404000, 1414407600, 1414411200, 1414414800, 1414418400, 
    1414422000, 1414425600, 1414429200, 1414432800, 1414436400, 1414440000, 
    1414443600, 1414447200, 1414450800, 1414454400, 1414458000, 1414461600, 
    1414465200, 1414468800, 1414472400, 1414476000, 1414479600, 1414483200, 
    1414486800, 1414490400, 1414494000, 1414497600, 1414501200, 1414504800, 
    1414508400, 1414512000, 1414515600, 1414519200, 1414522800, 1414526400, 
    1414530000, 1414533600, 1414537200, 1414540800, 1414544400, 1414548000, 
    1414551600, 1414555200, 1414558800, 1414562400, 1414566000, 1414569600, 
    1414573200, 1414576800, 1414580400, 1414584000, 1414587600, 1414591200, 
    1414594800, 1414598400, 1414602000, 1414605600, 1414609200, 1414612800, 
    1414616400, 1414620000, 1414623600, 1414627200, 1414630800, 1414634400, 
    1414638000, 1414641600, 1414645200, 1414648800, 1414652400, 1414656000, 
    1414659600, 1414663200, 1414666800, 1414670400, 1414674000, 1414677600, 
    1414681200, 1414684800, 1414688400, 1414692000, 1414695600, 1414699200, 
    1414702800, 1414706400, 1414710000, 1414713600, 1414717200, 1414720800, 
    1414724400, 1414728000, 1414731600, 1414735200, 1414738800, 1414742400, 
    1414746000, 1414749600, 1414753200, 1414756800, 1414760400, 1414764000, 
    1414767600, 1414771200, 1414774800, 1414778400, 1414782000, 1414785600, 
    1414789200, 1414792800, 1414796400, 1414800000, 1414803600, 1414807200, 
    1414810800, 1414814400, 1414818000, 1414821600, 1414825200, 1414828800, 
    1414832400, 1414836000, 1414839600, 1414843200, 1414846800, 1414850400, 
    1414854000, 1414857600, 1414861200, 1414864800, 1414868400, 1414872000, 
    1414875600, 1414879200, 1414882800, 1414886400, 1414890000, 1414893600, 
    1414897200, 1414900800, 1414904400, 1414908000, 1414911600, 1414915200, 
    1414918800, 1414922400, 1414926000, 1414929600, 1414933200, 1414936800, 
    1414940400, 1414944000, 1414947600, 1414951200, 1414954800, 1414958400, 
    1414962000, 1414965600, 1414969200, 1414972800, 1414976400, 1414980000, 
    1414983600, 1414987200, 1414990800, 1414994400, 1414998000, 1415001600, 
    1415005200, 1415008800, 1415012400, 1415016000, 1415019600, 1415023200, 
    1415026800, 1415030400, 1415034000, 1415037600, 1415041200, 1415044800, 
    1415048400, 1415052000, 1415055600, 1415059200, 1415062800, 1415066400, 
    1415070000, 1415073600, 1415077200, 1415080800, 1415084400, 1415088000, 
    1415091600, 1415095200, 1415098800, 1415102400, 1415106000, 1415109600, 
    1415113200, 1415116800, 1415120400, 1415124000, 1415127600, 1415131200, 
    1415134800, 1415138400, 1415142000, 1415145600, 1415149200, 1415152800, 
    1415156400, 1415160000, 1415163600, 1415167200, 1415170800, 1415174400, 
    1415178000, 1415181600, 1415185200, 1415188800, 1415192400, 1415196000, 
    1415199600, 1415203200, 1415206800, 1415210400, 1415214000, 1415217600, 
    1415221200, 1415224800, 1415228400, 1415232000, 1415235600, 1415239200, 
    1415242800, 1415246400, 1415250000, 1415253600, 1415257200, 1415260800, 
    1415264400, 1415268000, 1415271600, 1415275200, 1415278800, 1415282400, 
    1415286000, 1415289600, 1415293200, 1415296800, 1415300400, 1415304000, 
    1415307600, 1415311200, 1415314800, 1415318400, 1415322000, 1415325600, 
    1415329200, 1415332800, 1415336400, 1415340000, 1415343600, 1415347200, 
    1415350800, 1415354400, 1415358000, 1415361600, 1415365200, 1415368800, 
    1415372400, 1415376000, 1415379600, 1415383200, 1415386800, 1415390400, 
    1415394000, 1415397600, 1415401200, 1415404800, 1415408400, 1415412000, 
    1415415600, 1415419200, 1415422800, 1415426400, 1415430000, 1415433600, 
    1415437200, 1415440800, 1415444400, 1415448000, 1415451600, 1415455200, 
    1415458800, 1415462400, 1415466000, 1415469600, 1415473200, 1415476800, 
    1415480400, 1415484000, 1415487600, 1415491200, 1415494800, 1415498400, 
    1415502000, 1415505600, 1415509200, 1415512800, 1415516400, 1415520000, 
    1415523600, 1415527200, 1415530800, 1415534400, 1415538000, 1415541600, 
    1415545200, 1415548800, 1415552400, 1415556000, 1415559600, 1415563200, 
    1415566800, 1415570400, 1415574000, 1415577600, 1415581200, 1415584800, 
    1415588400, 1415592000, 1415595600, 1415599200, 1415602800, 1415606400, 
    1415610000, 1415613600, 1415617200, 1415620800, 1415624400, 1415628000, 
    1415631600, 1415635200, 1415638800, 1415642400, 1415646000, 1415649600, 
    1415653200, 1415656800, 1415660400, 1415664000, 1415667600, 1415671200, 
    1415674800, 1415678400, 1415682000, 1415685600, 1415689200, 1415692800, 
    1415696400, 1415700000, 1415703600, 1415707200, 1415710800, 1415714400, 
    1415718000, 1415721600, 1415725200, 1415728800, 1415732400, 1415736000, 
    1415739600, 1415743200, 1415746800, 1415750400, 1415754000, 1415757600, 
    1415761200, 1415764800, 1415768400, 1415772000, 1415775600, 1415779200, 
    1415782800, 1415786400, 1415790000, 1415793600, 1415797200, 1415800800, 
    1415804400, 1415808000, 1415811600, 1415815200, 1415818800, 1415822400, 
    1415826000, 1415829600, 1415833200, 1415836800, 1415840400, 1415844000, 
    1415847600, 1415851200, 1415854800, 1415858400, 1415862000, 1415865600, 
    1415869200, 1415872800, 1415876400, 1415880000, 1415883600, 1415887200, 
    1415890800, 1415894400, 1415898000, 1415901600, 1415905200, 1415908800, 
    1415912400, 1415916000, 1415919600, 1415923200, 1415926800, 1415930400, 
    1415934000, 1415937600, 1415941200, 1415944800, 1415948400, 1415952000, 
    1415955600, 1415959200, 1415962800, 1415966400, 1415970000, 1415973600, 
    1415977200, 1415980800, 1415984400, 1415988000, 1415991600, 1415995200, 
    1415998800, 1416002400, 1416006000, 1416009600, 1416013200, 1416016800, 
    1416020400, 1416024000, 1416027600, 1416031200, 1416034800, 1416038400, 
    1416042000, 1416045600, 1416049200, 1416052800, 1416056400, 1416060000, 
    1416063600, 1416067200, 1416070800, 1416074400, 1416078000, 1416081600, 
    1416085200, 1416088800, 1416092400, 1416096000, 1416099600, 1416103200, 
    1416106800, 1416110400, 1416114000, 1416117600, 1416121200, 1416124800, 
    1416128400, 1416132000, 1416135600, 1416139200, 1416142800, 1416146400, 
    1416150000, 1416153600, 1416157200, 1416160800, 1416164400, 1416168000, 
    1416171600, 1416175200, 1416178800, 1416182400, 1416186000, 1416189600, 
    1416193200, 1416196800, 1416200400, 1416204000, 1416207600, 1416211200, 
    1416214800, 1416218400, 1416222000, 1416225600, 1416229200, 1416232800, 
    1416236400, 1416240000, 1416243600, 1416247200, 1416250800, 1416254400, 
    1416258000, 1416261600, 1416265200, 1416268800, 1416272400, 1416276000, 
    1416279600, 1416283200, 1416286800, 1416290400, 1416294000, 1416297600, 
    1416301200, 1416304800, 1416308400, 1416312000, 1416315600, 1416319200, 
    1416322800, 1416326400, 1416330000, 1416333600, 1416337200, 1416340800, 
    1416344400, 1416348000, 1416351600, 1416355200, 1416358800, 1416362400, 
    1416366000, 1416369600, 1416373200, 1416376800, 1416380400, 1416384000, 
    1416387600, 1416391200, 1416394800, 1416398400, 1416402000, 1416405600, 
    1416409200, 1416412800, 1416416400, 1416420000, 1416423600, 1416427200, 
    1416430800, 1416434400, 1416438000, 1416441600, 1416445200, 1416448800, 
    1416452400, 1416456000, 1416459600, 1416463200, 1416466800, 1416470400, 
    1416474000, 1416477600, 1416481200, 1416484800, 1416488400, 1416492000, 
    1416495600, 1416499200, 1416502800, 1416506400, 1416510000, 1416513600, 
    1416517200, 1416520800, 1416524400, 1416528000, 1416531600, 1416535200, 
    1416538800, 1416542400, 1416546000, 1416549600, 1416553200, 1416556800, 
    1416560400, 1416564000, 1416567600, 1416571200, 1416574800, 1416578400, 
    1416582000, 1416585600, 1416589200, 1416592800, 1416596400, 1416600000, 
    1416603600, 1416607200, 1416610800, 1416614400, 1416618000, 1416621600, 
    1416625200, 1416628800, 1416632400, 1416636000, 1416639600, 1416643200, 
    1416646800, 1416650400, 1416654000, 1416657600, 1416661200, 1416664800, 
    1416668400, 1416672000, 1416675600, 1416679200, 1416682800, 1416686400, 
    1416690000, 1416693600, 1416697200, 1416700800, 1416704400, 1416708000, 
    1416711600, 1416715200, 1416718800, 1416722400, 1416726000, 1416729600, 
    1416733200, 1416736800, 1416740400, 1416744000, 1416747600, 1416751200, 
    1416754800, 1416758400, 1416762000, 1416765600, 1416769200, 1416772800, 
    1416776400, 1416780000, 1416783600, 1416787200, 1416790800, 1416794400, 
    1416798000, 1416801600, 1416805200, 1416808800, 1416812400, 1416816000, 
    1416819600, 1416823200, 1416826800, 1416830400, 1416834000, 1416837600, 
    1416841200, 1416844800, 1416848400, 1416852000, 1416855600, 1416859200, 
    1416862800, 1416866400, 1416870000, 1416873600, 1416877200, 1416880800, 
    1416884400, 1416888000, 1416891600, 1416895200, 1416898800, 1416902400, 
    1416906000, 1416909600, 1416913200, 1416916800, 1416920400, 1416924000, 
    1416927600, 1416931200, 1416934800, 1416938400, 1416942000, 1416945600, 
    1416949200, 1416952800, 1416956400, 1416960000, 1416963600, 1416967200, 
    1416970800, 1416974400, 1416978000, 1416981600, 1416985200, 1416988800, 
    1416992400, 1416996000, 1416999600, 1417003200, 1417006800, 1417010400, 
    1417014000, 1417017600, 1417021200, 1417024800, 1417028400, 1417032000, 
    1417035600, 1417039200, 1417042800, 1417046400, 1417050000, 1417053600, 
    1417057200, 1417060800, 1417064400, 1417068000, 1417071600, 1417075200, 
    1417078800, 1417082400, 1417086000, 1417089600, 1417093200, 1417096800, 
    1417100400, 1417104000, 1417107600, 1417111200, 1417114800, 1417118400, 
    1417122000, 1417125600, 1417129200, 1417132800, 1417136400, 1417140000, 
    1417143600, 1417147200, 1417150800, 1417154400, 1417158000, 1417161600, 
    1417165200, 1417168800, 1417172400, 1417176000, 1417179600, 1417183200, 
    1417186800, 1417190400, 1417194000, 1417197600, 1417201200, 1417204800, 
    1417208400, 1417212000, 1417215600, 1417219200, 1417222800, 1417226400, 
    1417230000, 1417233600, 1417237200, 1417240800, 1417244400, 1417248000, 
    1417251600, 1417255200, 1417258800, 1417262400, 1417266000, 1417269600, 
    1417273200, 1417276800, 1417280400, 1417284000, 1417287600, 1417291200, 
    1417294800, 1417298400, 1417302000, 1417305600, 1417309200, 1417312800, 
    1417316400, 1417320000, 1417323600, 1417327200, 1417330800, 1417334400, 
    1417338000, 1417341600, 1417345200, 1417348800, 1417352400, 1417356000, 
    1417359600, 1417363200, 1417366800, 1417370400, 1417374000, 1417377600, 
    1417381200, 1417384800, 1417388400, 1417392000, 1417395600, 1417399200, 
    1417402800, 1417406400, 1417410000, 1417413600, 1417417200, 1417420800, 
    1417424400, 1417428000, 1417431600, 1417435200, 1417438800, 1417442400, 
    1417446000, 1417449600, 1417453200, 1417456800, 1417460400, 1417464000, 
    1417467600, 1417471200, 1417474800, 1417478400, 1417482000, 1417485600, 
    1417489200, 1417492800, 1417496400, 1417500000, 1417503600, 1417507200, 
    1417510800, 1417514400, 1417518000, 1417521600, 1417525200, 1417528800, 
    1417532400, 1417536000, 1417539600, 1417543200, 1417546800, 1417550400, 
    1417554000, 1417557600, 1417561200, 1417564800, 1417568400, 1417572000, 
    1417575600, 1417579200, 1417582800, 1417586400, 1417590000, 1417593600, 
    1417597200, 1417600800, 1417604400, 1417608000, 1417611600, 1417615200, 
    1417618800, 1417622400, 1417626000, 1417629600, 1417633200, 1417636800, 
    1417640400, 1417644000, 1417647600, 1417651200, 1417654800, 1417658400, 
    1417662000, 1417665600, 1417669200, 1417672800, 1417676400, 1417680000, 
    1417683600, 1417687200, 1417690800, 1417694400, 1417698000, 1417701600, 
    1417705200, 1417708800, 1417712400, 1417716000, 1417719600, 1417723200, 
    1417726800, 1417730400, 1417734000, 1417737600, 1417741200, 1417744800, 
    1417748400, 1417752000, 1417755600, 1417759200, 1417762800, 1417766400, 
    1417770000, 1417773600, 1417777200, 1417780800, 1417784400, 1417788000, 
    1417791600, 1417795200, 1417798800, 1417802400, 1417806000, 1417809600, 
    1417813200, 1417816800, 1417820400, 1417824000, 1417827600, 1417831200, 
    1417834800, 1417838400, 1417842000, 1417845600, 1417849200, 1417852800, 
    1417856400, 1417860000, 1417863600, 1417867200, 1417870800, 1417874400, 
    1417878000, 1417881600, 1417885200, 1417888800, 1417892400, 1417896000, 
    1417899600, 1417903200, 1417906800, 1417910400, 1417914000, 1417917600, 
    1417921200, 1417924800, 1417928400, 1417932000, 1417935600, 1417939200, 
    1417942800, 1417946400, 1417950000, 1417953600, 1417957200, 1417960800, 
    1417964400, 1417968000, 1417971600, 1417975200, 1417978800, 1417982400, 
    1417986000, 1417989600, 1417993200, 1417996800, 1418000400, 1418004000, 
    1418007600, 1418011200, 1418014800, 1418018400, 1418022000, 1418025600, 
    1418029200, 1418032800, 1418036400, 1418040000, 1418043600, 1418047200, 
    1418050800, 1418054400, 1418058000, 1418061600, 1418065200, 1418068800, 
    1418072400, 1418076000, 1418079600, 1418083200, 1418086800, 1418090400, 
    1418094000, 1418097600, 1418101200, 1418104800, 1418108400, 1418112000, 
    1418115600, 1418119200, 1418122800, 1418126400, 1418130000, 1418133600, 
    1418137200, 1418140800, 1418144400, 1418148000, 1418151600, 1418155200, 
    1418158800, 1418162400, 1418166000, 1418169600, 1418173200, 1418176800, 
    1418180400, 1418184000, 1418187600, 1418191200, 1418194800, 1418198400, 
    1418202000, 1418205600, 1418209200, 1418212800, 1418216400, 1418220000, 
    1418223600, 1418227200, 1418230800, 1418234400, 1418238000, 1418241600, 
    1418245200, 1418248800, 1418252400, 1418256000, 1418259600, 1418263200, 
    1418266800, 1418270400, 1418274000, 1418277600, 1418281200, 1418284800, 
    1418288400, 1418292000, 1418295600, 1418299200, 1418302800, 1418306400, 
    1418310000, 1418313600, 1418317200, 1418320800, 1418324400, 1418328000, 
    1418331600, 1418335200, 1418338800, 1418342400, 1418346000, 1418349600, 
    1418353200, 1418356800, 1418360400, 1418364000, 1418367600, 1418371200, 
    1418374800, 1418378400, 1418382000, 1418385600, 1418389200, 1418392800, 
    1418396400, 1418400000, 1418403600, 1418407200, 1418410800, 1418414400, 
    1418418000, 1418421600, 1418425200, 1418428800, 1418432400, 1418436000, 
    1418439600, 1418443200, 1418446800, 1418450400, 1418454000, 1418457600, 
    1418461200, 1418464800, 1418468400, 1418472000, 1418475600, 1418479200, 
    1418482800, 1418486400, 1418490000, 1418493600, 1418497200, 1418500800, 
    1418504400, 1418508000, 1418511600, 1418515200, 1418518800, 1418522400, 
    1418526000, 1418529600, 1418533200, 1418536800, 1418540400, 1418544000, 
    1418547600, 1418551200, 1418554800, 1418558400, 1418562000, 1418565600, 
    1418569200, 1418572800, 1418576400, 1418580000, 1418583600, 1418587200, 
    1418590800, 1418594400, 1418598000, 1418601600, 1418605200, 1418608800, 
    1418612400, 1418616000, 1418619600, 1418623200, 1418626800, 1418630400, 
    1418634000, 1418637600, 1418641200, 1418644800, 1418648400, 1418652000, 
    1418655600, 1418659200, 1418662800, 1418666400, 1418670000, 1418673600, 
    1418677200, 1418680800, 1418684400, 1418688000, 1418691600, 1418695200, 
    1418698800, 1418702400, 1418706000, 1418709600, 1418713200, 1418716800, 
    1418720400, 1418724000, 1418727600, 1418731200, 1418734800, 1418738400, 
    1418742000, 1418745600, 1418749200, 1418752800, 1418756400, 1418760000, 
    1418763600, 1418767200, 1418770800, 1418774400, 1418778000, 1418781600, 
    1418785200, 1418788800, 1418792400, 1418796000, 1418799600, 1418803200, 
    1418806800, 1418810400, 1418814000, 1418817600, 1418821200, 1418824800, 
    1418828400, 1418832000, 1418835600, 1418839200, 1418842800, 1418846400, 
    1418850000, 1418853600, 1418857200, 1418860800, 1418864400, 1418868000, 
    1418871600, 1418875200, 1418878800, 1418882400, 1418886000, 1418889600, 
    1418893200, 1418896800, 1418900400, 1418904000, 1418907600, 1418911200, 
    1418914800, 1418918400, 1418922000, 1418925600, 1418929200, 1418932800, 
    1418936400, 1418940000, 1418943600, 1418947200, 1418950800, 1418954400, 
    1418958000, 1418961600, 1418965200, 1418968800, 1418972400, 1418976000, 
    1418979600, 1418983200, 1418986800, 1418990400, 1418994000, 1418997600, 
    1419001200, 1419004800, 1419008400, 1419012000, 1419015600, 1419019200, 
    1419022800, 1419026400, 1419030000, 1419033600, 1419037200, 1419040800, 
    1419044400, 1419048000, 1419051600, 1419055200, 1419058800, 1419062400, 
    1419066000, 1419069600, 1419073200, 1419076800, 1419080400, 1419084000, 
    1419087600, 1419091200, 1419094800, 1419098400, 1419102000, 1419105600, 
    1419109200, 1419112800, 1419116400, 1419120000, 1419123600, 1419127200, 
    1419130800, 1419134400, 1419138000, 1419141600, 1419145200, 1419148800, 
    1419152400, 1419156000, 1419159600, 1419163200, 1419166800, 1419170400, 
    1419174000, 1419177600, 1419181200, 1419184800, 1419188400, 1419192000, 
    1419195600, 1419199200, 1419202800, 1419206400, 1419210000, 1419213600, 
    1419217200, 1419220800, 1419224400, 1419228000, 1419231600, 1419235200, 
    1419238800, 1419242400, 1419246000, 1419249600, 1419253200, 1419256800, 
    1419260400, 1419264000, 1419267600, 1419271200, 1419274800, 1419278400, 
    1419282000, 1419285600, 1419289200, 1419292800, 1419296400, 1419300000, 
    1419303600, 1419307200, 1419310800, 1419314400, 1419318000, 1419321600, 
    1419325200, 1419328800, 1419332400, 1419336000, 1419339600, 1419343200, 
    1419346800, 1419350400, 1419354000, 1419357600, 1419361200, 1419364800, 
    1419368400, 1419372000, 1419375600, 1419379200, 1419382800, 1419386400, 
    1419390000, 1419393600, 1419397200, 1419400800, 1419404400, 1419408000, 
    1419411600, 1419415200, 1419418800, 1419422400, 1419426000, 1419429600, 
    1419433200, 1419436800, 1419440400, 1419444000, 1419447600, 1419451200, 
    1419454800, 1419458400, 1419462000, 1419465600, 1419469200, 1419472800, 
    1419476400, 1419480000, 1419483600, 1419487200, 1419490800, 1419494400, 
    1419498000, 1419501600, 1419505200, 1419508800, 1419512400, 1419516000, 
    1419519600, 1419523200, 1419526800, 1419530400, 1419534000, 1419537600, 
    1419541200, 1419544800, 1419548400, 1419552000, 1419555600, 1419559200, 
    1419562800, 1419566400, 1419570000, 1419573600, 1419577200, 1419580800, 
    1419584400, 1419588000, 1419591600, 1419595200, 1419598800, 1419602400, 
    1419606000, 1419609600, 1419613200, 1419616800, 1419620400, 1419624000, 
    1419627600, 1419631200, 1419634800, 1419638400, 1419642000, 1419645600, 
    1419649200, 1419652800, 1419656400, 1419660000, 1419663600, 1419667200, 
    1419670800, 1419674400, 1419678000, 1419681600, 1419685200, 1419688800, 
    1419692400, 1419696000, 1419699600, 1419703200, 1419706800, 1419710400, 
    1419714000, 1419717600, 1419721200, 1419724800, 1419728400, 1419732000, 
    1419735600, 1419739200, 1419742800, 1419746400, 1419750000, 1419753600, 
    1419757200, 1419760800, 1419764400, 1419768000, 1419771600, 1419775200, 
    1419778800, 1419782400, 1419786000, 1419789600, 1419793200, 1419796800, 
    1419800400, 1419804000, 1419807600, 1419811200, 1419814800, 1419818400, 
    1419822000, 1419825600, 1419829200, 1419832800, 1419836400, 1419840000, 
    1419843600, 1419847200, 1419850800, 1419854400, 1419858000, 1419861600, 
    1419865200, 1419868800, 1419872400, 1419876000, 1419879600, 1419883200, 
    1419886800, 1419890400, 1419894000, 1419897600, 1419901200, 1419904800, 
    1419908400, 1419912000, 1419915600, 1419919200, 1419922800, 1419926400, 
    1419930000, 1419933600, 1419937200, 1419940800, 1419944400, 1419948000, 
    1419951600, 1419955200, 1419958800, 1419962400, 1419966000, 1419969600, 
    1419973200, 1419976800, 1419980400, 1419984000, 1419987600, 1419991200, 
    1419994800, 1419998400, 1420002000, 1420005600, 1420009200, 1420012800, 
    1420016400, 1420020000, 1420023600, 1420027200, 1420030800, 1420034400, 
    1420038000, 1420041600, 1420045200, 1420048800, 1420052400, 1420056000, 
    1420059600, 1420063200, 1420066800, 1420070400, 1420074000, 1420077600, 
    1420081200, 1420084800, 1420088400, 1420092000, 1420095600, 1420099200, 
    1420102800, 1420106400, 1420110000, 1420113600, 1420117200, 1420120800, 
    1420124400, 1420128000, 1420131600, 1420135200, 1420138800, 1420142400, 
    1420146000, 1420149600, 1420153200, 1420156800, 1420160400, 1420164000, 
    1420167600, 1420171200, 1420174800, 1420178400, 1420182000, 1420185600, 
    1420189200, 1420192800, 1420196400, 1420200000, 1420203600, 1420207200, 
    1420210800, 1420214400, 1420218000, 1420221600, 1420225200, 1420228800, 
    1420232400, 1420236000, 1420239600, 1420243200, 1420246800, 1420250400, 
    1420254000, 1420257600, 1420261200, 1420264800, 1420268400, 1420272000, 
    1420275600, 1420279200, 1420282800, 1420286400, 1420290000, 1420293600, 
    1420297200, 1420300800, 1420304400, 1420308000, 1420311600, 1420315200, 
    1420318800, 1420322400, 1420326000, 1420329600, 1420333200, 1420336800, 
    1420340400, 1420344000, 1420347600, 1420351200, 1420354800, 1420358400, 
    1420362000, 1420365600, 1420369200, 1420372800, 1420376400, 1420380000, 
    1420383600, 1420387200, 1420390800, 1420394400, 1420398000, 1420401600, 
    1420405200, 1420408800, 1420412400, 1420416000, 1420419600, 1420423200, 
    1420426800, 1420430400, 1420434000, 1420437600, 1420441200, 1420444800, 
    1420448400, 1420452000, 1420455600, 1420459200, 1420462800, 1420466400, 
    1420470000, 1420473600, 1420477200, 1420480800, 1420484400, 1420488000, 
    1420491600, 1420495200, 1420498800, 1420502400, 1420506000, 1420509600, 
    1420513200, 1420516800, 1420520400, 1420524000, 1420527600, 1420531200, 
    1420534800, 1420538400, 1420542000, 1420545600, 1420549200, 1420552800, 
    1420556400, 1420560000, 1420563600, 1420567200, 1420570800, 1420574400, 
    1420578000, 1420581600, 1420585200, 1420588800, 1420592400, 1420596000, 
    1420599600, 1420603200, 1420606800, 1420610400, 1420614000, 1420617600, 
    1420621200, 1420624800, 1420628400, 1420632000, 1420635600, 1420639200, 
    1420642800, 1420646400, 1420650000, 1420653600, 1420657200, 1420660800, 
    1420664400, 1420668000, 1420671600, 1420675200, 1420678800, 1420682400, 
    1420686000, 1420689600, 1420693200, 1420696800, 1420700400, 1420704000, 
    1420707600, 1420711200, 1420714800, 1420718400, 1420722000, 1420725600, 
    1420729200, 1420732800, 1420736400, 1420740000, 1420743600, 1420747200, 
    1420750800, 1420754400, 1420758000, 1420761600, 1420765200, 1420768800, 
    1420772400, 1420776000, 1420779600, 1420783200, 1420786800, 1420790400, 
    1420794000, 1420797600, 1420801200, 1420804800, 1420808400, 1420812000, 
    1420815600, 1420819200, 1420822800, 1420826400, 1420830000, 1420833600, 
    1420837200, 1420840800, 1420844400, 1420848000, 1420851600, 1420855200, 
    1420858800, 1420862400, 1420866000, 1420869600, 1420873200, 1420876800, 
    1420880400, 1420884000, 1420887600, 1420891200, 1420894800, 1420898400, 
    1420902000, 1420905600, 1420909200, 1420912800, 1420916400, 1420920000, 
    1420923600, 1420927200, 1420930800, 1420934400, 1420938000, 1420941600, 
    1420945200, 1420948800, 1420952400, 1420956000, 1420959600, 1420963200, 
    1420966800, 1420970400, 1420974000, 1420977600, 1420981200, 1420984800, 
    1420988400, 1420992000, 1420995600, 1420999200, 1421002800, 1421006400, 
    1421010000, 1421013600, 1421017200, 1421020800, 1421024400, 1421028000, 
    1421031600, 1421035200, 1421038800, 1421042400, 1421046000, 1421049600, 
    1421053200, 1421056800, 1421060400, 1421064000, 1421067600, 1421071200, 
    1421074800, 1421078400, 1421082000, 1421085600, 1421089200, 1421092800, 
    1421096400, 1421100000, 1421103600, 1421107200, 1421110800, 1421114400, 
    1421118000, 1421121600, 1421125200, 1421128800, 1421132400, 1421136000, 
    1421139600, 1421143200, 1421146800, 1421150400, 1421154000, 1421157600, 
    1421161200, 1421164800, 1421168400, 1421172000, 1421175600, 1421179200, 
    1421182800, 1421186400, 1421190000, 1421193600, 1421197200, 1421200800, 
    1421204400, 1421208000, 1421211600, 1421215200, 1421218800, 1421222400, 
    1421226000, 1421229600, 1421233200, 1421236800, 1421240400, 1421244000, 
    1421247600, 1421251200, 1421254800, 1421258400, 1421262000, 1421265600, 
    1421269200, 1421272800, 1421276400, 1421280000, 1421283600, 1421287200, 
    1421290800, 1421294400, 1421298000, 1421301600, 1421305200, 1421308800, 
    1421312400, 1421316000, 1421319600, 1421323200, 1421326800, 1421330400, 
    1421334000, 1421337600, 1421341200, 1421344800, 1421348400, 1421352000, 
    1421355600, 1421359200, 1421362800, 1421366400, 1421370000, 1421373600, 
    1421377200, 1421380800, 1421384400, 1421388000, 1421391600, 1421395200, 
    1421398800, 1421402400, 1421406000, 1421409600, 1421413200, 1421416800, 
    1421420400, 1421424000, 1421427600, 1421431200, 1421434800, 1421438400, 
    1421442000, 1421445600, 1421449200, 1421452800, 1421456400, 1421460000, 
    1421463600, 1421467200, 1421470800, 1421474400, 1421478000, 1421481600, 
    1421485200, 1421488800, 1421492400, 1421496000, 1421499600, 1421503200, 
    1421506800, 1421510400, 1421514000, 1421517600, 1421521200, 1421524800, 
    1421528400, 1421532000, 1421535600, 1421539200, 1421542800, 1421546400, 
    1421550000, 1421553600, 1421557200, 1421560800, 1421564400, 1421568000, 
    1421571600, 1421575200, 1421578800, 1421582400, 1421586000, 1421589600, 
    1421593200, 1421596800, 1421600400, 1421604000, 1421607600, 1421611200, 
    1421614800, 1421618400, 1421622000, 1421625600, 1421629200, 1421632800, 
    1421636400, 1421640000, 1421643600, 1421647200, 1421650800, 1421654400, 
    1421658000, 1421661600, 1421665200, 1421668800, 1421672400, 1421676000, 
    1421679600, 1421683200, 1421686800, 1421690400, 1421694000, 1421697600, 
    1421701200, 1421704800, 1421708400, 1421712000, 1421715600, 1421719200, 
    1421722800, 1421726400, 1421730000, 1421733600, 1421737200, 1421740800, 
    1421744400, 1421748000, 1421751600, 1421755200, 1421758800, 1421762400, 
    1421766000, 1421769600, 1421773200, 1421776800, 1421780400, 1421784000, 
    1421787600, 1421791200, 1421794800, 1421798400, 1421802000, 1421805600, 
    1421809200, 1421812800, 1421816400, 1421820000, 1421823600, 1421827200, 
    1421830800, 1421834400, 1421838000, 1421841600, 1421845200, 1421848800, 
    1421852400, 1421856000, 1421859600, 1421863200, 1421866800, 1421870400, 
    1421874000, 1421877600, 1421881200, 1421884800, 1421888400, 1421892000, 
    1421895600, 1421899200, 1421902800, 1421906400, 1421910000, 1421913600, 
    1421917200, 1421920800, 1421924400, 1421928000, 1421931600, 1421935200, 
    1421938800, 1421942400, 1421946000, 1421949600, 1421953200, 1421956800, 
    1421960400, 1421964000, 1421967600, 1421971200, 1421974800, 1421978400, 
    1421982000, 1421985600, 1421989200, 1421992800, 1421996400, 1422000000, 
    1422003600, 1422007200, 1422010800, 1422014400, 1422018000, 1422021600, 
    1422025200, 1422028800, 1422032400, 1422036000, 1422039600, 1422043200, 
    1422046800, 1422050400, 1422054000, 1422057600, 1422061200, 1422064800, 
    1422068400, 1422072000, 1422075600, 1422079200, 1422082800, 1422086400, 
    1422090000, 1422093600, 1422097200, 1422100800, 1422104400, 1422108000, 
    1422111600, 1422115200, 1422118800, 1422122400, 1422126000, 1422129600, 
    1422133200, 1422136800, 1422140400, 1422144000, 1422147600, 1422151200, 
    1422154800, 1422158400, 1422162000, 1422165600, 1422169200, 1422172800, 
    1422176400, 1422180000, 1422183600, 1422187200, 1422190800, 1422194400, 
    1422198000, 1422201600, 1422205200, 1422208800, 1422212400, 1422216000, 
    1422219600, 1422223200, 1422226800, 1422230400, 1422234000, 1422237600, 
    1422241200, 1422244800, 1422248400, 1422252000, 1422255600, 1422259200, 
    1422262800, 1422266400, 1422270000, 1422273600, 1422277200, 1422280800, 
    1422284400, 1422288000, 1422291600, 1422295200, 1422298800, 1422302400, 
    1422306000, 1422309600, 1422313200, 1422316800, 1422320400, 1422324000, 
    1422327600, 1422331200, 1422334800, 1422338400, 1422342000, 1422345600, 
    1422349200, 1422352800, 1422356400, 1422360000, 1422363600, 1422367200, 
    1422370800, 1422374400, 1422378000, 1422381600, 1422385200, 1422388800, 
    1422392400, 1422396000, 1422399600, 1422403200, 1422406800, 1422410400, 
    1422414000, 1422417600, 1422421200, 1422424800, 1422428400, 1422432000, 
    1422435600, 1422439200, 1422442800, 1422446400, 1422450000, 1422453600, 
    1422457200, 1422460800, 1422464400, 1422468000, 1422471600, 1422475200, 
    1422478800, 1422482400, 1422486000, 1422489600, 1422493200, 1422496800, 
    1422500400, 1422504000, 1422507600, 1422511200, 1422514800, 1422518400, 
    1422522000, 1422525600, 1422529200, 1422532800, 1422536400, 1422540000, 
    1422543600, 1422547200, 1422550800, 1422554400, 1422558000, 1422561600, 
    1422565200, 1422568800, 1422572400, 1422576000, 1422579600, 1422583200, 
    1422586800, 1422590400, 1422594000, 1422597600, 1422601200, 1422604800, 
    1422608400, 1422612000, 1422615600, 1422619200, 1422622800, 1422626400, 
    1422630000, 1422633600, 1422637200, 1422640800, 1422644400, 1422648000, 
    1422651600, 1422655200, 1422658800, 1422662400, 1422666000, 1422669600, 
    1422673200, 1422676800, 1422680400, 1422684000, 1422687600, 1422691200, 
    1422694800, 1422698400, 1422702000, 1422705600, 1422709200, 1422712800, 
    1422716400, 1422720000, 1422723600, 1422727200, 1422730800, 1422734400, 
    1422738000, 1422741600, 1422745200, 1422748800, 1422752400, 1422756000, 
    1422759600, 1422763200, 1422766800, 1422770400, 1422774000, 1422777600, 
    1422781200, 1422784800, 1422788400, 1422792000, 1422795600, 1422799200, 
    1422802800, 1422806400, 1422810000, 1422813600, 1422817200, 1422820800, 
    1422824400, 1422828000, 1422831600, 1422835200, 1422838800, 1422842400, 
    1422846000, 1422849600, 1422853200, 1422856800, 1422860400, 1422864000, 
    1422867600, 1422871200, 1422874800, 1422878400, 1422882000, 1422885600, 
    1422889200, 1422892800, 1422896400, 1422900000, 1422903600, 1422907200, 
    1422910800, 1422914400, 1422918000, 1422921600, 1422925200, 1422928800, 
    1422932400, 1422936000, 1422939600, 1422943200, 1422946800, 1422950400, 
    1422954000, 1422957600, 1422961200, 1422964800, 1422968400, 1422972000, 
    1422975600, 1422979200, 1422982800, 1422986400, 1422990000, 1422993600, 
    1422997200, 1423000800, 1423004400, 1423008000, 1423011600, 1423015200, 
    1423018800, 1423022400, 1423026000, 1423029600, 1423033200, 1423036800, 
    1423040400, 1423044000, 1423047600, 1423051200, 1423054800, 1423058400, 
    1423062000, 1423065600, 1423069200, 1423072800, 1423076400, 1423080000, 
    1423083600, 1423087200, 1423090800, 1423094400, 1423098000, 1423101600, 
    1423105200, 1423108800, 1423112400, 1423116000, 1423119600, 1423123200, 
    1423126800, 1423130400, 1423134000, 1423137600, 1423141200, 1423144800, 
    1423148400, 1423152000, 1423155600, 1423159200, 1423162800, 1423166400, 
    1423170000, 1423173600, 1423177200, 1423180800, 1423184400, 1423188000, 
    1423191600, 1423195200, 1423198800, 1423202400, 1423206000, 1423209600, 
    1423213200, 1423216800, 1423220400, 1423224000, 1423227600, 1423231200, 
    1423234800, 1423238400, 1423242000, 1423245600, 1423249200, 1423252800, 
    1423256400, 1423260000, 1423263600, 1423267200, 1423270800, 1423274400, 
    1423278000, 1423281600, 1423285200, 1423288800, 1423292400, 1423296000, 
    1423299600, 1423303200, 1423306800, 1423310400, 1423314000, 1423317600, 
    1423321200, 1423324800, 1423328400, 1423332000, 1423335600, 1423339200, 
    1423342800, 1423346400, 1423350000, 1423353600, 1423357200, 1423360800, 
    1423364400, 1423368000, 1423371600, 1423375200, 1423378800, 1423382400, 
    1423386000, 1423389600, 1423393200, 1423396800, 1423400400, 1423404000, 
    1423407600, 1423411200, 1423414800, 1423418400, 1423422000, 1423425600, 
    1423429200, 1423432800, 1423436400, 1423440000, 1423443600, 1423447200, 
    1423450800, 1423454400, 1423458000, 1423461600, 1423465200, 1423468800, 
    1423472400, 1423476000, 1423479600, 1423483200, 1423486800, 1423490400, 
    1423494000, 1423497600, 1423501200, 1423504800, 1423508400, 1423512000, 
    1423515600, 1423519200, 1423522800, 1423526400, 1423530000, 1423533600, 
    1423537200, 1423540800, 1423544400, 1423548000, 1423551600, 1423555200, 
    1423558800, 1423562400, 1423566000, 1423569600, 1423573200, 1423576800, 
    1423580400, 1423584000, 1423587600, 1423591200, 1423594800, 1423598400, 
    1423602000, 1423605600, 1423609200, 1423612800, 1423616400, 1423620000, 
    1423623600, 1423627200, 1423630800, 1423634400, 1423638000, 1423641600, 
    1423645200, 1423648800, 1423652400, 1423656000, 1423659600, 1423663200, 
    1423666800, 1423670400, 1423674000, 1423677600, 1423681200, 1423684800, 
    1423688400, 1423692000, 1423695600, 1423699200, 1423702800, 1423706400, 
    1423710000, 1423713600, 1423717200, 1423720800, 1423724400, 1423728000, 
    1423731600, 1423735200, 1423738800, 1423742400, 1423746000, 1423749600, 
    1423753200, 1423756800, 1423760400, 1423764000, 1423767600, 1423771200, 
    1423774800, 1423778400, 1423782000, 1423785600, 1423789200, 1423792800, 
    1423796400, 1423800000, 1423803600, 1423807200, 1423810800, 1423814400, 
    1423818000, 1423821600, 1423825200, 1423828800, 1423832400, 1423836000, 
    1423839600, 1423843200, 1423846800, 1423850400, 1423854000, 1423857600, 
    1423861200, 1423864800, 1423868400, 1423872000, 1423875600, 1423879200, 
    1423882800, 1423886400, 1423890000, 1423893600, 1423897200, 1423900800, 
    1423904400, 1423908000, 1423911600, 1423915200, 1423918800, 1423922400, 
    1423926000, 1423929600, 1423933200, 1423936800, 1423940400, 1423944000, 
    1423947600, 1423951200, 1423954800, 1423958400, 1423962000, 1423965600, 
    1423969200, 1423972800, 1423976400, 1423980000, 1423983600, 1423987200, 
    1423990800, 1423994400, 1423998000, 1424001600, 1424005200, 1424008800, 
    1424012400, 1424016000, 1424019600, 1424023200, 1424026800, 1424030400, 
    1424034000, 1424037600, 1424041200, 1424044800, 1424048400, 1424052000, 
    1424055600, 1424059200, 1424062800, 1424066400, 1424070000, 1424073600, 
    1424077200, 1424080800, 1424084400, 1424088000, 1424091600, 1424095200, 
    1424098800, 1424102400, 1424106000, 1424109600, 1424113200, 1424116800, 
    1424120400, 1424124000, 1424127600, 1424131200, 1424134800, 1424138400, 
    1424142000, 1424145600, 1424149200, 1424152800, 1424156400, 1424160000, 
    1424163600, 1424167200, 1424170800, 1424174400, 1424178000, 1424181600, 
    1424185200, 1424188800, 1424192400, 1424196000, 1424199600, 1424203200, 
    1424206800, 1424210400, 1424214000, 1424217600, 1424221200, 1424224800, 
    1424228400, 1424232000, 1424235600, 1424239200, 1424242800, 1424246400, 
    1424250000, 1424253600, 1424257200, 1424260800, 1424264400, 1424268000, 
    1424271600, 1424275200, 1424278800, 1424282400, 1424286000, 1424289600, 
    1424293200, 1424296800, 1424300400, 1424304000, 1424307600, 1424311200, 
    1424314800, 1424318400, 1424322000, 1424325600, 1424329200, 1424332800, 
    1424336400, 1424340000, 1424343600, 1424347200, 1424350800, 1424354400, 
    1424358000, 1424361600, 1424365200, 1424368800, 1424372400, 1424376000, 
    1424379600, 1424383200, 1424386800, 1424390400, 1424394000, 1424397600, 
    1424401200, 1424404800, 1424408400, 1424412000, 1424415600, 1424419200, 
    1424422800, 1424426400, 1424430000, 1424433600, 1424437200, 1424440800, 
    1424444400, 1424448000, 1424451600, 1424455200, 1424458800, 1424462400, 
    1424466000, 1424469600, 1424473200, 1424476800, 1424480400, 1424484000, 
    1424487600, 1424491200, 1424494800, 1424498400, 1424502000, 1424505600, 
    1424509200, 1424512800, 1424516400, 1424520000, 1424523600, 1424527200, 
    1424530800, 1424534400, 1424538000, 1424541600, 1424545200, 1424548800, 
    1424552400, 1424556000, 1424559600, 1424563200, 1424566800, 1424570400, 
    1424574000, 1424577600, 1424581200, 1424584800, 1424588400, 1424592000, 
    1424595600, 1424599200, 1424602800, 1424606400, 1424610000, 1424613600, 
    1424617200, 1424620800, 1424624400, 1424628000, 1424631600, 1424635200, 
    1424638800, 1424642400, 1424646000, 1424649600, 1424653200, 1424656800, 
    1424660400, 1424664000, 1424667600, 1424671200, 1424674800, 1424678400, 
    1424682000, 1424685600, 1424689200, 1424692800, 1424696400, 1424700000, 
    1424703600, 1424707200, 1424710800, 1424714400, 1424718000, 1424721600, 
    1424725200, 1424728800, 1424732400, 1424736000, 1424739600, 1424743200, 
    1424746800, 1424750400, 1424754000, 1424757600, 1424761200, 1424764800, 
    1424768400, 1424772000, 1424775600, 1424779200, 1424782800, 1424786400, 
    1424790000, 1424793600, 1424797200, 1424800800, 1424804400, 1424808000, 
    1424811600, 1424815200, 1424818800, 1424822400, 1424826000, 1424829600, 
    1424833200, 1424836800, 1424840400, 1424844000, 1424847600, 1424851200, 
    1424854800, 1424858400, 1424862000, 1424865600, 1424869200, 1424872800, 
    1424876400, 1424880000, 1424883600, 1424887200, 1424890800, 1424894400, 
    1424898000, 1424901600, 1424905200, 1424908800, 1424912400, 1424916000, 
    1424919600, 1424923200, 1424926800, 1424930400, 1424934000, 1424937600, 
    1424941200, 1424944800, 1424948400, 1424952000, 1424955600, 1424959200, 
    1424962800, 1424966400, 1424970000, 1424973600, 1424977200, 1424980800, 
    1424984400, 1424988000, 1424991600, 1424995200, 1424998800, 1425002400, 
    1425006000, 1425009600, 1425013200, 1425016800, 1425020400, 1425024000, 
    1425027600, 1425031200, 1425034800, 1425038400, 1425042000, 1425045600, 
    1425049200, 1425052800, 1425056400, 1425060000, 1425063600, 1425067200, 
    1425070800, 1425074400, 1425078000, 1425081600, 1425085200, 1425088800, 
    1425092400, 1425096000, 1425099600, 1425103200, 1425106800, 1425110400, 
    1425114000, 1425117600, 1425121200, 1425124800, 1425128400, 1425132000, 
    1425135600, 1425139200, 1425142800, 1425146400, 1425150000, 1425153600, 
    1425157200, 1425160800, 1425164400, 1425168000, 1425171600, 1425175200, 
    1425178800, 1425182400, 1425186000, 1425189600, 1425193200, 1425196800, 
    1425200400, 1425204000, 1425207600, 1425211200, 1425214800, 1425218400, 
    1425222000, 1425225600, 1425229200, 1425232800, 1425236400, 1425240000, 
    1425243600, 1425247200, 1425250800, 1425254400, 1425258000, 1425261600, 
    1425265200, 1425268800, 1425272400, 1425276000, 1425279600, 1425283200, 
    1425286800, 1425290400, 1425294000, 1425297600, 1425301200, 1425304800, 
    1425308400, 1425312000, 1425315600, 1425319200, 1425322800, 1425326400, 
    1425330000, 1425333600, 1425337200, 1425340800, 1425344400, 1425348000, 
    1425351600, 1425355200, 1425358800, 1425362400, 1425366000, 1425369600, 
    1425373200, 1425376800, 1425380400, 1425384000, 1425387600, 1425391200, 
    1425394800, 1425398400, 1425402000, 1425405600, 1425409200, 1425412800, 
    1425416400, 1425420000, 1425423600, 1425427200, 1425430800, 1425434400, 
    1425438000, 1425441600, 1425445200, 1425448800, 1425452400, 1425456000, 
    1425459600, 1425463200, 1425466800, 1425470400, 1425474000, 1425477600, 
    1425481200, 1425484800, 1425488400, 1425492000, 1425495600, 1425499200, 
    1425502800, 1425506400, 1425510000, 1425513600, 1425517200, 1425520800, 
    1425524400, 1425528000, 1425531600, 1425535200, 1425538800, 1425542400, 
    1425546000, 1425549600, 1425553200, 1425556800, 1425560400, 1425564000, 
    1425567600, 1425571200, 1425574800, 1425578400, 1425582000, 1425585600, 
    1425589200, 1425592800, 1425596400, 1425600000, 1425603600, 1425607200, 
    1425610800, 1425614400, 1425618000, 1425621600, 1425625200, 1425628800, 
    1425632400, 1425636000, 1425639600, 1425643200, 1425646800, 1425650400, 
    1425654000, 1425657600, 1425661200, 1425664800, 1425668400, 1425672000, 
    1425675600, 1425679200, 1425682800, 1425686400, 1425690000, 1425693600, 
    1425697200, 1425700800, 1425704400, 1425708000, 1425711600, 1425715200, 
    1425718800, 1425722400, 1425726000, 1425729600, 1425733200, 1425736800, 
    1425740400, 1425744000, 1425747600, 1425751200, 1425754800, 1425758400, 
    1425762000, 1425765600, 1425769200, 1425772800, 1425776400, 1425780000, 
    1425783600, 1425787200, 1425790800, 1425794400, 1425798000, 1425801600, 
    1425805200, 1425808800, 1425812400, 1425816000, 1425819600, 1425823200, 
    1425826800, 1425830400, 1425834000, 1425837600, 1425841200, 1425844800, 
    1425848400, 1425852000, 1425855600, 1425859200, 1425862800, 1425866400, 
    1425870000, 1425873600, 1425877200, 1425880800, 1425884400, 1425888000, 
    1425891600, 1425895200, 1425898800, 1425902400, 1425906000, 1425909600, 
    1425913200, 1425916800, 1425920400, 1425924000, 1425927600, 1425931200, 
    1425934800, 1425938400, 1425942000, 1425945600, 1425949200, 1425952800, 
    1425956400, 1425960000, 1425963600, 1425967200, 1425970800, 1425974400, 
    1425981600, 1425985200, 1425988800, 1425992400, 1425996000, 1425999600, 
    1426003200, 1426006800, 1426010400, 1426014000, 1426017600, 1426021200, 
    1426024800, 1426028400, 1426032000, 1426035600, 1426039200, 1426042800, 
    1426046400, 1426050000, 1426053600, 1426057200, 1426060800, 1426064400, 
    1426068000, 1426071600, 1426075200, 1426078800, 1426082400, 1426086000, 
    1426089600, 1426093200, 1426096800, 1426100400, 1426104000, 1426107600, 
    1426111200, 1426114800, 1426118400, 1426122000, 1426125600, 1426129200, 
    1426132800, 1426136400, 1426140000, 1426143600, 1426147200, 1426150800, 
    1426154400, 1426158000, 1426161600, 1426165200, 1426168800, 1426172400, 
    1426176000, 1426179600, 1426183200, 1426186800, 1426190400, 1426194000, 
    1426197600, 1426201200, 1426204800, 1426208400, 1426212000, 1426215600, 
    1426219200, 1426222800, 1426226400, 1426230000, 1426233600, 1426237200, 
    1426240800, 1426244400, 1426248000, 1426251600, 1426255200, 1426258800, 
    1426262400, 1426266000, 1426269600, 1426273200, 1426276800, 1426280400, 
    1426284000, 1426287600, 1426291200, 1426294800, 1426298400, 1426302000, 
    1426305600, 1426309200, 1426312800, 1426316400, 1426320000, 1426323600, 
    1426327200, 1426330800, 1426334400, 1426338000, 1426341600, 1426345200, 
    1426348800, 1426352400, 1426356000, 1426359600, 1426363200, 1426366800, 
    1426370400, 1426374000, 1426377600, 1426381200, 1426384800, 1426388400, 
    1426392000, 1426395600, 1426399200, 1426402800, 1426406400, 1426410000, 
    1426413600, 1426417200, 1426420800, 1426424400, 1426428000, 1426431600, 
    1426435200, 1426438800, 1426442400, 1426446000, 1426449600, 1426453200, 
    1426456800, 1426460400, 1426464000, 1426467600, 1426471200, 1426474800, 
    1426478400, 1426482000, 1426485600, 1426489200, 1426492800, 1426496400, 
    1426500000, 1426503600, 1426507200, 1426510800, 1426514400, 1426518000, 
    1426521600, 1426525200, 1426528800, 1426532400, 1426536000, 1426539600, 
    1426543200, 1426546800, 1426550400, 1426554000, 1426557600, 1426561200, 
    1426564800, 1426568400, 1426572000, 1426575600, 1426579200, 1426582800, 
    1426586400, 1426590000, 1426593600, 1426597200, 1426600800, 1426604400, 
    1426608000, 1426611600, 1426615200, 1426618800, 1426622400, 1426626000, 
    1426629600, 1426633200, 1426636800, 1426640400, 1426644000, 1426647600, 
    1426651200, 1426654800, 1426658400, 1426662000, 1426665600, 1426669200, 
    1426672800, 1426676400, 1426680000, 1426683600, 1426687200, 1426690800, 
    1426694400, 1426698000, 1426701600, 1426705200, 1426708800, 1426712400, 
    1426716000, 1426719600, 1426723200, 1426726800, 1426730400, 1426734000, 
    1426737600, 1426741200, 1426744800, 1426748400, 1426752000, 1426755600, 
    1426759200, 1426762800, 1426766400, 1426770000, 1426773600, 1426777200, 
    1426780800, 1426784400, 1426788000, 1426791600, 1426795200, 1426798800, 
    1426802400, 1426806000, 1426809600, 1426813200, 1426816800, 1426820400, 
    1426824000, 1426827600, 1426831200, 1426834800, 1426838400, 1426842000, 
    1426845600, 1426849200, 1426852800, 1426856400, 1426860000, 1426863600, 
    1426867200, 1426870800, 1426874400, 1426878000, 1426881600, 1426885200, 
    1426888800, 1426892400, 1426896000, 1426899600, 1426903200, 1426906800, 
    1426910400, 1426914000, 1426917600, 1426921200, 1426924800, 1426928400, 
    1426932000, 1426935600, 1426939200, 1426942800, 1426946400, 1426950000, 
    1426953600, 1426957200, 1426960800, 1426964400, 1426968000, 1426971600, 
    1426975200, 1426978800, 1426982400, 1426986000, 1426989600, 1426993200, 
    1426996800, 1427000400, 1427004000, 1427007600, 1427011200, 1427014800, 
    1427018400, 1427022000, 1427025600, 1427029200, 1427032800, 1427036400, 
    1427040000, 1427043600, 1427047200, 1427050800, 1427054400, 1427058000, 
    1427061600, 1427065200, 1427068800, 1427072400, 1427076000, 1427079600, 
    1427083200, 1427086800, 1427090400, 1427094000, 1427097600, 1427101200, 
    1427104800, 1427108400, 1427112000, 1427115600, 1427119200, 1427122800, 
    1427126400, 1427130000, 1427133600, 1427137200, 1427140800, 1427144400, 
    1427148000, 1427151600, 1427155200, 1427158800, 1427162400, 1427166000, 
    1427169600, 1427173200, 1427176800, 1427180400, 1427184000, 1427187600, 
    1427191200, 1427194800, 1427198400, 1427202000, 1427205600, 1427209200, 
    1427212800, 1427216400, 1427220000, 1427223600, 1427227200, 1427230800, 
    1427234400, 1427238000, 1427252400, 1427256000, 1427263200, 1427266800, 
    1427270400, 1427274000, 1427277600, 1427281200, 1427284800, 1427288400, 
    1427292000, 1427295600, 1427299200, 1427302800, 1427306400, 1427310000, 
    1427313600, 1427317200, 1427320800, 1427324400, 1427328000, 1427331600, 
    1427335200, 1427338800, 1427342400, 1427346000, 1427349600, 1427353200, 
    1427356800, 1427360400, 1427364000, 1427367600, 1427371200, 1427374800, 
    1427378400, 1427382000, 1427385600, 1427389200, 1427392800, 1427396400, 
    1427400000, 1427403600, 1427407200, 1427410800, 1427414400, 1427418000, 
    1427421600, 1427425200, 1427428800, 1427432400, 1427436000, 1427439600, 
    1427443200, 1427446800, 1427450400, 1427454000, 1427457600, 1427461200, 
    1427464800, 1427468400, 1427472000, 1427475600, 1427479200, 1427482800, 
    1427486400, 1427490000, 1427493600, 1427497200, 1427500800, 1427504400, 
    1427508000, 1427511600, 1427515200, 1427518800, 1427522400, 1427526000, 
    1427529600, 1427533200, 1427536800, 1427540400, 1427544000, 1427547600, 
    1427551200, 1427554800, 1427558400, 1427562000, 1427565600, 1427569200, 
    1427572800, 1427576400, 1427580000, 1427583600, 1427587200, 1427590800, 
    1427594400, 1427598000, 1427601600, 1427605200, 1427608800, 1427612400, 
    1427616000, 1427619600, 1427623200, 1427626800, 1427630400, 1427634000, 
    1427637600, 1427641200, 1427644800, 1427648400, 1427652000, 1427655600, 
    1427659200, 1427662800, 1427666400, 1427670000, 1427673600, 1427677200, 
    1427680800, 1427684400, 1427688000, 1427691600, 1427695200, 1427698800, 
    1427702400, 1427706000, 1427709600, 1427713200, 1427716800, 1427720400, 
    1427724000, 1427727600, 1427731200, 1427734800, 1427738400, 1427742000, 
    1427745600, 1427749200, 1427752800, 1427756400, 1427760000, 1427763600, 
    1427767200, 1427770800, 1427774400, 1427778000, 1427781600, 1427785200, 
    1427788800, 1427792400, 1427796000, 1427799600, 1427803200, 1427806800, 
    1427810400, 1427814000, 1427817600, 1427821200, 1427824800, 1427828400, 
    1427832000, 1427835600, 1427839200, 1427842800, 1427846400, 1427850000, 
    1427853600, 1427857200, 1427860800, 1427864400, 1427868000, 1427871600, 
    1427875200, 1427878800, 1427882400, 1427886000, 1427889600, 1427893200, 
    1427896800, 1427900400, 1427904000, 1427907600, 1427911200, 1427914800, 
    1427918400, 1427922000, 1427925600, 1427929200, 1427932800, 1427936400, 
    1427940000, 1427943600, 1427947200, 1427950800, 1427954400, 1427958000, 
    1427961600, 1427965200, 1427968800, 1427972400, 1427976000, 1427979600, 
    1427983200, 1427986800, 1427990400, 1427994000, 1427997600, 1428001200, 
    1428004800, 1428008400, 1428012000, 1428015600, 1428019200, 1428022800, 
    1428026400, 1428030000, 1428033600, 1428037200, 1428040800, 1428044400, 
    1428048000, 1428051600, 1428055200, 1428058800, 1428062400, 1428066000, 
    1428069600, 1428073200, 1428076800, 1428080400, 1428084000, 1428087600, 
    1428091200, 1428094800, 1428098400, 1428102000, 1428105600, 1428109200, 
    1428112800, 1428116400, 1428120000, 1428123600, 1428127200, 1428130800, 
    1428134400, 1428138000, 1428141600, 1428145200, 1428148800, 1428152400, 
    1428156000, 1428159600, 1428163200, 1428166800, 1428170400, 1428174000, 
    1428177600, 1428181200, 1428184800, 1428188400, 1428192000, 1428195600, 
    1428199200, 1428202800, 1428206400, 1428210000, 1428213600, 1428217200, 
    1428220800, 1428224400, 1428228000, 1428231600, 1428235200, 1428238800, 
    1428242400, 1428246000, 1428249600, 1428253200, 1428256800, 1428260400, 
    1428264000, 1428267600, 1428271200, 1428274800, 1428278400, 1428282000, 
    1428285600, 1428289200, 1428292800, 1428296400, 1428300000, 1428303600, 
    1428307200, 1428310800, 1428314400, 1428318000, 1428321600, 1428325200, 
    1428328800, 1428332400, 1428336000, 1428339600, 1428343200, 1428346800, 
    1428350400, 1428354000, 1428357600, 1428361200, 1428364800, 1428368400, 
    1428372000, 1428375600, 1428379200, 1428382800, 1428386400, 1428390000, 
    1428393600, 1428397200, 1428400800, 1428404400, 1428408000, 1428411600, 
    1428415200, 1428418800, 1428422400, 1428426000, 1428429600, 1428433200, 
    1428436800, 1428440400, 1428444000, 1428447600, 1428451200, 1428454800, 
    1428458400, 1428462000, 1428465600, 1428469200, 1428472800, 1428476400, 
    1428480000, 1428483600, 1428487200, 1428490800, 1428494400, 1428498000, 
    1428501600, 1428505200, 1428508800, 1428512400, 1428516000, 1428519600, 
    1428523200, 1428526800, 1428530400, 1428534000, 1428537600, 1428541200, 
    1428544800, 1428548400, 1428552000, 1428555600, 1428559200, 1428562800, 
    1428566400, 1428570000, 1428573600, 1428577200, 1428580800, 1428584400, 
    1428588000, 1428591600, 1428595200, 1428598800, 1428602400, 1428606000, 
    1428609600, 1428613200, 1428616800, 1428620400, 1428624000, 1428627600, 
    1428631200, 1428634800, 1428638400, 1428642000, 1428645600, 1428649200, 
    1428652800, 1428656400, 1428660000, 1428663600, 1428667200, 1428670800, 
    1428674400, 1428678000, 1428681600, 1428685200, 1428688800, 1428692400, 
    1428696000, 1428699600, 1428703200, 1428706800, 1428717600, 1428721200, 
    1428724800, 1428728400, 1428732000, 1428735600, 1428739200, 1428742800, 
    1428746400, 1428750000, 1428753600, 1428757200, 1428760800, 1428764400, 
    1428768000, 1428771600, 1428775200, 1428778800, 1428782400, 1428786000, 
    1428789600, 1428796800, 1428800400, 1428804000, 1428807600, 1428811200, 
    1428814800, 1428822000, 1428825600, 1428829200, 1428832800, 1428836400, 
    1428840000, 1428843600, 1428847200, 1428850800, 1428854400, 1428858000, 
    1428861600, 1428865200, 1428872400, 1428876000, 1428879600, 1428883200, 
    1428886800, 1428890400, 1428894000, 1428901200, 1428904800, 1428908400, 
    1428912000, 1428915600, 1428922800, 1428926400, 1428930000, 1428933600, 
    1428937200, 1428940800, 1428944400, 1428948000, 1428951600, 1428955200, 
    1428958800, 1428962400, 1428966000, 1428987600, 1428991200, 1428994800, 
    1428998400, 1429002000, 1429005600, 1429009200, 1429012800, 1429016400, 
    1429020000, 1429023600, 1429027200, 1429030800, 1429034400, 1429038000, 
    1429041600, 1429045200, 1429048800, 1429056000, 1429059600, 1429063200, 
    1429066800, 1429070400, 1429074000, 1429081200, 1429084800, 1429088400, 
    1429092000, 1429095600, 1429099200, 1429102800, 1429185600, 1429189200, 
    1429192800, 1429196400, 1429200000, 1429203600, 1429207200, 1429210800, 
    1429214400, 1429218000, 1429221600, 1429225200, 1429236000, 1429239600, 
    1429243200, 1429246800, 1429250400, 1429254000, 1429257600, 1429261200, 
    1429264800, 1429268400, 1429272000, 1429275600, 1429279200, 1429282800, 
    1429286400, 1429290000, 1429293600, 1429297200, 1429300800, 1429304400, 
    1429308000, 1429315200, 1429318800, 1429322400, 1429326000, 1429329600, 
    1429333200, 1429336800, 1429340400, 1429344000, 1429347600, 1429351200, 
    1429354800, 1429358400, 1429362000, 1429365600, 1429369200, 1429372800, 
    1429376400, 1429380000, 1429383600, 1429387200, 1429390800, 1429394400, 
    1429398000, 1429401600, 1429405200, 1429408800, 1429412400, 1429416000, 
    1429419600, 1429423200, 1429426800, 1429430400, 1429434000, 1429437600, 
    1429441200, 1429444800, 1429448400, 1429452000, 1429455600, 1429459200, 
    1429462800, 1429466400, 1429470000, 1429473600, 1429477200, 1429480800, 
    1429484400, 1429488000, 1429491600, 1429495200, 1429498800, 1429502400, 
    1429506000, 1429509600, 1429513200, 1429516800, 1429520400, 1429524000, 
    1429527600, 1429531200, 1429534800, 1429538400, 1429542000, 1429545600, 
    1429549200, 1429552800, 1429556400, 1429560000, 1429563600, 1429567200, 
    1429574400, 1429581600, 1429585200, 1429588800, 1429592400, 1429596000, 
    1429599600, 1429603200, 1429606800, 1429610400, 1429614000, 1429617600, 
    1429621200, 1429628400, 1429635600, 1429639200, 1429646400, 1429650000, 
    1429653600, 1429657200, 1429664400, 1429668000, 1429671600, 1429682400, 
    1429689600, 1429696800, 1429700400, 1429707600, 1429711200, 1429714800, 
    1429718400, 1429722000, 1429725600, 1429729200, 1429736400, 1429740000, 
    1429747200, 1429754400, 1429761600, 1429765200, 1429772400, 1429776000, 
    1429779600, 1429786800, 1429794000, 1429797600, 1429801200, 1429804800, 
    1429812000, 1429815600, 1429819200, 1429822800, 1429826400, 1429833600, 
    1429837200, 1429840800, 1429844400, 1429848000, 1429851600, 1429855200, 
    1429858800, 1429862400, 1429866000, 1429876800, 1429880400, 1429887600, 
    1429891200, 1429898400, 1429912800, 1429916400, 1429923600, 1429927200, 
    1429945200, 1429948800, 1429956000, 1429959600, 1429966800, 1429970400, 
    1429974000, 1429977600, 1429984800, 1429988400, 1429992000, 1429995600, 
    1429999200, 1430002800, 1430006400, 1430017200, 1430020800, 1430028000, 
    1430031600, 1430042400, 1430046000, 1430049600, 1430053200, 1430056800, 
    1430064000, 1430067600, 1430071200, 1430074800, 1430078400, 1430082000, 
    1430085600, 1430096400, 1430103600, 1430110800, 1430121600, 1430132400, 
    1430136000, 1430143200, 1430146800, 1430150400, 1430154000, 1430157600, 
    1430168400, 1430172000, 1430175600, 1430179200, 1430182800, 1430186400, 
    1430190000, 1430197200, 1430204400, 1430208000, 1430211600, 1430218800, 
    1430226000, 1430233200, 1430236800, 1430240400, 1430244000, 1430247600, 
    1430251200, 1430262000, 1430265600, 1430272800, 1430280000, 1430283600, 
    1430287200, 1430290800, 1430294400, 1430298000, 1430301600, 1430305200, 
    1430316000, 1430323200, 1430326800, 1430330400, 1430334000, 1430337600, 
    1430344800, 1430362800, 1430366400, 1430370000, 1430373600, 1430377200, 
    1430380800, 1430388000, 1430402400, 1430406000, 1430409600, 1430413200, 
    1430420400, 1430434800, 1430438400, 1430442000, 1430445600, 1430449200, 
    1430456400, 1430460000, 1430463600, 1430467200, 1430474400, 1430478000, 
    1430481600, 1430488800, 1430492400, 1430496000, 1430499600, 1430503200, 
    1430506800, 1430510400, 1430514000, 1430546400, 1430550000, 1430553600, 
    1430557200, 1430560800, 1430564400, 1430568000, 1430571600, 1430575200, 
    1430578800, 1430582400, 1430586000, 1430589600, 1430593200, 1430596800, 
    1430604000, 1430614800, 1430618400, 1430622000, 1430625600, 1430629200, 
    1430632800, 1430636400, 1430640000, 1430643600, 1430647200, 1430650800, 
    1430654400, 1430658000, 1430661600, 1430665200, 1430668800, 1430672400, 
    1430683200, 1430722800, 1430726400, 1430730000, 1430733600, 1430737200, 
    1430740800, 1430744400, 1430748000, 1430755200, 1430758800, 1430762400, 
    1430766000, 1430769600, 1430773200, 1430776800, 1430780400, 1430784000, 
    1430787600, 1430791200, 1430794800, 1430798400, 1430802000, 1430805600, 
    1430809200, 1430812800, 1430816400, 1430820000, 1430823600, 1430827200, 
    1430830800, 1430834400, 1430838000, 1430841600, 1430845200, 1430848800, 
    1430852400, 1430856000, 1430863200, 1430874000, 1430877600, 1430881200, 
    1430884800, 1430892000, 1430895600, 1430899200, 1430902800, 1430906400, 
    1430910000, 1430913600, 1430917200, 1430920800, 1430924400, 1430928000, 
    1430931600, 1430935200, 1430938800, 1430942400, 1430946000, 1430949600, 
    1430953200, 1430956800, 1430960400, 1430964000, 1430967600, 1430971200, 
    1430974800, 1430978400, 1430982000, 1430985600, 1430989200, 1430992800, 
    1430996400, 1431000000, 1431003600, 1431007200, 1431010800, 1431014400, 
    1431018000, 1431021600, 1431025200, 1431028800, 1431032400, 1431036000, 
    1431039600, 1431043200, 1431050400, 1431054000, 1431057600, 1431061200, 
    1431064800, 1431068400, 1431072000, 1431075600, 1431079200, 1431082800, 
    1431086400, 1431090000, 1431093600, 1431097200, 1431100800, 1431104400, 
    1431108000, 1431111600, 1431115200, 1431122400, 1431133200, 1431136800, 
    1431140400, 1431144000, 1431147600, 1431151200, 1431154800, 1431158400, 
    1431162000, 1431165600, 1431169200, 1431172800, 1431176400, 1431180000, 
    1431183600, 1431187200, 1431194400, 1431198000, 1431201600, 1431205200, 
    1431208800, 1431212400, 1431216000, 1431219600, 1431223200, 1431226800, 
    1431230400, 1431234000, 1431237600, 1431241200, 1431244800, 1431248400, 
    1431252000, 1431255600, 1431259200, 1431262800, 1431266400, 1431270000, 
    1431273600, 1431277200, 1431280800, 1431284400, 1431288000, 1431291600, 
    1431295200, 1431298800, 1431302400, 1431313200, 1431316800, 1431320400, 
    1431324000, 1431327600, 1431331200, 1431334800, 1431338400, 1431342000, 
    1431345600, 1431349200, 1431352800, 1431356400, 1431360000, 1431363600, 
    1431367200, 1431370800, 1431374400, 1431378000, 1431381600, 1431392400, 
    1431396000, 1431399600, 1431403200, 1431406800, 1431410400, 1431414000, 
    1431417600, 1431421200, 1431424800, 1431428400, 1431432000, 1431435600, 
    1431439200, 1431442800, 1431446400, 1431450000, 1431453600, 1431457200, 
    1431460800, 1431464400, 1431468000, 1431471600, 1431475200, 1431478800, 
    1431482400, 1431486000, 1431489600, 1431493200, 1431496800, 1431500400, 
    1431504000, 1431507600, 1431511200, 1431514800, 1431518400, 1431522000, 
    1431525600, 1431529200, 1431532800, 1431536400, 1431550800, 1431554400, 
    1431558000, 1431561600, 1431565200, 1431568800, 1431572400, 1431576000, 
    1431579600, 1431583200, 1431586800, 1431590400, 1431594000, 1431597600, 
    1431601200, 1431604800, 1431608400, 1431612000, 1431615600, 1431619200, 
    1431622800, 1431626400, 1431630000, 1431633600, 1431637200, 1431640800, 
    1431651600, 1431655200, 1431658800, 1431662400, 1431666000, 1431669600, 
    1431673200, 1431676800, 1431680400, 1431684000, 1431687600, 1431691200, 
    1431694800, 1431698400, 1431702000, 1431705600, 1431709200, 1431712800, 
    1431716400, 1431723600, 1431727200, 1431730800, 1431734400, 1431738000, 
    1431741600, 1431745200, 1431748800, 1431752400, 1431756000, 1431759600, 
    1431763200, 1431766800, 1431770400, 1431774000, 1431777600, 1431781200, 
    1431784800, 1431788400, 1431792000, 1431795600, 1431810000, 1431813600, 
    1431817200, 1431820800, 1431824400, 1431828000, 1431831600, 1431835200, 
    1431838800, 1431842400, 1431846000, 1431849600, 1431853200, 1431856800, 
    1431860400, 1431864000, 1431867600, 1431871200, 1431874800, 1431878400, 
    1431882000, 1431885600, 1431889200, 1431892800, 1431896400, 1431900000, 
    1431910800, 1431914400, 1431918000, 1431921600, 1431925200, 1431928800, 
    1431932400, 1431936000, 1431939600, 1431943200, 1431946800, 1431950400, 
    1431954000, 1431957600, 1431961200, 1431964800, 1431968400, 1431972000, 
    1431975600, 1431982800, 1431986400, 1431990000, 1431993600, 1431997200, 
    1432000800, 1432004400, 1432008000, 1432011600, 1432015200, 1432018800, 
    1432022400, 1432026000, 1432029600, 1432033200, 1432036800, 1432040400, 
    1432044000, 1432047600, 1432051200, 1432054800, 1432062000, 1432069200, 
    1432072800, 1432076400, 1432083600, 1432087200, 1432090800, 1432098000, 
    1432101600, 1432105200, 1432108800, 1432112400, 1432116000, 1432119600, 
    1432123200, 1432126800, 1432130400, 1432134000, 1432137600, 1432141200, 
    1432144800, 1432148400, 1432152000, 1432155600, 1432159200, 1432162800, 
    1432170000, 1432173600, 1432177200, 1432180800, 1432184400, 1432188000, 
    1432191600, 1432195200, 1432198800, 1432202400, 1432206000, 1432209600, 
    1432213200, 1432216800, 1432220400, 1432224000, 1432227600, 1432231200, 
    1432234800, 1432242000, 1432249200, 1432252800, 1432256400, 1432260000, 
    1432263600, 1432267200, 1432270800, 1432274400, 1432278000, 1432281600, 
    1432285200, 1432288800, 1432292400, 1432296000, 1432299600, 1432303200, 
    1432306800, 1432310400, 1432314000, 1432321200, 1432328400, 1432332000, 
    1432335600, 1432342800, 1432346400, 1432350000, 1432353600, 1432357200, 
    1432360800, 1432364400, 1432368000, 1432371600, 1432375200, 1432378800, 
    1432382400, 1432386000, 1432389600, 1432393200, 1432396800, 1432411200, 
    1432414800, 1432418400, 1432422000, 1432432800, 1432436400, 1432458000, 
    1432461600, 1432465200, 1432468800, 1432472400, 1432479600, 1432483200, 
    1432490400, 1432501200, 1432508400, 1432512000, 1432515600, 1432519200, 
    1432522800, 1432533600, 1432537200, 1432540800, 1432544400, 1432548000, 
    1432555200, 1432558800, 1432562400, 1432566000, 1432569600, 1432573200, 
    1432580400, 1432587600, 1432591200, 1432594800, 1432598400, 1432602000, 
    1432605600, 1432609200, 1432616400, 1432620000, 1432627200, 1432630800, 
    1432634400, 1432638000, 1432641600, 1432645200, 1432648800, 1432652400, 
    1432656000, 1432659600, 1432666800, 1432670400, 1432674000, 1432677600, 
    1432681200, 1432692000, 1432695600, 1432699200, 1432702800, 1432706400, 
    1432710000, 1432713600, 1432717200, 1432720800, 1432724400, 1432728000, 
    1432731600, 1432735200, 1432738800, 1432742400, 1432746000, 1432749600, 
    1432753200, 1432756800, 1432760400, 1432764000, 1432767600, 1432771200, 
    1432774800, 1432778400, 1432782000, 1432785600, 1432789200, 1432792800, 
    1432796400, 1432800000, 1432803600, 1432807200, 1432810800, 1432814400, 
    1432818000, 1432821600, 1432825200, 1432828800, 1432832400, 1432836000, 
    1432839600, 1432843200, 1432846800, 1432850400, 1432854000, 1432857600, 
    1432861200, 1432864800, 1432868400, 1432872000, 1432875600, 1432879200, 
    1432882800, 1432886400, 1432890000, 1432893600, 1432897200, 1432900800, 
    1432904400, 1432908000, 1432911600, 1432915200, 1432918800, 1432922400, 
    1432926000, 1432929600, 1432933200, 1432936800, 1432940400, 1432944000, 
    1432947600, 1432951200, 1432954800, 1432958400, 1432962000, 1432965600, 
    1432969200, 1432972800, 1432976400, 1432980000, 1432983600, 1432987200, 
    1432990800, 1432994400, 1432998000, 1433001600, 1433005200, 1433008800, 
    1433012400, 1433016000, 1433019600, 1433023200, 1433026800, 1433030400, 
    1433034000, 1433037600, 1433041200, 1433044800, 1433048400, 1433052000, 
    1433055600, 1433059200, 1433062800, 1433066400, 1433070000, 1433073600, 
    1433077200, 1433080800, 1433084400, 1433088000, 1433091600, 1433095200, 
    1433098800, 1433102400, 1433106000, 1433109600, 1433113200, 1433116800, 
    1433120400, 1433124000, 1433127600, 1433131200, 1433134800, 1433138400, 
    1433142000, 1433145600, 1433149200, 1433152800, 1433156400, 1433160000, 
    1433163600, 1433167200, 1433170800, 1433174400, 1433178000, 1433181600, 
    1433185200, 1433188800, 1433192400, 1433196000, 1433199600, 1433203200, 
    1433206800, 1433210400, 1433214000, 1433217600, 1433221200, 1433224800, 
    1433228400, 1433232000, 1433235600, 1433239200, 1433242800, 1433246400, 
    1433250000, 1433253600, 1433257200, 1433260800, 1433264400, 1433268000, 
    1433271600, 1433275200, 1433278800, 1433282400, 1433286000, 1433289600, 
    1433293200, 1433296800, 1433300400, 1433304000, 1433307600, 1433311200, 
    1433314800, 1433318400, 1433322000, 1433325600, 1433329200, 1433332800, 
    1433336400, 1433340000, 1433343600, 1433347200, 1433350800, 1433354400, 
    1433358000, 1433361600, 1433365200, 1433368800, 1433372400, 1433376000, 
    1433379600, 1433383200, 1433386800, 1433390400, 1433394000, 1433397600, 
    1433401200, 1433404800, 1433408400, 1433412000, 1433415600, 1433419200, 
    1433422800, 1433426400, 1433430000, 1433433600, 1433437200, 1433440800, 
    1433444400, 1433448000, 1433451600, 1433455200, 1433458800, 1433462400, 
    1433466000, 1433469600, 1433473200, 1433476800, 1433480400, 1433484000, 
    1433487600, 1433491200, 1433494800, 1433498400, 1433502000, 1433505600, 
    1433509200, 1433512800, 1433516400, 1433520000, 1433523600, 1433527200, 
    1433530800, 1433534400, 1433538000, 1433541600, 1433545200, 1433548800, 
    1433552400, 1433556000, 1433559600, 1433563200, 1433566800, 1433570400, 
    1433574000, 1433577600, 1433581200, 1433584800, 1433588400, 1433592000, 
    1433595600, 1433599200, 1433602800, 1433606400, 1433610000, 1433613600, 
    1433617200, 1433620800, 1433624400, 1433628000, 1433631600, 1433635200, 
    1433638800, 1433642400, 1433646000, 1433649600, 1433653200, 1433656800, 
    1433660400, 1433664000, 1433667600, 1433671200, 1433674800, 1433678400, 
    1433682000, 1433685600, 1433689200, 1433692800, 1433696400, 1433700000, 
    1433703600, 1433707200, 1433710800, 1433714400, 1433718000, 1433721600, 
    1433725200, 1433728800, 1433732400, 1433736000, 1433739600, 1433743200, 
    1433746800, 1433750400, 1433754000, 1433757600, 1433761200, 1433764800, 
    1433768400, 1433772000, 1433775600, 1433779200, 1433782800, 1433786400, 
    1433790000, 1433793600, 1433797200, 1433800800, 1433804400, 1433808000, 
    1433811600, 1433815200, 1433818800, 1433822400, 1433826000, 1433829600, 
    1433833200, 1433836800, 1433840400, 1433844000, 1433847600, 1433851200, 
    1433854800, 1433858400, 1433862000, 1433865600, 1433869200, 1433872800, 
    1433876400, 1433880000, 1433883600, 1433887200, 1433890800, 1433894400, 
    1433898000, 1433901600, 1433905200, 1433908800, 1433912400, 1433916000, 
    1433919600, 1433923200, 1433926800, 1433930400, 1433934000, 1433937600, 
    1433941200, 1433944800, 1433948400, 1433952000, 1433955600, 1433959200, 
    1433962800, 1433966400, 1433970000, 1433973600, 1433977200, 1433980800, 
    1433984400, 1433988000, 1433991600, 1433995200, 1433998800, 1434002400, 
    1434006000, 1434009600, 1434013200, 1434016800, 1434020400, 1434024000, 
    1434027600, 1434031200, 1434034800, 1434038400, 1434042000, 1434045600, 
    1434049200, 1434052800, 1434056400, 1434060000, 1434063600, 1434067200, 
    1434070800, 1434074400, 1434078000, 1434081600, 1434085200, 1434088800, 
    1434092400, 1434096000, 1434099600, 1434103200, 1434106800, 1434110400, 
    1434114000, 1434117600, 1434121200, 1434124800, 1434128400, 1434132000, 
    1434135600, 1434139200, 1434142800, 1434146400, 1434150000, 1434153600, 
    1434157200, 1434160800, 1434164400, 1434168000, 1434171600, 1434175200, 
    1434178800, 1434182400, 1434186000, 1434189600, 1434193200, 1434196800, 
    1434200400, 1434204000, 1434207600, 1434211200, 1434214800, 1434218400, 
    1434222000, 1434225600, 1434229200, 1434232800, 1434236400, 1434240000, 
    1434243600, 1434247200, 1434250800, 1434254400, 1434258000, 1434261600, 
    1434265200, 1434268800, 1434272400, 1434276000, 1434279600, 1434283200, 
    1434286800, 1434290400, 1434294000, 1434297600, 1434301200, 1434304800, 
    1434308400, 1434312000, 1434315600, 1434319200, 1434322800, 1434326400, 
    1434330000, 1434333600, 1434337200, 1434340800, 1434344400, 1434348000, 
    1434351600, 1434355200, 1434358800, 1434362400, 1434366000, 1434369600, 
    1434373200, 1434376800, 1434380400, 1434384000, 1434387600, 1434391200, 
    1434394800, 1434398400, 1434402000, 1434405600, 1434409200, 1434412800, 
    1434416400, 1434420000, 1434423600, 1434427200, 1434430800, 1434434400, 
    1434438000, 1434441600, 1434445200, 1434448800, 1434452400, 1434456000, 
    1434459600, 1434463200, 1434466800, 1434470400, 1434474000, 1434477600, 
    1434481200, 1434484800, 1434488400, 1434492000, 1434495600, 1434499200, 
    1434502800, 1434506400, 1434510000, 1434513600, 1434517200, 1434520800, 
    1434524400, 1434528000, 1434531600, 1434535200, 1434538800, 1434542400, 
    1434546000, 1434549600, 1434553200, 1434556800, 1434560400, 1434564000, 
    1434567600, 1434571200, 1434574800, 1434578400, 1434582000, 1434585600, 
    1434589200, 1434592800, 1434596400, 1434600000, 1434603600, 1434607200, 
    1434610800, 1434614400, 1434618000, 1434621600, 1434625200, 1434628800, 
    1434632400, 1434636000, 1434639600, 1434643200, 1434646800, 1434650400, 
    1434654000, 1434657600, 1434661200, 1434664800, 1434668400, 1434672000, 
    1434675600, 1434679200, 1434682800, 1434686400, 1434690000, 1434693600, 
    1434697200, 1434700800, 1434704400, 1434708000, 1434711600, 1434715200, 
    1434718800, 1434722400, 1434726000, 1434729600, 1434733200, 1434736800, 
    1434740400, 1434744000, 1434747600, 1434751200, 1434754800, 1434758400, 
    1434762000, 1434765600, 1434769200, 1434772800, 1434776400, 1434780000, 
    1434783600, 1434787200, 1434790800, 1434794400, 1434798000, 1434801600, 
    1434805200, 1434808800, 1434812400, 1434816000, 1434819600, 1434823200, 
    1434826800, 1434830400, 1434834000, 1434837600, 1434841200, 1434844800, 
    1434848400, 1434852000, 1434855600, 1434859200, 1434862800, 1434866400, 
    1434870000, 1434873600, 1434877200, 1434880800, 1434884400, 1434888000, 
    1434891600, 1434895200, 1434898800, 1434902400, 1434906000, 1434909600, 
    1434913200, 1434916800, 1434920400, 1434924000, 1434927600, 1434931200, 
    1434934800, 1434938400, 1434942000, 1434945600, 1434949200, 1434952800, 
    1434956400, 1434960000, 1434963600, 1434967200, 1434970800, 1434974400, 
    1434978000, 1434981600, 1434985200, 1434988800, 1434992400, 1434996000, 
    1434999600, 1435003200, 1435006800, 1435010400, 1435014000, 1435017600, 
    1435021200, 1435024800, 1435028400, 1435032000, 1435035600, 1435039200, 
    1435042800, 1435046400, 1435050000, 1435053600, 1435057200, 1435060800, 
    1435064400, 1435068000, 1435071600, 1435075200, 1435078800, 1435082400, 
    1435086000, 1435089600, 1435093200, 1435096800, 1435100400, 1435104000, 
    1435107600, 1435111200, 1435114800, 1435118400, 1435122000, 1435125600, 
    1435129200, 1435132800, 1435136400, 1435140000, 1435143600, 1435147200, 
    1435150800, 1435154400, 1435158000, 1435161600, 1435165200, 1435168800, 
    1435172400, 1435176000, 1435179600, 1435183200, 1435186800, 1435190400, 
    1435194000, 1435197600, 1435201200, 1435204800, 1435208400, 1435212000, 
    1435215600, 1435219200, 1435222800, 1435226400, 1435230000, 1435233600, 
    1435237200, 1435240800, 1435244400, 1435248000, 1435251600, 1435255200, 
    1435258800, 1435262400, 1435266000, 1435269600, 1435273200, 1435276800, 
    1435280400, 1435284000, 1435287600, 1435291200, 1435294800, 1435298400, 
    1435302000, 1435305600, 1435309200, 1435312800, 1435316400, 1435320000, 
    1435323600, 1435327200, 1435330800, 1435334400, 1435338000, 1435341600, 
    1435345200, 1435348800, 1435352400, 1435356000, 1435359600, 1435363200, 
    1435366800, 1435370400, 1435374000, 1435377600, 1435381200, 1435384800, 
    1435388400, 1435392000, 1435395600, 1435399200, 1435402800, 1435406400, 
    1435410000, 1435413600, 1435417200, 1435420800, 1435424400, 1435428000, 
    1435431600, 1435435200, 1435438800, 1435442400, 1435446000, 1435449600, 
    1435453200, 1435456800, 1435460400, 1435464000, 1435467600, 1435471200, 
    1435474800, 1435478400, 1435482000, 1435485600, 1435489200, 1435492800, 
    1435496400, 1435500000, 1435503600, 1435507200, 1435510800, 1435514400, 
    1435518000, 1435521600, 1435525200, 1435528800, 1435532400, 1435536000, 
    1435539600, 1435543200, 1435546800, 1435550400, 1435554000, 1435557600, 
    1435561200, 1435564800, 1435568400, 1435572000, 1435575600, 1435579200, 
    1435582800, 1435586400, 1435590000, 1435593600, 1435597200, 1435600800, 
    1435604400, 1435608000, 1435611600, 1435615200, 1435618800, 1435622400, 
    1435626000, 1435629600, 1435633200, 1435636800, 1435640400, 1435644000, 
    1435647600, 1435651200, 1435654800, 1435658400, 1435662000, 1435665600, 
    1435669200, 1435672800, 1435676400, 1435680000, 1435683600, 1435687200, 
    1435690800, 1435694400, 1435698000, 1435701600, 1435705200, 1435708800, 
    1435712400, 1435716000, 1435719600, 1435723200, 1435726800, 1435730400, 
    1435734000, 1435737600, 1435741200, 1435744800, 1435748400, 1435752000, 
    1435755600, 1435759200, 1435762800, 1435766400, 1435770000, 1435773600, 
    1435777200, 1435780800, 1435784400, 1435788000, 1435791600, 1435795200, 
    1435798800, 1435802400, 1435806000, 1435809600, 1435813200, 1435816800, 
    1435820400, 1435824000, 1435827600, 1435831200, 1435834800, 1435838400, 
    1435842000, 1435845600, 1435849200, 1435852800, 1435856400, 1435860000, 
    1435863600, 1435867200, 1435870800, 1435874400, 1435878000, 1435881600, 
    1435885200, 1435888800, 1435892400, 1435896000, 1435899600, 1435903200, 
    1435906800, 1435910400, 1435914000, 1435917600, 1435921200, 1435924800, 
    1435928400, 1435932000, 1435935600, 1435939200, 1435942800, 1435946400, 
    1435950000, 1435953600, 1435957200, 1435960800, 1435964400, 1435968000, 
    1435971600, 1435975200, 1435978800, 1435982400, 1435986000, 1435989600, 
    1435993200, 1435996800, 1436000400, 1436004000, 1436007600, 1436011200, 
    1436014800, 1436018400, 1436022000, 1436025600, 1436029200, 1436032800, 
    1436036400, 1436040000, 1436043600, 1436047200, 1436050800, 1436054400, 
    1436058000, 1436061600, 1436065200, 1436068800, 1436072400, 1436076000, 
    1436079600, 1436083200, 1436086800, 1436090400, 1436094000, 1436097600, 
    1436101200, 1436104800, 1436108400, 1436112000, 1436115600, 1436119200, 
    1436122800, 1436126400, 1436130000, 1436133600, 1436137200, 1436140800, 
    1436144400, 1436148000, 1436151600, 1436155200, 1436158800, 1436162400, 
    1436166000, 1436169600, 1436173200, 1436176800, 1436180400, 1436184000, 
    1436187600, 1436191200, 1436194800, 1436198400, 1436202000, 1436205600, 
    1436209200, 1436212800, 1436216400, 1436220000, 1436223600, 1436227200, 
    1436230800, 1436234400, 1436238000, 1436241600, 1436245200, 1436248800, 
    1436252400, 1436256000, 1436259600, 1436263200, 1436266800, 1436270400, 
    1436274000, 1436277600, 1436281200, 1436284800, 1436288400, 1436292000, 
    1436295600, 1436299200, 1436302800, 1436306400, 1436310000, 1436313600, 
    1436317200, 1436320800, 1436324400, 1436328000, 1436331600, 1436335200, 
    1436338800, 1436342400, 1436346000, 1436349600, 1436353200, 1436356800, 
    1436360400, 1436364000, 1436367600, 1436371200, 1436374800, 1436378400, 
    1436382000, 1436385600, 1436389200, 1436392800, 1436396400, 1436400000, 
    1436403600, 1436407200, 1436410800, 1436414400, 1436418000, 1436421600, 
    1436425200, 1436428800, 1436432400, 1436436000, 1436439600, 1436443200, 
    1436446800, 1436450400, 1436454000, 1436457600, 1436461200, 1436464800, 
    1436468400, 1436472000, 1436475600, 1436479200, 1436482800, 1436486400, 
    1436490000, 1436493600, 1436497200, 1436500800, 1436504400, 1436508000, 
    1436511600, 1436515200, 1436518800, 1436522400, 1436526000, 1436529600, 
    1436533200, 1436536800, 1436540400, 1436544000, 1436547600, 1436551200, 
    1436554800, 1436558400, 1436562000, 1436565600, 1436569200, 1436572800, 
    1436576400, 1436580000, 1436583600, 1436587200, 1436590800, 1436594400, 
    1436598000, 1436601600, 1436605200, 1436608800, 1436612400, 1436616000, 
    1436619600, 1436623200, 1436626800, 1436630400, 1436634000, 1436637600, 
    1436641200, 1436644800, 1436648400, 1436652000, 1436655600, 1436659200, 
    1436662800, 1436666400, 1436670000, 1436673600, 1436677200, 1436680800, 
    1436684400, 1436688000, 1436691600, 1436695200, 1436698800, 1436702400, 
    1436706000, 1436709600, 1436713200, 1436716800, 1436720400, 1436724000, 
    1436727600, 1436731200, 1436734800, 1436738400, 1436742000, 1436745600, 
    1436749200, 1436752800, 1436756400, 1436760000, 1436763600, 1436767200, 
    1436770800, 1436774400, 1436778000, 1436781600, 1436785200, 1436788800, 
    1436792400, 1436796000, 1436799600, 1436803200, 1436806800, 1436810400, 
    1436814000, 1436817600, 1436821200, 1436824800, 1436828400, 1436832000, 
    1436835600, 1436839200, 1436842800, 1436846400, 1436850000, 1436853600, 
    1436857200, 1436860800, 1436864400, 1436868000, 1436871600, 1436875200, 
    1436878800, 1436882400, 1436886000, 1436889600, 1436893200, 1436896800, 
    1436900400, 1436904000, 1436907600, 1436911200, 1436914800, 1436918400, 
    1436922000, 1436925600, 1436929200, 1436932800, 1436936400, 1436940000, 
    1436943600, 1436947200, 1436950800, 1436954400, 1436958000, 1436961600, 
    1436965200, 1436968800, 1436972400, 1436976000, 1436979600, 1436983200, 
    1436986800, 1436990400, 1436994000, 1436997600, 1437001200, 1437004800, 
    1437008400, 1437012000, 1437015600, 1437019200, 1437022800, 1437026400, 
    1437030000, 1437033600, 1437037200, 1437040800, 1437044400, 1437048000, 
    1437051600, 1437055200, 1437058800, 1437062400, 1437066000, 1437069600, 
    1437073200, 1437076800, 1437080400, 1437084000, 1437087600, 1437091200, 
    1437094800, 1437098400, 1437102000, 1437105600, 1437109200, 1437112800, 
    1437116400, 1437120000, 1437123600, 1437127200, 1437130800, 1437134400, 
    1437138000, 1437141600, 1437145200, 1437148800, 1437152400, 1437156000, 
    1437159600, 1437163200, 1437166800, 1437170400, 1437174000, 1437177600, 
    1437181200, 1437184800, 1437188400, 1437192000, 1437195600, 1437199200, 
    1437202800, 1437206400, 1437210000, 1437213600, 1437217200, 1437220800, 
    1437224400, 1437228000, 1437231600, 1437235200, 1437238800, 1437242400, 
    1437246000, 1437249600, 1437253200, 1437256800, 1437260400, 1437264000, 
    1437267600, 1437271200, 1437274800, 1437278400, 1437282000, 1437285600, 
    1437289200, 1437292800, 1437296400, 1437300000, 1437303600, 1437307200, 
    1437310800, 1437314400, 1437318000, 1437321600, 1437325200, 1437328800, 
    1437332400, 1437336000, 1437339600, 1437343200, 1437346800, 1437350400, 
    1437354000, 1437357600, 1437361200, 1437364800, 1437368400, 1437372000, 
    1437375600, 1437379200, 1437382800, 1437386400, 1437390000, 1437393600, 
    1437397200, 1437400800, 1437404400, 1437408000, 1437411600, 1437415200, 
    1437418800, 1437422400, 1437426000, 1437429600, 1437433200, 1437436800, 
    1437440400, 1437444000, 1437447600, 1437451200, 1437454800, 1437458400, 
    1437462000, 1437465600, 1437469200, 1437472800, 1437476400, 1437480000, 
    1437483600, 1437487200, 1437490800, 1437494400, 1437498000, 1437501600, 
    1437505200, 1437508800, 1437512400, 1437516000, 1437519600, 1437523200, 
    1437526800, 1437530400, 1437534000, 1437537600, 1437541200, 1437544800, 
    1437548400, 1437552000, 1437555600, 1437559200, 1437562800, 1437566400, 
    1437570000, 1437573600, 1437577200, 1437580800, 1437584400, 1437588000, 
    1437591600, 1437595200, 1437598800, 1437602400, 1437606000, 1437609600, 
    1437613200, 1437616800, 1437620400, 1437624000, 1437627600, 1437631200, 
    1437634800, 1437638400, 1437642000, 1437645600, 1437649200, 1437652800, 
    1437656400, 1437660000, 1437663600, 1437667200, 1437670800, 1437674400, 
    1437678000, 1437681600, 1437685200, 1437688800, 1437692400, 1437696000, 
    1437699600, 1437703200, 1437706800, 1437710400, 1437714000, 1437717600, 
    1437721200, 1437724800, 1437728400, 1437732000, 1437735600, 1437739200, 
    1437742800, 1437746400, 1437750000, 1437753600, 1437757200, 1437760800, 
    1437764400, 1437768000, 1437771600, 1437775200, 1437778800, 1437782400, 
    1437786000, 1437789600, 1437793200, 1437796800, 1437800400, 1437804000, 
    1437807600, 1437811200, 1437814800, 1437818400, 1437822000, 1437825600, 
    1437829200, 1437832800, 1437836400, 1437840000, 1437843600, 1437847200, 
    1437850800, 1437854400, 1437858000, 1437861600, 1437865200, 1437868800, 
    1437872400, 1437876000, 1437879600, 1437883200, 1437886800, 1437890400, 
    1437894000, 1437897600, 1437901200, 1437904800, 1437908400, 1437912000, 
    1437915600, 1437919200, 1437922800, 1437926400, 1437930000, 1437933600, 
    1437937200, 1437940800, 1437944400, 1437948000, 1437951600, 1437955200, 
    1437958800, 1437962400, 1437966000, 1437969600, 1437973200, 1437976800, 
    1437980400, 1437984000, 1437987600, 1437991200, 1437994800, 1437998400, 
    1438002000, 1438005600, 1438009200, 1438012800, 1438016400, 1438020000, 
    1438023600, 1438027200, 1438030800, 1438034400, 1438038000, 1438041600, 
    1438045200, 1438048800, 1438052400, 1438056000, 1438059600, 1438063200, 
    1438066800, 1438070400, 1438074000, 1438077600, 1438081200, 1438084800, 
    1438088400, 1438092000, 1438095600, 1438099200, 1438102800, 1438106400, 
    1438110000, 1438113600, 1438117200, 1438120800, 1438124400, 1438128000, 
    1438131600, 1438135200, 1438138800, 1438142400, 1438146000, 1438149600, 
    1438153200, 1438156800, 1438160400, 1438164000, 1438167600, 1438171200, 
    1438174800, 1438178400, 1438182000, 1438185600, 1438189200, 1438192800, 
    1438196400, 1438200000, 1438203600, 1438207200, 1438210800, 1438214400, 
    1438218000, 1438221600, 1438225200, 1438228800, 1438232400, 1438236000, 
    1438239600, 1438243200, 1438246800, 1438250400, 1438254000, 1438257600, 
    1438261200, 1438264800, 1438268400, 1438272000, 1438275600, 1438279200, 
    1438282800, 1438286400, 1438290000, 1438293600, 1438297200, 1438300800, 
    1438304400, 1438308000, 1438311600, 1438315200, 1438318800, 1438322400, 
    1438326000, 1438329600, 1438333200, 1438336800, 1438340400, 1438344000, 
    1438347600, 1438351200, 1438354800, 1438358400, 1438362000, 1438365600, 
    1438369200, 1438372800, 1438376400, 1438380000, 1438383600, 1438387200, 
    1438390800, 1438394400, 1438398000, 1438401600, 1438405200, 1438408800, 
    1438412400, 1438416000, 1438419600, 1438423200, 1438426800, 1438430400, 
    1438434000, 1438437600, 1438441200, 1438444800, 1438448400, 1438452000, 
    1438455600, 1438459200, 1438462800, 1438466400, 1438470000, 1438473600, 
    1438477200, 1438480800, 1438484400, 1438488000, 1438491600, 1438495200, 
    1438498800, 1438502400, 1438506000, 1438509600, 1438513200, 1438516800, 
    1438520400, 1438524000, 1438527600, 1438531200, 1438534800, 1438538400, 
    1438542000, 1438545600, 1438549200, 1438552800, 1438556400, 1438560000, 
    1438563600, 1438567200, 1438570800, 1438574400, 1438578000, 1438581600, 
    1438585200, 1438588800, 1438592400, 1438596000, 1438599600, 1438603200, 
    1438606800, 1438610400, 1438614000, 1438617600, 1438621200, 1438624800, 
    1438628400, 1438632000, 1438635600, 1438639200, 1438642800, 1438646400, 
    1438650000, 1438653600, 1438657200, 1438660800, 1438664400, 1438668000, 
    1438671600, 1438675200, 1438678800, 1438682400, 1438686000, 1438689600, 
    1438693200, 1438696800, 1438700400, 1438704000, 1438707600, 1438711200, 
    1438714800, 1438718400, 1438722000, 1438725600, 1438729200, 1438732800, 
    1438736400, 1438740000, 1438743600, 1438747200, 1438750800, 1438754400, 
    1438758000, 1438761600, 1438765200, 1438768800, 1438772400, 1438776000, 
    1438779600, 1438783200, 1438786800, 1438790400, 1438794000, 1438797600, 
    1438801200, 1438804800, 1438808400, 1438812000, 1438815600, 1438819200, 
    1438822800, 1438826400, 1438830000, 1438833600, 1438837200, 1438840800, 
    1438844400, 1438848000, 1438851600, 1438855200, 1438858800, 1438862400, 
    1438866000, 1438869600, 1438873200, 1438876800, 1438880400, 1438884000, 
    1438887600, 1438891200, 1438894800, 1438898400, 1438902000, 1438905600, 
    1438909200, 1438912800, 1438916400, 1438920000, 1438923600, 1438927200, 
    1438930800, 1438934400, 1438938000, 1438941600, 1438945200, 1438948800, 
    1438952400, 1438956000, 1438959600, 1438963200, 1438966800, 1438970400, 
    1438974000, 1438977600, 1438981200, 1438984800, 1438988400, 1438992000, 
    1438995600, 1438999200, 1439002800, 1439006400, 1439010000, 1439013600, 
    1439017200, 1439020800, 1439024400, 1439028000, 1439031600, 1439035200, 
    1439038800, 1439042400, 1439046000, 1439049600, 1439053200, 1439056800, 
    1439060400, 1439064000, 1439067600, 1439071200, 1439074800, 1439078400, 
    1439082000, 1439085600, 1439089200, 1439092800, 1439096400, 1439100000, 
    1439103600, 1439107200, 1439110800, 1439114400, 1439118000, 1439121600, 
    1439125200, 1439128800, 1439132400, 1439136000, 1439139600, 1439143200, 
    1439146800, 1439150400, 1439154000, 1439157600, 1439161200, 1439164800, 
    1439168400, 1439172000, 1439175600, 1439179200, 1439182800, 1439186400, 
    1439190000, 1439193600, 1439197200, 1439200800, 1439204400, 1439208000, 
    1439211600, 1439215200, 1439218800, 1439222400, 1439226000, 1439229600, 
    1439233200, 1439236800, 1439240400, 1439244000, 1439247600, 1439251200, 
    1439254800, 1439258400, 1439262000, 1439265600, 1439269200, 1439272800, 
    1439276400, 1439280000, 1439283600, 1439287200, 1439290800, 1439294400, 
    1439298000, 1439301600, 1439305200, 1439308800, 1439312400, 1439316000, 
    1439319600, 1439323200, 1439326800, 1439330400, 1439334000, 1439337600, 
    1439341200, 1439344800, 1439348400, 1439352000, 1439355600, 1439359200, 
    1439362800, 1439366400, 1439370000, 1439373600, 1439377200, 1439380800, 
    1439384400, 1439388000, 1439391600, 1439395200, 1439398800, 1439402400, 
    1439406000, 1439409600, 1439413200, 1439416800, 1439420400, 1439424000, 
    1439427600, 1439431200, 1439434800, 1439438400, 1439442000, 1439445600, 
    1439449200, 1439452800, 1439456400, 1439460000, 1439463600, 1439467200, 
    1439470800, 1439474400, 1439478000, 1439481600, 1439485200, 1439488800, 
    1439492400, 1439496000, 1439499600, 1439503200, 1439506800, 1439510400, 
    1439514000, 1439517600, 1439521200, 1439524800, 1439528400, 1439532000, 
    1439535600, 1439539200, 1439542800, 1439546400, 1439550000, 1439553600, 
    1439557200, 1439560800, 1439564400, 1439568000, 1439571600, 1439575200, 
    1439578800, 1439582400, 1439586000, 1439589600, 1439593200, 1439596800, 
    1439600400, 1439604000, 1439607600, 1439611200, 1439614800, 1439618400, 
    1439622000, 1439625600, 1439629200, 1439632800, 1439636400, 1439640000, 
    1439643600, 1439647200, 1439650800, 1439654400, 1439658000, 1439661600, 
    1439665200, 1439668800, 1439672400, 1439676000, 1439679600, 1439683200, 
    1439686800, 1439690400, 1439694000, 1439697600, 1439701200, 1439704800, 
    1439708400, 1439712000, 1439715600, 1439719200, 1439722800, 1439726400, 
    1439730000, 1439733600, 1439737200, 1439740800, 1439744400, 1439748000, 
    1439751600, 1439755200, 1439758800, 1439762400, 1439766000, 1439769600, 
    1439773200, 1439776800, 1439780400, 1439784000, 1439787600, 1439791200, 
    1439794800, 1439798400, 1439802000, 1439805600, 1439809200, 1439812800, 
    1439816400, 1439820000, 1439823600, 1439827200, 1439830800, 1439834400, 
    1439838000, 1439841600, 1439845200, 1439848800, 1439852400, 1439856000, 
    1439859600, 1439863200, 1439866800, 1439870400, 1439874000, 1439877600, 
    1439881200, 1439884800, 1439888400, 1439892000, 1439895600, 1439899200, 
    1439902800, 1439906400, 1439910000, 1439913600, 1439917200, 1439920800, 
    1439924400, 1439928000, 1439931600, 1439935200, 1439938800, 1439942400, 
    1439946000, 1439949600, 1439953200, 1439956800, 1439960400, 1439964000, 
    1439967600, 1439971200, 1439974800, 1439978400, 1439982000, 1439985600, 
    1439989200, 1439992800, 1439996400, 1440000000, 1440003600, 1440007200, 
    1440010800, 1440014400, 1440018000, 1440021600, 1440025200, 1440028800, 
    1440032400, 1440036000, 1440039600, 1440043200, 1440046800, 1440050400, 
    1440054000, 1440057600, 1440061200, 1440064800, 1440068400, 1440072000, 
    1440075600, 1440079200, 1440082800, 1440086400, 1440090000, 1440093600, 
    1440097200, 1440100800, 1440104400, 1440108000, 1440111600, 1440115200, 
    1440118800, 1440122400, 1440126000, 1440129600, 1440133200, 1440136800, 
    1440140400, 1440144000, 1440147600, 1440151200, 1440154800, 1440158400, 
    1440162000, 1440165600, 1440169200, 1440172800, 1440176400, 1440180000, 
    1440183600, 1440187200, 1440190800, 1440194400, 1440198000, 1440201600, 
    1440205200, 1440208800, 1440212400, 1440216000, 1440219600, 1440223200, 
    1440226800, 1440230400, 1440234000, 1440237600, 1440241200, 1440244800, 
    1440248400, 1440252000, 1440255600, 1440259200, 1440262800, 1440266400, 
    1440270000, 1440273600, 1440277200, 1440280800, 1440284400, 1440288000, 
    1440291600, 1440295200, 1440298800, 1440302400, 1440306000, 1440309600, 
    1440313200, 1440316800, 1440320400, 1440324000, 1440327600, 1440331200, 
    1440334800, 1440338400, 1440342000, 1440345600, 1440349200, 1440352800, 
    1440356400, 1440360000, 1440363600, 1440367200, 1440370800, 1440374400, 
    1440378000, 1440381600, 1440385200, 1440388800, 1440392400, 1440396000, 
    1440399600, 1440403200, 1440406800, 1440410400, 1440414000, 1440417600, 
    1440421200, 1440424800, 1440428400, 1440432000, 1440435600, 1440439200, 
    1440442800, 1440446400, 1440450000, 1440453600, 1440457200, 1440460800, 
    1440464400, 1440468000, 1440471600, 1440475200, 1440478800, 1440482400, 
    1440486000, 1440489600, 1440493200, 1440496800, 1440500400, 1440504000, 
    1440507600, 1440511200, 1440514800, 1440518400, 1440522000, 1440525600, 
    1440529200, 1440532800, 1440536400, 1440540000, 1440543600, 1440547200, 
    1440550800, 1440554400, 1440558000, 1440561600, 1440565200, 1440568800, 
    1440572400, 1440576000, 1440579600, 1440583200, 1440586800, 1440590400, 
    1440594000, 1440597600, 1440601200, 1440604800, 1440608400, 1440612000, 
    1440615600, 1440619200, 1440622800, 1440626400, 1440630000, 1440633600, 
    1440637200, 1440640800, 1440644400, 1440648000, 1440651600, 1440655200, 
    1440658800, 1440662400, 1440666000, 1440669600, 1440673200, 1440676800, 
    1440680400, 1440684000, 1440687600, 1440691200, 1440694800, 1440698400, 
    1440702000, 1440705600, 1440709200, 1440712800, 1440716400, 1440720000, 
    1440723600, 1440727200, 1440730800, 1440734400, 1440738000, 1440741600, 
    1440745200, 1440748800, 1440752400, 1440756000, 1440759600, 1440763200, 
    1440766800, 1440770400, 1440774000, 1440777600, 1440781200, 1440784800, 
    1440788400, 1440792000, 1440795600, 1440799200, 1440802800, 1440806400, 
    1440810000, 1440813600, 1440817200, 1440820800, 1440824400, 1440828000, 
    1440831600, 1440835200, 1440838800, 1440842400, 1440846000, 1440849600, 
    1440853200, 1440856800, 1440860400, 1440864000, 1440867600, 1440871200, 
    1440874800, 1440878400, 1440882000, 1440885600, 1440889200, 1440892800, 
    1440896400, 1440900000, 1440903600, 1440907200, 1440910800, 1440914400, 
    1440918000, 1440921600, 1440925200, 1440928800, 1440932400, 1440936000, 
    1440939600, 1440943200, 1440946800, 1440950400, 1440954000, 1440957600, 
    1440961200, 1440964800, 1440968400, 1440972000, 1440975600, 1440979200, 
    1440982800, 1440986400, 1440990000, 1440993600, 1440997200, 1441000800, 
    1441004400, 1441008000, 1441011600, 1441015200, 1441018800, 1441022400, 
    1441026000, 1441029600, 1441033200, 1441036800, 1441040400, 1441044000, 
    1441047600, 1441051200, 1441054800, 1441058400, 1441062000, 1441065600, 
    1441069200, 1441072800, 1441076400, 1441080000, 1441083600, 1441087200, 
    1441090800, 1441094400, 1441098000, 1441101600, 1441105200, 1441108800, 
    1441112400, 1441116000, 1441119600, 1441123200, 1441126800, 1441130400, 
    1441134000, 1441137600, 1441141200, 1441144800, 1441148400, 1441152000, 
    1441155600, 1441159200, 1441162800, 1441166400, 1441170000, 1441173600, 
    1441177200, 1441180800, 1441184400, 1441188000, 1441191600, 1441195200, 
    1441198800, 1441202400, 1441206000, 1441209600, 1441213200, 1441216800, 
    1441220400, 1441224000, 1441227600, 1441231200, 1441234800, 1441238400, 
    1441242000, 1441245600, 1441249200, 1441252800, 1441256400, 1441260000, 
    1441263600, 1441267200, 1441270800, 1441274400, 1441278000, 1441281600, 
    1441285200, 1441288800, 1441292400, 1441296000, 1441299600, 1441303200, 
    1441306800, 1441310400, 1441314000, 1441317600, 1441321200, 1441324800, 
    1441328400, 1441332000, 1441335600, 1441339200, 1441342800, 1441346400, 
    1441350000, 1441353600, 1441357200, 1441360800, 1441364400, 1441368000, 
    1441371600, 1441375200, 1441378800, 1441382400, 1441386000, 1441389600, 
    1441393200, 1441396800, 1441400400, 1441404000, 1441407600, 1441411200, 
    1441414800, 1441418400, 1441422000, 1441425600, 1441429200, 1441432800, 
    1441436400, 1441440000, 1441443600, 1441447200, 1441450800, 1441454400, 
    1441458000, 1441461600, 1441465200, 1441468800, 1441472400, 1441476000, 
    1441479600, 1441483200, 1441486800, 1441490400, 1441494000, 1441497600, 
    1441501200, 1441504800, 1441508400, 1441512000, 1441515600, 1441519200, 
    1441522800, 1441526400, 1441530000, 1441533600, 1441537200, 1441540800, 
    1441544400, 1441548000, 1441551600, 1441555200, 1441558800, 1441562400, 
    1441566000, 1441569600, 1441573200, 1441576800, 1441580400, 1441584000, 
    1441587600, 1441591200, 1441594800, 1441598400, 1441602000, 1441605600, 
    1441609200, 1441612800, 1441616400, 1441620000, 1441623600, 1441627200, 
    1441630800, 1441634400, 1441638000, 1441641600, 1441645200, 1441648800, 
    1441652400, 1441656000, 1441659600, 1441663200, 1441666800, 1441670400, 
    1441674000, 1441677600, 1441681200, 1441684800, 1441688400, 1441692000, 
    1441695600, 1441699200, 1441702800, 1441706400, 1441710000, 1441713600, 
    1441717200, 1441720800, 1441724400, 1441728000, 1441731600, 1441735200, 
    1441738800, 1441742400, 1441746000, 1441749600, 1441753200, 1441756800, 
    1441760400, 1441764000, 1441767600, 1441771200, 1441774800, 1441778400, 
    1441782000, 1441785600, 1441789200, 1441792800, 1441796400, 1441800000, 
    1441803600, 1441807200, 1441810800, 1441814400, 1441818000, 1441821600, 
    1441825200, 1441828800, 1441832400, 1441836000, 1441839600, 1441843200, 
    1441846800, 1441850400, 1441854000, 1441857600, 1441861200, 1441864800, 
    1441868400, 1441872000, 1441875600, 1441879200, 1441882800, 1441886400, 
    1441890000, 1441893600, 1441897200, 1441900800, 1441904400, 1441908000, 
    1441911600, 1441915200, 1441918800, 1441922400, 1441926000, 1441929600, 
    1441933200, 1441936800, 1441940400, 1441944000, 1441947600, 1441951200, 
    1441954800, 1441958400, 1441962000, 1441965600, 1441969200, 1441972800, 
    1441976400, 1441980000, 1441983600, 1441987200, 1441990800, 1441994400, 
    1441998000, 1442001600, 1442005200, 1442008800, 1442012400, 1442016000, 
    1442019600, 1442023200, 1442026800, 1442030400, 1442034000, 1442037600, 
    1442041200, 1442044800, 1442048400, 1442052000, 1442055600, 1442059200, 
    1442062800, 1442066400, 1442070000, 1442073600, 1442077200, 1442080800, 
    1442084400, 1442088000, 1442091600, 1442095200, 1442098800, 1442102400, 
    1442106000, 1442109600, 1442113200, 1442116800, 1442120400, 1442124000, 
    1442127600, 1442131200, 1442134800, 1442138400, 1442142000, 1442145600, 
    1442149200, 1442152800, 1442156400, 1442160000, 1442163600, 1442167200, 
    1442170800, 1442174400, 1442178000, 1442181600, 1442185200, 1442188800, 
    1442192400, 1442196000, 1442199600, 1442203200, 1442206800, 1442210400, 
    1442214000, 1442217600, 1442221200, 1442224800, 1442228400, 1442232000, 
    1442235600, 1442239200, 1442242800, 1442246400, 1442250000, 1442253600, 
    1442257200, 1442260800, 1442264400, 1442268000, 1442271600, 1442275200, 
    1442278800, 1442282400, 1442286000, 1442289600, 1442293200, 1442296800, 
    1442300400, 1442304000, 1442307600, 1442311200, 1442314800, 1442318400, 
    1442322000, 1442325600, 1442329200, 1442332800, 1442336400, 1442340000, 
    1442343600, 1442347200, 1442350800, 1442354400, 1442358000, 1442361600, 
    1442365200, 1442368800, 1442372400, 1442376000, 1442379600, 1442383200, 
    1442386800, 1442390400, 1442394000, 1442397600, 1442401200, 1442404800, 
    1442408400, 1442412000, 1442415600, 1442419200, 1442422800, 1442426400, 
    1442430000, 1442433600, 1442437200, 1442440800, 1442444400, 1442448000, 
    1442451600, 1442455200, 1442458800, 1442462400, 1442466000, 1442469600, 
    1442473200, 1442476800, 1442480400, 1442484000, 1442487600, 1442491200, 
    1442494800, 1442498400, 1442502000, 1442505600, 1442509200, 1442512800, 
    1442516400, 1442520000, 1442523600, 1442527200, 1442530800, 1442534400, 
    1442538000, 1442541600, 1442545200, 1442548800, 1442552400, 1442556000, 
    1442559600, 1442563200, 1442566800, 1442570400, 1442574000, 1442577600, 
    1442581200, 1442584800, 1442588400, 1442592000, 1442595600, 1442599200, 
    1442602800, 1442606400, 1442610000, 1442613600, 1442617200, 1442620800, 
    1442624400, 1442628000, 1442631600, 1442635200, 1442638800, 1442642400, 
    1442646000, 1442649600, 1442653200, 1442656800, 1442660400, 1442664000, 
    1442667600, 1442671200, 1442674800, 1442678400, 1442682000, 1442685600, 
    1442689200, 1442692800, 1442696400, 1442700000, 1442703600, 1442707200, 
    1442710800, 1442714400, 1442718000, 1442721600, 1442725200, 1442728800, 
    1442732400, 1442736000, 1442739600, 1442743200, 1442746800, 1442750400, 
    1442754000, 1442757600, 1442761200, 1442764800, 1442768400, 1442772000, 
    1442775600, 1442779200, 1442782800, 1442786400, 1442790000, 1442793600, 
    1442797200, 1442800800, 1442804400, 1442808000, 1442811600, 1442815200, 
    1442818800, 1442822400, 1442826000, 1442829600, 1442833200, 1442836800, 
    1442840400, 1442844000, 1442847600, 1442851200, 1442854800, 1442858400, 
    1442862000, 1442865600, 1442869200, 1442872800, 1442876400, 1442880000, 
    1442883600, 1442887200, 1442890800, 1442894400, 1442898000, 1442901600, 
    1442905200, 1442908800, 1442912400, 1442916000, 1442919600, 1442923200, 
    1442926800, 1442930400, 1442934000, 1442937600, 1442941200, 1442944800, 
    1442948400, 1442952000, 1442955600, 1442959200, 1442962800, 1442966400, 
    1442970000, 1442973600, 1442977200, 1442980800, 1442984400, 1442988000, 
    1442991600, 1442995200, 1442998800, 1443002400, 1443006000, 1443009600, 
    1443013200, 1443016800, 1443020400, 1443024000, 1443027600, 1443031200, 
    1443034800, 1443038400, 1443042000, 1443045600, 1443049200, 1443052800, 
    1443056400, 1443060000, 1443063600, 1443067200, 1443070800, 1443074400, 
    1443078000, 1443081600, 1443085200, 1443088800, 1443092400, 1443096000, 
    1443099600, 1443103200, 1443106800, 1443110400, 1443114000, 1443117600, 
    1443121200, 1443124800, 1443128400, 1443132000, 1443135600, 1443139200, 
    1443142800, 1443146400, 1443150000, 1443153600, 1443157200, 1443160800, 
    1443164400, 1443168000, 1443171600, 1443175200, 1443178800, 1443182400, 
    1443186000, 1443189600, 1443193200, 1443196800, 1443200400, 1443204000, 
    1443207600, 1443211200, 1443214800, 1443218400, 1443222000, 1443225600, 
    1443229200, 1443232800, 1443236400, 1443240000, 1443243600, 1443247200, 
    1443250800, 1443254400, 1443258000, 1443261600, 1443265200, 1443268800, 
    1443272400, 1443276000, 1443279600, 1443283200, 1443286800, 1443290400, 
    1443294000, 1443297600, 1443301200, 1443304800, 1443308400, 1443312000, 
    1443315600, 1443319200, 1443322800, 1443326400, 1443330000, 1443333600, 
    1443337200, 1443340800, 1443344400, 1443348000, 1443351600, 1443355200, 
    1443358800, 1443362400, 1443366000, 1443369600, 1443373200, 1443376800, 
    1443380400, 1443384000, 1443387600, 1443391200, 1443394800, 1443398400, 
    1443402000, 1443405600, 1443409200, 1443412800, 1443416400, 1443420000, 
    1443423600, 1443427200, 1443430800, 1443434400, 1443438000, 1443441600, 
    1443445200, 1443448800, 1443452400, 1443456000, 1443459600, 1443463200, 
    1443466800, 1443470400, 1443474000, 1443477600, 1443481200, 1443484800, 
    1443488400, 1443492000, 1443495600, 1443499200, 1443502800, 1443506400, 
    1443510000, 1443513600, 1443517200, 1443520800, 1443524400, 1443528000, 
    1443531600, 1443535200, 1443538800, 1443542400, 1443546000, 1443549600, 
    1443553200, 1443556800, 1443560400, 1443564000, 1443567600, 1443571200, 
    1443574800, 1443578400, 1443582000, 1443585600, 1443589200, 1443592800, 
    1443596400, 1443600000, 1443603600, 1443607200, 1443610800, 1443614400, 
    1443618000, 1443621600, 1443625200, 1443628800, 1443632400, 1443636000, 
    1443639600, 1443643200, 1443646800, 1443650400, 1443654000, 1443657600, 
    1443661200, 1443664800, 1443668400, 1443672000, 1443675600, 1443679200, 
    1443682800, 1443686400, 1443690000, 1443693600, 1443697200, 1443700800, 
    1443704400, 1443708000, 1443711600, 1443715200, 1443718800, 1443722400, 
    1443726000, 1443729600, 1443733200, 1443736800, 1443740400, 1443744000, 
    1443747600, 1443751200, 1443754800, 1443758400, 1443762000, 1443765600, 
    1443769200, 1443772800, 1443776400, 1443780000, 1443783600, 1443787200, 
    1443790800, 1443794400, 1443798000, 1443801600, 1443805200, 1443808800, 
    1443812400, 1443816000, 1443819600, 1443823200, 1443826800, 1443830400, 
    1443834000, 1443837600, 1443841200, 1443844800, 1443848400, 1443852000, 
    1443855600, 1443859200, 1443862800, 1443866400, 1443870000, 1443873600, 
    1443877200, 1443880800, 1443884400, 1443888000, 1443891600, 1443895200, 
    1443898800, 1443902400, 1443906000, 1443909600, 1443913200, 1443916800, 
    1443920400, 1443924000, 1443927600, 1443931200, 1443934800, 1443938400, 
    1443942000, 1443945600, 1443949200, 1443952800, 1443956400, 1443960000, 
    1443963600, 1443967200, 1443970800, 1443974400, 1443978000, 1443981600, 
    1443985200, 1443988800, 1443992400, 1443996000, 1443999600, 1444003200, 
    1444006800, 1444010400, 1444014000, 1444017600, 1444021200, 1444024800, 
    1444028400, 1444032000, 1444035600, 1444039200, 1444042800, 1444046400, 
    1444050000, 1444053600, 1444057200, 1444060800, 1444064400, 1444068000, 
    1444071600, 1444075200, 1444078800, 1444082400, 1444086000, 1444089600, 
    1444093200, 1444096800, 1444100400, 1444104000, 1444107600, 1444111200, 
    1444114800, 1444118400, 1444122000, 1444125600, 1444129200, 1444132800, 
    1444136400, 1444140000, 1444143600, 1444147200, 1444150800, 1444154400, 
    1444158000, 1444161600, 1444165200, 1444168800, 1444172400, 1444176000, 
    1444179600, 1444183200, 1444186800, 1444190400, 1444194000, 1444197600, 
    1444201200, 1444204800, 1444208400, 1444212000, 1444215600, 1444219200, 
    1444222800, 1444226400, 1444230000, 1444233600, 1444237200, 1444240800, 
    1444244400, 1444248000, 1444251600, 1444255200, 1444258800, 1444262400, 
    1444266000, 1444269600, 1444273200, 1444276800, 1444280400, 1444284000, 
    1444287600, 1444291200, 1444294800, 1444298400, 1444302000, 1444305600, 
    1444309200, 1444312800, 1444316400, 1444320000, 1444323600, 1444327200, 
    1444330800, 1444334400, 1444338000, 1444341600, 1444345200, 1444348800, 
    1444352400, 1444356000, 1444359600, 1444363200, 1444366800, 1444370400, 
    1444374000, 1444377600, 1444381200, 1444384800, 1444388400, 1444392000, 
    1444395600, 1444399200, 1444402800, 1444406400, 1444410000, 1444413600, 
    1444417200, 1444420800, 1444424400, 1444428000, 1444431600, 1444435200, 
    1444438800, 1444442400, 1444446000, 1444449600, 1444453200, 1444456800, 
    1444460400, 1444464000, 1444467600, 1444471200, 1444474800, 1444478400, 
    1444482000, 1444485600, 1444489200, 1444492800, 1444496400, 1444500000, 
    1444503600, 1444507200, 1444510800, 1444514400, 1444518000, 1444521600, 
    1444525200, 1444528800, 1444532400, 1444536000, 1444539600, 1444543200, 
    1444546800, 1444550400, 1444554000, 1444557600, 1444561200, 1444564800, 
    1444568400, 1444572000, 1444575600, 1444579200, 1444582800, 1444586400, 
    1444590000, 1444593600, 1444597200, 1444600800, 1444604400, 1444608000, 
    1444611600, 1444615200, 1444618800, 1444622400, 1444626000, 1444629600, 
    1444633200, 1444636800, 1444640400, 1444644000, 1444647600, 1444651200, 
    1444654800, 1444658400, 1444662000, 1444665600, 1444669200, 1444672800, 
    1444676400, 1444680000, 1444683600, 1444687200, 1444690800, 1444694400, 
    1444698000, 1444701600, 1444705200, 1444708800, 1444712400, 1444716000, 
    1444719600, 1444723200, 1444726800, 1444730400, 1444734000, 1444737600, 
    1444741200, 1444744800, 1444748400, 1444752000, 1444755600, 1444759200, 
    1444762800, 1444766400, 1444770000, 1444773600, 1444777200, 1444780800, 
    1444784400, 1444788000, 1444791600, 1444795200, 1444798800, 1444802400, 
    1444806000, 1444809600, 1444813200, 1444816800, 1444820400, 1444824000, 
    1444827600, 1444831200, 1444834800, 1444838400, 1444842000, 1444845600, 
    1444849200, 1444852800, 1444856400, 1444860000, 1444863600, 1444867200, 
    1444870800, 1444874400, 1444878000, 1444881600, 1444885200, 1444888800, 
    1444892400, 1444896000, 1444899600, 1444903200, 1444906800, 1444910400, 
    1444914000, 1444917600, 1444921200, 1444924800, 1444928400, 1444932000, 
    1444935600, 1444939200, 1444942800, 1444946400, 1444950000, 1444953600, 
    1444957200, 1444960800, 1444964400, 1444968000, 1444971600, 1444975200, 
    1444978800, 1444982400, 1444986000, 1444989600, 1444993200, 1444996800, 
    1445000400, 1445004000, 1445007600, 1445011200, 1445014800, 1445018400, 
    1445022000, 1445025600, 1445029200, 1445032800, 1445036400, 1445040000, 
    1445043600, 1445047200, 1445050800, 1445054400, 1445058000, 1445061600, 
    1445065200, 1445068800, 1445072400, 1445076000, 1445079600, 1445083200, 
    1445086800, 1445090400, 1445094000, 1445097600, 1445101200, 1445104800, 
    1445108400, 1445112000, 1445115600, 1445119200, 1445122800, 1445126400, 
    1445130000, 1445133600, 1445137200, 1445140800, 1445144400, 1445148000, 
    1445151600, 1445155200, 1445158800, 1445162400, 1445166000, 1445169600, 
    1445173200, 1445176800, 1445180400, 1445184000, 1445187600, 1445191200, 
    1445194800, 1445198400, 1445202000, 1445205600, 1445209200, 1445212800, 
    1445216400, 1445220000, 1445223600, 1445227200, 1445230800, 1445234400, 
    1445238000, 1445241600, 1445245200, 1445248800, 1445252400, 1445256000, 
    1445259600, 1445263200, 1445266800, 1445270400, 1445274000, 1445277600, 
    1445281200, 1445284800, 1445288400, 1445292000, 1445295600, 1445299200, 
    1445302800, 1445306400, 1445310000, 1445313600, 1445317200, 1445320800, 
    1445324400, 1445328000, 1445331600, 1445335200, 1445338800, 1445342400, 
    1445346000, 1445349600, 1445353200, 1445356800, 1445360400, 1445364000, 
    1445367600, 1445371200, 1445374800, 1445378400, 1445382000, 1445385600, 
    1445389200, 1445392800, 1445396400, 1445400000, 1445403600, 1445407200, 
    1445410800, 1445414400, 1445418000, 1445421600, 1445425200, 1445428800, 
    1445432400, 1445436000, 1445439600, 1445443200, 1445446800, 1445450400, 
    1445454000, 1445457600, 1445461200, 1445464800, 1445468400, 1445472000, 
    1445475600, 1445479200, 1445482800, 1445486400, 1445490000, 1445493600, 
    1445497200, 1445500800, 1445504400, 1445508000, 1445511600, 1445515200, 
    1445518800, 1445522400, 1445526000, 1445529600, 1445533200, 1445536800, 
    1445540400, 1445544000, 1445547600, 1445551200, 1445554800, 1445558400, 
    1445562000, 1445565600, 1445569200, 1445572800, 1445576400, 1445580000, 
    1445583600, 1445587200, 1445590800, 1445594400, 1445598000, 1445601600, 
    1445605200, 1445608800, 1445612400, 1445616000, 1445619600, 1445623200, 
    1445626800, 1445630400, 1445634000, 1445637600, 1445641200, 1445644800, 
    1445648400, 1445652000, 1445655600, 1445659200, 1445662800, 1445666400, 
    1445670000, 1445673600, 1445677200, 1445680800, 1445684400, 1445688000, 
    1445691600, 1445695200, 1445698800, 1445702400, 1445706000, 1445709600, 
    1445713200, 1445716800, 1445720400, 1445724000, 1445727600, 1445731200, 
    1445734800, 1445738400, 1445742000, 1445745600, 1445749200, 1445752800, 
    1445756400, 1445760000, 1445763600, 1445767200, 1445770800, 1445774400, 
    1445778000, 1445781600, 1445785200, 1445788800, 1445792400, 1445796000, 
    1445799600, 1445803200, 1445806800, 1445810400, 1445814000, 1445817600, 
    1445821200, 1445824800, 1445828400, 1445832000, 1445835600, 1445839200, 
    1445842800, 1445846400, 1445850000, 1445853600, 1445857200, 1445860800, 
    1445864400, 1445868000, 1445871600, 1445875200, 1445878800, 1445882400, 
    1445886000, 1445889600, 1445893200, 1445896800, 1445900400, 1445904000, 
    1445907600, 1445911200, 1445914800, 1445918400, 1445922000, 1445925600, 
    1445929200, 1445932800, 1445936400, 1445940000, 1445943600, 1445947200, 
    1445950800, 1445954400, 1445958000, 1445961600, 1445965200, 1445968800, 
    1445972400, 1445976000, 1445979600, 1445983200, 1445986800, 1445990400, 
    1445994000, 1445997600, 1446001200, 1446004800, 1446008400, 1446012000, 
    1446015600, 1446019200, 1446022800, 1446026400, 1446030000, 1446033600, 
    1446037200, 1446040800, 1446044400, 1446048000, 1446051600, 1446055200, 
    1446058800, 1446062400, 1446066000, 1446069600, 1446073200, 1446076800, 
    1446080400, 1446084000, 1446087600, 1446091200, 1446094800, 1446098400, 
    1446102000, 1446105600, 1446109200, 1446112800, 1446116400, 1446120000, 
    1446123600, 1446127200, 1446130800, 1446134400, 1446138000, 1446141600, 
    1446145200, 1446148800, 1446152400, 1446156000, 1446159600, 1446163200, 
    1446166800, 1446170400, 1446174000, 1446177600, 1446181200, 1446184800, 
    1446188400, 1446192000, 1446195600, 1446199200, 1446202800, 1446206400, 
    1446210000, 1446213600, 1446217200, 1446220800, 1446224400, 1446228000, 
    1446231600, 1446235200, 1446238800, 1446242400, 1446246000, 1446249600, 
    1446253200, 1446256800, 1446260400, 1446264000, 1446267600, 1446271200, 
    1446274800, 1446278400, 1446282000, 1446285600, 1446289200, 1446292800, 
    1446296400, 1446300000, 1446303600, 1446307200, 1446310800, 1446314400, 
    1446318000, 1446321600, 1446325200, 1446328800, 1446332400, 1446336000, 
    1446339600, 1446343200, 1446346800, 1446350400, 1446354000, 1446357600, 
    1446361200, 1446364800, 1446368400, 1446372000, 1446375600, 1446379200, 
    1446382800, 1446386400, 1446390000, 1446393600, 1446397200, 1446400800, 
    1446404400, 1446408000, 1446411600, 1446415200, 1446418800, 1446422400, 
    1446426000, 1446429600, 1446433200, 1446436800, 1446440400, 1446444000, 
    1446447600, 1446451200, 1446454800, 1446458400, 1446462000, 1446465600, 
    1446469200, 1446472800, 1446476400, 1446480000, 1446483600, 1446487200, 
    1446490800, 1446494400, 1446498000, 1446501600, 1446505200, 1446508800, 
    1446512400, 1446516000, 1446519600, 1446523200, 1446526800, 1446530400, 
    1446534000, 1446537600, 1446541200, 1446544800, 1446548400, 1446552000, 
    1446555600, 1446559200, 1446562800, 1446566400, 1446570000, 1446573600, 
    1446577200, 1446580800, 1446584400, 1446588000, 1446591600, 1446595200, 
    1446598800, 1446602400, 1446606000, 1446609600, 1446613200, 1446616800, 
    1446620400, 1446624000, 1446627600, 1446631200, 1446634800, 1446638400, 
    1446642000, 1446645600, 1446649200, 1446652800, 1446656400, 1446660000, 
    1446663600, 1446667200, 1446670800, 1446674400, 1446678000, 1446681600, 
    1446685200, 1446688800, 1446692400, 1446696000, 1446699600, 1446703200, 
    1446706800, 1446710400, 1446714000, 1446717600, 1446721200, 1446724800, 
    1446728400, 1446732000, 1446735600, 1446739200, 1446742800, 1446746400, 
    1446750000, 1446753600, 1446757200, 1446760800, 1446764400, 1446768000, 
    1446771600, 1446775200, 1446778800, 1446782400, 1446786000, 1446789600, 
    1446793200, 1446796800, 1446800400, 1446804000, 1446807600, 1446811200, 
    1446814800, 1446818400, 1446822000, 1446825600, 1446829200, 1446832800, 
    1446836400, 1446840000, 1446843600, 1446847200, 1446850800, 1446854400, 
    1446858000, 1446861600, 1446865200, 1446868800, 1446872400, 1446876000, 
    1446879600, 1446883200, 1446886800, 1446890400, 1446894000, 1446897600, 
    1446901200, 1446904800, 1446908400, 1446912000, 1446915600, 1446919200, 
    1446922800, 1446926400, 1446930000, 1446933600, 1446937200, 1446940800, 
    1446944400, 1446948000, 1446951600, 1446955200, 1446958800, 1446962400, 
    1446966000, 1446969600, 1446973200, 1446976800, 1446980400, 1446984000, 
    1446987600, 1446991200, 1446994800, 1446998400, 1447002000, 1447005600, 
    1447009200, 1447012800, 1447016400, 1447020000, 1447023600, 1447027200, 
    1447030800, 1447034400, 1447038000, 1447041600, 1447045200, 1447048800, 
    1447052400, 1447056000, 1447059600, 1447063200, 1447066800, 1447070400, 
    1447074000, 1447077600, 1447081200, 1447084800, 1447088400, 1447092000, 
    1447095600, 1447099200, 1447102800, 1447106400, 1447110000, 1447113600, 
    1447117200, 1447120800, 1447124400, 1447128000, 1447131600, 1447135200, 
    1447138800, 1447142400, 1447146000, 1447149600, 1447153200, 1447156800, 
    1447160400, 1447164000, 1447167600, 1447171200, 1447174800, 1447178400, 
    1447182000, 1447185600, 1447189200, 1447192800, 1447196400, 1447200000, 
    1447203600, 1447207200, 1447210800, 1447214400, 1447218000, 1447221600, 
    1447225200, 1447228800, 1447232400, 1447236000, 1447239600, 1447243200, 
    1447246800, 1447250400, 1447254000, 1447257600, 1447261200, 1447264800, 
    1447268400, 1447272000, 1447275600, 1447279200, 1447282800, 1447286400, 
    1447290000, 1447293600, 1447297200, 1447300800, 1447304400, 1447308000, 
    1447311600, 1447315200, 1447318800, 1447322400, 1447326000, 1447329600, 
    1447333200, 1447336800, 1447340400, 1447344000, 1447347600, 1447351200, 
    1447354800, 1447358400, 1447362000, 1447365600, 1447369200, 1447372800, 
    1447376400, 1447380000, 1447383600, 1447387200, 1447390800, 1447394400, 
    1447398000, 1447401600, 1447405200, 1447408800, 1447412400, 1447416000, 
    1447419600, 1447423200, 1447426800, 1447430400, 1447434000, 1447437600, 
    1447441200, 1447444800, 1447448400, 1447452000, 1447455600, 1447459200, 
    1447462800, 1447466400, 1447470000, 1447473600, 1447477200, 1447480800, 
    1447484400, 1447488000, 1447491600, 1447495200, 1447498800, 1447502400, 
    1447506000, 1447509600, 1447513200, 1447516800, 1447520400, 1447524000, 
    1447527600, 1447531200, 1447534800, 1447538400, 1447542000, 1447545600, 
    1447549200, 1447552800, 1447556400, 1447560000, 1447563600, 1447567200, 
    1447570800, 1447574400, 1447578000, 1447581600, 1447585200, 1447588800, 
    1447592400, 1447596000, 1447599600, 1447603200, 1447606800, 1447610400, 
    1447614000, 1447617600, 1447621200, 1447624800, 1447628400, 1447632000, 
    1447635600, 1447639200, 1447642800, 1447646400, 1447650000, 1447653600, 
    1447657200, 1447660800, 1447664400, 1447668000, 1447671600, 1447675200, 
    1447678800, 1447682400, 1447686000, 1447689600, 1447693200, 1447696800, 
    1447700400, 1447704000, 1447707600, 1447711200, 1447714800, 1447718400, 
    1447722000, 1447725600, 1447729200, 1447732800, 1447736400, 1447740000, 
    1447743600, 1447747200, 1447750800, 1447754400, 1447758000, 1447761600, 
    1447765200, 1447768800, 1447772400, 1447776000, 1447779600, 1447783200, 
    1447786800, 1447790400, 1447794000, 1447797600, 1447801200, 1447804800, 
    1447808400, 1447812000, 1447815600, 1447819200, 1447822800, 1447826400, 
    1447830000, 1447833600, 1447837200, 1447840800, 1447844400, 1447848000, 
    1447851600, 1447855200, 1447858800, 1447862400, 1447866000, 1447869600, 
    1447873200, 1447876800, 1447880400, 1447884000, 1447887600, 1447891200, 
    1447894800, 1447898400, 1447902000, 1447905600, 1447909200, 1447912800, 
    1447916400, 1447920000, 1447923600, 1447927200, 1447930800, 1447934400, 
    1447938000, 1447941600, 1447945200, 1447948800, 1447952400, 1447956000, 
    1447959600, 1447963200, 1447966800, 1447970400, 1447974000, 1447977600, 
    1447981200, 1447984800, 1447988400, 1447992000, 1447995600, 1447999200, 
    1448002800, 1448006400, 1448010000, 1448013600, 1448017200, 1448020800, 
    1448024400, 1448028000, 1448031600, 1448035200, 1448038800, 1448042400, 
    1448046000, 1448049600, 1448053200, 1448056800, 1448060400, 1448064000, 
    1448067600, 1448071200, 1448074800, 1448078400, 1448082000, 1448085600, 
    1448089200, 1448092800, 1448096400, 1448100000, 1448103600, 1448107200, 
    1448110800, 1448114400, 1448118000, 1448121600, 1448125200, 1448128800, 
    1448132400, 1448136000, 1448139600, 1448143200, 1448146800, 1448150400, 
    1448154000, 1448157600, 1448161200, 1448164800, 1448168400, 1448172000, 
    1448175600, 1448179200, 1448182800, 1448186400, 1448190000, 1448193600, 
    1448197200, 1448200800, 1448204400, 1448208000, 1448211600, 1448215200, 
    1448218800, 1448222400, 1448226000, 1448229600, 1448233200, 1448236800, 
    1448240400, 1448244000, 1448247600, 1448251200, 1448254800, 1448258400, 
    1448262000, 1448265600, 1448269200, 1448272800, 1448276400, 1448280000, 
    1448283600, 1448287200, 1448290800, 1448294400, 1448298000, 1448301600, 
    1448305200, 1448308800, 1448312400, 1448316000, 1448319600, 1448323200, 
    1448326800, 1448330400, 1448334000, 1448337600, 1448341200, 1448344800, 
    1448348400, 1448352000, 1448355600, 1448359200, 1448362800, 1448366400, 
    1448370000, 1448373600, 1448377200, 1448380800, 1448384400, 1448388000, 
    1448391600, 1448395200, 1448398800, 1448402400, 1448406000, 1448409600, 
    1448413200, 1448416800, 1448420400, 1448424000, 1448427600, 1448431200, 
    1448434800, 1448438400, 1448442000, 1448445600, 1448449200, 1448452800, 
    1448456400, 1448460000, 1448463600, 1448467200, 1448470800, 1448474400, 
    1448478000, 1448481600, 1448485200, 1448488800, 1448492400, 1448496000, 
    1448499600, 1448503200, 1448506800, 1448510400, 1448514000, 1448517600, 
    1448521200, 1448524800, 1448528400, 1448532000, 1448535600, 1448539200, 
    1448542800, 1448546400, 1448550000, 1448553600, 1448557200, 1448560800, 
    1448564400, 1448568000, 1448571600, 1448575200, 1448578800, 1448582400, 
    1448586000, 1448589600, 1448593200, 1448596800, 1448600400, 1448604000, 
    1448607600, 1448611200, 1448614800, 1448618400, 1448622000, 1448625600, 
    1448629200, 1448632800, 1448636400, 1448640000, 1448643600, 1448647200, 
    1448650800, 1448654400, 1448658000, 1448661600, 1448665200, 1448668800, 
    1448672400, 1448676000, 1448679600, 1448683200, 1448686800, 1448690400, 
    1448694000, 1448697600, 1448701200, 1448704800, 1448708400, 1448712000, 
    1448715600, 1448719200, 1448722800, 1448726400, 1448730000, 1448733600, 
    1448737200, 1448740800, 1448744400, 1448748000, 1448751600, 1448755200, 
    1448758800, 1448762400, 1448766000, 1448769600, 1448773200, 1448776800, 
    1448780400, 1448784000, 1448787600, 1448791200, 1448794800, 1448798400, 
    1448802000, 1448805600, 1448809200, 1448812800, 1448816400, 1448820000, 
    1448823600, 1448827200, 1448830800, 1448834400, 1448838000, 1448841600, 
    1448845200, 1448848800, 1448852400, 1448856000, 1448859600, 1448863200, 
    1448866800, 1448870400, 1448874000, 1448877600, 1448881200, 1448884800, 
    1448888400, 1448892000, 1448895600, 1448899200, 1448902800, 1448906400, 
    1448910000, 1448913600, 1448917200, 1448920800, 1448924400, 1448928000, 
    1448931600, 1448935200, 1448938800, 1448942400, 1448946000, 1448949600, 
    1448953200, 1448956800, 1448960400, 1448964000, 1448967600, 1448971200, 
    1448974800, 1448978400, 1448982000, 1448985600, 1448989200, 1448992800, 
    1448996400, 1449000000, 1449003600, 1449007200, 1449010800, 1449014400, 
    1449018000, 1449021600, 1449025200, 1449028800, 1449032400, 1449036000, 
    1449039600, 1449043200, 1449046800, 1449050400, 1449054000, 1449057600, 
    1449061200, 1449064800, 1449068400, 1449072000, 1449075600, 1449079200, 
    1449082800, 1449086400, 1449090000, 1449093600, 1449097200, 1449100800, 
    1449104400, 1449108000, 1449111600, 1449115200, 1449118800, 1449122400, 
    1449126000, 1449129600, 1449133200, 1449136800, 1449140400, 1449144000, 
    1449147600, 1449151200, 1449154800, 1449158400, 1449162000, 1449165600, 
    1449169200, 1449172800, 1449176400, 1449180000, 1449183600, 1449187200, 
    1449190800, 1449194400, 1449198000, 1449201600, 1449205200, 1449208800, 
    1449212400, 1449216000, 1449219600, 1449223200, 1449226800, 1449230400, 
    1449234000, 1449237600, 1449241200, 1449244800, 1449248400, 1449252000, 
    1449255600, 1449259200, 1449262800, 1449266400, 1449270000, 1449273600, 
    1449277200, 1449280800, 1449284400, 1449288000, 1449291600, 1449295200, 
    1449298800, 1449302400, 1449306000, 1449309600, 1449313200, 1449316800, 
    1449320400, 1449324000, 1449327600, 1449331200, 1449334800, 1449338400, 
    1449342000, 1449345600, 1449349200, 1449352800, 1449356400, 1449360000, 
    1449363600, 1449367200, 1449370800, 1449374400, 1449378000, 1449381600, 
    1449385200, 1449388800, 1449392400, 1449396000, 1449399600, 1449403200, 
    1449406800, 1449410400, 1449414000, 1449417600, 1449421200, 1449424800, 
    1449428400, 1449432000, 1449435600, 1449439200, 1449442800, 1449446400, 
    1449450000, 1449453600, 1449457200, 1449460800, 1449464400, 1449468000, 
    1449471600, 1449475200, 1449478800, 1449482400, 1449486000, 1449489600, 
    1449493200, 1449496800, 1449500400, 1449504000, 1449507600, 1449511200, 
    1449514800, 1449518400, 1449522000, 1449525600, 1449529200, 1449532800, 
    1449536400, 1449540000, 1449543600, 1449547200, 1449550800, 1449554400, 
    1449558000, 1449561600, 1449565200, 1449568800, 1449572400, 1449576000, 
    1449579600, 1449583200, 1449586800, 1449590400, 1449594000, 1449597600, 
    1449601200, 1449604800, 1449608400, 1449612000, 1449615600, 1449619200, 
    1449622800, 1449626400, 1449630000, 1449633600, 1449637200, 1449640800, 
    1449644400, 1449648000, 1449651600, 1449655200, 1449658800, 1449662400, 
    1449666000, 1449669600, 1449673200, 1449676800, 1449680400, 1449684000, 
    1449687600, 1449691200, 1449694800, 1449698400, 1449702000, 1449705600, 
    1449709200, 1449712800, 1449716400, 1449720000, 1449723600, 1449727200, 
    1449730800, 1449734400, 1449738000, 1449741600, 1449745200, 1449748800, 
    1449752400, 1449756000, 1449759600, 1449763200, 1449766800, 1449770400, 
    1449774000, 1449777600, 1449781200, 1449784800, 1449788400, 1449792000, 
    1449795600, 1449799200, 1449802800, 1449806400, 1449810000, 1449813600, 
    1449817200, 1449820800, 1449824400, 1449828000, 1449831600, 1449835200, 
    1449838800, 1449842400, 1449846000, 1449849600, 1449853200, 1449856800, 
    1449860400, 1449864000, 1449867600, 1449871200, 1449874800, 1449878400, 
    1449882000, 1449885600, 1449889200, 1449892800, 1449896400, 1449900000, 
    1449903600, 1449907200, 1449910800, 1449914400, 1449918000, 1449921600, 
    1449925200, 1449928800, 1449932400, 1449936000, 1449939600, 1449943200, 
    1449946800, 1449950400, 1449954000, 1449957600, 1449961200, 1449964800, 
    1449968400, 1449972000, 1449975600, 1449979200, 1449982800, 1449986400, 
    1449990000, 1449993600, 1449997200, 1450000800, 1450004400, 1450008000, 
    1450011600, 1450015200, 1450018800, 1450022400, 1450026000, 1450029600, 
    1450033200, 1450036800, 1450040400, 1450044000, 1450047600, 1450051200, 
    1450054800, 1450058400, 1450062000, 1450065600, 1450069200, 1450072800, 
    1450076400, 1450080000, 1450083600, 1450087200, 1450090800, 1450094400, 
    1450098000, 1450101600, 1450105200, 1450108800, 1450112400, 1450116000, 
    1450119600, 1450123200, 1450126800, 1450130400, 1450134000, 1450137600, 
    1450141200, 1450144800, 1450148400, 1450152000, 1450155600, 1450159200, 
    1450162800, 1450166400, 1450170000, 1450173600, 1450177200, 1450180800, 
    1450184400, 1450188000, 1450191600, 1450195200, 1450198800, 1450202400, 
    1450206000, 1450209600, 1450213200, 1450216800, 1450220400, 1450224000, 
    1450227600, 1450231200, 1450234800, 1450238400, 1450242000, 1450245600, 
    1450249200, 1450252800, 1450256400, 1450260000, 1450263600, 1450267200, 
    1450270800, 1450274400, 1450278000, 1450281600, 1450285200, 1450288800, 
    1450292400, 1450296000, 1450299600, 1450303200, 1450306800, 1450310400, 
    1450314000, 1450317600, 1450321200, 1450324800, 1450328400, 1450332000, 
    1450335600, 1450339200, 1450342800, 1450346400, 1450350000, 1450353600, 
    1450357200, 1450360800, 1450364400, 1450368000, 1450371600, 1450375200, 
    1450378800, 1450382400, 1450386000, 1450389600, 1450393200, 1450396800, 
    1450400400, 1450404000, 1450407600, 1450411200, 1450414800, 1450418400, 
    1450422000, 1450425600, 1450429200, 1450432800, 1450436400, 1450440000, 
    1450443600, 1450447200, 1450450800, 1450454400, 1450458000, 1450461600, 
    1450465200, 1450468800, 1450472400, 1450476000, 1450479600, 1450483200, 
    1450486800, 1450490400, 1450494000, 1450497600, 1450501200, 1450504800, 
    1450508400, 1450512000, 1450515600, 1450519200, 1450522800, 1450526400, 
    1450530000, 1450533600, 1450537200, 1450540800, 1450544400, 1450548000, 
    1450551600, 1450555200, 1450558800, 1450562400, 1450566000, 1450569600, 
    1450573200, 1450576800, 1450580400, 1450584000, 1450587600, 1450591200, 
    1450594800, 1450598400, 1450602000, 1450605600, 1450609200, 1450612800, 
    1450616400, 1450620000, 1450623600, 1450627200, 1450630800, 1450634400, 
    1450638000, 1450641600, 1450645200, 1450648800, 1450652400, 1450656000, 
    1450659600, 1450663200, 1450666800, 1450670400, 1450674000, 1450677600, 
    1450681200, 1450684800, 1450688400, 1450692000, 1450695600, 1450699200, 
    1450702800, 1450706400, 1450710000, 1450713600, 1450717200, 1450720800, 
    1450724400, 1450728000, 1450731600, 1450735200, 1450738800, 1450742400, 
    1450746000, 1450749600, 1450753200, 1450756800, 1450760400, 1450764000, 
    1450767600, 1450771200, 1450774800, 1450778400, 1450782000, 1450785600, 
    1450789200, 1450792800, 1450796400, 1450800000, 1450803600, 1450807200, 
    1450810800, 1450814400, 1450818000, 1450821600, 1450825200, 1450828800, 
    1450832400, 1450836000, 1450839600, 1450843200, 1450846800, 1450850400, 
    1450854000, 1450857600, 1450861200, 1450864800, 1450868400, 1450872000, 
    1450875600, 1450879200, 1450882800, 1450886400, 1450890000, 1450893600, 
    1450897200, 1450900800, 1450904400, 1450908000, 1450911600, 1450915200, 
    1450918800, 1450922400, 1450926000, 1450929600, 1450933200, 1450936800, 
    1450940400, 1450944000, 1450947600, 1450951200, 1450954800, 1450958400, 
    1450962000, 1450965600, 1450969200, 1450972800, 1450976400, 1450980000, 
    1450983600, 1450987200, 1450990800, 1450994400, 1450998000, 1451001600, 
    1451005200, 1451008800, 1451012400, 1451016000, 1451019600, 1451023200, 
    1451026800, 1451030400, 1451034000, 1451037600, 1451041200, 1451044800, 
    1451048400, 1451052000, 1451055600, 1451059200, 1451062800, 1451066400, 
    1451070000, 1451073600, 1451077200, 1451080800, 1451084400, 1451088000, 
    1451091600, 1451095200, 1451098800, 1451102400, 1451106000, 1451109600, 
    1451113200, 1451116800, 1451120400, 1451124000, 1451127600, 1451131200, 
    1451134800, 1451138400, 1451142000, 1451145600, 1451149200, 1451152800, 
    1451156400, 1451160000, 1451163600, 1451167200, 1451170800, 1451174400, 
    1451178000, 1451181600, 1451185200, 1451188800, 1451192400, 1451196000, 
    1451199600, 1451203200, 1451206800, 1451210400, 1451214000, 1451217600, 
    1451221200, 1451224800, 1451228400, 1451232000, 1451235600, 1451239200, 
    1451242800, 1451246400, 1451250000, 1451253600, 1451257200, 1451260800, 
    1451264400, 1451268000, 1451271600, 1451275200, 1451278800, 1451282400, 
    1451286000, 1451289600, 1451293200, 1451296800, 1451300400, 1451304000, 
    1451307600, 1451311200, 1451314800, 1451318400, 1451322000, 1451325600, 
    1451329200, 1451332800, 1451336400, 1451340000, 1451343600, 1451347200, 
    1451350800, 1451354400, 1451358000, 1451361600, 1451365200, 1451368800, 
    1451372400, 1451376000, 1451379600, 1451383200, 1451386800, 1451390400, 
    1451394000, 1451397600, 1451401200, 1451404800, 1451408400, 1451412000, 
    1451415600, 1451419200, 1451422800, 1451426400, 1451430000, 1451433600, 
    1451437200, 1451440800, 1451444400, 1451448000, 1451451600, 1451455200, 
    1451458800, 1451462400, 1451466000, 1451469600, 1451473200, 1451476800, 
    1451480400, 1451484000, 1451487600, 1451491200, 1451494800, 1451498400, 
    1451502000, 1451505600, 1451509200, 1451512800, 1451516400, 1451520000, 
    1451523600, 1451527200, 1451530800, 1451534400, 1451538000, 1451541600, 
    1451545200, 1451548800, 1451552400, 1451556000, 1451559600, 1451563200, 
    1451566800, 1451570400, 1451574000, 1451577600, 1451581200, 1451584800, 
    1451588400, 1451592000, 1451595600, 1451599200, 1451602800, 1451606400, 
    1451610000, 1451613600, 1451617200, 1451620800, 1451624400, 1451628000, 
    1451631600, 1451635200, 1451638800, 1451642400, 1451646000, 1451649600, 
    1451653200, 1451656800, 1451660400, 1451664000, 1451667600, 1451671200, 
    1451674800, 1451678400, 1451682000, 1451685600, 1451689200, 1451692800, 
    1451696400, 1451700000, 1451703600, 1451707200, 1451710800, 1451714400, 
    1451718000, 1451721600, 1451725200, 1451728800, 1451732400, 1451736000, 
    1451739600, 1451743200, 1451746800, 1451750400, 1451754000, 1451757600, 
    1451761200, 1451764800, 1451768400, 1451772000, 1451775600, 1451779200, 
    1451782800, 1451786400, 1451790000, 1451793600, 1451797200, 1451800800, 
    1451804400, 1451808000, 1451811600, 1451815200, 1451818800, 1451822400, 
    1451826000, 1451829600, 1451833200, 1451836800, 1451840400, 1451844000, 
    1451847600, 1451851200, 1451854800, 1451858400, 1451862000, 1451865600, 
    1451869200, 1451872800, 1451876400, 1451880000, 1451883600, 1451887200, 
    1451890800, 1451894400, 1451898000, 1451901600, 1451905200, 1451908800, 
    1451912400, 1451916000, 1451919600, 1451923200, 1451926800, 1451930400, 
    1451934000, 1451937600, 1451941200, 1451944800, 1451948400, 1451952000, 
    1451955600, 1451959200, 1451962800, 1451966400, 1451970000, 1451973600, 
    1451977200, 1451980800, 1451984400, 1451988000, 1451991600, 1451995200, 
    1451998800, 1452002400, 1452006000, 1452009600, 1452013200, 1452016800, 
    1452020400, 1452024000, 1452027600, 1452031200, 1452034800, 1452038400, 
    1452042000, 1452045600, 1452049200, 1452052800, 1452056400, 1452060000, 
    1452063600, 1452067200, 1452070800, 1452074400, 1452078000, 1452081600, 
    1452085200, 1452088800, 1452092400, 1452096000, 1452099600, 1452103200, 
    1452106800, 1452110400, 1452114000, 1452117600, 1452121200, 1452124800, 
    1452128400, 1452132000, 1452135600, 1452139200, 1452142800, 1452146400, 
    1452150000, 1452153600, 1452157200, 1452160800, 1452164400, 1452168000, 
    1452171600, 1452175200, 1452178800, 1452182400, 1452186000, 1452189600, 
    1452193200, 1452196800, 1452200400, 1452204000, 1452207600, 1452211200, 
    1452214800, 1452218400, 1452222000, 1452225600, 1452229200, 1452232800, 
    1452236400, 1452240000, 1452243600, 1452247200, 1452250800, 1452254400, 
    1452258000, 1452261600, 1452265200, 1452268800, 1452272400, 1452276000, 
    1452279600, 1452283200, 1452286800, 1452290400, 1452294000, 1452297600, 
    1452301200, 1452304800, 1452308400, 1452312000, 1452315600, 1452319200, 
    1452322800, 1452326400, 1452330000, 1452333600, 1452337200, 1452340800, 
    1452344400, 1452348000, 1452351600, 1452355200, 1452358800, 1452362400, 
    1452366000, 1452369600, 1452373200, 1452376800, 1452380400, 1452384000, 
    1452387600, 1452391200, 1452394800, 1452398400, 1452402000, 1452405600, 
    1452409200, 1452412800, 1452416400, 1452420000, 1452423600, 1452427200, 
    1452430800, 1452434400, 1452438000, 1452441600, 1452445200, 1452448800, 
    1452452400, 1452456000, 1452459600, 1452463200, 1452466800, 1452470400, 
    1452474000, 1452477600, 1452481200, 1452484800, 1452488400, 1452492000, 
    1452495600, 1452499200, 1452502800, 1452506400, 1452510000, 1452513600, 
    1452517200, 1452520800, 1452524400, 1452528000, 1452531600, 1452535200, 
    1452538800, 1452542400, 1452546000, 1452549600, 1452553200, 1452556800, 
    1452560400, 1452564000, 1452567600, 1452571200, 1452574800, 1452578400, 
    1452582000, 1452585600, 1452589200, 1452592800, 1452596400, 1452600000, 
    1452603600, 1452607200, 1452610800, 1452614400, 1452618000, 1452621600, 
    1452625200, 1452628800, 1452632400, 1452636000, 1452639600, 1452643200, 
    1452646800, 1452650400, 1452654000, 1452657600, 1452661200, 1452664800, 
    1452668400, 1452672000, 1452675600, 1452679200, 1452682800, 1452686400, 
    1452690000, 1452693600, 1452697200, 1452700800, 1452704400, 1452708000, 
    1452711600, 1452715200, 1452718800, 1452722400, 1452726000, 1452729600, 
    1452733200, 1452736800, 1452740400, 1452744000, 1452747600, 1452751200, 
    1452754800, 1452758400, 1452762000, 1452765600, 1452769200, 1452772800, 
    1452776400, 1452780000, 1452783600, 1452787200, 1452790800, 1452794400, 
    1452798000, 1452801600, 1452805200, 1452808800, 1452812400, 1452816000, 
    1452819600, 1452823200, 1452826800, 1452830400, 1452834000, 1452837600, 
    1452841200, 1452844800, 1452848400, 1452852000, 1452855600, 1452859200, 
    1452862800, 1452866400, 1452870000, 1452873600, 1452877200, 1452880800, 
    1452884400, 1452888000, 1452891600, 1452895200, 1452898800, 1452902400, 
    1452906000, 1452909600, 1452913200, 1452916800, 1452920400, 1452924000, 
    1452927600, 1452931200, 1452934800, 1452938400, 1452942000, 1452945600, 
    1452949200, 1452952800, 1452956400, 1452960000, 1452963600, 1452967200, 
    1452970800, 1452974400, 1452978000, 1452981600, 1452985200, 1452988800, 
    1452992400, 1452996000, 1452999600, 1453003200, 1453006800, 1453010400, 
    1453014000, 1453017600, 1453021200, 1453024800, 1453028400, 1453032000, 
    1453035600, 1453039200, 1453042800, 1453046400, 1453050000, 1453053600, 
    1453057200, 1453060800, 1453064400, 1453068000, 1453071600, 1453075200, 
    1453078800, 1453082400, 1453086000, 1453089600, 1453093200, 1453096800, 
    1453100400, 1453104000, 1453107600, 1453111200, 1453114800, 1453118400, 
    1453122000, 1453125600, 1453129200, 1453132800, 1453136400, 1453140000, 
    1453143600, 1453147200, 1453150800, 1453154400, 1453158000, 1453161600, 
    1453165200, 1453168800, 1453172400, 1453176000, 1453179600, 1453183200, 
    1453186800, 1453190400, 1453194000, 1453197600, 1453201200, 1453204800, 
    1453208400, 1453212000, 1453215600, 1453219200, 1453222800, 1453226400, 
    1453230000, 1453233600, 1453237200, 1453240800, 1453244400, 1453248000, 
    1453251600, 1453255200, 1453258800, 1453262400, 1453266000, 1453269600, 
    1453273200, 1453276800, 1453280400, 1453284000, 1453287600, 1453291200, 
    1453294800, 1453298400, 1453302000, 1453305600, 1453309200, 1453312800, 
    1453316400, 1453320000, 1453323600, 1453327200, 1453330800, 1453334400, 
    1453338000, 1453341600, 1453345200, 1453348800, 1453352400, 1453356000, 
    1453359600, 1453363200, 1453366800, 1453370400, 1453374000, 1453377600, 
    1453381200, 1453384800, 1453388400, 1453392000, 1453395600, 1453399200, 
    1453402800, 1453406400, 1453410000, 1453413600, 1453417200, 1453420800, 
    1453424400, 1453428000, 1453431600, 1453435200, 1453438800, 1453442400, 
    1453446000, 1453449600, 1453453200, 1453456800, 1453460400, 1453464000, 
    1453467600, 1453471200, 1453474800, 1453478400, 1453482000, 1453485600, 
    1453489200, 1453492800, 1453496400, 1453500000, 1453503600, 1453507200, 
    1453510800, 1453514400, 1453518000, 1453521600, 1453525200, 1453528800, 
    1453532400, 1453536000, 1453539600, 1453543200, 1453546800, 1453550400, 
    1453554000, 1453557600, 1453561200, 1453564800, 1453568400, 1453572000, 
    1453575600, 1453579200, 1453582800, 1453586400, 1453590000, 1453593600, 
    1453597200, 1453600800, 1453604400, 1453608000, 1453611600, 1453615200, 
    1453618800, 1453622400, 1453626000, 1453629600, 1453633200, 1453636800, 
    1453640400, 1453644000, 1453647600, 1453651200, 1453654800, 1453658400, 
    1453662000, 1453665600, 1453669200, 1453672800, 1453676400, 1453680000, 
    1453683600, 1453687200, 1453690800, 1453694400, 1453698000, 1453701600, 
    1453705200, 1453708800, 1453712400, 1453716000, 1453719600, 1453723200, 
    1453726800, 1453730400, 1453734000, 1453737600, 1453741200, 1453744800, 
    1453748400, 1453752000, 1453755600, 1453759200, 1453762800, 1453766400, 
    1453770000, 1453773600, 1453777200, 1453780800, 1453784400, 1453788000, 
    1453791600, 1453795200, 1453798800, 1453802400, 1453806000, 1453809600, 
    1453813200, 1453816800, 1453820400, 1453824000, 1453827600, 1453831200, 
    1453834800, 1453838400, 1453842000, 1453845600, 1453849200, 1453852800, 
    1453856400, 1453860000, 1453863600, 1453867200, 1453870800, 1453874400, 
    1453878000, 1453881600, 1453885200, 1453888800, 1453892400, 1453896000, 
    1453899600, 1453903200, 1453906800, 1453910400, 1453914000, 1453917600, 
    1453921200, 1453924800, 1453928400, 1453932000, 1453935600, 1453939200, 
    1453942800, 1453946400, 1453950000, 1453953600, 1453957200, 1453960800, 
    1453964400, 1453968000, 1453971600, 1453975200, 1453978800, 1453982400, 
    1453986000, 1453989600, 1453993200, 1453996800, 1454000400, 1454004000, 
    1454007600, 1454011200, 1454014800, 1454018400, 1454022000, 1454025600, 
    1454029200, 1454032800, 1454036400, 1454040000, 1454043600, 1454047200, 
    1454050800, 1454054400, 1454058000, 1454061600, 1454065200, 1454068800, 
    1454072400, 1454076000, 1454079600, 1454083200, 1454086800, 1454090400, 
    1454094000, 1454097600, 1454101200, 1454104800, 1454108400, 1454112000, 
    1454115600, 1454119200, 1454122800, 1454126400, 1454130000, 1454133600, 
    1454137200, 1454140800, 1454144400, 1454148000, 1454151600, 1454155200, 
    1454158800, 1454162400, 1454166000, 1454169600, 1454173200, 1454176800, 
    1454180400, 1454184000, 1454187600, 1454191200, 1454194800, 1454198400, 
    1454202000, 1454205600, 1454209200, 1454212800, 1454216400, 1454220000, 
    1454223600, 1454227200, 1454230800, 1454234400, 1454238000, 1454241600, 
    1454245200, 1454248800, 1454252400, 1454256000, 1454259600, 1454263200, 
    1454266800, 1454270400, 1454274000, 1454277600, 1454281200, 1454284800, 
    1454288400, 1454292000, 1454295600, 1454299200, 1454302800, 1454306400, 
    1454310000, 1454313600, 1454317200, 1454320800, 1454324400, 1454328000, 
    1454331600, 1454335200, 1454338800, 1454342400, 1454346000, 1454349600, 
    1454353200, 1454356800, 1454360400, 1454364000, 1454367600, 1454371200, 
    1454374800, 1454378400, 1454382000, 1454385600, 1454389200, 1454392800, 
    1454396400, 1454400000, 1454403600, 1454407200, 1454410800, 1454414400, 
    1454418000, 1454421600, 1454425200, 1454428800, 1454432400, 1454436000, 
    1454439600, 1454443200, 1454446800, 1454450400, 1454454000, 1454457600, 
    1454461200, 1454464800, 1454468400, 1454472000, 1454475600, 1454479200, 
    1454482800, 1454486400, 1454490000, 1454493600, 1454497200, 1454500800, 
    1454504400, 1454508000, 1454511600, 1454515200, 1454518800, 1454522400, 
    1454526000, 1454529600, 1454533200, 1454536800, 1454540400, 1454544000, 
    1454547600, 1454551200, 1454554800, 1454558400, 1454562000, 1454565600, 
    1454569200, 1454572800, 1454576400, 1454580000, 1454583600, 1454587200, 
    1454590800, 1454594400, 1454598000, 1454601600, 1454605200, 1454608800, 
    1454612400, 1454616000, 1454619600, 1454623200, 1454626800, 1454630400, 
    1454634000, 1454637600, 1454641200, 1454644800, 1454648400, 1454652000, 
    1454655600, 1454659200, 1454662800, 1454666400, 1454670000, 1454673600, 
    1454677200, 1454680800, 1454684400, 1454688000, 1454691600, 1454695200, 
    1454698800, 1454702400, 1454706000, 1454709600, 1454713200, 1454716800, 
    1454720400, 1454724000, 1454727600, 1454731200, 1454734800, 1454738400, 
    1454742000, 1454745600, 1454749200, 1454752800, 1454756400, 1454760000, 
    1454763600, 1454767200, 1454770800, 1454774400, 1454778000, 1454781600, 
    1454785200, 1454788800, 1454792400, 1454796000, 1454799600, 1454803200, 
    1454806800, 1454810400, 1454814000, 1454817600, 1454821200, 1454824800, 
    1454828400, 1454832000, 1454835600, 1454839200, 1454842800, 1454846400, 
    1454850000, 1454853600, 1454857200, 1454860800, 1454864400, 1454868000, 
    1454871600, 1454875200, 1454878800, 1454882400, 1454886000, 1454889600, 
    1454893200, 1454896800, 1454900400, 1454904000, 1454907600, 1454911200, 
    1454914800, 1454918400, 1454922000, 1454925600, 1454929200, 1454932800, 
    1454936400, 1454940000, 1454943600, 1454947200, 1454950800, 1454954400, 
    1454958000, 1454961600, 1454965200, 1454968800, 1454972400, 1454976000, 
    1454979600, 1454983200, 1454986800, 1454990400, 1454994000, 1454997600, 
    1455001200, 1455004800, 1455008400, 1455012000, 1455015600, 1455019200, 
    1455022800, 1455026400, 1455030000, 1455033600, 1455037200, 1455040800, 
    1455044400, 1455048000, 1455051600, 1455055200, 1455058800, 1455062400, 
    1455066000, 1455069600, 1455073200, 1455076800, 1455080400, 1455084000, 
    1455087600, 1455091200, 1455094800, 1455098400, 1455102000, 1455105600, 
    1455109200, 1455112800, 1455116400, 1455120000, 1455123600, 1455127200, 
    1455130800, 1455134400, 1455138000, 1455141600, 1455145200, 1455148800, 
    1455152400, 1455156000, 1455159600, 1455163200, 1455166800, 1455170400, 
    1455174000, 1455177600, 1455181200, 1455184800, 1455188400, 1455192000, 
    1455195600, 1455199200, 1455202800, 1455206400, 1455210000, 1455213600, 
    1455217200, 1455220800, 1455224400, 1455228000, 1455231600, 1455235200, 
    1455238800, 1455242400, 1455246000, 1455249600, 1455253200, 1455256800, 
    1455260400, 1455264000, 1455267600, 1455271200, 1455274800, 1455278400, 
    1455282000, 1455285600, 1455289200, 1455292800, 1455296400, 1455300000, 
    1455303600, 1455307200, 1455310800, 1455314400, 1455318000, 1455321600, 
    1455325200, 1455328800, 1455332400, 1455336000, 1455339600, 1455343200, 
    1455346800, 1455350400, 1455354000, 1455357600, 1455361200, 1455364800, 
    1455368400, 1455372000, 1455375600, 1455379200, 1455382800, 1455386400, 
    1455390000, 1455393600, 1455397200, 1455400800, 1455404400, 1455408000, 
    1455411600, 1455415200, 1455418800, 1455422400, 1455426000, 1455429600, 
    1455433200, 1455436800, 1455440400, 1455444000, 1455447600, 1455451200, 
    1455454800, 1455458400, 1455462000, 1455465600, 1455469200, 1455472800, 
    1455476400, 1455480000, 1455483600, 1455487200, 1455490800, 1455494400, 
    1455498000, 1455501600, 1455505200, 1455508800, 1455512400, 1455516000, 
    1455519600, 1455523200, 1455526800, 1455530400, 1455534000, 1455537600, 
    1455541200, 1455544800, 1455548400, 1455552000, 1455555600, 1455559200, 
    1455562800, 1455566400, 1455570000, 1455573600, 1455577200, 1455580800, 
    1455584400, 1455588000, 1455591600, 1455595200, 1455598800, 1455602400, 
    1455606000, 1455609600, 1455613200, 1455616800, 1455620400, 1455624000, 
    1455627600, 1455631200, 1455634800, 1455638400, 1455642000, 1455645600, 
    1455649200, 1455652800, 1455656400, 1455660000, 1455663600, 1455667200, 
    1455670800, 1455674400, 1455678000, 1455681600, 1455685200, 1455688800, 
    1455692400, 1455696000, 1455699600, 1455703200, 1455706800, 1455710400, 
    1455714000, 1455717600, 1455721200, 1455724800, 1455728400, 1455732000, 
    1455735600, 1455739200, 1455742800, 1455746400, 1455750000, 1455753600, 
    1455757200, 1455760800, 1455764400, 1455768000, 1455771600, 1455775200, 
    1455778800, 1455782400, 1455786000, 1455789600, 1455793200, 1455796800, 
    1455800400, 1455804000, 1455807600, 1455811200, 1455814800, 1455818400, 
    1455822000, 1455825600, 1455829200, 1455832800, 1455836400, 1455840000, 
    1455843600, 1455847200, 1455850800, 1455854400, 1455858000, 1455861600, 
    1455865200, 1455868800, 1455872400, 1455876000, 1455879600, 1455883200, 
    1455886800, 1455890400, 1455894000, 1455897600, 1455901200, 1455904800, 
    1455908400, 1455912000, 1455915600, 1455919200, 1455922800, 1455926400, 
    1455930000, 1455933600, 1455937200, 1455940800, 1455944400, 1455948000, 
    1455951600, 1455955200, 1455958800, 1455962400, 1455966000, 1455969600, 
    1455973200, 1455976800, 1455980400, 1455984000, 1455987600, 1455991200, 
    1455994800, 1455998400, 1456002000, 1456005600, 1456009200, 1456012800, 
    1456016400, 1456020000, 1456023600, 1456027200, 1456030800, 1456034400, 
    1456038000, 1456041600, 1456045200, 1456048800, 1456052400, 1456056000, 
    1456059600, 1456063200, 1456066800, 1456070400, 1456074000, 1456077600, 
    1456081200, 1456084800, 1456088400, 1456092000, 1456095600, 1456099200, 
    1456102800, 1456106400, 1456110000, 1456113600, 1456117200, 1456120800, 
    1456124400, 1456128000, 1456131600, 1456135200, 1456138800, 1456142400, 
    1456146000, 1456149600, 1456153200, 1456156800, 1456160400, 1456164000, 
    1456167600, 1456171200, 1456174800, 1456178400, 1456182000, 1456185600, 
    1456189200, 1456192800, 1456196400, 1456200000, 1456203600, 1456207200, 
    1456210800, 1456214400, 1456218000, 1456221600, 1456225200, 1456228800, 
    1456232400, 1456236000, 1456239600, 1456243200, 1456246800, 1456250400, 
    1456254000, 1456257600, 1456261200, 1456264800, 1456268400, 1456272000, 
    1456275600, 1456279200, 1456282800, 1456286400, 1456290000, 1456293600, 
    1456297200, 1456300800, 1456304400, 1456308000, 1456311600, 1456315200, 
    1456318800, 1456322400, 1456326000, 1456329600, 1456333200, 1456336800, 
    1456340400, 1456344000, 1456347600, 1456351200, 1456354800, 1456358400, 
    1456362000, 1456365600, 1456369200, 1456372800, 1456376400, 1456380000, 
    1456383600, 1456387200, 1456390800, 1456394400, 1456398000, 1456401600, 
    1456405200, 1456408800, 1456412400, 1456416000, 1456419600, 1456423200, 
    1456426800, 1456430400, 1456434000, 1456437600, 1456441200, 1456444800, 
    1456448400, 1456452000, 1456455600, 1456459200, 1456462800, 1456466400, 
    1456470000, 1456473600, 1456477200, 1456480800, 1456484400, 1456488000, 
    1456491600, 1456495200, 1456498800, 1456502400, 1456506000, 1456509600, 
    1456513200, 1456516800, 1456520400, 1456524000, 1456527600, 1456531200, 
    1456534800, 1456538400, 1456542000, 1456545600, 1456549200, 1456552800, 
    1456556400, 1456560000, 1456563600, 1456567200, 1456570800, 1456574400, 
    1456578000, 1456581600, 1456585200, 1456588800, 1456592400, 1456596000, 
    1456599600, 1456603200, 1456606800, 1456610400, 1456614000, 1456617600, 
    1456621200, 1456624800, 1456628400, 1456632000, 1456635600, 1456639200, 
    1456642800, 1456646400, 1456650000, 1456653600, 1456657200, 1456660800, 
    1456664400, 1456668000, 1456671600, 1456675200, 1456678800, 1456682400, 
    1456686000, 1456689600, 1456693200, 1456696800, 1456700400, 1456704000, 
    1456707600, 1456711200, 1456714800, 1456718400, 1456722000, 1456725600, 
    1456729200, 1456732800, 1456736400, 1456740000, 1456743600, 1456747200, 
    1456750800, 1456754400, 1456758000, 1456761600, 1456765200, 1456768800, 
    1456772400, 1456776000, 1456779600, 1456783200, 1456786800, 1456790400, 
    1456794000, 1456797600, 1456801200, 1456804800, 1456808400, 1456812000, 
    1456815600, 1456819200, 1456822800, 1456826400, 1456830000, 1456833600, 
    1456837200, 1456840800, 1456844400, 1456848000, 1456851600, 1456855200, 
    1456858800, 1456862400, 1456866000, 1456869600, 1456873200, 1456876800, 
    1456880400, 1456884000, 1456887600, 1456891200, 1456894800, 1456898400, 
    1456902000, 1456905600, 1456909200, 1456912800, 1456916400, 1456920000, 
    1456923600, 1456927200, 1456930800, 1456934400, 1456938000, 1456941600, 
    1456945200, 1456948800, 1456952400, 1456956000, 1456959600, 1456963200, 
    1456966800, 1456970400, 1456974000, 1456977600, 1456981200, 1456984800, 
    1456988400, 1456992000, 1456995600, 1456999200, 1457002800, 1457006400, 
    1457010000, 1457013600, 1457017200, 1457020800, 1457024400, 1457028000, 
    1457031600, 1457035200, 1457038800, 1457042400, 1457046000, 1457049600, 
    1457053200, 1457056800, 1457060400, 1457064000, 1457067600, 1457071200, 
    1457074800, 1457078400, 1457082000, 1457085600, 1457089200, 1457092800, 
    1457096400, 1457100000, 1457103600, 1457107200, 1457110800, 1457114400, 
    1457118000, 1457121600, 1457125200, 1457128800, 1457132400, 1457136000, 
    1457139600, 1457143200, 1457146800, 1457150400, 1457154000, 1457157600, 
    1457161200, 1457164800, 1457168400, 1457172000, 1457175600, 1457179200, 
    1457182800, 1457186400, 1457190000, 1457193600, 1457197200, 1457200800, 
    1457204400, 1457208000, 1457211600, 1457215200, 1457218800, 1457222400, 
    1457226000, 1457229600, 1457233200, 1457236800, 1457240400, 1457244000, 
    1457247600, 1457251200, 1457254800, 1457258400, 1457262000, 1457265600, 
    1457269200, 1457272800, 1457276400, 1457280000, 1457283600, 1457287200, 
    1457290800, 1457294400, 1457298000, 1457301600, 1457305200, 1457308800, 
    1457312400, 1457316000, 1457319600, 1457323200, 1457326800, 1457330400, 
    1457334000, 1457337600, 1457341200, 1457344800, 1457348400, 1457352000, 
    1457355600, 1457359200, 1457362800, 1457366400, 1457370000, 1457373600, 
    1457377200, 1457380800, 1457384400, 1457388000, 1457391600, 1457395200, 
    1457398800, 1457402400, 1457406000, 1457409600, 1457413200, 1457416800, 
    1457420400, 1457424000, 1457427600, 1457431200, 1457434800, 1457438400, 
    1457442000, 1457445600, 1457449200, 1457452800, 1457456400, 1457460000, 
    1457463600, 1457467200, 1457470800, 1457474400, 1457478000, 1457481600, 
    1457485200, 1457488800, 1457492400, 1457496000, 1457499600, 1457503200, 
    1457506800, 1457510400, 1457514000, 1457517600, 1457521200, 1457524800, 
    1457528400, 1457532000, 1457535600, 1457539200, 1457542800, 1457546400, 
    1457550000, 1457553600, 1457557200, 1457560800, 1457564400, 1457568000, 
    1457571600, 1457575200, 1457578800, 1457582400, 1457586000, 1457589600, 
    1457593200, 1457596800, 1457600400, 1457604000, 1457607600, 1457611200, 
    1457614800, 1457618400, 1457622000, 1457625600, 1457629200, 1457632800, 
    1457636400, 1457640000, 1457643600, 1457647200, 1457650800, 1457654400, 
    1457658000, 1457661600, 1457665200, 1457668800, 1457672400, 1457676000, 
    1457679600, 1457683200, 1457686800, 1457690400, 1457694000, 1457697600, 
    1457701200, 1457704800, 1457708400, 1457712000, 1457715600, 1457719200, 
    1457722800, 1457726400, 1457730000, 1457733600, 1457737200, 1457740800, 
    1457744400, 1457748000, 1457751600, 1457755200, 1457758800, 1457762400, 
    1457766000, 1457769600, 1457773200, 1457776800, 1457780400, 1457784000, 
    1457787600, 1457791200, 1457794800, 1457798400, 1457802000, 1457805600, 
    1457809200, 1457812800, 1457816400, 1457820000, 1457823600, 1457827200, 
    1457830800, 1457834400, 1457838000, 1457841600, 1457845200, 1457848800, 
    1457852400, 1457856000, 1457859600, 1457863200, 1457866800, 1457870400, 
    1457874000, 1457877600, 1457881200, 1457884800, 1457888400, 1457892000, 
    1457895600, 1457899200, 1457902800, 1457906400, 1457910000, 1457913600, 
    1457917200, 1457920800, 1457924400, 1457928000, 1457931600, 1457935200, 
    1457938800, 1457942400, 1457946000, 1457949600, 1457953200, 1457956800, 
    1457960400, 1457964000, 1457967600, 1457971200, 1457974800, 1457978400, 
    1457982000, 1457985600, 1457989200, 1457992800, 1457996400, 1458000000, 
    1458003600, 1458007200, 1458010800, 1458014400, 1458018000, 1458021600, 
    1458025200, 1458028800, 1458032400, 1458036000, 1458039600, 1458043200, 
    1458046800, 1458050400, 1458054000, 1458057600, 1458061200, 1458064800, 
    1458068400, 1458072000, 1458075600, 1458079200, 1458082800, 1458086400, 
    1458090000, 1458093600, 1458097200, 1458100800, 1458104400, 1458108000, 
    1458111600, 1458115200, 1458118800, 1458122400, 1458126000, 1458129600, 
    1458133200, 1458136800, 1458140400, 1458144000, 1458147600, 1458151200, 
    1458154800, 1458158400, 1458162000, 1458165600, 1458169200, 1458172800, 
    1458176400, 1458180000, 1458183600, 1458187200, 1458190800, 1458194400, 
    1458198000, 1458201600, 1458205200, 1458208800, 1458212400, 1458216000, 
    1458219600, 1458223200, 1458226800, 1458230400, 1458234000, 1458237600, 
    1458241200, 1458244800, 1458248400, 1458252000, 1458255600, 1458259200, 
    1458262800, 1458266400, 1458270000, 1458273600, 1458277200, 1458280800, 
    1458284400, 1458288000, 1458291600, 1458295200, 1458298800, 1458302400, 
    1458306000, 1458309600, 1458313200, 1458316800, 1458320400, 1458324000, 
    1458327600, 1458331200, 1458334800, 1458338400, 1458342000, 1458345600, 
    1458349200, 1458352800, 1458356400, 1458360000, 1458363600, 1458367200, 
    1458370800, 1458374400, 1458378000, 1458381600, 1458385200, 1458388800, 
    1458392400, 1458396000, 1458399600, 1458403200, 1458406800, 1458410400, 
    1458414000, 1458417600, 1458421200, 1458424800, 1458428400, 1458432000, 
    1458435600, 1458439200, 1458442800, 1458446400, 1458450000, 1458453600, 
    1458457200, 1458460800, 1458464400, 1458468000, 1458471600, 1458475200, 
    1458478800, 1458482400, 1458486000, 1458489600, 1458493200, 1458496800, 
    1458500400, 1458504000, 1458507600, 1458511200, 1458514800, 1458518400, 
    1458522000, 1458525600, 1458529200, 1458532800, 1458536400, 1458540000, 
    1458543600, 1458547200, 1458550800, 1458554400, 1458558000, 1458561600, 
    1458565200, 1458568800, 1458572400, 1458576000, 1458579600, 1458583200, 
    1458586800, 1458590400, 1458594000, 1458597600, 1458601200, 1458604800, 
    1458608400, 1458612000, 1458615600, 1458619200, 1458622800, 1458626400, 
    1458630000, 1458633600, 1458637200, 1458640800, 1458644400, 1458648000, 
    1458651600, 1458655200, 1458658800, 1458662400, 1458666000, 1458669600, 
    1458673200, 1458676800, 1458680400, 1458684000, 1458687600, 1458691200, 
    1458694800, 1458698400, 1458702000, 1458705600, 1458709200, 1458712800, 
    1458716400, 1458720000, 1458723600, 1458727200, 1458730800, 1458734400, 
    1458738000, 1458741600, 1458745200, 1458748800, 1458752400, 1458756000, 
    1458759600, 1458763200, 1458766800, 1458770400, 1458774000, 1458777600, 
    1458781200, 1458784800, 1458788400, 1458792000, 1458795600, 1458799200, 
    1458802800, 1458806400, 1458810000, 1458813600, 1458817200, 1458820800, 
    1458824400, 1458828000, 1458831600, 1458835200, 1458838800, 1458842400, 
    1458846000, 1458849600, 1458853200, 1458856800, 1458860400, 1458864000, 
    1458867600, 1458871200, 1458874800, 1458878400, 1458882000, 1458885600, 
    1458889200, 1458892800, 1458896400, 1458900000, 1458903600, 1458907200, 
    1458910800, 1458914400, 1458918000, 1458921600, 1458925200, 1458928800, 
    1458932400, 1458936000, 1458939600, 1458943200, 1458946800, 1458950400, 
    1458954000, 1458957600, 1458961200, 1458964800, 1458968400, 1458972000, 
    1458975600, 1458979200, 1458982800, 1458986400, 1458990000, 1458993600, 
    1458997200, 1459000800, 1459004400, 1459008000, 1459011600, 1459015200, 
    1459018800, 1459022400, 1459026000, 1459029600, 1459033200, 1459036800, 
    1459040400, 1459044000, 1459047600, 1459051200, 1459054800, 1459058400, 
    1459062000, 1459065600, 1459069200, 1459072800, 1459076400, 1459080000, 
    1459083600, 1459087200, 1459090800, 1459094400, 1459098000, 1459101600, 
    1459105200, 1459108800, 1459112400, 1459116000, 1459119600, 1459123200, 
    1459126800, 1459130400, 1459134000, 1459137600, 1459141200, 1459144800, 
    1459148400, 1459152000, 1459155600, 1459159200, 1459162800, 1459166400, 
    1459170000, 1459173600, 1459177200, 1459180800, 1459184400, 1459188000, 
    1459191600, 1459195200, 1459198800, 1459202400, 1459206000, 1459209600, 
    1459213200, 1459216800, 1459220400, 1459224000, 1459227600, 1459231200, 
    1459234800, 1459238400, 1459242000, 1459245600, 1459249200, 1459252800, 
    1459256400, 1459260000, 1459263600, 1459267200, 1459270800, 1459274400, 
    1459278000, 1459281600, 1459285200, 1459288800, 1459292400, 1459296000, 
    1459299600, 1459303200, 1459306800, 1459310400, 1459314000, 1459317600, 
    1459321200, 1459324800, 1459328400, 1459332000, 1459335600, 1459339200, 
    1459342800, 1459346400, 1459350000, 1459353600, 1459357200, 1459360800, 
    1459364400, 1459368000, 1459371600, 1459375200, 1459378800, 1459382400, 
    1459386000, 1459389600, 1459393200, 1459396800, 1459400400, 1459404000, 
    1459407600, 1459411200, 1459414800, 1459418400, 1459422000, 1459425600, 
    1459429200, 1459432800, 1459436400, 1459440000, 1459443600, 1459447200, 
    1459450800, 1459454400, 1459458000, 1459461600, 1459465200, 1459468800, 
    1459472400, 1459476000, 1459479600, 1459483200, 1459486800, 1459490400, 
    1459494000, 1459497600, 1459501200, 1459504800, 1459508400, 1459512000, 
    1459515600, 1459519200, 1459522800, 1459526400, 1459530000, 1459533600, 
    1459537200, 1459540800, 1459544400, 1459548000, 1459551600, 1459555200, 
    1459558800, 1459562400, 1459566000, 1459569600, 1459573200, 1459576800, 
    1459580400, 1459584000, 1459587600, 1459591200, 1459594800, 1459598400, 
    1459602000, 1459605600, 1459609200, 1459612800, 1459616400, 1459620000, 
    1459623600, 1459627200, 1459630800, 1459634400, 1459638000, 1459641600, 
    1459645200, 1459648800, 1459652400, 1459656000, 1459659600, 1459663200, 
    1459666800, 1459670400, 1459674000, 1459677600, 1459681200, 1459684800, 
    1459688400, 1459692000, 1459695600, 1459699200, 1459702800, 1459706400, 
    1459710000, 1459713600, 1459717200, 1459720800, 1459724400, 1459728000, 
    1459731600, 1459735200, 1459738800, 1459742400, 1459746000, 1459749600, 
    1459753200, 1459756800, 1459760400, 1459764000, 1459767600, 1459771200, 
    1459774800, 1459778400, 1459782000, 1459785600, 1459789200, 1459792800, 
    1459796400, 1459800000, 1459803600, 1459807200, 1459810800, 1459814400, 
    1459818000, 1459821600, 1459825200, 1459828800, 1459832400, 1459836000, 
    1459839600, 1459843200, 1459846800, 1459850400, 1459854000, 1459857600, 
    1459861200, 1459864800, 1459868400, 1459872000, 1459875600, 1459879200, 
    1459882800, 1459886400, 1459890000, 1459893600, 1459897200, 1459900800, 
    1459904400, 1459908000, 1459911600, 1459915200, 1459918800, 1459922400, 
    1459926000, 1459929600, 1459933200, 1459936800, 1459940400, 1459944000, 
    1459947600, 1459951200, 1459954800, 1459958400, 1459962000, 1459965600, 
    1459969200, 1459972800, 1459976400, 1459980000, 1459983600, 1459987200, 
    1459990800, 1459994400, 1459998000, 1460001600, 1460005200, 1460008800, 
    1460012400, 1460016000, 1460019600, 1460023200, 1460026800, 1460030400, 
    1460034000, 1460037600, 1460041200, 1460044800, 1460048400, 1460052000, 
    1460055600, 1460059200, 1460062800, 1460066400, 1460070000, 1460073600, 
    1460077200, 1460080800, 1460084400, 1460088000, 1460091600, 1460095200, 
    1460098800, 1460102400, 1460106000, 1460109600, 1460113200, 1460116800, 
    1460120400, 1460124000, 1460127600, 1460131200, 1460134800, 1460138400, 
    1460142000, 1460145600, 1460149200, 1460152800, 1460156400, 1460160000, 
    1460163600, 1460167200, 1460170800, 1460174400, 1460178000, 1460181600, 
    1460185200, 1460188800, 1460192400, 1460196000, 1460199600, 1460203200, 
    1460206800, 1460210400, 1460214000, 1460217600, 1460221200, 1460224800, 
    1460228400, 1460232000, 1460235600, 1460239200, 1460242800, 1460246400, 
    1460250000, 1460253600, 1460257200, 1460260800, 1460264400, 1460268000, 
    1460271600, 1460275200, 1460278800, 1460282400, 1460286000, 1460289600, 
    1460293200, 1460296800, 1460300400, 1460304000, 1460307600, 1460311200, 
    1460314800, 1460318400, 1460322000, 1460325600, 1460329200, 1460332800, 
    1460336400, 1460340000, 1460343600, 1460347200, 1460350800, 1460354400, 
    1460358000, 1460361600, 1460365200, 1460368800, 1460372400, 1460376000, 
    1460379600, 1460383200, 1460386800, 1460390400, 1460394000, 1460397600, 
    1460401200, 1460404800, 1460408400, 1460412000, 1460415600, 1460419200, 
    1460422800, 1460426400, 1460430000, 1460433600, 1460437200, 1460440800, 
    1460444400, 1460448000, 1460451600, 1460455200, 1460458800, 1460462400, 
    1460466000, 1460469600, 1460473200, 1460476800, 1460480400, 1460484000, 
    1460487600, 1460491200, 1460494800, 1460498400, 1460502000, 1460505600, 
    1460509200, 1460512800, 1460516400, 1460520000, 1460523600, 1460527200, 
    1460530800, 1460534400, 1460538000, 1460541600, 1460545200, 1460548800, 
    1460552400, 1460556000, 1460559600, 1460563200, 1460566800, 1460570400, 
    1460574000, 1460577600, 1460581200, 1460584800, 1460588400, 1460592000, 
    1460595600, 1460599200, 1460602800, 1460606400, 1460610000, 1460613600, 
    1460617200, 1460620800, 1460624400, 1460628000, 1460631600, 1460635200, 
    1460638800, 1460642400, 1460646000, 1460649600, 1460653200, 1460656800, 
    1460660400, 1460664000, 1460667600, 1460671200, 1460674800, 1460678400, 
    1460682000, 1460685600, 1460689200, 1460692800, 1460696400, 1460700000, 
    1460703600, 1460707200, 1460710800, 1460714400, 1460718000, 1460721600, 
    1460725200, 1460728800, 1460732400, 1460736000, 1460739600, 1460743200, 
    1460746800, 1460750400, 1460754000, 1460757600, 1460761200, 1460764800, 
    1460768400, 1460772000, 1460775600, 1460779200, 1460782800, 1460786400, 
    1460790000, 1460793600, 1460797200, 1460800800, 1460804400, 1460808000, 
    1460811600, 1460815200, 1460818800, 1460822400, 1460826000, 1460829600, 
    1460833200, 1460836800, 1460840400, 1460844000, 1460847600, 1460851200, 
    1460854800, 1460858400, 1460862000, 1460865600, 1460869200, 1460872800, 
    1460876400, 1460880000, 1460883600, 1460887200, 1460890800, 1460894400, 
    1460898000, 1460901600, 1460905200, 1460908800, 1460912400, 1460916000, 
    1460919600, 1460923200, 1460926800, 1460930400, 1460934000, 1460937600, 
    1460941200, 1460944800, 1460948400, 1460952000, 1460955600, 1460959200, 
    1460962800, 1460966400, 1460970000, 1460973600, 1460977200, 1460980800, 
    1460984400, 1460988000, 1460991600, 1460995200, 1460998800, 1461002400, 
    1461006000, 1461009600, 1461013200, 1461016800, 1461020400, 1461024000, 
    1461027600, 1461031200, 1461034800, 1461038400, 1461042000, 1461045600, 
    1461049200, 1461052800, 1461056400, 1461060000, 1461063600, 1461067200, 
    1461070800, 1461074400, 1461078000, 1461081600, 1461085200, 1461088800, 
    1461092400, 1461096000, 1461099600, 1461103200, 1461106800, 1461110400, 
    1461114000, 1461117600, 1461121200, 1461124800, 1461128400, 1461132000, 
    1461135600, 1461139200, 1461142800, 1461146400, 1461150000, 1461153600, 
    1461157200, 1461160800, 1461164400, 1461168000, 1461171600, 1461175200, 
    1461178800, 1461182400, 1461186000, 1461189600, 1461193200, 1461196800, 
    1461200400, 1461204000, 1461207600, 1461211200, 1461214800, 1461218400, 
    1461222000, 1461225600, 1461229200, 1461232800, 1461236400, 1461240000, 
    1461243600, 1461247200, 1461250800, 1461254400, 1461258000, 1461261600, 
    1461265200, 1461268800, 1461272400, 1461276000, 1461279600, 1461283200, 
    1461286800, 1461290400, 1461294000, 1461297600, 1461301200, 1461304800, 
    1461308400, 1461312000, 1461315600, 1461319200, 1461322800, 1461326400, 
    1461330000, 1461333600, 1461337200, 1461340800, 1461344400, 1461348000, 
    1461351600, 1461355200, 1461358800, 1461362400, 1461366000, 1461369600, 
    1461373200, 1461376800, 1461380400, 1461384000, 1461387600, 1461391200, 
    1461394800, 1461398400, 1461402000, 1461405600, 1461409200, 1461412800, 
    1461416400, 1461420000, 1461423600, 1461427200, 1461430800, 1461434400, 
    1461438000, 1461441600, 1461445200, 1461448800, 1461452400, 1461456000, 
    1461459600, 1461463200, 1461466800, 1461470400, 1461474000, 1461477600, 
    1461481200, 1461484800, 1461488400, 1461492000, 1461495600, 1461499200, 
    1461502800, 1461506400, 1461510000, 1461513600, 1461517200, 1461520800, 
    1461524400, 1461528000, 1461531600, 1461535200, 1461538800, 1461542400, 
    1461546000, 1461549600, 1461553200, 1461556800, 1461560400, 1461564000, 
    1461567600, 1461571200, 1461574800, 1461578400, 1461582000, 1461585600, 
    1461589200, 1461592800, 1461596400, 1461600000, 1461603600, 1461607200, 
    1461610800, 1461614400, 1461618000, 1461621600, 1461625200, 1461628800, 
    1461632400, 1461636000, 1461639600, 1461643200, 1461646800, 1461650400, 
    1461654000, 1461657600, 1461661200, 1461664800, 1461668400, 1461672000, 
    1461675600, 1461679200, 1461682800, 1461686400, 1461690000, 1461693600, 
    1461697200, 1461700800, 1461704400, 1461708000, 1461711600, 1461715200, 
    1461718800, 1461722400, 1461726000, 1461729600, 1461733200, 1461736800, 
    1461740400, 1461744000, 1461747600, 1461751200, 1461754800, 1461758400, 
    1461762000, 1461765600, 1461769200, 1461772800, 1461776400, 1461780000, 
    1461783600, 1461787200, 1461790800, 1461794400, 1461798000, 1461801600, 
    1461805200, 1461808800, 1461812400, 1461816000, 1461819600, 1461823200, 
    1461826800, 1461830400, 1461834000, 1461837600, 1461841200, 1461844800, 
    1461848400, 1461852000, 1461855600, 1461859200, 1461862800, 1461866400, 
    1461870000, 1461873600, 1461877200, 1461880800, 1461884400, 1461888000, 
    1461891600, 1461895200, 1461898800, 1461902400, 1461906000, 1461909600, 
    1461913200, 1461916800, 1461920400, 1461924000, 1461927600, 1461931200, 
    1461934800, 1461938400, 1461942000, 1461945600, 1461949200, 1461952800, 
    1461956400, 1461960000, 1461963600, 1461967200, 1461970800, 1461974400, 
    1461978000, 1461981600, 1461985200, 1461988800, 1461992400, 1461996000, 
    1461999600, 1462003200, 1462006800, 1462010400, 1462014000, 1462017600, 
    1462021200, 1462024800, 1462028400, 1462032000, 1462035600, 1462039200, 
    1462042800, 1462046400, 1462050000, 1462053600, 1462057200, 1462060800, 
    1462064400, 1462068000, 1462071600, 1462075200, 1462078800, 1462082400, 
    1462086000, 1462089600, 1462093200, 1462096800, 1462100400, 1462104000, 
    1462107600, 1462111200, 1462114800, 1462118400, 1462122000, 1462125600, 
    1462129200, 1462132800, 1462136400, 1462140000, 1462143600, 1462147200, 
    1462150800, 1462154400, 1462158000, 1462161600, 1462165200, 1462168800, 
    1462172400, 1462176000, 1462179600, 1462183200, 1462186800, 1462190400, 
    1462194000, 1462197600, 1462201200, 1462204800, 1462208400, 1462212000, 
    1462215600, 1462219200, 1462222800, 1462226400, 1462230000, 1462233600, 
    1462237200, 1462240800, 1462244400, 1462248000, 1462251600, 1462255200, 
    1462258800, 1462262400, 1462266000, 1462269600, 1462273200, 1462276800, 
    1462280400, 1462284000, 1462287600, 1462291200, 1462294800, 1462298400, 
    1462302000, 1462305600, 1462309200, 1462312800, 1462316400, 1462320000, 
    1462323600, 1462327200, 1462330800, 1462334400, 1462338000, 1462341600, 
    1462345200, 1462348800, 1462352400, 1462356000, 1462359600, 1462363200, 
    1462366800, 1462370400, 1462374000, 1462377600, 1462381200, 1462384800, 
    1462388400, 1462392000, 1462395600, 1462399200, 1462402800, 1462406400, 
    1462410000, 1462413600, 1462417200, 1462420800, 1462424400, 1462428000, 
    1462431600, 1462435200, 1462438800, 1462442400, 1462446000, 1462449600, 
    1462453200, 1462456800, 1462460400, 1462464000, 1462467600, 1462471200, 
    1462474800, 1462478400, 1462482000, 1462485600, 1462489200, 1462492800, 
    1462496400, 1462500000, 1462503600, 1462507200, 1462510800, 1462514400, 
    1462518000, 1462521600, 1462525200, 1462528800, 1462532400, 1462536000, 
    1462539600, 1462543200, 1462546800, 1462550400, 1462554000, 1462557600, 
    1462561200, 1462564800, 1462568400, 1462572000, 1462575600, 1462579200, 
    1462582800, 1462586400, 1462590000, 1462593600, 1462597200, 1462600800, 
    1462604400, 1462608000, 1462611600, 1462615200, 1462618800, 1462622400, 
    1462626000, 1462629600, 1462633200, 1462636800, 1462640400, 1462644000, 
    1462647600, 1462651200, 1462654800, 1462658400, 1462662000, 1462665600, 
    1462669200, 1462672800, 1462676400, 1462680000, 1462683600, 1462687200, 
    1462690800, 1462694400, 1462698000, 1462701600, 1462705200, 1462708800, 
    1462712400, 1462716000, 1462719600, 1462723200, 1462726800, 1462730400, 
    1462734000, 1462737600, 1462741200, 1462744800, 1462748400, 1462752000, 
    1462755600, 1462759200, 1462762800, 1462766400, 1462770000, 1462773600, 
    1462777200, 1462780800, 1462784400, 1462788000, 1462791600, 1462795200, 
    1462798800, 1462802400, 1462806000, 1462809600, 1462813200, 1462816800, 
    1462820400, 1462824000, 1462827600, 1462831200, 1462834800, 1462838400, 
    1462842000, 1462845600, 1462849200, 1462852800, 1462856400, 1462860000, 
    1462863600, 1462867200, 1462870800, 1462874400, 1462878000, 1462881600, 
    1462885200, 1462888800, 1462892400, 1462896000, 1462899600, 1462903200, 
    1462906800, 1462910400, 1462914000, 1462917600, 1462921200, 1462924800, 
    1462928400, 1462932000, 1462935600, 1462939200, 1462942800, 1462946400, 
    1462950000, 1462953600, 1462957200, 1462960800, 1462964400, 1462968000, 
    1462971600, 1462975200, 1462978800, 1462982400, 1462986000, 1462989600, 
    1462993200, 1462996800, 1463000400, 1463004000, 1463007600, 1463011200, 
    1463014800, 1463018400, 1463022000, 1463025600, 1463029200, 1463032800, 
    1463036400, 1463040000, 1463043600, 1463047200, 1463050800, 1463054400, 
    1463058000, 1463061600, 1463065200, 1463068800, 1463072400, 1463076000, 
    1463079600, 1463083200, 1463086800, 1463090400, 1463094000, 1463097600, 
    1463101200, 1463104800, 1463108400, 1463112000, 1463115600, 1463119200, 
    1463122800, 1463126400, 1463130000, 1463133600, 1463137200, 1463140800, 
    1463144400, 1463148000, 1463151600, 1463155200, 1463158800, 1463162400, 
    1463166000, 1463169600, 1463173200, 1463176800, 1463180400, 1463184000, 
    1463187600, 1463191200, 1463194800, 1463198400, 1463202000, 1463205600, 
    1463209200, 1463212800, 1463216400, 1463220000, 1463223600, 1463227200, 
    1463230800, 1463234400, 1463238000, 1463241600, 1463245200, 1463248800, 
    1463252400, 1463256000, 1463259600, 1463263200, 1463266800, 1463270400, 
    1463274000, 1463277600, 1463281200, 1463284800, 1463288400, 1463292000, 
    1463295600, 1463299200, 1463302800, 1463306400, 1463310000, 1463313600, 
    1463317200, 1463320800, 1463324400, 1463328000, 1463331600, 1463335200, 
    1463338800, 1463342400, 1463346000, 1463349600, 1463353200, 1463356800, 
    1463360400, 1463364000, 1463367600, 1463371200, 1463374800, 1463378400, 
    1463382000, 1463385600, 1463389200, 1463392800, 1463396400, 1463400000, 
    1463403600, 1463407200, 1463410800, 1463414400, 1463418000, 1463421600, 
    1463425200, 1463428800, 1463432400, 1463436000, 1463439600, 1463443200, 
    1463446800, 1463450400, 1463454000, 1463457600, 1463461200, 1463464800, 
    1463468400, 1463472000, 1463475600, 1463479200, 1463482800, 1463486400, 
    1463490000, 1463493600, 1463497200, 1463500800, 1463504400, 1463508000, 
    1463511600, 1463515200, 1463518800, 1463522400, 1463526000, 1463529600, 
    1463533200, 1463536800, 1463540400, 1463544000, 1463547600, 1463551200, 
    1463554800, 1463558400, 1463562000, 1463565600, 1463569200, 1463572800, 
    1463576400, 1463580000, 1463583600, 1463587200, 1463590800, 1463594400, 
    1463598000, 1463601600, 1463605200, 1463608800, 1463612400, 1463616000, 
    1463619600, 1463623200, 1463626800, 1463630400, 1463634000, 1463637600, 
    1463641200, 1463644800, 1463648400, 1463652000, 1463655600, 1463659200, 
    1463662800, 1463666400, 1463670000, 1463673600, 1463677200, 1463680800, 
    1463684400, 1463688000, 1463691600, 1463695200, 1463698800, 1463702400, 
    1463706000, 1463709600, 1463713200, 1463716800, 1463720400, 1463724000, 
    1463727600, 1463731200, 1463734800, 1463738400, 1463742000, 1463745600, 
    1463749200, 1463752800, 1463756400, 1463760000, 1463763600, 1463767200, 
    1463770800, 1463774400, 1463778000, 1463781600, 1463785200, 1463788800, 
    1463792400, 1463796000, 1463799600, 1463803200, 1463806800, 1463810400, 
    1463814000, 1463817600, 1463821200, 1463824800, 1463828400, 1463832000, 
    1463835600, 1463839200, 1463842800, 1463846400, 1463850000, 1463853600, 
    1463857200, 1463860800, 1463864400, 1463868000, 1463871600, 1463875200, 
    1463878800, 1463882400, 1463886000, 1463889600, 1463893200, 1463896800, 
    1463900400, 1463904000, 1463907600, 1463911200, 1463914800, 1463918400, 
    1463922000, 1463925600, 1463929200, 1463932800, 1463936400, 1463940000, 
    1463943600, 1463947200, 1463950800, 1463954400, 1463958000, 1463961600, 
    1463965200, 1463968800, 1463972400, 1463976000, 1463979600, 1463983200, 
    1463986800, 1463990400, 1463994000, 1463997600, 1464001200, 1464004800, 
    1464008400, 1464012000, 1464015600, 1464019200, 1464022800, 1464026400, 
    1464030000, 1464033600, 1464037200, 1464040800, 1464044400, 1464048000, 
    1464051600, 1464055200, 1464058800, 1464062400, 1464066000, 1464069600, 
    1464073200, 1464076800, 1464080400, 1464084000, 1464087600, 1464091200, 
    1464094800, 1464098400, 1464102000, 1464105600, 1464109200, 1464112800, 
    1464116400, 1464120000, 1464123600, 1464127200, 1464130800, 1464134400, 
    1464138000, 1464141600, 1464145200, 1464148800, 1464152400, 1464156000, 
    1464159600, 1464163200, 1464166800, 1464170400, 1464174000, 1464177600, 
    1464181200, 1464184800, 1464188400, 1464192000, 1464195600, 1464199200, 
    1464202800, 1464206400, 1464210000, 1464213600, 1464217200, 1464220800, 
    1464224400, 1464228000, 1464231600, 1464235200, 1464238800, 1464242400, 
    1464246000, 1464249600, 1464253200, 1464256800, 1464260400, 1464264000, 
    1464267600, 1464271200, 1464274800, 1464278400, 1464282000, 1464285600, 
    1464289200, 1464292800, 1464296400, 1464300000, 1464303600, 1464307200, 
    1464310800, 1464314400, 1464318000, 1464321600, 1464325200, 1464328800, 
    1464332400, 1464336000, 1464339600, 1464343200, 1464346800, 1464350400, 
    1464354000, 1464357600, 1464361200, 1464364800, 1464368400, 1464372000, 
    1464375600, 1464379200, 1464382800, 1464386400, 1464390000, 1464393600, 
    1464397200, 1464400800, 1464404400, 1464408000, 1464411600, 1464415200, 
    1464418800, 1464422400, 1464426000, 1464429600, 1464433200, 1464436800, 
    1464440400, 1464444000, 1464447600, 1464451200, 1464454800, 1464458400, 
    1464462000, 1464465600, 1464469200, 1464472800, 1464476400, 1464480000, 
    1464483600, 1464487200, 1464490800, 1464494400, 1464498000, 1464501600, 
    1464505200, 1464508800, 1464512400, 1464516000, 1464519600, 1464523200, 
    1464526800, 1464530400, 1464534000, 1464537600, 1464541200, 1464544800, 
    1464548400, 1464552000, 1464555600, 1464559200, 1464562800, 1464566400, 
    1464570000, 1464573600, 1464577200, 1464580800, 1464584400, 1464588000, 
    1464591600, 1464595200, 1464598800, 1464602400, 1464606000, 1464609600, 
    1464613200, 1464616800, 1464620400, 1464624000, 1464627600, 1464631200, 
    1464634800, 1464638400, 1464642000, 1464645600, 1464649200, 1464652800, 
    1464656400, 1464660000, 1464663600, 1464667200, 1464670800, 1464674400, 
    1464678000, 1464681600, 1464685200, 1464688800, 1464692400, 1464696000, 
    1464699600, 1464703200, 1464706800, 1464710400, 1464714000, 1464717600, 
    1464721200, 1464724800, 1464728400, 1464732000, 1464735600, 1464739200, 
    1464742800, 1464746400, 1464750000, 1464753600, 1464757200, 1464760800, 
    1464764400, 1464768000, 1464771600, 1464775200, 1464778800, 1464782400, 
    1464786000, 1464789600, 1464793200, 1464796800, 1464800400, 1464804000, 
    1464807600, 1464811200, 1464814800, 1464818400, 1464822000, 1464825600, 
    1464829200, 1464832800, 1464836400, 1464840000, 1464843600, 1464847200, 
    1464850800, 1464854400, 1464858000, 1464861600, 1464865200, 1464868800, 
    1464872400, 1464876000, 1464879600, 1464883200, 1464886800, 1464890400, 
    1464894000, 1464897600, 1464901200, 1464904800, 1464908400, 1464912000, 
    1464915600, 1464919200, 1464922800, 1464926400, 1464930000, 1464933600, 
    1464937200, 1464940800, 1464944400, 1464948000, 1464951600, 1464955200, 
    1464958800, 1464962400, 1464966000, 1464969600, 1464973200, 1464976800, 
    1464980400, 1464984000, 1464987600, 1464991200, 1464994800, 1464998400, 
    1465002000, 1465005600, 1465009200, 1465012800, 1465016400, 1465020000, 
    1465023600, 1465027200, 1465030800, 1465034400, 1465038000, 1465041600, 
    1465045200, 1465048800, 1465052400, 1465056000, 1465059600, 1465063200, 
    1465066800, 1465070400, 1465074000, 1465077600, 1465081200, 1465084800, 
    1465088400, 1465092000, 1465095600, 1465099200, 1465102800, 1465106400, 
    1465110000, 1465113600, 1465117200, 1465120800, 1465124400, 1465128000, 
    1465131600, 1465135200, 1465138800, 1465142400, 1465146000, 1465149600, 
    1465153200, 1465156800, 1465160400, 1465164000, 1465167600, 1465171200, 
    1465174800, 1465178400, 1465182000, 1465185600, 1465189200, 1465192800, 
    1465196400, 1465200000, 1465203600, 1465207200, 1465210800, 1465214400, 
    1465218000, 1465221600, 1465225200, 1465228800, 1465232400, 1465236000, 
    1465239600, 1465243200, 1465246800, 1465250400, 1465254000, 1465257600, 
    1465261200, 1465264800, 1465268400, 1465272000, 1465275600, 1465279200, 
    1465282800, 1465286400, 1465290000, 1465293600, 1465297200, 1465300800, 
    1465304400, 1465308000, 1465311600, 1465315200, 1465318800, 1465322400, 
    1465326000, 1465329600, 1465333200, 1465336800, 1465340400, 1465344000, 
    1465347600, 1465351200, 1465354800, 1465358400, 1465362000, 1465365600, 
    1465369200, 1465372800, 1465376400, 1465380000, 1465383600, 1465387200, 
    1465390800, 1465394400, 1465398000, 1465401600, 1465405200, 1465408800, 
    1465412400, 1465416000, 1465419600, 1465423200, 1465426800, 1465430400, 
    1465434000, 1465437600, 1465441200, 1465444800, 1465448400, 1465452000, 
    1465455600, 1465459200, 1465462800, 1465466400, 1465470000, 1465473600, 
    1465477200, 1465480800, 1465484400, 1465488000, 1465491600, 1465495200, 
    1465498800, 1465502400, 1465506000, 1465509600, 1465513200, 1465516800, 
    1465520400, 1465524000, 1465527600, 1465531200, 1465534800, 1465538400, 
    1465542000, 1465545600, 1465549200, 1465552800, 1465556400, 1465560000, 
    1465563600, 1465567200, 1465570800, 1465574400, 1465578000, 1465581600, 
    1465585200, 1465588800, 1465592400, 1465596000, 1465599600, 1465603200, 
    1465606800, 1465610400, 1465614000, 1465617600, 1465621200, 1465624800, 
    1465628400, 1465632000, 1465635600, 1465639200, 1465642800, 1465646400, 
    1465650000, 1465653600, 1465657200, 1465660800, 1465664400, 1465668000, 
    1465671600, 1465675200, 1465678800, 1465682400, 1465686000, 1465689600, 
    1465693200, 1465696800, 1465700400, 1465704000, 1465707600, 1465711200, 
    1465714800, 1465718400, 1465722000, 1465725600, 1465729200, 1465732800, 
    1465736400, 1465740000, 1465743600, 1465747200, 1465750800, 1465754400, 
    1465758000, 1465761600, 1465765200, 1465768800, 1465772400, 1465776000, 
    1465779600, 1465783200, 1465786800, 1465790400, 1465794000, 1465797600, 
    1465801200, 1465804800, 1465808400, 1465812000, 1465815600, 1465819200, 
    1465822800, 1465826400, 1465830000, 1465833600, 1465837200, 1465840800, 
    1465844400, 1465848000, 1465851600, 1465855200, 1465858800, 1465862400, 
    1465866000, 1465869600, 1465873200, 1465876800, 1465880400, 1465884000, 
    1465887600, 1465891200, 1465894800, 1465898400, 1465902000, 1465905600, 
    1465909200, 1465912800, 1465916400, 1465920000, 1465923600, 1465927200, 
    1465930800, 1465934400, 1465938000, 1465941600, 1465945200, 1465948800, 
    1465952400, 1465956000, 1465959600, 1465963200, 1465966800, 1465970400, 
    1465974000, 1465977600, 1465981200, 1465984800, 1465988400, 1465992000, 
    1465995600, 1465999200, 1466002800, 1466006400, 1466010000, 1466013600, 
    1466017200, 1466020800, 1466024400, 1466028000, 1466031600, 1466035200, 
    1466038800, 1466042400, 1466046000, 1466049600, 1466053200, 1466056800, 
    1466060400, 1466064000, 1466067600, 1466071200, 1466074800, 1466078400, 
    1466082000, 1466085600, 1466089200, 1466092800, 1466096400, 1466100000, 
    1466103600, 1466107200, 1466110800, 1466114400, 1466118000, 1466121600, 
    1466125200, 1466128800, 1466132400, 1466136000, 1466139600, 1466143200, 
    1466146800, 1466150400, 1466154000, 1466157600, 1466161200, 1466164800, 
    1466168400, 1466172000, 1466175600, 1466179200, 1466182800, 1466186400, 
    1466190000, 1466193600, 1466197200, 1466200800, 1466204400, 1466208000, 
    1466211600, 1466215200, 1466218800, 1466222400, 1466226000, 1466229600, 
    1466233200, 1466236800, 1466240400, 1466244000, 1466247600, 1466251200, 
    1466254800, 1466258400, 1466262000, 1466265600, 1466269200, 1466272800, 
    1466276400, 1466280000, 1466283600, 1466287200, 1466290800, 1466294400, 
    1466298000, 1466301600, 1466305200, 1466308800, 1466312400, 1466316000, 
    1466319600, 1466323200, 1466326800, 1466330400, 1466334000, 1466337600, 
    1466341200, 1466344800, 1466348400, 1466352000, 1466355600, 1466359200, 
    1466362800, 1466366400, 1466370000, 1466373600, 1466377200, 1466380800, 
    1466384400, 1466388000, 1466391600, 1466395200, 1466398800, 1466402400, 
    1466406000, 1466409600, 1466413200, 1466416800, 1466420400, 1466424000, 
    1466427600, 1466431200, 1466434800, 1466438400, 1466442000, 1466445600, 
    1466449200, 1466452800, 1466456400, 1466460000, 1466463600, 1466467200, 
    1466470800, 1466474400, 1466478000, 1466481600, 1466485200, 1466488800, 
    1466492400, 1466496000, 1466499600, 1466503200, 1466506800, 1466510400, 
    1466514000, 1466517600, 1466521200, 1466524800, 1466528400, 1466532000, 
    1466535600, 1466539200, 1466542800, 1466546400, 1466550000, 1466553600, 
    1466557200, 1466560800, 1466564400, 1466568000, 1466571600, 1466575200, 
    1466578800, 1466582400, 1466586000, 1466589600, 1466593200, 1466596800, 
    1466600400, 1466604000, 1466607600, 1466611200, 1466614800, 1466618400, 
    1466622000, 1466625600, 1466629200, 1466632800, 1466636400, 1466640000, 
    1466643600, 1466647200, 1466650800, 1466654400, 1466658000, 1466661600, 
    1466665200, 1466668800, 1466672400, 1466676000, 1466679600, 1466683200, 
    1466686800, 1466690400, 1466694000, 1466697600, 1466701200, 1466704800, 
    1466708400, 1466712000, 1466715600, 1466719200, 1466722800, 1466726400, 
    1466730000, 1466733600, 1466737200, 1466740800, 1466744400, 1466748000, 
    1466751600, 1466755200, 1466758800, 1466762400, 1466766000, 1466769600, 
    1466773200, 1466776800, 1466780400, 1466784000, 1466787600, 1466791200, 
    1466794800, 1466798400, 1466802000, 1466805600, 1466809200, 1466812800, 
    1466816400, 1466820000, 1466823600, 1466827200, 1466830800, 1466834400, 
    1466838000, 1466841600, 1466845200, 1466848800, 1466852400, 1466856000, 
    1466859600, 1466863200, 1466866800, 1466870400, 1466874000, 1466877600, 
    1466881200, 1466884800, 1466888400, 1466892000, 1466895600, 1466899200, 
    1466902800, 1466906400, 1466910000, 1466913600, 1466917200, 1466920800, 
    1466924400, 1466928000, 1466931600, 1466935200, 1466938800, 1466942400, 
    1466946000, 1466949600, 1466953200, 1466956800, 1466960400, 1466964000, 
    1466967600, 1466971200, 1466974800, 1466978400, 1466982000, 1466985600, 
    1466989200, 1466992800, 1466996400, 1467000000, 1467003600, 1467007200, 
    1467010800, 1467014400, 1467018000, 1467021600, 1467025200, 1467028800, 
    1467032400, 1467036000, 1467039600, 1467043200, 1467046800, 1467050400, 
    1467054000, 1467057600, 1467061200, 1467064800, 1467068400, 1467072000, 
    1467075600, 1467079200, 1467082800, 1467086400, 1467090000, 1467093600, 
    1467097200, 1467100800, 1467104400, 1467108000, 1467111600, 1467115200, 
    1467118800, 1467122400, 1467126000, 1467129600, 1467133200, 1467136800, 
    1467140400, 1467144000, 1467147600, 1467151200, 1467154800, 1467158400, 
    1467162000, 1467165600, 1467169200, 1467172800, 1467176400, 1467180000, 
    1467183600, 1467187200, 1467190800, 1467194400, 1467198000, 1467201600, 
    1467205200, 1467208800, 1467212400, 1467216000, 1467219600, 1467223200, 
    1467226800, 1467230400, 1467234000, 1467237600, 1467241200, 1467244800, 
    1467248400, 1467252000, 1467255600, 1467259200, 1467262800, 1467266400, 
    1467270000, 1467273600, 1467277200, 1467280800, 1467284400, 1467288000, 
    1467291600, 1467295200, 1467298800, 1467302400, 1467306000, 1467309600, 
    1467313200, 1467316800, 1467320400, 1467324000, 1467327600, 1467331200, 
    1467334800, 1467338400, 1467342000, 1467345600, 1467349200, 1467352800, 
    1467356400, 1467360000, 1467363600, 1467367200, 1467370800, 1467374400, 
    1467378000, 1467381600, 1467385200, 1467388800, 1467392400, 1467396000, 
    1467399600, 1467403200, 1467406800, 1467410400, 1467414000, 1467417600, 
    1467421200, 1467424800, 1467428400, 1467432000, 1467435600, 1467439200, 
    1467442800, 1467446400, 1467450000, 1467453600, 1467457200, 1467460800, 
    1467464400, 1467468000, 1467471600, 1467475200, 1467478800, 1467482400, 
    1467486000, 1467489600, 1467493200, 1467496800, 1467500400, 1467504000, 
    1467507600, 1467511200, 1467514800, 1467518400, 1467522000, 1467525600, 
    1467529200, 1467532800, 1467536400, 1467540000, 1467543600, 1467547200, 
    1467550800, 1467554400, 1467558000, 1467561600, 1467565200, 1467568800, 
    1467572400, 1467576000, 1467579600, 1467583200, 1467586800, 1467590400, 
    1467594000, 1467597600, 1467601200, 1467604800, 1467608400, 1467612000, 
    1467615600, 1467619200, 1467622800, 1467626400, 1467630000, 1467633600, 
    1467637200, 1467640800, 1467644400, 1467648000, 1467651600, 1467655200, 
    1467658800, 1467662400, 1467666000, 1467669600, 1467673200, 1467676800, 
    1467680400, 1467684000, 1467687600, 1467691200, 1467694800, 1467698400, 
    1467702000, 1467705600, 1467709200, 1467712800, 1467716400, 1467720000, 
    1467723600, 1467727200, 1467730800, 1467734400, 1467738000, 1467741600, 
    1467745200, 1467748800, 1467752400, 1467756000, 1467759600, 1467763200, 
    1467766800, 1467770400, 1467774000, 1467777600, 1467781200, 1467784800, 
    1467788400, 1467792000, 1467795600, 1467799200, 1467802800, 1467806400, 
    1467810000, 1467813600, 1467817200, 1467820800, 1467824400, 1467828000, 
    1467831600, 1467835200, 1467838800, 1467842400, 1467846000, 1467849600, 
    1467853200, 1467856800, 1467860400, 1467864000, 1467867600, 1467871200, 
    1467874800, 1467878400, 1467882000, 1467885600, 1467889200, 1467892800, 
    1467896400, 1467900000, 1467903600, 1467907200, 1467910800, 1467914400, 
    1467918000, 1467921600, 1467925200, 1467928800, 1467932400, 1467936000, 
    1467939600, 1467943200, 1467946800, 1467950400, 1467954000, 1467957600, 
    1467961200, 1467964800, 1467968400, 1467972000, 1467975600, 1467979200, 
    1467982800, 1467986400, 1467990000, 1467993600, 1467997200, 1468000800, 
    1468004400, 1468008000, 1468011600, 1468015200, 1468018800, 1468022400, 
    1468026000, 1468029600, 1468033200, 1468036800, 1468040400, 1468044000, 
    1468047600, 1468051200, 1468054800, 1468058400, 1468062000, 1468065600, 
    1468069200, 1468072800, 1468076400, 1468080000, 1468083600, 1468087200, 
    1468090800, 1468094400, 1468098000, 1468101600, 1468105200, 1468108800, 
    1468112400, 1468116000, 1468119600, 1468123200, 1468126800, 1468130400, 
    1468134000, 1468137600, 1468141200, 1468144800, 1468148400, 1468152000, 
    1468155600, 1468159200, 1468162800, 1468166400, 1468170000, 1468173600, 
    1468177200, 1468180800, 1468184400, 1468188000, 1468191600, 1468195200, 
    1468198800, 1468202400, 1468206000, 1468209600, 1468213200, 1468216800, 
    1468220400, 1468224000, 1468227600, 1468231200, 1468234800, 1468238400, 
    1468242000, 1468245600, 1468249200, 1468252800, 1468256400, 1468260000, 
    1468263600, 1468267200, 1468270800, 1468274400, 1468278000, 1468281600, 
    1468285200, 1468288800, 1468292400, 1468296000, 1468299600, 1468303200, 
    1468306800, 1468310400, 1468314000, 1468317600, 1468321200, 1468324800, 
    1468328400, 1468332000, 1468335600, 1468339200, 1468342800, 1468346400, 
    1468350000, 1468353600, 1468357200, 1468360800, 1468364400, 1468368000, 
    1468371600, 1468375200, 1468378800, 1468382400, 1468386000, 1468389600, 
    1468393200, 1468396800, 1468400400, 1468404000, 1468407600, 1468411200, 
    1468414800, 1468418400, 1468422000, 1468425600, 1468429200, 1468432800, 
    1468436400, 1468440000, 1468443600, 1468447200, 1468450800, 1468454400, 
    1468458000, 1468461600, 1468465200, 1468468800, 1468472400, 1468476000, 
    1468479600, 1468483200, 1468486800, 1468490400, 1468494000, 1468497600, 
    1468501200, 1468504800, 1468508400, 1468512000, 1468515600, 1468519200, 
    1468522800, 1468526400, 1468530000, 1468533600, 1468537200, 1468540800, 
    1468544400, 1468548000, 1468551600, 1468555200, 1468558800, 1468562400, 
    1468566000, 1468569600, 1468573200, 1468576800, 1468580400, 1468584000, 
    1468587600, 1468591200, 1468594800, 1468598400, 1468602000, 1468605600, 
    1468609200, 1468612800, 1468616400, 1468620000, 1468623600, 1468627200, 
    1468630800, 1468634400, 1468638000, 1468641600, 1468645200, 1468648800, 
    1468652400, 1468656000, 1468659600, 1468663200, 1468666800, 1468670400, 
    1468674000, 1468677600, 1468681200, 1468684800, 1468688400, 1468692000, 
    1468695600, 1468699200, 1468702800, 1468706400, 1468710000, 1468713600, 
    1468717200, 1468720800, 1468724400, 1468728000, 1468731600, 1468735200, 
    1468738800, 1468742400, 1468746000, 1468749600, 1468753200, 1468756800, 
    1468760400, 1468764000, 1468767600, 1468771200, 1468774800, 1468778400, 
    1468782000, 1468785600, 1468789200, 1468792800, 1468796400, 1468800000, 
    1468803600, 1468807200, 1468810800, 1468814400, 1468818000, 1468821600, 
    1468825200, 1468828800, 1468832400, 1468836000, 1468839600, 1468843200, 
    1468846800, 1468850400, 1468854000, 1468857600, 1468861200, 1468864800, 
    1468868400, 1468872000, 1468875600, 1468879200, 1468882800, 1468886400, 
    1468890000, 1468893600, 1468897200, 1468900800, 1468904400, 1468908000, 
    1468911600, 1468915200, 1468918800, 1468922400, 1468926000, 1468929600, 
    1468933200, 1468936800, 1468940400, 1468944000, 1468947600, 1468951200, 
    1468954800, 1468958400, 1468962000, 1468965600, 1468969200, 1468972800, 
    1468976400, 1468980000, 1468983600, 1468987200, 1468990800, 1468994400, 
    1468998000, 1469001600, 1469005200, 1469008800, 1469012400, 1469016000, 
    1469019600, 1469023200, 1469026800, 1469030400, 1469034000, 1469037600, 
    1469041200, 1469044800, 1469048400, 1469052000, 1469055600, 1469059200, 
    1469062800, 1469066400, 1469070000, 1469073600, 1469077200, 1469080800, 
    1469084400, 1469088000, 1469091600, 1469095200, 1469098800, 1469102400, 
    1469106000, 1469109600, 1469113200, 1469116800, 1469120400, 1469124000, 
    1469127600, 1469131200, 1469134800, 1469138400, 1469142000, 1469145600, 
    1469149200, 1469152800, 1469156400, 1469160000, 1469163600, 1469167200, 
    1469170800, 1469174400, 1469178000, 1469181600, 1469185200, 1469188800, 
    1469192400, 1469196000, 1469199600, 1469203200, 1469206800, 1469210400, 
    1469214000, 1469217600, 1469221200, 1469224800, 1469228400, 1469232000, 
    1469235600, 1469239200, 1469242800, 1469246400, 1469250000, 1469253600, 
    1469257200, 1469260800, 1469264400, 1469268000, 1469271600, 1469275200, 
    1469278800, 1469282400, 1469286000, 1469289600, 1469293200, 1469296800, 
    1469300400, 1469304000, 1469307600, 1469311200, 1469314800, 1469318400, 
    1469322000, 1469325600, 1469329200, 1469332800, 1469336400, 1469340000, 
    1469343600, 1469347200, 1469350800, 1469354400, 1469358000, 1469361600, 
    1469365200, 1469368800, 1469372400, 1469376000, 1469379600, 1469383200, 
    1469386800, 1469390400, 1469394000, 1469397600, 1469401200, 1469404800, 
    1469408400, 1469412000, 1469415600, 1469419200, 1469422800, 1469426400, 
    1469430000, 1469433600, 1469437200, 1469440800, 1469444400, 1469448000, 
    1469451600, 1469455200, 1469458800, 1469462400, 1469466000, 1469469600, 
    1469473200, 1469476800, 1469480400, 1469484000, 1469487600, 1469491200, 
    1469494800, 1469498400, 1469502000, 1469505600, 1469509200, 1469512800, 
    1469516400, 1469520000, 1469523600, 1469527200, 1469530800, 1469534400, 
    1469538000, 1469541600, 1469545200, 1469548800, 1469552400, 1469556000, 
    1469559600, 1469563200, 1469566800, 1469570400, 1469574000, 1469577600, 
    1469581200, 1469584800, 1469588400, 1469592000, 1469595600, 1469599200, 
    1469602800, 1469606400, 1469610000, 1469613600, 1469617200, 1469620800, 
    1469624400, 1469628000, 1469631600, 1469635200, 1469638800, 1469642400, 
    1469646000, 1469649600, 1469653200, 1469656800, 1469660400, 1469664000, 
    1469667600, 1469671200, 1469674800, 1469678400, 1469682000, 1469685600, 
    1469689200, 1469692800, 1469696400, 1469700000, 1469703600, 1469707200, 
    1469710800, 1469714400, 1469718000, 1469721600, 1469725200, 1469728800, 
    1469732400, 1469736000, 1469739600, 1469743200, 1469746800, 1469750400, 
    1469754000, 1469757600, 1469761200, 1469764800, 1469768400, 1469772000, 
    1469775600, 1469779200, 1469782800, 1469786400, 1469790000, 1469793600, 
    1469797200, 1469800800, 1469804400, 1469808000, 1469811600, 1469815200, 
    1469818800, 1469822400, 1469826000, 1469829600, 1469833200, 1469836800, 
    1469840400, 1469844000, 1469847600, 1469851200, 1469854800, 1469858400, 
    1469862000, 1469865600, 1469869200, 1469872800, 1469876400, 1469880000, 
    1469883600, 1469887200, 1469890800, 1469894400, 1469898000, 1469901600, 
    1469905200, 1469908800, 1469912400, 1469916000, 1469919600, 1469923200, 
    1469926800, 1469930400, 1469934000, 1469937600, 1469941200, 1469944800, 
    1469948400, 1469952000, 1469955600, 1469959200, 1469962800, 1469966400, 
    1469970000, 1469973600, 1469977200, 1469980800, 1469984400, 1469988000, 
    1469991600, 1469995200, 1469998800, 1470002400, 1470006000, 1470009600, 
    1470013200, 1470016800, 1470020400, 1470024000, 1470027600, 1470031200, 
    1470034800, 1470038400, 1470042000, 1470045600, 1470049200, 1470052800, 
    1470056400, 1470060000, 1470063600, 1470067200, 1470070800, 1470074400, 
    1470078000, 1470081600, 1470085200, 1470088800, 1470092400, 1470096000, 
    1470099600, 1470103200, 1470106800, 1470110400, 1470114000, 1470117600, 
    1470121200, 1470124800, 1470128400, 1470132000, 1470135600, 1470139200, 
    1470142800, 1470146400, 1470150000, 1470153600, 1470157200, 1470160800, 
    1470164400, 1470168000, 1470171600, 1470175200, 1470178800, 1470182400, 
    1470186000, 1470189600, 1470193200, 1470196800, 1470200400, 1470204000, 
    1470207600, 1470211200, 1470214800, 1470218400, 1470222000, 1470225600, 
    1470229200, 1470232800, 1470236400, 1470240000, 1470243600, 1470247200, 
    1470250800, 1470254400, 1470258000, 1470261600, 1470265200, 1470268800, 
    1470272400, 1470276000, 1470279600, 1470283200, 1470286800, 1470290400, 
    1470294000, 1470297600, 1470301200, 1470304800, 1470308400, 1470312000, 
    1470315600, 1470319200, 1470322800, 1470326400, 1470330000, 1470333600, 
    1470337200, 1470340800, 1470344400, 1470348000, 1470351600, 1470355200, 
    1470358800, 1470362400, 1470366000, 1470369600, 1470373200, 1470376800, 
    1470380400, 1470384000, 1470387600, 1470391200, 1470394800, 1470398400, 
    1470402000, 1470405600, 1470409200, 1470412800, 1470416400, 1470420000, 
    1470423600, 1470427200, 1470430800, 1470434400, 1470438000, 1470441600, 
    1470445200, 1470448800, 1470452400, 1470456000, 1470459600, 1470463200, 
    1470466800, 1470470400, 1470474000, 1470477600, 1470481200, 1470484800, 
    1470488400, 1470492000, 1470495600, 1470499200, 1470502800, 1470506400, 
    1470510000, 1470513600, 1470517200, 1470520800, 1470524400, 1470528000, 
    1470531600, 1470535200, 1470538800, 1470542400, 1470546000, 1470549600, 
    1470553200, 1470556800, 1470560400, 1470564000, 1470567600, 1470571200, 
    1470574800, 1470578400, 1470582000, 1470585600, 1470589200, 1470592800, 
    1470596400, 1470600000, 1470603600, 1470607200, 1470610800, 1470614400, 
    1470618000, 1470621600, 1470625200, 1470628800, 1470632400, 1470636000, 
    1470639600, 1470643200, 1470646800, 1470650400, 1470654000, 1470657600, 
    1470661200, 1470664800, 1470668400, 1470672000, 1470675600, 1470679200, 
    1470682800, 1470686400, 1470690000, 1470693600, 1470697200, 1470700800, 
    1470704400, 1470708000, 1470711600, 1470715200, 1470718800, 1470722400, 
    1470726000, 1470729600, 1470736800, 1470740400, 1470744000, 1470747600, 
    1470751200, 1470754800, 1470758400, 1470762000, 1470765600, 1470769200, 
    1470772800, 1470776400, 1470780000, 1470783600, 1470787200, 1470790800, 
    1470794400, 1470798000, 1470801600, 1470805200, 1470808800, 1470812400, 
    1470816000, 1470819600, 1470823200, 1470826800, 1470830400, 1470834000, 
    1470837600, 1470841200, 1470844800, 1470848400, 1470852000, 1470855600, 
    1470859200, 1470862800, 1470866400, 1470870000, 1470873600, 1470877200, 
    1470880800, 1470884400, 1470888000, 1470891600, 1470895200, 1470898800, 
    1470902400, 1470906000, 1470909600, 1470913200, 1470916800, 1470920400, 
    1470924000, 1470927600, 1470931200, 1470934800, 1470938400, 1470942000, 
    1470945600, 1470949200, 1470952800, 1470956400, 1470960000, 1470963600, 
    1470967200, 1470970800, 1470974400, 1470978000, 1470981600, 1470985200, 
    1470988800, 1470992400, 1470996000, 1470999600, 1471003200, 1471006800, 
    1471010400, 1471014000, 1471017600, 1471021200, 1471024800, 1471028400, 
    1471032000, 1471035600, 1471039200, 1471042800, 1471046400, 1471050000, 
    1471053600, 1471057200, 1471060800, 1471064400, 1471068000, 1471071600, 
    1471075200, 1471078800, 1471082400, 1471086000, 1471089600, 1471093200, 
    1471096800, 1471100400, 1471104000, 1471107600, 1471111200, 1471114800, 
    1471118400, 1471122000, 1471125600, 1471129200, 1471132800, 1471136400, 
    1471140000, 1471143600, 1471147200, 1471150800, 1471154400, 1471158000, 
    1471161600, 1471165200, 1471168800, 1471172400, 1471176000, 1471179600, 
    1471183200, 1471186800, 1471190400, 1471194000, 1471197600, 1471201200, 
    1471204800, 1471208400, 1471212000, 1471215600, 1471219200, 1471222800, 
    1471226400, 1471230000, 1471233600, 1471237200, 1471240800, 1471244400, 
    1471248000, 1471251600, 1471255200, 1471258800, 1471262400, 1471266000, 
    1471269600, 1471273200, 1471276800, 1471280400, 1471284000, 1471287600, 
    1471291200, 1471294800, 1471298400, 1471302000, 1471305600, 1471309200, 
    1471312800, 1471316400, 1471320000, 1471323600, 1471327200, 1471330800, 
    1471334400, 1471338000, 1471341600, 1471345200, 1471348800, 1471352400, 
    1471356000, 1471359600, 1471363200, 1471366800, 1471370400, 1471374000, 
    1471377600, 1471381200, 1471384800, 1471388400, 1471392000, 1471395600, 
    1471399200, 1471402800, 1471406400, 1471410000, 1471413600, 1471417200, 
    1471420800, 1471424400, 1471428000, 1471431600, 1471435200, 1471438800, 
    1471442400, 1471446000, 1471449600, 1471453200, 1471456800, 1471460400, 
    1471464000, 1471467600, 1471471200, 1471474800, 1471478400, 1471482000, 
    1471485600, 1471489200, 1471492800, 1471496400, 1471500000, 1471503600, 
    1471507200, 1471510800, 1471514400, 1471518000, 1471521600, 1471525200, 
    1471528800, 1471532400, 1471536000, 1471539600, 1471543200, 1471546800, 
    1471550400, 1471554000, 1471557600, 1471561200, 1471564800, 1471568400, 
    1471572000, 1471575600, 1471579200, 1471582800, 1471586400, 1471590000, 
    1471593600, 1471597200, 1471600800, 1471604400, 1471608000, 1471611600, 
    1471615200, 1471618800, 1471622400, 1471626000, 1471629600, 1471633200, 
    1471636800, 1471640400, 1471644000, 1471647600, 1471651200, 1471654800, 
    1471658400, 1471662000, 1471665600, 1471669200, 1471672800, 1471676400, 
    1471680000, 1471683600, 1471687200, 1471690800, 1471694400, 1471698000, 
    1471701600, 1471705200, 1471708800, 1471712400, 1471716000, 1471719600, 
    1471723200, 1471726800, 1471730400, 1471734000, 1471737600, 1471741200, 
    1471744800, 1471748400, 1471752000, 1471755600, 1471759200, 1471762800, 
    1471766400, 1471770000, 1471773600, 1471777200, 1471780800, 1471784400, 
    1471788000, 1471791600, 1471795200, 1471798800, 1471802400, 1471806000, 
    1471809600, 1471813200, 1471816800, 1471820400, 1471824000, 1471827600, 
    1471831200, 1471834800, 1471838400, 1471842000, 1471845600, 1471849200, 
    1471852800, 1471856400, 1471860000, 1471863600, 1471867200, 1471870800, 
    1471874400, 1471878000, 1471881600, 1471885200, 1471888800, 1471892400, 
    1471896000, 1471899600, 1471903200, 1471906800, 1471910400, 1471914000, 
    1471917600, 1471921200, 1471924800, 1471928400, 1471932000, 1471935600, 
    1471939200, 1471942800, 1471946400, 1471950000, 1471953600, 1471957200, 
    1471960800, 1471964400, 1471968000, 1471971600, 1471975200, 1471978800, 
    1471982400, 1471986000, 1471989600, 1471993200, 1471996800, 1472000400, 
    1472004000, 1472007600, 1472011200, 1472014800, 1472018400, 1472022000, 
    1472025600, 1472029200, 1472032800, 1472036400, 1472040000, 1472043600, 
    1472047200, 1472050800, 1472054400, 1472058000, 1472061600, 1472065200, 
    1472068800, 1472072400, 1472076000, 1472079600, 1472083200, 1472086800, 
    1472090400, 1472094000, 1472097600, 1472101200, 1472104800, 1472108400, 
    1472112000, 1472115600, 1472119200, 1472122800, 1472126400, 1472130000, 
    1472133600, 1472137200, 1472140800, 1472144400, 1472148000, 1472151600, 
    1472155200, 1472158800, 1472162400, 1472166000, 1472169600, 1472173200, 
    1472176800, 1472180400, 1472184000, 1472187600, 1472191200, 1472194800, 
    1472198400, 1472202000, 1472205600, 1472209200, 1472212800, 1472216400, 
    1472220000, 1472223600, 1472227200, 1472230800, 1472234400, 1472238000, 
    1472241600, 1472245200, 1472248800, 1472252400, 1472256000, 1472259600, 
    1472263200, 1472266800, 1472270400, 1472274000, 1472277600, 1472281200, 
    1472284800, 1472288400, 1472292000, 1472295600, 1472299200, 1472302800, 
    1472306400, 1472310000, 1472313600, 1472317200, 1472320800, 1472324400, 
    1472328000, 1472331600, 1472335200, 1472338800, 1472342400, 1472346000, 
    1472349600, 1472353200, 1472356800, 1472360400, 1472364000, 1472367600, 
    1472371200, 1472374800, 1472378400, 1472382000, 1472385600, 1472389200, 
    1472392800, 1472396400, 1472400000, 1472403600, 1472407200, 1472410800, 
    1472414400, 1472418000, 1472421600, 1472425200, 1472428800, 1472432400, 
    1472436000, 1472439600, 1472443200, 1472446800, 1472450400, 1472454000, 
    1472457600, 1472461200, 1472464800, 1472468400, 1472472000, 1472475600, 
    1472479200, 1472482800, 1472486400, 1472490000, 1472493600, 1472497200, 
    1472500800, 1472504400, 1472508000, 1472511600, 1472515200, 1472518800, 
    1472522400, 1472526000, 1472529600, 1472533200, 1472536800, 1472540400, 
    1472544000, 1472547600, 1472551200, 1472554800, 1472558400, 1472562000, 
    1472565600, 1472569200, 1472572800, 1472576400, 1472580000, 1472583600, 
    1472587200, 1472590800, 1472594400, 1472598000, 1472601600, 1472605200, 
    1472608800, 1472612400, 1472616000, 1472619600, 1472623200, 1472626800, 
    1472630400, 1472634000, 1472637600, 1472641200, 1472644800, 1472648400, 
    1472652000, 1472655600, 1472659200, 1472662800, 1472666400, 1472670000, 
    1472673600, 1472677200, 1472680800, 1472684400, 1472688000, 1472691600, 
    1472695200, 1472698800, 1472702400, 1472706000, 1472709600, 1472713200, 
    1472716800, 1472720400, 1472724000, 1472727600, 1472731200, 1472734800, 
    1472738400, 1472742000, 1472745600, 1472749200, 1472752800, 1472756400, 
    1472760000, 1472763600, 1472767200, 1472770800, 1472774400, 1472778000, 
    1472781600, 1472785200, 1472788800, 1472792400, 1472796000, 1472799600, 
    1472803200, 1472806800, 1472810400, 1472814000, 1472817600, 1472821200, 
    1472824800, 1472828400, 1472832000, 1472835600, 1472839200, 1472842800, 
    1472846400, 1472850000, 1472853600, 1472857200, 1472860800, 1472864400, 
    1472868000, 1472871600, 1472875200, 1472878800, 1472882400, 1472886000, 
    1472889600, 1472893200, 1472896800, 1472900400, 1472904000, 1472907600, 
    1472911200, 1472914800, 1472918400, 1472922000, 1472925600, 1472929200, 
    1472932800, 1472936400, 1472940000, 1472943600, 1472947200, 1472950800, 
    1472954400, 1472958000, 1472961600, 1472965200, 1472968800, 1472972400, 
    1472976000, 1472979600, 1472983200, 1472986800, 1472990400, 1472994000, 
    1472997600, 1473001200, 1473004800, 1473008400, 1473012000, 1473015600, 
    1473019200, 1473022800, 1473026400, 1473030000, 1473033600, 1473037200, 
    1473040800, 1473044400, 1473048000, 1473051600, 1473055200, 1473058800, 
    1473062400, 1473066000, 1473069600, 1473073200, 1473076800, 1473080400, 
    1473084000, 1473087600, 1473091200, 1473094800, 1473098400, 1473102000, 
    1473105600, 1473109200, 1473112800, 1473116400, 1473120000, 1473123600, 
    1473127200, 1473130800, 1473134400, 1473138000, 1473141600, 1473145200, 
    1473148800, 1473152400, 1473156000, 1473159600, 1473163200, 1473166800, 
    1473170400, 1473174000, 1473177600, 1473181200, 1473184800, 1473188400, 
    1473192000, 1473195600, 1473199200, 1473202800, 1473206400, 1473210000, 
    1473213600, 1473217200, 1473220800, 1473224400, 1473228000, 1473231600, 
    1473235200, 1473238800, 1473242400, 1473246000, 1473249600, 1473253200, 
    1473256800, 1473260400, 1473264000, 1473267600, 1473271200, 1473274800, 
    1473278400, 1473282000, 1473285600, 1473289200, 1473292800, 1473296400, 
    1473300000, 1473303600, 1473307200, 1473310800, 1473314400, 1473318000, 
    1473321600, 1473325200, 1473328800, 1473332400, 1473336000, 1473339600, 
    1473343200, 1473346800, 1473350400, 1473354000, 1473357600, 1473361200, 
    1473364800, 1473368400, 1473372000, 1473375600, 1473379200, 1473382800, 
    1473386400, 1473390000, 1473393600, 1473397200, 1473400800, 1473404400, 
    1473408000, 1473411600, 1473415200, 1473418800, 1473422400, 1473426000, 
    1473429600, 1473433200, 1473436800, 1473440400, 1473444000, 1473447600, 
    1473451200, 1473454800, 1473458400, 1473462000, 1473465600, 1473469200, 
    1473472800, 1473476400, 1473480000, 1473483600, 1473487200, 1473490800, 
    1473494400, 1473498000, 1473501600, 1473505200, 1473508800, 1473512400, 
    1473516000, 1473519600, 1473523200, 1473526800, 1473530400, 1473534000, 
    1473537600, 1473541200, 1473544800, 1473548400, 1473552000, 1473555600, 
    1473559200, 1473562800, 1473566400, 1473570000, 1473573600, 1473577200, 
    1473580800, 1473584400, 1473588000, 1473591600, 1473595200, 1473598800, 
    1473602400, 1473606000, 1473609600, 1473613200, 1473616800, 1473620400, 
    1473624000, 1473627600, 1473631200, 1473634800, 1473638400, 1473642000, 
    1473645600, 1473649200, 1473652800, 1473656400, 1473660000, 1473663600, 
    1473667200, 1473670800, 1473674400, 1473678000, 1473681600, 1473685200, 
    1473688800, 1473692400, 1473696000, 1473699600, 1473703200, 1473706800, 
    1473710400, 1473714000, 1473717600, 1473721200, 1473724800, 1473728400, 
    1473732000, 1473735600, 1473739200, 1473742800, 1473746400, 1473750000, 
    1473753600, 1473757200, 1473760800, 1473764400, 1473768000, 1473771600, 
    1473775200, 1473778800, 1473782400, 1473786000, 1473789600, 1473793200, 
    1473796800, 1473800400, 1473804000, 1473807600, 1473811200, 1473814800, 
    1473818400, 1473822000, 1473825600, 1473829200, 1473832800, 1473836400, 
    1473840000, 1473843600, 1473847200, 1473850800, 1473854400, 1473858000, 
    1473861600, 1473865200, 1473868800, 1473872400, 1473876000, 1473879600, 
    1473883200, 1473886800, 1473890400, 1473894000, 1473897600, 1473901200, 
    1473904800, 1473908400, 1473912000, 1473915600, 1473919200, 1473922800, 
    1473926400, 1473930000, 1473933600, 1473937200, 1473940800, 1473944400, 
    1473948000, 1473951600, 1473955200, 1473958800, 1473962400, 1473966000, 
    1473969600, 1473973200, 1473976800, 1473980400, 1473984000, 1473987600, 
    1473991200, 1473994800, 1473998400, 1474002000, 1474005600, 1474009200, 
    1474012800, 1474016400, 1474020000, 1474023600, 1474027200, 1474030800, 
    1474034400, 1474038000, 1474041600, 1474045200, 1474048800, 1474052400, 
    1474056000, 1474059600, 1474063200, 1474066800, 1474070400, 1474074000, 
    1474077600, 1474081200, 1474084800, 1474088400, 1474092000, 1474095600, 
    1474099200, 1474102800, 1474106400, 1474110000, 1474113600, 1474117200, 
    1474120800, 1474124400, 1474128000, 1474131600, 1474135200, 1474138800, 
    1474142400, 1474146000, 1474149600, 1474153200, 1474156800, 1474160400, 
    1474164000, 1474167600, 1474171200, 1474174800, 1474178400, 1474182000, 
    1474185600, 1474189200, 1474192800, 1474196400, 1474200000, 1474203600, 
    1474207200, 1474210800, 1474214400, 1474218000, 1474221600, 1474225200, 
    1474228800, 1474232400, 1474236000, 1474239600, 1474243200, 1474246800, 
    1474250400, 1474254000, 1474257600, 1474261200, 1474264800, 1474268400, 
    1474272000, 1474275600, 1474279200, 1474282800, 1474286400, 1474290000, 
    1474293600, 1474297200, 1474300800, 1474304400, 1474308000, 1474311600, 
    1474315200, 1474318800, 1474322400, 1474326000, 1474329600, 1474333200, 
    1474336800, 1474340400, 1474344000, 1474347600, 1474351200, 1474354800, 
    1474358400, 1474362000, 1474365600, 1474369200, 1474372800, 1474376400, 
    1474380000, 1474383600, 1474387200, 1474390800, 1474394400, 1474398000, 
    1474401600, 1474405200, 1474408800, 1474412400, 1474416000, 1474419600, 
    1474423200, 1474426800, 1474430400, 1474434000, 1474437600, 1474441200, 
    1474444800, 1474448400, 1474452000, 1474455600, 1474459200, 1474462800, 
    1474466400, 1474470000, 1474473600, 1474477200, 1474480800, 1474484400, 
    1474488000, 1474491600, 1474495200, 1474498800, 1474502400, 1474506000, 
    1474509600, 1474513200, 1474516800, 1474520400, 1474524000, 1474527600, 
    1474531200, 1474534800, 1474538400, 1474542000, 1474545600, 1474549200, 
    1474552800, 1474556400, 1474560000, 1474563600, 1474567200, 1474570800, 
    1474574400, 1474578000, 1474581600, 1474585200, 1474588800, 1474592400, 
    1474596000, 1474599600, 1474603200, 1474606800, 1474610400, 1474614000, 
    1474617600, 1474621200, 1474624800, 1474628400, 1474632000, 1474635600, 
    1474639200, 1474642800, 1474646400, 1474650000, 1474653600, 1474657200, 
    1474660800, 1474664400, 1474668000, 1474671600, 1474675200, 1474678800, 
    1474682400, 1474686000, 1474689600, 1474693200, 1474696800, 1474700400, 
    1474704000, 1474707600, 1474711200, 1474714800, 1474718400, 1474722000, 
    1474725600, 1474729200, 1474732800, 1474736400, 1474740000, 1474743600, 
    1474747200, 1474750800, 1474754400, 1474758000, 1474761600, 1474765200, 
    1474768800, 1474772400, 1474776000, 1474779600, 1474783200, 1474786800, 
    1474790400, 1474794000, 1474797600, 1474801200, 1474804800, 1474808400, 
    1474812000, 1474815600, 1474819200, 1474822800, 1474826400, 1474830000, 
    1474833600, 1474837200, 1474840800, 1474844400, 1474848000, 1474851600, 
    1474855200, 1474858800, 1474862400, 1474866000, 1474869600, 1474873200, 
    1474876800, 1474880400, 1474884000, 1474887600, 1474891200, 1474894800, 
    1474898400, 1474902000, 1474905600, 1474909200, 1474912800, 1474916400, 
    1474920000, 1474923600, 1474927200, 1474930800, 1474934400, 1474938000, 
    1474941600, 1474945200, 1474948800, 1474952400, 1474956000, 1474959600, 
    1474963200, 1474966800, 1474970400, 1474974000, 1474977600, 1474981200, 
    1474984800, 1474988400, 1474992000, 1474995600, 1474999200, 1475002800, 
    1475006400, 1475010000, 1475013600, 1475017200, 1475020800, 1475024400, 
    1475028000, 1475031600, 1475035200, 1475038800, 1475042400, 1475046000, 
    1475049600, 1475053200, 1475056800, 1475060400, 1475064000, 1475067600, 
    1475071200, 1475074800, 1475078400, 1475082000, 1475085600, 1475089200, 
    1475092800, 1475096400, 1475100000, 1475103600, 1475107200, 1475110800, 
    1475114400, 1475118000, 1475121600, 1475125200, 1475128800, 1475132400, 
    1475136000, 1475139600, 1475143200, 1475146800, 1475150400, 1475154000, 
    1475157600, 1475161200, 1475164800, 1475168400, 1475172000, 1475175600, 
    1475179200, 1475182800, 1475186400, 1475190000, 1475193600, 1475197200, 
    1475200800, 1475204400, 1475208000, 1475211600, 1475215200, 1475218800, 
    1475222400, 1475226000, 1475229600, 1475233200, 1475236800, 1475240400, 
    1475244000, 1475247600, 1475251200, 1475254800, 1475258400, 1475262000, 
    1475265600, 1475269200, 1475272800, 1475276400, 1475280000, 1475283600, 
    1475287200, 1475290800, 1475294400, 1475298000, 1475301600, 1475305200, 
    1475308800, 1475312400, 1475316000, 1475319600, 1475323200, 1475326800, 
    1475330400, 1475334000, 1475337600, 1475341200, 1475344800, 1475348400, 
    1475352000, 1475355600, 1475359200, 1475362800, 1475366400, 1475370000, 
    1475373600, 1475377200, 1475380800, 1475384400, 1475388000, 1475391600, 
    1475395200, 1475398800, 1475402400, 1475406000, 1475409600, 1475413200, 
    1475416800, 1475420400, 1475424000, 1475427600, 1475431200, 1475434800, 
    1475438400, 1475442000, 1475445600, 1475449200, 1475452800, 1475456400, 
    1475460000, 1475463600, 1475467200, 1475470800, 1475474400, 1475478000, 
    1475481600, 1475485200, 1475488800, 1475492400, 1475496000, 1475499600, 
    1475503200, 1475506800, 1475510400, 1475514000, 1475517600, 1475521200, 
    1475524800, 1475528400, 1475532000, 1475535600, 1475539200, 1475542800, 
    1475546400, 1475550000, 1475553600, 1475557200, 1475560800, 1475564400, 
    1475568000, 1475571600, 1475575200, 1475578800, 1475582400, 1475586000, 
    1475589600, 1475593200, 1475596800, 1475600400, 1475604000, 1475607600, 
    1475611200, 1475614800, 1475618400, 1475622000, 1475625600, 1475629200, 
    1475632800, 1475636400, 1475640000, 1475643600, 1475647200, 1475650800, 
    1475654400, 1475658000, 1475661600, 1475665200, 1475668800, 1475672400, 
    1475676000, 1475679600, 1475683200, 1475686800, 1475690400, 1475694000, 
    1475697600, 1475701200, 1475704800, 1475708400, 1475712000, 1475715600, 
    1475719200, 1475722800, 1475726400, 1475730000, 1475733600, 1475737200, 
    1475740800, 1475744400, 1475748000, 1475751600, 1475755200, 1475758800, 
    1475762400, 1475766000, 1475769600, 1475773200, 1475776800, 1475780400, 
    1475784000, 1475787600, 1475791200, 1475794800, 1475798400, 1475802000, 
    1475805600, 1475809200, 1475812800, 1475816400, 1475820000, 1475823600, 
    1475827200, 1475830800, 1475834400, 1475838000, 1475841600, 1475845200, 
    1475848800, 1475852400, 1475856000, 1475859600, 1475863200, 1475866800, 
    1475870400, 1475874000, 1475877600, 1475881200, 1475884800, 1475888400, 
    1475892000, 1475895600, 1475899200, 1475902800, 1475906400, 1475910000, 
    1475913600, 1475917200, 1475920800, 1475924400, 1475928000, 1475931600, 
    1475935200, 1475938800, 1475942400, 1475946000, 1475949600, 1475953200, 
    1475956800, 1475960400, 1475964000, 1475967600, 1475971200, 1475974800, 
    1475978400, 1475982000, 1475985600, 1475989200, 1475992800, 1475996400, 
    1476000000, 1476003600, 1476007200, 1476010800, 1476014400, 1476018000, 
    1476021600, 1476025200, 1476028800, 1476032400, 1476036000, 1476039600, 
    1476043200, 1476046800, 1476050400, 1476054000, 1476057600, 1476061200, 
    1476064800, 1476068400, 1476072000, 1476075600, 1476079200, 1476082800, 
    1476086400, 1476090000, 1476093600, 1476097200, 1476100800, 1476104400, 
    1476108000, 1476111600, 1476115200, 1476118800, 1476122400, 1476126000, 
    1476129600, 1476133200, 1476136800, 1476140400, 1476144000, 1476147600, 
    1476151200, 1476154800, 1476158400, 1476162000, 1476165600, 1476169200, 
    1476172800, 1476176400, 1476180000, 1476183600, 1476187200, 1476190800, 
    1476194400, 1476198000, 1476201600, 1476205200, 1476208800, 1476212400, 
    1476216000, 1476219600, 1476223200, 1476226800, 1476230400, 1476234000, 
    1476237600, 1476241200, 1476244800, 1476248400, 1476252000, 1476255600, 
    1476259200, 1476262800, 1476266400, 1476270000, 1476273600, 1476277200, 
    1476280800, 1476284400, 1476288000, 1476291600, 1476295200, 1476298800, 
    1476302400, 1476306000, 1476309600, 1476313200, 1476316800, 1476320400, 
    1476324000, 1476327600, 1476331200, 1476334800, 1476338400, 1476342000, 
    1476345600, 1476349200, 1476352800, 1476356400, 1476360000, 1476363600, 
    1476367200, 1476370800, 1476374400, 1476378000, 1476381600, 1476385200, 
    1476388800, 1476392400, 1476396000, 1476399600, 1476403200, 1476406800, 
    1476410400, 1476414000, 1476417600, 1476421200, 1476424800, 1476428400, 
    1476432000, 1476435600, 1476439200, 1476442800, 1476446400, 1476450000, 
    1476453600, 1476457200, 1476460800, 1476464400, 1476468000, 1476471600, 
    1476475200, 1476478800, 1476482400, 1476486000, 1476489600, 1476493200, 
    1476496800, 1476500400, 1476504000, 1476507600, 1476511200, 1476514800, 
    1476518400, 1476522000, 1476525600, 1476529200, 1476532800, 1476536400, 
    1476540000, 1476543600, 1476547200, 1476550800, 1476554400, 1476558000, 
    1476561600, 1476565200, 1476568800, 1476572400, 1476576000, 1476579600, 
    1476583200, 1476586800, 1476590400, 1476594000, 1476597600, 1476601200, 
    1476604800, 1476608400, 1476612000, 1476615600, 1476619200, 1476622800, 
    1476626400, 1476630000, 1476633600, 1476637200, 1476640800, 1476644400, 
    1476648000, 1476651600, 1476655200, 1476658800, 1476662400, 1476666000, 
    1476669600, 1476673200, 1476676800, 1476680400, 1476684000, 1476687600, 
    1476691200, 1476694800, 1476698400, 1476702000, 1476705600, 1476709200, 
    1476712800, 1476716400, 1476720000, 1476723600, 1476727200, 1476730800, 
    1476734400, 1476738000, 1476741600, 1476745200, 1476748800, 1476752400, 
    1476756000, 1476759600, 1476763200, 1476766800, 1476770400, 1476774000, 
    1476777600, 1476781200, 1476784800, 1476788400, 1476792000, 1476795600, 
    1476799200, 1476802800, 1476806400, 1476810000, 1476813600, 1476817200, 
    1476820800, 1476824400, 1476828000, 1476831600, 1476835200, 1476838800, 
    1476842400, 1476846000, 1476849600, 1476853200, 1476856800, 1476860400, 
    1476864000, 1476867600, 1476871200, 1476874800, 1476878400, 1476882000, 
    1476885600, 1476889200, 1476892800, 1476896400, 1476900000, 1476903600, 
    1476907200, 1476910800, 1476914400, 1476918000, 1476921600, 1476925200, 
    1476928800, 1476932400, 1476936000, 1476939600, 1476943200, 1476946800, 
    1476950400, 1476954000, 1476957600, 1476961200, 1476964800, 1476968400, 
    1476972000, 1476975600, 1476979200, 1476982800, 1476986400, 1476990000, 
    1476993600, 1476997200, 1477000800, 1477004400, 1477008000, 1477011600, 
    1477015200, 1477018800, 1477022400, 1477026000, 1477029600, 1477033200, 
    1477036800, 1477040400, 1477044000, 1477047600, 1477051200, 1477054800, 
    1477058400, 1477062000, 1477065600, 1477069200, 1477072800, 1477076400, 
    1477080000, 1477083600, 1477087200, 1477090800, 1477094400, 1477098000, 
    1477101600, 1477105200, 1477108800, 1477112400, 1477116000, 1477119600, 
    1477123200, 1477126800, 1477130400, 1477134000, 1477137600, 1477141200, 
    1477144800, 1477148400, 1477152000, 1477155600, 1477159200, 1477162800, 
    1477166400, 1477170000, 1477173600, 1477177200, 1477180800, 1477184400, 
    1477188000, 1477191600, 1477195200, 1477198800, 1477202400, 1477206000, 
    1477209600, 1477213200, 1477216800, 1477220400, 1477224000, 1477227600, 
    1477231200, 1477234800, 1477238400, 1477242000, 1477245600, 1477249200, 
    1477252800, 1477256400, 1477260000, 1477263600, 1477267200, 1477270800, 
    1477274400, 1477278000, 1477281600, 1477285200, 1477288800, 1477292400, 
    1477296000, 1477299600, 1477303200, 1477306800, 1477310400, 1477314000, 
    1477317600, 1477321200, 1477324800, 1477328400, 1477332000, 1477335600, 
    1477339200, 1477342800, 1477346400, 1477350000, 1477353600, 1477357200, 
    1477360800, 1477364400, 1477368000, 1477371600, 1477375200, 1477378800, 
    1477382400, 1477386000, 1477389600, 1477393200, 1477396800, 1477400400, 
    1477404000, 1477407600, 1477411200, 1477414800, 1477418400, 1477422000, 
    1477425600, 1477429200, 1477432800, 1477436400, 1477440000, 1477443600, 
    1477447200, 1477450800, 1477454400, 1477458000, 1477461600, 1477465200, 
    1477468800, 1477472400, 1477476000, 1477479600, 1477483200, 1477486800, 
    1477490400, 1477494000, 1477497600, 1477501200, 1477504800, 1477508400, 
    1477512000, 1477515600, 1477519200, 1477522800, 1477526400, 1477530000, 
    1477533600, 1477537200, 1477540800, 1477544400, 1477548000, 1477551600, 
    1477555200, 1477558800, 1477562400, 1477566000, 1477569600, 1477573200, 
    1477576800, 1477580400, 1477584000, 1477587600, 1477591200, 1477594800, 
    1477598400, 1477602000, 1477605600, 1477609200, 1477612800, 1477616400, 
    1477620000, 1477623600, 1477627200, 1477630800, 1477634400, 1477638000, 
    1477641600, 1477645200, 1477648800, 1477652400, 1477656000, 1477659600, 
    1477663200, 1477666800, 1477670400, 1477674000, 1477677600, 1477681200, 
    1477684800, 1477688400, 1477692000, 1477695600, 1477699200, 1477702800, 
    1477706400, 1477710000, 1477713600, 1477717200, 1477720800, 1477724400, 
    1477728000, 1477731600, 1477735200, 1477738800, 1477742400, 1477746000, 
    1477749600, 1477753200, 1477756800, 1477760400, 1477764000, 1477767600, 
    1477771200, 1477774800, 1477778400, 1477782000, 1477785600, 1477789200, 
    1477792800, 1477796400, 1477800000, 1477803600, 1477807200, 1477810800, 
    1477814400, 1477818000, 1477821600, 1477825200, 1477828800, 1477832400, 
    1477836000, 1477839600, 1477843200, 1477846800, 1477850400, 1477854000, 
    1477857600, 1477861200, 1477864800, 1477868400, 1477872000, 1477875600, 
    1477879200, 1477882800, 1477886400, 1477890000, 1477893600, 1477897200, 
    1477900800, 1477904400, 1477908000, 1477911600, 1477915200, 1477918800, 
    1477922400, 1477926000, 1477929600, 1477933200, 1477936800, 1477940400, 
    1477944000, 1477947600, 1477951200, 1477954800, 1477958400, 1477962000, 
    1477965600, 1477969200, 1477972800, 1477976400, 1477980000, 1477983600, 
    1477987200, 1477990800, 1477994400, 1477998000, 1478001600, 1478005200, 
    1478008800, 1478012400, 1478016000, 1478019600, 1478023200, 1478026800, 
    1478030400, 1478034000, 1478037600, 1478041200, 1478044800, 1478048400, 
    1478052000, 1478055600, 1478059200, 1478062800, 1478066400, 1478070000, 
    1478073600, 1478077200, 1478080800, 1478084400, 1478088000, 1478091600, 
    1478095200, 1478098800, 1478102400, 1478106000, 1478109600, 1478113200, 
    1478116800, 1478120400, 1478124000, 1478127600, 1478131200, 1478134800, 
    1478138400, 1478142000, 1478145600, 1478149200, 1478152800, 1478156400, 
    1478160000, 1478163600, 1478167200, 1478170800, 1478174400, 1478178000, 
    1478181600, 1478185200, 1478188800, 1478192400, 1478196000, 1478199600, 
    1478203200, 1478206800, 1478210400, 1478214000, 1478217600, 1478221200, 
    1478224800, 1478228400, 1478232000, 1478235600, 1478239200, 1478242800, 
    1478246400, 1478250000, 1478253600, 1478257200, 1478260800, 1478264400, 
    1478268000, 1478271600, 1478275200, 1478278800, 1478282400, 1478286000, 
    1478289600, 1478293200, 1478296800, 1478300400, 1478304000, 1478307600, 
    1478311200, 1478314800, 1478318400, 1478322000, 1478325600, 1478329200, 
    1478332800, 1478336400, 1478340000, 1478343600, 1478347200, 1478350800, 
    1478354400, 1478358000, 1478361600, 1478365200, 1478368800, 1478372400, 
    1478376000, 1478379600, 1478383200, 1478386800, 1478390400, 1478394000, 
    1478397600, 1478401200, 1478404800, 1478408400, 1478412000, 1478415600, 
    1478419200, 1478422800, 1478426400, 1478430000, 1478433600, 1478437200, 
    1478440800, 1478444400, 1478448000, 1478451600, 1478455200, 1478458800, 
    1478462400, 1478466000, 1478469600, 1478473200, 1478476800, 1478480400, 
    1478484000, 1478487600, 1478491200, 1478494800, 1478498400, 1478502000, 
    1478505600, 1478509200, 1478512800, 1478516400, 1478520000, 1478523600, 
    1478527200, 1478530800, 1478534400, 1478538000, 1478541600, 1478545200, 
    1478548800, 1478552400, 1478556000, 1478559600, 1478563200, 1478566800, 
    1478570400, 1478574000, 1478577600, 1478581200, 1478584800, 1478588400, 
    1478592000, 1478595600, 1478599200, 1478602800, 1478606400, 1478610000, 
    1478613600, 1478617200, 1478620800, 1478624400, 1478628000, 1478631600, 
    1478635200, 1478638800, 1478642400, 1478646000, 1478649600, 1478653200, 
    1478656800, 1478660400, 1478664000, 1478667600, 1478671200, 1478674800, 
    1478678400, 1478682000, 1478685600, 1478689200, 1478692800, 1478696400, 
    1478700000, 1478703600, 1478707200, 1478710800, 1478714400, 1478718000, 
    1478721600, 1478725200, 1478728800, 1478732400, 1478736000, 1478739600, 
    1478743200, 1478746800, 1478750400, 1478754000, 1478757600, 1478761200, 
    1478764800, 1478768400, 1478772000, 1478775600, 1478779200, 1478782800, 
    1478786400, 1478790000, 1478793600, 1478797200, 1478800800, 1478804400, 
    1478808000, 1478811600, 1478815200, 1478818800, 1478822400, 1478826000, 
    1478829600, 1478833200, 1478836800, 1478840400, 1478844000, 1478847600, 
    1478851200, 1478854800, 1478858400, 1478862000, 1478865600, 1478869200, 
    1478872800, 1478876400, 1478880000, 1478883600, 1478887200, 1478890800, 
    1478894400, 1478898000, 1478901600, 1478905200, 1478908800, 1478912400, 
    1478916000, 1478919600, 1478923200, 1478926800, 1478930400, 1478934000, 
    1478937600, 1478941200, 1478944800, 1478948400, 1478952000, 1478955600, 
    1478959200, 1478962800, 1478966400, 1478970000, 1478973600, 1478977200, 
    1478980800, 1478984400, 1478988000, 1478991600, 1478995200, 1478998800, 
    1479002400, 1479006000, 1479009600, 1479013200, 1479016800, 1479020400, 
    1479024000, 1479027600, 1479031200, 1479034800, 1479038400, 1479042000, 
    1479045600, 1479049200, 1479052800, 1479056400, 1479060000, 1479063600, 
    1479067200, 1479070800, 1479074400, 1479078000, 1479081600, 1479085200, 
    1479088800, 1479092400, 1479096000, 1479099600, 1479103200, 1479106800, 
    1479110400, 1479114000, 1479117600, 1479121200, 1479124800, 1479128400, 
    1479132000, 1479135600, 1479139200, 1479142800, 1479146400, 1479150000, 
    1479153600, 1479157200, 1479160800, 1479164400, 1479168000, 1479171600, 
    1479175200, 1479178800, 1479182400, 1479186000, 1479189600, 1479193200, 
    1479196800, 1479200400, 1479204000, 1479207600, 1479211200, 1479214800, 
    1479218400, 1479222000, 1479225600, 1479229200, 1479232800, 1479236400, 
    1479240000, 1479243600, 1479247200, 1479250800, 1479254400, 1479258000, 
    1479261600, 1479265200, 1479268800, 1479272400, 1479276000, 1479279600, 
    1479283200, 1479286800, 1479290400, 1479294000, 1479297600, 1479301200, 
    1479304800, 1479308400, 1479312000, 1479315600, 1479319200, 1479322800, 
    1479326400, 1479330000, 1479333600, 1479337200, 1479340800, 1479344400, 
    1479348000, 1479351600, 1479355200, 1479358800, 1479362400, 1479366000, 
    1479369600, 1479373200, 1479376800, 1479380400, 1479384000, 1479387600, 
    1479391200, 1479394800, 1479398400, 1479402000, 1479405600, 1479409200, 
    1479412800, 1479416400, 1479420000, 1479423600, 1479427200, 1479430800, 
    1479434400, 1479438000, 1479441600, 1479445200, 1479448800, 1479452400, 
    1479456000, 1479459600, 1479463200, 1479466800, 1479470400, 1479474000, 
    1479477600, 1479481200, 1479484800, 1479488400, 1479492000, 1479495600, 
    1479499200, 1479502800, 1479506400, 1479510000, 1479513600, 1479517200, 
    1479520800, 1479524400, 1479528000, 1479531600, 1479535200, 1479538800, 
    1479542400, 1479546000, 1479549600, 1479553200, 1479556800, 1479560400, 
    1479564000, 1479567600, 1479571200, 1479574800, 1479578400, 1479582000, 
    1479585600, 1479589200, 1479592800, 1479596400, 1479600000, 1479603600, 
    1479607200, 1479610800, 1479614400, 1479618000, 1479621600, 1479625200, 
    1479628800, 1479632400, 1479636000, 1479639600, 1479643200, 1479646800, 
    1479650400, 1479654000, 1479657600, 1479661200, 1479664800, 1479668400, 
    1479672000, 1479675600, 1479679200, 1479682800, 1479686400, 1479690000, 
    1479693600, 1479697200, 1479700800, 1479704400, 1479708000, 1479711600, 
    1479715200, 1479718800, 1479722400, 1479726000, 1479729600, 1479733200, 
    1479736800, 1479740400, 1479744000, 1479747600, 1479751200, 1479754800, 
    1479758400, 1479762000, 1479765600, 1479769200, 1479772800, 1479776400, 
    1479780000, 1479783600, 1479787200, 1479790800, 1479794400, 1479798000, 
    1479801600, 1479805200, 1479808800, 1479812400, 1479816000, 1479819600, 
    1479823200, 1479826800, 1479830400, 1479834000, 1479837600, 1479841200, 
    1479844800, 1479848400, 1479852000, 1479855600, 1479859200, 1479862800, 
    1479866400, 1479870000, 1479873600, 1479877200, 1479880800, 1479884400, 
    1479888000, 1479891600, 1479895200, 1479898800, 1479902400, 1479906000, 
    1479909600, 1479913200, 1479916800, 1479920400, 1479924000, 1479927600, 
    1479931200, 1479934800, 1479938400, 1479942000, 1479945600, 1479949200, 
    1479952800, 1479956400, 1479960000, 1479963600, 1479967200, 1479970800, 
    1479974400, 1479978000, 1479981600, 1479985200, 1479988800, 1479992400, 
    1479996000, 1479999600, 1480003200, 1480006800, 1480010400, 1480014000, 
    1480017600, 1480021200, 1480024800, 1480028400, 1480032000, 1480035600, 
    1480039200, 1480042800, 1480046400, 1480050000, 1480053600, 1480057200, 
    1480060800, 1480064400, 1480068000, 1480071600, 1480075200, 1480078800, 
    1480082400, 1480086000, 1480089600, 1480093200, 1480096800, 1480100400, 
    1480104000, 1480107600, 1480111200, 1480114800, 1480118400, 1480122000, 
    1480125600, 1480129200, 1480132800, 1480136400, 1480140000, 1480143600, 
    1480147200, 1480150800, 1480154400, 1480158000, 1480161600, 1480165200, 
    1480168800, 1480172400, 1480176000, 1480179600, 1480183200, 1480186800, 
    1480190400, 1480194000, 1480197600, 1480201200, 1480204800, 1480208400, 
    1480212000, 1480215600, 1480219200, 1480222800, 1480226400, 1480230000, 
    1480233600, 1480237200, 1480240800, 1480244400, 1480248000, 1480251600, 
    1480255200, 1480258800, 1480262400, 1480266000, 1480269600, 1480273200, 
    1480276800, 1480280400, 1480284000, 1480287600, 1480291200, 1480294800, 
    1480298400, 1480302000, 1480305600, 1480309200, 1480312800, 1480316400, 
    1480320000, 1480323600, 1480327200, 1480330800, 1480334400, 1480338000, 
    1480341600, 1480345200, 1480348800, 1480352400, 1480356000, 1480359600, 
    1480363200, 1480366800, 1480370400, 1480374000, 1480377600, 1480381200, 
    1480384800, 1480388400, 1480392000, 1480395600, 1480399200, 1480402800, 
    1480406400, 1480410000, 1480413600, 1480417200, 1480420800, 1480424400, 
    1480428000, 1480431600, 1480435200, 1480438800, 1480442400, 1480446000, 
    1480449600, 1480453200, 1480456800, 1480460400, 1480464000, 1480467600, 
    1480471200, 1480474800, 1480478400, 1480482000, 1480485600, 1480489200, 
    1480492800, 1480496400, 1480500000, 1480503600, 1480507200, 1480510800, 
    1480514400, 1480518000, 1480521600, 1480525200, 1480528800, 1480532400, 
    1480536000, 1480539600, 1480543200, 1480546800, 1480550400, 1480554000, 
    1480557600, 1480561200, 1480564800, 1480568400, 1480572000, 1480575600, 
    1480579200, 1480582800, 1480586400, 1480590000, 1480593600, 1480597200, 
    1480600800, 1480604400, 1480608000, 1480611600, 1480615200, 1480618800, 
    1480622400, 1480626000, 1480629600, 1480633200, 1480636800, 1480640400, 
    1480644000, 1480647600, 1480651200, 1480654800, 1480658400, 1480662000, 
    1480665600, 1480669200, 1480672800, 1480676400, 1480680000, 1480683600, 
    1480687200, 1480690800, 1480694400, 1480698000, 1480701600, 1480705200, 
    1480708800, 1480712400, 1480716000, 1480719600, 1480723200, 1480726800, 
    1480730400, 1480734000, 1480737600, 1480741200, 1480744800, 1480748400, 
    1480752000, 1480755600, 1480759200, 1480762800, 1480766400, 1480770000, 
    1480773600, 1480777200, 1480780800, 1480784400, 1480788000, 1480791600, 
    1480795200, 1480798800, 1480802400, 1480806000, 1480809600, 1480813200, 
    1480816800, 1480820400, 1480824000, 1480827600, 1480831200, 1480834800, 
    1480838400, 1480842000, 1480845600, 1480849200, 1480852800, 1480856400, 
    1480860000, 1480863600, 1480867200, 1480870800, 1480874400, 1480878000, 
    1480881600, 1480885200, 1480888800, 1480892400, 1480896000, 1480899600, 
    1480903200, 1480906800, 1480910400, 1480914000, 1480917600, 1480921200, 
    1480924800, 1480928400, 1480932000, 1480935600, 1480939200, 1480942800, 
    1480946400, 1480950000, 1480953600, 1480957200, 1480960800, 1480964400, 
    1480968000, 1480971600, 1480975200, 1480978800, 1480982400, 1480986000, 
    1480989600, 1480993200, 1480996800, 1481000400, 1481004000, 1481007600, 
    1481011200, 1481014800, 1481018400, 1481022000, 1481025600, 1481029200, 
    1481032800, 1481036400, 1481040000, 1481043600, 1481047200, 1481050800, 
    1481054400, 1481058000, 1481061600, 1481065200, 1481068800, 1481072400, 
    1481076000, 1481079600, 1481083200, 1481086800, 1481090400, 1481094000, 
    1481097600, 1481101200, 1481104800, 1481108400, 1481112000, 1481115600, 
    1481119200, 1481122800, 1481126400, 1481130000, 1481133600, 1481137200, 
    1481140800, 1481144400, 1481148000, 1481151600, 1481155200, 1481158800, 
    1481162400, 1481166000, 1481169600, 1481173200, 1481176800, 1481180400, 
    1481184000, 1481187600, 1481191200, 1481194800, 1481198400, 1481202000, 
    1481205600, 1481209200, 1481212800, 1481216400, 1481220000, 1481223600, 
    1481227200, 1481230800, 1481234400, 1481238000, 1481241600, 1481245200, 
    1481248800, 1481252400, 1481256000, 1481259600, 1481263200, 1481266800, 
    1481270400, 1481274000, 1481277600, 1481281200, 1481284800, 1481288400, 
    1481292000, 1481295600, 1481299200, 1481302800, 1481306400, 1481310000, 
    1481313600, 1481317200, 1481320800, 1481324400, 1481328000, 1481331600, 
    1481335200, 1481338800, 1481342400, 1481346000, 1481349600, 1481353200, 
    1481356800, 1481360400, 1481364000, 1481367600, 1481371200, 1481374800, 
    1481378400, 1481382000, 1481385600, 1481389200, 1481392800, 1481396400, 
    1481400000, 1481403600, 1481407200, 1481410800, 1481414400, 1481418000, 
    1481421600, 1481425200, 1481428800, 1481432400, 1481436000, 1481439600, 
    1481443200, 1481446800, 1481450400, 1481454000, 1481457600, 1481461200, 
    1481464800, 1481468400, 1481472000, 1481475600, 1481479200, 1481482800, 
    1481486400, 1481490000, 1481493600, 1481497200, 1481500800, 1481504400, 
    1481508000, 1481511600, 1481515200, 1481518800, 1481522400, 1481526000, 
    1481529600, 1481533200, 1481536800, 1481540400, 1481544000, 1481547600, 
    1481551200, 1481554800, 1481558400, 1481562000, 1481565600, 1481569200, 
    1481572800, 1481576400, 1481580000, 1481583600, 1481587200, 1481590800, 
    1481594400, 1481598000, 1481601600, 1481605200, 1481608800, 1481612400, 
    1481616000, 1481619600, 1481623200, 1481626800, 1481630400, 1481634000, 
    1481637600, 1481641200, 1481644800, 1481648400, 1481652000, 1481655600, 
    1481659200, 1481662800, 1481666400, 1481670000, 1481673600, 1481677200, 
    1481680800, 1481684400, 1481688000, 1481691600, 1481695200, 1481698800, 
    1481702400, 1481706000, 1481709600, 1481713200, 1481716800, 1481720400, 
    1481724000, 1481727600, 1481731200, 1481734800, 1481738400, 1481742000, 
    1481745600, 1481749200, 1481752800, 1481756400, 1481760000, 1481763600, 
    1481767200, 1481770800, 1481774400, 1481778000, 1481781600, 1481785200, 
    1481788800, 1481792400, 1481796000, 1481799600, 1481803200, 1481806800, 
    1481810400, 1481814000, 1481817600, 1481821200, 1481824800, 1481828400, 
    1481832000, 1481835600, 1481839200, 1481842800, 1481846400, 1481850000, 
    1481853600, 1481857200, 1481860800, 1481864400, 1481868000, 1481871600, 
    1481875200, 1481878800, 1481882400, 1481886000, 1481889600, 1481893200, 
    1481896800, 1481900400, 1481904000, 1481907600, 1481911200, 1481914800, 
    1481918400, 1481922000, 1481925600, 1481929200, 1481932800, 1481936400, 
    1481940000, 1481943600, 1481947200, 1481950800, 1481954400, 1481958000, 
    1481961600, 1481965200, 1481968800, 1481972400, 1481976000, 1481979600, 
    1481983200, 1481986800, 1481990400, 1481994000, 1481997600, 1482001200, 
    1482004800, 1482008400, 1482012000, 1482015600, 1482019200, 1482022800, 
    1482026400, 1482030000, 1482033600, 1482037200, 1482040800, 1482044400, 
    1482048000, 1482051600, 1482055200, 1482058800, 1482062400, 1482066000, 
    1482069600, 1482073200, 1482076800, 1482080400, 1482084000, 1482087600, 
    1482091200, 1482094800, 1482098400, 1482102000, 1482105600, 1482109200, 
    1482112800, 1482116400, 1482120000, 1482123600, 1482127200, 1482130800, 
    1482134400, 1482138000, 1482141600, 1482145200, 1482148800, 1482152400, 
    1482156000, 1482159600, 1482163200, 1482166800, 1482170400, 1482174000, 
    1482177600, 1482181200, 1482184800, 1482188400, 1482192000, 1482195600, 
    1482199200, 1482202800, 1482206400, 1482210000, 1482213600, 1482217200, 
    1482220800, 1482224400, 1482228000, 1482231600, 1482235200, 1482238800, 
    1482242400, 1482246000, 1482249600, 1482253200, 1482256800, 1482260400, 
    1482264000, 1482267600, 1482271200, 1482274800, 1482278400, 1482282000, 
    1482285600, 1482289200, 1482292800, 1482296400, 1482300000, 1482303600, 
    1482307200, 1482310800, 1482314400, 1482318000, 1482321600, 1482325200, 
    1482328800, 1482332400, 1482336000, 1482339600, 1482343200, 1482346800, 
    1482350400, 1482354000, 1482357600, 1482361200, 1482364800, 1482368400, 
    1482372000, 1482375600, 1482379200, 1482382800, 1482386400, 1482390000, 
    1482393600, 1482397200, 1482400800, 1482404400, 1482408000, 1482411600, 
    1482415200, 1482418800, 1482422400, 1482426000, 1482429600, 1482433200, 
    1482436800, 1482440400, 1482444000, 1482447600, 1482451200, 1482454800, 
    1482458400, 1482462000, 1482465600, 1482469200, 1482472800, 1482476400, 
    1482480000, 1482483600, 1482487200, 1482490800, 1482494400, 1482498000, 
    1482501600, 1482505200, 1482508800, 1482512400, 1482516000, 1482519600, 
    1482523200, 1482526800, 1482530400, 1482534000, 1482537600, 1482541200, 
    1482544800, 1482548400, 1482552000, 1482555600, 1482559200, 1482562800, 
    1482566400, 1482570000, 1482573600, 1482577200, 1482580800, 1482584400, 
    1482588000, 1482591600, 1482595200, 1482598800, 1482602400, 1482606000, 
    1482609600, 1482613200, 1482616800, 1482620400, 1482624000, 1482627600, 
    1482631200, 1482634800, 1482638400, 1482642000, 1482645600, 1482649200, 
    1482652800, 1482656400, 1482660000, 1482663600, 1482667200, 1482670800, 
    1482674400, 1482678000, 1482681600, 1482685200, 1482688800, 1482692400, 
    1482696000, 1482699600, 1482703200, 1482706800, 1482710400, 1482714000, 
    1482717600, 1482721200, 1482724800, 1482728400, 1482732000, 1482735600, 
    1482739200, 1482742800, 1482746400, 1482750000, 1482753600, 1482757200, 
    1482760800, 1482764400, 1482768000, 1482771600, 1482775200, 1482778800, 
    1482782400, 1482786000, 1482789600, 1482793200, 1482796800, 1482800400, 
    1482804000, 1482807600, 1482811200, 1482814800, 1482818400, 1482822000, 
    1482825600, 1482829200, 1482832800, 1482836400, 1482840000, 1482843600, 
    1482847200, 1482850800, 1482854400, 1482858000, 1482861600, 1482865200, 
    1482868800, 1482872400, 1482876000, 1482879600, 1482883200, 1482886800, 
    1482890400, 1482894000, 1482897600, 1482901200, 1482904800, 1482908400, 
    1482912000, 1482915600, 1482919200, 1482922800, 1482926400, 1482930000, 
    1482933600, 1482937200, 1482940800, 1482944400, 1482948000, 1482951600, 
    1482955200, 1482958800, 1482962400, 1482966000, 1482969600, 1482973200, 
    1482976800, 1482980400, 1482984000, 1482987600, 1482991200, 1482994800, 
    1482998400, 1483002000, 1483005600, 1483009200, 1483012800, 1483016400, 
    1483020000, 1483023600, 1483027200, 1483030800, 1483034400, 1483038000, 
    1483041600, 1483045200, 1483048800, 1483052400, 1483056000, 1483059600, 
    1483063200, 1483066800, 1483070400, 1483074000, 1483077600, 1483081200, 
    1483084800, 1483088400, 1483092000, 1483095600, 1483099200, 1483102800, 
    1483106400, 1483110000, 1483113600, 1483117200, 1483120800, 1483124400, 
    1483128000, 1483131600, 1483135200, 1483138800, 1483142400, 1483146000, 
    1483149600, 1483153200, 1483156800, 1483160400, 1483164000, 1483167600, 
    1483171200, 1483174800, 1483178400, 1483182000, 1483185600, 1483189200, 
    1483192800, 1483196400, 1483200000, 1483203600, 1483207200, 1483210800, 
    1483214400, 1483218000, 1483221600, 1483225200, 1483228800, 1483232400, 
    1483236000, 1483239600, 1483243200, 1483246800, 1483250400, 1483254000, 
    1483257600, 1483261200, 1483264800, 1483268400, 1483272000, 1483275600, 
    1483279200, 1483282800, 1483286400, 1483290000, 1483293600, 1483297200, 
    1483300800, 1483304400, 1483308000, 1483311600, 1483315200, 1483318800, 
    1483322400, 1483326000, 1483329600, 1483333200, 1483336800, 1483340400, 
    1483344000, 1483347600, 1483351200, 1483354800, 1483358400, 1483362000, 
    1483365600, 1483369200, 1483372800, 1483376400, 1483380000, 1483383600, 
    1483387200, 1483390800, 1483394400, 1483398000, 1483401600, 1483405200, 
    1483408800, 1483412400, 1483416000, 1483419600, 1483423200, 1483426800, 
    1483430400, 1483434000, 1483437600, 1483441200, 1483444800, 1483448400, 
    1483452000, 1483455600, 1483459200, 1483462800, 1483466400, 1483470000, 
    1483473600, 1483477200, 1483480800, 1483484400, 1483488000, 1483491600, 
    1483495200, 1483498800, 1483502400, 1483506000, 1483509600, 1483513200, 
    1483516800, 1483520400, 1483524000, 1483527600, 1483531200, 1483534800, 
    1483538400, 1483542000, 1483545600, 1483549200, 1483552800, 1483556400, 
    1483560000, 1483563600, 1483567200, 1483570800, 1483574400, 1483578000, 
    1483581600, 1483585200, 1483588800, 1483592400, 1483596000, 1483599600, 
    1483603200, 1483606800, 1483610400, 1483614000, 1483617600, 1483621200, 
    1483624800, 1483628400, 1483632000, 1483635600, 1483639200, 1483642800, 
    1483646400, 1483650000, 1483653600, 1483657200, 1483660800, 1483664400, 
    1483668000, 1483671600, 1483675200, 1483678800, 1483682400, 1483686000, 
    1483689600, 1483693200, 1483696800, 1483700400, 1483704000, 1483707600, 
    1483711200, 1483714800, 1483718400, 1483722000, 1483725600, 1483729200, 
    1483732800, 1483736400, 1483740000, 1483743600, 1483747200, 1483750800, 
    1483754400, 1483758000, 1483761600, 1483765200, 1483768800, 1483772400, 
    1483776000, 1483779600, 1483783200, 1483786800, 1483790400, 1483794000, 
    1483797600, 1483801200, 1483804800, 1483808400, 1483812000, 1483815600, 
    1483819200, 1483822800, 1483826400, 1483830000, 1483833600, 1483837200, 
    1483840800, 1483844400, 1483848000, 1483851600, 1483855200, 1483858800, 
    1483862400, 1483866000, 1483869600, 1483873200, 1483876800, 1483880400, 
    1483884000, 1483887600, 1483891200, 1483894800, 1483898400, 1483902000, 
    1483905600, 1483909200, 1483912800, 1483916400, 1483920000, 1483923600, 
    1483927200, 1483930800, 1483934400, 1483938000, 1483941600, 1483945200, 
    1483948800, 1483952400, 1483956000, 1483959600, 1483963200, 1483966800, 
    1483970400, 1483974000, 1483977600, 1483981200, 1483984800, 1483988400, 
    1483992000, 1483995600, 1483999200, 1484002800, 1484006400, 1484010000, 
    1484013600, 1484017200, 1484020800, 1484024400, 1484028000, 1484031600, 
    1484035200, 1484038800, 1484042400, 1484046000, 1484049600, 1484053200, 
    1484056800, 1484060400, 1484064000, 1484067600, 1484071200, 1484074800, 
    1484078400, 1484082000, 1484085600, 1484089200, 1484092800, 1484096400, 
    1484100000, 1484103600, 1484107200, 1484110800, 1484114400, 1484118000, 
    1484121600, 1484125200, 1484128800, 1484132400, 1484136000, 1484139600, 
    1484143200, 1484146800, 1484150400, 1484154000, 1484157600, 1484161200, 
    1484164800, 1484168400, 1484172000, 1484175600, 1484179200, 1484182800, 
    1484186400, 1484190000, 1484193600, 1484197200, 1484200800, 1484204400, 
    1484208000, 1484211600, 1484215200, 1484218800, 1484222400, 1484226000, 
    1484229600, 1484233200, 1484236800, 1484240400, 1484244000, 1484247600, 
    1484251200, 1484254800, 1484258400, 1484262000, 1484265600, 1484269200, 
    1484272800, 1484276400, 1484280000, 1484283600, 1484287200, 1484290800, 
    1484294400, 1484298000, 1484301600, 1484305200, 1484308800, 1484312400, 
    1484316000, 1484319600, 1484323200, 1484326800, 1484330400, 1484334000, 
    1484337600, 1484341200, 1484344800, 1484348400, 1484352000, 1484355600, 
    1484359200, 1484362800, 1484366400, 1484370000, 1484373600, 1484377200, 
    1484380800, 1484384400, 1484388000, 1484391600, 1484395200, 1484398800, 
    1484402400, 1484406000, 1484409600, 1484413200, 1484416800, 1484420400, 
    1484424000, 1484427600, 1484431200, 1484434800, 1484438400, 1484442000, 
    1484445600, 1484449200, 1484452800, 1484456400, 1484460000, 1484463600, 
    1484467200, 1484470800, 1484474400, 1484478000, 1484481600, 1484485200, 
    1484488800, 1484492400, 1484496000, 1484499600, 1484503200, 1484506800, 
    1484510400, 1484514000, 1484517600, 1484521200, 1484524800, 1484528400, 
    1484532000, 1484535600, 1484539200, 1484542800, 1484546400, 1484550000, 
    1484553600, 1484557200, 1484560800, 1484564400, 1484568000, 1484571600, 
    1484575200, 1484578800, 1484582400, 1484586000, 1484589600, 1484593200, 
    1484596800, 1484600400, 1484604000, 1484607600, 1484611200, 1484614800, 
    1484618400, 1484622000, 1484625600, 1484629200, 1484632800, 1484636400, 
    1484640000, 1484643600, 1484647200, 1484650800, 1484654400, 1484658000, 
    1484661600, 1484665200, 1484668800, 1484672400, 1484676000, 1484679600, 
    1484683200, 1484686800, 1484690400, 1484694000, 1484697600, 1484701200, 
    1484704800, 1484708400, 1484712000, 1484715600, 1484719200, 1484722800, 
    1484726400, 1484730000, 1484733600, 1484737200, 1484740800, 1484744400, 
    1484748000, 1484751600, 1484755200, 1484758800, 1484762400, 1484766000, 
    1484769600, 1484773200, 1484776800, 1484780400, 1484784000, 1484787600, 
    1484791200, 1484794800, 1484798400, 1484802000, 1484805600, 1484809200, 
    1484812800, 1484816400, 1484820000, 1484823600, 1484827200, 1484830800, 
    1484834400, 1484838000, 1484841600, 1484845200, 1484848800, 1484852400, 
    1484856000, 1484859600, 1484863200, 1484866800, 1484870400, 1484874000, 
    1484877600, 1484881200, 1484884800, 1484888400, 1484892000, 1484895600, 
    1484899200, 1484902800, 1484906400, 1484910000, 1484913600, 1484917200, 
    1484920800, 1484924400, 1484928000, 1484931600, 1484935200, 1484938800, 
    1484942400, 1484946000, 1484949600, 1484953200, 1484956800, 1484960400, 
    1484964000, 1484967600, 1484971200, 1484974800, 1484978400, 1484982000, 
    1484985600, 1484989200, 1484992800, 1484996400, 1485000000, 1485003600, 
    1485007200, 1485010800, 1485014400, 1485018000, 1485021600, 1485025200, 
    1485028800, 1485032400, 1485036000, 1485039600, 1485043200, 1485046800, 
    1485050400, 1485054000, 1485057600, 1485061200, 1485064800, 1485068400, 
    1485072000, 1485075600, 1485079200, 1485082800, 1485086400, 1485090000, 
    1485093600, 1485097200, 1485100800, 1485104400, 1485108000, 1485111600, 
    1485115200, 1485118800, 1485122400, 1485126000, 1485129600, 1485133200, 
    1485136800, 1485140400, 1485144000, 1485147600, 1485151200, 1485154800, 
    1485158400, 1485162000, 1485165600, 1485169200, 1485172800, 1485176400, 
    1485180000, 1485183600, 1485187200, 1485190800, 1485194400, 1485198000, 
    1485201600, 1485205200, 1485208800, 1485212400, 1485216000, 1485219600, 
    1485223200, 1485226800, 1485230400, 1485234000, 1485237600, 1485241200, 
    1485244800, 1485248400, 1485252000, 1485255600, 1485259200, 1485262800, 
    1485266400, 1485270000, 1485273600, 1485277200, 1485280800, 1485284400, 
    1485288000, 1485291600, 1485295200, 1485298800, 1485302400, 1485306000, 
    1485309600, 1485313200, 1485316800, 1485320400, 1485324000, 1485327600, 
    1485331200, 1485334800, 1485338400, 1485342000, 1485345600, 1485349200, 
    1485352800, 1485356400, 1485360000, 1485363600, 1485367200, 1485370800, 
    1485374400, 1485378000, 1485381600, 1485385200, 1485388800, 1485392400, 
    1485396000, 1485399600, 1485403200, 1485406800, 1485410400, 1485414000, 
    1485417600, 1485421200, 1485424800, 1485428400, 1485432000, 1485435600, 
    1485439200, 1485442800, 1485446400, 1485450000, 1485453600, 1485457200, 
    1485460800, 1485464400, 1485468000, 1485471600, 1485475200, 1485478800, 
    1485482400, 1485486000, 1485489600, 1485493200, 1485496800, 1485500400, 
    1485504000, 1485507600, 1485511200, 1485514800, 1485518400, 1485522000, 
    1485525600, 1485529200, 1485532800, 1485536400, 1485540000, 1485543600, 
    1485547200, 1485550800, 1485554400, 1485558000, 1485561600, 1485565200, 
    1485568800, 1485572400, 1485576000, 1485579600, 1485583200, 1485586800, 
    1485590400, 1485594000, 1485597600, 1485601200, 1485604800, 1485608400, 
    1485612000, 1485615600, 1485619200, 1485622800, 1485626400, 1485630000, 
    1485633600, 1485637200, 1485640800, 1485644400, 1485648000, 1485651600, 
    1485655200, 1485658800, 1485662400, 1485666000, 1485669600, 1485673200, 
    1485676800, 1485680400, 1485684000, 1485687600, 1485691200, 1485694800, 
    1485698400, 1485702000, 1485705600, 1485709200, 1485712800, 1485716400, 
    1485720000, 1485723600, 1485727200, 1485730800, 1485734400, 1485738000, 
    1485741600, 1485745200, 1485748800, 1485752400, 1485756000, 1485759600, 
    1485763200, 1485766800, 1485770400, 1485774000, 1485777600, 1485781200, 
    1485784800, 1485788400, 1485792000, 1485795600, 1485799200, 1485802800, 
    1485806400, 1485810000, 1485813600, 1485817200, 1485820800, 1485824400, 
    1485828000, 1485831600, 1485835200, 1485838800, 1485842400, 1485846000, 
    1485849600, 1485853200, 1485856800, 1485860400, 1485864000, 1485867600, 
    1485871200, 1485874800, 1485878400, 1485882000, 1485885600, 1485889200, 
    1485892800, 1485896400, 1485900000, 1485903600, 1485907200, 1485910800, 
    1485914400, 1485918000, 1485921600, 1485925200, 1485928800, 1485932400, 
    1485936000, 1485939600, 1485943200, 1485946800, 1485950400, 1485954000, 
    1485957600, 1485961200, 1485964800, 1485968400, 1485972000, 1485975600, 
    1485979200, 1485982800, 1485986400, 1485990000, 1485993600, 1485997200, 
    1486000800, 1486004400, 1486008000, 1486011600, 1486015200, 1486018800, 
    1486022400, 1486026000, 1486029600, 1486033200, 1486036800, 1486040400, 
    1486044000, 1486047600, 1486051200, 1486054800, 1486058400, 1486062000, 
    1486065600, 1486069200, 1486072800, 1486076400, 1486080000, 1486083600, 
    1486087200, 1486090800, 1486094400, 1486098000, 1486101600, 1486105200, 
    1486108800, 1486112400, 1486116000, 1486119600, 1486123200, 1486126800, 
    1486130400, 1486134000, 1486137600, 1486141200, 1486144800, 1486148400, 
    1486152000, 1486155600, 1486159200, 1486162800, 1486166400, 1486170000, 
    1486173600, 1486177200, 1486180800, 1486184400, 1486188000, 1486191600, 
    1486195200, 1486198800, 1486202400, 1486206000, 1486209600, 1486213200, 
    1486216800, 1486220400, 1486224000, 1486227600, 1486231200, 1486234800, 
    1486238400, 1486242000, 1486245600, 1486249200, 1486252800, 1486256400, 
    1486260000, 1486263600, 1486267200, 1486270800, 1486274400, 1486278000, 
    1486281600, 1486285200, 1486288800, 1486292400, 1486296000, 1486299600, 
    1486303200, 1486306800, 1486310400, 1486314000, 1486317600, 1486321200, 
    1486324800, 1486328400, 1486332000, 1486335600, 1486339200, 1486342800, 
    1486346400, 1486350000, 1486353600, 1486357200, 1486360800, 1486364400, 
    1486368000, 1486371600, 1486375200, 1486378800, 1486382400, 1486386000, 
    1486389600, 1486393200, 1486396800, 1486400400, 1486404000, 1486407600, 
    1486411200, 1486414800, 1486418400, 1486422000, 1486425600, 1486429200, 
    1486432800, 1486436400, 1486440000, 1486443600, 1486447200, 1486450800, 
    1486454400, 1486458000, 1486461600, 1486465200, 1486468800, 1486472400, 
    1486476000, 1486479600, 1486483200, 1486486800, 1486490400, 1486494000, 
    1486497600, 1486501200, 1486504800, 1486508400, 1486512000, 1486515600, 
    1486519200, 1486522800, 1486526400, 1486530000, 1486533600, 1486537200, 
    1486540800, 1486544400, 1486548000, 1486551600, 1486555200, 1486558800, 
    1486562400, 1486566000, 1486569600, 1486573200, 1486576800, 1486580400, 
    1486584000, 1486587600, 1486591200, 1486594800, 1486598400, 1486602000, 
    1486605600, 1486609200, 1486612800, 1486616400, 1486620000, 1486623600, 
    1486627200, 1486630800, 1486634400, 1486638000, 1486641600, 1486645200, 
    1486648800, 1486652400, 1486656000, 1486659600, 1486663200, 1486666800, 
    1486670400, 1486674000, 1486677600, 1486681200, 1486684800, 1486688400, 
    1486692000, 1486695600, 1486699200, 1486702800, 1486706400, 1486710000, 
    1486713600, 1486717200, 1486720800, 1486724400, 1486728000, 1486731600, 
    1486735200, 1486738800, 1486742400, 1486746000, 1486749600, 1486753200, 
    1486756800, 1486760400, 1486764000, 1486767600, 1486771200, 1486774800, 
    1486778400, 1486782000, 1486785600, 1486789200, 1486792800, 1486796400, 
    1486800000, 1486803600, 1486807200, 1486810800, 1486814400, 1486818000, 
    1486821600, 1486825200, 1486828800, 1486832400, 1486836000, 1486839600, 
    1486843200, 1486846800, 1486850400, 1486854000, 1486857600, 1486861200, 
    1486864800, 1486868400, 1486872000, 1486875600, 1486879200, 1486882800, 
    1486886400, 1486890000, 1486893600, 1486897200, 1486900800, 1486904400, 
    1486908000, 1486911600, 1486915200, 1486918800, 1486922400, 1486926000, 
    1486929600, 1486933200, 1486936800, 1486940400, 1486944000, 1486947600, 
    1486951200, 1486954800, 1486958400, 1486962000, 1486965600, 1486969200, 
    1486972800, 1486976400, 1486980000, 1486983600, 1486987200, 1486990800, 
    1486994400, 1486998000, 1487001600, 1487005200, 1487008800, 1487012400, 
    1487016000, 1487019600, 1487023200, 1487026800, 1487030400, 1487034000, 
    1487037600, 1487041200, 1487044800, 1487048400, 1487052000, 1487055600, 
    1487059200, 1487062800, 1487066400, 1487070000, 1487073600, 1487077200, 
    1487080800, 1487084400, 1487088000, 1487091600, 1487095200, 1487098800, 
    1487102400, 1487106000, 1487109600, 1487113200, 1487116800, 1487120400, 
    1487124000, 1487127600, 1487131200, 1487134800, 1487138400, 1487142000, 
    1487145600, 1487149200, 1487152800, 1487156400, 1487160000, 1487163600, 
    1487167200, 1487170800, 1487174400, 1487178000, 1487181600, 1487185200, 
    1487188800, 1487192400, 1487196000, 1487199600, 1487203200, 1487206800, 
    1487210400, 1487214000, 1487217600, 1487221200, 1487224800, 1487228400, 
    1487232000, 1487235600, 1487239200, 1487242800, 1487246400, 1487250000, 
    1487253600, 1487257200, 1487260800, 1487264400, 1487268000, 1487271600, 
    1487275200, 1487278800, 1487282400, 1487286000, 1487289600, 1487293200, 
    1487296800, 1487300400, 1487304000, 1487307600, 1487311200, 1487314800, 
    1487318400, 1487322000, 1487325600, 1487329200, 1487332800, 1487336400, 
    1487340000, 1487343600, 1487347200, 1487350800, 1487354400, 1487358000, 
    1487361600, 1487365200, 1487368800, 1487372400, 1487376000, 1487379600, 
    1487383200, 1487386800, 1487390400, 1487394000, 1487397600, 1487401200, 
    1487404800, 1487408400, 1487412000, 1487415600, 1487419200, 1487422800, 
    1487426400, 1487430000, 1487433600, 1487437200, 1487440800, 1487444400, 
    1487448000, 1487451600, 1487455200, 1487458800, 1487462400, 1487466000, 
    1487469600, 1487473200, 1487476800, 1487480400, 1487484000, 1487487600, 
    1487491200, 1487494800, 1487498400, 1487502000, 1487505600, 1487509200, 
    1487512800, 1487516400, 1487520000, 1487523600, 1487527200, 1487530800, 
    1487534400, 1487538000, 1487541600, 1487545200, 1487548800, 1487552400, 
    1487556000, 1487559600, 1487563200, 1487566800, 1487570400, 1487574000, 
    1487577600, 1487581200, 1487584800, 1487588400, 1487592000, 1487595600, 
    1487599200, 1487602800, 1487606400, 1487610000, 1487613600, 1487617200, 
    1487620800, 1487624400, 1487628000, 1487631600, 1487635200, 1487638800, 
    1487642400, 1487646000, 1487649600, 1487653200, 1487656800, 1487660400, 
    1487664000, 1487667600, 1487671200, 1487674800, 1487678400, 1487682000, 
    1487685600, 1487689200, 1487692800, 1487696400, 1487700000, 1487703600, 
    1487707200, 1487710800, 1487714400, 1487718000, 1487721600, 1487725200, 
    1487728800, 1487732400, 1487736000, 1487739600, 1487743200, 1487746800, 
    1487750400, 1487754000, 1487757600, 1487761200, 1487764800, 1487768400, 
    1487772000, 1487775600, 1487779200, 1487782800, 1487786400, 1487790000, 
    1487793600, 1487797200, 1487800800, 1487804400, 1487808000, 1487811600, 
    1487815200, 1487818800, 1487822400, 1487826000, 1487829600, 1487833200, 
    1487836800, 1487840400, 1487844000, 1487847600, 1487851200, 1487854800, 
    1487858400, 1487862000, 1487865600, 1487869200, 1487872800, 1487876400, 
    1487880000, 1487883600, 1487887200, 1487890800, 1487894400, 1487898000, 
    1487901600, 1487905200, 1487908800, 1487912400, 1487916000, 1487919600, 
    1487923200, 1487926800, 1487930400, 1487934000, 1487937600, 1487941200, 
    1487944800, 1487948400, 1487952000, 1487955600, 1487959200, 1487962800, 
    1487966400, 1487970000, 1487973600, 1487977200, 1487980800, 1487984400, 
    1487988000, 1487991600, 1487995200, 1487998800, 1488002400, 1488006000, 
    1488009600, 1488013200, 1488016800, 1488020400, 1488024000, 1488027600, 
    1488031200, 1488034800, 1488038400, 1488042000, 1488045600, 1488049200, 
    1488052800, 1488056400, 1488060000, 1488063600, 1488067200, 1488070800, 
    1488074400, 1488078000, 1488081600, 1488085200, 1488088800, 1488092400, 
    1488096000, 1488099600, 1488103200, 1488106800, 1488110400, 1488114000, 
    1488117600, 1488121200, 1488124800, 1488128400, 1488132000, 1488135600, 
    1488139200, 1488142800, 1488146400, 1488150000, 1488153600, 1488157200, 
    1488160800, 1488164400, 1488168000, 1488171600, 1488175200, 1488178800, 
    1488182400, 1488186000, 1488189600, 1488193200, 1488196800, 1488200400, 
    1488204000, 1488207600, 1488211200, 1488214800, 1488218400, 1488222000, 
    1488225600, 1488229200, 1488232800, 1488236400, 1488240000, 1488243600, 
    1488247200, 1488250800, 1488254400, 1488258000, 1488261600, 1488265200, 
    1488268800, 1488272400, 1488276000, 1488279600, 1488283200, 1488286800, 
    1488290400, 1488294000, 1488297600, 1488301200, 1488304800, 1488308400, 
    1488312000, 1488315600, 1488319200, 1488322800, 1488326400, 1488330000, 
    1488333600, 1488337200, 1488340800, 1488344400, 1488348000, 1488351600, 
    1488355200, 1488358800, 1488362400, 1488366000, 1488369600, 1488373200, 
    1488376800, 1488380400, 1488384000, 1488387600, 1488391200, 1488394800, 
    1488398400, 1488402000, 1488405600, 1488409200, 1488412800, 1488416400, 
    1488420000, 1488423600, 1488427200, 1488430800, 1488434400, 1488438000, 
    1488441600, 1488445200, 1488448800, 1488452400, 1488456000, 1488459600, 
    1488463200, 1488466800, 1488470400, 1488474000, 1488477600, 1488481200, 
    1488484800, 1488488400, 1488492000, 1488495600, 1488499200, 1488502800, 
    1488506400, 1488510000, 1488513600, 1488517200, 1488520800, 1488524400, 
    1488528000, 1488531600, 1488535200, 1488538800, 1488542400, 1488546000, 
    1488549600, 1488553200, 1488556800, 1488560400, 1488564000, 1488567600, 
    1488571200, 1488574800, 1488578400, 1488582000, 1488585600, 1488589200, 
    1488592800, 1488596400, 1488600000, 1488603600, 1488607200, 1488610800, 
    1488614400, 1488618000, 1488621600, 1488625200, 1488628800, 1488632400, 
    1488636000, 1488639600, 1488643200, 1488646800, 1488650400, 1488654000, 
    1488657600, 1488661200, 1488664800, 1488668400, 1488672000, 1488675600, 
    1488679200, 1488682800, 1488686400, 1488690000, 1488693600, 1488697200, 
    1488700800, 1488704400, 1488708000, 1488711600, 1488715200, 1488718800, 
    1488722400, 1488726000, 1488729600, 1488733200, 1488736800, 1488740400, 
    1488744000, 1488747600, 1488751200, 1488754800, 1488758400, 1488762000, 
    1488765600, 1488769200, 1488772800, 1488776400, 1488780000, 1488783600, 
    1488787200, 1488790800, 1488794400, 1488798000, 1488801600, 1488805200, 
    1488808800, 1488812400, 1488816000, 1488819600, 1488823200, 1488826800, 
    1488830400, 1488834000, 1488837600, 1488841200, 1488844800, 1488848400, 
    1488852000, 1488855600, 1488859200, 1488862800, 1488866400, 1488870000, 
    1488873600, 1488877200, 1488880800, 1488884400, 1488888000, 1488891600, 
    1488895200, 1488898800, 1488902400, 1488906000, 1488909600, 1488913200, 
    1488916800, 1488920400, 1488924000, 1488927600, 1488931200, 1488934800, 
    1488938400, 1488942000, 1488945600, 1488949200, 1488952800, 1488956400, 
    1488960000, 1488963600, 1488967200, 1488970800, 1488974400, 1488978000, 
    1488981600, 1488985200, 1488988800, 1488992400, 1488996000, 1488999600, 
    1489003200, 1489006800, 1489010400, 1489014000, 1489017600, 1489021200, 
    1489024800, 1489028400, 1489032000, 1489035600, 1489039200, 1489042800, 
    1489046400, 1489050000, 1489053600, 1489057200, 1489060800, 1489064400, 
    1489068000, 1489071600, 1489075200, 1489078800, 1489082400, 1489086000, 
    1489089600, 1489093200, 1489096800, 1489100400, 1489104000, 1489107600, 
    1489111200, 1489114800, 1489118400, 1489122000, 1489125600, 1489129200, 
    1489132800, 1489136400, 1489140000, 1489143600, 1489147200, 1489150800, 
    1489154400, 1489158000, 1489161600, 1489165200, 1489168800, 1489172400, 
    1489176000, 1489179600, 1489183200, 1489186800, 1489190400, 1489194000, 
    1489197600, 1489201200, 1489204800, 1489208400, 1489212000, 1489215600, 
    1489219200, 1489222800, 1489226400, 1489230000, 1489233600, 1489237200, 
    1489240800, 1489244400, 1489248000, 1489251600, 1489255200, 1489258800, 
    1489262400, 1489266000, 1489269600, 1489273200, 1489276800, 1489280400, 
    1489284000, 1489287600, 1489291200, 1489294800, 1489298400, 1489302000, 
    1489305600, 1489309200, 1489312800, 1489316400, 1489320000, 1489323600, 
    1489327200, 1489330800, 1489334400, 1489338000, 1489341600, 1489345200, 
    1489348800, 1489352400, 1489356000, 1489359600, 1489363200, 1489366800, 
    1489370400, 1489374000, 1489377600, 1489381200, 1489384800, 1489388400, 
    1489392000, 1489395600, 1489399200, 1489402800, 1489406400, 1489410000, 
    1489413600, 1489417200, 1489420800, 1489424400, 1489428000, 1489431600, 
    1489435200, 1489438800, 1489442400, 1489446000, 1489449600, 1489453200, 
    1489456800, 1489460400, 1489464000, 1489467600, 1489471200, 1489474800, 
    1489478400, 1489482000, 1489485600, 1489489200, 1489492800, 1489496400, 
    1489500000, 1489503600, 1489507200, 1489510800, 1489514400, 1489518000, 
    1489521600, 1489525200, 1489528800, 1489532400, 1489536000, 1489539600, 
    1489543200, 1489546800, 1489550400, 1489554000, 1489557600, 1489561200, 
    1489564800, 1489568400, 1489572000, 1489575600, 1489579200, 1489582800, 
    1489586400, 1489590000, 1489593600, 1489597200, 1489600800, 1489604400, 
    1489608000, 1489611600, 1489615200, 1489618800, 1489622400, 1489626000, 
    1489629600, 1489633200, 1489636800, 1489640400, 1489644000, 1489647600, 
    1489651200, 1489654800, 1489658400, 1489662000, 1489665600, 1489669200, 
    1489672800, 1489676400, 1489680000, 1489683600, 1489687200, 1489690800, 
    1489694400, 1489698000, 1489701600, 1489705200, 1489708800, 1489712400, 
    1489716000, 1489719600, 1489723200, 1489726800, 1489730400, 1489734000, 
    1489737600, 1489741200, 1489744800, 1489748400, 1489752000, 1489755600, 
    1489759200, 1489762800, 1489766400, 1489770000, 1489773600, 1489777200, 
    1489780800, 1489784400, 1489788000, 1489791600, 1489795200, 1489798800, 
    1489802400, 1489806000, 1489809600, 1489813200, 1489816800, 1489820400, 
    1489824000, 1489827600, 1489831200, 1489834800, 1489838400, 1489842000, 
    1489845600, 1489849200, 1489852800, 1489856400, 1489860000, 1489863600, 
    1489867200, 1489870800, 1489874400, 1489878000, 1489881600, 1489885200, 
    1489888800, 1489892400, 1489896000, 1489899600, 1489903200, 1489906800, 
    1489910400, 1489914000, 1489917600, 1489921200, 1489924800, 1489928400, 
    1489932000, 1489935600, 1489939200, 1489942800, 1489946400, 1489950000, 
    1489953600, 1489957200, 1489960800, 1489964400, 1489968000, 1489971600, 
    1489975200, 1489978800, 1489982400, 1489986000, 1489989600, 1489993200, 
    1489996800, 1490000400, 1490004000, 1490007600, 1490011200, 1490014800, 
    1490018400, 1490022000, 1490025600, 1490029200, 1490032800, 1490036400, 
    1490040000, 1490043600, 1490047200, 1490050800, 1490054400, 1490058000, 
    1490061600, 1490065200, 1490068800, 1490072400, 1490076000, 1490079600, 
    1490083200, 1490086800, 1490090400, 1490094000, 1490097600, 1490101200, 
    1490104800, 1490108400, 1490112000, 1490115600, 1490119200, 1490122800, 
    1490126400, 1490130000, 1490133600, 1490137200, 1490140800, 1490144400, 
    1490148000, 1490151600, 1490155200, 1490158800, 1490162400, 1490166000, 
    1490169600, 1490173200, 1490176800, 1490180400, 1490184000, 1490187600, 
    1490191200, 1490194800, 1490198400, 1490202000, 1490205600, 1490209200, 
    1490212800, 1490216400, 1490220000, 1490223600, 1490227200, 1490230800, 
    1490234400, 1490238000, 1490241600, 1490245200, 1490248800, 1490252400, 
    1490256000, 1490259600, 1490263200, 1490266800, 1490270400, 1490274000, 
    1490277600, 1490281200, 1490284800, 1490288400, 1490292000, 1490295600, 
    1490299200, 1490302800, 1490306400, 1490310000, 1490313600, 1490317200, 
    1490320800, 1490324400, 1490328000, 1490331600, 1490335200, 1490338800, 
    1490342400, 1490346000, 1490349600, 1490353200, 1490356800, 1490360400, 
    1490364000, 1490367600, 1490371200, 1490374800, 1490378400, 1490382000, 
    1490385600, 1490389200, 1490392800, 1490396400, 1490400000, 1490403600, 
    1490407200, 1490410800, 1490414400, 1490418000, 1490421600, 1490425200, 
    1490428800, 1490432400, 1490436000, 1490439600, 1490443200, 1490446800, 
    1490450400, 1490454000, 1490457600, 1490461200, 1490464800, 1490468400, 
    1490472000, 1490475600, 1490479200, 1490482800, 1490486400, 1490490000, 
    1490493600, 1490497200, 1490500800, 1490504400, 1490508000, 1490511600, 
    1490515200, 1490518800, 1490522400, 1490526000, 1490529600, 1490533200, 
    1490536800, 1490540400, 1490544000, 1490547600, 1490551200, 1490554800, 
    1490558400, 1490562000, 1490565600, 1490569200, 1490572800, 1490576400, 
    1490580000, 1490583600, 1490587200, 1490590800, 1490594400, 1490598000, 
    1490601600, 1490605200, 1490608800, 1490612400, 1490616000, 1490619600, 
    1490623200, 1490626800, 1490630400, 1490634000, 1490637600, 1490641200, 
    1490644800, 1490648400, 1490652000, 1490655600, 1490659200, 1490662800, 
    1490666400, 1490670000, 1490673600, 1490677200, 1490680800, 1490684400, 
    1490688000, 1490691600, 1490695200, 1490698800, 1490702400, 1490706000, 
    1490709600, 1490713200, 1490716800, 1490720400, 1490724000, 1490727600, 
    1490731200, 1490734800, 1490738400, 1490742000, 1490745600, 1490749200, 
    1490752800, 1490756400, 1490760000, 1490763600, 1490767200, 1490770800, 
    1490774400, 1490778000, 1490781600, 1490785200, 1490788800, 1490792400, 
    1490796000, 1490799600, 1490803200, 1490806800, 1490810400, 1490814000, 
    1490817600, 1490821200, 1490824800, 1490828400, 1490832000, 1490835600, 
    1490839200, 1490842800, 1490846400, 1490850000, 1490853600, 1490857200, 
    1490860800, 1490864400, 1490868000, 1490871600, 1490875200, 1490878800, 
    1490882400, 1490886000, 1490889600, 1490893200, 1490896800, 1490900400, 
    1490904000, 1490907600, 1490911200, 1490914800, 1490918400, 1490922000, 
    1490925600, 1490929200, 1490932800, 1490936400, 1490940000, 1490943600, 
    1490947200, 1490950800, 1490954400, 1490958000, 1490961600, 1490965200, 
    1490968800, 1490972400, 1490976000, 1490979600, 1490983200, 1490986800, 
    1490990400, 1490994000, 1490997600, 1491001200, 1491004800, 1491008400, 
    1491012000, 1491015600, 1491019200, 1491022800, 1491026400, 1491030000, 
    1491033600, 1491037200, 1491040800, 1491044400, 1491048000, 1491051600, 
    1491055200, 1491058800, 1491062400, 1491066000, 1491069600, 1491073200, 
    1491076800, 1491080400, 1491084000, 1491087600, 1491091200, 1491094800, 
    1491098400, 1491102000, 1491105600, 1491109200, 1491112800, 1491116400, 
    1491120000, 1491123600, 1491127200, 1491130800, 1491134400, 1491138000, 
    1491141600, 1491145200, 1491148800, 1491152400, 1491156000, 1491159600, 
    1491163200, 1491166800, 1491170400, 1491174000, 1491177600, 1491181200, 
    1491184800, 1491188400, 1491192000, 1491195600, 1491199200, 1491202800, 
    1491206400, 1491210000, 1491213600, 1491217200, 1491220800, 1491224400, 
    1491228000, 1491231600, 1491235200, 1491238800, 1491242400, 1491246000, 
    1491249600, 1491253200, 1491256800, 1491260400, 1491264000, 1491267600, 
    1491271200, 1491274800, 1491278400, 1491282000, 1491285600, 1491289200, 
    1491292800, 1491296400, 1491300000, 1491303600, 1491307200, 1491310800, 
    1491314400, 1491318000, 1491321600, 1491325200, 1491328800, 1491332400, 
    1491336000, 1491339600, 1491343200, 1491346800, 1491350400, 1491354000, 
    1491357600, 1491361200, 1491364800, 1491368400, 1491372000, 1491375600, 
    1491379200, 1491382800, 1491386400, 1491390000, 1491393600, 1491397200, 
    1491400800, 1491404400, 1491408000, 1491411600, 1491415200, 1491418800, 
    1491422400, 1491426000, 1491429600, 1491433200, 1491436800, 1491440400, 
    1491444000, 1491447600, 1491451200, 1491454800, 1491458400, 1491462000, 
    1491465600, 1491469200, 1491472800, 1491476400, 1491480000, 1491483600, 
    1491487200, 1491490800, 1491494400, 1491498000, 1491501600, 1491505200, 
    1491508800, 1491512400, 1491516000, 1491519600, 1491523200, 1491526800, 
    1491530400, 1491534000, 1491537600, 1491541200, 1491544800, 1491548400, 
    1491552000, 1491555600, 1491559200, 1491562800, 1491566400, 1491570000, 
    1491573600, 1491577200, 1491580800, 1491584400, 1491588000, 1491591600, 
    1491595200, 1491598800, 1491602400, 1491606000, 1491609600, 1491613200, 
    1491616800, 1491620400, 1491624000, 1491627600, 1491631200, 1491634800, 
    1491638400, 1491642000, 1491645600, 1491649200, 1491652800, 1491656400, 
    1491660000, 1491663600, 1491667200, 1491670800, 1491674400, 1491678000, 
    1491681600, 1491685200, 1491688800, 1491692400, 1491696000, 1491699600, 
    1491703200, 1491706800, 1491710400, 1491714000, 1491717600, 1491721200, 
    1491724800, 1491728400, 1491732000, 1491735600, 1491739200, 1491742800, 
    1491746400, 1491750000, 1491753600, 1491757200, 1491760800, 1491764400, 
    1491768000, 1491771600, 1491775200, 1491778800, 1491782400, 1491786000, 
    1491789600, 1491793200, 1491796800, 1491800400, 1491804000, 1491807600, 
    1491811200, 1491814800, 1491818400, 1491822000, 1491825600, 1491829200, 
    1491832800, 1491836400, 1491840000, 1491843600, 1491847200, 1491850800, 
    1491854400, 1491858000, 1491861600, 1491865200, 1491868800, 1491872400, 
    1491876000, 1491879600, 1491883200, 1491886800, 1491890400, 1491894000, 
    1491897600, 1491901200, 1491904800, 1491908400, 1491912000, 1491915600, 
    1491919200, 1491922800, 1491926400, 1491930000, 1491933600, 1491937200, 
    1491940800, 1491944400, 1491948000, 1491951600, 1491955200, 1491958800, 
    1491962400, 1491966000, 1491969600, 1491973200, 1491976800, 1491980400, 
    1491984000, 1491987600, 1491991200, 1491994800, 1491998400, 1492002000, 
    1492005600, 1492009200, 1492012800, 1492016400, 1492020000, 1492023600, 
    1492027200, 1492030800, 1492034400, 1492038000, 1492041600, 1492045200, 
    1492048800, 1492052400, 1492056000, 1492059600, 1492063200, 1492066800, 
    1492070400, 1492074000, 1492077600, 1492081200, 1492084800, 1492088400, 
    1492092000, 1492095600, 1492099200, 1492102800, 1492106400, 1492110000, 
    1492113600, 1492117200, 1492120800, 1492124400, 1492128000, 1492131600, 
    1492135200, 1492138800, 1492142400, 1492146000, 1492149600, 1492153200, 
    1492156800, 1492160400, 1492164000, 1492167600, 1492171200, 1492174800, 
    1492178400, 1492182000, 1492185600, 1492189200, 1492192800, 1492196400, 
    1492200000, 1492203600, 1492207200, 1492210800, 1492214400, 1492218000, 
    1492221600, 1492225200, 1492228800, 1492232400, 1492236000, 1492239600, 
    1492243200, 1492246800, 1492250400, 1492254000, 1492257600, 1492261200, 
    1492264800, 1492268400, 1492272000, 1492275600, 1492279200, 1492282800, 
    1492286400, 1492290000, 1492293600, 1492297200, 1492300800, 1492304400, 
    1492308000, 1492311600, 1492315200, 1492318800, 1492322400, 1492326000, 
    1492329600, 1492333200, 1492336800, 1492340400, 1492344000, 1492347600, 
    1492351200, 1492354800, 1492358400, 1492362000, 1492365600, 1492369200, 
    1492372800, 1492376400, 1492380000, 1492383600, 1492387200, 1492390800, 
    1492394400, 1492398000, 1492401600, 1492405200, 1492408800, 1492412400, 
    1492416000, 1492419600, 1492423200, 1492426800, 1492430400, 1492434000, 
    1492437600, 1492441200, 1492444800, 1492448400, 1492452000, 1492455600, 
    1492459200, 1492462800, 1492466400, 1492470000, 1492473600, 1492477200, 
    1492480800, 1492484400, 1492488000, 1492491600, 1492495200, 1492498800, 
    1492502400, 1492506000, 1492509600, 1492513200, 1492516800, 1492520400, 
    1492524000, 1492527600, 1492531200, 1492534800, 1492538400, 1492542000, 
    1492545600, 1492549200, 1492552800, 1492556400, 1492560000, 1492563600, 
    1492567200, 1492570800, 1492574400, 1492578000, 1492581600, 1492585200, 
    1492588800, 1492592400, 1492596000, 1492599600, 1492603200, 1492606800, 
    1492610400, 1492614000, 1492617600, 1492621200, 1492624800, 1492628400, 
    1492632000, 1492635600, 1492639200, 1492642800, 1492646400, 1492650000, 
    1492653600, 1492657200, 1492660800, 1492664400, 1492668000, 1492671600, 
    1492675200, 1492678800, 1492682400, 1492686000, 1492689600, 1492693200, 
    1492696800, 1492700400, 1492704000, 1492707600, 1492711200, 1492714800, 
    1492718400, 1492722000, 1492725600, 1492729200, 1492732800, 1492736400, 
    1492740000, 1492743600, 1492747200, 1492750800, 1492754400, 1492758000, 
    1492761600, 1492765200, 1492768800, 1492772400, 1492776000, 1492779600, 
    1492783200, 1492786800, 1492790400, 1492794000, 1492797600, 1492801200, 
    1492804800, 1492808400, 1492812000, 1492815600, 1492819200, 1492822800, 
    1492826400, 1492830000, 1492833600, 1492837200, 1492840800, 1492844400, 
    1492848000, 1492851600, 1492855200, 1492858800, 1492862400, 1492866000, 
    1492869600, 1492873200, 1492876800, 1492880400, 1492884000, 1492887600, 
    1492891200, 1492894800, 1492898400, 1492902000, 1492905600, 1492909200, 
    1492912800, 1492916400, 1492920000, 1492923600, 1492927200, 1492930800, 
    1492934400, 1492938000, 1492941600, 1492945200, 1492948800, 1492952400, 
    1492956000, 1492959600, 1492963200, 1492966800, 1492970400, 1492974000, 
    1492977600, 1492981200, 1492984800, 1492988400, 1492992000, 1492995600, 
    1492999200, 1493002800, 1493006400, 1493010000, 1493013600, 1493017200, 
    1493020800, 1493024400, 1493028000, 1493031600, 1493035200, 1493038800, 
    1493042400, 1493046000, 1493049600, 1493053200, 1493056800, 1493060400, 
    1493064000, 1493067600, 1493071200, 1493074800, 1493078400, 1493082000, 
    1493085600, 1493089200, 1493092800, 1493096400, 1493100000, 1493103600, 
    1493107200, 1493110800, 1493114400, 1493118000, 1493121600, 1493125200, 
    1493128800, 1493132400, 1493136000, 1493139600, 1493143200, 1493146800, 
    1493150400, 1493154000, 1493157600, 1493161200, 1493164800, 1493168400, 
    1493172000, 1493175600, 1493179200, 1493182800, 1493186400, 1493190000, 
    1493193600, 1493197200, 1493200800, 1493204400, 1493208000, 1493211600, 
    1493215200, 1493218800, 1493222400, 1493226000, 1493229600, 1493233200, 
    1493236800, 1493240400, 1493244000, 1493247600, 1493251200, 1493254800, 
    1493258400, 1493262000, 1493265600, 1493269200, 1493272800, 1493276400, 
    1493280000, 1493283600, 1493287200, 1493290800, 1493294400, 1493298000, 
    1493301600, 1493305200, 1493308800, 1493312400, 1493316000, 1493319600, 
    1493323200, 1493326800, 1493330400, 1493334000, 1493337600, 1493341200, 
    1493344800, 1493348400, 1493352000, 1493355600, 1493359200, 1493362800, 
    1493366400, 1493370000, 1493373600, 1493377200, 1493380800, 1493384400, 
    1493388000, 1493391600, 1493395200, 1493398800, 1493402400, 1493406000, 
    1493409600, 1493413200, 1493416800, 1493420400, 1493424000, 1493427600, 
    1493431200, 1493434800, 1493438400, 1493442000, 1493445600, 1493449200, 
    1493452800, 1493456400, 1493460000, 1493463600, 1493467200, 1493470800, 
    1493474400, 1493478000, 1493481600, 1493485200, 1493488800, 1493492400, 
    1493496000, 1493499600, 1493503200, 1493506800, 1493510400, 1493514000, 
    1493517600, 1493521200, 1493524800, 1493528400, 1493532000, 1493535600, 
    1493539200, 1493542800, 1493546400, 1493550000, 1493553600, 1493557200, 
    1493560800, 1493564400, 1493568000, 1493571600, 1493575200, 1493578800, 
    1493582400, 1493586000, 1493589600, 1493593200, 1493596800, 1493600400, 
    1493604000, 1493607600, 1493611200, 1493614800, 1493618400, 1493622000, 
    1493625600, 1493629200, 1493632800, 1493636400, 1493640000, 1493643600, 
    1493647200, 1493650800, 1493654400, 1493658000, 1493661600, 1493665200, 
    1493668800, 1493672400, 1493676000, 1493679600, 1493683200, 1493686800, 
    1493690400, 1493694000, 1493697600, 1493701200, 1493704800, 1493708400, 
    1493712000, 1493715600, 1493719200, 1493722800, 1493726400, 1493730000, 
    1493733600, 1493737200, 1493740800, 1493744400, 1493748000, 1493751600, 
    1493755200, 1493758800, 1493762400, 1493766000, 1493769600, 1493773200, 
    1493776800, 1493780400, 1493784000, 1493787600, 1493791200, 1493794800, 
    1493798400, 1493802000, 1493805600, 1493809200, 1493812800, 1493816400, 
    1493820000, 1493823600, 1493827200, 1493830800, 1493834400, 1493838000, 
    1493841600, 1493845200, 1493848800, 1493852400, 1493856000, 1493859600, 
    1493863200, 1493866800, 1493870400, 1493874000, 1493877600, 1493881200, 
    1493884800, 1493888400, 1493892000, 1493895600, 1493899200, 1493902800, 
    1493906400, 1493910000, 1493913600, 1493917200, 1493920800, 1493924400, 
    1493928000, 1493931600, 1493935200, 1493938800, 1493942400, 1493946000, 
    1493949600, 1493953200, 1493956800, 1493960400, 1493964000, 1493967600, 
    1493971200, 1493974800, 1493978400, 1493982000, 1493985600, 1493989200, 
    1493992800, 1493996400, 1494000000, 1494003600, 1494007200, 1494010800, 
    1494014400, 1494018000, 1494021600, 1494025200, 1494028800, 1494032400, 
    1494036000, 1494039600, 1494043200, 1494046800, 1494050400, 1494054000, 
    1494057600, 1494061200, 1494064800, 1494068400, 1494072000, 1494075600, 
    1494079200, 1494082800, 1494086400, 1494090000, 1494093600, 1494097200, 
    1494100800, 1494104400, 1494108000, 1494111600, 1494115200, 1494118800, 
    1494122400, 1494126000, 1494129600, 1494133200, 1494136800, 1494140400, 
    1494144000, 1494147600, 1494151200, 1494154800, 1494158400, 1494162000, 
    1494165600, 1494169200, 1494172800, 1494176400, 1494180000, 1494183600, 
    1494187200, 1494190800, 1494194400, 1494198000, 1494201600, 1494205200, 
    1494208800, 1494212400, 1494216000, 1494219600, 1494223200, 1494226800, 
    1494230400, 1494234000, 1494237600, 1494241200, 1494244800, 1494248400, 
    1494252000, 1494255600, 1494259200, 1494262800, 1494266400, 1494270000, 
    1494273600, 1494277200, 1494280800, 1494284400, 1494288000, 1494291600, 
    1494295200, 1494298800, 1494302400, 1494306000, 1494309600, 1494313200, 
    1494316800, 1494320400, 1494324000, 1494327600, 1494331200, 1494334800, 
    1494338400, 1494342000, 1494345600, 1494349200, 1494352800, 1494356400, 
    1494360000, 1494363600, 1494367200, 1494370800, 1494374400, 1494378000, 
    1494381600, 1494385200, 1494388800, 1494392400, 1494396000, 1494399600, 
    1494403200, 1494406800, 1494410400, 1494414000, 1494417600, 1494421200, 
    1494424800, 1494428400, 1494432000, 1494435600, 1494439200, 1494442800, 
    1494446400, 1494450000, 1494453600, 1494457200, 1494460800, 1494464400, 
    1494468000, 1494471600, 1494475200, 1494478800, 1494482400, 1494486000, 
    1494489600, 1494493200, 1494496800, 1494500400, 1494504000, 1494507600, 
    1494511200, 1494514800, 1494518400, 1494522000, 1494525600, 1494529200, 
    1494532800, 1494536400, 1494540000, 1494543600, 1494547200, 1494550800, 
    1494554400, 1494558000, 1494561600, 1494565200, 1494568800, 1494572400, 
    1494576000, 1494579600, 1494583200, 1494586800, 1494590400, 1494594000, 
    1494597600, 1494601200, 1494604800, 1494608400, 1494612000, 1494615600, 
    1494619200, 1494622800, 1494626400, 1494630000, 1494633600, 1494637200, 
    1494640800, 1494644400, 1494648000, 1494651600, 1494655200, 1494658800, 
    1494662400, 1494666000, 1494669600, 1494673200, 1494676800, 1494680400, 
    1494684000, 1494687600, 1494691200, 1494694800, 1494698400, 1494702000, 
    1494705600, 1494709200, 1494712800, 1494716400, 1494720000, 1494723600, 
    1494727200, 1494730800, 1494734400, 1494738000, 1494741600, 1494745200, 
    1494748800, 1494752400, 1494756000, 1494759600, 1494763200, 1494766800, 
    1494770400, 1494774000, 1494777600, 1494781200, 1494784800, 1494788400, 
    1494792000, 1494795600, 1494799200, 1494802800, 1494806400, 1494810000, 
    1494813600, 1494817200, 1494820800, 1494824400, 1494828000, 1494831600, 
    1494835200, 1494838800, 1494842400, 1494846000, 1494849600, 1494853200, 
    1494856800, 1494860400, 1494864000, 1494867600, 1494871200, 1494874800, 
    1494878400, 1494882000, 1494885600, 1494889200, 1494892800, 1494896400, 
    1494900000, 1494903600, 1494907200, 1494910800, 1494914400, 1494918000, 
    1494921600, 1494925200, 1494928800, 1494932400, 1494936000, 1494939600, 
    1494943200, 1494946800, 1494950400, 1494954000, 1494957600, 1494961200, 
    1494964800, 1494968400, 1494972000, 1494975600, 1494979200, 1494982800, 
    1494986400, 1494990000, 1494993600, 1494997200, 1495000800, 1495004400, 
    1495008000, 1495011600, 1495015200, 1495018800, 1495022400, 1495026000, 
    1495029600, 1495033200, 1495036800, 1495040400, 1495044000, 1495047600, 
    1495051200, 1495054800, 1495058400, 1495062000, 1495065600, 1495069200, 
    1495072800, 1495076400, 1495080000, 1495083600, 1495087200, 1495090800, 
    1495094400, 1495098000, 1495101600, 1495105200, 1495108800, 1495112400, 
    1495116000, 1495119600, 1495123200, 1495126800, 1495130400, 1495134000, 
    1495137600, 1495141200, 1495144800, 1495148400, 1495152000, 1495155600, 
    1495159200, 1495162800, 1495166400, 1495170000, 1495173600, 1495177200, 
    1495180800, 1495184400, 1495188000, 1495191600, 1495195200, 1495198800, 
    1495202400, 1495206000, 1495209600, 1495213200, 1495216800, 1495220400, 
    1495224000, 1495227600, 1495231200, 1495234800, 1495238400, 1495242000, 
    1495245600, 1495249200, 1495252800, 1495256400, 1495260000, 1495263600, 
    1495267200, 1495270800, 1495274400, 1495278000, 1495281600, 1495285200, 
    1495288800, 1495292400, 1495296000, 1495299600, 1495303200, 1495306800, 
    1495310400, 1495314000, 1495317600, 1495321200, 1495324800, 1495328400, 
    1495332000, 1495335600, 1495339200, 1495342800, 1495346400, 1495350000, 
    1495353600, 1495357200, 1495360800, 1495364400, 1495368000, 1495371600, 
    1495375200, 1495378800, 1495382400, 1495386000, 1495389600, 1495393200, 
    1495396800, 1495400400, 1495404000, 1495407600, 1495411200, 1495414800, 
    1495418400, 1495422000, 1495425600, 1495429200, 1495432800, 1495436400, 
    1495440000, 1495443600, 1495447200, 1495450800, 1495454400, 1495458000, 
    1495461600, 1495465200, 1495468800, 1495472400, 1495476000, 1495479600, 
    1495483200, 1495486800, 1495490400, 1495494000, 1495497600, 1495501200, 
    1495504800, 1495508400, 1495512000, 1495515600, 1495519200, 1495522800, 
    1495526400, 1495530000, 1495533600, 1495537200, 1495540800, 1495544400, 
    1495548000, 1495551600, 1495555200, 1495558800, 1495562400, 1495566000, 
    1495569600, 1495573200, 1495576800, 1495580400, 1495584000, 1495587600, 
    1495591200, 1495594800, 1495598400, 1495602000, 1495605600, 1495609200, 
    1495612800, 1495616400, 1495620000, 1495623600, 1495627200, 1495630800, 
    1495634400, 1495638000, 1495641600, 1495645200, 1495648800, 1495652400, 
    1495656000, 1495659600, 1495663200, 1495666800, 1495670400, 1495674000, 
    1495677600, 1495681200, 1495684800, 1495688400, 1495692000, 1495695600, 
    1495699200, 1495702800, 1495706400, 1495710000, 1495713600, 1495717200, 
    1495720800, 1495724400, 1495728000, 1495731600, 1495735200, 1495738800, 
    1495742400, 1495746000, 1495749600, 1495753200, 1495756800, 1495760400, 
    1495764000, 1495767600, 1495771200, 1495774800, 1495778400, 1495782000, 
    1495785600, 1495789200, 1495792800, 1495796400, 1495800000, 1495803600, 
    1495807200, 1495810800, 1495814400, 1495818000, 1495821600, 1495825200, 
    1495828800, 1495832400, 1495836000, 1495839600, 1495843200, 1495846800, 
    1495850400, 1495854000, 1495857600, 1495861200, 1495864800, 1495868400, 
    1495872000, 1495875600, 1495879200, 1495882800, 1495886400, 1495890000, 
    1495893600, 1495897200, 1495900800, 1495904400, 1495908000, 1495911600, 
    1495915200, 1495918800, 1495922400, 1495926000, 1495929600, 1495933200, 
    1495936800, 1495940400, 1495944000, 1495947600, 1495951200, 1495954800, 
    1495958400, 1495962000, 1495965600, 1495969200, 1495972800, 1495976400, 
    1495980000, 1495983600, 1495987200, 1495990800, 1495994400, 1495998000, 
    1496001600, 1496005200, 1496008800, 1496012400, 1496016000, 1496019600, 
    1496023200, 1496026800, 1496030400, 1496034000, 1496037600, 1496041200, 
    1496044800, 1496048400, 1496052000, 1496055600, 1496059200, 1496062800, 
    1496066400, 1496070000, 1496073600, 1496077200, 1496080800, 1496084400, 
    1496088000, 1496091600, 1496095200, 1496098800, 1496102400, 1496106000, 
    1496109600, 1496113200, 1496116800, 1496120400, 1496124000, 1496127600, 
    1496131200, 1496134800, 1496138400, 1496142000, 1496145600, 1496149200, 
    1496152800, 1496156400, 1496160000, 1496163600, 1496167200, 1496170800, 
    1496174400, 1496178000, 1496181600, 1496185200, 1496188800, 1496192400, 
    1496196000, 1496199600, 1496203200, 1496206800, 1496210400, 1496214000, 
    1496217600, 1496221200, 1496224800, 1496228400, 1496232000, 1496235600, 
    1496239200, 1496242800, 1496246400, 1496250000, 1496253600, 1496257200, 
    1496260800, 1496264400, 1496268000, 1496271600, 1496275200, 1496278800, 
    1496282400, 1496286000, 1496289600, 1496293200, 1496296800, 1496300400, 
    1496304000, 1496307600, 1496311200, 1496314800, 1496318400, 1496322000, 
    1496325600, 1496329200, 1496332800, 1496336400, 1496340000, 1496343600, 
    1496347200, 1496350800, 1496354400, 1496358000, 1496361600, 1496365200, 
    1496368800, 1496372400, 1496376000, 1496379600, 1496383200, 1496386800, 
    1496390400, 1496394000, 1496397600, 1496401200, 1496404800, 1496408400, 
    1496412000, 1496415600, 1496419200, 1496422800, 1496426400, 1496430000, 
    1496433600, 1496437200, 1496440800, 1496444400, 1496448000, 1496451600, 
    1496455200, 1496458800, 1496462400, 1496466000, 1496469600, 1496473200, 
    1496476800, 1496480400, 1496484000, 1496487600, 1496491200, 1496494800, 
    1496498400, 1496502000, 1496505600, 1496509200, 1496512800, 1496516400, 
    1496520000, 1496523600, 1496527200, 1496530800, 1496534400, 1496538000, 
    1496541600, 1496545200, 1496548800, 1496552400, 1496556000, 1496559600, 
    1496563200, 1496566800, 1496570400, 1496574000, 1496577600, 1496581200, 
    1496584800, 1496588400, 1496592000, 1496595600, 1496599200, 1496602800, 
    1496606400, 1496610000, 1496613600, 1496617200, 1496620800, 1496624400, 
    1496628000, 1496631600, 1496635200, 1496638800, 1496642400, 1496646000, 
    1496649600, 1496653200, 1496656800, 1496660400, 1496664000, 1496667600, 
    1496671200, 1496674800, 1496678400, 1496682000, 1496685600, 1496689200, 
    1496692800, 1496696400, 1496700000, 1496703600, 1496707200, 1496710800, 
    1496714400, 1496718000, 1496721600, 1496725200, 1496728800, 1496732400, 
    1496736000, 1496739600, 1496743200, 1496746800, 1496750400, 1496754000, 
    1496757600, 1496761200, 1496764800, 1496768400, 1496772000, 1496775600, 
    1496779200, 1496782800, 1496786400, 1496790000, 1496793600, 1496797200, 
    1496800800, 1496804400, 1496808000, 1496811600, 1496815200, 1496818800, 
    1496822400, 1496826000, 1496829600, 1496833200, 1496836800, 1496840400, 
    1496844000, 1496847600, 1496851200, 1496854800, 1496858400, 1496862000, 
    1496865600, 1496869200, 1496872800, 1496876400, 1496880000, 1496883600, 
    1496887200, 1496890800, 1496894400, 1496898000, 1496901600, 1496905200, 
    1496908800, 1496912400, 1496916000, 1496919600, 1496923200, 1496926800, 
    1496930400, 1496934000, 1496937600, 1496941200, 1496944800, 1496948400, 
    1496952000, 1496955600, 1496959200, 1496962800, 1496966400, 1496970000, 
    1496973600, 1496977200, 1496980800, 1496984400, 1496988000, 1496991600, 
    1496995200, 1496998800, 1497002400, 1497006000, 1497009600, 1497013200, 
    1497016800, 1497020400, 1497024000, 1497027600, 1497031200, 1497034800, 
    1497038400, 1497042000, 1497045600, 1497049200, 1497052800, 1497056400, 
    1497060000, 1497063600, 1497067200, 1497070800, 1497074400, 1497078000, 
    1497081600, 1497085200, 1497088800, 1497092400, 1497096000, 1497099600, 
    1497103200, 1497106800, 1497110400, 1497114000, 1497117600, 1497121200, 
    1497124800, 1497128400, 1497132000, 1497135600, 1497139200, 1497142800, 
    1497146400, 1497150000, 1497153600, 1497157200, 1497160800, 1497164400, 
    1497168000, 1497171600, 1497175200, 1497178800, 1497182400, 1497186000, 
    1497189600, 1497193200, 1497196800, 1497200400, 1497204000, 1497207600, 
    1497211200, 1497214800, 1497218400, 1497222000, 1497225600, 1497229200, 
    1497232800, 1497236400, 1497240000, 1497243600, 1497247200, 1497250800, 
    1497254400, 1497258000, 1497261600, 1497265200, 1497268800, 1497272400, 
    1497276000, 1497279600, 1497283200, 1497286800, 1497290400, 1497294000, 
    1497297600, 1497301200, 1497304800, 1497308400, 1497312000, 1497315600, 
    1497319200, 1497322800, 1497326400, 1497330000, 1497333600, 1497337200, 
    1497340800, 1497344400, 1497348000, 1497351600, 1497355200, 1497358800, 
    1497362400, 1497366000, 1497369600, 1497373200, 1497376800, 1497380400, 
    1497384000, 1497387600, 1497391200, 1497394800, 1497398400, 1497402000, 
    1497405600, 1497409200, 1497412800, 1497416400, 1497420000, 1497423600, 
    1497427200, 1497430800, 1497434400, 1497438000, 1497441600, 1497445200, 
    1497448800, 1497452400, 1497456000, 1497459600, 1497463200, 1497466800, 
    1497470400, 1497474000, 1497477600, 1497481200, 1497484800, 1497488400, 
    1497492000, 1497495600, 1497499200, 1497502800, 1497506400, 1497510000, 
    1497513600, 1497517200, 1497520800, 1497524400, 1497528000, 1497531600, 
    1497535200, 1497538800, 1497542400, 1497546000, 1497549600, 1497553200, 
    1497556800, 1497560400, 1497564000, 1497567600, 1497571200, 1497574800, 
    1497578400, 1497582000, 1497585600, 1497589200, 1497592800, 1497596400, 
    1497600000, 1497603600, 1497607200, 1497610800, 1497614400, 1497618000, 
    1497621600, 1497625200, 1497628800, 1497632400, 1497636000, 1497639600, 
    1497643200, 1497646800, 1497650400, 1497654000, 1497657600, 1497661200, 
    1497664800, 1497668400, 1497672000, 1497675600, 1497679200, 1497682800, 
    1497686400, 1497690000, 1497693600, 1497697200, 1497700800, 1497704400, 
    1497708000, 1497711600, 1497715200, 1497718800, 1497722400, 1497726000, 
    1497729600, 1497733200, 1497736800, 1497740400, 1497744000, 1497747600, 
    1497751200, 1497754800, 1497758400, 1497762000, 1497765600, 1497769200, 
    1497772800, 1497776400, 1497780000, 1497783600, 1497787200, 1497790800, 
    1497794400, 1497798000, 1497801600, 1497805200, 1497808800, 1497812400, 
    1497816000, 1497819600, 1497823200, 1497826800, 1497830400, 1497834000, 
    1497837600, 1497841200, 1497844800, 1497848400, 1497852000, 1497855600, 
    1497859200, 1497862800, 1497866400, 1497870000, 1497873600, 1497877200, 
    1497880800, 1497884400, 1497888000, 1497891600, 1497895200, 1497898800, 
    1497902400, 1497906000, 1497909600, 1497913200, 1497916800, 1497920400, 
    1497924000, 1497927600, 1497931200, 1497934800, 1497938400, 1497942000, 
    1497945600, 1497949200, 1497952800, 1497956400, 1497960000, 1497963600, 
    1497967200, 1497970800, 1497974400, 1497978000, 1497981600, 1497985200, 
    1497988800, 1497992400, 1497996000, 1497999600, 1498003200, 1498006800, 
    1498010400, 1498014000, 1498017600, 1498021200, 1498024800, 1498028400, 
    1498032000, 1498035600, 1498039200, 1498042800, 1498046400, 1498050000, 
    1498053600, 1498057200, 1498060800, 1498064400, 1498068000, 1498071600, 
    1498075200, 1498078800, 1498082400, 1498086000, 1498089600, 1498093200, 
    1498096800, 1498100400, 1498104000, 1498107600, 1498111200, 1498114800, 
    1498118400, 1498122000, 1498125600, 1498129200, 1498132800, 1498136400, 
    1498140000, 1498143600, 1498147200, 1498150800, 1498154400, 1498158000, 
    1498161600, 1498165200, 1498168800, 1498172400, 1498176000, 1498179600, 
    1498183200, 1498186800, 1498190400, 1498194000, 1498197600, 1498201200, 
    1498204800, 1498208400, 1498212000, 1498215600, 1498219200, 1498222800, 
    1498226400, 1498230000, 1498233600, 1498237200, 1498240800, 1498244400, 
    1498248000, 1498251600, 1498255200, 1498258800, 1498262400, 1498266000, 
    1498269600, 1498273200, 1498276800, 1498280400, 1498284000, 1498287600, 
    1498291200, 1498294800, 1498298400, 1498302000, 1498305600, 1498309200, 
    1498312800, 1498316400, 1498320000, 1498323600, 1498327200, 1498330800, 
    1498334400, 1498338000, 1498341600, 1498345200, 1498348800, 1498352400, 
    1498356000, 1498359600, 1498363200, 1498366800, 1498370400, 1498374000, 
    1498377600, 1498381200, 1498384800, 1498388400, 1498392000, 1498395600, 
    1498399200, 1498402800, 1498406400, 1498410000, 1498413600, 1498417200, 
    1498420800, 1498424400, 1498428000, 1498431600, 1498435200, 1498438800, 
    1498442400, 1498446000, 1498449600, 1498453200, 1498456800, 1498460400, 
    1498464000, 1498467600, 1498471200, 1498474800, 1498478400, 1498482000, 
    1498485600, 1498489200, 1498492800, 1498496400, 1498500000, 1498503600, 
    1498507200, 1498510800, 1498514400, 1498518000, 1498521600, 1498525200, 
    1498528800, 1498532400, 1498536000, 1498539600, 1498543200, 1498546800, 
    1498550400, 1498554000, 1498557600, 1498561200, 1498564800, 1498568400, 
    1498572000, 1498575600, 1498579200, 1498582800, 1498586400, 1498590000, 
    1498593600, 1498597200, 1498600800, 1498604400, 1498608000, 1498611600, 
    1498615200, 1498618800, 1498622400, 1498626000, 1498629600, 1498633200, 
    1498636800, 1498640400, 1498644000, 1498647600, 1498651200, 1498654800, 
    1498658400, 1498662000, 1498665600, 1498669200, 1498672800, 1498676400, 
    1498680000, 1498683600, 1498687200, 1498690800, 1498694400, 1498698000, 
    1498701600, 1498705200, 1498708800, 1498712400, 1498716000, 1498719600, 
    1498723200, 1498726800, 1498730400, 1498734000, 1498737600, 1498741200, 
    1498744800, 1498748400, 1498752000, 1498755600, 1498759200, 1498762800, 
    1498766400, 1498770000, 1498773600, 1498777200, 1498780800, 1498784400, 
    1498788000, 1498791600, 1498795200, 1498798800, 1498802400, 1498806000, 
    1498809600, 1498813200, 1498816800, 1498820400, 1498824000, 1498827600, 
    1498831200, 1498834800, 1498838400, 1498842000, 1498845600, 1498849200, 
    1498852800, 1498856400, 1498860000, 1498863600, 1498867200, 1498870800, 
    1498874400, 1498878000, 1498881600, 1498885200, 1498888800, 1498892400, 
    1498896000, 1498899600, 1498903200, 1498906800, 1498910400, 1498914000, 
    1498917600, 1498921200, 1498924800, 1498928400, 1498932000, 1498935600, 
    1498939200, 1498942800, 1498946400, 1498950000, 1498953600, 1498957200, 
    1498960800, 1498964400, 1498968000, 1498971600, 1498975200, 1498978800, 
    1498982400, 1498986000, 1498989600, 1498993200, 1498996800, 1499000400, 
    1499004000, 1499007600, 1499011200, 1499014800, 1499018400, 1499022000, 
    1499025600, 1499029200, 1499032800, 1499036400, 1499040000, 1499043600, 
    1499047200, 1499050800, 1499054400, 1499058000, 1499061600, 1499065200, 
    1499068800, 1499072400, 1499076000, 1499079600, 1499083200, 1499086800, 
    1499090400, 1499094000, 1499097600, 1499101200, 1499104800, 1499108400, 
    1499112000, 1499115600, 1499119200, 1499122800, 1499126400, 1499130000, 
    1499133600, 1499137200, 1499140800, 1499144400, 1499148000, 1499151600, 
    1499155200, 1499158800, 1499162400, 1499166000, 1499169600, 1499173200, 
    1499176800, 1499180400, 1499184000, 1499187600, 1499191200, 1499194800, 
    1499198400, 1499202000, 1499205600, 1499209200, 1499212800, 1499216400, 
    1499220000, 1499223600, 1499227200, 1499230800, 1499234400, 1499238000, 
    1499241600, 1499245200, 1499248800, 1499252400, 1499256000, 1499259600, 
    1499263200, 1499266800, 1499270400, 1499274000, 1499277600, 1499281200, 
    1499284800, 1499288400, 1499292000, 1499295600, 1499299200, 1499302800, 
    1499306400, 1499310000, 1499313600, 1499317200, 1499320800, 1499324400, 
    1499328000, 1499331600, 1499335200, 1499338800, 1499342400, 1499346000, 
    1499349600, 1499353200, 1499356800, 1499360400, 1499364000, 1499367600, 
    1499371200, 1499374800, 1499378400, 1499382000, 1499385600, 1499389200, 
    1499392800, 1499396400, 1499400000, 1499403600, 1499407200, 1499410800, 
    1499414400, 1499418000, 1499421600, 1499425200, 1499428800, 1499432400, 
    1499436000, 1499439600, 1499443200, 1499446800, 1499450400, 1499454000, 
    1499457600, 1499461200, 1499464800, 1499468400, 1499472000, 1499475600, 
    1499479200, 1499482800, 1499486400, 1499490000, 1499493600, 1499497200, 
    1499500800, 1499504400, 1499508000, 1499511600, 1499515200, 1499518800, 
    1499522400, 1499526000, 1499529600, 1499533200, 1499536800, 1499540400, 
    1499544000, 1499547600, 1499551200, 1499554800, 1499558400, 1499562000, 
    1499565600, 1499569200, 1499572800, 1499576400, 1499580000, 1499583600, 
    1499587200, 1499590800, 1499594400, 1499598000, 1499601600, 1499605200, 
    1499608800, 1499612400, 1499616000, 1499619600, 1499623200, 1499626800, 
    1499630400, 1499634000, 1499637600, 1499641200, 1499644800, 1499648400, 
    1499652000, 1499655600, 1499659200, 1499662800, 1499666400, 1499670000, 
    1499673600, 1499677200, 1499680800, 1499684400, 1499688000, 1499691600, 
    1499695200, 1499698800, 1499702400, 1499706000, 1499709600, 1499713200, 
    1499716800, 1499720400, 1499724000, 1499727600, 1499731200, 1499734800, 
    1499738400, 1499742000, 1499745600, 1499749200, 1499752800, 1499756400, 
    1499760000, 1499763600, 1499767200, 1499770800, 1499774400, 1499778000, 
    1499781600, 1499785200, 1499788800, 1499792400, 1499796000, 1499799600, 
    1499803200, 1499806800, 1499810400, 1499814000, 1499817600, 1499821200, 
    1499824800, 1499828400, 1499832000, 1499835600, 1499839200, 1499842800, 
    1499846400, 1499850000, 1499853600, 1499857200, 1499860800, 1499864400, 
    1499868000, 1499871600, 1499875200, 1499878800, 1499882400, 1499886000, 
    1499889600, 1499893200, 1499896800, 1499900400, 1499904000, 1499907600, 
    1499911200, 1499914800, 1499918400, 1499922000, 1499925600, 1499929200, 
    1499932800, 1499936400, 1499940000, 1499943600, 1499947200, 1499950800, 
    1499954400, 1499958000, 1499961600, 1499965200, 1499968800, 1499972400, 
    1499976000, 1499979600, 1499983200, 1499986800, 1499990400, 1499994000, 
    1499997600, 1500001200, 1500004800, 1500008400, 1500012000, 1500015600, 
    1500019200, 1500022800, 1500026400, 1500030000, 1500033600, 1500037200, 
    1500040800, 1500044400, 1500048000, 1500051600, 1500055200, 1500058800, 
    1500062400, 1500066000, 1500069600, 1500073200, 1500076800, 1500080400, 
    1500084000, 1500087600, 1500091200, 1500094800, 1500098400, 1500102000, 
    1500105600, 1500109200, 1500112800, 1500116400, 1500120000, 1500123600, 
    1500127200, 1500130800, 1500134400, 1500138000, 1500141600, 1500145200, 
    1500148800, 1500152400, 1500156000, 1500159600, 1500163200, 1500166800, 
    1500170400, 1500174000, 1500177600, 1500181200, 1500184800, 1500188400, 
    1500192000, 1500195600, 1500199200, 1500202800, 1500206400, 1500210000, 
    1500213600, 1500217200, 1500220800, 1500224400, 1500228000, 1500231600, 
    1500235200, 1500238800, 1500242400, 1500246000, 1500249600, 1500253200, 
    1500256800, 1500260400, 1500264000, 1500267600, 1500271200, 1500274800, 
    1500278400, 1500282000, 1500285600, 1500289200, 1500292800, 1500296400, 
    1500300000, 1500303600, 1500307200, 1500310800, 1500314400, 1500318000, 
    1500321600, 1500325200, 1500328800, 1500332400, 1500336000, 1500339600, 
    1500343200, 1500346800, 1500350400, 1500354000, 1500357600, 1500361200, 
    1500364800, 1500368400, 1500372000, 1500375600, 1500379200, 1500382800, 
    1500386400, 1500390000, 1500393600, 1500397200, 1500400800, 1500404400, 
    1500408000, 1500411600, 1500415200, 1500418800, 1500422400, 1500426000, 
    1500429600, 1500433200, 1500436800, 1500440400, 1500444000, 1500447600, 
    1500451200, 1500454800, 1500458400, 1500462000, 1500465600, 1500469200, 
    1500472800, 1500476400, 1500480000, 1500483600, 1500487200, 1500490800, 
    1500494400, 1500498000, 1500501600, 1500505200, 1500508800, 1500512400, 
    1500516000, 1500519600, 1500523200, 1500526800, 1500530400, 1500534000, 
    1500537600, 1500541200, 1500544800, 1500548400, 1500552000, 1500555600, 
    1500559200, 1500562800, 1500566400, 1500570000, 1500573600, 1500577200, 
    1500580800, 1500584400, 1500588000, 1500591600, 1500595200, 1500598800, 
    1500602400, 1500606000, 1500609600, 1500613200, 1500616800, 1500620400, 
    1500624000, 1500627600, 1500631200, 1500634800, 1500638400, 1500642000, 
    1500645600, 1500649200, 1500652800, 1500656400, 1500660000, 1500663600, 
    1500667200, 1500670800, 1500674400, 1500678000, 1500681600, 1500685200, 
    1500688800, 1500692400, 1500696000, 1500699600, 1500703200, 1500706800, 
    1500710400, 1500714000, 1500717600, 1500721200, 1500724800, 1500728400, 
    1500732000, 1500735600, 1500739200, 1500742800, 1500746400, 1500750000, 
    1500753600, 1500757200, 1500760800, 1500764400, 1500768000, 1500771600, 
    1500775200, 1500778800, 1500782400, 1500786000, 1500789600, 1500793200, 
    1500796800, 1500800400, 1500804000, 1500807600, 1500811200, 1500814800, 
    1500818400, 1500822000, 1500825600, 1500829200, 1500832800, 1500836400, 
    1500840000, 1500843600, 1500847200, 1500850800, 1500854400, 1500858000, 
    1500861600, 1500865200, 1500868800, 1500872400, 1500876000, 1500879600, 
    1500883200, 1500886800, 1500890400, 1500894000, 1500897600, 1500901200, 
    1500904800, 1500908400, 1500912000, 1500915600, 1500919200, 1500922800, 
    1500926400, 1500930000, 1500933600, 1500937200, 1500940800, 1500944400, 
    1500948000, 1500951600, 1500955200, 1500958800, 1500962400, 1500966000, 
    1500969600, 1500973200, 1500976800, 1500980400, 1500984000, 1500987600, 
    1500991200, 1500994800, 1500998400, 1501002000, 1501005600, 1501009200, 
    1501012800, 1501016400, 1501020000, 1501023600, 1501027200, 1501030800, 
    1501034400, 1501038000, 1501041600, 1501045200, 1501048800, 1501052400, 
    1501056000, 1501059600, 1501063200, 1501066800, 1501070400, 1501074000, 
    1501077600, 1501081200, 1501084800, 1501088400, 1501092000, 1501095600, 
    1501099200, 1501102800, 1501106400, 1501110000, 1501113600, 1501117200, 
    1501120800, 1501124400, 1501128000, 1501131600, 1501135200, 1501138800, 
    1501142400, 1501146000, 1501149600, 1501153200, 1501156800, 1501160400, 
    1501164000, 1501167600, 1501171200, 1501174800, 1501178400, 1501182000, 
    1501185600, 1501189200, 1501192800, 1501196400, 1501200000, 1501203600, 
    1501207200, 1501210800, 1501214400, 1501218000, 1501221600, 1501225200, 
    1501228800, 1501232400, 1501236000, 1501239600, 1501243200, 1501246800, 
    1501250400, 1501254000, 1501257600, 1501261200, 1501264800, 1501268400, 
    1501272000, 1501275600, 1501279200, 1501282800, 1501286400, 1501290000, 
    1501293600, 1501297200, 1501300800, 1501304400, 1501308000, 1501311600, 
    1501315200, 1501318800, 1501322400, 1501326000, 1501329600, 1501333200, 
    1501336800, 1501340400, 1501344000, 1501347600, 1501351200, 1501354800, 
    1501358400, 1501362000, 1501365600, 1501369200, 1501372800, 1501376400, 
    1501380000, 1501383600, 1501387200, 1501390800, 1501394400, 1501398000, 
    1501401600, 1501405200, 1501408800, 1501412400, 1501416000, 1501419600, 
    1501423200, 1501426800, 1501430400, 1501434000, 1501437600, 1501441200, 
    1501444800, 1501448400, 1501452000, 1501455600, 1501459200, 1501462800, 
    1501466400, 1501470000, 1501473600, 1501477200, 1501480800, 1501484400, 
    1501488000, 1501491600, 1501495200, 1501498800, 1501502400, 1501506000, 
    1501509600, 1501513200, 1501516800, 1501520400, 1501524000, 1501527600, 
    1501531200, 1501534800, 1501538400, 1501542000, 1501545600, 1501549200, 
    1501552800, 1501556400, 1501560000, 1501563600, 1501567200, 1501570800, 
    1501574400, 1501578000, 1501581600, 1501585200, 1501588800, 1501592400, 
    1501596000, 1501599600, 1501603200, 1501606800, 1501610400, 1501614000, 
    1501617600, 1501621200, 1501624800, 1501628400, 1501632000, 1501635600, 
    1501639200, 1501642800, 1501646400, 1501650000, 1501653600, 1501657200, 
    1501660800, 1501664400, 1501668000, 1501671600, 1501675200, 1501678800, 
    1501682400, 1501686000, 1501689600, 1501693200, 1501696800, 1501700400, 
    1501704000, 1501707600, 1501711200, 1501714800, 1501718400, 1501722000, 
    1501725600, 1501729200, 1501732800, 1501736400, 1501740000, 1501743600, 
    1501747200, 1501750800, 1501754400, 1501758000, 1501761600, 1501765200, 
    1501768800, 1501772400, 1501776000, 1501779600, 1501783200, 1501786800, 
    1501790400, 1501794000, 1501797600, 1501801200, 1501804800, 1501808400, 
    1501812000, 1501815600, 1501819200, 1501822800, 1501826400, 1501830000, 
    1501833600, 1501837200, 1501840800, 1501844400, 1501848000, 1501851600, 
    1501855200, 1501858800, 1501862400, 1501866000, 1501869600, 1501873200, 
    1501876800, 1501880400, 1501884000, 1501887600, 1501891200, 1501894800, 
    1501898400, 1501902000, 1501905600, 1501909200, 1501912800, 1501916400, 
    1501920000, 1501923600, 1501927200, 1501930800, 1501934400, 1501938000, 
    1501941600, 1501945200, 1501948800, 1501952400, 1501956000, 1501959600, 
    1501963200, 1501966800, 1501970400, 1501974000, 1501977600, 1501981200, 
    1501984800, 1501988400, 1501992000, 1501995600, 1501999200, 1502002800, 
    1502006400, 1502010000, 1502013600, 1502017200, 1502020800, 1502024400, 
    1502028000, 1502031600, 1502035200, 1502038800, 1502042400, 1502046000, 
    1502049600, 1502053200, 1502056800, 1502060400, 1502064000, 1502067600, 
    1502071200, 1502074800, 1502078400, 1502082000, 1502085600, 1502089200, 
    1502092800, 1502096400, 1502100000, 1502103600, 1502107200, 1502110800, 
    1502114400, 1502118000, 1502121600, 1502125200, 1502128800, 1502132400, 
    1502136000, 1502139600, 1502143200, 1502146800, 1502150400, 1502154000, 
    1502157600, 1502161200, 1502164800, 1502168400, 1502172000, 1502175600, 
    1502179200, 1502182800, 1502186400, 1502190000, 1502193600, 1502197200, 
    1502200800, 1502204400, 1502208000, 1502211600, 1502215200, 1502218800, 
    1502222400, 1502226000, 1502229600, 1502233200, 1502236800, 1502240400, 
    1502244000, 1502247600, 1502251200, 1502254800, 1502258400, 1502262000, 
    1502265600, 1502269200, 1502272800, 1502276400, 1502280000, 1502283600, 
    1502287200, 1502290800, 1502294400, 1502298000, 1502301600, 1502305200, 
    1502308800, 1502312400, 1502316000, 1502319600, 1502323200, 1502326800, 
    1502330400, 1502334000, 1502337600, 1502341200, 1502344800, 1502348400, 
    1502352000, 1502355600, 1502359200, 1502362800, 1502366400, 1502370000, 
    1502373600, 1502377200, 1502380800, 1502384400, 1502388000, 1502391600, 
    1502395200, 1502398800, 1502402400, 1502406000, 1502409600, 1502413200, 
    1502416800, 1502420400, 1502424000, 1502427600, 1502431200, 1502434800, 
    1502438400, 1502442000, 1502445600, 1502449200, 1502452800, 1502456400, 
    1502460000, 1502463600, 1502467200, 1502470800, 1502474400, 1502478000, 
    1502481600, 1502485200, 1502488800, 1502492400, 1502496000, 1502499600, 
    1502503200, 1502506800, 1502510400, 1502514000, 1502517600, 1502521200, 
    1502524800, 1502528400, 1502532000, 1502535600, 1502539200, 1502542800, 
    1502546400, 1502550000, 1502553600, 1502557200, 1502560800, 1502564400, 
    1502568000, 1502571600, 1502575200, 1502578800, 1502582400, 1502586000, 
    1502589600, 1502593200, 1502596800, 1502600400, 1502604000, 1502607600, 
    1502611200, 1502614800, 1502618400, 1502622000, 1502625600, 1502629200, 
    1502632800, 1502636400, 1502640000, 1502643600, 1502647200, 1502650800, 
    1502654400, 1502658000, 1502661600, 1502665200, 1502668800, 1502672400, 
    1502676000, 1502679600, 1502683200, 1502686800, 1502690400, 1502694000, 
    1502697600, 1502701200, 1502704800, 1502708400, 1502712000, 1502715600, 
    1502719200, 1502722800, 1502726400, 1502730000, 1502733600, 1502737200, 
    1502740800, 1502744400, 1502748000, 1502751600, 1502755200, 1502758800, 
    1502762400, 1502766000, 1502769600, 1502773200, 1502776800, 1502780400, 
    1502784000, 1502787600, 1502791200, 1502794800, 1502798400, 1502802000, 
    1502805600, 1502809200, 1502812800, 1502816400, 1502820000, 1502823600, 
    1502827200, 1502830800, 1502834400, 1502838000, 1502841600, 1502845200, 
    1502848800, 1502852400, 1502856000, 1502859600, 1502863200, 1502866800, 
    1502870400, 1502874000, 1502877600, 1502881200, 1502884800, 1502888400, 
    1502892000, 1502895600, 1502899200, 1502902800, 1502906400, 1502910000, 
    1502913600, 1502917200, 1502920800, 1502924400, 1502928000, 1502931600, 
    1502935200, 1502938800, 1502942400, 1502946000, 1502949600, 1502953200, 
    1502956800, 1502960400, 1502964000, 1502967600, 1502971200, 1502974800, 
    1502978400, 1502982000, 1502985600, 1502989200, 1502992800, 1502996400, 
    1503000000, 1503003600, 1503007200, 1503010800, 1503014400, 1503018000, 
    1503021600, 1503025200, 1503028800, 1503032400, 1503036000, 1503039600, 
    1503043200, 1503046800, 1503050400, 1503054000, 1503057600, 1503061200, 
    1503064800, 1503068400, 1503072000, 1503075600, 1503079200, 1503082800, 
    1503086400, 1503090000, 1503093600, 1503097200, 1503100800, 1503104400, 
    1503108000, 1503111600, 1503115200, 1503118800, 1503122400, 1503126000, 
    1503129600, 1503133200, 1503136800, 1503140400, 1503144000, 1503147600, 
    1503151200, 1503154800, 1503158400, 1503162000, 1503165600, 1503169200, 
    1503172800, 1503176400, 1503180000, 1503183600, 1503187200, 1503190800, 
    1503194400, 1503198000, 1503201600, 1503205200, 1503208800, 1503212400, 
    1503216000, 1503219600, 1503223200, 1503226800, 1503230400, 1503234000, 
    1503237600, 1503241200, 1503244800, 1503248400, 1503252000, 1503255600, 
    1503259200, 1503262800, 1503266400, 1503270000, 1503273600, 1503277200, 
    1503280800, 1503284400, 1503288000, 1503291600, 1503295200, 1503298800, 
    1503302400, 1503306000, 1503309600, 1503313200, 1503316800, 1503320400, 
    1503324000, 1503327600, 1503331200, 1503334800, 1503338400, 1503342000, 
    1503345600, 1503349200, 1503352800, 1503356400, 1503360000, 1503363600, 
    1503367200, 1503370800, 1503374400, 1503378000, 1503381600, 1503385200, 
    1503388800, 1503392400, 1503396000, 1503399600, 1503403200, 1503406800, 
    1503410400, 1503414000, 1503417600, 1503421200, 1503424800, 1503428400, 
    1503432000, 1503435600, 1503439200, 1503442800, 1503446400, 1503450000, 
    1503453600, 1503457200, 1503460800, 1503464400, 1503468000, 1503471600, 
    1503475200, 1503478800, 1503482400, 1503486000, 1503489600, 1503493200, 
    1503496800, 1503500400, 1503504000, 1503507600, 1503511200, 1503514800, 
    1503518400, 1503522000, 1503525600, 1503529200, 1503532800, 1503536400, 
    1503540000, 1503543600, 1503547200, 1503550800, 1503554400, 1503558000, 
    1503561600, 1503565200, 1503568800, 1503572400, 1503576000, 1503579600, 
    1503583200, 1503586800, 1503590400, 1503594000, 1503597600, 1503601200, 
    1503604800, 1503608400, 1503612000, 1503615600, 1503619200, 1503622800, 
    1503626400, 1503630000, 1503633600, 1503637200, 1503640800, 1503644400, 
    1503648000, 1503651600, 1503655200, 1503658800, 1503662400, 1503666000, 
    1503669600, 1503673200, 1503676800, 1503680400, 1503684000, 1503687600, 
    1503691200, 1503694800, 1503698400, 1503702000, 1503705600, 1503709200, 
    1503712800, 1503716400, 1503720000, 1503723600, 1503727200, 1503730800, 
    1503734400, 1503738000, 1503741600, 1503745200, 1503748800, 1503752400, 
    1503756000, 1503759600, 1503763200, 1503766800, 1503770400, 1503774000, 
    1503777600, 1503781200, 1503784800, 1503788400, 1503792000, 1503795600, 
    1503799200, 1503802800, 1503806400, 1503810000, 1503813600, 1503817200, 
    1503820800, 1503824400, 1503828000, 1503831600, 1503835200, 1503838800, 
    1503842400, 1503846000, 1503849600, 1503853200, 1503856800, 1503860400, 
    1503864000, 1503867600, 1503871200, 1503874800, 1503878400, 1503882000, 
    1503885600, 1503889200, 1503892800, 1503896400, 1503900000, 1503903600, 
    1503907200, 1503910800, 1503914400, 1503918000, 1503921600, 1503925200, 
    1503928800, 1503932400, 1503936000, 1503939600, 1503943200, 1503946800, 
    1503950400, 1503954000, 1503957600, 1503961200, 1503964800, 1503968400, 
    1503972000, 1503975600, 1503979200, 1503982800, 1503986400, 1503990000, 
    1503993600, 1503997200, 1504000800, 1504004400, 1504008000, 1504011600, 
    1504015200, 1504018800, 1504022400, 1504026000, 1504029600, 1504033200, 
    1504036800, 1504040400, 1504044000, 1504047600, 1504051200, 1504054800, 
    1504058400, 1504062000, 1504065600, 1504069200, 1504072800, 1504076400, 
    1504080000, 1504083600, 1504087200, 1504090800, 1504094400, 1504098000, 
    1504101600, 1504105200, 1504108800, 1504112400, 1504116000, 1504119600, 
    1504123200, 1504126800, 1504130400, 1504134000, 1504137600, 1504141200, 
    1504144800, 1504148400, 1504152000, 1504155600, 1504159200, 1504162800, 
    1504166400, 1504170000, 1504173600, 1504177200, 1504180800, 1504184400, 
    1504188000, 1504191600, 1504195200, 1504198800, 1504202400, 1504206000, 
    1504209600, 1504213200, 1504216800, 1504220400, 1504224000, 1504227600, 
    1504231200, 1504234800, 1504238400, 1504242000, 1504245600, 1504249200, 
    1504252800, 1504256400, 1504260000, 1504263600, 1504267200, 1504270800, 
    1504274400, 1504278000, 1504281600, 1504285200, 1504288800, 1504292400, 
    1504296000, 1504299600, 1504303200, 1504306800, 1504310400, 1504314000, 
    1504317600, 1504321200, 1504324800, 1504328400, 1504332000, 1504335600, 
    1504339200, 1504342800, 1504346400, 1504350000, 1504353600, 1504357200, 
    1504360800, 1504364400, 1504368000, 1504371600, 1504375200, 1504378800, 
    1504382400, 1504386000, 1504389600, 1504393200, 1504396800, 1504400400, 
    1504404000, 1504407600, 1504411200, 1504414800, 1504418400, 1504422000, 
    1504425600, 1504429200, 1504432800, 1504436400, 1504440000, 1504443600, 
    1504447200, 1504450800, 1504454400, 1504458000, 1504461600, 1504465200, 
    1504468800, 1504472400, 1504476000, 1504479600, 1504483200, 1504486800, 
    1504490400, 1504494000, 1504497600, 1504501200, 1504504800, 1504508400, 
    1504512000, 1504515600, 1504519200, 1504522800, 1504526400, 1504530000, 
    1504533600, 1504537200, 1504540800, 1504544400, 1504548000, 1504551600, 
    1504555200, 1504558800, 1504562400, 1504566000, 1504569600, 1504573200, 
    1504576800, 1504580400, 1504584000, 1504587600, 1504591200, 1504594800, 
    1504598400, 1504602000, 1504605600, 1504609200, 1504612800, 1504616400, 
    1504620000, 1504623600, 1504627200, 1504630800, 1504634400, 1504638000, 
    1504641600, 1504645200, 1504648800, 1504652400, 1504656000, 1504659600, 
    1504663200, 1504666800, 1504670400, 1504674000, 1504677600, 1504681200, 
    1504684800, 1504688400, 1504692000, 1504695600, 1504699200, 1504702800, 
    1504706400, 1504710000, 1504713600, 1504717200, 1504720800, 1504724400, 
    1504728000, 1504731600, 1504735200, 1504738800, 1504742400, 1504746000, 
    1504749600, 1504753200, 1504756800, 1504760400, 1504764000, 1504767600, 
    1504771200, 1504774800, 1504778400, 1504782000, 1504785600, 1504789200, 
    1504792800, 1504796400, 1504800000, 1504803600, 1504807200, 1504810800, 
    1504814400, 1504818000, 1504821600, 1504825200, 1504828800, 1504832400, 
    1504836000, 1504839600, 1504843200, 1504846800, 1504850400, 1504854000, 
    1504857600, 1504861200, 1504864800, 1504868400, 1504872000, 1504875600, 
    1504879200, 1504882800, 1504886400, 1504890000, 1504893600, 1504897200, 
    1504900800, 1504904400, 1504908000, 1504911600, 1504915200, 1504918800, 
    1504922400, 1504926000, 1504929600, 1504933200, 1504936800, 1504940400, 
    1504944000, 1504947600, 1504951200, 1504954800, 1504958400, 1504962000, 
    1504965600, 1504969200, 1504972800, 1504976400, 1504980000, 1504983600, 
    1504987200, 1504990800, 1504994400, 1504998000, 1505001600, 1505005200, 
    1505008800, 1505012400, 1505016000, 1505019600, 1505023200, 1505026800, 
    1505030400, 1505034000, 1505037600, 1505041200, 1505044800, 1505048400, 
    1505052000, 1505055600, 1505059200, 1505062800, 1505066400, 1505070000, 
    1505073600, 1505077200, 1505080800, 1505084400, 1505088000, 1505091600, 
    1505095200, 1505098800, 1505102400, 1505106000, 1505109600, 1505113200, 
    1505116800, 1505120400, 1505124000, 1505127600, 1505131200, 1505134800, 
    1505138400, 1505142000, 1505145600, 1505149200, 1505152800, 1505156400, 
    1505160000, 1505163600, 1505167200, 1505170800, 1505174400, 1505178000, 
    1505181600, 1505185200, 1505188800, 1505192400, 1505196000, 1505199600, 
    1505203200, 1505206800, 1505210400, 1505214000, 1505217600, 1505221200, 
    1505224800, 1505228400, 1505232000, 1505235600, 1505239200, 1505242800, 
    1505246400, 1505250000, 1505253600, 1505257200, 1505260800, 1505264400, 
    1505268000, 1505271600, 1505275200, 1505278800, 1505282400, 1505286000, 
    1505289600, 1505293200, 1505296800, 1505300400, 1505304000, 1505307600, 
    1505311200, 1505314800, 1505318400, 1505322000, 1505325600, 1505329200, 
    1505332800, 1505336400, 1505340000, 1505343600, 1505347200, 1505350800, 
    1505354400, 1505358000, 1505361600, 1505365200, 1505368800, 1505372400, 
    1505376000, 1505379600, 1505383200, 1505386800, 1505390400, 1505394000, 
    1505397600, 1505401200, 1505404800, 1505408400, 1505412000, 1505415600, 
    1505419200, 1505422800, 1505426400, 1505430000, 1505433600, 1505437200, 
    1505440800, 1505444400, 1505448000, 1505451600, 1505455200, 1505458800, 
    1505462400, 1505466000, 1505469600, 1505473200, 1505476800, 1505480400, 
    1505484000, 1505487600, 1505491200, 1505494800, 1505498400, 1505502000, 
    1505505600, 1505509200, 1505512800, 1505516400, 1505520000, 1505523600, 
    1505527200, 1505530800, 1505534400, 1505538000, 1505541600, 1505545200, 
    1505548800, 1505552400, 1505556000, 1505559600, 1505563200, 1505566800, 
    1505570400, 1505574000, 1505577600, 1505581200, 1505584800, 1505588400, 
    1505592000, 1505595600, 1505599200, 1505602800, 1505606400, 1505610000, 
    1505613600, 1505617200, 1505620800, 1505624400, 1505628000, 1505631600, 
    1505635200, 1505638800, 1505642400, 1505646000, 1505649600, 1505653200, 
    1505656800, 1505660400, 1505664000, 1505667600, 1505671200, 1505674800, 
    1505678400, 1505682000, 1505685600, 1505689200, 1505692800, 1505696400, 
    1505700000, 1505703600, 1505707200, 1505710800, 1505714400, 1505718000, 
    1505721600, 1505725200, 1505728800, 1505732400, 1505736000, 1505739600, 
    1505743200, 1505746800, 1505750400, 1505754000, 1505757600, 1505761200, 
    1505764800, 1505768400, 1505772000, 1505775600, 1505779200, 1505782800, 
    1505786400, 1505790000, 1505793600, 1505797200, 1505800800, 1505804400, 
    1505808000, 1505811600, 1505815200, 1505818800, 1505822400, 1505826000, 
    1505829600, 1505833200, 1505836800, 1505840400, 1505844000, 1505847600, 
    1505851200, 1505854800, 1505858400, 1505862000, 1505865600, 1505869200, 
    1505872800, 1505876400, 1505880000, 1505883600, 1505887200, 1505890800, 
    1505894400, 1505898000, 1505901600, 1505905200, 1505908800, 1505912400, 
    1505916000, 1505919600, 1505923200, 1505926800, 1505930400, 1505934000, 
    1505937600, 1505941200, 1505944800, 1505948400, 1505952000, 1505955600, 
    1505959200, 1505962800, 1505966400, 1505970000, 1505973600, 1505977200, 
    1505980800, 1505984400, 1505988000, 1505991600, 1505995200, 1505998800, 
    1506002400, 1506006000, 1506009600, 1506013200, 1506016800, 1506020400, 
    1506024000, 1506027600, 1506031200, 1506034800, 1506038400, 1506042000, 
    1506045600, 1506049200, 1506052800, 1506056400, 1506060000, 1506063600, 
    1506067200, 1506070800, 1506074400, 1506078000, 1506081600, 1506085200, 
    1506088800, 1506092400, 1506096000, 1506099600, 1506103200, 1506106800, 
    1506110400, 1506114000, 1506117600, 1506121200, 1506124800, 1506128400, 
    1506132000, 1506135600, 1506139200, 1506142800, 1506146400, 1506150000, 
    1506153600, 1506157200, 1506160800, 1506164400, 1506168000, 1506171600, 
    1506175200, 1506178800, 1506182400, 1506186000, 1506189600, 1506193200, 
    1506196800, 1506200400, 1506204000, 1506207600, 1506211200, 1506214800, 
    1506218400, 1506222000, 1506225600, 1506229200, 1506232800, 1506236400, 
    1506240000, 1506243600, 1506247200, 1506250800, 1506254400, 1506258000, 
    1506261600, 1506265200, 1506268800, 1506272400, 1506276000, 1506279600, 
    1506283200, 1506286800, 1506290400, 1506294000, 1506297600, 1506301200, 
    1506304800, 1506308400, 1506312000, 1506315600, 1506319200, 1506322800, 
    1506326400, 1506330000, 1506333600, 1506337200, 1506340800, 1506344400, 
    1506348000, 1506351600, 1506355200, 1506358800, 1506362400, 1506366000, 
    1506369600, 1506373200, 1506376800, 1506380400, 1506384000, 1506387600, 
    1506391200, 1506394800, 1506398400, 1506402000, 1506405600, 1506409200, 
    1506412800, 1506416400, 1506420000, 1506423600, 1506427200, 1506430800, 
    1506434400, 1506438000, 1506441600, 1506445200, 1506448800, 1506452400, 
    1506456000, 1506459600, 1506463200, 1506466800, 1506470400, 1506474000, 
    1506477600, 1506481200, 1506484800, 1506488400, 1506492000, 1506495600, 
    1506499200, 1506502800, 1506506400, 1506510000, 1506513600, 1506517200, 
    1506520800, 1506524400, 1506528000, 1506531600, 1506535200, 1506538800, 
    1506542400, 1506546000, 1506549600, 1506553200, 1506556800, 1506560400, 
    1506564000, 1506567600, 1506571200, 1506574800, 1506578400, 1506582000, 
    1506585600, 1506589200, 1506592800, 1506596400, 1506600000, 1506603600, 
    1506607200, 1506610800, 1506614400, 1506618000, 1506621600, 1506625200, 
    1506628800, 1506632400, 1506636000, 1506639600, 1506643200, 1506646800, 
    1506650400, 1506654000, 1506657600, 1506661200, 1506664800, 1506668400, 
    1506672000, 1506675600, 1506679200, 1506682800, 1506686400, 1506690000, 
    1506693600, 1506697200, 1506700800, 1506704400, 1506708000, 1506711600, 
    1506715200, 1506718800, 1506722400, 1506726000, 1506729600, 1506733200, 
    1506736800, 1506740400, 1506744000, 1506747600, 1506751200, 1506754800, 
    1506758400, 1506762000, 1506765600, 1506769200, 1506772800, 1506776400, 
    1506780000, 1506783600, 1506787200, 1506790800, 1506794400, 1506798000, 
    1506801600, 1506805200, 1506808800, 1506812400, 1506816000, 1506819600, 
    1506823200, 1506826800, 1506830400, 1506834000, 1506837600, 1506841200, 
    1506844800, 1506848400, 1506852000, 1506855600, 1506859200, 1506862800, 
    1506866400, 1506870000, 1506873600, 1506877200, 1506880800, 1506884400, 
    1506888000, 1506891600, 1506895200, 1506898800, 1506902400, 1506906000, 
    1506909600, 1506913200, 1506916800, 1506920400, 1506924000, 1506927600, 
    1506931200, 1506934800, 1506938400, 1506942000, 1506945600, 1506949200, 
    1506952800, 1506956400, 1506960000, 1506963600, 1506967200, 1506970800, 
    1506974400, 1506978000, 1506981600, 1506985200, 1506988800, 1506992400, 
    1506996000, 1506999600, 1507003200, 1507006800, 1507010400, 1507014000, 
    1507017600, 1507021200, 1507024800, 1507028400, 1507032000, 1507035600, 
    1507039200, 1507042800, 1507046400, 1507050000, 1507053600, 1507057200, 
    1507060800, 1507064400, 1507068000, 1507071600, 1507075200, 1507078800, 
    1507082400, 1507086000, 1507089600, 1507093200, 1507096800, 1507100400, 
    1507104000, 1507107600, 1507111200, 1507114800, 1507118400, 1507122000, 
    1507125600, 1507129200, 1507132800, 1507136400, 1507140000, 1507143600, 
    1507147200, 1507150800, 1507154400, 1507158000, 1507161600, 1507165200, 
    1507168800, 1507172400, 1507176000, 1507179600, 1507183200, 1507186800, 
    1507190400, 1507194000, 1507197600, 1507201200, 1507204800, 1507208400, 
    1507212000, 1507215600, 1507219200, 1507222800, 1507226400, 1507230000, 
    1507233600, 1507237200, 1507240800, 1507244400, 1507248000, 1507251600, 
    1507255200, 1507258800, 1507262400, 1507266000, 1507269600, 1507273200, 
    1507276800, 1507280400, 1507284000, 1507287600, 1507291200, 1507294800, 
    1507298400, 1507302000, 1507305600, 1507309200, 1507312800, 1507316400, 
    1507320000, 1507323600, 1507327200, 1507330800, 1507334400, 1507338000, 
    1507341600, 1507345200, 1507348800, 1507352400, 1507356000, 1507359600, 
    1507363200, 1507366800, 1507370400, 1507374000, 1507377600, 1507381200, 
    1507384800, 1507388400, 1507392000, 1507395600, 1507399200, 1507402800, 
    1507406400, 1507410000, 1507413600, 1507417200, 1507420800, 1507424400, 
    1507428000, 1507431600, 1507435200, 1507438800, 1507442400, 1507446000, 
    1507449600, 1507453200, 1507456800, 1507460400, 1507464000, 1507467600, 
    1507471200, 1507474800, 1507478400, 1507482000, 1507485600, 1507489200, 
    1507492800, 1507496400, 1507500000, 1507503600, 1507507200, 1507510800, 
    1507514400, 1507518000, 1507521600, 1507525200, 1507528800, 1507532400, 
    1507536000, 1507539600, 1507543200, 1507546800, 1507550400, 1507554000, 
    1507557600, 1507561200, 1507564800, 1507568400, 1507572000, 1507575600, 
    1507579200, 1507582800, 1507586400, 1507590000, 1507593600, 1507597200, 
    1507600800, 1507604400, 1507608000, 1507611600, 1507615200, 1507618800, 
    1507622400, 1507626000, 1507629600, 1507633200, 1507636800, 1507640400, 
    1507644000, 1507647600, 1507651200, 1507654800, 1507658400, 1507662000, 
    1507665600, 1507669200, 1507672800, 1507676400, 1507680000, 1507683600, 
    1507687200, 1507690800, 1507694400, 1507698000, 1507701600, 1507705200, 
    1507708800, 1507712400, 1507716000, 1507719600, 1507723200, 1507726800, 
    1507730400, 1507734000, 1507737600, 1507741200, 1507744800, 1507748400, 
    1507752000, 1507755600, 1507759200, 1507762800, 1507766400, 1507770000, 
    1507773600, 1507777200, 1507780800, 1507784400, 1507788000, 1507791600, 
    1507795200, 1507798800, 1507802400, 1507806000, 1507809600, 1507813200, 
    1507816800, 1507820400, 1507824000, 1507827600, 1507831200, 1507834800, 
    1507838400, 1507842000, 1507845600, 1507849200, 1507852800, 1507856400, 
    1507860000, 1507863600, 1507867200, 1507870800, 1507874400, 1507878000, 
    1507881600, 1507885200, 1507888800, 1507892400, 1507896000, 1507899600, 
    1507903200, 1507906800, 1507910400, 1507914000, 1507917600, 1507921200, 
    1507924800, 1507928400, 1507932000, 1507935600, 1507939200, 1507942800, 
    1507946400, 1507950000, 1507953600, 1507957200, 1507960800, 1507964400, 
    1507968000, 1507971600, 1507975200, 1507978800, 1507982400, 1507986000, 
    1507989600, 1507993200, 1507996800, 1508000400, 1508004000, 1508007600, 
    1508011200, 1508014800, 1508018400, 1508022000, 1508025600, 1508029200, 
    1508032800, 1508036400, 1508040000, 1508043600, 1508047200, 1508050800, 
    1508054400, 1508058000, 1508061600, 1508065200, 1508068800, 1508072400, 
    1508076000, 1508079600, 1508083200, 1508086800, 1508090400, 1508094000, 
    1508097600, 1508101200, 1508104800, 1508108400, 1508112000, 1508115600, 
    1508119200, 1508122800, 1508126400, 1508130000, 1508133600, 1508137200, 
    1508140800, 1508144400, 1508148000, 1508151600, 1508155200, 1508158800, 
    1508162400, 1508166000, 1508169600, 1508173200, 1508176800, 1508180400, 
    1508184000, 1508187600, 1508191200, 1508194800, 1508198400, 1508202000, 
    1508205600, 1508209200, 1508212800, 1508216400, 1508220000, 1508223600, 
    1508227200, 1508230800, 1508234400, 1508238000, 1508241600, 1508245200, 
    1508248800, 1508252400, 1508256000, 1508259600, 1508263200, 1508266800, 
    1508270400, 1508274000, 1508277600, 1508281200, 1508284800, 1508288400, 
    1508292000, 1508295600, 1508299200, 1508302800, 1508306400, 1508310000, 
    1508313600, 1508317200, 1508320800, 1508324400, 1508328000, 1508331600, 
    1508335200, 1508338800, 1508342400, 1508346000, 1508349600, 1508353200, 
    1508356800, 1508360400, 1508364000, 1508367600, 1508371200, 1508374800, 
    1508378400, 1508382000, 1508385600, 1508389200, 1508392800, 1508396400, 
    1508400000, 1508403600, 1508407200, 1508410800, 1508414400, 1508418000, 
    1508421600, 1508425200, 1508428800, 1508432400, 1508436000, 1508439600, 
    1508443200, 1508446800, 1508450400, 1508454000, 1508457600, 1508461200, 
    1508464800, 1508468400, 1508472000, 1508475600, 1508479200, 1508482800, 
    1508486400, 1508490000, 1508493600, 1508497200, 1508500800, 1508504400, 
    1508508000, 1508511600, 1508515200, 1508518800, 1508522400, 1508526000, 
    1508529600, 1508533200, 1508536800, 1508540400, 1508544000, 1508547600, 
    1508551200, 1508554800, 1508558400, 1508562000, 1508565600, 1508569200, 
    1508572800, 1508576400, 1508580000, 1508583600, 1508587200, 1508590800, 
    1508594400, 1508598000, 1508601600, 1508605200, 1508608800, 1508612400, 
    1508616000, 1508619600, 1508623200, 1508626800, 1508630400, 1508634000, 
    1508637600, 1508641200, 1508644800, 1508648400, 1508652000, 1508655600, 
    1508659200, 1508662800, 1508666400, 1508670000, 1508673600, 1508677200, 
    1508680800, 1508684400, 1508688000, 1508691600, 1508695200, 1508698800, 
    1508702400, 1508706000, 1508709600, 1508713200, 1508716800, 1508720400, 
    1508724000, 1508727600, 1508731200, 1508734800, 1508738400, 1508742000, 
    1508745600, 1508749200, 1508752800, 1508756400, 1508760000, 1508763600, 
    1508767200, 1508770800, 1508774400, 1508778000, 1508781600, 1508785200, 
    1508788800, 1508792400, 1508796000, 1508799600, 1508803200, 1508806800, 
    1508810400, 1508814000, 1508817600, 1508821200, 1508824800, 1508828400, 
    1508832000, 1508835600, 1508839200, 1508842800, 1508846400, 1508850000, 
    1508853600, 1508857200, 1508860800, 1508864400, 1508868000, 1508871600, 
    1508875200, 1508878800, 1508882400, 1508886000, 1508889600, 1508893200, 
    1508896800, 1508900400, 1508904000, 1508907600, 1508911200, 1508914800, 
    1508918400, 1508922000, 1508925600, 1508929200, 1508932800, 1508936400, 
    1508940000, 1508943600, 1508947200, 1508950800, 1508954400, 1508958000, 
    1508961600, 1508965200, 1508968800, 1508972400, 1508976000, 1508979600, 
    1508983200, 1508986800, 1508990400, 1508994000, 1508997600, 1509001200, 
    1509004800, 1509008400, 1509012000, 1509015600, 1509019200, 1509022800, 
    1509026400, 1509030000, 1509033600, 1509037200, 1509040800, 1509044400, 
    1509048000, 1509051600, 1509055200, 1509058800, 1509062400, 1509066000, 
    1509069600, 1509073200, 1509076800, 1509080400, 1509084000, 1509087600, 
    1509091200, 1509094800, 1509098400, 1509102000, 1509105600, 1509109200, 
    1509112800, 1509116400, 1509120000, 1509123600, 1509127200, 1509130800, 
    1509134400, 1509138000, 1509141600, 1509145200, 1509148800, 1509152400, 
    1509156000, 1509159600, 1509163200, 1509166800, 1509170400, 1509174000, 
    1509177600, 1509181200, 1509184800, 1509188400, 1509192000, 1509195600, 
    1509199200, 1509202800, 1509206400, 1509210000, 1509213600, 1509217200, 
    1509220800, 1509224400, 1509228000, 1509231600, 1509235200, 1509238800, 
    1509242400, 1509246000, 1509249600, 1509253200, 1509256800, 1509260400, 
    1509264000, 1509267600, 1509271200, 1509274800, 1509278400, 1509282000, 
    1509285600, 1509289200, 1509292800, 1509296400, 1509300000, 1509303600, 
    1509307200, 1509310800, 1509314400, 1509318000, 1509321600, 1509325200, 
    1509328800, 1509332400, 1509336000, 1509339600, 1509343200, 1509346800, 
    1509350400, 1509354000, 1509357600, 1509361200, 1509364800, 1509368400, 
    1509372000, 1509375600, 1509379200, 1509382800, 1509386400, 1509390000, 
    1509393600, 1509397200, 1509400800, 1509404400, 1509408000, 1509411600, 
    1509415200, 1509418800, 1509422400, 1509426000, 1509429600, 1509433200, 
    1509436800, 1509440400, 1509444000, 1509447600, 1509451200, 1509454800, 
    1509458400, 1509462000, 1509465600, 1509469200, 1509472800, 1509476400, 
    1509480000, 1509483600, 1509487200, 1509490800, 1509494400, 1509498000, 
    1509501600, 1509505200, 1509508800, 1509512400, 1509516000, 1509519600, 
    1509523200, 1509526800, 1509530400, 1509534000, 1509537600, 1509541200, 
    1509544800, 1509548400, 1509552000, 1509555600, 1509559200, 1509562800, 
    1509566400, 1509570000, 1509573600, 1509577200, 1509580800, 1509584400, 
    1509588000, 1509591600, 1509595200, 1509598800, 1509602400, 1509606000, 
    1509609600, 1509613200, 1509616800, 1509620400, 1509624000, 1509627600, 
    1509631200, 1509634800, 1509638400, 1509642000, 1509645600, 1509649200, 
    1509652800, 1509656400, 1509660000, 1509663600, 1509667200, 1509670800, 
    1509674400, 1509678000, 1509681600, 1509685200, 1509688800, 1509692400, 
    1509696000, 1509699600, 1509703200, 1509706800, 1509710400, 1509714000, 
    1509717600, 1509721200, 1509724800, 1509728400, 1509732000, 1509735600, 
    1509739200, 1509742800, 1509746400, 1509750000, 1509753600, 1509757200, 
    1509760800, 1509764400, 1509768000, 1509771600, 1509775200, 1509778800, 
    1509782400, 1509786000, 1509789600, 1509793200, 1509796800, 1509800400, 
    1509804000, 1509807600, 1509811200, 1509814800, 1509818400, 1509822000, 
    1509825600, 1509829200, 1509832800, 1509836400, 1509840000, 1509843600, 
    1509847200, 1509850800, 1509854400, 1509858000, 1509861600, 1509865200, 
    1509868800, 1509872400, 1509876000, 1509879600, 1509883200, 1509886800, 
    1509890400, 1509894000, 1509897600, 1509901200, 1509904800, 1509908400, 
    1509912000, 1509915600, 1509919200, 1509922800, 1509926400, 1509930000, 
    1509933600, 1509937200, 1509940800, 1509944400, 1509948000, 1509951600, 
    1509955200, 1509958800, 1509962400, 1509966000, 1509969600, 1509973200, 
    1509976800, 1509980400, 1509984000, 1509987600, 1509991200, 1509994800, 
    1509998400, 1510002000, 1510005600, 1510009200, 1510012800, 1510016400, 
    1510020000, 1510023600, 1510027200, 1510030800, 1510034400, 1510038000, 
    1510041600, 1510045200, 1510048800, 1510052400, 1510056000, 1510059600, 
    1510063200, 1510066800, 1510070400, 1510074000, 1510077600, 1510081200, 
    1510084800, 1510088400, 1510092000, 1510095600, 1510099200, 1510102800, 
    1510106400, 1510110000, 1510113600, 1510117200, 1510120800, 1510124400, 
    1510128000, 1510131600, 1510135200, 1510138800, 1510142400, 1510146000, 
    1510149600, 1510153200, 1510156800, 1510160400, 1510164000, 1510167600, 
    1510171200, 1510174800, 1510178400, 1510182000, 1510185600, 1510189200, 
    1510192800, 1510196400, 1510200000, 1510203600, 1510207200, 1510210800, 
    1510214400, 1510218000, 1510221600, 1510225200, 1510228800, 1510232400, 
    1510236000, 1510239600, 1510243200, 1510246800, 1510250400, 1510254000, 
    1510257600, 1510261200, 1510264800, 1510268400, 1510272000, 1510275600, 
    1510279200, 1510282800, 1510286400, 1510290000, 1510293600, 1510297200, 
    1510300800, 1510304400, 1510308000, 1510311600, 1510315200, 1510318800, 
    1510322400, 1510326000, 1510329600, 1510333200, 1510336800, 1510340400, 
    1510344000, 1510347600, 1510351200, 1510354800, 1510358400, 1510362000, 
    1510365600, 1510369200, 1510372800, 1510376400, 1510380000, 1510383600, 
    1510387200, 1510390800, 1510394400, 1510398000, 1510401600, 1510405200, 
    1510408800, 1510412400, 1510416000, 1510419600, 1510423200, 1510426800, 
    1510430400, 1510434000, 1510437600, 1510441200, 1510444800, 1510448400, 
    1510452000, 1510455600, 1510459200, 1510462800, 1510466400, 1510470000, 
    1510473600, 1510477200, 1510480800, 1510484400, 1510488000, 1510491600, 
    1510495200, 1510498800, 1510502400, 1510506000, 1510509600, 1510513200, 
    1510516800, 1510520400, 1510524000, 1510527600, 1510531200, 1510534800, 
    1510538400, 1510542000, 1510545600, 1510549200, 1510552800, 1510556400, 
    1510560000, 1510563600, 1510567200, 1510570800, 1510574400, 1510578000, 
    1510581600, 1510585200, 1510588800, 1510592400, 1510596000, 1510599600, 
    1510603200, 1510606800, 1510610400, 1510614000, 1510617600, 1510621200, 
    1510624800, 1510628400, 1510632000, 1510635600, 1510639200, 1510642800, 
    1510646400, 1510650000, 1510653600, 1510657200, 1510660800, 1510664400, 
    1510668000, 1510671600, 1510675200, 1510678800, 1510682400, 1510686000, 
    1510689600, 1510693200, 1510696800, 1510700400, 1510704000, 1510707600, 
    1510711200, 1510714800, 1510718400, 1510722000, 1510725600, 1510729200, 
    1510732800, 1510736400, 1510740000, 1510743600, 1510747200, 1510750800, 
    1510754400, 1510758000, 1510761600, 1510765200, 1510768800, 1510772400, 
    1510776000, 1510779600, 1510783200, 1510786800, 1510790400, 1510794000, 
    1510797600, 1510801200, 1510804800, 1510808400, 1510812000, 1510815600, 
    1510819200, 1510822800, 1510826400, 1510830000, 1510833600, 1510837200, 
    1510840800, 1510844400, 1510848000, 1510851600, 1510855200, 1510858800, 
    1510862400, 1510866000, 1510869600, 1510873200, 1510876800, 1510880400, 
    1510884000, 1510887600, 1510891200, 1510894800, 1510898400, 1510902000, 
    1510905600, 1510909200, 1510912800, 1510916400, 1510920000, 1510923600, 
    1510927200, 1510930800, 1510934400, 1510938000, 1510941600, 1510945200, 
    1510948800, 1510952400, 1510956000, 1510959600, 1510963200, 1510966800, 
    1510970400, 1510974000, 1510977600, 1510981200, 1510984800, 1510988400, 
    1510992000, 1510995600, 1510999200, 1511002800, 1511006400, 1511010000, 
    1511013600, 1511017200, 1511020800, 1511024400, 1511028000, 1511031600, 
    1511035200, 1511038800, 1511042400, 1511046000, 1511049600, 1511053200, 
    1511056800, 1511060400, 1511064000, 1511067600, 1511071200, 1511074800, 
    1511078400, 1511082000, 1511085600, 1511089200, 1511092800, 1511096400, 
    1511100000, 1511103600, 1511107200, 1511110800, 1511114400, 1511118000, 
    1511121600, 1511125200, 1511128800, 1511132400, 1511136000, 1511139600, 
    1511143200, 1511146800, 1511150400, 1511154000, 1511157600, 1511161200, 
    1511164800, 1511168400, 1511172000, 1511175600, 1511179200, 1511182800, 
    1511186400, 1511190000, 1511193600, 1511197200, 1511200800, 1511204400, 
    1511208000, 1511211600, 1511215200, 1511218800, 1511222400, 1511226000, 
    1511229600, 1511233200, 1511236800, 1511240400, 1511244000, 1511247600, 
    1511251200, 1511254800, 1511258400, 1511262000, 1511265600, 1511269200, 
    1511272800, 1511276400, 1511280000, 1511283600, 1511287200, 1511290800, 
    1511294400, 1511298000, 1511301600, 1511305200, 1511308800, 1511312400, 
    1511316000, 1511319600, 1511323200, 1511326800, 1511330400, 1511334000, 
    1511337600, 1511341200, 1511344800, 1511348400, 1511352000, 1511355600, 
    1511359200, 1511362800, 1511366400, 1511370000, 1511373600, 1511377200, 
    1511380800, 1511384400, 1511388000, 1511391600, 1511395200, 1511398800, 
    1511402400, 1511406000, 1511409600, 1511413200, 1511416800, 1511420400, 
    1511424000, 1511427600, 1511431200, 1511434800, 1511438400, 1511442000, 
    1511445600, 1511449200, 1511452800, 1511456400, 1511460000, 1511463600, 
    1511467200, 1511470800, 1511474400, 1511478000, 1511481600, 1511485200, 
    1511488800, 1511492400, 1511496000, 1511499600, 1511503200, 1511506800, 
    1511510400, 1511514000, 1511517600, 1511521200, 1511524800, 1511528400, 
    1511532000, 1511535600, 1511539200, 1511542800, 1511546400, 1511550000, 
    1511553600, 1511557200, 1511560800, 1511564400, 1511568000, 1511571600, 
    1511575200, 1511578800, 1511582400, 1511586000, 1511589600, 1511593200, 
    1511596800, 1511600400, 1511604000, 1511607600, 1511611200, 1511614800, 
    1511618400, 1511622000, 1511625600, 1511629200, 1511632800, 1511636400, 
    1511640000, 1511643600, 1511647200, 1511650800, 1511654400, 1511658000, 
    1511661600, 1511665200, 1511668800, 1511672400, 1511676000, 1511679600, 
    1511683200, 1511686800, 1511690400, 1511694000, 1511697600, 1511701200, 
    1511704800, 1511708400, 1511712000, 1511715600, 1511719200, 1511722800, 
    1511726400, 1511730000, 1511733600, 1511737200, 1511740800, 1511744400, 
    1511748000, 1511751600, 1511755200, 1511758800, 1511762400, 1511766000, 
    1511769600, 1511773200, 1511776800, 1511780400, 1511784000, 1511787600, 
    1511791200, 1511794800, 1511798400, 1511802000, 1511805600, 1511809200, 
    1511812800, 1511816400, 1511820000, 1511823600, 1511827200, 1511830800, 
    1511834400, 1511838000, 1511841600, 1511845200, 1511848800, 1511852400, 
    1511856000, 1511859600, 1511863200, 1511866800, 1511870400, 1511874000, 
    1511877600, 1511881200, 1511884800, 1511888400, 1511892000, 1511895600, 
    1511899200, 1511902800, 1511906400, 1511910000, 1511913600, 1511917200, 
    1511920800, 1511924400, 1511928000, 1511931600, 1511935200, 1511938800, 
    1511942400, 1511946000, 1511949600, 1511953200, 1511956800, 1511960400, 
    1511964000, 1511967600, 1511971200, 1511974800, 1511978400, 1511982000, 
    1511985600, 1511989200, 1511992800, 1511996400, 1512000000, 1512003600, 
    1512007200, 1512010800, 1512014400, 1512018000, 1512021600, 1512025200, 
    1512028800, 1512032400, 1512036000, 1512039600, 1512043200, 1512046800, 
    1512050400, 1512054000, 1512057600, 1512061200, 1512064800, 1512068400, 
    1512072000, 1512075600, 1512079200, 1512082800, 1512086400, 1512090000, 
    1512093600, 1512097200, 1512100800, 1512104400, 1512108000, 1512111600, 
    1512115200, 1512118800, 1512122400, 1512126000, 1512129600, 1512133200, 
    1512136800, 1512140400, 1512144000, 1512147600, 1512151200, 1512154800, 
    1512158400, 1512162000, 1512165600, 1512169200, 1512172800, 1512176400, 
    1512180000, 1512183600, 1512187200, 1512190800, 1512194400, 1512198000, 
    1512201600, 1512205200, 1512208800, 1512212400, 1512216000, 1512219600, 
    1512223200, 1512226800, 1512230400, 1512234000, 1512237600, 1512241200, 
    1512244800, 1512248400, 1512252000, 1512255600, 1512259200, 1512262800, 
    1512266400, 1512270000, 1512273600, 1512277200, 1512280800, 1512284400, 
    1512288000, 1512291600, 1512295200, 1512298800, 1512302400, 1512306000, 
    1512309600, 1512313200, 1512316800, 1512320400, 1512324000, 1512327600, 
    1512331200, 1512334800, 1512338400, 1512342000, 1512345600, 1512349200, 
    1512352800, 1512356400, 1512360000, 1512363600, 1512367200, 1512370800, 
    1512374400, 1512378000, 1512381600, 1512385200, 1512388800, 1512392400, 
    1512396000, 1512399600, 1512403200, 1512406800, 1512410400, 1512414000, 
    1512417600, 1512421200, 1512424800, 1512428400, 1512432000, 1512435600, 
    1512439200, 1512442800, 1512446400, 1512450000, 1512453600, 1512457200, 
    1512460800, 1512464400, 1512468000, 1512471600, 1512475200, 1512478800, 
    1512482400, 1512486000, 1512489600, 1512493200, 1512496800, 1512500400, 
    1512504000, 1512507600, 1512511200, 1512514800, 1512518400, 1512522000, 
    1512525600, 1512529200, 1512532800, 1512536400, 1512540000, 1512543600, 
    1512547200, 1512550800, 1512554400, 1512558000, 1512561600, 1512565200, 
    1512568800, 1512572400, 1512576000, 1512579600, 1512583200, 1512586800, 
    1512590400, 1512594000, 1512597600, 1512601200, 1512604800, 1512608400, 
    1512612000, 1512615600, 1512619200, 1512622800, 1512626400, 1512630000, 
    1512633600, 1512637200, 1512640800, 1512644400, 1512648000, 1512651600, 
    1512655200, 1512658800, 1512662400, 1512666000, 1512669600, 1512673200, 
    1512676800, 1512680400, 1512684000, 1512687600, 1512691200, 1512694800, 
    1512698400, 1512702000, 1512705600, 1512709200, 1512712800, 1512716400, 
    1512720000, 1512723600, 1512727200, 1512730800, 1512734400, 1512738000, 
    1512741600, 1512745200, 1512748800, 1512752400, 1512756000, 1512759600, 
    1512763200, 1512766800, 1512770400, 1512774000, 1512777600, 1512781200, 
    1512784800, 1512788400, 1512792000, 1512795600, 1512799200, 1512802800, 
    1512806400, 1512810000, 1512813600, 1512817200, 1512820800, 1512824400, 
    1512828000, 1512831600, 1512835200, 1512838800, 1512842400, 1512846000, 
    1512849600, 1512853200, 1512856800, 1512860400, 1512864000, 1512867600, 
    1512871200, 1512874800, 1512878400, 1512882000, 1512885600, 1512889200, 
    1512892800, 1512896400, 1512900000, 1512903600, 1512907200, 1512910800, 
    1512914400, 1512918000, 1512921600, 1512925200, 1512928800, 1512932400, 
    1512936000, 1512939600, 1512943200, 1512946800, 1512950400, 1512954000, 
    1512957600, 1512961200, 1512964800, 1512968400, 1512972000, 1512975600, 
    1512979200, 1512982800, 1512986400, 1512990000, 1512993600, 1512997200, 
    1513000800, 1513004400, 1513008000, 1513011600, 1513015200, 1513018800, 
    1513022400, 1513026000, 1513029600, 1513033200, 1513036800, 1513040400, 
    1513044000, 1513047600, 1513051200, 1513054800, 1513058400, 1513062000, 
    1513065600, 1513069200, 1513072800, 1513076400, 1513080000, 1513083600, 
    1513087200, 1513090800, 1513094400, 1513098000, 1513101600, 1513105200, 
    1513108800, 1513112400, 1513116000, 1513119600, 1513123200, 1513126800, 
    1513130400, 1513134000, 1513137600, 1513141200, 1513144800, 1513148400, 
    1513152000, 1513155600, 1513159200, 1513162800, 1513166400, 1513170000, 
    1513173600, 1513177200, 1513180800, 1513184400, 1513188000, 1513191600, 
    1513195200, 1513198800, 1513202400, 1513206000, 1513209600, 1513213200, 
    1513216800, 1513220400, 1513224000, 1513227600, 1513231200, 1513234800, 
    1513238400, 1513242000, 1513245600, 1513249200, 1513252800, 1513256400, 
    1513260000, 1513263600, 1513267200, 1513270800, 1513274400, 1513278000, 
    1513281600, 1513285200, 1513288800, 1513292400, 1513296000, 1513299600, 
    1513303200, 1513306800, 1513310400, 1513314000, 1513317600, 1513321200, 
    1513324800, 1513328400, 1513332000, 1513335600, 1513339200, 1513342800, 
    1513346400, 1513350000, 1513353600, 1513357200, 1513360800, 1513364400, 
    1513368000, 1513371600, 1513375200, 1513378800, 1513382400, 1513386000, 
    1513389600, 1513393200, 1513396800, 1513400400, 1513404000, 1513407600, 
    1513411200, 1513414800, 1513418400, 1513422000, 1513425600, 1513429200, 
    1513432800, 1513436400, 1513440000, 1513443600, 1513447200, 1513450800, 
    1513454400, 1513458000, 1513461600, 1513465200, 1513468800, 1513472400, 
    1513476000, 1513479600, 1513483200, 1513486800, 1513490400, 1513494000, 
    1513497600, 1513501200, 1513504800, 1513508400, 1513512000, 1513515600, 
    1513519200, 1513522800, 1513526400, 1513530000, 1513533600, 1513537200, 
    1513540800, 1513544400, 1513548000, 1513551600, 1513555200, 1513558800, 
    1513562400, 1513566000, 1513569600, 1513573200, 1513576800, 1513580400, 
    1513584000, 1513587600, 1513591200, 1513594800, 1513598400, 1513602000, 
    1513605600, 1513609200, 1513612800, 1513616400, 1513620000, 1513623600, 
    1513627200, 1513630800, 1513634400, 1513638000, 1513641600, 1513645200, 
    1513648800, 1513652400, 1513656000, 1513659600, 1513663200, 1513666800, 
    1513670400, 1513674000, 1513677600, 1513681200, 1513684800, 1513688400, 
    1513692000, 1513695600, 1513699200, 1513702800, 1513706400, 1513710000, 
    1513713600, 1513717200, 1513720800, 1513724400, 1513728000, 1513731600, 
    1513735200, 1513738800, 1513742400, 1513746000, 1513749600, 1513753200, 
    1513756800, 1513760400, 1513764000, 1513767600, 1513771200, 1513774800, 
    1513778400, 1513782000, 1513785600, 1513789200, 1513792800, 1513796400, 
    1513800000, 1513803600, 1513807200, 1513810800, 1513814400, 1513818000, 
    1513821600, 1513825200, 1513828800, 1513832400, 1513836000, 1513839600, 
    1513843200, 1513846800, 1513850400, 1513854000, 1513857600, 1513861200, 
    1513864800, 1513868400, 1513872000, 1513875600, 1513879200, 1513882800, 
    1513886400, 1513890000, 1513893600, 1513897200, 1513900800, 1513904400, 
    1513908000, 1513911600, 1513915200, 1513918800, 1513922400, 1513926000, 
    1513929600, 1513933200, 1513936800, 1513940400, 1513944000, 1513947600, 
    1513951200, 1513954800, 1513958400, 1513962000, 1513965600, 1513969200, 
    1513972800, 1513976400, 1513980000, 1513983600, 1513987200, 1513990800, 
    1513994400, 1513998000, 1514001600, 1514005200, 1514008800, 1514012400, 
    1514016000, 1514019600, 1514023200, 1514026800, 1514030400, 1514034000, 
    1514037600, 1514041200, 1514044800, 1514048400, 1514052000, 1514055600, 
    1514059200, 1514062800, 1514066400, 1514070000, 1514073600, 1514077200, 
    1514080800, 1514084400, 1514088000, 1514091600, 1514095200, 1514098800, 
    1514102400, 1514106000, 1514109600, 1514113200, 1514116800, 1514120400, 
    1514124000, 1514127600, 1514131200, 1514134800, 1514138400, 1514142000, 
    1514145600, 1514149200, 1514152800, 1514156400, 1514160000, 1514163600, 
    1514167200, 1514170800, 1514174400, 1514178000, 1514181600, 1514185200, 
    1514188800, 1514192400, 1514196000, 1514199600, 1514203200, 1514206800, 
    1514210400, 1514214000, 1514217600, 1514221200, 1514224800, 1514228400, 
    1514232000, 1514235600, 1514239200, 1514242800, 1514246400, 1514250000, 
    1514253600, 1514257200, 1514260800, 1514264400, 1514268000, 1514271600, 
    1514275200, 1514278800, 1514282400, 1514286000, 1514289600, 1514293200, 
    1514296800, 1514300400, 1514304000, 1514307600, 1514311200, 1514314800, 
    1514318400, 1514322000, 1514325600, 1514329200, 1514332800, 1514336400, 
    1514340000, 1514343600, 1514347200, 1514350800, 1514354400, 1514358000, 
    1514361600, 1514365200, 1514368800, 1514372400, 1514376000, 1514379600, 
    1514383200, 1514386800, 1514390400, 1514394000, 1514397600, 1514401200, 
    1514404800, 1514408400, 1514412000, 1514415600, 1514419200, 1514422800, 
    1514426400, 1514430000, 1514433600, 1514437200, 1514440800, 1514444400, 
    1514448000, 1514451600, 1514455200, 1514458800, 1514462400, 1514466000, 
    1514469600, 1514473200, 1514476800, 1514480400, 1514484000, 1514487600, 
    1514491200, 1514494800, 1514498400, 1514502000, 1514505600, 1514509200, 
    1514512800, 1514516400, 1514520000, 1514523600, 1514527200, 1514530800, 
    1514534400, 1514538000, 1514541600, 1514545200, 1514548800, 1514552400, 
    1514556000, 1514559600, 1514563200, 1514566800, 1514570400, 1514574000, 
    1514577600, 1514581200, 1514584800, 1514588400, 1514592000, 1514595600, 
    1514599200, 1514602800, 1514606400, 1514610000, 1514613600, 1514617200, 
    1514620800, 1514624400, 1514628000, 1514631600, 1514635200, 1514638800, 
    1514642400, 1514646000, 1514649600, 1514653200, 1514656800, 1514660400, 
    1514664000, 1514667600, 1514671200, 1514674800, 1514678400, 1514682000, 
    1514685600, 1514689200, 1514692800, 1514696400, 1514700000, 1514703600, 
    1514707200, 1514710800, 1514714400, 1514718000, 1514721600, 1514725200, 
    1514728800, 1514732400, 1514736000, 1514739600, 1514743200, 1514746800, 
    1514750400, 1514754000, 1514757600, 1514761200, 1514764800, 1514768400, 
    1514772000, 1514775600, 1514779200, 1514782800, 1514786400, 1514790000, 
    1514793600, 1514797200, 1514800800, 1514804400, 1514808000, 1514811600, 
    1514815200, 1514818800, 1514822400, 1514826000, 1514829600, 1514833200, 
    1514836800, 1514840400, 1514844000, 1514847600, 1514851200, 1514854800, 
    1514858400, 1514862000, 1514865600, 1514869200, 1514872800, 1514876400, 
    1514880000, 1514883600, 1514887200, 1514890800, 1514894400, 1514898000, 
    1514901600, 1514905200, 1514908800, 1514912400, 1514916000, 1514919600, 
    1514923200, 1514926800, 1514930400, 1514934000, 1514937600, 1514941200, 
    1514944800, 1514948400, 1514952000, 1514955600, 1514959200, 1514962800, 
    1514966400, 1514970000, 1514973600, 1514977200, 1514980800, 1514984400, 
    1514988000, 1514991600, 1514995200, 1514998800, 1515002400, 1515006000, 
    1515009600, 1515013200, 1515016800, 1515020400, 1515024000, 1515027600, 
    1515031200, 1515034800, 1515038400, 1515042000, 1515045600, 1515049200, 
    1515052800, 1515056400, 1515060000, 1515063600, 1515067200, 1515070800, 
    1515074400, 1515078000, 1515081600, 1515085200, 1515088800, 1515092400, 
    1515096000, 1515099600, 1515103200, 1515106800, 1515110400, 1515114000, 
    1515117600, 1515121200, 1515124800, 1515128400, 1515132000, 1515135600, 
    1515139200, 1515142800, 1515146400, 1515150000, 1515153600, 1515157200, 
    1515160800, 1515164400, 1515168000, 1515171600, 1515175200, 1515178800, 
    1515182400, 1515186000, 1515189600, 1515193200, 1515196800, 1515200400, 
    1515204000, 1515207600, 1515211200, 1515214800, 1515218400, 1515222000, 
    1515225600, 1515229200, 1515232800, 1515236400, 1515240000, 1515243600, 
    1515247200, 1515250800, 1515254400, 1515258000, 1515261600, 1515265200, 
    1515268800, 1515272400, 1515276000, 1515279600, 1515283200, 1515286800, 
    1515290400, 1515294000, 1515297600, 1515301200, 1515304800, 1515308400, 
    1515312000, 1515315600, 1515319200, 1515322800, 1515326400, 1515330000, 
    1515333600, 1515337200, 1515340800, 1515344400, 1515348000, 1515351600, 
    1515355200, 1515358800, 1515362400, 1515366000, 1515369600, 1515373200, 
    1515376800, 1515380400, 1515384000, 1515387600, 1515391200, 1515394800, 
    1515398400, 1515402000, 1515405600, 1515409200, 1515412800, 1515416400, 
    1515420000, 1515423600, 1515427200, 1515430800, 1515434400, 1515438000, 
    1515441600, 1515445200, 1515448800, 1515452400, 1515456000, 1515459600, 
    1515463200, 1515466800, 1515470400, 1515474000, 1515477600, 1515481200, 
    1515484800, 1515488400, 1515492000, 1515495600, 1515499200, 1515502800, 
    1515506400, 1515510000, 1515513600, 1515517200, 1515520800, 1515524400, 
    1515528000, 1515531600, 1515535200, 1515538800, 1515542400, 1515546000, 
    1515549600, 1515553200, 1515556800, 1515560400, 1515564000, 1515567600, 
    1515571200, 1515574800, 1515578400, 1515582000, 1515585600, 1515589200, 
    1515592800, 1515596400, 1515600000, 1515603600, 1515607200, 1515610800, 
    1515614400, 1515618000, 1515621600, 1515625200, 1515628800, 1515632400, 
    1515636000, 1515639600, 1515643200, 1515646800, 1515650400, 1515654000, 
    1515657600, 1515661200, 1515664800, 1515668400, 1515672000, 1515675600, 
    1515679200, 1515682800, 1515686400, 1515690000, 1515693600, 1515697200, 
    1515700800, 1515704400, 1515708000, 1515711600, 1515715200, 1515718800, 
    1515722400, 1515726000, 1515729600, 1515733200, 1515736800, 1515740400, 
    1515744000, 1515747600, 1515751200, 1515754800, 1515758400, 1515762000, 
    1515765600, 1515769200, 1515772800, 1515776400, 1515780000, 1515783600, 
    1515787200, 1515790800, 1515794400, 1515798000, 1515801600, 1515805200, 
    1515808800, 1515812400, 1515816000, 1515819600, 1515823200, 1515826800, 
    1515830400, 1515834000, 1515837600, 1515841200, 1515844800, 1515848400, 
    1515852000, 1515855600, 1515859200, 1515862800, 1515866400, 1515870000, 
    1515873600, 1515877200, 1515880800, 1515884400, 1515888000, 1515891600, 
    1515895200, 1515898800, 1515902400, 1515906000, 1515909600, 1515913200, 
    1515916800, 1515920400, 1515924000, 1515927600, 1515931200, 1515934800, 
    1515938400, 1515942000, 1515945600, 1515949200, 1515952800, 1515956400, 
    1515960000, 1515963600, 1515967200, 1515970800, 1515974400, 1515978000, 
    1515981600, 1515985200, 1515988800, 1515992400, 1515996000, 1515999600, 
    1516003200, 1516006800, 1516010400, 1516014000, 1516017600, 1516021200, 
    1516024800, 1516028400, 1516032000, 1516035600, 1516039200, 1516042800, 
    1516046400, 1516050000, 1516053600, 1516057200, 1516060800, 1516064400, 
    1516068000, 1516071600, 1516075200, 1516078800, 1516082400, 1516086000, 
    1516089600, 1516093200, 1516096800, 1516100400, 1516104000, 1516107600, 
    1516111200, 1516114800, 1516118400, 1516122000, 1516125600, 1516129200, 
    1516132800, 1516136400, 1516140000, 1516143600, 1516147200, 1516150800, 
    1516154400, 1516158000, 1516161600, 1516165200, 1516168800, 1516172400, 
    1516176000, 1516179600, 1516183200, 1516186800, 1516190400, 1516194000, 
    1516197600, 1516201200, 1516204800, 1516208400, 1516212000, 1516215600, 
    1516219200, 1516222800, 1516226400, 1516230000, 1516233600, 1516237200, 
    1516240800, 1516244400, 1516248000, 1516251600, 1516255200, 1516258800, 
    1516262400, 1516266000, 1516269600, 1516273200, 1516276800, 1516280400, 
    1516284000, 1516287600, 1516291200, 1516294800, 1516298400, 1516302000, 
    1516305600, 1516309200, 1516312800, 1516316400, 1516320000, 1516323600, 
    1516327200, 1516330800, 1516334400, 1516338000, 1516341600, 1516345200, 
    1516348800, 1516352400, 1516356000, 1516359600, 1516363200, 1516366800, 
    1516370400, 1516374000, 1516377600, 1516381200, 1516384800, 1516388400, 
    1516392000, 1516395600, 1516399200, 1516402800, 1516406400, 1516410000, 
    1516413600, 1516417200, 1516420800, 1516424400, 1516428000, 1516431600, 
    1516435200, 1516438800, 1516442400, 1516446000, 1516449600, 1516453200, 
    1516456800, 1516460400, 1516464000, 1516467600, 1516471200, 1516474800, 
    1516478400, 1516482000, 1516485600, 1516489200, 1516492800, 1516496400, 
    1516500000, 1516503600, 1516507200, 1516510800, 1516514400, 1516518000, 
    1516521600, 1516525200, 1516528800, 1516532400, 1516536000, 1516539600, 
    1516543200, 1516546800, 1516550400, 1516554000, 1516557600, 1516561200, 
    1516564800, 1516568400, 1516572000, 1516575600, 1516579200, 1516582800, 
    1516586400, 1516590000, 1516593600, 1516597200, 1516600800, 1516604400, 
    1516608000, 1516611600, 1516615200, 1516618800, 1516622400, 1516626000, 
    1516629600, 1516633200, 1516636800, 1516640400, 1516644000, 1516647600, 
    1516651200, 1516654800, 1516658400, 1516662000, 1516665600, 1516669200, 
    1516672800, 1516676400, 1516680000, 1516683600, 1516687200, 1516690800, 
    1516694400, 1516698000, 1516701600, 1516705200, 1516708800, 1516712400, 
    1516716000, 1516719600, 1516723200, 1516726800, 1516730400, 1516734000, 
    1516737600, 1516741200, 1516744800, 1516748400, 1516752000, 1516755600, 
    1516759200, 1516762800, 1516766400, 1516770000, 1516773600, 1516777200, 
    1516780800, 1516784400, 1516788000, 1516791600, 1516795200, 1516798800, 
    1516802400, 1516806000, 1516809600, 1516813200, 1516816800, 1516820400, 
    1516824000, 1516827600, 1516831200, 1516834800, 1516838400, 1516842000, 
    1516845600, 1516849200, 1516852800, 1516856400, 1516860000, 1516863600, 
    1516867200, 1516870800, 1516874400, 1516878000, 1516881600, 1516885200, 
    1516888800, 1516892400, 1516896000, 1516899600, 1516903200, 1516906800, 
    1516910400, 1516914000, 1516917600, 1516921200, 1516924800, 1516928400, 
    1516932000, 1516935600, 1516939200, 1516942800, 1516946400, 1516950000, 
    1516953600, 1516957200, 1516960800, 1516964400, 1516968000, 1516971600, 
    1516975200, 1516978800, 1516982400, 1516986000, 1516989600, 1516993200, 
    1516996800, 1517000400, 1517004000, 1517007600, 1517011200, 1517014800, 
    1517018400, 1517022000, 1517025600, 1517029200, 1517032800, 1517036400, 
    1517040000, 1517043600, 1517047200, 1517050800, 1517054400, 1517058000, 
    1517061600, 1517065200, 1517068800, 1517072400, 1517076000, 1517079600, 
    1517083200, 1517086800, 1517090400, 1517094000, 1517097600, 1517101200, 
    1517104800, 1517108400, 1517112000, 1517115600, 1517119200, 1517122800, 
    1517126400, 1517130000, 1517133600, 1517137200, 1517140800, 1517144400, 
    1517148000, 1517151600, 1517155200, 1517158800, 1517162400, 1517166000, 
    1517169600, 1517173200, 1517176800, 1517180400, 1517184000, 1517187600, 
    1517191200, 1517194800, 1517198400, 1517202000, 1517205600, 1517209200, 
    1517212800, 1517216400, 1517220000, 1517223600, 1517227200, 1517230800, 
    1517234400, 1517238000, 1517241600, 1517245200, 1517248800, 1517252400, 
    1517256000, 1517259600, 1517263200, 1517266800, 1517270400, 1517274000, 
    1517277600, 1517281200, 1517284800, 1517288400, 1517292000, 1517295600, 
    1517299200, 1517302800, 1517306400, 1517310000, 1517313600, 1517317200, 
    1517320800, 1517324400, 1517328000, 1517331600, 1517335200, 1517338800, 
    1517342400, 1517346000, 1517349600, 1517353200, 1517356800, 1517360400, 
    1517364000, 1517367600, 1517371200, 1517374800, 1517378400, 1517382000, 
    1517385600, 1517389200, 1517392800, 1517396400, 1517400000, 1517403600, 
    1517407200, 1517410800, 1517414400, 1517418000, 1517421600, 1517425200, 
    1517428800, 1517432400, 1517436000, 1517439600, 1517443200, 1517446800, 
    1517450400, 1517454000, 1517457600, 1517461200, 1517464800, 1517468400, 
    1517472000, 1517475600, 1517479200, 1517482800, 1517486400, 1517490000, 
    1517493600, 1517497200, 1517500800, 1517504400, 1517508000, 1517511600, 
    1517515200, 1517518800, 1517522400, 1517526000, 1517529600, 1517533200, 
    1517536800, 1517540400, 1517544000, 1517547600, 1517551200, 1517554800, 
    1517558400, 1517562000, 1517565600, 1517569200, 1517572800, 1517576400, 
    1517580000, 1517583600, 1517587200, 1517590800, 1517594400, 1517598000, 
    1517601600, 1517605200, 1517608800, 1517612400, 1517616000, 1517619600, 
    1517623200, 1517626800, 1517630400, 1517634000, 1517637600, 1517641200, 
    1517644800, 1517648400, 1517652000, 1517655600, 1517659200, 1517662800, 
    1517666400, 1517670000, 1517673600, 1517677200, 1517680800, 1517684400, 
    1517688000, 1517691600, 1517695200, 1517698800, 1517702400, 1517706000, 
    1517709600, 1517713200, 1517716800, 1517720400, 1517724000, 1517727600, 
    1517731200, 1517734800, 1517738400, 1517742000, 1517745600, 1517749200, 
    1517752800, 1517756400, 1517760000, 1517763600, 1517767200, 1517770800, 
    1517774400, 1517778000, 1517781600, 1517785200, 1517788800, 1517792400, 
    1517796000, 1517799600, 1517803200, 1517806800, 1517810400, 1517814000, 
    1517817600, 1517821200, 1517824800, 1517828400, 1517832000, 1517835600, 
    1517839200, 1517842800, 1517846400, 1517850000, 1517853600, 1517857200, 
    1517860800, 1517864400, 1517868000, 1517871600, 1517875200, 1517878800, 
    1517882400, 1517886000, 1517889600, 1517893200, 1517896800, 1517900400, 
    1517904000, 1517907600, 1517911200, 1517914800, 1517918400, 1517922000, 
    1517925600, 1517929200, 1517932800, 1517936400, 1517940000, 1517943600, 
    1517947200, 1517950800, 1517954400, 1517958000, 1517961600, 1517965200, 
    1517968800, 1517972400, 1517976000, 1517979600, 1517983200, 1517986800, 
    1517990400, 1517994000, 1517997600, 1518001200, 1518004800, 1518008400, 
    1518012000, 1518015600, 1518019200, 1518022800, 1518026400, 1518030000, 
    1518033600, 1518037200, 1518040800, 1518044400, 1518048000, 1518051600, 
    1518055200, 1518058800, 1518062400, 1518066000, 1518069600, 1518073200, 
    1518076800, 1518080400, 1518084000, 1518087600, 1518091200, 1518094800, 
    1518098400, 1518102000, 1518105600, 1518109200, 1518112800, 1518116400, 
    1518120000, 1518123600, 1518127200, 1518130800, 1518134400, 1518138000, 
    1518141600, 1518145200, 1518148800, 1518152400, 1518156000, 1518159600, 
    1518163200, 1518166800, 1518170400, 1518174000, 1518177600, 1518181200, 
    1518184800, 1518188400, 1518192000, 1518195600, 1518199200, 1518202800, 
    1518206400, 1518210000, 1518213600, 1518217200, 1518220800, 1518224400, 
    1518228000, 1518231600, 1518235200, 1518238800, 1518242400, 1518246000, 
    1518249600, 1518253200, 1518256800, 1518260400, 1518264000, 1518267600, 
    1518271200, 1518274800, 1518278400, 1518282000, 1518285600, 1518289200, 
    1518292800, 1518296400, 1518300000, 1518303600, 1518307200, 1518310800, 
    1518314400, 1518318000, 1518321600, 1518325200, 1518328800, 1518332400, 
    1518336000, 1518339600, 1518343200, 1518346800, 1518350400, 1518354000, 
    1518357600, 1518361200, 1518364800, 1518368400, 1518372000, 1518375600, 
    1518379200, 1518382800, 1518386400, 1518390000, 1518393600, 1518397200, 
    1518400800, 1518404400, 1518408000, 1518411600, 1518415200, 1518418800, 
    1518422400, 1518426000, 1518429600, 1518433200, 1518436800, 1518440400, 
    1518444000, 1518447600, 1518451200, 1518454800, 1518458400, 1518462000, 
    1518465600, 1518469200, 1518472800, 1518476400, 1518480000, 1518483600, 
    1518487200, 1518490800, 1518494400, 1518498000, 1518501600, 1518505200, 
    1518508800, 1518512400, 1518516000, 1518519600, 1518523200, 1518526800, 
    1518530400, 1518534000, 1518537600, 1518541200, 1518544800, 1518548400, 
    1518552000, 1518555600, 1518559200, 1518562800, 1518566400, 1518570000, 
    1518573600, 1518577200, 1518580800, 1518584400, 1518588000, 1518591600, 
    1518595200, 1518598800, 1518602400, 1518606000, 1518609600, 1518613200, 
    1518616800, 1518620400, 1518624000, 1518627600, 1518631200, 1518634800, 
    1518638400, 1518642000, 1518645600, 1518649200, 1518652800, 1518656400, 
    1518660000, 1518663600, 1518667200, 1518670800, 1518674400, 1518678000, 
    1518681600, 1518685200, 1518688800, 1518692400, 1518696000, 1518699600, 
    1518703200, 1518706800, 1518710400, 1518714000, 1518717600, 1518721200, 
    1518724800, 1518728400, 1518732000, 1518735600, 1518739200, 1518742800, 
    1518746400, 1518750000, 1518753600, 1518757200, 1518760800, 1518764400, 
    1518768000, 1518771600, 1518775200, 1518778800, 1518782400, 1518786000, 
    1518789600, 1518793200, 1518796800, 1518800400, 1518804000, 1518807600, 
    1518811200, 1518814800, 1518818400, 1518822000, 1518825600, 1518829200, 
    1518832800, 1518836400, 1518840000, 1518843600, 1518847200, 1518850800, 
    1518854400, 1518858000, 1518861600, 1518865200, 1518868800, 1518872400, 
    1518876000, 1518879600, 1518883200, 1518886800, 1518890400, 1518894000, 
    1518897600, 1518901200, 1518904800, 1518908400, 1518912000, 1518915600, 
    1518919200, 1518922800, 1518926400, 1518930000, 1518933600, 1518937200, 
    1518940800, 1518944400, 1518948000, 1518951600, 1518955200, 1518958800, 
    1518962400, 1518966000, 1518969600, 1518973200, 1518976800, 1518980400, 
    1518984000, 1518987600, 1518991200, 1518994800, 1518998400, 1519002000, 
    1519005600, 1519009200, 1519012800, 1519016400, 1519020000, 1519023600, 
    1519027200, 1519030800, 1519034400, 1519038000, 1519041600, 1519045200, 
    1519048800, 1519052400, 1519056000, 1519059600, 1519063200, 1519066800, 
    1519070400, 1519074000, 1519077600, 1519081200, 1519084800, 1519088400, 
    1519092000, 1519095600, 1519099200, 1519102800, 1519106400, 1519110000, 
    1519113600, 1519117200, 1519120800, 1519124400, 1519128000, 1519131600, 
    1519135200, 1519138800, 1519142400, 1519146000, 1519149600, 1519153200, 
    1519156800, 1519160400, 1519164000, 1519167600, 1519171200, 1519174800, 
    1519178400, 1519182000, 1519185600, 1519189200, 1519192800, 1519196400, 
    1519200000, 1519203600, 1519207200, 1519210800, 1519214400, 1519218000, 
    1519221600, 1519225200, 1519228800, 1519232400, 1519236000, 1519239600, 
    1519243200, 1519246800, 1519250400, 1519254000, 1519257600, 1519261200, 
    1519264800, 1519268400, 1519272000, 1519275600, 1519279200, 1519282800, 
    1519286400, 1519290000, 1519293600, 1519297200, 1519300800, 1519304400, 
    1519308000, 1519311600, 1519315200, 1519318800, 1519322400, 1519326000, 
    1519329600, 1519333200, 1519336800, 1519340400, 1519344000, 1519347600, 
    1519351200, 1519354800, 1519358400, 1519362000, 1519365600, 1519369200, 
    1519372800, 1519376400, 1519380000, 1519383600, 1519387200, 1519390800, 
    1519394400, 1519398000, 1519401600, 1519405200, 1519408800, 1519412400, 
    1519416000, 1519419600, 1519423200, 1519426800, 1519430400, 1519434000, 
    1519437600, 1519441200, 1519444800, 1519448400, 1519452000, 1519455600, 
    1519459200, 1519462800, 1519466400, 1519470000, 1519473600, 1519477200, 
    1519480800, 1519484400, 1519488000, 1519491600, 1519495200, 1519498800, 
    1519502400, 1519506000, 1519509600, 1519513200, 1519516800, 1519520400, 
    1519524000, 1519527600, 1519531200, 1519534800, 1519538400, 1519542000, 
    1519545600, 1519549200, 1519552800, 1519556400, 1519560000, 1519563600, 
    1519567200, 1519570800, 1519574400, 1519578000, 1519581600, 1519585200, 
    1519588800, 1519592400, 1519596000, 1519599600, 1519603200, 1519606800, 
    1519610400, 1519614000, 1519617600, 1519621200, 1519624800, 1519628400, 
    1519632000, 1519635600, 1519639200, 1519642800, 1519646400, 1519650000, 
    1519653600, 1519657200, 1519660800, 1519664400, 1519668000, 1519671600, 
    1519675200, 1519678800, 1519682400, 1519686000, 1519689600, 1519693200, 
    1519696800, 1519700400, 1519704000, 1519707600, 1519711200, 1519714800, 
    1519718400, 1519722000, 1519725600, 1519729200, 1519732800, 1519736400, 
    1519740000, 1519743600, 1519747200, 1519750800, 1519754400, 1519758000, 
    1519761600, 1519765200, 1519768800, 1519772400, 1519776000, 1519779600, 
    1519783200, 1519786800, 1519790400, 1519794000, 1519797600, 1519801200, 
    1519804800, 1519808400, 1519812000, 1519815600, 1519819200, 1519822800, 
    1519826400, 1519830000, 1519833600, 1519837200, 1519840800, 1519844400, 
    1519848000, 1519851600, 1519855200, 1519858800, 1519862400, 1519866000, 
    1519869600, 1519873200, 1519876800, 1519880400, 1519884000, 1519887600, 
    1519891200, 1519894800, 1519898400, 1519902000, 1519905600, 1519909200, 
    1519912800, 1519916400, 1519920000, 1519923600, 1519927200, 1519930800, 
    1519934400, 1519938000, 1519941600, 1519945200, 1519948800, 1519952400, 
    1519956000, 1519959600, 1519963200, 1519966800, 1519970400, 1519974000, 
    1519977600, 1519981200, 1519984800, 1519988400, 1519992000, 1519995600, 
    1519999200, 1520002800, 1520006400, 1520010000, 1520013600, 1520017200, 
    1520020800, 1520024400, 1520028000, 1520031600, 1520035200, 1520038800, 
    1520042400, 1520046000, 1520049600, 1520053200, 1520056800, 1520060400, 
    1520064000, 1520067600, 1520071200, 1520074800, 1520078400, 1520082000, 
    1520085600, 1520089200, 1520092800, 1520096400, 1520100000, 1520103600, 
    1520107200, 1520110800, 1520114400, 1520118000, 1520121600, 1520125200, 
    1520128800, 1520132400, 1520136000, 1520139600, 1520143200, 1520146800, 
    1520150400, 1520154000, 1520157600, 1520161200, 1520164800, 1520168400, 
    1520172000, 1520175600, 1520179200, 1520182800, 1520186400, 1520190000, 
    1520193600, 1520197200, 1520200800, 1520204400, 1520208000, 1520211600, 
    1520215200, 1520218800, 1520222400, 1520226000, 1520229600, 1520233200, 
    1520236800, 1520240400, 1520244000, 1520247600, 1520251200, 1520254800, 
    1520258400, 1520262000, 1520265600, 1520269200, 1520272800, 1520276400, 
    1520280000, 1520283600, 1520287200, 1520290800, 1520294400, 1520298000, 
    1520301600, 1520305200, 1520308800, 1520312400, 1520316000, 1520319600, 
    1520323200, 1520326800, 1520330400, 1520334000, 1520337600, 1520341200, 
    1520344800, 1520348400, 1520352000, 1520355600, 1520359200, 1520362800, 
    1520366400, 1520370000, 1520373600, 1520377200, 1520380800, 1520384400, 
    1520388000, 1520391600, 1520395200, 1520398800, 1520402400, 1520406000, 
    1520409600, 1520413200, 1520416800, 1520420400, 1520424000, 1520427600, 
    1520431200, 1520434800, 1520438400, 1520442000, 1520445600, 1520449200, 
    1520452800, 1520456400, 1520460000, 1520463600, 1520467200, 1520470800, 
    1520474400, 1520478000, 1520481600, 1520485200, 1520488800, 1520492400, 
    1520496000, 1520499600, 1520503200, 1520506800, 1520510400, 1520514000, 
    1520517600, 1520521200, 1520524800, 1520528400, 1520532000, 1520535600, 
    1520539200, 1520542800, 1520546400, 1520550000, 1520553600, 1520557200, 
    1520560800, 1520564400, 1520568000, 1520571600, 1520575200, 1520578800, 
    1520582400, 1520586000, 1520589600, 1520593200, 1520596800, 1520600400, 
    1520604000, 1520607600, 1520611200, 1520614800, 1520618400, 1520622000, 
    1520625600, 1520629200, 1520632800, 1520636400, 1520640000, 1520643600, 
    1520647200, 1520650800, 1520654400, 1520658000, 1520661600, 1520665200, 
    1520668800, 1520672400, 1520676000, 1520679600, 1520683200, 1520686800, 
    1520690400, 1520694000, 1520697600, 1520701200, 1520704800, 1520708400, 
    1520712000, 1520715600, 1520719200, 1520722800, 1520726400, 1520730000, 
    1520733600, 1520737200, 1520740800, 1520744400, 1520748000, 1520751600, 
    1520755200, 1520758800, 1520762400, 1520766000, 1520769600, 1520773200, 
    1520776800, 1520780400, 1520784000, 1520787600, 1520791200, 1520794800, 
    1520798400, 1520802000, 1520805600, 1520809200, 1520812800, 1520816400, 
    1520820000, 1520823600, 1520827200, 1520830800, 1520834400, 1520838000, 
    1520841600, 1520845200, 1520848800, 1520852400, 1520856000, 1520859600, 
    1520863200, 1520866800, 1520870400, 1520874000, 1520877600, 1520881200, 
    1520884800, 1520888400, 1520892000, 1520895600, 1520899200, 1520902800, 
    1520906400, 1520910000, 1520913600, 1520917200, 1520920800, 1520924400, 
    1520928000, 1520931600, 1520935200, 1520938800, 1520942400, 1520946000, 
    1520949600, 1520953200, 1520956800, 1520960400, 1520964000, 1520967600, 
    1520971200, 1520974800, 1520978400, 1520982000, 1520985600, 1520989200, 
    1520992800, 1520996400, 1521000000, 1521003600, 1521007200, 1521010800, 
    1521014400, 1521018000, 1521021600, 1521025200, 1521028800, 1521032400, 
    1521036000, 1521039600, 1521043200, 1521046800, 1521050400, 1521054000, 
    1521057600, 1521061200, 1521064800, 1521068400, 1521072000, 1521075600, 
    1521079200, 1521082800, 1521086400, 1521090000, 1521093600, 1521097200, 
    1521100800, 1521104400, 1521108000, 1521111600, 1521115200, 1521118800, 
    1521122400, 1521126000, 1521129600, 1521133200, 1521136800, 1521140400, 
    1521144000, 1521147600, 1521151200, 1521154800, 1521158400, 1521162000, 
    1521165600, 1521169200, 1521172800, 1521176400, 1521180000, 1521183600, 
    1521187200, 1521190800, 1521194400, 1521198000, 1521201600, 1521205200, 
    1521208800, 1521212400, 1521216000, 1521219600, 1521223200, 1521226800, 
    1521230400, 1521234000, 1521237600, 1521241200, 1521244800, 1521248400, 
    1521252000, 1521255600, 1521259200, 1521262800, 1521266400, 1521270000, 
    1521273600, 1521277200, 1521280800, 1521284400, 1521288000, 1521291600, 
    1521295200, 1521298800, 1521302400, 1521306000, 1521309600, 1521313200, 
    1521316800, 1521320400, 1521324000, 1521327600, 1521331200, 1521334800, 
    1521338400, 1521342000, 1521345600, 1521349200, 1521352800, 1521356400, 
    1521360000, 1521363600, 1521367200, 1521370800, 1521374400, 1521378000, 
    1521381600, 1521385200, 1521388800, 1521392400, 1521396000, 1521399600, 
    1521403200, 1521406800, 1521410400, 1521414000, 1521417600, 1521421200, 
    1521424800, 1521428400, 1521432000, 1521435600, 1521439200, 1521442800, 
    1521446400, 1521450000, 1521453600, 1521457200, 1521460800, 1521464400, 
    1521468000, 1521471600, 1521475200, 1521478800, 1521482400, 1521486000, 
    1521489600, 1521493200, 1521496800, 1521500400, 1521504000, 1521507600, 
    1521511200, 1521514800, 1521518400, 1521522000, 1521525600, 1521529200, 
    1521532800, 1521536400, 1521540000, 1521543600, 1521547200, 1521550800, 
    1521554400, 1521558000, 1521561600, 1521565200, 1521568800, 1521572400, 
    1521576000, 1521579600, 1521583200, 1521586800, 1521590400, 1521594000, 
    1521597600, 1521601200, 1521604800, 1521608400, 1521612000, 1521615600, 
    1521619200, 1521622800, 1521626400, 1521630000, 1521633600, 1521637200, 
    1521640800, 1521644400, 1521648000, 1521651600, 1521655200, 1521658800, 
    1521662400, 1521666000, 1521669600, 1521673200, 1521676800, 1521680400, 
    1521684000, 1521687600, 1521691200, 1521694800, 1521698400, 1521702000, 
    1521705600, 1521709200, 1521712800, 1521716400, 1521720000, 1521723600, 
    1521727200, 1521730800, 1521734400, 1521738000, 1521741600, 1521745200, 
    1521748800, 1521752400, 1521756000, 1521759600, 1521763200, 1521766800, 
    1521770400, 1521774000, 1521777600, 1521781200, 1521784800, 1521788400, 
    1521792000, 1521795600, 1521799200, 1521802800, 1521806400, 1521810000, 
    1521813600, 1521817200, 1521820800, 1521824400, 1521828000, 1521831600, 
    1521835200, 1521838800, 1521842400, 1521846000, 1521849600, 1521853200, 
    1521856800, 1521860400, 1521864000, 1521867600, 1521871200, 1521874800, 
    1521878400, 1521882000, 1521885600, 1521889200, 1521892800, 1521896400, 
    1521900000, 1521903600, 1521907200, 1521910800, 1521914400, 1521918000, 
    1521921600, 1521925200, 1521928800, 1521932400, 1521936000, 1521939600, 
    1521943200, 1521946800, 1521950400, 1521954000, 1521957600, 1521961200, 
    1521964800, 1521968400, 1521972000, 1521975600, 1521979200, 1521982800, 
    1521986400, 1521990000, 1521993600, 1521997200, 1522000800, 1522004400, 
    1522008000, 1522011600, 1522015200, 1522018800, 1522022400, 1522026000, 
    1522029600, 1522033200, 1522036800, 1522040400, 1522044000, 1522047600, 
    1522051200, 1522054800, 1522058400, 1522062000, 1522065600, 1522069200, 
    1522072800, 1522076400, 1522080000, 1522083600, 1522087200, 1522090800, 
    1522094400, 1522098000, 1522101600, 1522105200, 1522108800, 1522112400, 
    1522116000, 1522119600, 1522123200, 1522126800, 1522130400, 1522134000, 
    1522137600, 1522141200, 1522144800, 1522148400, 1522152000, 1522155600, 
    1522159200, 1522162800, 1522166400, 1522170000, 1522173600, 1522177200, 
    1522180800, 1522184400, 1522188000, 1522191600, 1522195200, 1522198800, 
    1522202400, 1522206000, 1522209600, 1522213200, 1522216800, 1522220400, 
    1522224000, 1522227600, 1522231200, 1522234800, 1522238400, 1522242000, 
    1522245600, 1522249200, 1522252800, 1522256400, 1522260000, 1522263600, 
    1522267200, 1522270800, 1522274400, 1522278000, 1522281600, 1522285200, 
    1522288800, 1522292400, 1522296000, 1522299600, 1522303200, 1522306800, 
    1522310400, 1522314000, 1522317600, 1522321200, 1522324800, 1522328400, 
    1522332000, 1522335600, 1522339200, 1522342800, 1522346400, 1522350000, 
    1522353600, 1522357200, 1522360800, 1522364400, 1522368000, 1522371600, 
    1522375200, 1522378800, 1522382400, 1522386000, 1522389600, 1522393200, 
    1522396800, 1522400400, 1522404000, 1522407600, 1522411200, 1522414800, 
    1522418400, 1522422000, 1522425600, 1522429200, 1522432800, 1522436400, 
    1522440000, 1522443600, 1522447200, 1522450800, 1522454400, 1522458000, 
    1522461600, 1522465200, 1522468800, 1522472400, 1522476000, 1522479600, 
    1522483200, 1522486800, 1522490400, 1522494000, 1522497600, 1522501200, 
    1522504800, 1522508400, 1522512000, 1522515600, 1522519200, 1522522800, 
    1522526400, 1522530000, 1522533600, 1522537200, 1522540800, 1522544400, 
    1522548000, 1522551600, 1522555200, 1522558800, 1522562400, 1522566000, 
    1522569600, 1522573200, 1522576800, 1522580400, 1522584000, 1522587600, 
    1522591200, 1522594800, 1522598400, 1522602000, 1522605600, 1522609200, 
    1522612800, 1522616400, 1522620000, 1522623600, 1522627200, 1522630800, 
    1522634400, 1522638000, 1522641600, 1522645200, 1522648800, 1522652400, 
    1522656000, 1522659600, 1522663200, 1522666800, 1522670400, 1522674000, 
    1522677600, 1522681200, 1522684800, 1522688400, 1522692000, 1522695600, 
    1522699200, 1522702800, 1522706400, 1522710000, 1522713600, 1522717200, 
    1522720800, 1522724400, 1522728000, 1522731600, 1522735200, 1522738800, 
    1522742400, 1522746000, 1522749600, 1522753200, 1522756800, 1522760400, 
    1522764000, 1522767600, 1522771200, 1522774800, 1522778400, 1522782000, 
    1522785600, 1522789200, 1522792800, 1522796400, 1522800000, 1522803600, 
    1522807200, 1522810800, 1522814400, 1522818000, 1522821600, 1522825200, 
    1522828800, 1522832400, 1522836000, 1522839600, 1522843200, 1522846800, 
    1522850400, 1522854000, 1522857600, 1522861200, 1522864800, 1522868400, 
    1522872000, 1522875600, 1522879200, 1522882800, 1522886400, 1522890000, 
    1522893600, 1522897200, 1522900800, 1522904400, 1522908000, 1522911600, 
    1522915200, 1522918800, 1522922400, 1522926000, 1522929600, 1522933200, 
    1522936800, 1522940400, 1522944000, 1522947600, 1522951200, 1522954800, 
    1522958400, 1522962000, 1522965600, 1522969200, 1522972800, 1522976400, 
    1522980000, 1522983600, 1522987200, 1522990800, 1522994400, 1522998000, 
    1523001600, 1523005200, 1523008800, 1523012400, 1523016000, 1523019600, 
    1523023200, 1523026800, 1523030400, 1523034000, 1523037600, 1523041200, 
    1523044800, 1523048400, 1523052000, 1523055600, 1523059200, 1523062800, 
    1523066400, 1523070000, 1523073600, 1523077200, 1523080800, 1523084400, 
    1523088000, 1523091600, 1523095200, 1523098800, 1523102400, 1523106000, 
    1523109600, 1523113200, 1523116800, 1523120400, 1523124000, 1523127600, 
    1523131200, 1523134800, 1523138400, 1523142000, 1523145600, 1523149200, 
    1523152800, 1523156400, 1523160000, 1523163600, 1523167200, 1523170800, 
    1523174400, 1523178000, 1523181600, 1523185200, 1523188800, 1523192400, 
    1523196000, 1523199600, 1523203200, 1523206800, 1523210400, 1523214000, 
    1523217600, 1523221200, 1523224800, 1523228400, 1523232000, 1523235600, 
    1523239200, 1523242800, 1523246400, 1523250000, 1523253600, 1523257200, 
    1523260800, 1523264400, 1523268000, 1523271600, 1523275200, 1523278800, 
    1523282400, 1523286000, 1523289600, 1523293200, 1523296800, 1523300400, 
    1523304000, 1523307600, 1523311200, 1523314800, 1523318400, 1523322000, 
    1523325600, 1523329200, 1523332800, 1523336400, 1523340000, 1523343600, 
    1523347200, 1523350800, 1523354400, 1523358000, 1523361600, 1523365200, 
    1523368800, 1523372400, 1523376000, 1523379600, 1523383200, 1523386800, 
    1523390400, 1523394000, 1523397600, 1523401200, 1523404800, 1523408400, 
    1523412000, 1523415600, 1523419200, 1523422800, 1523426400, 1523430000, 
    1523433600, 1523437200, 1523440800, 1523444400, 1523448000, 1523451600, 
    1523455200, 1523458800, 1523462400, 1523466000, 1523469600, 1523473200, 
    1523476800, 1523480400, 1523484000, 1523487600, 1523491200, 1523494800, 
    1523498400, 1523502000, 1523505600, 1523509200, 1523512800, 1523516400, 
    1523520000, 1523523600, 1523527200, 1523530800, 1523534400, 1523538000, 
    1523541600, 1523545200, 1523548800, 1523552400, 1523556000, 1523559600, 
    1523563200, 1523566800, 1523570400, 1523574000, 1523577600, 1523581200, 
    1523584800, 1523588400, 1523592000, 1523595600, 1523599200, 1523602800, 
    1523606400, 1523610000, 1523613600, 1523617200, 1523620800, 1523624400, 
    1523628000, 1523631600, 1523635200, 1523638800, 1523642400, 1523646000, 
    1523649600, 1523653200, 1523656800, 1523660400, 1523664000, 1523667600, 
    1523671200, 1523674800, 1523678400, 1523682000, 1523685600, 1523689200, 
    1523692800, 1523696400, 1523700000, 1523703600, 1523707200, 1523710800, 
    1523714400, 1523718000, 1523721600, 1523725200, 1523728800, 1523732400, 
    1523736000, 1523739600, 1523743200, 1523746800, 1523750400, 1523754000, 
    1523757600, 1523761200, 1523764800, 1523768400, 1523772000, 1523775600, 
    1523779200, 1523782800, 1523786400, 1523790000, 1523793600, 1523797200, 
    1523800800, 1523804400, 1523808000, 1523811600, 1523815200, 1523818800, 
    1523822400, 1523826000, 1523829600, 1523833200, 1523836800, 1523840400, 
    1523844000, 1523847600, 1523851200, 1523854800, 1523858400, 1523862000, 
    1523865600, 1523869200, 1523872800, 1523876400, 1523880000, 1523883600, 
    1523887200, 1523890800, 1523894400, 1523898000, 1523901600, 1523905200, 
    1523908800, 1523912400, 1523916000, 1523919600, 1523923200, 1523926800, 
    1523930400, 1523934000, 1523937600, 1523941200, 1523944800, 1523948400, 
    1523952000, 1523955600, 1523959200, 1523962800, 1523966400, 1523970000, 
    1523973600, 1523977200, 1523980800, 1523984400, 1523988000, 1523991600, 
    1523995200, 1523998800, 1524002400, 1524006000, 1524009600, 1524013200, 
    1524016800, 1524020400, 1524024000, 1524027600, 1524031200, 1524034800, 
    1524038400, 1524042000, 1524045600, 1524049200, 1524052800, 1524056400, 
    1524060000, 1524063600, 1524067200, 1524070800, 1524074400, 1524078000, 
    1524081600, 1524085200, 1524088800, 1524092400, 1524096000, 1524099600, 
    1524103200, 1524106800, 1524110400, 1524114000, 1524117600, 1524121200, 
    1524124800, 1524128400, 1524132000, 1524135600, 1524139200, 1524142800, 
    1524146400, 1524150000, 1524153600, 1524157200, 1524160800, 1524164400, 
    1524168000, 1524171600, 1524175200, 1524178800, 1524182400, 1524186000, 
    1524189600, 1524193200, 1524196800, 1524200400, 1524204000, 1524207600, 
    1524211200, 1524214800, 1524218400, 1524222000, 1524225600, 1524229200, 
    1524232800, 1524236400, 1524240000, 1524243600, 1524247200, 1524250800, 
    1524254400, 1524258000, 1524261600, 1524265200, 1524268800, 1524272400, 
    1524276000, 1524279600, 1524283200, 1524286800, 1524290400, 1524294000, 
    1524297600, 1524301200, 1524304800, 1524308400, 1524312000, 1524315600, 
    1524319200, 1524322800, 1524326400, 1524330000, 1524333600, 1524337200, 
    1524340800, 1524344400, 1524348000, 1524351600, 1524355200, 1524358800, 
    1524362400, 1524366000, 1524369600, 1524373200, 1524376800, 1524380400, 
    1524384000, 1524387600, 1524391200, 1524394800, 1524398400, 1524402000, 
    1524405600, 1524409200, 1524412800, 1524416400, 1524420000, 1524423600, 
    1524427200, 1524430800, 1524434400, 1524438000, 1524441600, 1524445200, 
    1524448800, 1524452400, 1524456000, 1524459600, 1524463200, 1524466800, 
    1524470400, 1524474000, 1524477600, 1524481200, 1524484800, 1524488400, 
    1524492000, 1524495600, 1524499200, 1524502800, 1524506400, 1524510000, 
    1524513600, 1524517200, 1524520800, 1524524400, 1524528000, 1524531600, 
    1524535200, 1524538800, 1524542400, 1524546000, 1524549600, 1524553200, 
    1524556800, 1524560400, 1524564000, 1524567600, 1524571200, 1524574800, 
    1524578400, 1524582000, 1524585600, 1524589200, 1524592800, 1524596400, 
    1524600000, 1524603600, 1524607200, 1524610800, 1524614400, 1524618000, 
    1524621600, 1524625200, 1524628800, 1524632400, 1524636000, 1524639600, 
    1524643200, 1524646800, 1524650400, 1524654000, 1524657600, 1524661200, 
    1524664800, 1524668400, 1524672000, 1524675600, 1524679200, 1524682800, 
    1524686400, 1524690000, 1524693600, 1524697200, 1524700800, 1524704400, 
    1524708000, 1524711600, 1524715200, 1524718800, 1524722400, 1524726000, 
    1524729600, 1524733200, 1524736800, 1524740400, 1524744000, 1524747600, 
    1524751200, 1524754800, 1524758400, 1524762000, 1524765600, 1524769200, 
    1524772800, 1524776400, 1524780000, 1524783600, 1524787200, 1524790800, 
    1524794400, 1524798000, 1524801600, 1524805200, 1524808800, 1524812400, 
    1524816000, 1524819600, 1524823200, 1524826800, 1524830400, 1524834000, 
    1524837600, 1524841200, 1524844800, 1524848400, 1524852000, 1524855600, 
    1524859200, 1524862800, 1524866400, 1524870000, 1524873600, 1524877200, 
    1524880800, 1524884400, 1524888000, 1524891600, 1524895200, 1524898800, 
    1524902400, 1524906000, 1524909600, 1524913200, 1524916800, 1524920400, 
    1524924000, 1524927600, 1524931200, 1524934800, 1524938400, 1524942000, 
    1524945600, 1524949200, 1524952800, 1524956400, 1524960000, 1524963600, 
    1524967200, 1524970800, 1524974400, 1524978000, 1524981600, 1524985200, 
    1524988800, 1524992400, 1524996000, 1524999600, 1525003200, 1525006800, 
    1525010400, 1525014000, 1525017600, 1525021200, 1525024800, 1525028400, 
    1525032000, 1525035600, 1525039200, 1525042800, 1525046400, 1525050000, 
    1525053600, 1525057200, 1525060800, 1525064400, 1525068000, 1525071600, 
    1525075200, 1525078800, 1525082400, 1525086000, 1525089600, 1525093200, 
    1525096800, 1525100400, 1525104000, 1525107600, 1525111200, 1525114800, 
    1525118400, 1525122000, 1525125600, 1525129200, 1525132800, 1525136400, 
    1525140000, 1525143600, 1525147200, 1525150800, 1525154400, 1525158000, 
    1525161600, 1525165200, 1525168800, 1525172400, 1525176000, 1525179600, 
    1525183200, 1525186800, 1525190400, 1525194000, 1525197600, 1525201200, 
    1525204800, 1525208400, 1525212000, 1525215600, 1525219200, 1525222800, 
    1525226400, 1525230000, 1525233600, 1525237200, 1525240800, 1525244400, 
    1525248000, 1525251600, 1525255200, 1525258800, 1525262400, 1525266000, 
    1525269600, 1525273200, 1525276800, 1525280400, 1525284000, 1525287600, 
    1525291200, 1525294800, 1525298400, 1525302000, 1525305600, 1525309200, 
    1525312800, 1525316400, 1525320000, 1525323600, 1525327200, 1525330800, 
    1525334400, 1525338000, 1525341600, 1525345200, 1525348800, 1525352400, 
    1525356000, 1525359600, 1525363200, 1525366800, 1525370400, 1525374000, 
    1525377600, 1525381200, 1525384800, 1525388400, 1525392000, 1525395600, 
    1525399200, 1525402800, 1525406400, 1525410000, 1525413600, 1525417200, 
    1525420800, 1525424400, 1525428000, 1525431600, 1525435200, 1525438800, 
    1525442400, 1525446000, 1525449600, 1525453200, 1525456800, 1525460400, 
    1525464000, 1525467600, 1525471200, 1525474800, 1525478400, 1525482000, 
    1525485600, 1525489200, 1525492800, 1525496400, 1525500000, 1525503600, 
    1525507200, 1525510800, 1525514400, 1525518000, 1525521600, 1525525200, 
    1525528800, 1525532400, 1525536000, 1525539600, 1525543200, 1525546800, 
    1525550400, 1525554000, 1525557600, 1525561200, 1525564800, 1525568400, 
    1525572000, 1525575600, 1525579200, 1525582800, 1525586400, 1525590000, 
    1525593600, 1525597200, 1525600800, 1525604400, 1525608000, 1525611600, 
    1525615200, 1525618800, 1525622400, 1525626000, 1525629600, 1525633200, 
    1525636800, 1525640400, 1525644000, 1525647600, 1525651200, 1525654800, 
    1525658400, 1525662000, 1525665600, 1525669200, 1525672800, 1525676400, 
    1525680000, 1525683600, 1525687200, 1525690800, 1525694400, 1525698000, 
    1525701600, 1525705200, 1525708800, 1525712400, 1525716000, 1525719600, 
    1525723200, 1525726800, 1525730400, 1525734000, 1525737600, 1525741200, 
    1525744800, 1525748400, 1525752000, 1525755600, 1525759200, 1525762800, 
    1525766400, 1525770000, 1525773600, 1525777200, 1525780800, 1525784400, 
    1525788000, 1525791600, 1525795200, 1525798800, 1525802400, 1525806000, 
    1525809600, 1525813200, 1525816800, 1525820400, 1525824000, 1525827600, 
    1525831200, 1525834800, 1525838400, 1525842000, 1525845600, 1525849200, 
    1525852800, 1525856400, 1525860000, 1525863600, 1525867200, 1525870800, 
    1525874400, 1525878000, 1525881600, 1525885200, 1525888800, 1525892400, 
    1525896000, 1525899600, 1525903200, 1525906800, 1525910400, 1525914000, 
    1525917600, 1525921200, 1525924800, 1525928400, 1525932000, 1525935600, 
    1525939200, 1525942800, 1525946400, 1525950000, 1525953600, 1525957200, 
    1525960800, 1525964400, 1525968000, 1525971600, 1525975200, 1525978800, 
    1525982400, 1525986000, 1525989600, 1525993200, 1525996800, 1526000400, 
    1526004000, 1526007600, 1526011200, 1526014800, 1526018400, 1526022000, 
    1526025600, 1526029200, 1526032800, 1526036400, 1526040000, 1526043600, 
    1526047200, 1526050800, 1526054400, 1526058000, 1526061600, 1526065200, 
    1526068800, 1526072400, 1526076000, 1526079600, 1526083200, 1526086800, 
    1526090400, 1526094000, 1526097600, 1526101200, 1526104800, 1526108400, 
    1526112000, 1526115600, 1526119200, 1526122800, 1526126400, 1526130000, 
    1526133600, 1526137200, 1526140800, 1526144400, 1526148000, 1526151600, 
    1526155200, 1526158800, 1526162400, 1526166000, 1526169600, 1526173200, 
    1526176800, 1526180400, 1526184000, 1526187600, 1526191200, 1526194800, 
    1526198400, 1526202000, 1526205600, 1526209200, 1526212800, 1526216400, 
    1526220000, 1526223600, 1526227200, 1526230800, 1526234400, 1526238000, 
    1526241600, 1526245200, 1526248800, 1526252400, 1526256000, 1526259600, 
    1526263200, 1526266800, 1526270400, 1526274000, 1526277600, 1526281200, 
    1526284800, 1526288400, 1526292000, 1526295600, 1526299200, 1526302800, 
    1526306400, 1526310000, 1526313600, 1526317200, 1526320800, 1526324400, 
    1526328000, 1526331600, 1526335200, 1526338800, 1526342400, 1526346000, 
    1526349600, 1526353200, 1526356800, 1526360400, 1526364000, 1526367600, 
    1526371200, 1526374800, 1526378400, 1526382000, 1526385600, 1526389200, 
    1526392800, 1526396400, 1526400000, 1526403600, 1526407200, 1526410800, 
    1526414400, 1526418000, 1526421600, 1526425200, 1526428800, 1526432400, 
    1526436000, 1526439600, 1526443200, 1526446800, 1526450400, 1526454000, 
    1526457600, 1526461200, 1526464800, 1526468400, 1526472000, 1526475600, 
    1526479200, 1526482800, 1526486400, 1526490000, 1526493600, 1526497200, 
    1526500800, 1526504400, 1526508000, 1526511600, 1526515200, 1526518800, 
    1526522400, 1526526000, 1526529600, 1526533200, 1526536800, 1526540400, 
    1526544000, 1526547600, 1526551200, 1526554800, 1526558400, 1526562000, 
    1526565600, 1526569200, 1526572800, 1526576400, 1526580000, 1526583600, 
    1526587200, 1526590800, 1526594400, 1526598000, 1526601600, 1526605200, 
    1526608800, 1526612400, 1526616000, 1526619600, 1526623200, 1526626800, 
    1526630400, 1526634000, 1526637600, 1526641200, 1526644800, 1526648400, 
    1526652000, 1526655600, 1526659200, 1526662800, 1526666400, 1526670000, 
    1526673600, 1526677200, 1526680800, 1526684400, 1526688000, 1526691600, 
    1526695200, 1526698800, 1526702400, 1526706000, 1526709600, 1526713200, 
    1526716800, 1526720400, 1526724000, 1526727600, 1526731200, 1526734800, 
    1526738400, 1526742000, 1526745600, 1526749200, 1526752800, 1526756400, 
    1526760000, 1526763600, 1526767200, 1526770800, 1526774400, 1526778000, 
    1526781600, 1526785200, 1526788800, 1526792400, 1526796000, 1526799600, 
    1526803200, 1526806800, 1526810400, 1526814000, 1526817600, 1526821200, 
    1526824800, 1526828400, 1526832000, 1526835600, 1526839200, 1526842800, 
    1526846400, 1526850000, 1526853600, 1526857200, 1526860800, 1526864400, 
    1526868000, 1526871600, 1526875200, 1526878800, 1526882400, 1526886000, 
    1526889600, 1526893200, 1526896800, 1526900400, 1526904000, 1526907600, 
    1526911200, 1526914800, 1526918400, 1526922000, 1526925600, 1526929200, 
    1526932800, 1526936400, 1526940000, 1526943600, 1526947200, 1526950800, 
    1526954400, 1526958000, 1526961600, 1526965200, 1526968800, 1526972400, 
    1526976000, 1526979600, 1526983200, 1526986800, 1526990400, 1526994000, 
    1526997600, 1527001200, 1527004800, 1527008400, 1527012000, 1527015600, 
    1527019200, 1527022800, 1527026400, 1527030000, 1527033600, 1527037200, 
    1527040800, 1527044400, 1527048000, 1527051600, 1527055200, 1527058800, 
    1527062400, 1527066000, 1527069600, 1527073200, 1527076800, 1527080400, 
    1527084000, 1527087600, 1527091200, 1527094800, 1527098400, 1527102000, 
    1527105600, 1527109200, 1527112800, 1527116400, 1527120000, 1527123600, 
    1527127200, 1527130800, 1527134400, 1527138000, 1527141600, 1527145200, 
    1527148800, 1527152400, 1527156000, 1527159600, 1527163200, 1527166800, 
    1527170400, 1527174000, 1527177600, 1527181200, 1527184800, 1527188400, 
    1527192000, 1527195600, 1527199200, 1527202800, 1527206400, 1527210000, 
    1527213600, 1527217200, 1527220800, 1527224400, 1527228000, 1527231600, 
    1527235200, 1527238800, 1527242400, 1527246000, 1527249600, 1527253200, 
    1527256800, 1527260400, 1527264000, 1527267600, 1527271200, 1527274800, 
    1527278400, 1527282000, 1527285600, 1527289200, 1527292800, 1527296400, 
    1527300000, 1527303600, 1527307200, 1527310800, 1527314400, 1527318000, 
    1527321600, 1527325200, 1527328800, 1527332400, 1527336000, 1527339600, 
    1527343200, 1527346800, 1527350400, 1527354000, 1527357600, 1527361200, 
    1527364800, 1527368400, 1527372000, 1527375600, 1527379200, 1527382800, 
    1527386400, 1527390000, 1527393600, 1527397200, 1527400800, 1527404400, 
    1527408000, 1527411600, 1527415200, 1527418800, 1527422400, 1527426000, 
    1527429600, 1527433200, 1527436800, 1527440400, 1527444000, 1527447600, 
    1527451200, 1527454800, 1527458400, 1527462000, 1527465600, 1527469200, 
    1527472800, 1527476400, 1527480000, 1527483600, 1527487200, 1527490800, 
    1527494400, 1527498000, 1527501600, 1527505200, 1527508800, 1527512400, 
    1527516000, 1527519600, 1527523200, 1527526800, 1527530400, 1527534000, 
    1527537600, 1527541200, 1527544800, 1527548400, 1527552000, 1527555600, 
    1527559200, 1527562800, 1527566400, 1527570000, 1527573600, 1527577200, 
    1527580800, 1527584400, 1527588000, 1527591600, 1527595200, 1527598800, 
    1527602400, 1527606000, 1527609600, 1527613200, 1527616800, 1527620400, 
    1527624000, 1527627600, 1527631200, 1527634800, 1527638400, 1527642000, 
    1527645600, 1527649200, 1527652800, 1527656400, 1527660000, 1527663600, 
    1527667200, 1527670800, 1527674400, 1527678000, 1527681600, 1527685200, 
    1527688800, 1527692400, 1527696000, 1527699600, 1527703200, 1527706800, 
    1527710400, 1527714000, 1527717600, 1527721200, 1527724800, 1527728400, 
    1527732000, 1527735600, 1527739200, 1527742800, 1527746400, 1527750000, 
    1527753600, 1527757200, 1527760800, 1527764400, 1527768000, 1527771600, 
    1527775200, 1527778800, 1527782400, 1527786000, 1527789600, 1527793200, 
    1527796800, 1527800400, 1527804000, 1527807600, 1527811200, 1527814800, 
    1527818400, 1527822000, 1527825600, 1527829200, 1527832800, 1527836400, 
    1527840000, 1527843600, 1527847200, 1527850800, 1527854400, 1527858000, 
    1527861600, 1527865200, 1527868800, 1527872400, 1527876000, 1527879600, 
    1527883200, 1527886800, 1527890400, 1527894000, 1527897600, 1527901200, 
    1527904800, 1527908400, 1527912000, 1527915600, 1527919200, 1527922800, 
    1527926400, 1527930000, 1527933600, 1527937200, 1527940800, 1527944400, 
    1527948000, 1527951600, 1527955200, 1527958800, 1527962400, 1527966000, 
    1527969600, 1527973200, 1527976800, 1527980400, 1527984000, 1527987600, 
    1527991200, 1527994800, 1527998400, 1528002000, 1528005600, 1528009200, 
    1528012800, 1528016400, 1528020000, 1528023600, 1528027200, 1528030800, 
    1528034400, 1528038000, 1528041600, 1528045200, 1528048800, 1528052400, 
    1528056000, 1528059600, 1528063200, 1528066800, 1528070400, 1528074000, 
    1528077600, 1528081200, 1528084800, 1528088400, 1528092000, 1528095600, 
    1528099200, 1528102800, 1528106400, 1528110000, 1528113600, 1528117200, 
    1528120800, 1528124400, 1528128000, 1528131600, 1528135200, 1528138800, 
    1528142400, 1528146000, 1528149600, 1528153200, 1528156800, 1528160400, 
    1528164000, 1528167600, 1528171200, 1528174800, 1528178400, 1528182000, 
    1528185600, 1528189200, 1528192800, 1528196400, 1528200000, 1528203600, 
    1528207200, 1528210800, 1528214400, 1528218000, 1528221600, 1528225200, 
    1528228800, 1528232400, 1528236000, 1528239600, 1528243200, 1528246800, 
    1528250400, 1528254000, 1528257600, 1528261200, 1528264800, 1528268400, 
    1528272000, 1528275600, 1528279200, 1528282800, 1528286400, 1528290000, 
    1528293600, 1528297200, 1528300800, 1528304400, 1528308000, 1528311600, 
    1528315200, 1528318800, 1528322400, 1528326000, 1528329600, 1528333200, 
    1528336800, 1528340400, 1528344000, 1528347600, 1528351200, 1528354800, 
    1528358400, 1528362000, 1528365600, 1528369200, 1528372800, 1528376400, 
    1528380000, 1528383600, 1528387200, 1528390800, 1528394400, 1528398000, 
    1528401600, 1528405200, 1528408800, 1528412400, 1528416000, 1528419600, 
    1528423200, 1528426800, 1528430400, 1528434000, 1528437600, 1528441200, 
    1528444800, 1528448400, 1528452000, 1528455600, 1528459200, 1528462800, 
    1528466400, 1528470000, 1528473600, 1528477200, 1528480800, 1528484400, 
    1528488000, 1528491600, 1528495200, 1528498800, 1528502400, 1528506000, 
    1528509600, 1528513200, 1528516800, 1528520400, 1528524000, 1528527600, 
    1528531200, 1528534800, 1528538400, 1528542000, 1528545600, 1528549200, 
    1528552800, 1528556400, 1528560000, 1528563600, 1528567200, 1528570800, 
    1528574400, 1528578000, 1528581600, 1528585200, 1528588800, 1528592400, 
    1528596000, 1528599600, 1528603200, 1528606800, 1528610400, 1528614000, 
    1528617600, 1528621200, 1528624800, 1528628400, 1528632000, 1528635600, 
    1528639200, 1528642800, 1528646400, 1528650000, 1528653600, 1528657200, 
    1528660800, 1528664400, 1528668000, 1528671600, 1528675200, 1528678800, 
    1528682400, 1528686000, 1528689600, 1528693200, 1528696800, 1528700400, 
    1528704000, 1528707600, 1528711200, 1528714800, 1528718400, 1528722000, 
    1528725600, 1528729200, 1528732800, 1528736400, 1528740000, 1528743600, 
    1528747200, 1528750800, 1528754400, 1528758000, 1528761600, 1528765200, 
    1528768800, 1528772400, 1528776000, 1528779600, 1528783200, 1528786800, 
    1528790400, 1528794000, 1528797600, 1528801200, 1528804800, 1528808400, 
    1528812000, 1528815600, 1528819200, 1528822800, 1528826400, 1528830000, 
    1528833600, 1528837200, 1528840800, 1528844400, 1528848000, 1528851600, 
    1528855200, 1528858800, 1528862400, 1528866000, 1528869600, 1528873200, 
    1528876800, 1528880400, 1528884000, 1528887600, 1528891200, 1528894800, 
    1528898400, 1528902000, 1528905600, 1528909200, 1528912800, 1528916400, 
    1528920000, 1528923600, 1528927200, 1528930800, 1528934400, 1528938000, 
    1528941600, 1528945200, 1528948800, 1528952400, 1528956000, 1528959600, 
    1528963200, 1528966800, 1528970400, 1528974000, 1528977600, 1528981200, 
    1528984800, 1528988400, 1528992000, 1528995600, 1528999200, 1529002800, 
    1529006400, 1529010000, 1529013600, 1529017200, 1529020800, 1529024400, 
    1529028000, 1529031600, 1529035200, 1529038800, 1529042400, 1529046000, 
    1529049600, 1529053200, 1529056800, 1529060400, 1529064000, 1529067600, 
    1529071200, 1529074800, 1529078400, 1529082000, 1529085600, 1529089200, 
    1529092800, 1529096400, 1529100000, 1529103600, 1529107200, 1529110800, 
    1529114400, 1529118000, 1529121600, 1529125200, 1529128800, 1529132400, 
    1529136000, 1529139600, 1529143200, 1529146800, 1529150400, 1529154000, 
    1529157600, 1529161200, 1529164800, 1529168400, 1529172000, 1529175600, 
    1529179200, 1529182800, 1529186400, 1529190000, 1529193600, 1529197200, 
    1529200800, 1529204400, 1529208000, 1529211600, 1529215200, 1529218800, 
    1529222400, 1529226000, 1529229600, 1529233200, 1529236800, 1529240400, 
    1529244000, 1529247600, 1529251200, 1529254800, 1529258400, 1529262000, 
    1529265600, 1529269200, 1529272800, 1529276400, 1529280000, 1529283600, 
    1529287200, 1529290800, 1529294400, 1529298000, 1529301600, 1529305200, 
    1529308800, 1529312400, 1529316000, 1529319600, 1529323200, 1529326800, 
    1529330400, 1529334000, 1529337600, 1529341200, 1529344800, 1529348400, 
    1529352000, 1529355600, 1529359200, 1529362800, 1529366400, 1529370000, 
    1529373600, 1529377200, 1529380800, 1529384400, 1529388000, 1529391600, 
    1529395200, 1529398800, 1529402400, 1529406000, 1529409600, 1529413200, 
    1529416800, 1529420400, 1529424000, 1529427600, 1529431200, 1529434800, 
    1529438400, 1529442000, 1529445600, 1529449200, 1529452800, 1529456400, 
    1529460000, 1529463600, 1529467200, 1529470800, 1529474400, 1529478000, 
    1529481600, 1529485200, 1529488800, 1529492400, 1529496000, 1529499600, 
    1529503200, 1529506800, 1529510400, 1529514000, 1529517600, 1529521200, 
    1529524800, 1529528400, 1529532000, 1529535600, 1529539200, 1529542800, 
    1529546400, 1529550000, 1529553600, 1529557200, 1529560800, 1529564400, 
    1529568000, 1529571600, 1529575200, 1529578800, 1529582400, 1529586000, 
    1529589600, 1529593200, 1529596800, 1529600400, 1529604000, 1529607600, 
    1529611200, 1529614800, 1529618400, 1529622000, 1529625600, 1529629200, 
    1529632800, 1529636400, 1529640000, 1529643600, 1529647200, 1529650800, 
    1529654400, 1529658000, 1529661600, 1529665200, 1529668800, 1529672400, 
    1529676000, 1529679600, 1529683200, 1529686800, 1529690400, 1529694000, 
    1529697600, 1529701200, 1529704800, 1529708400, 1529712000, 1529715600, 
    1529719200, 1529722800, 1529726400, 1529730000, 1529733600, 1529737200, 
    1529740800, 1529744400, 1529748000, 1529751600, 1529755200, 1529758800, 
    1529762400, 1529766000, 1529769600, 1529773200, 1529776800, 1529780400, 
    1529784000, 1529787600, 1529791200, 1529794800, 1529798400, 1529802000, 
    1529805600, 1529809200, 1529812800, 1529816400, 1529820000, 1529823600, 
    1529827200, 1529830800, 1529834400, 1529838000, 1529841600, 1529845200, 
    1529848800, 1529852400, 1529856000, 1529859600, 1529863200, 1529866800, 
    1529870400, 1529874000, 1529877600, 1529881200, 1529884800, 1529888400, 
    1529892000, 1529895600, 1529899200, 1529902800, 1529906400, 1529910000, 
    1529913600, 1529917200, 1529920800, 1529924400, 1529928000, 1529931600, 
    1529935200, 1529938800, 1529942400, 1529946000, 1529949600, 1529953200, 
    1529956800, 1529960400, 1529964000, 1529967600, 1529971200, 1529974800, 
    1529978400, 1529982000, 1529985600, 1529989200, 1529992800, 1529996400, 
    1530000000, 1530003600, 1530007200, 1530010800, 1530014400, 1530018000, 
    1530021600, 1530025200, 1530028800, 1530032400, 1530036000, 1530039600, 
    1530043200, 1530046800, 1530050400, 1530054000, 1530057600, 1530061200, 
    1530064800, 1530068400, 1530072000, 1530075600, 1530079200, 1530082800, 
    1530086400, 1530090000, 1530093600, 1530097200, 1530100800, 1530104400, 
    1530108000, 1530111600, 1530115200, 1530118800, 1530122400, 1530126000, 
    1530129600, 1530133200, 1530136800, 1530140400, 1530144000, 1530147600, 
    1530151200, 1530154800, 1530158400, 1530162000, 1530165600, 1530169200, 
    1530172800, 1530176400, 1530180000, 1530183600, 1530187200, 1530190800, 
    1530194400, 1530198000, 1530201600, 1530205200, 1530208800, 1530212400, 
    1530216000, 1530219600, 1530223200, 1530226800, 1530230400, 1530234000, 
    1530237600, 1530241200, 1530244800, 1530248400, 1530252000, 1530255600, 
    1530259200, 1530262800, 1530266400, 1530270000, 1530273600, 1530277200, 
    1530280800, 1530284400, 1530288000, 1530291600, 1530295200, 1530298800, 
    1530302400, 1530306000, 1530309600, 1530313200, 1530316800, 1530320400, 
    1530324000, 1530327600, 1530331200, 1530334800, 1530338400, 1530342000, 
    1530345600, 1530349200, 1530352800, 1530356400, 1530360000, 1530363600, 
    1530367200, 1530370800, 1530374400, 1530378000, 1530381600, 1530385200, 
    1530388800, 1530392400, 1530396000, 1530399600, 1530403200, 1530406800, 
    1530410400, 1530414000, 1530417600, 1530421200, 1530424800, 1530428400, 
    1530432000, 1530435600, 1530439200, 1530442800, 1530446400, 1530450000, 
    1530453600, 1530457200, 1530460800, 1530464400, 1530468000, 1530471600, 
    1530475200, 1530478800, 1530482400, 1530486000, 1530489600, 1530493200, 
    1530496800, 1530500400, 1530504000, 1530507600, 1530511200, 1530514800, 
    1530518400, 1530522000, 1530525600, 1530529200, 1530532800, 1530536400, 
    1530540000, 1530543600, 1530547200, 1530550800, 1530554400, 1530558000, 
    1530561600, 1530565200, 1530568800, 1530572400, 1530576000, 1530579600, 
    1530583200, 1530586800, 1530590400, 1530594000, 1530597600, 1530601200, 
    1530604800, 1530608400, 1530612000, 1530615600, 1530619200, 1530622800, 
    1530626400, 1530630000, 1530633600, 1530637200, 1530640800, 1530644400, 
    1530648000, 1530651600, 1530655200, 1530658800, 1530662400, 1530666000, 
    1530669600, 1530673200, 1530676800, 1530680400, 1530684000, 1530687600, 
    1530691200, 1530694800, 1530698400, 1530702000, 1530705600, 1530709200, 
    1530712800, 1530716400, 1530720000, 1530723600, 1530727200, 1530730800, 
    1530734400, 1530738000, 1530741600, 1530745200, 1530748800, 1530752400, 
    1530756000, 1530759600, 1530763200, 1530766800, 1530770400, 1530774000, 
    1530777600, 1530781200, 1530784800, 1530788400, 1530792000, 1530795600, 
    1530799200, 1530802800, 1530806400, 1530810000, 1530813600, 1530817200, 
    1530820800, 1530824400, 1530828000, 1530831600, 1530835200, 1530838800, 
    1530842400, 1530846000, 1530849600, 1530853200, 1530856800, 1530860400, 
    1530864000, 1530867600, 1530871200, 1530874800, 1530878400, 1530882000, 
    1530885600, 1530889200, 1530892800, 1530896400, 1530900000, 1530903600, 
    1530907200, 1530910800, 1530914400, 1530918000, 1530921600, 1530925200, 
    1530928800, 1530932400, 1530936000, 1530939600, 1530943200, 1530946800, 
    1530950400, 1530954000, 1530957600, 1530961200, 1530964800, 1530968400, 
    1530972000, 1530975600, 1530979200, 1530982800, 1530986400, 1530990000, 
    1530993600, 1530997200, 1531000800, 1531004400, 1531008000, 1531011600, 
    1531015200, 1531018800, 1531022400, 1531026000, 1531029600, 1531033200, 
    1531036800, 1531040400, 1531044000, 1531047600, 1531051200, 1531054800, 
    1531058400, 1531062000, 1531065600, 1531069200, 1531072800, 1531076400, 
    1531080000, 1531083600, 1531087200, 1531090800, 1531094400, 1531098000, 
    1531101600, 1531105200, 1531108800, 1531112400, 1531116000, 1531119600, 
    1531123200, 1531126800, 1531130400, 1531134000, 1531137600, 1531141200, 
    1531144800, 1531148400, 1531152000, 1531155600, 1531159200, 1531162800, 
    1531166400, 1531170000, 1531173600, 1531177200, 1531180800, 1531184400, 
    1531188000, 1531191600, 1531195200, 1531198800, 1531202400, 1531206000, 
    1531209600, 1531213200, 1531216800, 1531220400, 1531224000, 1531227600, 
    1531231200, 1531234800, 1531238400, 1531242000, 1531245600, 1531249200, 
    1531252800, 1531256400, 1531260000, 1531263600, 1531267200, 1531270800, 
    1531274400, 1531278000, 1531281600, 1531285200, 1531288800, 1531292400, 
    1531296000, 1531299600, 1531303200, 1531306800, 1531310400, 1531314000, 
    1531317600, 1531321200, 1531324800, 1531328400, 1531332000, 1531335600, 
    1531339200, 1531342800, 1531346400, 1531350000, 1531353600, 1531357200, 
    1531360800, 1531364400, 1531368000, 1531371600, 1531375200, 1531378800, 
    1531382400, 1531386000, 1531389600, 1531393200, 1531396800, 1531400400, 
    1531404000, 1531407600, 1531411200, 1531414800, 1531418400, 1531422000, 
    1531425600, 1531429200, 1531432800, 1531436400, 1531440000, 1531443600, 
    1531447200, 1531450800, 1531454400, 1531458000, 1531461600, 1531465200, 
    1531468800, 1531472400, 1531476000, 1531479600, 1531483200, 1531486800, 
    1531490400, 1531494000, 1531497600, 1531501200, 1531504800, 1531508400, 
    1531512000, 1531515600, 1531519200, 1531522800, 1531526400, 1531530000, 
    1531533600, 1531537200, 1531540800, 1531544400, 1531548000, 1531551600, 
    1531555200, 1531558800, 1531562400, 1531566000, 1531569600, 1531573200, 
    1531576800, 1531580400, 1531584000, 1531587600, 1531591200, 1531594800, 
    1531598400, 1531602000, 1531605600, 1531609200, 1531612800, 1531616400, 
    1531620000, 1531623600, 1531627200, 1531630800, 1531634400, 1531638000, 
    1531641600, 1531645200, 1531648800, 1531652400, 1531656000, 1531659600, 
    1531663200, 1531666800, 1531670400, 1531674000, 1531677600, 1531681200, 
    1531684800, 1531688400, 1531692000, 1531695600, 1531699200, 1531702800, 
    1531706400, 1531710000, 1531713600, 1531717200, 1531720800, 1531724400, 
    1531728000, 1531731600, 1531735200, 1531738800, 1531742400, 1531746000, 
    1531749600, 1531753200, 1531756800, 1531760400, 1531764000, 1531767600, 
    1531771200, 1531774800, 1531778400, 1531782000, 1531785600, 1531789200, 
    1531792800, 1531796400, 1531800000, 1531803600, 1531807200, 1531810800, 
    1531814400, 1531818000, 1531821600, 1531825200, 1531828800, 1531832400, 
    1531836000, 1531839600, 1531843200, 1531846800, 1531850400, 1531854000, 
    1531857600, 1531861200, 1531864800, 1531868400, 1531872000, 1531875600, 
    1531879200, 1531882800, 1531886400, 1531890000, 1531893600, 1531897200, 
    1531900800, 1531904400, 1531908000, 1531911600, 1531915200, 1531918800, 
    1531922400, 1531926000, 1531929600, 1531933200, 1531936800, 1531940400, 
    1531944000, 1531947600, 1531951200, 1531954800, 1531958400, 1531962000, 
    1531965600, 1531969200, 1531972800, 1531976400, 1531980000, 1531983600, 
    1531987200, 1531990800, 1531994400, 1531998000, 1532001600, 1532005200, 
    1532008800, 1532012400, 1532016000, 1532019600, 1532023200, 1532026800, 
    1532030400, 1532034000, 1532037600, 1532041200, 1532044800, 1532048400, 
    1532052000, 1532055600, 1532059200, 1532062800, 1532066400, 1532070000, 
    1532073600, 1532077200, 1532080800, 1532084400, 1532088000, 1532091600, 
    1532095200, 1532098800, 1532102400, 1532106000, 1532109600, 1532113200, 
    1532116800, 1532120400, 1532124000, 1532127600, 1532131200, 1532134800, 
    1532138400, 1532142000, 1532145600, 1532149200, 1532152800, 1532156400, 
    1532160000, 1532163600, 1532167200, 1532170800, 1532174400, 1532178000, 
    1532181600, 1532185200, 1532188800, 1532192400, 1532196000, 1532199600, 
    1532203200, 1532206800, 1532210400, 1532214000, 1532217600, 1532221200, 
    1532224800, 1532228400, 1532232000, 1532235600, 1532239200, 1532242800, 
    1532246400, 1532250000, 1532253600, 1532257200, 1532260800, 1532264400, 
    1532268000, 1532271600, 1532275200, 1532278800, 1532282400, 1532286000, 
    1532289600, 1532293200, 1532296800, 1532300400, 1532304000, 1532307600, 
    1532311200, 1532314800, 1532318400, 1532322000, 1532325600, 1532329200, 
    1532332800, 1532336400, 1532340000, 1532343600, 1532347200, 1532350800, 
    1532354400, 1532358000, 1532361600, 1532365200, 1532368800, 1532372400, 
    1532376000, 1532379600, 1532383200, 1532386800, 1532390400, 1532394000, 
    1532397600, 1532401200, 1532404800, 1532408400, 1532412000, 1532415600, 
    1532419200, 1532422800, 1532426400, 1532430000, 1532433600, 1532437200, 
    1532440800, 1532444400, 1532448000, 1532451600, 1532455200, 1532458800, 
    1532462400, 1532466000, 1532469600, 1532473200, 1532476800, 1532480400, 
    1532484000, 1532487600, 1532491200, 1532494800, 1532498400, 1532502000, 
    1532505600, 1532509200, 1532512800, 1532516400, 1532520000, 1532523600, 
    1532527200, 1532530800, 1532534400, 1532538000, 1532541600, 1532545200, 
    1532548800, 1532552400, 1532556000, 1532559600, 1532563200, 1532566800, 
    1532570400, 1532574000, 1532577600, 1532581200, 1532584800, 1532588400, 
    1532592000, 1532595600, 1532599200, 1532602800, 1532606400, 1532610000, 
    1532613600, 1532617200, 1532620800, 1532624400, 1532628000, 1532631600, 
    1532635200, 1532638800, 1532642400, 1532646000, 1532649600, 1532653200, 
    1532656800, 1532660400, 1532664000, 1532667600, 1532671200, 1532674800, 
    1532678400, 1532682000, 1532685600, 1532689200, 1532692800, 1532696400, 
    1532700000, 1532703600, 1532707200, 1532710800, 1532714400, 1532718000, 
    1532721600, 1532725200, 1532728800, 1532732400, 1532736000, 1532739600, 
    1532743200, 1532746800, 1532750400, 1532754000, 1532757600, 1532761200, 
    1532764800, 1532768400, 1532772000, 1532775600, 1532779200, 1532782800, 
    1532786400, 1532790000, 1532793600, 1532797200, 1532800800, 1532804400, 
    1532808000, 1532811600, 1532815200, 1532818800, 1532822400, 1532826000, 
    1532829600, 1532833200, 1532836800, 1532840400, 1532844000, 1532847600, 
    1532851200, 1532854800, 1532858400, 1532862000, 1532865600, 1532869200, 
    1532872800, 1532876400, 1532880000, 1532883600, 1532887200, 1532890800, 
    1532894400, 1532898000, 1532901600, 1532905200, 1532908800, 1532912400, 
    1532916000, 1532919600, 1532923200, 1532926800, 1532930400, 1532934000, 
    1532937600, 1532941200, 1532944800, 1532948400, 1532952000, 1532955600, 
    1532959200, 1532962800, 1532966400, 1532970000, 1532973600, 1532977200, 
    1532980800, 1532984400, 1532988000, 1532991600, 1532995200, 1532998800, 
    1533002400, 1533006000, 1533009600, 1533013200, 1533016800, 1533020400, 
    1533024000, 1533027600, 1533031200, 1533034800, 1533038400, 1533042000, 
    1533045600, 1533049200, 1533052800, 1533056400, 1533060000, 1533063600, 
    1533067200, 1533070800, 1533074400, 1533078000, 1533081600, 1533085200, 
    1533088800, 1533092400, 1533096000, 1533099600, 1533103200, 1533106800, 
    1533110400, 1533114000, 1533117600, 1533121200, 1533124800, 1533128400, 
    1533132000, 1533135600, 1533139200, 1533142800, 1533146400, 1533150000, 
    1533153600, 1533157200, 1533160800, 1533164400, 1533168000, 1533171600, 
    1533175200, 1533178800, 1533182400, 1533186000, 1533189600, 1533193200, 
    1533196800, 1533200400, 1533204000, 1533207600, 1533211200, 1533214800, 
    1533218400, 1533222000, 1533225600, 1533229200, 1533232800, 1533236400, 
    1533240000, 1533243600, 1533247200, 1533250800, 1533254400, 1533258000, 
    1533261600, 1533265200, 1533268800, 1533272400, 1533276000, 1533279600, 
    1533283200, 1533286800, 1533290400, 1533294000, 1533297600, 1533301200, 
    1533304800, 1533308400, 1533312000, 1533315600, 1533319200, 1533322800, 
    1533326400, 1533330000, 1533333600, 1533337200, 1533340800, 1533344400, 
    1533348000, 1533351600, 1533355200, 1533358800, 1533362400, 1533366000, 
    1533369600, 1533373200, 1533376800, 1533380400, 1533384000, 1533387600, 
    1533391200, 1533394800, 1533398400, 1533402000, 1533405600, 1533409200, 
    1533412800, 1533416400, 1533420000, 1533423600, 1533427200, 1533430800, 
    1533434400, 1533438000, 1533441600, 1533445200, 1533448800, 1533452400, 
    1533456000, 1533459600, 1533463200, 1533466800, 1533470400, 1533474000, 
    1533477600, 1533481200, 1533484800, 1533488400, 1533492000, 1533495600, 
    1533499200, 1533502800, 1533506400, 1533510000, 1533513600, 1533517200, 
    1533520800, 1533524400, 1533528000, 1533531600, 1533535200, 1533538800, 
    1533542400, 1533546000, 1533549600, 1533553200, 1533556800, 1533560400, 
    1533564000, 1533567600, 1533571200, 1533574800, 1533578400, 1533582000, 
    1533585600, 1533589200, 1533592800, 1533596400, 1533600000, 1533603600, 
    1533607200, 1533610800, 1533614400, 1533618000, 1533621600, 1533625200, 
    1533628800, 1533632400, 1533636000, 1533639600, 1533643200, 1533646800, 
    1533650400, 1533654000, 1533657600, 1533661200, 1533664800, 1533668400, 
    1533672000, 1533675600, 1533679200, 1533682800, 1533686400, 1533690000, 
    1533693600, 1533697200, 1533700800, 1533704400, 1533708000, 1533711600, 
    1533715200, 1533718800, 1533722400, 1533726000, 1533729600, 1533733200, 
    1533736800, 1533740400, 1533744000, 1533747600, 1533751200, 1533754800, 
    1533758400, 1533762000, 1533765600, 1533769200, 1533772800, 1533776400, 
    1533780000, 1533783600, 1533787200, 1533790800, 1533794400, 1533798000, 
    1533801600, 1533805200, 1533808800, 1533812400, 1533816000, 1533819600, 
    1533823200, 1533826800, 1533830400, 1533834000, 1533837600, 1533841200, 
    1533844800, 1533848400, 1533852000, 1533855600, 1533859200, 1533862800, 
    1533866400, 1533870000, 1533873600, 1533877200, 1533880800, 1533884400, 
    1533888000, 1533891600, 1533895200, 1533898800, 1533902400, 1533906000, 
    1533909600, 1533913200, 1533916800, 1533920400, 1533924000, 1533927600, 
    1533931200, 1533934800, 1533938400, 1533942000, 1533945600, 1533949200, 
    1533952800, 1533956400, 1533960000, 1533963600, 1533967200, 1533970800, 
    1533974400, 1533978000, 1533981600, 1533985200, 1533988800, 1533992400, 
    1533996000, 1533999600, 1534003200, 1534006800, 1534010400, 1534014000, 
    1534017600, 1534021200, 1534024800, 1534028400, 1534032000, 1534035600, 
    1534039200, 1534042800, 1534046400, 1534050000, 1534053600, 1534057200, 
    1534060800, 1534064400, 1534068000, 1534071600, 1534075200, 1534078800, 
    1534082400, 1534086000, 1534089600, 1534093200, 1534096800, 1534100400, 
    1534104000, 1534107600, 1534111200, 1534114800, 1534118400, 1534122000, 
    1534125600, 1534129200, 1534132800, 1534136400, 1534140000, 1534143600, 
    1534147200, 1534150800, 1534154400, 1534158000, 1534161600, 1534165200, 
    1534168800, 1534172400, 1534176000, 1534179600, 1534183200, 1534186800, 
    1534190400, 1534194000, 1534197600, 1534201200, 1534204800, 1534208400, 
    1534212000, 1534215600, 1534219200, 1534222800, 1534226400, 1534230000, 
    1534233600, 1534237200, 1534240800, 1534244400, 1534248000, 1534251600, 
    1534255200, 1534258800, 1534262400, 1534266000, 1534269600, 1534273200, 
    1534276800, 1534280400, 1534284000, 1534287600, 1534291200, 1534294800, 
    1534298400, 1534302000, 1534305600, 1534309200, 1534312800, 1534316400, 
    1534320000, 1534323600, 1534327200, 1534330800, 1534334400, 1534338000, 
    1534341600, 1534345200, 1534348800, 1534352400, 1534356000, 1534359600, 
    1534363200, 1534366800, 1534370400, 1534374000, 1534377600, 1534381200, 
    1534384800, 1534388400, 1534392000, 1534395600, 1534399200, 1534402800, 
    1534406400, 1534410000, 1534413600, 1534417200, 1534420800, 1534424400, 
    1534428000, 1534431600, 1534435200, 1534438800, 1534442400, 1534446000, 
    1534449600, 1534453200, 1534456800, 1534460400, 1534464000, 1534467600, 
    1534471200, 1534474800, 1534478400, 1534482000, 1534485600, 1534489200, 
    1534492800, 1534496400, 1534500000, 1534503600, 1534507200, 1534510800, 
    1534514400, 1534518000, 1534521600, 1534525200, 1534528800, 1534532400, 
    1534536000, 1534539600, 1534543200, 1534546800, 1534550400, 1534554000, 
    1534557600, 1534561200, 1534564800, 1534568400, 1534572000, 1534575600, 
    1534579200, 1534582800, 1534586400, 1534590000, 1534593600, 1534597200, 
    1534600800, 1534604400, 1534608000, 1534611600, 1534615200, 1534618800, 
    1534622400, 1534626000, 1534629600, 1534633200, 1534636800, 1534640400, 
    1534644000, 1534647600, 1534651200, 1534654800, 1534658400, 1534662000, 
    1534665600, 1534669200, 1534672800, 1534676400, 1534680000, 1534683600, 
    1534687200, 1534690800, 1534694400, 1534698000, 1534701600, 1534705200, 
    1534708800, 1534712400, 1534716000, 1534719600, 1534723200, 1534726800, 
    1534730400, 1534734000, 1534737600, 1534741200, 1534744800, 1534748400, 
    1534752000, 1534755600, 1534759200, 1534762800, 1534766400, 1534770000, 
    1534773600, 1534777200, 1534780800, 1534784400, 1534788000, 1534791600, 
    1534795200, 1534798800, 1534802400, 1534806000, 1534809600, 1534813200, 
    1534816800, 1534820400, 1534824000, 1534827600, 1534831200, 1534834800, 
    1534838400, 1534842000, 1534845600, 1534849200, 1534852800, 1534856400, 
    1534860000, 1534863600, 1534867200, 1534870800, 1534874400, 1534878000, 
    1534881600, 1534885200, 1534888800, 1534892400, 1534896000, 1534899600, 
    1534903200, 1534906800, 1534910400, 1534914000, 1534917600, 1534921200, 
    1534924800, 1534928400, 1534932000, 1534935600, 1534939200, 1534942800, 
    1534946400, 1534950000, 1534953600, 1534957200, 1534960800, 1534964400, 
    1534968000, 1534971600, 1534975200, 1534978800, 1534982400, 1534986000, 
    1534989600, 1534993200, 1534996800, 1535000400, 1535004000, 1535007600, 
    1535011200, 1535014800, 1535018400, 1535022000, 1535025600, 1535029200, 
    1535032800, 1535036400, 1535040000, 1535043600, 1535047200, 1535050800, 
    1535054400, 1535058000, 1535061600, 1535065200, 1535068800, 1535072400, 
    1535076000, 1535079600, 1535083200, 1535086800, 1535090400, 1535094000, 
    1535097600, 1535101200, 1535104800, 1535108400, 1535112000, 1535115600, 
    1535119200, 1535122800, 1535126400, 1535130000, 1535133600, 1535137200, 
    1535140800, 1535144400, 1535148000, 1535151600, 1535155200, 1535158800, 
    1535162400, 1535166000, 1535169600, 1535173200, 1535176800, 1535180400, 
    1535184000, 1535187600, 1535191200, 1535194800, 1535198400, 1535202000, 
    1535205600, 1535209200, 1535212800, 1535216400, 1535220000, 1535223600, 
    1535227200, 1535230800, 1535234400, 1535238000, 1535241600, 1535245200, 
    1535248800, 1535252400, 1535256000, 1535259600, 1535263200, 1535266800, 
    1535270400, 1535274000, 1535277600, 1535281200, 1535284800, 1535288400, 
    1535292000, 1535295600, 1535299200, 1535302800, 1535306400, 1535310000, 
    1535313600, 1535317200, 1535320800, 1535324400, 1535328000, 1535331600, 
    1535335200, 1535338800, 1535342400, 1535346000, 1535349600, 1535353200, 
    1535356800, 1535360400, 1535364000, 1535367600, 1535371200, 1535374800, 
    1535378400, 1535382000, 1535385600, 1535389200, 1535392800, 1535396400, 
    1535400000, 1535403600, 1535407200, 1535410800, 1535414400, 1535418000, 
    1535421600, 1535425200, 1535428800, 1535432400, 1535436000, 1535439600, 
    1535443200, 1535446800, 1535450400, 1535454000, 1535457600, 1535461200, 
    1535464800, 1535468400, 1535472000, 1535475600, 1535479200, 1535482800, 
    1535486400, 1535490000, 1535493600, 1535497200, 1535500800, 1535504400, 
    1535508000, 1535511600, 1535515200, 1535518800, 1535522400, 1535526000, 
    1535529600, 1535533200, 1535536800, 1535540400, 1535544000, 1535547600, 
    1535551200, 1535554800, 1535558400, 1535562000, 1535565600, 1535569200, 
    1535572800, 1535576400, 1535580000, 1535583600, 1535587200, 1535590800, 
    1535594400, 1535598000, 1535601600, 1535605200, 1535608800, 1535612400, 
    1535616000, 1535619600, 1535623200, 1535626800, 1535630400, 1535634000, 
    1535637600, 1535641200, 1535644800, 1535648400, 1535652000, 1535655600, 
    1535659200, 1535662800, 1535666400, 1535670000, 1535673600, 1535677200, 
    1535680800, 1535684400, 1535688000, 1535691600, 1535695200, 1535698800, 
    1535702400, 1535706000, 1535709600, 1535713200, 1535716800, 1535720400, 
    1535724000, 1535727600, 1535731200, 1535734800, 1535738400, 1535742000, 
    1535745600, 1535749200, 1535752800, 1535756400, 1535760000, 1535763600, 
    1535767200, 1535770800, 1535774400, 1535778000, 1535781600, 1535785200, 
    1535788800, 1535792400, 1535796000, 1535799600, 1535803200, 1535806800, 
    1535810400, 1535814000, 1535817600, 1535821200, 1535824800, 1535828400, 
    1535832000, 1535835600, 1535839200, 1535842800, 1535846400, 1535850000, 
    1535853600, 1535857200, 1535860800, 1535864400, 1535868000, 1535871600, 
    1535875200, 1535878800, 1535882400, 1535886000, 1535889600, 1535893200, 
    1535896800, 1535900400, 1535904000, 1535907600, 1535911200, 1535914800, 
    1535918400, 1535922000, 1535925600, 1535929200, 1535932800, 1535936400, 
    1535940000, 1535943600, 1535947200, 1535950800, 1535954400, 1535958000, 
    1535961600, 1535965200, 1535968800, 1535972400, 1535976000, 1535979600, 
    1535983200, 1535986800, 1535990400, 1535994000, 1535997600, 1536001200, 
    1536004800, 1536008400, 1536012000, 1536015600, 1536019200, 1536022800, 
    1536026400, 1536030000, 1536033600, 1536037200, 1536040800, 1536044400, 
    1536048000, 1536051600, 1536055200, 1536058800, 1536062400, 1536066000, 
    1536069600, 1536073200, 1536076800, 1536080400, 1536084000, 1536087600, 
    1536091200, 1536094800, 1536098400, 1536102000, 1536105600, 1536109200, 
    1536112800, 1536116400, 1536120000, 1536123600, 1536127200, 1536130800, 
    1536134400, 1536138000, 1536141600, 1536145200, 1536148800, 1536152400, 
    1536156000, 1536159600, 1536163200, 1536166800, 1536170400, 1536174000, 
    1536177600, 1536181200, 1536184800, 1536188400, 1536192000, 1536195600, 
    1536199200, 1536202800, 1536206400, 1536210000, 1536213600, 1536217200, 
    1536220800, 1536224400, 1536228000, 1536231600, 1536235200, 1536238800, 
    1536242400, 1536246000, 1536249600, 1536253200, 1536256800, 1536260400, 
    1536264000, 1536267600, 1536271200, 1536274800, 1536278400, 1536282000, 
    1536285600, 1536289200, 1536292800, 1536296400, 1536300000, 1536303600, 
    1536307200, 1536310800, 1536314400, 1536318000, 1536321600, 1536325200, 
    1536328800, 1536332400, 1536336000, 1536339600, 1536343200, 1536346800, 
    1536350400, 1536354000, 1536357600, 1536361200, 1536364800, 1536368400, 
    1536372000, 1536375600, 1536379200, 1536382800, 1536386400, 1536390000, 
    1536393600, 1536397200, 1536400800, 1536404400, 1536408000, 1536411600, 
    1536415200, 1536418800, 1536422400, 1536426000, 1536429600, 1536433200, 
    1536436800, 1536440400, 1536444000, 1536447600, 1536451200, 1536454800, 
    1536458400, 1536462000, 1536465600, 1536469200, 1536472800, 1536476400, 
    1536480000, 1536483600, 1536487200, 1536490800, 1536494400, 1536498000, 
    1536501600, 1536505200, 1536508800, 1536512400, 1536516000, 1536519600, 
    1536523200, 1536526800, 1536530400, 1536534000, 1536537600, 1536541200, 
    1536544800, 1536548400, 1536552000, 1536555600, 1536559200, 1536562800, 
    1536566400, 1536570000, 1536573600, 1536577200, 1536580800, 1536584400, 
    1536588000, 1536591600, 1536595200, 1536598800, 1536602400, 1536606000, 
    1536609600, 1536613200, 1536616800, 1536620400, 1536624000, 1536627600, 
    1536631200, 1536634800, 1536638400, 1536642000, 1536645600, 1536649200, 
    1536652800, 1536656400, 1536660000, 1536663600, 1536667200, 1536670800, 
    1536674400, 1536678000, 1536681600, 1536685200, 1536688800, 1536692400, 
    1536696000, 1536699600, 1536703200, 1536706800, 1536710400, 1536714000, 
    1536717600, 1536721200, 1536724800, 1536728400, 1536732000, 1536735600, 
    1536739200, 1536742800, 1536746400, 1536750000, 1536753600, 1536757200, 
    1536760800, 1536764400, 1536768000, 1536771600, 1536775200, 1536778800, 
    1536782400, 1536786000, 1536789600, 1536793200, 1536796800, 1536800400, 
    1536804000, 1536807600, 1536811200, 1536814800, 1536818400, 1536822000, 
    1536825600, 1536829200, 1536832800, 1536836400, 1536840000, 1536843600, 
    1536847200, 1536850800, 1536854400, 1536858000, 1536861600, 1536865200, 
    1536868800, 1536872400, 1536876000, 1536879600, 1536883200, 1536886800, 
    1536890400, 1536894000, 1536897600, 1536901200, 1536904800, 1536908400, 
    1536912000, 1536915600, 1536919200, 1536922800, 1536926400, 1536930000, 
    1536933600, 1536937200, 1536940800, 1536944400, 1536948000, 1536951600, 
    1536955200, 1536958800, 1536962400, 1536966000, 1536969600, 1536973200, 
    1536976800, 1536980400, 1536984000, 1536987600, 1536991200, 1536994800, 
    1536998400, 1537002000, 1537005600, 1537009200, 1537012800, 1537016400, 
    1537020000, 1537023600, 1537027200, 1537030800, 1537034400, 1537038000, 
    1537041600, 1537045200, 1537048800, 1537052400, 1537056000, 1537059600, 
    1537063200, 1537066800, 1537070400, 1537074000, 1537077600, 1537081200, 
    1537084800, 1537088400, 1537092000, 1537095600, 1537099200, 1537102800, 
    1537106400, 1537110000, 1537113600, 1537117200, 1537120800, 1537124400, 
    1537128000, 1537131600, 1537135200, 1537138800, 1537142400, 1537146000, 
    1537149600, 1537153200, 1537156800, 1537160400, 1537164000, 1537167600, 
    1537171200, 1537174800, 1537178400, 1537182000, 1537185600, 1537189200, 
    1537192800, 1537196400, 1537200000, 1537203600, 1537207200, 1537210800, 
    1537214400, 1537218000, 1537221600, 1537225200, 1537228800, 1537232400, 
    1537236000, 1537239600, 1537243200, 1537246800, 1537250400, 1537254000, 
    1537257600, 1537261200, 1537264800, 1537268400, 1537272000, 1537275600, 
    1537279200, 1537282800, 1537286400, 1537290000, 1537293600, 1537297200, 
    1537300800, 1537304400, 1537308000, 1537311600, 1537315200, 1537318800, 
    1537322400, 1537326000, 1537329600, 1537333200, 1537336800, 1537340400, 
    1537344000, 1537347600, 1537351200, 1537354800, 1537358400, 1537362000, 
    1537365600, 1537369200, 1537372800, 1537376400, 1537380000, 1537383600, 
    1537387200, 1537390800, 1537394400, 1537398000, 1537401600, 1537405200, 
    1537408800, 1537412400, 1537416000, 1537419600, 1537423200, 1537426800, 
    1537430400, 1537434000, 1537437600, 1537441200, 1537444800, 1537448400, 
    1537452000, 1537455600, 1537459200, 1537462800, 1537466400, 1537470000, 
    1537473600, 1537477200, 1537480800, 1537484400, 1537488000, 1537491600, 
    1537495200, 1537498800, 1537502400, 1537506000, 1537509600, 1537513200, 
    1537516800, 1537520400, 1537524000, 1537527600, 1537531200, 1537534800, 
    1537538400, 1537542000, 1537545600, 1537549200, 1537552800, 1537556400, 
    1537560000, 1537563600, 1537567200, 1537570800, 1537574400, 1537578000, 
    1537581600, 1537585200, 1537588800, 1537592400, 1537596000, 1537599600, 
    1537603200, 1537606800, 1537610400, 1537614000, 1537617600, 1537621200, 
    1537624800, 1537628400, 1537632000, 1537635600, 1537639200, 1537642800, 
    1537646400, 1537650000, 1537653600, 1537657200, 1537660800, 1537664400, 
    1537668000, 1537671600, 1537675200, 1537678800, 1537682400, 1537686000, 
    1537689600, 1537693200, 1537696800, 1537700400, 1537704000, 1537707600, 
    1537711200, 1537714800, 1537718400, 1537722000, 1537725600, 1537729200, 
    1537732800, 1537736400, 1537740000, 1537743600, 1537747200, 1537750800, 
    1537754400, 1537758000, 1537761600, 1537765200, 1537768800, 1537772400, 
    1537776000, 1537779600, 1537783200, 1537786800, 1537790400, 1537794000, 
    1537797600, 1537801200, 1537804800, 1537808400, 1537812000, 1537815600, 
    1537819200, 1537822800, 1537826400, 1537830000, 1537833600, 1537837200, 
    1537840800, 1537844400, 1537848000, 1537851600, 1537855200, 1537858800, 
    1537862400, 1537866000, 1537869600, 1537873200, 1537876800, 1537880400, 
    1537884000, 1537887600, 1537891200, 1537894800, 1537898400, 1537902000, 
    1537905600, 1537909200, 1537912800, 1537916400, 1537920000, 1537923600, 
    1537927200, 1537930800, 1537934400, 1537938000, 1537941600, 1537945200, 
    1537948800, 1537952400, 1537956000, 1537959600, 1537963200, 1537966800, 
    1537970400, 1537974000, 1537977600, 1537981200, 1537984800, 1537988400, 
    1537992000, 1537995600, 1537999200, 1538002800, 1538006400, 1538010000, 
    1538013600, 1538017200, 1538020800, 1538024400, 1538028000, 1538031600, 
    1538035200, 1538038800, 1538042400, 1538046000, 1538049600, 1538053200, 
    1538056800, 1538060400, 1538064000, 1538067600, 1538071200, 1538074800, 
    1538078400, 1538082000, 1538085600, 1538089200, 1538092800, 1538096400, 
    1538100000, 1538103600, 1538107200, 1538110800, 1538114400, 1538118000, 
    1538121600, 1538125200, 1538128800, 1538132400, 1538136000, 1538139600, 
    1538143200, 1538146800, 1538150400, 1538154000, 1538157600, 1538161200, 
    1538164800, 1538168400, 1538172000, 1538175600, 1538179200, 1538182800, 
    1538186400, 1538190000, 1538193600, 1538197200, 1538200800, 1538204400, 
    1538208000, 1538211600, 1538215200, 1538218800, 1538222400, 1538226000, 
    1538229600, 1538233200, 1538236800, 1538240400, 1538244000, 1538247600, 
    1538251200, 1538254800, 1538258400, 1538262000, 1538265600, 1538269200, 
    1538272800, 1538276400, 1538280000, 1538283600, 1538287200, 1538290800, 
    1538294400, 1538298000, 1538301600, 1538305200, 1538308800, 1538312400, 
    1538316000, 1538319600, 1538323200, 1538326800, 1538330400, 1538334000, 
    1538337600, 1538341200, 1538344800, 1538348400, 1538352000, 1538355600, 
    1538359200, 1538362800, 1538366400, 1538370000, 1538373600, 1538377200, 
    1538380800, 1538384400, 1538388000, 1538391600, 1538395200, 1538398800, 
    1538402400, 1538406000, 1538409600, 1538413200, 1538416800, 1538420400, 
    1538424000, 1538427600, 1538431200, 1538434800, 1538438400, 1538442000, 
    1538445600, 1538449200, 1538452800, 1538456400, 1538460000, 1538463600, 
    1538467200, 1538470800, 1538474400, 1538478000, 1538481600, 1538485200, 
    1538488800, 1538492400, 1538496000, 1538499600, 1538503200, 1538506800, 
    1538510400, 1538514000, 1538517600, 1538521200, 1538524800, 1538528400, 
    1538532000, 1538535600, 1538539200, 1538542800, 1538546400, 1538550000, 
    1538553600, 1538557200, 1538560800, 1538564400, 1538568000, 1538571600, 
    1538575200, 1538578800, 1538582400, 1538586000, 1538589600, 1538593200, 
    1538596800, 1538600400, 1538604000, 1538607600, 1538611200, 1538614800, 
    1538618400, 1538622000, 1538625600, 1538629200, 1538632800, 1538636400, 
    1538640000, 1538643600, 1538647200, 1538650800, 1538654400, 1538658000, 
    1538661600, 1538665200, 1538668800, 1538672400, 1538676000, 1538679600, 
    1538683200, 1538686800, 1538690400, 1538694000, 1538697600, 1538701200, 
    1538704800, 1538708400, 1538712000, 1538715600, 1538719200, 1538722800, 
    1538726400, 1538730000, 1538733600, 1538737200, 1538740800, 1538744400, 
    1538748000, 1538751600, 1538755200, 1538758800, 1538762400, 1538766000, 
    1538769600, 1538773200, 1538776800, 1538780400, 1538784000, 1538787600, 
    1538791200, 1538794800, 1538798400, 1538802000, 1538805600, 1538809200, 
    1538812800, 1538816400, 1538820000, 1538823600, 1538827200, 1538830800, 
    1538834400, 1538838000, 1538841600, 1538845200, 1538848800, 1538852400, 
    1538856000, 1538859600, 1538863200, 1538866800, 1538870400, 1538874000, 
    1538877600, 1538881200, 1538884800, 1538888400, 1538892000, 1538895600, 
    1538899200, 1538902800, 1538906400, 1538910000, 1538913600, 1538917200, 
    1538920800, 1538924400, 1538928000, 1538931600, 1538935200, 1538938800, 
    1538942400, 1538946000, 1538949600, 1538953200, 1538956800, 1538960400, 
    1538964000, 1538967600, 1538971200, 1538974800, 1538978400, 1538982000, 
    1538985600, 1538989200, 1538992800, 1538996400, 1539000000, 1539003600, 
    1539007200, 1539010800, 1539014400, 1539018000, 1539021600, 1539025200, 
    1539028800, 1539032400, 1539036000, 1539039600, 1539043200, 1539046800, 
    1539050400, 1539054000, 1539057600, 1539061200, 1539064800, 1539068400, 
    1539072000, 1539075600, 1539079200, 1539082800, 1539086400, 1539090000, 
    1539093600, 1539097200, 1539100800, 1539104400, 1539108000, 1539111600, 
    1539115200, 1539118800, 1539122400, 1539126000, 1539129600, 1539133200, 
    1539136800, 1539140400, 1539144000, 1539147600, 1539151200, 1539154800, 
    1539158400, 1539162000, 1539165600, 1539169200, 1539172800, 1539176400, 
    1539180000, 1539183600, 1539187200, 1539190800, 1539194400, 1539198000, 
    1539201600, 1539205200, 1539208800, 1539212400, 1539216000, 1539219600, 
    1539223200, 1539226800, 1539230400, 1539234000, 1539237600, 1539241200, 
    1539244800, 1539248400, 1539252000, 1539255600, 1539259200, 1539262800, 
    1539266400, 1539270000, 1539273600, 1539277200, 1539280800, 1539284400, 
    1539288000, 1539291600, 1539295200, 1539298800, 1539302400, 1539306000, 
    1539309600, 1539313200, 1539316800, 1539320400, 1539324000, 1539327600, 
    1539331200, 1539334800, 1539338400, 1539342000, 1539345600, 1539349200, 
    1539352800, 1539356400, 1539360000, 1539363600, 1539367200, 1539370800, 
    1539374400, 1539378000, 1539381600, 1539385200, 1539388800, 1539392400, 
    1539396000, 1539399600, 1539403200, 1539406800, 1539410400, 1539414000, 
    1539417600, 1539421200, 1539424800, 1539428400, 1539432000, 1539435600, 
    1539439200, 1539442800, 1539446400, 1539450000, 1539453600, 1539457200, 
    1539460800, 1539464400, 1539468000, 1539471600, 1539475200, 1539478800, 
    1539482400, 1539486000, 1539489600, 1539493200, 1539496800, 1539500400, 
    1539504000, 1539507600, 1539511200, 1539514800, 1539518400, 1539522000, 
    1539525600, 1539529200, 1539532800, 1539536400, 1539540000, 1539543600, 
    1539547200, 1539550800, 1539554400, 1539558000, 1539561600, 1539565200, 
    1539568800, 1539572400, 1539576000, 1539579600, 1539583200, 1539586800, 
    1539590400, 1539594000, 1539597600, 1539601200, 1539604800, 1539608400, 
    1539612000, 1539615600, 1539619200, 1539622800, 1539626400, 1539630000, 
    1539633600, 1539637200, 1539640800, 1539644400, 1539648000, 1539651600, 
    1539655200, 1539658800, 1539662400, 1539666000, 1539669600, 1539673200, 
    1539676800, 1539680400, 1539684000, 1539687600, 1539691200, 1539694800, 
    1539698400, 1539702000, 1539705600, 1539709200, 1539712800, 1539716400, 
    1539720000, 1539723600, 1539727200, 1539730800, 1539734400, 1539738000, 
    1539741600, 1539745200, 1539748800, 1539752400, 1539756000, 1539759600, 
    1539763200, 1539766800, 1539770400, 1539774000, 1539777600, 1539781200, 
    1539784800, 1539788400, 1539792000, 1539795600, 1539799200, 1539802800, 
    1539806400, 1539810000, 1539813600, 1539817200, 1539820800, 1539824400, 
    1539828000, 1539831600, 1539835200, 1539838800, 1539842400, 1539846000, 
    1539849600, 1539853200, 1539856800, 1539860400, 1539864000, 1539867600, 
    1539871200, 1539874800, 1539878400, 1539882000, 1539885600, 1539889200, 
    1539892800, 1539896400, 1539900000, 1539903600, 1539907200, 1539910800, 
    1539914400, 1539918000, 1539921600, 1539925200, 1539928800, 1539932400, 
    1539936000, 1539939600, 1539943200, 1539946800, 1539950400, 1539954000, 
    1539957600, 1539961200, 1539964800, 1539968400, 1539972000, 1539975600, 
    1539979200, 1539982800, 1539986400, 1539990000, 1539993600, 1539997200, 
    1540000800, 1540004400, 1540008000, 1540011600, 1540015200, 1540018800, 
    1540022400, 1540026000, 1540029600, 1540033200, 1540036800, 1540040400, 
    1540044000, 1540047600, 1540051200, 1540054800, 1540058400, 1540062000, 
    1540065600, 1540069200, 1540072800, 1540076400, 1540080000, 1540083600, 
    1540087200, 1540090800, 1540094400, 1540098000, 1540101600, 1540105200, 
    1540108800, 1540112400, 1540116000, 1540119600, 1540123200, 1540126800, 
    1540130400, 1540134000, 1540137600, 1540141200, 1540144800, 1540148400, 
    1540152000, 1540155600, 1540159200, 1540162800, 1540166400, 1540170000, 
    1540173600, 1540177200, 1540180800, 1540184400, 1540188000, 1540191600, 
    1540195200, 1540198800, 1540202400, 1540206000, 1540209600, 1540213200, 
    1540216800, 1540220400, 1540224000, 1540227600, 1540231200, 1540234800, 
    1540238400, 1540242000, 1540245600, 1540249200, 1540252800, 1540256400, 
    1540260000, 1540263600, 1540267200, 1540270800, 1540274400, 1540278000, 
    1540281600, 1540285200, 1540288800, 1540292400, 1540296000, 1540299600, 
    1540303200, 1540306800, 1540310400, 1540314000, 1540317600, 1540321200, 
    1540324800, 1540328400, 1540332000, 1540335600, 1540339200, 1540342800, 
    1540346400, 1540350000, 1540353600, 1540357200, 1540360800, 1540364400, 
    1540368000, 1540371600, 1540375200, 1540378800, 1540382400, 1540386000, 
    1540389600, 1540393200, 1540396800, 1540400400, 1540404000, 1540407600, 
    1540411200, 1540414800, 1540418400, 1540422000, 1540425600, 1540429200, 
    1540432800, 1540436400, 1540440000, 1540443600, 1540447200, 1540450800, 
    1540454400, 1540458000, 1540461600, 1540465200, 1540468800, 1540472400, 
    1540476000, 1540479600, 1540483200, 1540486800, 1540490400, 1540494000, 
    1540497600, 1540501200, 1540504800, 1540508400, 1540512000, 1540515600, 
    1540519200, 1540522800, 1540526400, 1540530000, 1540533600, 1540537200, 
    1540540800, 1540544400, 1540548000, 1540551600, 1540555200, 1540558800, 
    1540562400, 1540566000, 1540569600, 1540573200, 1540576800, 1540580400, 
    1540584000, 1540587600, 1540591200, 1540594800, 1540598400, 1540602000, 
    1540605600, 1540609200, 1540612800, 1540616400, 1540620000, 1540623600, 
    1540627200, 1540630800, 1540634400, 1540638000, 1540641600, 1540645200, 
    1540648800, 1540652400, 1540656000, 1540659600, 1540663200, 1540666800, 
    1540670400, 1540674000, 1540677600, 1540681200, 1540684800, 1540688400, 
    1540692000, 1540695600, 1540699200, 1540702800, 1540706400, 1540710000, 
    1540713600, 1540717200, 1540720800, 1540724400, 1540728000, 1540731600, 
    1540735200, 1540738800, 1540742400, 1540746000, 1540749600, 1540753200, 
    1540756800, 1540760400, 1540764000, 1540767600, 1540771200, 1540774800, 
    1540778400, 1540782000, 1540785600, 1540789200, 1540792800, 1540796400, 
    1540800000, 1540803600, 1540807200, 1540810800, 1540814400, 1540818000, 
    1540821600, 1540825200, 1540828800, 1540832400, 1540836000, 1540839600, 
    1540843200, 1540846800, 1540850400, 1540854000, 1540857600, 1540861200, 
    1540864800, 1540868400, 1540872000, 1540875600, 1540879200, 1540882800, 
    1540886400, 1540890000, 1540893600, 1540897200, 1540900800, 1540904400, 
    1540908000, 1540911600, 1540915200, 1540918800, 1540922400, 1540926000, 
    1540929600, 1540933200, 1540936800, 1540940400, 1540944000, 1540947600, 
    1540951200, 1540954800, 1540958400, 1540962000, 1540965600, 1540969200, 
    1540972800, 1540976400, 1540980000, 1540983600, 1540987200, 1540990800, 
    1540994400, 1540998000, 1541001600, 1541005200, 1541008800, 1541012400, 
    1541016000, 1541019600, 1541023200, 1541026800, 1541030400, 1541034000, 
    1541037600, 1541041200, 1541044800, 1541048400, 1541052000, 1541055600, 
    1541059200, 1541062800, 1541066400, 1541070000, 1541073600, 1541077200, 
    1541080800, 1541084400, 1541088000, 1541091600, 1541095200, 1541098800, 
    1541102400, 1541106000, 1541109600, 1541113200, 1541116800, 1541120400, 
    1541124000, 1541127600, 1541131200, 1541134800, 1541138400, 1541142000, 
    1541145600, 1541149200, 1541152800, 1541156400, 1541160000, 1541163600, 
    1541167200, 1541170800, 1541174400, 1541178000, 1541181600, 1541185200, 
    1541188800, 1541192400, 1541196000, 1541199600, 1541203200, 1541206800, 
    1541210400, 1541214000, 1541217600, 1541221200, 1541224800, 1541228400, 
    1541232000, 1541235600, 1541239200, 1541242800, 1541246400, 1541250000, 
    1541253600, 1541257200, 1541260800, 1541264400, 1541268000, 1541271600, 
    1541275200, 1541278800, 1541282400, 1541286000, 1541289600, 1541293200, 
    1541296800, 1541300400, 1541304000, 1541307600, 1541311200, 1541314800, 
    1541318400, 1541322000, 1541325600, 1541329200, 1541332800, 1541336400, 
    1541340000, 1541343600, 1541347200, 1541350800, 1541354400, 1541358000, 
    1541361600, 1541365200, 1541368800, 1541372400, 1541376000, 1541379600, 
    1541383200, 1541386800, 1541390400, 1541394000, 1541397600, 1541401200, 
    1541404800, 1541408400, 1541412000, 1541415600, 1541419200, 1541422800, 
    1541426400, 1541430000, 1541433600, 1541437200, 1541440800, 1541444400, 
    1541448000, 1541451600, 1541455200, 1541458800, 1541462400, 1541466000, 
    1541469600, 1541473200, 1541476800, 1541480400, 1541484000, 1541487600, 
    1541491200, 1541494800, 1541498400, 1541502000, 1541505600, 1541509200, 
    1541512800, 1541516400, 1541520000, 1541523600, 1541527200, 1541530800, 
    1541534400, 1541538000, 1541541600, 1541545200, 1541548800, 1541552400, 
    1541556000, 1541559600, 1541563200, 1541566800, 1541570400, 1541574000, 
    1541577600, 1541581200, 1541584800, 1541588400, 1541592000, 1541595600, 
    1541599200, 1541602800, 1541606400, 1541610000, 1541613600, 1541617200, 
    1541620800, 1541624400, 1541628000, 1541631600, 1541635200, 1541638800, 
    1541642400, 1541646000, 1541649600, 1541653200, 1541656800, 1541660400, 
    1541664000, 1541667600, 1541671200, 1541674800, 1541678400, 1541682000, 
    1541685600, 1541689200, 1541692800, 1541696400, 1541700000, 1541703600, 
    1541707200, 1541710800, 1541714400, 1541718000, 1541721600, 1541725200, 
    1541728800, 1541732400, 1541736000, 1541739600, 1541743200, 1541746800, 
    1541750400, 1541754000, 1541757600, 1541761200, 1541764800, 1541768400, 
    1541772000, 1541775600, 1541779200, 1541782800, 1541786400, 1541790000, 
    1541793600, 1541797200, 1541800800, 1541804400, 1541808000, 1541811600, 
    1541815200, 1541818800, 1541822400, 1541826000, 1541829600, 1541833200, 
    1541836800, 1541840400, 1541844000, 1541847600, 1541851200, 1541854800, 
    1541858400, 1541862000, 1541865600, 1541869200, 1541872800, 1541876400, 
    1541880000, 1541883600, 1541887200, 1541890800, 1541894400, 1541898000, 
    1541901600, 1541905200, 1541908800, 1541912400, 1541916000, 1541919600, 
    1541923200, 1541926800, 1541930400, 1541934000, 1541937600, 1541941200, 
    1541944800, 1541948400, 1541952000, 1541955600, 1541959200, 1541962800, 
    1541966400, 1541970000, 1541973600, 1541977200, 1541980800, 1541984400, 
    1541988000, 1541991600, 1541995200, 1541998800, 1542002400, 1542006000, 
    1542009600, 1542013200, 1542016800, 1542020400, 1542024000, 1542027600, 
    1542031200, 1542034800, 1542038400, 1542042000, 1542045600, 1542049200, 
    1542052800, 1542056400, 1542060000, 1542063600, 1542067200, 1542070800, 
    1542074400, 1542078000, 1542081600, 1542085200, 1542088800, 1542092400, 
    1542096000, 1542099600, 1542103200, 1542106800, 1542110400, 1542114000, 
    1542117600, 1542121200, 1542124800, 1542128400, 1542132000, 1542135600, 
    1542139200, 1542142800, 1542146400, 1542150000, 1542153600, 1542157200, 
    1542160800, 1542164400, 1542168000, 1542171600, 1542175200, 1542178800, 
    1542182400, 1542186000, 1542189600, 1542193200, 1542196800, 1542200400, 
    1542204000, 1542207600, 1542211200, 1542214800, 1542218400, 1542222000, 
    1542225600, 1542229200, 1542232800, 1542236400, 1542240000, 1542243600, 
    1542247200, 1542250800, 1542254400, 1542258000, 1542261600, 1542265200, 
    1542268800, 1542272400, 1542276000, 1542279600, 1542283200, 1542286800, 
    1542290400, 1542294000, 1542297600, 1542301200, 1542304800, 1542308400, 
    1542312000, 1542315600, 1542319200, 1542322800, 1542326400, 1542330000, 
    1542333600, 1542337200, 1542340800, 1542344400, 1542348000, 1542351600, 
    1542355200, 1542358800, 1542362400, 1542366000, 1542369600, 1542373200, 
    1542376800, 1542380400, 1542384000, 1542387600, 1542391200, 1542394800, 
    1542398400, 1542402000, 1542405600, 1542409200, 1542412800, 1542416400, 
    1542420000, 1542423600, 1542427200, 1542430800, 1542434400, 1542438000, 
    1542441600, 1542445200, 1542448800, 1542452400, 1542456000, 1542459600, 
    1542463200, 1542466800, 1542470400, 1542474000, 1542477600, 1542481200, 
    1542484800, 1542488400, 1542492000, 1542495600, 1542499200, 1542502800, 
    1542506400, 1542510000, 1542513600, 1542517200, 1542520800, 1542524400, 
    1542528000, 1542531600, 1542535200, 1542538800, 1542542400, 1542546000, 
    1542549600, 1542553200, 1542556800, 1542560400, 1542564000, 1542567600, 
    1542571200, 1542574800, 1542578400, 1542582000, 1542585600, 1542589200, 
    1542592800, 1542596400, 1542600000, 1542603600, 1542607200, 1542610800, 
    1542614400, 1542618000, 1542621600, 1542625200, 1542628800, 1542632400, 
    1542636000, 1542639600, 1542643200, 1542646800, 1542650400, 1542654000, 
    1542657600, 1542661200, 1542664800, 1542668400, 1542672000, 1542675600, 
    1542679200, 1542682800, 1542686400, 1542690000, 1542693600, 1542697200, 
    1542700800, 1542704400, 1542708000, 1542711600, 1542715200, 1542718800, 
    1542722400, 1542726000, 1542729600, 1542733200, 1542736800, 1542740400, 
    1542744000, 1542747600, 1542751200, 1542754800, 1542758400, 1542762000, 
    1542765600, 1542769200, 1542772800, 1542776400, 1542780000, 1542783600, 
    1542787200, 1542790800, 1542794400, 1542798000, 1542801600, 1542805200, 
    1542808800, 1542812400, 1542816000, 1542819600, 1542823200, 1542826800, 
    1542830400, 1542834000, 1542837600, 1542841200, 1542844800, 1542848400, 
    1542852000, 1542855600, 1542859200, 1542862800, 1542866400, 1542870000, 
    1542873600, 1542877200, 1542880800, 1542884400, 1542888000, 1542891600, 
    1542895200, 1542898800, 1542902400, 1542906000, 1542909600, 1542913200, 
    1542916800, 1542920400, 1542924000, 1542927600, 1542931200, 1542934800, 
    1542938400, 1542942000, 1542945600, 1542949200, 1542952800, 1542956400, 
    1542960000, 1542963600, 1542967200, 1542970800, 1542974400, 1542978000, 
    1542981600, 1542985200, 1542988800, 1542992400, 1542996000, 1542999600, 
    1543003200, 1543006800, 1543010400, 1543014000, 1543017600, 1543021200, 
    1543024800, 1543028400, 1543032000, 1543035600, 1543039200, 1543042800, 
    1543046400, 1543050000, 1543053600, 1543057200, 1543060800, 1543064400, 
    1543068000, 1543071600, 1543075200, 1543078800, 1543082400, 1543086000, 
    1543089600, 1543093200, 1543096800, 1543100400, 1543104000, 1543107600, 
    1543111200, 1543114800, 1543118400, 1543122000, 1543125600, 1543129200, 
    1543132800, 1543136400, 1543140000, 1543143600, 1543147200, 1543150800, 
    1543154400, 1543158000, 1543161600, 1543165200, 1543168800, 1543172400, 
    1543176000, 1543179600, 1543183200, 1543186800, 1543190400, 1543194000, 
    1543197600, 1543201200, 1543204800, 1543208400, 1543212000, 1543215600, 
    1543219200, 1543222800, 1543226400, 1543230000, 1543233600, 1543237200, 
    1543240800, 1543244400, 1543248000, 1543251600, 1543255200, 1543258800, 
    1543262400, 1543266000, 1543269600, 1543273200, 1543276800, 1543280400, 
    1543284000, 1543287600, 1543291200, 1543294800, 1543298400, 1543302000, 
    1543305600, 1543309200, 1543312800, 1543316400, 1543320000, 1543323600, 
    1543327200, 1543330800, 1543334400, 1543338000, 1543341600, 1543345200, 
    1543348800, 1543352400, 1543356000, 1543359600, 1543363200, 1543366800, 
    1543370400, 1543374000, 1543377600, 1543381200, 1543384800, 1543388400, 
    1543392000, 1543395600, 1543399200, 1543402800, 1543406400, 1543410000, 
    1543413600, 1543417200, 1543420800, 1543424400, 1543428000, 1543431600, 
    1543435200, 1543438800, 1543442400, 1543446000, 1543449600, 1543453200, 
    1543456800, 1543460400, 1543464000, 1543467600, 1543471200, 1543474800, 
    1543478400, 1543482000, 1543485600, 1543489200, 1543492800, 1543496400, 
    1543500000, 1543503600, 1543507200, 1543510800, 1543514400, 1543518000, 
    1543521600, 1543525200, 1543528800, 1543532400, 1543536000, 1543539600, 
    1543543200, 1543546800, 1543550400, 1543554000, 1543557600, 1543561200, 
    1543564800, 1543568400, 1543572000, 1543575600, 1543579200, 1543582800, 
    1543586400, 1543590000, 1543593600, 1543597200, 1543600800, 1543604400, 
    1543608000, 1543611600, 1543615200, 1543618800, 1543622400, 1543626000, 
    1543629600, 1543633200, 1543636800, 1543640400, 1543644000, 1543647600, 
    1543651200, 1543654800, 1543658400, 1543662000, 1543665600, 1543669200, 
    1543672800, 1543676400, 1543680000, 1543683600, 1543687200, 1543690800, 
    1543694400, 1543698000, 1543701600, 1543705200, 1543708800, 1543712400, 
    1543716000, 1543719600, 1543723200, 1543726800, 1543730400, 1543734000, 
    1543737600, 1543741200, 1543744800, 1543748400, 1543752000, 1543755600, 
    1543759200, 1543762800, 1543766400, 1543770000, 1543773600, 1543777200, 
    1543780800, 1543784400, 1543788000, 1543791600, 1543795200, 1543798800, 
    1543802400, 1543806000, 1543809600, 1543813200, 1543816800, 1543820400, 
    1543824000, 1543827600, 1543831200, 1543834800, 1543838400, 1543842000, 
    1543845600, 1543849200, 1543852800, 1543856400, 1543860000, 1543863600, 
    1543867200, 1543870800, 1543874400, 1543878000, 1543881600, 1543885200, 
    1543888800, 1543892400, 1543896000, 1543899600, 1543903200, 1543906800, 
    1543910400, 1543914000, 1543917600, 1543921200, 1543924800, 1543928400, 
    1543932000, 1543935600, 1543939200, 1543942800, 1543946400, 1543950000, 
    1543953600, 1543957200, 1543960800, 1543964400, 1543968000, 1543971600, 
    1543975200, 1543978800, 1543982400, 1543986000, 1543989600, 1543993200, 
    1543996800, 1544000400, 1544004000, 1544007600, 1544011200, 1544014800, 
    1544018400, 1544022000, 1544025600, 1544029200, 1544032800, 1544036400, 
    1544040000, 1544043600, 1544047200, 1544050800, 1544054400, 1544058000, 
    1544061600, 1544065200, 1544068800, 1544072400, 1544076000, 1544079600, 
    1544083200, 1544086800, 1544090400, 1544094000, 1544097600, 1544101200, 
    1544104800, 1544108400, 1544112000, 1544115600, 1544119200, 1544122800, 
    1544126400, 1544130000, 1544133600, 1544137200, 1544140800, 1544144400, 
    1544148000, 1544151600, 1544155200, 1544158800, 1544162400, 1544166000, 
    1544169600, 1544173200, 1544176800, 1544180400, 1544184000, 1544187600, 
    1544191200, 1544194800, 1544198400, 1544202000, 1544205600, 1544209200, 
    1544212800, 1544216400, 1544220000, 1544223600, 1544227200, 1544230800, 
    1544234400, 1544238000, 1544241600, 1544245200, 1544248800, 1544252400, 
    1544256000, 1544259600, 1544263200, 1544266800, 1544270400, 1544274000, 
    1544277600, 1544281200, 1544284800, 1544288400, 1544292000, 1544295600, 
    1544299200, 1544302800, 1544306400, 1544310000, 1544313600, 1544317200, 
    1544320800, 1544324400, 1544328000, 1544331600, 1544335200, 1544338800, 
    1544342400, 1544346000, 1544349600, 1544353200, 1544356800, 1544360400, 
    1544364000, 1544367600, 1544371200, 1544374800, 1544378400, 1544382000, 
    1544385600, 1544389200, 1544392800, 1544396400, 1544400000, 1544403600, 
    1544407200, 1544410800, 1544414400, 1544418000, 1544421600, 1544425200, 
    1544428800, 1544432400, 1544436000, 1544439600, 1544443200, 1544446800, 
    1544450400, 1544454000, 1544457600, 1544461200, 1544464800, 1544468400, 
    1544472000, 1544475600, 1544479200, 1544482800, 1544486400, 1544490000, 
    1544493600, 1544497200, 1544500800, 1544504400, 1544508000, 1544511600, 
    1544515200, 1544518800, 1544522400, 1544526000, 1544529600, 1544533200, 
    1544536800, 1544540400, 1544544000, 1544547600, 1544551200, 1544554800, 
    1544558400, 1544562000, 1544565600, 1544569200, 1544572800, 1544576400, 
    1544580000, 1544583600, 1544587200, 1544590800, 1544594400, 1544598000, 
    1544601600, 1544605200, 1544608800, 1544612400, 1544616000, 1544619600, 
    1544623200, 1544626800, 1544630400, 1544634000, 1544637600, 1544641200, 
    1544644800, 1544648400, 1544652000, 1544655600, 1544659200, 1544662800, 
    1544666400, 1544670000, 1544673600, 1544677200, 1544680800, 1544684400, 
    1544688000, 1544691600, 1544695200, 1544698800, 1544702400, 1544706000, 
    1544709600, 1544713200, 1544716800, 1544720400, 1544724000, 1544727600, 
    1544731200, 1544734800, 1544738400, 1544742000, 1544745600, 1544749200, 
    1544752800, 1544756400, 1544760000, 1544763600, 1544767200, 1544770800, 
    1544774400, 1544778000, 1544781600, 1544785200, 1544788800, 1544792400, 
    1544796000, 1544799600, 1544803200, 1544806800, 1544810400, 1544814000, 
    1544817600, 1544821200, 1544824800, 1544828400, 1544832000, 1544835600, 
    1544839200, 1544842800, 1544846400, 1544850000, 1544853600, 1544857200, 
    1544860800, 1544864400, 1544868000, 1544871600, 1544875200, 1544878800, 
    1544882400, 1544886000, 1544889600, 1544893200, 1544896800, 1544900400, 
    1544904000, 1544907600, 1544911200, 1544914800, 1544918400, 1544922000, 
    1544925600, 1544929200, 1544932800, 1544936400, 1544940000, 1544943600, 
    1544947200, 1544950800, 1544954400, 1544958000, 1544961600, 1544965200, 
    1544968800, 1544972400, 1544976000, 1544979600, 1544983200, 1544986800, 
    1544990400, 1544994000, 1544997600, 1545001200, 1545004800, 1545008400, 
    1545012000, 1545015600, 1545019200, 1545022800, 1545026400, 1545030000, 
    1545033600, 1545037200, 1545040800, 1545044400, 1545048000, 1545051600, 
    1545055200, 1545058800, 1545062400, 1545066000, 1545069600, 1545073200, 
    1545076800, 1545080400, 1545084000, 1545087600, 1545091200, 1545094800, 
    1545098400, 1545102000, 1545105600, 1545109200, 1545112800, 1545116400, 
    1545120000, 1545123600, 1545127200, 1545130800, 1545134400, 1545138000, 
    1545141600, 1545145200, 1545148800, 1545152400, 1545156000, 1545159600, 
    1545163200, 1545166800, 1545170400, 1545174000, 1545177600, 1545181200, 
    1545184800, 1545188400, 1545192000, 1545195600, 1545199200, 1545202800, 
    1545206400, 1545210000, 1545213600, 1545217200, 1545220800, 1545224400, 
    1545228000, 1545231600, 1545235200, 1545238800, 1545242400, 1545246000, 
    1545249600, 1545253200, 1545256800, 1545260400, 1545264000, 1545267600, 
    1545271200, 1545274800, 1545278400, 1545282000, 1545285600, 1545289200, 
    1545292800, 1545296400, 1545300000, 1545303600, 1545307200, 1545310800, 
    1545314400, 1545318000, 1545321600, 1545325200, 1545328800, 1545332400, 
    1545336000, 1545339600, 1545343200, 1545346800, 1545350400, 1545354000, 
    1545357600, 1545361200, 1545364800, 1545368400, 1545372000, 1545375600, 
    1545379200, 1545382800, 1545386400, 1545390000, 1545393600, 1545397200, 
    1545400800, 1545404400, 1545408000, 1545411600, 1545415200, 1545418800, 
    1545422400, 1545426000, 1545429600, 1545433200, 1545436800, 1545440400, 
    1545444000, 1545447600, 1545451200, 1545454800, 1545458400, 1545462000, 
    1545465600, 1545469200, 1545472800, 1545476400, 1545480000, 1545483600, 
    1545487200, 1545490800, 1545494400, 1545498000, 1545501600, 1545505200, 
    1545508800, 1545512400, 1545516000, 1545519600, 1545523200, 1545526800, 
    1545530400, 1545534000, 1545537600, 1545541200, 1545544800, 1545548400, 
    1545552000, 1545555600, 1545559200, 1545562800, 1545566400, 1545570000, 
    1545573600, 1545577200, 1545580800, 1545584400, 1545588000, 1545591600, 
    1545595200, 1545598800, 1545602400, 1545606000, 1545609600, 1545613200, 
    1545616800, 1545620400, 1545624000, 1545627600, 1545631200, 1545634800, 
    1545638400, 1545642000, 1545645600, 1545649200, 1545652800, 1545656400, 
    1545660000, 1545663600, 1545667200, 1545670800, 1545674400, 1545678000, 
    1545681600, 1545685200, 1545688800, 1545692400, 1545696000, 1545699600, 
    1545703200, 1545706800, 1545710400, 1545714000, 1545717600, 1545721200, 
    1545724800, 1545728400, 1545732000, 1545735600, 1545739200, 1545742800, 
    1545746400, 1545750000, 1545753600, 1545757200, 1545760800, 1545764400, 
    1545768000, 1545771600, 1545775200, 1545778800, 1545782400, 1545786000, 
    1545789600, 1545793200, 1545796800, 1545800400, 1545804000, 1545807600, 
    1545811200, 1545814800, 1545818400, 1545822000, 1545825600, 1545829200, 
    1545832800, 1545836400, 1545840000, 1545843600, 1545847200, 1545850800, 
    1545854400, 1545858000, 1545861600, 1545865200, 1545868800, 1545872400, 
    1545876000, 1545879600, 1545883200, 1545886800, 1545890400, 1545894000, 
    1545897600, 1545901200, 1545904800, 1545908400, 1545912000, 1545915600, 
    1545919200, 1545922800, 1545926400, 1545930000, 1545933600, 1545937200, 
    1545940800, 1545944400, 1545948000, 1545951600, 1545955200, 1545958800, 
    1545962400, 1545966000, 1545969600, 1545973200, 1545976800, 1545980400, 
    1545984000, 1545987600, 1545991200, 1545994800, 1545998400, 1546002000, 
    1546005600, 1546009200, 1546012800, 1546016400, 1546020000, 1546023600, 
    1546027200, 1546030800, 1546034400, 1546038000, 1546041600, 1546045200, 
    1546048800, 1546052400, 1546056000, 1546059600, 1546063200, 1546066800, 
    1546070400, 1546074000, 1546077600, 1546081200, 1546084800, 1546088400, 
    1546092000, 1546095600, 1546099200, 1546102800, 1546106400, 1546110000, 
    1546113600, 1546117200, 1546120800, 1546124400, 1546128000, 1546131600, 
    1546135200, 1546138800, 1546142400, 1546146000, 1546149600, 1546153200, 
    1546156800, 1546160400, 1546164000, 1546167600, 1546171200, 1546174800, 
    1546178400, 1546182000, 1546185600, 1546189200, 1546192800, 1546196400, 
    1546200000, 1546203600, 1546207200, 1546210800, 1546214400, 1546218000, 
    1546221600, 1546225200, 1546228800, 1546232400, 1546236000, 1546239600, 
    1546243200, 1546246800, 1546250400, 1546254000, 1546257600, 1546261200, 
    1546264800, 1546268400, 1546272000, 1546275600, 1546279200, 1546282800, 
    1546286400, 1546290000, 1546293600, 1546297200, 1546300800, 1546304400, 
    1546308000, 1546311600, 1546315200, 1546318800, 1546322400, 1546326000, 
    1546329600, 1546333200, 1546336800, 1546340400, 1546344000, 1546347600, 
    1546351200, 1546354800, 1546358400, 1546362000, 1546365600, 1546369200, 
    1546372800, 1546376400, 1546380000, 1546383600, 1546387200, 1546390800, 
    1546394400, 1546398000, 1546401600, 1546405200, 1546408800, 1546412400, 
    1546416000, 1546419600, 1546423200, 1546426800, 1546430400, 1546434000, 
    1546437600, 1546441200, 1546444800, 1546448400, 1546452000, 1546455600, 
    1546459200, 1546462800, 1546466400, 1546470000, 1546473600, 1546477200, 
    1546480800, 1546484400, 1546488000, 1546491600, 1546495200, 1546498800, 
    1546502400, 1546506000, 1546509600, 1546513200, 1546516800, 1546520400, 
    1546524000, 1546527600, 1546531200, 1546534800, 1546538400, 1546542000, 
    1546545600, 1546549200, 1546552800, 1546556400, 1546560000, 1546563600, 
    1546567200, 1546570800, 1546574400, 1546578000, 1546581600, 1546585200, 
    1546588800, 1546592400, 1546596000, 1546599600, 1546603200, 1546606800, 
    1546610400, 1546614000, 1546617600, 1546621200, 1546624800, 1546628400, 
    1546632000, 1546635600, 1546639200, 1546642800, 1546646400, 1546650000, 
    1546653600, 1546657200, 1546660800, 1546664400, 1546668000, 1546671600, 
    1546675200, 1546678800, 1546682400, 1546686000, 1546689600, 1546693200, 
    1546696800, 1546700400, 1546704000, 1546707600, 1546711200, 1546714800, 
    1546718400, 1546722000, 1546725600, 1546729200, 1546732800, 1546736400, 
    1546740000, 1546743600, 1546747200, 1546750800, 1546754400, 1546758000, 
    1546761600, 1546765200, 1546768800, 1546772400, 1546776000, 1546779600, 
    1546783200, 1546786800, 1546790400, 1546794000, 1546797600, 1546801200, 
    1546804800, 1546808400, 1546812000, 1546815600, 1546819200, 1546822800, 
    1546826400, 1546830000, 1546833600, 1546837200, 1546840800, 1546844400, 
    1546848000, 1546851600, 1546855200, 1546858800, 1546862400, 1546866000, 
    1546869600, 1546873200, 1546876800, 1546880400, 1546884000, 1546887600, 
    1546891200, 1546894800, 1546898400, 1546902000, 1546905600, 1546909200, 
    1546912800, 1546916400, 1546920000, 1546923600, 1546927200, 1546930800, 
    1546934400, 1546938000, 1546941600, 1546945200, 1546948800, 1546952400, 
    1546956000, 1546959600, 1546963200, 1546966800, 1546970400, 1546974000, 
    1546977600, 1546981200, 1546984800, 1546988400, 1546992000, 1546995600, 
    1546999200, 1547002800, 1547006400, 1547010000, 1547013600, 1547017200, 
    1547020800, 1547024400, 1547028000, 1547031600, 1547035200, 1547038800, 
    1547042400, 1547046000, 1547049600, 1547053200, 1547056800, 1547060400, 
    1547064000, 1547067600, 1547071200, 1547074800, 1547078400, 1547082000, 
    1547085600, 1547089200, 1547092800, 1547096400, 1547100000, 1547103600, 
    1547107200, 1547110800, 1547114400, 1547118000, 1547121600, 1547125200, 
    1547128800, 1547132400, 1547136000, 1547139600, 1547143200, 1547146800, 
    1547150400, 1547154000, 1547157600, 1547161200, 1547164800, 1547168400, 
    1547172000, 1547175600, 1547179200, 1547182800, 1547186400, 1547190000, 
    1547193600, 1547197200, 1547200800, 1547204400, 1547208000, 1547211600, 
    1547215200, 1547218800, 1547222400, 1547226000, 1547229600, 1547233200, 
    1547236800, 1547240400, 1547244000, 1547247600, 1547251200, 1547254800, 
    1547258400, 1547262000, 1547265600, 1547269200, 1547272800, 1547276400, 
    1547280000, 1547283600, 1547287200, 1547290800, 1547294400, 1547298000, 
    1547301600, 1547305200, 1547308800, 1547312400, 1547316000, 1547319600, 
    1547323200, 1547326800, 1547330400, 1547334000, 1547337600, 1547341200, 
    1547344800, 1547348400, 1547352000, 1547355600, 1547359200, 1547362800, 
    1547366400, 1547370000, 1547373600, 1547377200, 1547380800, 1547384400, 
    1547388000, 1547391600, 1547395200, 1547398800, 1547402400, 1547406000, 
    1547409600, 1547413200, 1547416800, 1547420400, 1547424000, 1547427600, 
    1547431200, 1547434800, 1547438400, 1547442000, 1547445600, 1547449200, 
    1547452800, 1547456400, 1547460000, 1547463600, 1547467200, 1547470800, 
    1547474400, 1547478000, 1547481600, 1547485200, 1547488800, 1547492400, 
    1547496000, 1547499600, 1547503200, 1547506800, 1547510400, 1547514000, 
    1547517600, 1547521200, 1547524800, 1547528400, 1547532000, 1547535600, 
    1547539200, 1547542800, 1547546400, 1547550000, 1547553600, 1547557200, 
    1547560800, 1547564400, 1547568000, 1547571600, 1547575200, 1547578800, 
    1547582400, 1547586000, 1547589600, 1547593200, 1547596800, 1547600400, 
    1547604000, 1547607600, 1547611200, 1547614800, 1547618400, 1547622000, 
    1547625600, 1547629200, 1547632800, 1547636400, 1547640000, 1547643600, 
    1547647200, 1547650800, 1547654400, 1547658000, 1547661600, 1547665200, 
    1547668800, 1547672400, 1547676000, 1547679600, 1547683200, 1547686800, 
    1547690400, 1547694000, 1547697600, 1547701200, 1547704800, 1547708400, 
    1547712000, 1547715600, 1547719200, 1547722800, 1547726400, 1547730000, 
    1547733600, 1547737200, 1547740800, 1547744400, 1547748000, 1547751600, 
    1547755200, 1547758800, 1547762400, 1547766000, 1547769600, 1547773200, 
    1547776800, 1547780400, 1547784000, 1547787600, 1547791200, 1547794800, 
    1547798400, 1547802000, 1547805600, 1547809200, 1547812800, 1547816400, 
    1547820000, 1547823600, 1547827200, 1547830800, 1547834400, 1547838000, 
    1547841600, 1547845200, 1547848800, 1547852400, 1547856000, 1547859600, 
    1547863200, 1547866800, 1547870400, 1547874000, 1547877600, 1547881200, 
    1547884800, 1547888400, 1547892000, 1547895600, 1547899200, 1547902800, 
    1547906400, 1547910000, 1547913600, 1547917200, 1547920800, 1547924400, 
    1547928000, 1547931600, 1547935200, 1547938800, 1547942400, 1547946000, 
    1547949600, 1547953200, 1547956800, 1547960400, 1547964000, 1547967600, 
    1547971200, 1547974800, 1547978400, 1547982000, 1547985600, 1547989200, 
    1547992800, 1547996400, 1548000000, 1548003600, 1548007200, 1548010800, 
    1548014400, 1548018000, 1548021600, 1548025200, 1548028800, 1548032400, 
    1548036000, 1548039600, 1548043200, 1548046800, 1548050400, 1548054000, 
    1548057600, 1548061200, 1548064800, 1548068400, 1548072000, 1548075600, 
    1548079200, 1548082800, 1548086400, 1548090000, 1548093600, 1548097200, 
    1548100800, 1548104400, 1548108000, 1548111600, 1548115200, 1548118800, 
    1548122400, 1548126000, 1548129600, 1548133200, 1548136800, 1548140400, 
    1548144000, 1548147600, 1548151200, 1548154800, 1548158400, 1548162000, 
    1548165600, 1548169200, 1548172800, 1548176400, 1548180000, 1548183600, 
    1548187200, 1548190800, 1548194400, 1548198000, 1548201600, 1548205200, 
    1548208800, 1548212400, 1548216000, 1548219600, 1548223200, 1548226800, 
    1548230400, 1548234000, 1548237600, 1548241200, 1548244800, 1548248400, 
    1548252000, 1548255600, 1548259200, 1548262800, 1548266400, 1548270000, 
    1548273600, 1548277200, 1548280800, 1548284400, 1548288000, 1548291600, 
    1548295200, 1548298800, 1548302400, 1548306000, 1548309600, 1548313200, 
    1548316800, 1548320400, 1548324000, 1548327600, 1548331200, 1548334800, 
    1548338400, 1548342000, 1548345600, 1548349200, 1548352800, 1548356400, 
    1548360000, 1548363600, 1548367200, 1548370800, 1548374400, 1548378000, 
    1548381600, 1548385200, 1548388800, 1548392400, 1548396000, 1548399600, 
    1548403200, 1548406800, 1548410400, 1548414000, 1548417600, 1548421200, 
    1548424800, 1548428400, 1548432000, 1548435600, 1548439200, 1548442800, 
    1548446400, 1548450000, 1548453600, 1548457200, 1548460800, 1548464400, 
    1548468000, 1548471600, 1548475200, 1548478800, 1548482400, 1548486000, 
    1548489600, 1548493200, 1548496800, 1548500400, 1548504000, 1548507600, 
    1548511200, 1548514800, 1548518400, 1548522000, 1548525600, 1548529200, 
    1548532800, 1548536400, 1548540000, 1548543600, 1548547200, 1548550800, 
    1548554400, 1548558000, 1548561600, 1548565200, 1548568800, 1548572400, 
    1548576000, 1548579600, 1548583200, 1548586800, 1548590400, 1548594000, 
    1548597600, 1548601200, 1548604800, 1548608400, 1548612000, 1548615600, 
    1548619200, 1548622800, 1548626400, 1548630000, 1548633600, 1548637200, 
    1548640800, 1548644400, 1548648000, 1548651600, 1548655200, 1548658800, 
    1548662400, 1548666000, 1548669600, 1548673200, 1548676800, 1548680400, 
    1548684000, 1548687600, 1548691200, 1548694800, 1548698400, 1548702000, 
    1548705600, 1548709200, 1548712800, 1548716400, 1548720000, 1548723600, 
    1548727200, 1548730800, 1548734400, 1548738000, 1548741600, 1548745200, 
    1548748800, 1548752400, 1548756000, 1548759600, 1548763200, 1548766800, 
    1548770400, 1548774000, 1548777600, 1548781200, 1548784800, 1548788400, 
    1548792000, 1548795600, 1548799200, 1548802800, 1548806400, 1548810000, 
    1548813600, 1548817200, 1548820800, 1548824400, 1548828000, 1548831600, 
    1548835200, 1548838800, 1548842400, 1548846000, 1548849600, 1548853200, 
    1548856800, 1548860400, 1548864000, 1548867600, 1548871200, 1548874800, 
    1548878400, 1548882000, 1548885600, 1548889200, 1548892800, 1548896400, 
    1548900000, 1548903600, 1548907200, 1548910800, 1548914400, 1548918000, 
    1548921600, 1548925200, 1548928800, 1548932400, 1548936000, 1548939600, 
    1548943200, 1548946800, 1548950400, 1548954000, 1548957600, 1548961200, 
    1548964800, 1548968400, 1548972000, 1548975600, 1548979200, 1548982800, 
    1548986400, 1548990000, 1548993600, 1548997200, 1549000800, 1549004400, 
    1549008000, 1549011600, 1549015200, 1549018800, 1549022400, 1549026000, 
    1549029600, 1549033200, 1549036800, 1549040400, 1549044000, 1549047600, 
    1549051200, 1549054800, 1549058400, 1549062000, 1549065600, 1549069200, 
    1549072800, 1549076400, 1549080000, 1549083600, 1549087200, 1549090800, 
    1549094400, 1549098000, 1549101600, 1549105200, 1549108800, 1549112400, 
    1549116000, 1549119600, 1549123200, 1549126800, 1549130400, 1549134000, 
    1549137600, 1549141200, 1549144800, 1549148400, 1549152000, 1549155600, 
    1549159200, 1549162800, 1549166400, 1549170000, 1549173600, 1549177200, 
    1549180800, 1549184400, 1549188000, 1549191600, 1549195200, 1549198800, 
    1549202400, 1549206000, 1549209600, 1549213200, 1549216800, 1549220400, 
    1549224000, 1549227600, 1549231200, 1549234800, 1549238400, 1549242000, 
    1549245600, 1549249200, 1549252800, 1549256400, 1549260000, 1549263600, 
    1549267200, 1549270800, 1549274400, 1549278000, 1549281600, 1549285200, 
    1549288800, 1549292400, 1549296000, 1549299600, 1549303200, 1549306800, 
    1549310400, 1549314000, 1549317600, 1549321200, 1549324800, 1549328400, 
    1549332000, 1549335600, 1549339200, 1549342800, 1549346400, 1549350000, 
    1549353600, 1549357200, 1549360800, 1549364400, 1549368000, 1549371600, 
    1549375200, 1549378800, 1549382400, 1549386000, 1549389600, 1549393200, 
    1549396800, 1549400400, 1549404000, 1549407600, 1549411200, 1549414800, 
    1549418400, 1549422000, 1549425600, 1549429200, 1549432800, 1549436400, 
    1549440000, 1549443600, 1549447200, 1549450800, 1549454400, 1549458000, 
    1549461600, 1549465200, 1549468800, 1549472400, 1549476000, 1549479600, 
    1549483200, 1549486800, 1549490400, 1549494000, 1549497600, 1549501200, 
    1549504800, 1549508400, 1549512000, 1549515600, 1549519200, 1549522800, 
    1549526400, 1549530000, 1549533600, 1549537200, 1549540800, 1549544400, 
    1549548000, 1549551600, 1549555200, 1549558800, 1549562400, 1549566000, 
    1549569600, 1549573200, 1549576800, 1549580400, 1549584000, 1549587600, 
    1549591200, 1549594800, 1549598400, 1549602000, 1549605600, 1549609200, 
    1549612800, 1549616400, 1549620000, 1549623600, 1549627200, 1549630800, 
    1549634400, 1549638000, 1549641600, 1549645200, 1549648800, 1549652400, 
    1549656000, 1549659600, 1549663200, 1549666800, 1549670400, 1549674000, 
    1549677600, 1549681200, 1549684800, 1549688400, 1549692000, 1549695600, 
    1549699200, 1549702800, 1549706400, 1549710000, 1549713600, 1549717200, 
    1549720800, 1549724400, 1549728000, 1549731600, 1549735200, 1549738800, 
    1549742400, 1549746000, 1549749600, 1549753200, 1549756800, 1549760400, 
    1549764000, 1549767600, 1549771200, 1549774800, 1549778400, 1549782000, 
    1549785600, 1549789200, 1549792800, 1549796400, 1549800000, 1549803600, 
    1549807200, 1549810800, 1549814400, 1549818000, 1549821600, 1549825200, 
    1549828800, 1549832400, 1549836000, 1549839600, 1549843200, 1549846800, 
    1549850400, 1549854000, 1549857600, 1549861200, 1549864800, 1549868400, 
    1549872000, 1549875600, 1549879200, 1549882800, 1549886400, 1549890000, 
    1549893600, 1549897200, 1549900800, 1549904400, 1549908000, 1549911600, 
    1549915200, 1549918800, 1549922400, 1549926000, 1549929600, 1549933200, 
    1549936800, 1549940400, 1549944000, 1549947600, 1549951200, 1549954800, 
    1549958400, 1549962000, 1549965600, 1549969200, 1549972800, 1549976400, 
    1549980000, 1549983600, 1549987200, 1549990800, 1549994400, 1549998000, 
    1550001600, 1550005200, 1550008800, 1550012400, 1550016000, 1550019600, 
    1550023200, 1550026800, 1550030400, 1550034000, 1550037600, 1550041200, 
    1550044800, 1550048400, 1550052000, 1550055600, 1550059200, 1550062800, 
    1550066400, 1550070000, 1550073600, 1550077200, 1550080800, 1550084400, 
    1550088000, 1550091600, 1550095200, 1550098800, 1550102400, 1550106000, 
    1550109600, 1550113200, 1550116800, 1550120400, 1550124000, 1550127600, 
    1550131200, 1550134800, 1550138400, 1550142000, 1550145600, 1550149200, 
    1550152800, 1550156400, 1550160000, 1550163600, 1550167200, 1550170800, 
    1550174400, 1550178000, 1550181600, 1550185200, 1550188800, 1550192400, 
    1550196000, 1550199600, 1550203200, 1550206800, 1550210400, 1550214000, 
    1550217600, 1550221200, 1550224800, 1550228400, 1550232000, 1550235600, 
    1550239200, 1550242800, 1550246400, 1550250000, 1550253600, 1550257200, 
    1550260800, 1550264400, 1550268000, 1550271600, 1550275200, 1550278800, 
    1550282400, 1550286000, 1550289600, 1550293200, 1550296800, 1550300400, 
    1550304000, 1550307600, 1550311200, 1550314800, 1550318400, 1550322000, 
    1550325600, 1550329200, 1550332800, 1550336400, 1550340000, 1550343600, 
    1550347200, 1550350800, 1550354400, 1550358000, 1550361600, 1550365200, 
    1550368800, 1550372400, 1550376000, 1550379600, 1550383200, 1550386800, 
    1550390400, 1550394000, 1550397600, 1550401200, 1550404800, 1550408400, 
    1550412000, 1550415600, 1550419200, 1550422800, 1550426400, 1550430000, 
    1550433600, 1550437200, 1550440800, 1550444400, 1550448000, 1550451600, 
    1550455200, 1550458800, 1550462400, 1550466000, 1550469600, 1550473200, 
    1550476800, 1550480400, 1550484000, 1550487600, 1550491200, 1550494800, 
    1550498400, 1550502000, 1550505600, 1550509200, 1550512800, 1550516400, 
    1550520000, 1550523600, 1550527200, 1550530800, 1550534400, 1550538000, 
    1550541600, 1550545200, 1550548800, 1550552400, 1550556000, 1550559600, 
    1550563200, 1550566800, 1550570400, 1550574000, 1550577600, 1550581200, 
    1550584800, 1550588400, 1550592000, 1550595600, 1550599200, 1550602800, 
    1550606400, 1550610000, 1550613600, 1550617200, 1550620800, 1550624400, 
    1550628000, 1550631600, 1550635200, 1550638800, 1550642400, 1550646000, 
    1550649600, 1550653200, 1550656800, 1550660400, 1550664000, 1550667600, 
    1550671200, 1550674800, 1550678400, 1550682000, 1550685600, 1550689200, 
    1550692800, 1550696400, 1550700000, 1550703600, 1550707200, 1550710800, 
    1550714400, 1550718000, 1550721600, 1550725200, 1550728800, 1550732400, 
    1550736000, 1550739600, 1550743200, 1550746800, 1550750400, 1550754000, 
    1550757600, 1550761200, 1550764800, 1550768400, 1550772000, 1550775600, 
    1550779200, 1550782800, 1550786400, 1550790000, 1550793600, 1550797200, 
    1550800800, 1550804400, 1550808000, 1550811600, 1550815200, 1550818800, 
    1550822400, 1550826000, 1550829600, 1550833200, 1550836800, 1550840400, 
    1550844000, 1550847600, 1550851200, 1550854800, 1550858400, 1550862000, 
    1550865600, 1550869200, 1550872800, 1550876400, 1550880000, 1550883600, 
    1550887200, 1550890800, 1550894400, 1550898000, 1550901600, 1550905200, 
    1550908800, 1550912400, 1550916000, 1550919600, 1550923200, 1550926800, 
    1550930400, 1550934000, 1550937600, 1550941200, 1550944800, 1550948400, 
    1550952000, 1550955600, 1550959200, 1550962800, 1550966400, 1550970000, 
    1550973600, 1550977200, 1550980800, 1550984400, 1550988000, 1550991600, 
    1550995200, 1550998800, 1551002400, 1551006000, 1551009600, 1551013200, 
    1551016800, 1551020400, 1551024000, 1551027600, 1551031200, 1551034800, 
    1551038400, 1551042000, 1551045600, 1551049200, 1551052800, 1551056400, 
    1551060000, 1551063600, 1551067200, 1551070800, 1551074400, 1551078000, 
    1551081600, 1551085200, 1551088800, 1551092400, 1551096000, 1551099600, 
    1551103200, 1551106800, 1551110400, 1551114000, 1551117600, 1551121200, 
    1551124800, 1551128400, 1551132000, 1551135600, 1551139200, 1551142800, 
    1551146400, 1551150000, 1551153600, 1551157200, 1551160800, 1551164400, 
    1551168000, 1551171600, 1551175200, 1551178800, 1551182400, 1551186000, 
    1551189600, 1551193200, 1551196800, 1551200400, 1551204000, 1551207600, 
    1551211200, 1551214800, 1551218400, 1551222000, 1551225600, 1551229200, 
    1551232800, 1551236400, 1551240000, 1551243600, 1551247200, 1551250800, 
    1551254400, 1551258000, 1551261600, 1551265200, 1551268800, 1551272400, 
    1551276000, 1551279600, 1551283200, 1551286800, 1551290400, 1551294000, 
    1551297600, 1551301200, 1551304800, 1551308400, 1551312000, 1551315600, 
    1551319200, 1551322800, 1551326400, 1551330000, 1551333600, 1551337200, 
    1551340800, 1551344400, 1551348000, 1551351600, 1551355200, 1551358800, 
    1551362400, 1551366000, 1551369600, 1551373200, 1551376800, 1551380400, 
    1551384000, 1551387600, 1551391200, 1551394800, 1551398400, 1551402000, 
    1551405600, 1551409200, 1551412800, 1551416400, 1551420000, 1551423600, 
    1551427200, 1551430800, 1551434400, 1551438000, 1551441600, 1551445200, 
    1551448800, 1551452400, 1551456000, 1551459600, 1551463200, 1551466800, 
    1551470400, 1551474000, 1551477600, 1551481200, 1551484800, 1551488400, 
    1551492000, 1551495600, 1551499200, 1551502800, 1551506400, 1551510000, 
    1551513600, 1551517200, 1551520800, 1551524400, 1551528000, 1551531600, 
    1551535200, 1551538800, 1551542400, 1551546000, 1551549600, 1551553200, 
    1551556800, 1551560400, 1551564000, 1551567600, 1551571200, 1551574800, 
    1551578400, 1551582000, 1551585600, 1551589200, 1551592800, 1551596400, 
    1551600000, 1551603600, 1551607200, 1551610800, 1551614400, 1551618000, 
    1551621600, 1551625200, 1551628800, 1551632400, 1551636000, 1551639600, 
    1551643200, 1551646800, 1551650400, 1551654000, 1551657600, 1551661200, 
    1551664800, 1551668400, 1551672000, 1551675600, 1551679200, 1551682800, 
    1551686400, 1551690000, 1551693600, 1551697200, 1551700800, 1551704400, 
    1551708000, 1551711600, 1551715200, 1551718800, 1551722400, 1551726000, 
    1551729600, 1551733200, 1551736800, 1551740400, 1551744000, 1551747600, 
    1551751200, 1551754800, 1551758400, 1551762000, 1551765600, 1551769200, 
    1551772800, 1551776400, 1551780000, 1551783600, 1551787200, 1551790800, 
    1551794400, 1551798000, 1551801600, 1551805200, 1551808800, 1551812400, 
    1551816000, 1551819600, 1551823200, 1551826800, 1551830400, 1551834000, 
    1551837600, 1551841200, 1551844800, 1551848400, 1551852000, 1551855600, 
    1551859200, 1551862800, 1551866400, 1551870000, 1551873600, 1551877200, 
    1551880800, 1551884400, 1551888000, 1551891600, 1551895200, 1551898800, 
    1551902400, 1551906000, 1551909600, 1551913200, 1551916800, 1551920400, 
    1551924000, 1551927600, 1551931200, 1551934800, 1551938400, 1551942000, 
    1551945600, 1551949200, 1551952800, 1551956400, 1551960000, 1551963600, 
    1551967200, 1551970800, 1551974400, 1551978000, 1551981600, 1551985200, 
    1551988800, 1551992400, 1551996000, 1551999600, 1552003200, 1552006800, 
    1552010400, 1552014000, 1552017600, 1552021200, 1552024800, 1552028400, 
    1552032000, 1552035600, 1552039200, 1552042800, 1552046400, 1552050000, 
    1552053600, 1552057200, 1552060800, 1552064400, 1552068000, 1552071600, 
    1552075200, 1552078800, 1552082400, 1552086000, 1552089600, 1552093200, 
    1552096800, 1552100400, 1552104000, 1552107600, 1552111200, 1552114800, 
    1552118400, 1552122000, 1552125600, 1552129200, 1552132800, 1552136400, 
    1552140000, 1552143600, 1552147200, 1552150800, 1552154400, 1552158000, 
    1552161600, 1552165200, 1552168800, 1552172400, 1552176000, 1552179600, 
    1552183200, 1552186800, 1552190400, 1552194000, 1552197600, 1552201200, 
    1552204800, 1552208400, 1552212000, 1552215600, 1552219200, 1552222800, 
    1552226400, 1552230000, 1552233600, 1552237200, 1552240800, 1552244400, 
    1552248000, 1552251600, 1552255200, 1552258800, 1552262400, 1552266000, 
    1552269600, 1552273200, 1552276800, 1552280400, 1552284000, 1552287600, 
    1552291200, 1552294800, 1552298400, 1552302000, 1552305600, 1552309200, 
    1552312800, 1552316400, 1552320000, 1552323600, 1552327200, 1552330800, 
    1552334400, 1552338000, 1552341600, 1552345200, 1552348800, 1552352400, 
    1552356000, 1552359600, 1552363200, 1552366800, 1552370400, 1552374000, 
    1552377600, 1552381200, 1552384800, 1552388400, 1552392000, 1552395600, 
    1552399200, 1552402800, 1552406400, 1552410000, 1552413600, 1552417200, 
    1552420800, 1552424400, 1552428000, 1552431600, 1552435200, 1552438800, 
    1552442400, 1552446000, 1552449600, 1552453200, 1552456800, 1552460400, 
    1552464000, 1552467600, 1552471200, 1552474800, 1552478400, 1552482000, 
    1552485600, 1552489200, 1552492800, 1552496400, 1552500000, 1552503600, 
    1552507200, 1552510800, 1552514400, 1552518000, 1552521600, 1552525200, 
    1552528800, 1552532400, 1552536000, 1552539600, 1552543200, 1552546800, 
    1552550400, 1552554000, 1552557600, 1552561200, 1552564800, 1552568400, 
    1552572000, 1552575600, 1552579200, 1552582800, 1552586400, 1552590000, 
    1552593600, 1552597200, 1552600800, 1552604400, 1552608000, 1552611600, 
    1552615200, 1552618800, 1552622400, 1552626000, 1552629600, 1552633200, 
    1552636800, 1552640400, 1552644000, 1552647600, 1552651200, 1552654800, 
    1552658400, 1552662000, 1552665600, 1552669200, 1552672800, 1552676400, 
    1552680000, 1552683600, 1552687200, 1552690800, 1552694400, 1552698000, 
    1552701600, 1552705200, 1552708800, 1552712400, 1552716000, 1552719600, 
    1552723200, 1552726800, 1552730400, 1552734000, 1552737600, 1552741200, 
    1552744800, 1552748400, 1552752000, 1552755600, 1552759200, 1552762800, 
    1552766400, 1552770000, 1552773600, 1552777200, 1552780800, 1552784400, 
    1552788000, 1552791600, 1552795200, 1552798800, 1552802400, 1552806000, 
    1552809600, 1552813200, 1552816800, 1552820400, 1552824000, 1552827600, 
    1552831200, 1552834800, 1552838400, 1552842000, 1552845600, 1552849200, 
    1552852800, 1552856400, 1552860000, 1552863600, 1552867200, 1552870800, 
    1552874400, 1552878000, 1552881600, 1552885200, 1552888800, 1552892400, 
    1552896000, 1552899600, 1552903200, 1552906800, 1552910400, 1552914000, 
    1552917600, 1552921200, 1552924800, 1552928400, 1552932000, 1552935600, 
    1552939200, 1552942800, 1552946400, 1552950000, 1552953600, 1552957200, 
    1552960800, 1552964400, 1552968000, 1552971600, 1552975200, 1552978800, 
    1552982400, 1552986000, 1552989600, 1552993200, 1552996800, 1553000400, 
    1553004000, 1553007600, 1553011200, 1553014800, 1553018400, 1553022000, 
    1553025600, 1553029200, 1553032800, 1553036400, 1553040000, 1553043600, 
    1553047200, 1553050800, 1553054400, 1553058000, 1553061600, 1553065200, 
    1553068800, 1553072400, 1553076000, 1553079600, 1553083200, 1553086800, 
    1553090400, 1553094000, 1553097600, 1553101200, 1553104800, 1553108400, 
    1553112000, 1553115600, 1553119200, 1553122800, 1553126400, 1553130000, 
    1553133600, 1553137200, 1553140800, 1553144400, 1553148000, 1553151600, 
    1553155200, 1553158800, 1553162400, 1553166000, 1553169600, 1553173200, 
    1553176800, 1553180400, 1553184000, 1553187600, 1553191200, 1553194800, 
    1553198400, 1553202000, 1553205600, 1553209200, 1553212800, 1553216400, 
    1553220000, 1553223600, 1553227200, 1553230800, 1553234400, 1553238000, 
    1553241600, 1553245200, 1553248800, 1553252400, 1553256000, 1553259600, 
    1553263200, 1553266800, 1553270400, 1553274000, 1553277600, 1553281200, 
    1553284800, 1553288400, 1553292000, 1553295600, 1553299200, 1553302800, 
    1553306400, 1553310000, 1553313600, 1553317200, 1553320800, 1553324400, 
    1553328000, 1553331600, 1553335200, 1553338800, 1553342400, 1553346000, 
    1553349600, 1553353200, 1553356800, 1553360400, 1553364000, 1553367600, 
    1553371200, 1553374800, 1553378400, 1553382000, 1553385600, 1553389200, 
    1553392800, 1553396400, 1553400000, 1553403600, 1553407200, 1553410800, 
    1553414400, 1553418000, 1553421600, 1553425200, 1553428800, 1553432400, 
    1553436000, 1553439600, 1553443200, 1553446800, 1553450400, 1553454000, 
    1553457600, 1553461200, 1553464800, 1553468400, 1553472000, 1553475600, 
    1553479200, 1553482800, 1553486400, 1553490000, 1553493600, 1553497200, 
    1553500800, 1553504400, 1553508000, 1553511600, 1553515200, 1553518800, 
    1553522400, 1553526000, 1553529600, 1553533200, 1553536800, 1553540400, 
    1553544000, 1553547600, 1553551200, 1553554800, 1553558400, 1553562000, 
    1553565600, 1553569200, 1553572800, 1553576400, 1553580000, 1553583600, 
    1553587200, 1553590800, 1553594400, 1553598000, 1553601600, 1553605200, 
    1553608800, 1553612400, 1553616000, 1553619600, 1553623200, 1553626800, 
    1553630400, 1553634000, 1553637600, 1553641200, 1553644800, 1553648400, 
    1553652000, 1553655600, 1553659200, 1553662800, 1553666400, 1553670000, 
    1553673600, 1553677200, 1553680800, 1553684400, 1553688000, 1553691600, 
    1553695200, 1553698800, 1553702400, 1553706000, 1553709600, 1553713200, 
    1553716800, 1553720400, 1553724000, 1553727600, 1553731200, 1553734800, 
    1553738400, 1553742000, 1553745600, 1553749200, 1553752800, 1553756400, 
    1553760000, 1553763600, 1553767200, 1553770800, 1553774400, 1553778000, 
    1553781600, 1553785200, 1553788800, 1553792400, 1553796000, 1553799600, 
    1553803200, 1553806800, 1553810400, 1553814000, 1553817600, 1553821200, 
    1553824800, 1553828400, 1553832000, 1553835600, 1553839200, 1553842800, 
    1553846400, 1553850000, 1553853600, 1553857200, 1553860800, 1553864400, 
    1553868000, 1553871600, 1553875200, 1553878800, 1553882400, 1553886000, 
    1553889600, 1553893200, 1553896800, 1553900400, 1553904000, 1553907600, 
    1553911200, 1553914800, 1553918400, 1553922000, 1553925600, 1553929200, 
    1553932800, 1553936400, 1553940000, 1553943600, 1553947200, 1553950800, 
    1553954400, 1553958000, 1553961600, 1553965200, 1553968800, 1553972400, 
    1553976000, 1553979600, 1553983200, 1553986800, 1553990400, 1553994000, 
    1553997600, 1554001200, 1554004800, 1554008400, 1554012000, 1554015600, 
    1554019200, 1554022800, 1554026400, 1554030000, 1554033600, 1554037200, 
    1554040800, 1554044400, 1554048000, 1554051600, 1554055200, 1554058800, 
    1554062400, 1554066000, 1554069600, 1554073200, 1554076800, 1554080400, 
    1554084000, 1554087600, 1554091200, 1554094800, 1554098400, 1554102000, 
    1554105600, 1554109200, 1554112800, 1554116400, 1554120000, 1554123600, 
    1554127200, 1554130800, 1554134400, 1554138000, 1554141600, 1554145200, 
    1554148800, 1554152400, 1554156000, 1554159600, 1554163200, 1554166800, 
    1554170400, 1554174000, 1554177600, 1554181200, 1554184800, 1554188400, 
    1554192000, 1554195600, 1554199200, 1554202800, 1554206400, 1554210000, 
    1554213600, 1554217200, 1554220800, 1554224400, 1554228000, 1554231600, 
    1554235200, 1554238800, 1554242400, 1554246000, 1554249600, 1554253200, 
    1554256800, 1554260400, 1554264000, 1554267600, 1554271200, 1554274800, 
    1554278400, 1554282000, 1554285600, 1554289200, 1554292800, 1554296400, 
    1554300000, 1554303600, 1554307200, 1554310800, 1554314400, 1554318000, 
    1554321600, 1554325200, 1554328800, 1554332400, 1554336000, 1554339600, 
    1554343200, 1554346800, 1554350400, 1554354000, 1554357600, 1554361200, 
    1554364800, 1554368400, 1554372000, 1554375600, 1554379200, 1554382800, 
    1554386400, 1554390000, 1554393600, 1554397200, 1554400800, 1554404400, 
    1554408000, 1554411600, 1554415200, 1554418800, 1554422400, 1554426000, 
    1554429600, 1554433200, 1554436800, 1554440400, 1554444000, 1554447600, 
    1554451200, 1554454800, 1554458400, 1554462000, 1554465600, 1554469200, 
    1554472800, 1554476400, 1554480000, 1554483600, 1554487200, 1554490800, 
    1554494400, 1554498000, 1554501600, 1554505200, 1554508800, 1554512400, 
    1554516000, 1554519600, 1554523200, 1554526800, 1554530400, 1554534000, 
    1554537600, 1554541200, 1554544800, 1554548400, 1554552000, 1554555600, 
    1554559200, 1554562800, 1554566400, 1554570000, 1554573600, 1554577200, 
    1554580800, 1554584400, 1554588000, 1554591600, 1554595200, 1554598800, 
    1554602400, 1554606000, 1554609600, 1554613200, 1554616800, 1554620400, 
    1554624000, 1554627600, 1554631200, 1554634800, 1554638400, 1554642000, 
    1554645600, 1554649200, 1554652800, 1554656400, 1554660000, 1554663600, 
    1554667200, 1554670800, 1554674400, 1554678000, 1554681600, 1554685200, 
    1554688800, 1554692400, 1554696000, 1554699600, 1554703200, 1554706800, 
    1554710400, 1554714000, 1554717600, 1554721200, 1554724800, 1554728400, 
    1554732000, 1554735600, 1554739200, 1554742800, 1554746400, 1554750000, 
    1554753600, 1554757200, 1554760800, 1554764400, 1554768000, 1554771600, 
    1554775200, 1554778800, 1554782400, 1554786000, 1554789600, 1554793200, 
    1554796800, 1554800400, 1554804000, 1554807600, 1554811200, 1554814800, 
    1554818400, 1554822000, 1554825600, 1554829200, 1554832800, 1554836400, 
    1554840000, 1554843600, 1554847200, 1554850800, 1554854400, 1554858000, 
    1554861600, 1554865200, 1554868800, 1554872400, 1554876000, 1554879600, 
    1554883200, 1554886800, 1554890400, 1554894000, 1554897600, 1554901200, 
    1554904800, 1554908400, 1554912000, 1554915600, 1554919200, 1554922800, 
    1554926400, 1554930000, 1554933600, 1554937200, 1554940800, 1554944400, 
    1554948000, 1554951600, 1554955200, 1554958800, 1554962400, 1554966000, 
    1554969600, 1554973200, 1554976800, 1554980400, 1554984000, 1554987600, 
    1554991200, 1554994800, 1554998400, 1555002000, 1555005600, 1555009200, 
    1555012800, 1555016400, 1555020000, 1555023600, 1555027200, 1555030800, 
    1555034400, 1555038000, 1555041600, 1555045200, 1555048800, 1555052400, 
    1555056000, 1555059600, 1555063200, 1555066800, 1555070400, 1555074000, 
    1555077600, 1555081200, 1555084800, 1555088400, 1555092000, 1555095600, 
    1555099200, 1555102800, 1555106400, 1555110000, 1555113600, 1555117200, 
    1555120800, 1555124400, 1555128000, 1555131600, 1555135200, 1555138800, 
    1555142400, 1555146000, 1555149600, 1555153200, 1555156800, 1555160400, 
    1555164000, 1555167600, 1555171200, 1555174800, 1555178400, 1555182000, 
    1555185600, 1555189200, 1555192800, 1555196400, 1555200000, 1555203600, 
    1555207200, 1555210800, 1555214400, 1555218000, 1555221600, 1555225200, 
    1555228800, 1555232400, 1555236000, 1555239600, 1555243200, 1555246800, 
    1555250400, 1555254000, 1555257600, 1555261200, 1555264800, 1555268400, 
    1555272000, 1555275600, 1555279200, 1555282800, 1555286400, 1555290000, 
    1555293600, 1555297200, 1555300800, 1555304400, 1555308000, 1555311600, 
    1555315200, 1555318800, 1555322400, 1555326000, 1555329600, 1555333200, 
    1555336800, 1555340400, 1555344000, 1555347600, 1555351200, 1555354800, 
    1555358400, 1555362000, 1555365600, 1555369200, 1555372800, 1555376400, 
    1555380000, 1555383600, 1555387200, 1555390800, 1555394400, 1555398000, 
    1555401600, 1555405200, 1555408800, 1555412400, 1555416000, 1555419600, 
    1555423200, 1555426800, 1555430400, 1555434000, 1555437600, 1555441200, 
    1555444800, 1555448400, 1555452000, 1555455600, 1555459200, 1555462800, 
    1555466400, 1555470000, 1555473600, 1555477200, 1555480800, 1555484400, 
    1555488000, 1555491600, 1555495200, 1555498800, 1555502400, 1555506000, 
    1555509600, 1555513200, 1555516800, 1555520400, 1555524000, 1555527600, 
    1555531200, 1555534800, 1555538400, 1555542000, 1555545600, 1555549200, 
    1555552800, 1555556400, 1555560000, 1555563600, 1555567200, 1555570800, 
    1555574400, 1555578000, 1555581600, 1555585200, 1555588800, 1555592400, 
    1555596000, 1555599600, 1555603200, 1555606800, 1555610400, 1555614000, 
    1555617600, 1555621200, 1555624800, 1555628400, 1555632000, 1555635600, 
    1555639200, 1555642800, 1555646400, 1555650000, 1555653600, 1555657200, 
    1555660800, 1555664400, 1555668000, 1555671600, 1555675200, 1555678800, 
    1555682400, 1555686000, 1555689600, 1555693200, 1555696800, 1555700400, 
    1555704000, 1555707600, 1555711200, 1555714800, 1555718400, 1555722000, 
    1555725600, 1555729200, 1555732800, 1555736400, 1555740000, 1555743600, 
    1555747200, 1555750800, 1555754400, 1555758000, 1555761600, 1555765200, 
    1555768800, 1555772400, 1555776000, 1555779600, 1555783200, 1555786800, 
    1555790400, 1555794000, 1555797600, 1555801200, 1555804800, 1555808400, 
    1555812000, 1555815600, 1555819200, 1555822800, 1555826400, 1555830000, 
    1555833600, 1555837200, 1555840800, 1555844400, 1555848000, 1555851600, 
    1555855200, 1555858800, 1555862400, 1555866000, 1555869600, 1555873200, 
    1555876800, 1555880400, 1555884000, 1555887600, 1555891200, 1555894800, 
    1555898400, 1555902000, 1555905600, 1555909200, 1555912800, 1555916400, 
    1555920000, 1555923600, 1555927200, 1555930800, 1555934400, 1555938000, 
    1555941600, 1555945200, 1555948800, 1555952400, 1555956000, 1555959600, 
    1555963200, 1555966800, 1555970400, 1555974000, 1555977600, 1555981200, 
    1555984800, 1555988400, 1555992000, 1555995600, 1555999200, 1556002800, 
    1556006400, 1556010000, 1556013600, 1556017200, 1556020800, 1556024400, 
    1556028000, 1556031600, 1556035200, 1556038800, 1556042400, 1556046000, 
    1556049600, 1556053200, 1556056800, 1556060400, 1556064000, 1556067600, 
    1556071200, 1556074800, 1556078400, 1556082000, 1556085600, 1556089200, 
    1556092800, 1556096400, 1556100000, 1556103600, 1556107200, 1556110800, 
    1556114400, 1556118000, 1556121600, 1556125200, 1556128800, 1556132400, 
    1556136000, 1556139600, 1556143200, 1556146800, 1556150400, 1556154000, 
    1556157600, 1556161200, 1556164800, 1556168400, 1556172000, 1556175600, 
    1556179200, 1556182800, 1556186400, 1556190000, 1556193600, 1556197200, 
    1556200800, 1556204400, 1556208000, 1556211600, 1556215200, 1556218800, 
    1556222400, 1556226000, 1556229600, 1556233200, 1556236800, 1556240400, 
    1556244000, 1556247600, 1556251200, 1556254800, 1556258400, 1556262000, 
    1556265600, 1556269200, 1556272800, 1556276400, 1556280000, 1556283600, 
    1556287200, 1556290800, 1556294400, 1556298000, 1556301600, 1556305200, 
    1556308800, 1556312400, 1556316000, 1556319600, 1556323200, 1556326800, 
    1556330400, 1556334000, 1556337600, 1556341200, 1556344800, 1556348400, 
    1556352000, 1556355600, 1556359200, 1556362800, 1556366400, 1556370000, 
    1556373600, 1556377200, 1556380800, 1556384400, 1556388000, 1556391600, 
    1556395200, 1556398800, 1556402400, 1556406000, 1556409600, 1556413200, 
    1556416800, 1556420400, 1556424000, 1556427600, 1556431200, 1556434800, 
    1556438400, 1556442000, 1556445600, 1556449200, 1556452800, 1556456400, 
    1556460000, 1556463600, 1556467200, 1556470800, 1556474400, 1556478000, 
    1556481600, 1556485200, 1556488800, 1556492400, 1556496000, 1556499600, 
    1556503200, 1556506800, 1556510400, 1556514000, 1556517600, 1556521200, 
    1556524800, 1556528400, 1556532000, 1556535600, 1556539200, 1556542800, 
    1556546400, 1556550000, 1556553600, 1556557200, 1556560800, 1556564400, 
    1556568000, 1556571600, 1556575200, 1556578800, 1556582400, 1556586000, 
    1556589600, 1556593200, 1556596800, 1556600400, 1556604000, 1556607600, 
    1556611200, 1556614800, 1556618400, 1556622000, 1556625600, 1556629200, 
    1556632800, 1556636400, 1556640000, 1556643600, 1556647200, 1556650800, 
    1556654400, 1556658000, 1556661600, 1556665200, 1556668800, 1556672400, 
    1556676000, 1556679600, 1556683200, 1556686800, 1556690400, 1556694000, 
    1556697600, 1556701200, 1556704800, 1556708400, 1556712000, 1556715600, 
    1556719200, 1556722800, 1556726400, 1556730000, 1556733600, 1556737200, 
    1556740800, 1556744400, 1556748000, 1556751600, 1556755200, 1556758800, 
    1556762400, 1556766000, 1556769600, 1556773200, 1556776800, 1556780400, 
    1556784000, 1556787600, 1556791200, 1556794800, 1556798400, 1556802000, 
    1556805600, 1556809200, 1556812800, 1556816400, 1556820000, 1556823600, 
    1556827200, 1556830800, 1556834400, 1556838000, 1556841600, 1556845200, 
    1556848800, 1556852400, 1556856000, 1556859600, 1556863200, 1556866800, 
    1556870400, 1556874000, 1556877600, 1556881200, 1556884800, 1556888400, 
    1556892000, 1556895600, 1556899200, 1556902800, 1556906400, 1556910000, 
    1556913600, 1556917200, 1556920800, 1556924400, 1556928000, 1556931600, 
    1556935200, 1556938800, 1556942400, 1556946000, 1556949600, 1556953200, 
    1556956800, 1556960400, 1556964000, 1556967600, 1556971200, 1556974800, 
    1556978400, 1556982000, 1556985600, 1556989200, 1556992800, 1556996400, 
    1557000000, 1557003600, 1557007200, 1557010800, 1557014400, 1557018000, 
    1557021600, 1557025200, 1557028800, 1557032400, 1557036000, 1557039600, 
    1557043200, 1557046800, 1557050400, 1557054000, 1557057600, 1557061200, 
    1557064800, 1557068400, 1557072000, 1557075600, 1557079200, 1557082800, 
    1557086400, 1557090000, 1557093600, 1557097200, 1557100800, 1557104400, 
    1557108000, 1557111600, 1557115200, 1557118800, 1557122400, 1557126000, 
    1557129600, 1557133200, 1557136800, 1557140400, 1557144000, 1557147600, 
    1557151200, 1557154800, 1557158400, 1557162000, 1557165600, 1557169200, 
    1557172800, 1557176400, 1557180000, 1557183600, 1557187200, 1557190800, 
    1557194400, 1557198000, 1557201600, 1557205200, 1557208800, 1557212400, 
    1557216000, 1557219600, 1557223200, 1557226800, 1557230400, 1557234000, 
    1557237600, 1557241200, 1557244800, 1557248400, 1557252000, 1557255600, 
    1557259200, 1557262800, 1557266400, 1557270000, 1557273600, 1557277200, 
    1557280800, 1557284400, 1557288000, 1557291600, 1557295200, 1557298800, 
    1557302400, 1557306000, 1557309600, 1557313200, 1557316800, 1557320400, 
    1557324000, 1557327600, 1557331200, 1557334800, 1557338400, 1557342000, 
    1557345600, 1557349200, 1557352800, 1557356400, 1557360000, 1557363600, 
    1557367200, 1557370800, 1557374400, 1557378000, 1557381600, 1557385200, 
    1557388800, 1557392400, 1557396000, 1557399600, 1557403200, 1557406800, 
    1557410400, 1557414000, 1557417600, 1557421200, 1557424800, 1557428400, 
    1557432000, 1557435600, 1557439200, 1557442800, 1557446400, 1557450000, 
    1557453600, 1557457200, 1557460800, 1557464400, 1557468000, 1557471600, 
    1557475200, 1557478800, 1557482400, 1557486000, 1557489600, 1557493200, 
    1557496800, 1557500400, 1557504000, 1557507600, 1557511200, 1557514800, 
    1557518400, 1557522000, 1557525600, 1557529200, 1557532800, 1557536400, 
    1557540000, 1557543600, 1557547200, 1557550800, 1557554400, 1557558000, 
    1557561600, 1557565200, 1557568800, 1557572400, 1557576000, 1557579600, 
    1557583200, 1557586800, 1557590400, 1557594000, 1557597600, 1557601200, 
    1557604800, 1557608400, 1557612000, 1557615600, 1557619200, 1557622800, 
    1557626400, 1557630000, 1557633600, 1557637200, 1557640800, 1557644400, 
    1557648000, 1557651600, 1557655200, 1557658800, 1557662400, 1557666000, 
    1557669600, 1557673200, 1557676800, 1557680400, 1557684000, 1557687600, 
    1557691200, 1557694800, 1557698400, 1557702000, 1557705600, 1557709200, 
    1557712800, 1557716400, 1557720000, 1557723600, 1557727200, 1557730800, 
    1557734400, 1557738000, 1557741600, 1557745200, 1557748800, 1557752400, 
    1557756000, 1557759600, 1557763200, 1557766800, 1557770400, 1557774000, 
    1557777600, 1557781200, 1557784800, 1557788400, 1557792000, 1557795600, 
    1557799200, 1557802800, 1557806400, 1557810000, 1557813600, 1557817200, 
    1557820800, 1557824400, 1557828000, 1557831600, 1557835200, 1557838800, 
    1557842400, 1557846000, 1557849600, 1557853200, 1557856800, 1557860400, 
    1557864000, 1557867600, 1557871200, 1557874800, 1557878400, 1557882000, 
    1557885600, 1557889200, 1557892800, 1557896400, 1557900000, 1557903600, 
    1557907200, 1557910800, 1557914400, 1557918000, 1557921600, 1557925200, 
    1557928800, 1557932400, 1557936000, 1557939600, 1557943200, 1557946800, 
    1557950400, 1557954000, 1557957600, 1557961200, 1557964800, 1557968400, 
    1557972000, 1557975600, 1557979200, 1557982800, 1557986400, 1557990000, 
    1557993600, 1557997200, 1558000800, 1558004400, 1558008000, 1558011600, 
    1558015200, 1558018800, 1558022400, 1558026000, 1558029600, 1558033200, 
    1558036800, 1558040400, 1558044000, 1558047600, 1558051200, 1558054800, 
    1558058400, 1558062000, 1558065600, 1558069200, 1558072800, 1558076400, 
    1558080000, 1558083600, 1558087200, 1558090800, 1558094400, 1558098000, 
    1558101600, 1558105200, 1558108800, 1558112400, 1558116000, 1558119600, 
    1558123200, 1558126800, 1558130400, 1558134000, 1558137600, 1558141200, 
    1558144800, 1558148400, 1558152000, 1558155600, 1558159200, 1558162800, 
    1558166400, 1558170000, 1558173600, 1558177200, 1558180800, 1558184400, 
    1558188000, 1558191600, 1558195200, 1558198800, 1558202400, 1558206000, 
    1558209600, 1558213200, 1558216800, 1558220400, 1558224000, 1558227600, 
    1558231200, 1558234800, 1558238400, 1558242000, 1558245600, 1558249200, 
    1558252800, 1558256400, 1558260000, 1558263600, 1558267200, 1558270800, 
    1558274400, 1558278000, 1558281600, 1558285200, 1558288800, 1558292400, 
    1558296000, 1558299600, 1558303200, 1558306800, 1558310400, 1558314000, 
    1558317600, 1558321200, 1558324800, 1558328400, 1558332000, 1558335600, 
    1558339200, 1558342800, 1558346400, 1558350000, 1558353600, 1558357200, 
    1558360800, 1558364400, 1558368000, 1558371600, 1558375200, 1558378800, 
    1558382400, 1558386000, 1558389600, 1558393200, 1558396800, 1558400400, 
    1558404000, 1558407600, 1558411200, 1558414800, 1558418400, 1558422000, 
    1558425600, 1558429200, 1558432800, 1558436400, 1558440000, 1558443600, 
    1558447200, 1558450800, 1558454400, 1558458000, 1558461600, 1558465200, 
    1558468800, 1558472400, 1558476000, 1558479600, 1558483200, 1558486800, 
    1558490400, 1558494000, 1558497600, 1558501200, 1558504800, 1558508400, 
    1558512000, 1558515600, 1558519200, 1558522800, 1558526400, 1558530000, 
    1558533600, 1558537200, 1558540800, 1558544400, 1558548000, 1558551600, 
    1558555200, 1558558800, 1558562400, 1558566000, 1558569600, 1558573200, 
    1558576800, 1558580400, 1558584000, 1558587600, 1558591200, 1558594800, 
    1558598400, 1558602000, 1558605600, 1558609200, 1558612800, 1558616400, 
    1558620000, 1558623600, 1558627200, 1558630800, 1558634400, 1558638000, 
    1558641600, 1558645200, 1558648800, 1558652400, 1558656000, 1558659600, 
    1558663200, 1558666800, 1558670400, 1558674000, 1558677600, 1558681200, 
    1558684800, 1558688400, 1558692000, 1558695600, 1558699200, 1558702800, 
    1558706400, 1558710000, 1558713600, 1558717200, 1558720800, 1558724400, 
    1558728000, 1558731600, 1558735200, 1558738800, 1558742400, 1558746000, 
    1558749600, 1558753200, 1558756800, 1558760400, 1558764000, 1558767600, 
    1558771200, 1558774800, 1558778400, 1558782000, 1558785600, 1558789200, 
    1558792800, 1558796400, 1558800000, 1558803600, 1558807200, 1558810800, 
    1558814400, 1558818000, 1558821600, 1558825200, 1558828800, 1558832400, 
    1558836000, 1558839600, 1558843200, 1558846800, 1558850400, 1558854000, 
    1558857600, 1558861200, 1558864800, 1558868400, 1558872000, 1558875600, 
    1558879200, 1558882800, 1558886400, 1558890000, 1558893600, 1558897200, 
    1558900800, 1558904400, 1558908000, 1558911600, 1558915200, 1558918800, 
    1558922400, 1558926000, 1558929600, 1558933200, 1558936800, 1558940400, 
    1558944000, 1558947600, 1558951200, 1558954800, 1558958400, 1558962000, 
    1558965600, 1558969200, 1558972800, 1558976400, 1558980000, 1558983600, 
    1558987200, 1558990800, 1558994400, 1558998000, 1559001600, 1559005200, 
    1559008800, 1559012400, 1559016000, 1559019600, 1559023200, 1559026800, 
    1559030400, 1559034000, 1559037600, 1559041200, 1559044800, 1559048400, 
    1559052000, 1559055600, 1559059200, 1559062800, 1559066400, 1559070000, 
    1559073600, 1559077200, 1559080800, 1559084400, 1559088000, 1559091600, 
    1559095200, 1559098800, 1559102400, 1559106000, 1559109600, 1559113200, 
    1559116800, 1559120400, 1559124000, 1559127600, 1559131200, 1559134800, 
    1559138400, 1559142000, 1559145600, 1559149200, 1559152800, 1559156400, 
    1559160000, 1559163600, 1559167200, 1559170800, 1559174400, 1559178000, 
    1559181600, 1559185200, 1559188800, 1559192400, 1559196000, 1559199600, 
    1559203200, 1559206800, 1559210400, 1559214000, 1559217600, 1559221200, 
    1559224800, 1559228400, 1559232000, 1559235600, 1559239200, 1559246400, 
    1559250000, 1559253600, 1559257200, 1559260800, 1559264400, 1559268000, 
    1559271600, 1559275200, 1559278800, 1559242800, 1559282400, 1559286000, 
    1559289600, 1559293200, 1559296800, 1559300400, 1559304000, 1559307600, 
    1559311200, 1559314800, 1559318400, 1559322000, 1559325600, 1559329200, 
    1559332800, 1559336400, 1559340000, 1559343600, 1559347200, 1559350800, 
    1559354400, 1559358000, 1559361600, 1559365200, 1559368800, 1559372400, 
    1559376000, 1559379600, 1559383200, 1559386800, 1559390400, 1559394000, 
    1559397600, 1559401200, 1559404800, 1559408400, 1559412000, 1559415600, 
    1559419200, 1559422800, 1559426400, 1559430000, 1559433600, 1559437200, 
    1559440800, 1559444400, 1559448000, 1559451600, 1559455200, 1559458800, 
    1559462400, 1559466000, 1559469600, 1559473200, 1559476800, 1559480400, 
    1559484000, 1559487600, 1559491200, 1559494800, 1559498400, 1559502000, 
    1559505600, 1559509200, 1559512800, 1559516400, 1559520000, 1559523600, 
    1559527200, 1559530800, 1559534400, 1559538000, 1559545200, 1559541600, 
    1559548800, 1559552400, 1559556000, 1559559600, 1559563200, 1559566800, 
    1559570400, 1559574000, 1559577600, 1559581200, 1559584800, 1559588400, 
    1559592000, 1559595600, 1559599200, 1559602800, 1559606400, 1559610000, 
    1559613600, 1559617200, 1559620800, 1559624400, 1559628000, 1559631600, 
    1559635200, 1559638800, 1559642400, 1559646000, 1559649600, 1559653200, 
    1559656800, 1559660400, 1559664000, 1559667600, 1559671200, 1559674800, 
    1559678400, 1559682000, 1559685600, 1559689200, 1559692800, 1559696400, 
    1559700000, 1559703600, 1559707200, 1559710800, 1559714400, 1559718000, 
    1559721600, 1559725200, 1559728800, 1559732400, 1559736000, 1559743200, 
    1559746800, 1559750400, 1559754000, 1559757600, 1559761200, 1559764800, 
    1559768400, 1559772000, 1559775600, 1559779200, 1559782800, 1559739600, 
    1559786400, 1559790000, 1559793600, 1559797200, 1559800800, 1559804400, 
    1559808000, 1559811600, 1559815200, 1559818800, 1559822400, 1559826000, 
    1559829600, 1559833200, 1559836800, 1559840400, 1559844000, 1559847600, 
    1559851200, 1559854800, 1559858400, 1559862000, 1559865600, 1559869200, 
    1559872800, 1559876400, 1559880000, 1559883600, 1559887200, 1559890800, 
    1559894400, 1559898000, 1559901600, 1559905200, 1559908800, 1559912400, 
    1559916000, 1559919600, 1559923200, 1559926800, 1559930400, 1559934000, 
    1559937600, 1559941200, 1559944800, 1559948400, 1559952000, 1559955600, 
    1559959200, 1559962800, 1559966400, 1559970000, 1559973600, 1559977200, 
    1559980800, 1559984400, 1559988000, 1559991600, 1559995200, 1559998800, 
    1560002400, 1560006000, 1560009600, 1560013200, 1560016800, 1560020400, 
    1560024000, 1560027600, 1560031200, 1560034800, 1560038400, 1560042000, 
    1560045600, 1560049200, 1560052800, 1560056400, 1560060000, 1560063600, 
    1560067200, 1560070800, 1560074400, 1560078000, 1560081600, 1560085200, 
    1560088800, 1560092400, 1560096000, 1560099600, 1560103200, 1560106800, 
    1560110400, 1560114000, 1560117600, 1560121200, 1560124800, 1560128400, 
    1560132000, 1560135600, 1560139200, 1560142800, 1560146400, 1560150000, 
    1560153600, 1560157200, 1560160800, 1560164400, 1560168000, 1560171600, 
    1560175200, 1560178800, 1560182400, 1560186000, 1560189600, 1560193200, 
    1560196800, 1560200400, 1560204000, 1560207600, 1560211200, 1560214800, 
    1560218400, 1560222000, 1560225600, 1560229200, 1560232800, 1560236400, 
    1560240000, 1560243600, 1560247200, 1560250800, 1560254400, 1560258000, 
    1560261600, 1560265200, 1560268800, 1560272400, 1560276000, 1560279600, 
    1560283200, 1560286800, 1560290400, 1560294000, 1560297600, 1560301200, 
    1560304800, 1560308400, 1560312000, 1560315600, 1560319200, 1560322800, 
    1560326400, 1560330000, 1560333600, 1560337200, 1560340800, 1560344400, 
    1560348000, 1560351600, 1560355200, 1560358800, 1560362400, 1560366000, 
    1560369600, 1560373200, 1560376800, 1560380400, 1560384000, 1560387600, 
    1560391200, 1560394800, 1560398400, 1560402000, 1560405600, 1560409200, 
    1560412800, 1560416400, 1560420000, 1560423600, 1560427200, 1560430800, 
    1560434400, 1560438000, 1560441600, 1560445200, 1560448800, 1560452400, 
    1560456000, 1560459600, 1560463200, 1560466800, 1560470400, 1560474000, 
    1560477600, 1560481200, 1560484800, 1560488400, 1560492000, 1560495600, 
    1560499200, 1560502800, 1560506400, 1560510000, 1560513600, 1560517200, 
    1560520800, 1560524400, 1560528000, 1560531600, 1560535200, 1560538800, 
    1560542400, 1560546000, 1560549600, 1560553200, 1560556800, 1560560400, 
    1560564000, 1560567600, 1560571200, 1560574800, 1560582000, 1560585600, 
    1560589200, 1560592800, 1560596400, 1560600000, 1560603600, 1560607200, 
    1560610800, 1560614400, 1560618000, 1560621600, 1560625200, 1560628800, 
    1560632400, 1560636000, 1560639600, 1560643200, 1560646800, 1560650400, 
    1560654000, 1560657600, 1560661200, 1560664800, 1560578400, 1560668400, 
    1560672000, 1560675600, 1560679200, 1560682800, 1560686400, 1560690000, 
    1560693600, 1560697200, 1560700800, 1560704400, 1560708000, 1560711600, 
    1560715200, 1560718800, 1560722400, 1560726000, 1560729600, 1560733200, 
    1560736800, 1560740400, 1560744000, 1560747600, 1560751200, 1560754800, 
    1560758400, 1560762000, 1560765600, 1560769200, 1560772800, 1560776400, 
    1560780000, 1560783600, 1560787200, 1560790800, 1560794400, 1560798000, 
    1560801600, 1560805200, 1560808800, 1560812400, 1560816000, 1560819600, 
    1560823200, 1560826800, 1560830400, 1560834000, 1560837600, 1560841200, 
    1560844800, 1560848400, 1560852000, 1560855600, 1560859200, 1560862800, 
    1560866400, 1560870000, 1560873600, 1560877200, 1560880800, 1560884400, 
    1560888000, 1560891600, 1560895200, 1560898800, 1560902400, 1560906000, 
    1560909600, 1560913200, 1560916800, 1560920400, 1560924000, 1560927600, 
    1560931200, 1560934800, 1560938400, 1560942000, 1560945600, 1560949200, 
    1560952800, 1560956400, 1560960000, 1560963600, 1560967200, 1560970800, 
    1560974400, 1560978000, 1560981600, 1560985200, 1560988800, 1560992400, 
    1560996000, 1560999600, 1561003200, 1561006800, 1561010400, 1561014000, 
    1561017600, 1561021200, 1561024800, 1561028400, 1561032000, 1561035600, 
    1561039200, 1561042800, 1561046400, 1561050000, 1561053600, 1561057200, 
    1561060800, 1561064400, 1561068000, 1561071600, 1561075200, 1561078800, 
    1561082400, 1561086000, 1561089600, 1561093200, 1561096800, 1561100400, 
    1561104000, 1561107600, 1561111200, 1561114800, 1561118400, 1561122000, 
    1561125600, 1561129200, 1561132800, 1561136400, 1561140000, 1561143600, 
    1561147200, 1561150800, 1561154400, 1561158000, 1561161600, 1561165200, 
    1561168800, 1561172400, 1561176000, 1561179600, 1561183200, 1561186800, 
    1561190400, 1561194000, 1561197600, 1561201200, 1561204800, 1561208400, 
    1561212000, 1561215600, 1561219200, 1561222800, 1561226400, 1561230000, 
    1561233600, 1561237200, 1561240800, 1561244400, 1561248000, 1561251600, 
    1561255200, 1561258800, 1561262400, 1561266000, 1561269600, 1561273200, 
    1561276800, 1561280400, 1561284000, 1561287600, 1561291200, 1561294800, 
    1561298400, 1561302000, 1561305600, 1561309200, 1561312800, 1561316400, 
    1561320000, 1561323600, 1561327200, 1561330800, 1561334400, 1561338000, 
    1561341600, 1561345200, 1561348800, 1561352400, 1561356000, 1561359600, 
    1561363200, 1561366800, 1561370400, 1561374000, 1561377600, 1561381200, 
    1561384800, 1561388400, 1561392000, 1561395600, 1561399200, 1561402800, 
    1561406400, 1561410000, 1561413600, 1561417200, 1561420800, 1561424400, 
    1561428000, 1561431600, 1561435200, 1561438800, 1561442400, 1561446000, 
    1561449600, 1561453200, 1561456800, 1561460400, 1561464000, 1561467600, 
    1561471200, 1561474800, 1561478400, 1561482000, 1561485600, 1561489200, 
    1561492800, 1561496400, 1561500000, 1561503600, 1561507200, 1561510800, 
    1561514400, 1561518000, 1561521600, 1561525200, 1561528800, 1561532400, 
    1561536000, 1561539600, 1561543200, 1561546800, 1561550400, 1561554000, 
    1561557600, 1561561200, 1561564800, 1561568400, 1561572000, 1561575600, 
    1561579200, 1561582800, 1561586400, 1561590000, 1561593600, 1561597200, 
    1561600800, 1561604400, 1561608000, 1561611600, 1561615200, 1561618800, 
    1561622400, 1561626000, 1561629600, 1561633200, 1561636800, 1561640400, 
    1561644000, 1561647600, 1561651200, 1561654800, 1561658400, 1561662000, 
    1561665600, 1561669200, 1561672800, 1561676400, 1561680000, 1561683600, 
    1561687200, 1561690800, 1561694400, 1561698000, 1561701600, 1561705200, 
    1561708800, 1561712400, 1561716000, 1561719600, 1561723200, 1561726800, 
    1561730400, 1561734000, 1561737600, 1561741200, 1561744800, 1561748400, 
    1561752000, 1561755600, 1561759200, 1561762800, 1561766400, 1561770000, 
    1561773600, 1561777200, 1561780800, 1561784400, 1561788000, 1561791600, 
    1561795200, 1561798800, 1561802400, 1561806000, 1561809600, 1561813200, 
    1561816800, 1561820400, 1561824000, 1561827600, 1561831200, 1561834800, 
    1561838400, 1561842000, 1561845600, 1561849200, 1561852800, 1561856400, 
    1561860000, 1561863600, 1561867200, 1561870800, 1561874400, 1561878000, 
    1561881600, 1561885200, 1561888800, 1561892400, 1561896000, 1561899600, 
    1561903200, 1561906800, 1561910400, 1561914000, 1561917600, 1561921200, 
    1561924800, 1561928400, 1561932000, 1561935600, 1561939200, 1561942800, 
    1561946400, 1561950000, 1561953600, 1561957200, 1561960800, 1561964400, 
    1561968000, 1561971600, 1561975200, 1561978800, 1561982400, 1561986000, 
    1561989600, 1561993200, 1561996800, 1562000400, 1562004000, 1562007600, 
    1562011200, 1562014800, 1562018400, 1562022000, 1562025600, 1562029200, 
    1562032800, 1562036400, 1562040000, 1562043600, 1562047200, 1562050800, 
    1562054400, 1562058000, 1562061600, 1562065200, 1562068800, 1562072400, 
    1562076000, 1562079600, 1562083200, 1562086800, 1562090400, 1562094000, 
    1562097600, 1562101200, 1562104800, 1562108400, 1562112000, 1562115600, 
    1562119200, 1562122800, 1562126400, 1562130000, 1562133600, 1562137200, 
    1562140800, 1562144400, 1562148000, 1562151600, 1562155200, 1562158800, 
    1562162400, 1562166000, 1562169600, 1562173200, 1562176800, 1562180400, 
    1562184000, 1562187600, 1562191200, 1562194800, 1562198400, 1562202000, 
    1562205600, 1562209200, 1562212800, 1562216400, 1562220000, 1562223600, 
    1562227200, 1562230800, 1562234400, 1562238000, 1562241600, 1562245200, 
    1562248800, 1562252400, 1562256000, 1562259600, 1562263200, 1562266800, 
    1562270400, 1562274000, 1562277600, 1562281200, 1562284800, 1562288400, 
    1562292000, 1562295600, 1562299200, 1562302800, 1562306400, 1562310000, 
    1562313600, 1562317200, 1562320800, 1562324400, 1562328000, 1562331600, 
    1562335200, 1562338800, 1562342400, 1562346000, 1562349600, 1562353200, 
    1562356800, 1562360400, 1562364000, 1562367600, 1562371200, 1562374800, 
    1562378400, 1562382000, 1562385600, 1562389200, 1562392800, 1562396400, 
    1562400000, 1562403600, 1562407200, 1562410800, 1562414400, 1562418000, 
    1562421600, 1562425200, 1562428800, 1562432400, 1562436000, 1562439600, 
    1562443200, 1562446800, 1562450400, 1562454000, 1562457600, 1562461200, 
    1562464800, 1562468400, 1562472000, 1562475600, 1562479200, 1562482800, 
    1562486400, 1562490000, 1562493600, 1562497200, 1562500800, 1562504400, 
    1562508000, 1562511600, 1562515200, 1562518800, 1562522400, 1562526000, 
    1562529600, 1562533200, 1562536800, 1562540400, 1562544000, 1562547600, 
    1562554800, 1562558400, 1562562000, 1562565600, 1562569200, 1562572800, 
    1562576400, 1562580000, 1562583600, 1562587200, 1562590800, 1562594400, 
    1562598000, 1562601600, 1562605200, 1562608800, 1562612400, 1562616000, 
    1562619600, 1562623200, 1562626800, 1562630400, 1562634000, 1562637600, 
    1562641200, 1562644800, 1562648400, 1562652000, 1562551200, 1562655600, 
    1562659200, 1562662800, 1562666400, 1562670000, 1562673600, 1562677200, 
    1562680800, 1562684400, 1562688000, 1562691600, 1562695200, 1562698800, 
    1562702400, 1562706000, 1562709600, 1562713200, 1562716800, 1562720400, 
    1562724000, 1562727600, 1562731200, 1562734800, 1562738400, 1562742000, 
    1562745600, 1562749200, 1562756400, 1562760000, 1562763600, 1562767200, 
    1562770800, 1562774400, 1562778000, 1562781600, 1562785200, 1562788800, 
    1562792400, 1562796000, 1562799600, 1562803200, 1562806800, 1562810400, 
    1562814000, 1562817600, 1562821200, 1562824800, 1562828400, 1562832000, 
    1562835600, 1562839200, 1562842800, 1562846400, 1562850000, 1562853600, 
    1562857200, 1562860800, 1562864400, 1562868000, 1562871600, 1562875200, 
    1562878800, 1562882400, 1562886000, 1562889600, 1562893200, 1562896800, 
    1562900400, 1562904000, 1562907600, 1562911200, 1562914800, 1562918400, 
    1562922000, 1562925600, 1562929200, 1562932800, 1562936400, 1562940000, 
    1562943600, 1562947200, 1562950800, 1562954400, 1562958000, 1562961600, 
    1562965200, 1562968800, 1562972400, 1562976000, 1562979600, 1562983200, 
    1562986800, 1562990400, 1562994000, 1562997600, 1563001200, 1563004800, 
    1563008400, 1563012000, 1563015600, 1563019200, 1563022800, 1563026400, 
    1563030000, 1563033600, 1563037200, 1563040800, 1563044400, 1563048000, 
    1563051600, 1563055200, 1563058800, 1563062400, 1563066000, 1563069600, 
    1563073200, 1563076800, 1563080400, 1563084000, 1563087600, 1563091200, 
    1563094800, 1563098400, 1563102000, 1563105600, 1563109200, 1563112800, 
    1563116400, 1563120000, 1563123600, 1563127200, 1563130800, 1563134400, 
    1563138000, 1563141600, 1563145200, 1563148800, 1563152400, 1563156000, 
    1563159600, 1563163200, 1563166800, 1563170400, 1563174000, 1563177600, 
    1563181200, 1563184800, 1563188400, 1563192000, 1563195600, 1563199200, 
    1563202800, 1563206400, 1563210000, 1563213600, 1563217200, 1563220800, 
    1563224400, 1563228000, 1563231600, 1563235200, 1563238800, 1563242400, 
    1563246000, 1563249600, 1563253200, 1563256800, 1563260400, 1563264000, 
    1563267600, 1563271200, 1563274800, 1562752800, 1563278400, 1563282000, 
    1563285600, 1563289200, 1563292800, 1563296400, 1563300000, 1563303600, 
    1563307200, 1563310800, 1563314400, 1563318000, 1563321600, 1563325200, 
    1563328800, 1563332400, 1563336000, 1563339600, 1563343200, 1563346800, 
    1563350400, 1563354000, 1563357600, 1563361200, 1563364800, 1563368400, 
    1563372000, 1563375600, 1563379200, 1563382800, 1563386400, 1563390000, 
    1563393600, 1563397200, 1563400800, 1563404400, 1563408000, 1563411600, 
    1563415200, 1563418800, 1563422400, 1563426000, 1563429600, 1563433200, 
    1563436800, 1563440400, 1563444000, 1563447600, 1563451200, 1563454800, 
    1563458400, 1563462000, 1563465600, 1563469200, 1563472800, 1563476400, 
    1563480000, 1563483600, 1563487200, 1563490800, 1563494400, 1563498000, 
    1563501600, 1563505200, 1563508800, 1563512400, 1563516000, 1563519600, 
    1563523200, 1563526800, 1563530400, 1563534000, 1563537600, 1563541200, 
    1563544800, 1563548400, 1563552000, 1563555600, 1563559200, 1563562800, 
    1563566400, 1563570000, 1563573600, 1563577200, 1563580800, 1563584400, 
    1563588000, 1563591600, 1563595200, 1563598800, 1563602400, 1563606000, 
    1563609600, 1563613200, 1563616800, 1563620400, 1563624000, 1563627600, 
    1563631200, 1563634800, 1563638400, 1563642000, 1563645600, 1563649200, 
    1563652800, 1563656400, 1563660000, 1563663600, 1563667200, 1563670800, 
    1563674400, 1563678000, 1563681600, 1563685200, 1563688800, 1563692400, 
    1563696000, 1563699600, 1563703200, 1563706800, 1563710400, 1563714000, 
    1563717600, 1563721200, 1563724800, 1563728400, 1563732000, 1563735600, 
    1563739200, 1563742800, 1563746400, 1563750000, 1563753600, 1563757200, 
    1563760800, 1563764400, 1563768000, 1563771600, 1563775200, 1563778800, 
    1563782400, 1563786000, 1563789600, 1563793200, 1563796800, 1563800400, 
    1563804000, 1563807600, 1563811200, 1563814800, 1563818400, 1563822000, 
    1563825600, 1563829200, 1563832800, 1563836400, 1563840000, 1563843600, 
    1563847200, 1563850800, 1563854400, 1563858000, 1563861600, 1563865200, 
    1563868800, 1563872400, 1563876000, 1563879600, 1563883200, 1563886800, 
    1563890400, 1563894000, 1563897600, 1563901200, 1563904800, 1563908400, 
    1563912000, 1563915600, 1563919200, 1563922800, 1563926400, 1563930000, 
    1563933600, 1563937200, 1563940800, 1563944400, 1563948000, 1563951600, 
    1563955200, 1563958800, 1563962400, 1563966000, 1563969600, 1563973200, 
    1563976800, 1563980400, 1563984000, 1563987600, 1563991200, 1563994800, 
    1563998400, 1564002000, 1564005600, 1564009200, 1564012800, 1564016400, 
    1564020000, 1564023600, 1564027200, 1564030800, 1564034400, 1564038000, 
    1564041600, 1564045200, 1564048800, 1564052400, 1564056000, 1564059600, 
    1564063200, 1564066800, 1564070400, 1564074000, 1564077600, 1564081200, 
    1564084800, 1564088400, 1564092000, 1564095600, 1564099200, 1564102800, 
    1564106400, 1564110000, 1564113600, 1564117200, 1564120800, 1564124400, 
    1564128000, 1564131600, 1564135200, 1564138800, 1564142400, 1564146000, 
    1564149600, 1564153200, 1564156800, 1564160400, 1564164000, 1564167600, 
    1564171200, 1564174800, 1564178400, 1564182000, 1564185600, 1564189200, 
    1564192800, 1564196400, 1564200000, 1564203600, 1564207200, 1564210800, 
    1564214400, 1564218000, 1564221600, 1564225200, 1564228800, 1564232400, 
    1564236000, 1564239600, 1564243200, 1564246800, 1564250400, 1564254000, 
    1564257600, 1564261200, 1564264800, 1564268400, 1564272000, 1564275600, 
    1564279200, 1564282800, 1564286400, 1564290000, 1564293600, 1564297200, 
    1564300800, 1564304400, 1564308000, 1564311600, 1564315200, 1564318800, 
    1564322400, 1564326000, 1564329600, 1564333200, 1564336800, 1564340400, 
    1564344000, 1564347600, 1564351200, 1564354800, 1564358400, 1564362000, 
    1564365600, 1564369200, 1564372800, 1564376400, 1564380000, 1564383600, 
    1564387200, 1564390800, 1564394400, 1564398000, 1564401600, 1564405200, 
    1564408800, 1564412400, 1564416000, 1564419600, 1564423200, 1564426800, 
    1564430400, 1564434000, 1564437600, 1564441200, 1564444800, 1564448400, 
    1564452000, 1564455600, 1564459200, 1564462800, 1564466400, 1564470000, 
    1564473600, 1564477200, 1564480800, 1564484400, 1564488000, 1564491600, 
    1564495200, 1564498800, 1564502400, 1564506000, 1564509600, 1564513200, 
    1564516800, 1564520400, 1564524000, 1564527600, 1564531200, 1564534800, 
    1564538400, 1564542000, 1564545600, 1564549200, 1564552800, 1564556400, 
    1564560000, 1564563600, 1564567200, 1564570800, 1564574400, 1564578000, 
    1564581600, 1564585200, 1564588800, 1564592400, 1564596000, 1564599600, 
    1564603200, 1564606800, 1564610400, 1564614000, 1564617600, 1564621200, 
    1564624800, 1564628400, 1564632000, 1564635600, 1564639200, 1564642800, 
    1564646400, 1564650000, 1564653600, 1564657200, 1564660800, 1564664400, 
    1564668000, 1564671600, 1564675200, 1564678800, 1564682400, 1564686000, 
    1564689600, 1564693200, 1564696800, 1564700400, 1564704000, 1564707600, 
    1564711200, 1564714800, 1564718400, 1564722000, 1564725600, 1564729200, 
    1564732800, 1564736400, 1564740000, 1564743600, 1564747200, 1564750800, 
    1564754400, 1564758000, 1564761600, 1564765200, 1564768800, 1564772400, 
    1564776000, 1564779600, 1564783200, 1564786800, 1564790400, 1564794000, 
    1564797600, 1564801200, 1564804800, 1564808400, 1564812000, 1564815600, 
    1564819200, 1564822800, 1564826400, 1564830000, 1564833600, 1564837200, 
    1564840800, 1564844400, 1564848000, 1564851600, 1564855200, 1564858800, 
    1564862400, 1564866000, 1564869600, 1564873200, 1564876800, 1564880400, 
    1564884000, 1564887600, 1564891200, 1564894800, 1564898400, 1564902000, 
    1564905600, 1564909200, 1564912800, 1564916400, 1564920000, 1564923600, 
    1564927200, 1564930800, 1564934400, 1564938000, 1564941600, 1564945200, 
    1564948800, 1564952400, 1564956000, 1564959600, 1564963200, 1564966800, 
    1564970400, 1564974000, 1564977600, 1564981200, 1564984800, 1564988400, 
    1564992000, 1564995600, 1564999200, 1565002800, 1565006400, 1565010000, 
    1565013600, 1565017200, 1565020800, 1565024400, 1565028000, 1565031600, 
    1565035200, 1565038800, 1565042400, 1565046000, 1565049600, 1565053200, 
    1565056800, 1565060400, 1565064000, 1565067600, 1565071200, 1565074800, 
    1565078400, 1565082000, 1565085600, 1565089200, 1565092800, 1565096400, 
    1565100000, 1565103600, 1565107200, 1565110800, 1565114400, 1565118000, 
    1565121600, 1565125200, 1565128800, 1565132400, 1565136000, 1565139600, 
    1565143200, 1565146800, 1565150400, 1565154000, 1565157600, 1565161200, 
    1565164800, 1565168400, 1565172000, 1565175600, 1565179200, 1565182800, 
    1565186400, 1565190000, 1565193600, 1565197200, 1565200800, 1565204400, 
    1565208000, 1565211600, 1565215200, 1565218800, 1565222400, 1565226000, 
    1565229600, 1565233200, 1565236800, 1565240400, 1565244000, 1565247600, 
    1565251200, 1565254800, 1565258400, 1565262000, 1565265600, 1565269200, 
    1565272800, 1565276400, 1565280000, 1565283600, 1565287200, 1565290800, 
    1565294400, 1565298000, 1565301600, 1565305200, 1565308800, 1565312400, 
    1565316000, 1565319600, 1565323200, 1565326800, 1565330400, 1565334000, 
    1565337600, 1565341200, 1565344800, 1565348400, 1565352000, 1565355600, 
    1565359200, 1565362800, 1565366400, 1565370000, 1565373600, 1565377200, 
    1565380800, 1565384400, 1565388000, 1565391600, 1565395200, 1565398800, 
    1565402400, 1565406000, 1565409600, 1565413200, 1565416800, 1565420400, 
    1565424000, 1565427600, 1565431200, 1565434800, 1565438400, 1565442000, 
    1565445600, 1565449200, 1565452800, 1565456400, 1565460000, 1565463600, 
    1565467200, 1565470800, 1565474400, 1565478000, 1565481600, 1565485200, 
    1565488800, 1565492400, 1565496000, 1565499600, 1565503200, 1565506800, 
    1565510400, 1565514000, 1565517600, 1565521200, 1565524800, 1565528400, 
    1565532000, 1565535600, 1565539200, 1565542800, 1565546400, 1565550000, 
    1565553600, 1565557200, 1565560800, 1565564400, 1565568000, 1565571600, 
    1565575200, 1565578800, 1565582400, 1565586000, 1565589600, 1565593200, 
    1565596800, 1565600400, 1565604000, 1565607600, 1565611200, 1565614800, 
    1565618400, 1565622000, 1565625600, 1565629200, 1565632800, 1565636400, 
    1565640000, 1565643600, 1565647200, 1565650800, 1565654400, 1565658000, 
    1565661600, 1565665200, 1565668800, 1565672400, 1565676000, 1565679600, 
    1565683200, 1565686800, 1565690400, 1565694000, 1565697600, 1565701200, 
    1565704800, 1565708400, 1565712000, 1565715600, 1565719200, 1565722800, 
    1565726400, 1565730000, 1565733600, 1565737200, 1565740800, 1565744400, 
    1565748000, 1565751600, 1565755200, 1565758800, 1565762400, 1565766000, 
    1565769600, 1565773200, 1565776800, 1565780400, 1565784000, 1565787600, 
    1565791200, 1565794800, 1565798400, 1565802000, 1565805600, 1565809200, 
    1565812800, 1565816400, 1565820000, 1565823600, 1565827200, 1565830800, 
    1565834400, 1565838000, 1565841600, 1565845200, 1565848800, 1565852400, 
    1565856000, 1565859600, 1565863200, 1565866800, 1565870400, 1565874000, 
    1565877600, 1565881200, 1565884800, 1565888400, 1565892000, 1565895600, 
    1565899200, 1565902800, 1565906400, 1565910000, 1565913600, 1565917200, 
    1565920800, 1565924400, 1565928000, 1565931600, 1565935200, 1565938800, 
    1565942400, 1565946000, 1565949600, 1565953200, 1565956800, 1565960400, 
    1565964000, 1565967600, 1565971200, 1565974800, 1565978400, 1565982000, 
    1565985600, 1565989200, 1565992800, 1565996400, 1566000000, 1566003600, 
    1566007200, 1566010800, 1566014400, 1566018000, 1566021600, 1566025200, 
    1566028800, 1566032400, 1566036000, 1566039600, 1566043200, 1566046800, 
    1566050400, 1566054000, 1566057600, 1566061200, 1566064800, 1566068400, 
    1566072000, 1566075600, 1566079200, 1566082800, 1566086400, 1566090000, 
    1566093600, 1566097200, 1566100800, 1566104400, 1566108000, 1566111600, 
    1566115200, 1566118800, 1566122400, 1566126000, 1566129600, 1566133200, 
    1566136800, 1566140400, 1566144000, 1566147600, 1566151200, 1566154800, 
    1566158400, 1566162000, 1566165600, 1566169200, 1566172800, 1566176400, 
    1566180000, 1566183600, 1566187200, 1566190800, 1566194400, 1566198000, 
    1566201600, 1566205200, 1566208800, 1566212400, 1566216000, 1566219600, 
    1566223200, 1566226800, 1566230400, 1566234000, 1566237600, 1566241200, 
    1566244800, 1566248400, 1566252000, 1566255600, 1566259200, 1566262800, 
    1566266400, 1566270000, 1566273600, 1566277200, 1566280800, 1566284400, 
    1566288000, 1566291600, 1566295200, 1566298800, 1566302400, 1566306000, 
    1566309600, 1566313200, 1566316800, 1566320400, 1566324000, 1566327600, 
    1566331200, 1566334800, 1566338400, 1566342000, 1566345600, 1566349200, 
    1566352800, 1566356400, 1566360000, 1566363600, 1566367200, 1566370800, 
    1566374400, 1566378000, 1566381600, 1566385200, 1566388800, 1566392400, 
    1566396000, 1566399600, 1566403200, 1566406800, 1566410400, 1566414000, 
    1566417600, 1566421200, 1566424800, 1566428400, 1566432000, 1566435600, 
    1566439200, 1566442800, 1566446400, 1566450000, 1566453600, 1566457200, 
    1566460800, 1566464400, 1566468000, 1566471600, 1566475200, 1566478800, 
    1566482400, 1566486000, 1566489600, 1566493200, 1566496800, 1566500400, 
    1566504000, 1566511200, 1566514800, 1566518400, 1566522000, 1566529200, 
    1566532800, 1566536400, 1566507600, 1566525600, 1566543600, 1566547200, 
    1566550800, 1566554400, 1566561600, 1566565200, 1566568800, 1566572400, 
    1566576000, 1566579600, 1566586800, 1566590400, 1566594000, 1566604800, 
    1566608400, 1566612000, 1566615600, 1566619200, 1566622800, 1566626400, 
    1566540000, 1566558000, 1566583200, 1566597600, 1566601200, 1566630000, 
    1566633600, 1566637200, 1566640800, 1566644400, 1566648000, 1566651600, 
    1566655200, 1566658800, 1566662400, 1566669600, 1566673200, 1566676800, 
    1566680400, 1566684000, 1566687600, 1566691200, 1566694800, 1566698400, 
    1566702000, 1566705600, 1566709200, 1566712800, 1566666000, 1566716400, 
    1566720000, 1566723600, 1566730800, 1566734400, 1566738000, 1566741600, 
    1566745200, 1566748800, 1566752400, 1566756000, 1566759600, 1566763200, 
    1566770400, 1566774000, 1566777600, 1566781200, 1566784800, 1566788400, 
    1566792000, 1566795600, 1566799200, 1566727200, 1566766800, 1566802800, 
    1566806400, 1566813600, 1566817200, 1566824400, 1566828000, 1566831600, 
    1566835200, 1566838800, 1566846000, 1566849600, 1566853200, 1566860400, 
    1566867600, 1566871200, 1566874800, 1566878400, 1566882000, 1566810000, 
    1566820800, 1566842400, 1566856800, 1566864000, 1566885600, 1566892800, 
    1566896400, 1566900000, 1566903600, 1566907200, 1566910800, 1566914400, 
    1566918000, 1566921600, 1566928800, 1566932400, 1566936000, 1566939600, 
    1566943200, 1566946800, 1566950400, 1566954000, 1566957600, 1566961200, 
    1566964800, 1566968400, 1566972000, 1566889200, 1566925200, 1566975600, 
    1566979200, 1566982800, 1566986400, 1566990000, 1566993600, 1566997200, 
    1567000800, 1567004400, 1567008000, 1567011600, 1567015200, 1567018800, 
    1567022400, 1567026000, 1567029600, 1567033200, 1567036800, 1567040400, 
    1567044000, 1567047600, 1567051200, 1567054800, 1567058400, 1567062000, 
    1567065600, 1567069200, 1567072800, 1567076400, 1567080000, 1567083600, 
    1567087200, 1567090800, 1567094400, 1567098000, 1567101600, 1567105200, 
    1567108800, 1567112400, 1567116000, 1567119600, 1567123200, 1567126800, 
    1567130400, 1567134000, 1567137600, 1567141200, 1567144800, 1567148400, 
    1567152000, 1567155600, 1567159200, 1567162800, 1567166400, 1567170000, 
    1567173600, 1567177200, 1567180800, 1567184400, 1567188000, 1567191600, 
    1567195200, 1567198800, 1567202400, 1567206000, 1567209600, 1567213200, 
    1567216800, 1567220400, 1567224000, 1567227600, 1567231200, 1567234800, 
    1567238400, 1567242000, 1567245600, 1567249200, 1567252800, 1567256400, 
    1567260000, 1567263600, 1567267200, 1567270800, 1567274400, 1567278000, 
    1567281600, 1567285200, 1567288800, 1567292400, 1567296000, 1567299600, 
    1567303200, 1567306800, 1567310400, 1567314000, 1567317600, 1567321200, 
    1567324800, 1567328400, 1567332000, 1567335600, 1567339200, 1567342800, 
    1567346400, 1567350000, 1567353600, 1567357200, 1567360800, 1567364400, 
    1567368000, 1567371600, 1567375200, 1567378800, 1567382400, 1567386000, 
    1567389600, 1567393200, 1567396800, 1567400400, 1567404000, 1567407600, 
    1567411200, 1567414800, 1567418400, 1567422000, 1567425600, 1567429200, 
    1567432800, 1567436400, 1567440000, 1567443600, 1567447200, 1567450800, 
    1567454400, 1567458000, 1567461600, 1567465200, 1567468800, 1567472400, 
    1567476000, 1567479600, 1567483200, 1567486800, 1567490400, 1567494000, 
    1567497600, 1567501200, 1567504800 ;

 latitude = 78.6557 ;

 longitude = 16.3603 ;

 station_id = "SN99880" ;

 air_temperature_2m = 254.45, 254.25, 254.05, 253.85, 253.95, 254.35, 255.15, 
    256.15, 255.85, 256.85, 257.05, 256.95, 257.15, 257.15, 257.05, 256.95, 
    257.15, 257.15, 256.45, 255.95, 259.25, 259.05, 258.85, 259.45, 260.95, 
    261.65, 262.15, 262.75, 263.75, 264.65, 265.45, 266.05, 265.05, 264.95, 
    265.05, 265.25, 265.25, 265.15, 265.15, 265.35, 265.25, 265.15, 264.95, 
    264.65, 263.65, 263.45, 263.45, 263.75, 264.15, 264.35, 264.15, 263.75, 
    263.55, 263.25, 263.25, 263.05, 262.05, 261.45, 261.15, 261.25, 260.85, 
    260.65, 260.45, 260.15, 259.95, 259.45, 259.25, 258.95, 257.65, 257.45, 
    257.25, 265.95, 265.75, 265.35, 264.95, 264.55, 265.15, 265.35, 264.35, 
    264.35, 264.05, 264.55, 264.85, 264.05, 264.45, 265.55, 264.75, 265.35, 
    266.15, 264.65, 265.55, 266.05, 265.65, 266.05, 265.95, 265.75, 265.95, 
    265.65, 265.95, 266.15, 266.15, 266.15, 266.85, 267.15, 266.75, 266.65, 
    266.65, 266.35, 266.65, 266.35, 265.85, 266.05, 265.95, 264.95, 264.85, 
    265.15, 264.85, 264.65, 264.55, 264.65, 264.55, 264.85, 264.95, 265.05, 
    264.75, 264.65, 264.65, 264.65, 264.25, 263.85, 263.45, 261.35, 261.35, 
    260.25, 260.05, 261.55, 260.95, 259.05, 260.75, 261.55, 259.65, 258.25, 
    259.65, 256.85, 255.65, 255.85, 256.15, 256.75, 257.55, 257.45, 257.55, 
    256.95, 256.95, 256.85, 257.95, 256.65, 256.35, 256.15, 255.95, 255.75, 
    255.65, 255.65, 255.45, 255.35, 255.25, 255.05, 255.05, 256.35, 256.65, 
    255.65, 255.35, 255.85, 255.65, 255.45, 255.55, 255.45, 255.65, 256.15, 
    256.15, 255.85, 256.05, 255.75, 256.25, 256.45, 255.15, 256.15, 257.05, 
    255.75, 257.55, 257.65, 257.15, 259.15, 257.85, 258.85, 259.65, 259.45, 
    258.95, 259.85, 261.35, 260.95, 260.75, 261.95, 264.25, 265.55, 265.45, 
    265.55, 265.95, 267.15, 267.75, 267.55, 267.75, 268.45, 268.75, 268.95, 
    268.95, 269.35, 269.25, 269.15, 269.05, 269.05, 269.15, 269.15, 269.15, 
    269.45, 269.45, 269.05, 269.25, 269.65, 269.55, 269.35, 269.35, 269.55, 
    269.05, 268.95, 269.25, 269.25, 269.35, 269.15, 269.25, 269.15, 269.15, 
    269.45, 269.65, 269.75, 269.75, 269.85, 270.15, 270.25, 270.45, 270.55, 
    270.35, 270.15, 269.75, 269.75, 269.35, 268.95, 268.95, 268.55, 267.95, 
    267.55, 267.15, 267.05, 266.75, 266.75, 266.95, 266.85, 266.75, 266.75, 
    263.05, 263.15, 266.25, 266.15, 266.25, 266.05, 266.15, 266.85, 265.45, 
    265.65, 267.45, 267.85, 266.65, 267.55, 268.15, 268.25, 268.35, 268.25, 
    269.05, 269.05, 268.95, 268.95, 268.95, 269.05, 269.65, 269.65, 268.15, 
    269.45, 269.55, 269.65, 269.65, 269.35, 269.05, 268.95, 268.95, 268.75, 
    268.45, 268.55, 268.35, 268.15, 268.05, 267.95, 268.05, 267.95, 268.05, 
    267.35, 265.95, 265.25, 263.85, 262.95, 264.45, 263.85, 266.75, 263.95, 
    264.85, 265.75, 264.25, 265.05, 265.15, 265.25, 265.45, 265.85, 267.15, 
    268.55, 269.45, 269.45, 269.35, 269.25, 268.95, 268.85, 268.85, 269.05, 
    268.75, 268.95, 269.55, 269.65, 269.65, 269.55, 269.75, 270.15, 269.95, 
    270.05, 270.35, 269.75, 268.45, 268.55, 267.75, 269.15, 267.65, 268.45, 
    268.25, 268.25, 266.15, 267.55, 268.35, 268.85, 268.95, 268.55, 269.45, 
    269.35, 268.85, 268.95, 269.65, 270.05, 270.05, 270.15, 269.45, 269.75, 
    269.45, 269.75, 268.15, 266.85, 267.15, 267.55, 269.05, 269.25, 269.15, 
    268.85, 268.95, 269.25, 268.45, 269.05, 269.75, 269.15, 268.95, 268.05, 
    267.05, 267.45, 268.05, 266.65, 266.45, 265.85, 268.05, 267.25, 267.15, 
    267.25, 267.85, 268.75, 269.35, 270.15, 270.15, 270.35, 270.45, 270.45, 
    270.55, 269.95, 266.75, 266.95, 266.85, 266.15, 265.45, 266.15, 266.85, 
    267.85, 266.95, 267.15, 266.75, 265.25, 265.65, 265.85, 265.15, 263.95, 
    264.95, 263.85, 262.75, 262.25, 263.05, 262.75, 262.55, 262.95, 262.85, 
    261.75, 262.75, 260.85, 261.95, 262.15, 261.55, 260.15, 262.25, 261.25, 
    261.35, 260.75, 260.35, 261.15, 261.45, 261.05, 260.45, 260.15, 260.15, 
    261.65, 260.75, 260.25, 259.35, 259.75, 260.25, 260.35, 258.65, 260.65, 
    262.45, 262.95, 263.25, 263.25, 263.75, 264.45, 264.15, 264.55, 265.15, 
    265.55, 265.75, 265.85, 266.65, 266.25, 266.85, 266.35, 266.95, 266.85, 
    266.75, 266.85, 266.95, 267.05, 267.65, 268.55, 267.75, 269.95, 268.65, 
    268.45, 268.15, 267.95, 267.55, 267.15, 266.25, 266.25, 265.75, 263.95, 
    264.45, 263.65, 264.25, 264.55, 265.35, 266.15, 266.45, 266.45, 266.85, 
    267.05, 267.15, 267.15, 267.55, 267.65, 267.85, 267.45, 267.35, 267.85, 
    267.25, 268.75, 268.35, 268.65, 267.95, 268.05, 268.45, 269.05, 269.65, 
    269.45, 269.65, 266.85, 266.95, 266.45, 267.05, 266.85, 266.95, 269.75, 
    272.65, 272.35, 272.75, 272.45, 272.55, 273.15, 272.65, 273.05, 273.85, 
    273.95, 274.05, 274.15, 273.45, 273.35, 272.45, 272.35, 272.25, 271.75, 
    272.05, 272.05, 272.05, 272.05, 272.55, 272.15, 271.95, 272.35, 272.75, 
    272.95, 273.25, 272.65, 272.35, 272.05, 271.35, 271.55, 270.95, 271.55, 
    271.95, 272.15, 272.05, 272.75, 274.05, 273.75, 273.25, 273.55, 274.15, 
    273.75, 274.05, 274.15, 273.85, 271.95, 270.85, 271.95, 271.65, 271.85, 
    272.45, 272.75, 273.25, 273.25, 273.25, 271.25, 271.45, 269.25, 270.55, 
    271.55, 271.55, 271.45, 272.45, 271.65, 271.65, 271.05, 269.75, 268.35, 
    268.25, 268.25, 266.55, 267.15, 267.75, 268.95, 269.75, 270.15, 270.55, 
    270.45, 270.15, 270.15, 270.35, 268.55, 267.75, 267.85, 266.45, 267.45, 
    267.35, 267.45, 267.65, 268.15, 268.55, 268.55, 268.95, 266.65, 264.15, 
    265.15, 267.15, 265.45, 265.85, 264.65, 264.65, 264.35, 265.15, 264.05, 
    263.25, 263.55, 264.45, 264.45, 264.45, 266.35, 266.05, 265.95, 266.65, 
    267.15, 266.85, 266.95, 266.75, 267.95, 267.25, 266.75, 268.05, 267.25, 
    264.45, 267.15, 266.35, 265.65, 266.75, 266.45, 265.45, 264.85, 264.95, 
    266.95, 267.45, 267.05, 267.05, 266.05, 267.35, 265.95, 267.05, 268.95, 
    270.25, 270.65, 270.55, 271.55, 271.25, 271.55, 271.05, 271.25, 270.15, 
    269.35, 267.45, 270.15, 269.65, 267.35, 267.65, 267.55, 267.45, 265.55, 
    267.45, 267.15, 266.65, 265.75, 267.75, 266.65, 267.35, 267.35, 268.45, 
    268.45, 268.85, 268.25, 268.15, 270.05, 269.65, 269.15, 267.85, 267.05, 
    265.95, 265.95, 265.75, 265.55, 264.95, 264.15, 263.95, 263.35, 262.85, 
    262.05, 261.55, 261.65, 260.95, 261.05, 260.95, 260.45, 260.95, 259.45, 
    257.85, 258.45, 257.45, 258.25, 257.05, 256.35, 256.35, 256.95, 257.45, 
    256.35, 256.75, 256.95, 256.45, 254.95, 256.55, 255.15, 255.95, 255.95, 
    256.15, 256.45, 256.95, 257.05, 257.85, 257.95, 257.75, 258.45, 259.25, 
    259.25, 259.65, 260.05, 260.65, 261.45, 262.85, 263.55, 264.45, 264.45, 
    264.65, 265.25, 267.05, 267.85, 266.45, 263.65, 262.45, 261.65, 260.65, 
    260.35, 260.65, 258.25, 257.25, 258.85, 258.95, 258.65, 258.65, 257.25, 
    257.65, 257.05, 256.55, 256.65, 255.85, 255.05, 257.15, 256.75, 258.35, 
    256.45, 256.45, 256.95, 258.15, 258.05, 257.15, 257.25, 257.45, 257.45, 
    258.25, 259.55, 261.05, 260.75, 261.35, 261.35, 261.65, 262.35, 263.05, 
    263.55, 264.05, 264.95, 266.15, 266.65, 267.35, 267.85, 268.35, 268.15, 
    268.45, 269.55, 270.05, 270.05, 271.75, 272.65, 271.55, 270.35, 269.25, 
    268.25, 267.25, 265.45, 264.35, 263.55, 263.25, 262.45, 263.25, 263.05, 
    263.45, 263.05, 262.55, 262.45, 262.15, 262.15, 262.45, 263.25, 263.45, 
    264.25, 264.75, 264.05, 263.25, 262.75, 263.25, 262.35, 260.55, 260.35, 
    262.55, 263.65, 263.85, 263.25, 262.45, 261.75, 261.35, 261.15, 262.15, 
    261.25, 260.95, 258.95, 258.45, 259.45, 258.85, 258.95, 260.05, 258.85, 
    261.35, 261.95, 261.65, 261.65, 260.85, 261.05, 261.35, 261.45, 260.95, 
    260.25, 260.05, 258.95, 257.95, 258.25, 259.35, 257.45, 257.85, 258.85, 
    255.95, 257.95, 260.15, 259.45, 259.05, 258.65, 258.25, 257.15, 256.75, 
    256.95, 255.85, 255.85, 255.75, 255.55, 255.75, 254.05, 254.05, 253.45, 
    254.35, 254.85, 251.75, 252.05, 252.75, 253.05, 252.65, 252.65, 253.15, 
    253.25, 253.75, 253.35, 253.45, 252.95, 252.45, 251.45, 251.65, 251.65, 
    251.75, 249.25, 251.45, 249.95, 250.85, 251.55, 251.35, 251.95, 251.75, 
    251.25, 252.55, 252.15, 259.15, 259.85, 260.35, 260.55, 260.85, 260.75, 
    260.55, 260.25, 259.65, 259.15, 258.45, 257.95, 257.65, 257.75, 257.35, 
    255.55, 255.65, 255.75, 255.75, 255.75, 255.55, 256.25, 256.15, 255.05, 
    255.65, 255.75, 255.35, 254.45, 254.95, 255.05, 254.85, 254.85, 254.75, 
    255.15, 255.55, 255.85, 255.65, 255.95, 255.35, 255.45, 256.65, 256.45, 
    257.45, 257.55, 256.85, 256.55, 257.15, 256.55, 257.35, 257.65, 256.45, 
    257.85, 257.25, 256.75, 256.45, 256.35, 257.25, 257.75, 258.25, 259.75, 
    258.25, 259.95, 260.25, 258.55, 261.15, 260.85, 262.85, 263.35, 264.75, 
    265.35, 264.95, 265.25, 264.05, 264.35, 264.45, 264.75, 264.85, 265.05, 
    265.15, 264.35, 263.25, 263.55, 263.55, 263.95, 266.15, 266.25, 265.85, 
    265.75, 265.85, 266.15, 266.15, 265.95, 265.75, 265.95, 265.55, 264.95, 
    264.35, 263.65, 263.05, 262.65, 262.65, 263.05, 263.15, 263.45, 264.35, 
    265.55, 266.75, 267.75, 268.75, 268.45, 272.15, 272.25, 271.55, 271.25, 
    271.25, 270.65, 270.95, 271.85, 273.45, 273.05, 273.55, 272.95, 272.85, 
    272.75, 272.75, 273.25, 272.75, 272.65, 272.35, 272.15, 272.05, 272.05, 
    272.25, 272.35, 272.25, 272.15, 271.85, 271.55, 271.35, 271.75, 272.15, 
    272.35, 273.15, 273.15, 273.25, 273.35, 273.65, 273.55, 273.15, 273.25, 
    273.15, 273.25, 273.45, 273.75, 273.95, 274.05, 273.95, 274.25, 274.35, 
    274.15, 274.55, 274.75, 274.35, 274.25, 274.55, 274.35, 274.25, 274.45, 
    274.45, 274.05, 274.05, 274.35, 274.55, 274.75, 274.35, 274.05, 274.65, 
    274.35, 273.85, 273.55, 273.85, 273.45, 274.25, 274.75, 274.25, 274.65, 
    274.85, 274.75, 274.45, 274.65, 274.75, 274.25, 274.25, 274.55, 274.75, 
    273.85, 273.95, 274.35, 273.95, 273.85, 274.15, 274.55, 273.95, 273.05, 
    274.25, 273.35, 272.25, 271.85, 271.95, 271.65, 271.85, 271.35, 271.15, 
    271.55, 271.65, 271.65, 272.55, 273.15, 272.95, 272.75, 272.35, 272.15, 
    271.85, 271.25, 271.35, 270.95, 271.05, 270.85, 270.85, 270.35, 269.35, 
    267.65, 267.45, 268.75, 267.85, 268.35, 267.95, 268.05, 267.45, 266.55, 
    266.95, 266.25, 264.75, 265.45, 265.55, 265.85, 266.55, 265.45, 266.05, 
    266.95, 267.45, 268.25, 268.05, 267.75, 268.85, 268.85, 268.05, 268.05, 
    268.95, 268.65, 268.75, 269.05, 270.15, 270.75, 270.45, 272.15, 272.35, 
    272.25, 273.05, 272.95, 272.65, 272.25, 273.25, 274.25, 275.15, 276.05, 
    275.35, 276.35, 274.75, 274.55, 274.95, 274.85, 275.05, 274.55, 274.45, 
    273.65, 273.25, 273.25, 273.25, 273.25, 272.95, 272.95, 272.45, 272.85, 
    274.75, 274.05, 273.65, 273.85, 273.85, 273.55, 273.05, 272.95, 272.85, 
    272.75, 272.85, 272.55, 271.65, 270.55, 269.85, 268.65, 266.95, 266.55, 
    267.05, 266.65, 266.55, 265.95, 265.65, 266.35, 265.95, 266.35, 265.85, 
    266.15, 265.35, 266.65, 265.65, 265.05, 264.75, 263.95, 263.75, 262.85, 
    262.55, 262.75, 261.35, 262.25, 263.35, 263.15, 264.55, 264.35, 264.25, 
    265.25, 265.55, 264.55, 264.25, 263.45, 263.15, 262.95, 263.25, 264.05, 
    264.55, 262.55, 263.55, 262.95, 263.05, 264.55, 264.95, 265.05, 265.85, 
    266.05, 266.05, 267.05, 267.35, 267.65, 269.95, 269.75, 269.85, 270.55, 
    270.05, 270.25, 270.25, 271.45, 270.95, 271.25, 272.15, 271.65, 271.65, 
    271.55, 271.35, 271.55, 274.05, 274.25, 274.45, 274.25, 274.05, 274.75, 
    274.85, 274.05, 274.15, 274.65, 274.65, 274.55, 274.15, 273.65, 273.35, 
    273.05, 272.75, 271.35, 271.65, 271.55, 268.85, 266.95, 267.15, 266.85, 
    266.35, 266.45, 265.85, 265.25, 265.15, 265.15, 265.45, 265.75, 266.35, 
    266.35, 266.05, 266.05, 266.35, 266.15, 264.75, 265.95, 265.35, 264.25, 
    263.75, 264.65, 263.55, 263.55, 262.65, 262.15, 263.75, 263.35, 263.25, 
    262.65, 262.15, 262.75, 262.05, 261.65, 261.75, 261.85, 263.35, 262.55, 
    261.65, 261.45, 261.55, 260.85, 263.75, 262.15, 262.55, 262.65, 262.45, 
    261.35, 260.55, 261.75, 260.65, 260.15, 260.25, 260.55, 260.75, 261.25, 
    260.75, 259.95, 260.15, 260.75, 262.25, 260.95, 260.05, 261.05, 258.95, 
    260.55, 260.35, 258.55, 261.45, 259.85, 260.45, 260.15, 259.55, 258.05, 
    259.85, 260.45, 258.65, 259.35, 259.55, 260.05, 259.35, 258.85, 259.25, 
    258.65, 259.45, 259.85, 260.25, 259.15, 257.55, 258.45, 259.05, 259.75, 
    261.55, 261.15, 260.95, 260.95, 260.65, 261.35, 260.45, 259.45, 260.45, 
    258.85, 261.15, 260.95, 262.65, 263.25, 263.65, 263.45, 264.05, 266.65, 
    265.25, 265.65, 267.85, 267.95, 268.05, 267.75, 268.15, 268.45, 268.55, 
    268.35, 267.95, 267.35, 267.15, 266.75, 266.75, 266.45, 266.35, 265.75, 
    265.95, 265.45, 265.45, 265.85, 265.85, 265.95, 265.55, 264.95, 265.95, 
    264.95, 264.15, 263.55, 264.75, 264.55, 264.15, 261.95, 261.25, 263.45, 
    264.85, 266.55, 265.75, 265.65, 262.25, 259.85, 263.15, 263.35, 267.45, 
    267.75, 268.35, 268.45, 268.55, 268.05, 267.45, 266.95, 266.25, 265.35, 
    262.05, 261.65, 260.55, 262.55, 259.35, 260.55, 260.45, 259.25, 261.65, 
    261.35, 261.55, 262.05, 263.45, 263.65, 264.05, 263.75, 263.55, 263.35, 
    262.05, 261.35, 261.95, 263.75, 262.65, 261.95, 260.35, 261.05, 261.45, 
    261.85, 261.95, 260.85, 261.45, 261.65, 262.85, 262.85, 263.05, 262.85, 
    264.15, 263.95, 263.65, 263.75, 263.75, 263.95, 264.05, 263.95, 263.95, 
    264.25, 264.75, 265.35, 265.55, 266.45, 266.85, 267.65, 267.85, 267.95, 
    268.15, 268.35, 269.25, 269.25, 268.45, 267.15, 266.25, 264.85, 265.65, 
    266.55, 266.25, 266.95, 266.85, 266.35, 265.65, 264.35, 263.85, 263.25, 
    262.55, 261.85, 261.85, 261.15, 260.35, 259.95, 258.65, 258.55, 258.45, 
    255.75, 254.25, 255.35, 256.45, 255.05, 257.35, 258.65, 258.75, 259.15, 
    261.15, 259.95, 261.45, 261.55, 262.15, 262.45, 262.25, 262.35, 261.45, 
    262.55, 262.05, 262.25, 263.15, 263.15, 263.15, 262.95, 262.65, 262.25, 
    262.05, 261.25, 260.55, 260.85, 261.25, 261.45, 258.35, 258.85, 259.05, 
    260.55, 262.65, 264.55, 265.15, 265.35, 265.15, 263.85, 263.45, 264.85, 
    264.95, 265.15, 265.55, 265.75, 265.35, 264.95, 264.75, 264.35, 263.85, 
    261.95, 260.25, 259.55, 260.05, 258.75, 258.75, 258.15, 257.75, 257.35, 
    256.95, 257.95, 257.85, 258.45, 259.15, 257.85, 260.25, 259.05, 260.85, 
    261.45, 260.75, 260.75, 260.05, 260.35, 259.95, 259.45, 258.45, 259.95, 
    259.25, 257.85, 258.05, 258.55, 258.35, 260.65, 259.35, 257.05, 257.35, 
    256.85, 256.25, 257.05, 256.35, 257.35, 256.55, 255.75, 255.35, 255.25, 
    256.25, 255.45, 256.85, 257.35, 257.45, 256.35, 256.95, 254.55, 256.15, 
    255.55, 255.75, 255.85, 255.75, 256.95, 257.05, 256.55, 256.35, 255.45, 
    256.85, 256.85, 256.15, 255.95, 256.85, 256.35, 255.25, 256.95, 256.55, 
    256.35, 255.85, 255.25, 255.15, 256.45, 255.75, 255.75, 256.05, 256.55, 
    256.85, 256.55, 255.65, 256.65, 256.35, 254.55, 256.65, 257.05, 254.85, 
    256.45, 255.25, 255.55, 255.15, 256.55, 256.25, 256.65, 256.25, 257.25, 
    255.55, 255.85, 254.65, 256.05, 255.25, 255.05, 254.25, 256.85, 256.05, 
    256.05, 255.55, 256.15, 254.85, 255.95, 254.85, 255.45, 256.15, 257.05, 
    255.45, 256.15, 256.85, 256.65, 256.25, 254.85, 254.65, 254.45, 255.35, 
    255.95, 256.05, 256.15, 255.05, 255.55, 255.75, 256.25, 255.25, 256.45, 
    255.65, 255.65, 256.35, 254.95, 256.65, 255.75, 254.85, 254.45, 255.55, 
    255.45, 254.45, 255.55, 255.75, 255.65, 255.15, 254.35, 253.85, 254.35, 
    255.25, 255.75, 255.75, 255.65, 255.45, 256.55, 256.85, 256.95, 256.85, 
    256.25, 256.65, 257.55, 258.05, 257.25, 258.05, 258.65, 259.05, 258.95, 
    257.45, 256.85, 258.85, 257.85, 259.85, 260.35, 260.25, 262.05, 263.45, 
    262.25, 261.45, 261.15, 261.85, 263.15, 263.75, 261.55, 265.55, 261.25, 
    266.05, 264.25, 265.45, 264.95, 264.55, 264.35, 264.55, 264.55, 264.55, 
    265.05, 265.35, 265.55, 265.55, 265.45, 265.05, 264.95, 264.85, 264.75, 
    264.35, 263.85, 264.15, 261.05, 257.85, 261.15, 259.35, 258.35, 259.55, 
    258.95, 258.75, 260.45, 257.85, 259.55, 258.85, 260.25, 258.75, 257.25, 
    259.25, 258.75, 259.15, 257.85, 258.85, 258.25, 259.25, 258.95, 260.25, 
    258.65, 258.55, 259.15, 260.15, 259.55, 258.45, 258.45, 257.35, 258.15, 
    258.25, 257.45, 258.65, 258.65, 258.35, 257.85, 258.55, 257.95, 259.25, 
    257.65, 258.35, 258.05, 258.25, 257.85, 257.55, 259.45, 257.55, 257.75, 
    256.85, 258.25, 256.55, 257.75, 258.35, 258.05, 257.45, 258.05, 258.25, 
    258.55, 258.35, 258.75, 259.15, 259.35, 259.65, 260.15, 261.25, 262.25, 
    262.75, 263.05, 263.95, 265.25, 267.15, 266.95, 268.95, 269.65, 269.85, 
    269.85, 268.25, 268.95, 269.35, 270.15, 270.35, 269.55, 268.85, 268.95, 
    268.85, 268.65, 268.05, 267.75, 264.95, 265.75, 267.95, 269.05, 267.35, 
    267.75, 268.85, 267.25, 268.15, 267.15, 267.25, 268.05, 267.85, 266.75, 
    266.85, 264.05, 265.65, 266.35, 265.25, 267.15, 265.15, 265.55, 266.15, 
    267.55, 265.05, 265.75, 266.05, 264.35, 264.85, 263.75, 263.35, 262.95, 
    263.35, 261.65, 261.75, 262.55, 262.55, 262.25, 261.65, 261.95, 262.95, 
    262.35, 263.05, 262.75, 263.35, 263.65, 263.75, 263.75, 263.55, 263.65, 
    263.45, 263.05, 263.55, 266.05, 266.65, 266.35, 267.05, 266.45, 267.35, 
    266.15, 265.85, 264.25, 264.95, 265.85, 265.65, 265.65, 266.55, 266.05, 
    266.45, 266.85, 268.35, 268.25, 268.15, 267.45, 268.55, 268.85, 268.75, 
    268.15, 267.35, 268.05, 268.95, 268.75, 268.85, 268.75, 268.55, 269.05, 
    268.35, 269.35, 269.35, 269.35, 269.75, 269.55, 268.75, 269.05, 268.75, 
    270.55, 271.05, 270.85, 271.35, 269.85, 270.15, 270.45, 268.95, 269.65, 
    269.55, 268.35, 268.75, 269.45, 270.05, 269.25, 269.05, 268.35, 268.45, 
    268.55, 268.65, 268.75, 268.05, 269.65, 270.15, 270.35, 270.05, 270.35, 
    270.75, 270.05, 269.75, 271.55, 273.15, 272.85, 272.95, 271.85, 271.05, 
    270.65, 267.75, 268.05, 267.15, 264.65, 264.75, 265.35, 266.15, 266.65, 
    266.85, 267.25, 267.45, 268.05, 268.25, 268.25, 268.15, 268.25, 268.85, 
    268.75, 268.95, 268.75, 269.05, 269.15, 269.65, 271.15, 272.65, 272.45, 
    271.75, 271.35, 270.35, 271.25, 271.35, 271.75, 271.85, 271.65, 271.95, 
    272.05, 271.95, 271.25, 271.55, 271.15, 271.25, 270.75, 271.45, 269.55, 
    270.55, 270.45, 270.05, 271.25, 272.05, 272.85, 274.75, 274.65, 274.45, 
    274.25, 274.15, 273.95, 274.35, 274.55, 274.65, 274.75, 274.85, 274.45, 
    274.25, 274.25, 274.05, 274.35, 273.15, 272.95, 272.85, 272.55, 272.95, 
    272.65, 272.05, 271.95, 271.35, 271.35, 271.05, 270.65, 271.85, 270.95, 
    270.75, 270.65, 270.75, 270.15, 269.85, 269.85, 270.05, 269.65, 269.45, 
    269.15, 269.75, 268.75, 268.35, 267.95, 267.85, 268.25, 268.65, 267.95, 
    268.95, 268.45, 268.55, 267.65, 266.15, 265.85, 265.55, 265.45, 264.25, 
    262.75, 262.05, 261.35, 260.75, 260.35, 259.35, 256.85, 257.15, 257.25, 
    256.75, 257.75, 257.45, 257.65, 256.95, 257.15, 256.65, 256.15, 256.05, 
    255.85, 255.35, 255.85, 256.65, 256.05, 255.05, 254.75, 255.05, 255.65, 
    258.35, 258.85, 259.85, 259.55, 260.05, 259.55, 260.45, 260.65, 260.95, 
    261.25, 262.95, 263.25, 263.65, 264.45, 264.45, 263.95, 263.85, 263.95, 
    264.05, 264.05, 264.35, 264.05, 264.35, 264.65, 264.75, 264.75, 264.95, 
    265.05, 265.05, 264.75, 262.95, 262.35, 262.25, 261.55, 261.85, 263.65, 
    264.45, 264.85, 264.95, 264.55, 264.25, 263.95, 263.75, 263.55, 263.45, 
    263.45, 263.05, 262.85, 262.45, 262.55, 262.25, 262.35, 261.75, 261.75, 
    261.85, 261.65, 261.65, 261.85, 261.25, 262.25, 261.85, 261.35, 260.95, 
    259.05, 259.05, 258.85, 258.75, 258.35, 257.85, 257.75, 257.25, 256.55, 
    255.85, 255.85, 256.15, 257.95, 258.35, 257.85, 258.25, 258.75, 257.55, 
    258.05, 258.55, 259.05, 258.75, 258.45, 258.15, 258.25, 258.15, 257.85, 
    257.65, 257.65, 257.35, 257.35, 257.35, 257.15, 257.35, 256.85, 256.55, 
    255.45, 255.25, 255.15, 254.85, 253.95, 253.65, 252.05, 250.25, 251.45, 
    250.95, 250.45, 250.35, 250.55, 248.95, 249.85, 248.75, 250.15, 248.65, 
    248.55, 248.45, 248.35, 248.65, 247.55, 248.45, 248.55, 248.35, 249.05, 
    248.15, 248.95, 249.75, 249.65, 249.85, 250.35, 251.15, 252.45, 252.15, 
    253.65, 254.35, 254.55, 254.65, 254.65, 254.85, 254.65, 254.85, 254.95, 
    254.75, 254.75, 254.25, 254.45, 254.35, 254.45, 254.85, 255.05, 254.45, 
    254.35, 254.25, 253.05, 251.85, 251.75, 250.65, 250.95, 249.75, 250.45, 
    251.15, 249.65, 250.55, 250.55, 249.95, 249.85, 249.85, 249.75, 250.95, 
    249.65, 251.15, 249.55, 251.15, 251.05, 251.15, 249.85, 249.75, 250.05, 
    250.45, 248.45, 251.05, 249.75, 249.35, 249.55, 251.15, 250.65, 248.75, 
    250.25, 249.25, 248.15, 250.35, 251.05, 250.25, 249.45, 249.25, 250.55, 
    249.05, 249.55, 249.45, 251.75, 251.15, 252.05, 251.45, 253.15, 252.65, 
    253.15, 255.75, 255.55, 255.85, 256.05, 256.15, 256.35, 256.85, 256.85, 
    256.65, 256.35, 256.15, 255.75, 254.75, 253.95, 251.35, 253.15, 252.85, 
    252.05, 252.45, 252.05, 251.55, 250.85, 250.65, 250.45, 250.15, 249.85, 
    250.35, 251.45, 250.85, 250.65, 249.85, 249.85, 250.45, 248.55, 249.25, 
    250.15, 249.75, 250.35, 250.65, 250.15, 250.35, 251.55, 250.35, 250.85, 
    252.85, 252.05, 252.45, 252.95, 253.85, 255.65, 257.15, 257.25, 257.05, 
    256.45, 256.35, 256.45, 256.65, 256.55, 256.55, 256.35, 256.15, 256.45, 
    255.95, 255.25, 255.45, 255.65, 255.35, 255.45, 254.85, 253.75, 251.15, 
    251.85, 252.95, 253.25, 251.95, 252.95, 251.75, 252.15, 252.55, 251.95, 
    251.35, 251.55, 250.55, 249.55, 250.85, 252.25, 252.25, 252.15, 252.85, 
    252.95, 253.75, 254.15, 254.55, 255.05, 255.35, 254.95, 253.65, 252.95, 
    254.85, 254.05, 254.45, 255.85, 255.45, 254.35, 255.15, 255.95, 256.35, 
    256.75, 256.55, 256.85, 256.65, 256.85, 256.85, 257.15, 258.65, 258.05, 
    258.25, 258.25, 258.25, 258.35, 258.45, 258.05, 258.25, 257.55, 257.55, 
    257.25, 257.35, 257.85, 257.95, 257.75, 258.05, 258.35, 256.95, 257.25, 
    258.35, 257.95, 257.55, 256.05, 255.45, 255.65, 254.95, 253.25, 253.95, 
    253.25, 252.55, 252.05, 250.45, 252.45, 250.75, 254.05, 253.05, 252.85, 
    252.55, 255.45, 254.55, 254.05, 253.85, 253.35, 253.35, 252.55, 252.45, 
    252.25, 250.55, 250.75, 250.95, 250.75, 250.55, 250.65, 250.05, 250.15, 
    248.55, 250.45, 251.85, 252.95, 254.45, 255.75, 255.95, 255.25, 256.55, 
    255.95, 255.65, 256.15, 256.55, 257.65, 260.15, 259.35, 258.55, 257.35, 
    256.45, 255.15, 253.05, 251.55, 250.35, 250.35, 250.45, 250.45, 250.65, 
    251.05, 251.15, 250.15, 249.95, 249.95, 250.85, 251.95, 251.95, 250.65, 
    251.75, 252.75, 252.75, 253.95, 253.95, 254.35, 254.15, 253.85, 254.25, 
    254.65, 254.45, 253.35, 253.85, 254.15, 254.35, 253.85, 253.55, 252.75, 
    252.95, 251.25, 251.55, 251.75, 251.95, 251.65, 251.55, 251.55, 252.35, 
    251.75, 250.65, 250.25, 250.95, 251.75, 252.55, 252.55, 252.75, 252.75, 
    252.95, 252.55, 252.95, 252.65, 251.85, 251.65, 250.75, 250.95, 250.95, 
    250.75, 249.75, 250.25, 250.85, 249.25, 250.65, 249.45, 248.75, 248.45, 
    250.25, 248.95, 249.75, 250.55, 249.45, 251.15, 249.25, 249.45, 251.05, 
    250.85, 249.85, 249.65, 250.55, 250.35, 250.05, 251.65, 251.35, 251.95, 
    252.15, 252.25, 251.85, 255.45, 252.45, 253.55, 254.05, 255.75, 257.25, 
    257.95, 258.45, 259.65, 260.45, 261.45, 261.45, 261.25, 261.45, 261.55, 
    260.15, 263.65, 263.65, 263.95, 262.75, 262.45, 262.35, 262.35, 262.05, 
    261.95, 258.75, 259.65, 261.75, 263.05, 262.75, 259.95, 261.95, 261.15, 
    260.75, 259.85, 259.25, 259.15, 259.15, 259.05, 258.65, 257.75, 257.55, 
    257.65, 257.35, 256.45, 255.35, 255.25, 255.75, 253.35, 253.85, 252.85, 
    251.55, 250.75, 250.45, 250.35, 250.55, 250.85, 251.15, 251.65, 252.15, 
    252.35, 251.25, 251.55, 252.55, 252.75, 252.35, 251.85, 252.95, 256.95, 
    255.25, 256.15, 258.25, 258.65, 259.05, 259.25, 259.25, 258.95, 259.15, 
    258.85, 258.55, 257.75, 257.95, 258.95, 257.85, 256.75, 256.15, 255.35, 
    256.45, 256.15, 256.05, 257.15, 256.65, 255.35, 256.15, 256.25, 257.05, 
    256.55, 255.65, 255.55, 255.65, 255.85, 255.95, 256.45, 255.65, 255.55, 
    255.35, 256.55, 256.95, 256.65, 257.55, 257.35, 257.45, 257.45, 257.65, 
    257.25, 257.55, 258.45, 258.85, 258.75, 258.95, 259.55, 259.35, 259.15, 
    258.15, 257.35, 257.45, 257.75, 257.45, 255.95, 255.35, 256.95, 256.05, 
    255.35, 256.05, 256.15, 255.65, 255.65, 255.95, 255.55, 255.75, 255.45, 
    254.45, 254.65, 256.05, 255.25, 253.95, 254.85, 256.15, 255.05, 255.75, 
    257.15, 257.05, 257.35, 257.85, 259.35, 258.25, 259.05, 258.85, 259.55, 
    257.75, 258.75, 259.05, 259.45, 258.95, 259.45, 257.85, 258.25, 258.65, 
    258.25, 257.45, 256.75, 256.05, 256.25, 259.15, 258.35, 257.55, 258.55, 
    260.45, 260.85, 261.45, 260.95, 261.25, 261.25, 260.25, 260.85, 258.95, 
    261.75, 261.25, 261.15, 262.05, 263.15, 263.65, 265.75, 263.15, 263.65, 
    265.35, 263.45, 263.25, 263.45, 264.25, 263.55, 264.15, 266.05, 264.75, 
    266.25, 265.45, 264.25, 265.25, 263.05, 265.35, 264.55, 263.15, 267.05, 
    266.55, 266.25, 265.45, 264.75, 267.25, 267.05, 266.95, 267.05, 267.45, 
    266.35, 266.85, 266.85, 266.65, 267.45, 266.85, 267.55, 265.85, 265.55, 
    265.45, 264.65, 264.45, 264.95, 263.75, 264.45, 264.85, 264.65, 262.95, 
    262.35, 261.95, 261.55, 261.15, 260.55, 260.55, 261.15, 261.05, 261.45, 
    260.95, 261.35, 262.05, 262.35, 264.05, 262.95, 262.95, 260.45, 260.35, 
    259.45, 259.45, 259.45, 259.05, 259.75, 259.35, 259.45, 259.25, 259.65, 
    256.75, 258.25, 257.85, 259.55, 258.85, 259.05, 258.75, 261.25, 259.35, 
    260.45, 260.55, 261.05, 260.25, 258.35, 260.05, 259.45, 259.85, 260.15, 
    257.35, 258.75, 257.75, 258.75, 258.75, 258.75, 258.65, 256.25, 257.75, 
    258.65, 258.05, 258.85, 258.65, 260.65, 258.75, 260.65, 262.75, 259.95, 
    260.05, 260.25, 259.95, 259.85, 257.25, 257.65, 258.45, 258.55, 257.95, 
    258.85, 258.35, 258.35, 258.55, 258.95, 260.65, 258.25, 259.55, 259.75, 
    259.15, 260.25, 260.45, 261.95, 261.55, 262.35, 261.95, 261.15, 263.25, 
    260.65, 262.65, 263.45, 262.05, 261.55, 262.35, 261.45, 261.25, 262.05, 
    262.45, 266.05, 265.85, 265.85, 264.85, 265.55, 265.15, 265.15, 264.95, 
    264.05, 263.85, 263.85, 263.85, 262.65, 262.75, 262.75, 262.35, 261.95, 
    261.55, 261.05, 259.95, 258.55, 260.05, 260.05, 259.95, 259.75, 259.45, 
    258.75, 257.45, 257.35, 258.55, 257.45, 257.25, 258.25, 257.85, 256.65, 
    257.75, 256.45, 255.35, 255.45, 254.95, 254.55, 254.15, 253.15, 252.75, 
    251.75, 251.25, _, 250.85, 251.15, 251.75, 252.05, 253.05, 252.95, 
    253.15, 253.55, 253.65, 255.15, 254.75, 256.45, 255.25, 254.85, 254.45, 
    254.35, 252.05, 251.55, 252.05, 252.45, 251.35, 253.45, 254.05, 254.95, 
    255.65, 254.45, 254.55, 255.45, 256.45, 257.15, 257.45, 257.95, 258.15, 
    259.45, 258.75, 259.75, 258.85, 259.15, 258.55, 258.95, 257.85, 257.75, 
    258.25, 257.75, 257.15, 257.95, 259.35, 262.15, 264.65, 265.45, 265.85, 
    267.05, 266.45, 266.25, 266.75, 267.75, 268.55, 268.75, 268.35, 269.05, 
    268.55, 269.55, 268.75, 268.35, 269.35, 268.95, 269.55, 270.15, 269.75, 
    270.65, 270.25, 270.95, 271.45, 271.25, 270.95, 271.05, 271.45, 271.75, 
    271.15, 271.35, 271.15, 269.85, 269.65, 269.65, 269.55, 268.65, 268.75, 
    268.75, 267.85, 267.65, 265.75, 264.25, 264.25, 263.25, 263.45, 262.65, 
    262.25, 261.25, 261.75, 262.05, 261.65, 261.85, 261.65, 262.45, 262.05, 
    261.45, 260.95, 262.65, 261.05, 261.85, 261.35, 260.35, 260.55, 260.05, 
    260.05, 259.55, 259.75, 261.35, 261.65, 261.05, 260.35, 259.25, 260.25, 
    261.05, 260.75, 260.05, 261.35, 261.65, 261.45, 263.75, 265.25, 265.25, 
    265.55, 265.25, 264.35, 263.95, 262.95, 261.25, 260.05, 260.05, 259.75, 
    260.75, 261.65, 262.25, 262.15, 261.15, 259.85, 258.65, 260.45, 262.05, 
    262.05, 261.55, 261.85, 262.05, 262.65, 262.35, 261.75, 261.15, 260.45, 
    258.55, 257.55, 258.05, 257.95, 256.15, 256.35, 257.65, 258.05, 255.55, 
    255.95, 255.85, 257.25, 256.15, 256.85, 258.15, 258.35, 260.45, 259.75, 
    260.45, 262.65, 260.95, 260.85, 260.15, 260.05, 259.35, 258.45, 258.25, 
    258.85, 259.55, 257.85, 258.05, 257.95, 258.35, 258.65, 258.45, 258.55, 
    259.55, 259.15, 258.55, 261.55, 260.75, 262.95, 262.15, 263.05, 264.35, 
    263.25, 262.45, 261.55, 262.35, 261.05, 261.15, 260.35, 259.65, 262.55, 
    263.05, 262.15, 262.65, 261.65, 259.85, 259.35, 260.65, 262.05, 263.05, 
    265.05, 264.15, 262.95, 265.45, 265.05, 263.05, 264.35, 264.35, 262.15, 
    262.65, 261.45, 259.45, 261.35, 258.95, 259.25, 260.45, 259.35, 261.75, 
    260.95, 262.75, 262.75, 262.35, 262.65, 262.25, 262.85, 265.05, 266.05, 
    266.55, 266.55, 266.35, 265.25, 266.75, 266.95, 266.95, 267.85, 267.35, 
    266.45, 267.05, 266.75, 266.95, 266.55, 266.35, 266.25, 266.05, 264.75, 
    264.95, 265.15, 265.05, 264.55, 264.15, 264.65, 265.35, 265.15, 264.85, 
    263.95, 262.85, 262.65, 260.95, 260.25, 259.85, 259.05, 258.75, 258.55, 
    258.35, 258.05, 257.95, 257.95, 257.35, 259.35, 259.85, 259.95, 260.35, 
    260.65, 260.55, 260.85, 261.05, 261.25, 261.05, 260.75, 260.65, 260.35, 
    259.95, 259.55, 258.55, 257.85, 257.35, 257.55, 257.35, 256.95, 256.45, 
    255.95, 256.05, 255.95, 255.75, 255.85, 255.65, 256.05, 256.65, 257.25, 
    256.85, 257.15, 257.15, 257.05, 256.95, 256.15, 257.25, 256.45, 256.05, 
    255.25, 255.65, 256.45, 257.45, 257.55, 257.75, 257.85, 256.85, 257.15, 
    257.15, 257.25, 257.65, 258.55, 258.75, 259.15, 258.95, 258.95, 259.45, 
    258.75, 258.65, 257.75, 257.75, 257.35, 256.75, 256.35, 256.25, 255.45, 
    254.75, 254.05, 254.35, 253.85, 253.05, 252.75, 253.25, 253.55, 255.05, 
    255.35, 256.75, 255.75, 256.05, 255.85, 255.95, 255.85, 256.05, 255.85, 
    254.95, 255.35, 253.25, 253.85, 253.25, 253.25, 252.85, 253.65, 253.55, 
    253.45, 253.25, 253.45, 252.25, 254.75, 255.05, 256.95, 257.85, 259.55, 
    259.05, 258.65, 259.75, 259.85, 259.95, 258.25, 258.65, 257.95, 258.95, 
    258.15, 257.85, 259.45, 260.85, 260.15, 257.65, 257.05, 257.25, 257.55, 
    257.95, 259.35, 260.05, 261.05, 261.75, 262.35, 262.35, 263.05, 263.15, 
    261.35, 261.85, 260.45, 259.05, 258.25, 256.75, 256.05, 257.05, 257.15, 
    257.15, 256.15, 255.45, 255.65, 254.95, 255.95, 255.65, 258.15, 259.65, 
    258.85, 261.35, 261.65, 261.55, 262.35, 262.85, 261.95, 262.45, 262.15, 
    260.45, 260.25, 258.85, 259.15, 258.85, 258.25, 257.25, 256.25, 256.05, 
    257.05, 257.95, 257.05, 257.75, 258.85, 259.85, 262.25, 261.25, 262.35, 
    263.45, 263.25, 261.85, 264.65, 263.65, 262.75, 262.15, 261.45, 260.45, 
    259.55, 259.05, 259.75, 257.65, 258.65, 257.75, 258.45, 257.55, 257.55, 
    258.35, 260.55, 261.35, 260.95, 262.25, 261.75, 262.65, 261.35, 261.85, 
    263.65, 262.35, 263.45, 262.35, 260.95, 259.35, 258.45, 258.75, 258.55, 
    258.35, 258.45, 257.75, 256.95, 256.45, 258.15, 257.35, 259.05, 260.35, 
    261.05, 261.35, 261.75, 263.35, 261.55, 261.45, 262.25, 262.35, 259.65, 
    261.35, 261.05, 259.85, 258.65, 259.35, 260.05, 257.95, 257.85, 259.75, 
    257.75, 256.85, 258.05, 260.45, 260.65, 262.75, 261.85, 263.35, 263.45, 
    265.75, 264.35, 264.95, 264.15, 264.65, 264.05, 263.85, 262.85, 262.55, 
    260.45, 261.95, 259.25, 259.55, 259.25, 259.25, 259.65, 261.15, 261.55, 
    262.85, 265.65, 265.25, 266.35, 266.25, 266.55, 266.75, 266.95, 266.25, 
    266.55, 265.75, 265.15, 264.45, 263.65, 262.85, 261.85, 261.65, 261.15, 
    260.75, 260.05, 260.05, 259.45, 259.25, 259.35, 259.45, 260.85, 261.05, 
    261.35, 262.05, 261.05, 261.35, 262.15, 261.85, 260.35, 260.95, 260.65, 
    259.85, 258.75, 256.75, 256.05, 256.45, 256.85, 254.25, 256.35, 255.65, 
    255.45, 256.35, 257.85, 257.75, 258.65, 259.55, 262.25, 261.55, 264.45, 
    261.65, 262.75, 262.75, 261.85, 261.95, 261.55, 261.85, 261.25, 260.15, 
    259.05, 258.55, 258.45, 258.35, 258.45, 258.45, 258.35, 257.95, 258.15, 
    259.85, 261.35, 262.95, 264.55, 264.95, 266.35, 264.65, 267.85, 264.95, 
    264.75, 265.45, 264.65, 263.65, 263.15, 264.45, 264.15, 263.85, 264.15, 
    264.85, 264.25, 264.05, 263.55, 264.05, 264.15, 264.55, 266.45, 267.65, 
    269.25, 268.05, 270.15, 268.25, 268.15, 269.35, 267.25, 266.85, 267.85, 
    269.85, 268.95, 270.25, 271.05, 270.95, 272.05, 272.65, 273.05, 273.25, 
    273.05, 274.05, 275.35, 275.05, 275.25, 275.55, 276.05, 277.45, 277.35, 
    277.95, 278.05, 276.75, 275.65, 275.85, 275.25, 274.15, 275.05, 273.75, 
    273.55, 274.05, 274.25, 274.55, 276.05, 274.75, 274.35, 274.65, 275.05, 
    275.15, 275.15, 275.15, 275.15, 275.15, 276.05, 276.15, 275.95, 275.65, 
    275.05, 276.15, 275.95, 274.35, 276.65, 274.05, _, 274.35, 274.75, 
    274.55, 274.85, 273.55, 274.25, 275.85, 275.55, 275.75, 275.15, 275.25, 
    275.35, 275.25, 275.25, 274.95, 274.75, 274.45, 274.35, 273.95, 273.35, 
    273.45, 273.55, 273.75, 273.85, 273.45, 273.45, 273.25, 273.15, 273.45, 
    272.95, 273.45, 273.05, 273.05, 273.25, 274.25, 274.45, 274.45, 275.45, 
    274.75, 275.45, 275.15, 274.55, 274.15, 273.35, 273.45, 272.95, 272.55, 
    271.85, 271.85, 271.55, 271.45, 271.45, 271.15, 271.05, 271.05, 271.05, 
    271.15, 271.05, 271.95, 272.65, 271.95, 272.15, 272.65, 272.45, 270.95, 
    271.35, 271.15, 270.95, 270.35, 269.85, 269.55, 269.35, 268.75, 268.25, 
    268.25, 267.85, 267.65, 267.95, 267.75, 267.65, 267.75, 268.35, 268.85, 
    268.45, 269.25, 268.75, 269.45, 268.75, 269.05, 268.55, 268.95, 267.65, 
    267.95, 267.25, 266.65, 266.25, 265.85, 265.55, 265.65, 265.75, 265.45, 
    265.05, 264.95, 265.65, 266.65, 267.05, 267.75, 268.15, 269.55, 271.45, 
    271.95, 271.95, 271.15, 271.75, 270.75, 270.45, 270.75, 269.95, 270.25, 
    270.55, 270.25, 269.25, 269.75, 269.95, 269.15, 268.75, 268.55, 268.55, 
    268.65, 270.05, 270.65, 270.55, 269.65, 268.65, 268.05, 269.55, 269.25, 
    268.75, 268.45, 268.25, 268.95, 267.85, 267.05, 265.45, 266.15, 266.05, 
    264.15, 263.45, 264.35, 263.85, 264.55, 265.05, 266.35, 268.15, 269.95, 
    270.25, 269.05, 269.55, 272.75, 268.65, 269.25, 271.05, 269.95, 270.35, 
    269.65, 269.85, 269.85, 269.95, 271.95, 272.35, 272.55, 272.75, 272.55, 
    273.05, 273.15, 272.95, 272.95, 273.65, 274.25, 274.55, 273.65, 274.55, 
    273.35, 274.25, 273.65, 273.75, 272.65, 273.05, 273.35, 272.55, 270.95, 
    269.05, 268.75, 267.15, 265.95, 267.35, 265.55, 265.15, 265.15, 266.85, 
    266.85, 267.85, 269.65, 268.95, 269.35, 271.75, 271.85, 271.45, 274.75, 
    272.25, 270.55, 270.15, 270.25, 269.75, 268.15, 265.35, 265.25, 263.85, 
    263.15, 263.95, 263.65, 263.85, 264.15, 266.15, 265.25, 267.55, 269.25, 
    267.75, 271.95, 268.65, 269.05, 267.95, 269.15, 268.55, 268.05, 267.95, 
    268.25, 267.75, 267.45, 266.95, 266.35, 265.95, 265.35, 264.65, 264.05, 
    263.65, 263.45, 263.35, 263.75, 263.85, 263.75, 264.75, 264.85, 267.75, 
    266.05, 267.35, 267.45, 267.55, 268.15, 266.75, 266.75, 266.75, 266.95, 
    266.45, 266.65, 265.95, 266.15, 266.75, 267.35, 268.35, 269.25, 269.15, 
    269.25, 269.35, 269.45, 270.15, 270.65, 270.95, 271.45, 271.15, 270.75, 
    270.55, 270.55, 270.35, 269.65, 270.65, 270.15, 268.75, 267.55, 267.05, 
    268.15, 267.85, 267.85, 267.65, 266.95, 266.85, 267.25, 268.15, 268.75, 
    267.75, 267.65, 268.45, 268.05, 268.75, 267.85, 268.25, 268.45, 267.95, 
    266.55, 267.25, 266.55, 264.35, 264.15, 262.65, 263.35, 261.05, 263.45, 
    261.75, 263.45, 263.25, 264.75, 266.55, 266.15, 268.45, 270.35, 269.75, 
    274.25, 272.05, 271.45, 271.45, 272.45, 272.85, 272.15, 271.45, 272.15, 
    272.05, 271.85, 271.45, 270.45, 270.25, 268.55, 270.25, 270.45, 270.85, 
    269.85, 270.45, 272.05, 274.55, 272.85, 272.05, 272.15, 272.75, 272.55, 
    272.95, 274.05, 272.05, 272.45, 270.95, 270.35, 270.25, 269.85, 269.45, 
    269.35, 269.05, 269.15, 269.25, 269.45, 268.15, 268.05, 269.35, 270.45, 
    270.25, 269.65, 269.55, 269.65, 269.75, 270.05, 270.25, 270.35, 270.95, 
    271.15, 270.75, 269.75, 270.55, 270.95, 270.95, 270.85, 270.45, 270.15, 
    270.75, 271.45, 271.45, 271.75, 272.65, 272.85, 272.85, 272.45, 272.95, 
    273.45, 273.65, 273.45, 273.85, 274.15, 273.65, 273.25, 273.95, 273.45, 
    273.25, 272.95, 272.55, 272.25, 271.85, 271.95, 271.25, 271.75, 271.75, 
    271.95, 272.55, 272.75, 273.35, 276.05, 273.85, 274.05, 274.25, 272.55, 
    272.05, 272.45, 272.25, 271.55, 271.15, 270.75, 270.55, 270.35, 268.45, 
    267.35, 265.95, 265.95, 267.55, 267.35, 269.65, 268.35, 269.75, 270.65, 
    269.85, 270.95, 271.15, 271.15, 272.35, 272.85, 272.15, 271.35, 271.65, 
    270.85, 270.65, 269.85, 268.65, 267.45, 266.65, 266.55, 266.05, 266.05, 
    265.75, 265.65, 267.35, 267.95, 269.55, 270.55, 269.75, 269.95, 270.45, 
    270.35, 270.75, 270.55, 271.05, 270.55, 270.15, 270.15, 269.85, 269.65, 
    269.45, 269.25, 268.95, 268.65, 268.35, 268.25, 267.85, 268.15, 268.05, 
    268.35, 268.65, 268.85, 268.95, 269.65, 269.85, 269.55, 269.75, 270.15, 
    270.25, 270.05, 269.95, 269.85, 269.65, 269.75, 269.45, 269.15, 269.05, 
    269.05, 269.15, 268.95, 268.95, 269.15, 269.25, 269.15, 269.65, 269.55, 
    270.35, 270.05, 270.55, 270.35, 270.35, 270.75, 270.55, 270.65, 270.65, 
    270.15, 270.05, 269.95, 269.45, 269.45, 269.55, 269.35, 269.15, 269.15, 
    269.25, 269.35, 269.25, 269.25, 269.65, 269.65, 269.95, 270.05, 270.45, 
    270.85, 270.55, 270.85, 270.35, 271.15, 270.15, 270.35, 270.05, 270.05, 
    269.95, 269.75, 269.15, 268.95, 269.25, 269.25, 269.65, 270.15, 270.25, 
    270.65, 271.55, 270.05, 270.95, 272.05, 272.15, 270.85, 271.45, 271.85, 
    272.45, 272.55, 273.15, 273.45, 273.15, 274.05, 274.45, 274.65, 274.65, 
    275.35, 275.35, 276.05, 276.35, 274.85, 275.35, 276.05, 275.85, 275.25, 
    275.85, 275.45, 278.25, 277.05, 277.05, 277.05, 276.75, 276.55, 276.25, 
    275.45, 275.35, 274.95, 274.95, 274.15, 273.85, 273.65, 273.25, 272.85, 
    272.35, 273.15, 271.55, 272.15, 272.85, 273.65, 273.55, 274.55, 274.35, 
    274.35, 274.55, 274.85, 274.55, 274.75, 274.55, 274.15, 274.25, 273.95, 
    273.95, 273.85, 273.45, 273.55, 273.85, 273.75, 273.45, 273.65, 273.35, 
    274.05, 274.75, 274.75, 274.95, 275.15, 274.85, 275.15, 275.05, 275.25, 
    274.95, 274.75, 274.75, 274.55, 274.35, 274.25, 274.05, 273.85, 273.95, 
    273.95, 274.05, 274.25, 274.05, 274.35, 273.75, 273.45, 273.55, 274.05, 
    274.15, 274.85, 274.75, 275.15, 274.55, 275.25, 275.85, 276.15, 275.95, 
    275.05, 274.55, 274.35, 273.95, 273.65, 273.25, 272.55, 272.85, 272.65, 
    272.65, 272.25, 272.15, 272.65, 272.35, 272.55, 272.45, 272.65, 273.25, 
    273.15, 273.65, 273.55, 273.05, 272.95, 272.85, 272.85, 272.85, 272.25, 
    272.05, 271.95, 271.75, 271.85, 272.05, 271.65, 271.95, 272.95, 272.15, 
    272.65, 271.85, 270.95, 271.15, 271.65, 271.75, 272.05, 271.35, 271.95, 
    271.25, 271.25, 271.75, 272.05, 271.75, 271.35, 271.15, 271.05, 271.05, 
    271.45, 271.35, 271.35, 271.75, 271.85, 271.75, 271.85, 272.35, 272.35, 
    272.55, 272.65, 273.55, 274.65, 274.45, 274.25, 273.35, 274.65, 274.55, 
    274.65, 274.35, 273.85, 273.15, 272.55, 271.85, 271.05, 270.15, 269.55, 
    270.05, 270.25, 269.95, 269.95, 269.85, 270.15, 270.05, 269.95, 269.85, 
    269.75, 269.85, 269.45, 269.05, 268.65, 267.95, 268.35, 267.85, 268.05, 
    267.65, 267.05, 265.85, 266.05, 266.45, 265.05, 265.85, 265.35, 265.95, 
    267.95, 267.95, 268.45, 268.65, 269.85, 270.15, 269.95, 270.35, 271.05, 
    272.25, 270.25, 270.75, 270.75, 270.55, 270.15, 269.35, 268.45, 268.05, 
    268.45, 268.55, 268.55, 268.15, 270.15, 269.75, 270.65, 271.15, 271.25, 
    271.45, 271.05, 271.25, 272.05, 272.15, 272.45, 271.95, 272.05, 272.05, 
    272.05, 272.95, 271.95, 271.75, 271.45, 271.35, 270.85, 270.55, 271.45, 
    270.25, 271.45, 270.75, 270.75, 271.15, 272.45, 272.75, 273.25, 273.65, 
    273.55, 273.85, 274.55, 275.15, 274.75, 274.45, 273.75, 273.25, 272.75, 
    272.45, 272.65, 273.35, 273.85, 273.35, 273.05, 272.05, 272.85, 274.85, 
    274.75, 274.95, 274.95, 275.65, 275.85, 275.85, 275.45, 275.75, 275.95, 
    274.45, 274.95, 275.45, 274.65, 274.45, 274.35, 274.55, 274.35, 274.35, 
    273.65, 273.15, 273.15, 273.15, 273.45, 274.05, 273.55, 273.45, 273.55, 
    274.15, 274.15, 274.35, 274.65, 275.05, 275.55, 276.45, 275.85, 275.45, 
    275.85, 275.35, 275.75, 275.55, 275.85, 274.45, 274.95, 274.45, 274.65, 
    274.65, 274.85, 274.55, 274.75, 274.65, 274.95, 274.55, 275.35, 275.05, 
    275.25, 275.85, 274.65, 274.95, 274.45, 274.65, 274.25, 274.15, 274.25, 
    274.45, 274.55, 274.35, 274.35, 274.35, 274.25, 273.85, 273.95, 274.25, 
    274.35, 274.45, 275.05, 275.55, 275.85, 276.05, 276.25, 277.45, 277.25, 
    276.85, 276.75, 276.65, 276.75, 276.65, 276.35, 275.75, 274.75, 274.05, 
    273.95, 273.35, 272.95, 273.75, 274.95, 275.45, 275.45, 274.15, 275.35, 
    276.35, 276.35, 277.15, 276.35, 276.55, 277.35, 276.75, 277.15, 277.05, 
    276.95, 277.25, 276.65, 276.15, 275.65, 276.25, 276.25, 275.55, 276.45, 
    275.05, 276.95, 278.25, 277.85, 278.35, 278.15, 278.25, 277.75, 278.55, 
    278.35, 277.55, 277.75, 276.75, 277.25, 276.25, 276.95, 275.55, 278.65, 
    276.95, 275.35, 275.85, 277.05, 276.35, 275.95, 275.95, 276.35, 275.85, 
    276.15, 276.65, 276.45, 276.15, 275.35, 275.65, 275.75, 276.55, 276.45, 
    276.15, 276.25, 276.05, 276.15, 276.15, 275.95, 275.95, 275.65, 275.25, 
    274.95, 274.45, 274.65, 274.85, 274.95, 274.75, 277.45, 277.75, 278.15, 
    278.95, 278.25, 277.45, 278.25, 277.75, 278.55, 277.55, 277.45, 277.35, 
    277.35, 277.55, 277.65, 276.55, 276.85, 276.75, 276.25, 276.35, 276.35, 
    276.35, 276.55, 277.15, 276.65, 276.45, 276.15, 276.25, 276.65, 277.05, 
    277.75, 277.45, 277.45, 277.55, 277.15, 277.25, 276.65, 276.25, 276.15, 
    275.85, 275.35, 275.55, 274.55, 274.75, 275.05, 274.65, 274.85, 276.15, 
    276.25, 276.75, 277.25, 277.75, 278.15, 276.45, 276.25, 276.95, 275.85, 
    275.95, 275.45, 276.15, 275.55, 275.55, 275.35, 274.05, 273.35, 273.65, 
    273.15, 272.85, 272.75, 272.85, 273.45, 273.45, 273.75, 274.45, 274.55, 
    275.05, 275.65, 275.95, 276.35, 276.25, 276.55, 276.35, 276.25, 276.45, 
    276.55, 276.65, 276.65, 276.55, 276.05, 276.05, 275.95, 276.15, 276.15, 
    276.15, 276.05, 276.25, 276.15, 275.85, 275.55, 275.55, 275.95, 276.55, 
    275.95, 274.95, 274.95, 275.05, 275.05, 275.45, 275.65, 275.05, 274.55, 
    273.95, 272.65, 272.35, 271.45, 271.35, 271.55, 271.85, 272.35, 272.15, 
    272.25, 272.95, 273.25, 273.65, 273.65, 274.25, 274.85, 274.85, 274.65, 
    274.35, 274.25, 274.45, 274.35, 274.55, 274.35, 274.05, 274.25, 274.35, 
    273.65, 274.05, 274.05, 274.15, 274.55, 274.75, 274.75, 275.45, 276.35, 
    276.35, 275.75, 275.85, 275.85, 276.15, 276.45, 276.45, 277.15, 277.95, 
    278.25, 277.65, 276.95, 276.35, 276.05, 276.15, 275.85, 275.55, 275.65, 
    275.65, 275.85, 275.85, 276.15, 276.75, 276.75, 277.75, 278.05, 277.85, 
    277.65, 277.65, 277.85, 276.65, 275.65, 274.75, 274.45, 274.05, 274.45, 
    273.25, 272.75, 273.25, 272.55, 272.35, 272.75, 273.45, 273.65, 273.55, 
    273.75, 273.65, 274.15, 274.25, 275.35, 275.65, 276.35, 276.05, 275.25, 
    274.95, 275.25, 274.75, 274.55, 274.95, 274.55, 274.25, 274.45, 274.65, 
    274.65, 274.45, 274.55, 274.55, 274.75, 275.15, 275.75, 276.55, 276.85, 
    276.35, 276.75, 276.85, 276.65, 276.95, 277.05, 276.45, 276.55, 276.55, 
    276.75, 276.45, 276.15, 276.15, 275.95, 275.95, 275.65, 274.85, 274.75, 
    274.65, 274.55, 275.15, 274.75, 273.75, 273.35, 273.35, 273.95, 273.85, 
    273.65, 274.05, 273.35, 273.75, 273.45, 273.25, 273.35, 273.05, 273.05, 
    272.95, 272.95, 272.95, 272.45, 272.75, 272.45, 272.85, 272.85, 272.85, 
    273.15, 273.95, 273.55, 273.45, 273.35, 273.35, 273.15, 273.05, 273.35, 
    273.75, 273.65, 274.45, 275.05, 275.65, 275.25, 275.25, 275.55, 275.35, 
    275.15, 275.35, 275.35, 275.45, 275.95, 275.65, 275.75, 275.85, 276.35, 
    276.85, 276.95, 277.15, 277.15, 277.45, 277.65, 277.75, 277.45, 277.85, 
    277.15, 277.15, 277.05, 276.85, 276.65, 276.55, 276.25, 276.35, 276.55, 
    276.15, 276.45, 276.15, 276.55, 276.55, 275.55, 275.85, 275.85, 276.45, 
    276.45, 277.35, 276.55, 276.95, 276.85, 277.45, 277.75, 277.25, 277.45, 
    277.45, 277.35, 276.65, 276.75, 276.25, 276.25, 276.15, 276.25, 275.85, 
    275.85, 275.45, 275.55, 275.75, 276.25, 277.45, 279.95, 279.25, 279.45, 
    279.55, 280.05, 278.95, 279.75, 278.65, 279.35, 279.65, 279.35, 278.95, 
    278.65, 277.75, 278.55, 278.25, 277.75, 277.55, 277.65, 278.05, 279.75, 
    279.65, 279.65, 279.75, 280.65, 282.05, 281.55, 281.55, 281.55, 281.25, 
    280.55, 280.65, 280.75, 280.45, 280.35, 280.35, 280.35, 280.35, 280.35, 
    280.45, 280.75, 280.25, 279.85, 279.95, 280.85, 281.05, 280.15, 281.25, 
    281.45, 282.25, 282.45, 283.05, 282.95, 283.25, 281.95, 279.95, 279.65, 
    278.65, 279.15, 279.05, 278.85, 279.25, 279.55, 279.35, 279.45, 279.85, 
    279.95, 281.65, 281.15, 280.85, 281.55, 281.35, 281.45, 282.15, 281.45, 
    282.15, 281.45, 281.15, 281.35, 281.05, 281.45, 280.55, 280.65, 280.55, 
    280.95, 280.85, 279.85, 279.95, 279.25, 279.45, 280.25, 280.35, 280.95, 
    280.15, 279.85, 278.75, 279.65, 279.25, 280.65, 281.15, 280.95, 280.85, 
    280.55, 280.55, 280.55, 280.45, 280.35, 280.05, 279.55, 279.25, 279.05, 
    278.75, 278.15, 277.85, 278.95, 278.95, 278.35, 277.65, 278.45, 278.95, 
    279.15, 279.55, 279.05, 277.85, 278.15, 277.85, 277.75, 277.65, 277.55, 
    277.35, 277.25, 277.15, 277.15, 277.05, 276.95, 277.05, 277.25, 277.05, 
    277.25, 277.35, 277.45, 277.65, 277.55, 277.65, 277.45, 277.65, 277.55, 
    277.95, 277.85, 278.05, 278.15, 277.95, 277.75, 277.45, 277.25, 277.15, 
    277.25, 277.35, 277.15, 277.05, 277.45, 277.75, 277.75, 277.65, 278.35, 
    278.45, 277.85, 277.45, 277.35, 277.55, 277.55, 277.95, 278.35, 278.65, 
    278.95, 279.05, 278.55, 277.85, 277.75, 277.95, 278.05, 278.05, 277.85, 
    278.15, 277.85, 278.15, 278.05, 278.35, 278.65, 278.95, 279.25, 278.95, 
    278.55, 278.25, 278.55, 278.75, 278.95, 279.25, 279.15, 279.35, 279.25, 
    279.65, 279.65, 279.95, 279.95, 280.35, 278.95, 279.35, 280.15, 280.05, 
    279.95, 279.95, 279.75, 279.75, 280.75, 281.15, 280.65, 280.65, 280.85, 
    281.35, 280.85, 281.35, 282.05, 281.45, 282.45, 281.85, 282.55, 282.05, 
    280.75, 281.35, 280.75, 281.85, 281.25, 281.85, 281.25, 283.05, 282.15, 
    282.35, 284.25, 285.85, 286.05, 285.75, 284.45, 284.75, 284.45, 284.05, 
    284.35, 284.15, 282.45, 282.55, 281.85, 281.85, 281.25, 280.95, 280.95, 
    281.45, 281.55, 281.05, 281.05, 281.55, 282.15, 281.65, 281.05, 280.75, 
    281.05, 281.05, 281.65, 281.15, 280.95, 281.05, 281.65, 282.55, 281.95, 
    280.45, 280.05, 279.95, 279.75, 279.65, 280.05, 280.25, 279.65, 279.55, 
    280.35, 280.35, 280.45, 281.05, 281.35, 281.55, 281.45, 283.15, 281.65, 
    281.45, 281.45, 280.75, 280.25, 281.05, 281.15, 281.15, 279.85, 280.05, 
    281.05, 280.65, 280.55, 280.95, 280.95, 280.15, 279.95, 279.65, 280.55, 
    280.55, 281.25, 281.95, 282.15, 282.35, 283.25, 284.55, 284.25, 283.25, 
    282.55, 282.85, 282.35, 282.35, 282.35, 282.25, 282.45, 283.15, 281.05, 
    282.05, 281.65, 282.15, 282.35, 283.45, 285.25, 285.25, 284.55, 284.55, 
    285.45, 286.35, 286.15, 284.65, 284.45, 284.25, 283.85, 285.45, 283.45, 
    284.15, 282.55, 283.05, 283.35, 283.35, 283.05, 282.75, 283.25, 283.05, 
    283.05, 283.45, 283.65, 283.45, 284.05, 282.65, 283.05, 282.25, 282.05, 
    281.85, 281.45, 280.85, 280.05, 279.75, 279.75, 279.55, 279.25, 279.25, 
    279.15, 279.25, 279.05, 279.05, 279.05, 278.85, 279.05, 279.15, 279.45, 
    279.35, 279.55, 279.55, 279.75, 279.75, 279.55, 279.55, 279.65, 279.55, 
    279.55, 279.05, 279.85, 281.05, 280.55, 281.35, 281.95, 281.55, 282.65, 
    281.45, 281.25, 281.95, 281.75, 281.55, 281.45, 281.65, 281.55, 281.45, 
    280.95, 281.25, 283.35, 283.65, 283.45, 283.25, 284.15, 283.65, 283.25, 
    282.75, 281.75, 282.05, 281.05, 280.85, 280.65, 280.85, 280.35, 280.85, 
    280.35, 280.65, 282.75, 281.85, 282.65, 282.85, 282.95, 283.05, 282.85, 
    282.95, 282.85, 282.75, 282.15, 283.45, 283.05, 282.85, 282.65, 281.85, 
    281.55, 281.45, 280.65, 280.85, 280.75, 282.05, 282.25, 281.25, 281.65, 
    282.65, 282.75, 282.55, 282.95, 282.95, 283.35, 283.65, 282.35, 282.25, 
    281.95, 281.55, 281.25, 280.75, 280.75, 280.35, 280.15, 280.15, 280.35, 
    280.25, 279.85, 280.15, 280.45, 280.25, 280.25, 280.55, 280.75, 280.25, 
    280.05, 280.85, 281.35, 282.65, 282.85, 282.55, 281.75, 281.55, 281.25, 
    280.75, 280.25, 279.35, 278.55, 278.05, 277.55, 277.65, 277.95, 278.25, 
    278.25, 278.35, 278.15, 278.45, 278.45, 278.25, 277.65, 277.85, 277.85, 
    278.35, 279.05, 279.05, 278.85, 278.45, 278.65, 278.15, 278.35, 278.65, 
    279.15, 279.55, 279.95, 279.95, 280.65, 280.35, 280.35, 280.05, 279.95, 
    279.85, 280.25, 281.05, 280.25, 279.25, 279.75, 280.45, 281.25, 280.95, 
    280.95, 280.55, 279.55, 279.55, 279.15, 278.85, 278.65, 278.65, 278.45, 
    279.15, 279.15, 279.45, 279.85, 280.15, 280.65, 281.05, 281.25, 281.35, 
    281.55, 282.05, 282.15, 282.05, 281.95, 281.95, 282.45, 282.35, 282.25, 
    281.55, 281.05, 280.85, 280.35, 280.35, 279.95, 280.35, 280.55, 280.95, 
    280.75, 280.75, 282.05, 281.75, 282.65, 283.85, 283.95, 284.15, 284.35, 
    283.95, 284.05, 284.35, 284.95, 284.25, 283.55, 283.35, 282.75, 282.05, 
    281.55, 281.15, 281.35, 281.15, 282.85, 282.45, 282.65, 283.35, 283.95, 
    283.95, 283.95, 284.85, 284.15, 284.25, 284.35, 283.85, 284.05, 284.25, 
    283.85, 282.75, 282.35, 281.15, 281.35, 280.55, 280.35, 280.15, 278.85, 
    279.95, 279.85, 279.95, 278.85, 279.25, 279.35, 280.35, 279.35, 279.65, 
    278.25, 278.85, 278.75, 278.95, 278.65, 278.25, 278.15, 277.75, 277.45, 
    277.75, 277.85, 278.15, 277.95, 278.05, 277.95, 277.75, 278.25, 278.45, 
    278.55, 279.55, 280.15, 279.15, 279.05, 279.15, 278.65, 278.55, 278.45, 
    278.35, 278.35, 278.35, 279.35, 278.65, 278.65, 278.25, 278.35, 278.45, 
    278.05, 278.25, 278.55, 278.35, 278.75, 278.55, 278.35, 278.65, 279.45, 
    279.45, 279.55, 279.65, 280.15, 280.65, 280.15, 280.35, 280.75, 280.65, 
    280.35, 280.95, 281.55, 281.35, 279.65, 279.75, 280.25, 279.35, 279.85, 
    280.45, 281.55, 284.05, 281.75, 283.75, 283.45, 283.05, 282.55, 283.15, 
    283.15, 283.75, 283.65, 283.45, 283.25, 283.05, 283.25, 283.05, 282.55, 
    282.05, 281.15, 280.45, 280.65, 279.75, 279.25, 279.25, 280.65, 280.85, 
    280.75, 281.95, 283.05, 284.65, 284.75, 285.15, 285.25, 284.75, 284.05, 
    283.45, 283.05, 282.85, 283.55, 282.95, 282.45, 282.35, 282.35, 282.25, 
    282.15, 282.85, 282.25, 282.65, 282.75, 283.15, 283.35, 283.15, 284.65, 
    283.15, 281.85, 281.95, 282.45, 281.15, 279.85, 279.85, 279.65, 279.65, 
    279.55, 279.35, 279.35, 279.05, 278.95, 278.75, 278.65, 278.85, 278.85, 
    278.75, 278.75, 278.95, 279.75, 279.85, 279.95, 279.95, 279.35, 279.25, 
    279.55, 279.85, 280.05, 279.95, 280.05, 280.05, 279.55, 278.85, 279.15, 
    278.25, 277.95, 278.25, 278.25, 278.05, 278.05, 278.25, 278.25, 278.05, 
    278.05, 277.85, 278.65, 278.65, 278.85, 279.75, 279.95, 280.25, 279.75, 
    279.15, 279.35, 279.35, 278.95, 278.55, 277.75, 278.05, 278.05, 278.05, 
    277.75, 278.05, 278.15, 278.35, 278.05, 278.25, 278.55, 278.85, 279.05, 
    278.95, 279.05, 279.35, 279.25, 279.35, 279.45, 279.55, 279.45, 279.65, 
    279.55, 279.65, 279.65, 279.55, 279.65, 279.85, 279.35, 279.45, 279.25, 
    279.45, 279.55, 279.55, 279.65, 279.65, 280.15, 280.15, 280.05, 280.25, 
    279.95, 279.85, 280.05, 279.95, 279.85, 279.85, 280.35, 279.65, 279.55, 
    279.45, 279.35, 279.15, 279.35, 279.25, 279.25, 279.35, 279.45, 279.65, 
    280.25, 279.95, 280.35, 280.85, 281.05, 281.15, 281.35, 281.75, 281.85, 
    281.75, 281.65, 281.35, 280.45, 280.15, 280.45, 279.85, 279.95, 279.25, 
    279.45, 279.35, 279.25, 278.75, 278.75, 278.95, 279.05, 279.05, 279.05, 
    279.05, 279.25, 279.25, 279.15, 279.15, 279.45, 279.55, 279.65, 280.05, 
    280.15, 280.15, 279.85, 280.05, 280.15, 280.05, 280.25, 280.15, 280.05, 
    279.95, 279.85, 279.75, 279.75, 279.95, 280.05, 280.25, 280.65, 280.45, 
    281.25, 281.35, 281.55, 281.75, 281.55, 281.35, 282.45, 282.15, 281.45, 
    280.75, 280.35, 280.25, 279.85, 279.55, 279.35, 279.25, 279.05, 279.15, 
    279.55, 279.85, 279.85, 279.95, 280.05, 280.55, 280.45, 281.15, 281.45, 
    281.35, 281.65, 281.55, 281.15, 281.05, 280.45, 280.55, 280.15, 280.15, 
    280.05, 279.95, 279.95, 280.15, 280.65, 281.75, 281.45, 281.95, 282.55, 
    282.15, 281.75, 281.35, 281.55, 281.75, 281.95, 282.25, 281.85, 281.95, 
    282.35, 281.75, 281.45, 281.45, 281.05, 280.95, 280.75, 280.35, 280.05, 
    280.15, 280.45, 281.15, 281.55, 280.35, 280.65, 282.15, 282.85, 281.25, 
    284.15, 283.45, 284.25, 285.05, 285.05, 285.05, 284.85, 285.15, 285.15, 
    284.35, 283.15, 282.75, 282.75, 282.05, 282.25, 282.05, 281.65, 281.85, 
    281.55, 281.65, 281.05, 281.75, 281.55, 282.15, 282.05, 282.25, 282.25, 
    282.15, 282.05, 281.85, 281.35, 281.35, 281.05, 281.45, 281.95, 282.05, 
    282.05, 282.45, 282.55, 282.65, 282.55, 282.45, 281.95, 281.65, 282.25, 
    282.35, 282.45, 282.15, 282.85, 283.65, 283.75, 284.15, 283.65, 283.45, 
    282.95, 282.95, 282.65, 281.95, 281.35, 280.75, 280.25, 280.05, 280.15, 
    280.15, 279.85, 279.85, 280.25, 279.85, 280.05, 280.75, 280.85, 280.75, 
    280.25, 281.35, 280.85, 281.25, 280.75, 280.65, 280.65, 281.25, 281.05, 
    281.45, 280.85, 280.55, 280.45, 280.25, 280.25, 280.05, 280.35, 280.45, 
    280.75, 281.25, 281.65, 281.95, 282.45, 283.85, 282.85, 281.65, 281.75, 
    282.35, 282.45, 282.45, 281.85, 281.55, 281.65, 281.35, 280.95, 281.25, 
    280.75, 280.35, 280.35, 280.55, 280.25, 280.95, 280.95, 281.05, 281.05, 
    280.95, 280.95, 281.25, 280.95, 281.45, 281.65, 281.25, 282.65, 281.75, 
    281.35, 281.45, 281.25, 281.85, 281.75, 281.65, 281.85, 281.75, 281.55, 
    281.35, 280.55, 280.75, 280.85, 280.05, 279.95, 280.35, 280.45, 281.35, 
    281.35, 281.25, 281.25, 281.55, 281.55, 281.35, 281.05, 280.85, 280.55, 
    280.45, 280.65, 280.35, 280.35, 280.25, 280.35, 280.45, 280.55, 280.45, 
    280.05, 280.15, 280.35, 280.65, 280.55, 280.65, 282.05, 281.95, 282.55, 
    283.05, 282.75, 282.45, 282.75, 283.15, 283.55, 282.45, 282.25, 282.15, 
    281.55, 281.05, 281.55, 281.65, 282.15, 281.55, 282.15, 282.25, 282.05, 
    282.45, 281.95, 282.05, 282.55, 283.05, 282.95, 282.55, 282.75, 282.05, 
    281.75, 281.45, 281.05, 280.95, 280.85, 280.75, 280.45, 280.55, 280.75, 
    281.15, 280.55, 280.35, 280.35, 280.25, 280.15, 279.95, 279.95, 279.85, 
    280.05, 280.15, 279.75, 279.45, 279.45, 279.05, 278.05, 277.95, 277.55, 
    277.25, 276.95, 276.85, 276.85, 276.65, 276.95, 277.15, 277.25, 277.15, 
    276.95, 277.15, 277.65, 277.95, 278.75, 278.35, 278.85, 278.85, 278.65, 
    278.65, 278.55, 278.35, 278.15, 277.75, 277.75, 277.65, 277.15, 276.95, 
    277.25, 277.15, 276.95, 277.15, 277.45, 277.45, 277.45, 277.05, 277.65, 
    278.35, 278.35, 277.95, 277.85, 278.75, 279.35, 279.55, 278.15, 277.65, 
    278.45, 276.85, 276.25, 276.25, 275.45, 275.05, 274.95, 274.65, 273.25, 
    273.65, 273.85, 275.65, 275.25, 276.05, 276.25, 276.15, 275.85, 276.95, 
    276.45, 276.55, 276.65, 276.45, 276.55, 277.35, 276.65, 276.95, 276.85, 
    276.65, 276.45, 276.55, 276.55, 276.45, 276.55, 277.05, 277.55, 277.35, 
    277.45, 277.75, 277.55, 277.75, 277.75, 277.05, 276.85, 276.65, 277.05, 
    278.05, 277.95, 277.55, 277.05, 276.85, 276.55, 276.25, 276.25, 276.25, 
    276.25, 275.95, 275.95, 276.05, 275.65, 275.35, 275.35, 275.25, 274.75, 
    274.65, 274.25, 274.35, 274.45, 274.55, 274.55, 274.65, 275.65, 275.75, 
    275.15, 275.05, 275.05, 274.95, 274.95, 274.95, 275.05, 274.95, 275.05, 
    275.15, 274.95, 274.95, 274.95, 275.15, 275.05, 274.95, 274.45, 274.25, 
    274.35, 275.85, 276.55, 276.65, 277.25, 275.95, 276.15, 278.45, 279.45, 
    280.05, 279.45, 279.75, 279.45, 279.15, 278.95, 278.65, 278.85, 278.95, 
    279.05, 279.15, 279.45, 279.15, 278.45, 278.65, 278.75, 279.35, 279.45, 
    279.35, 279.45, 279.35, 279.85, 279.95, 279.75, 279.55, 278.85, 279.05, 
    278.95, 279.15, 279.55, 279.55, 279.55, 280.15, 280.05, 279.85, 280.15, 
    280.45, 280.65, 280.65, 280.85, 280.65, 280.95, 281.15, 280.85, 280.35, 
    280.75, 281.05, 280.75, 280.05, 280.55, 280.55, 279.55, 279.85, 280.15, 
    280.25, 280.55, 281.25, 281.35, 280.25, 280.55, 280.15, 281.15, 281.95, 
    284.45, 285.15, 283.55, 283.55, 284.25, 287.45, 283.35, 285.45, 284.05, 
    284.15, 284.15, 283.25, 283.55, 283.95, 284.25, 284.75, 283.95, 284.35, 
    283.55, 283.75, 283.65, 283.95, 282.95, 282.85, 282.75, 282.75, 282.25, 
    281.85, 282.45, 282.55, 282.55, 282.65, 282.05, 281.85, 281.35, 281.65, 
    280.55, 279.15, 279.25, 279.85, 279.85, 279.85, 280.05, 279.75, 281.05, 
    280.35, 282.55, 283.15, 282.85, 285.25, 286.75, 287.25, 285.15, 285.05, 
    285.35, 285.25, 285.15, 283.85, 282.85, 282.95, 282.35, 282.15, 282.05, 
    282.05, 281.65, 280.75, 280.85, 281.45, 281.75, 281.35, 281.45, 281.25, 
    281.65, 281.95, 282.15, 280.75, 280.65, 280.75, 280.85, 281.85, 281.75, 
    281.65, 281.25, 281.55, 281.25, 281.35, 281.35, 281.35, 280.55, 279.55, 
    280.65, 281.65, 281.25, 281.75, 282.05, 282.25, 281.65, 282.05, 284.15, 
    284.15, 284.15, 283.45, 282.45, 282.15, 282.15, 281.65, 281.75, 280.75, 
    280.25, 280.05, 279.95, 279.85, 279.85, 280.35, 280.45, 280.15, 280.65, 
    281.35, 281.95, 281.45, 281.55, 281.55, 281.55, 281.45, 281.15, 280.65, 
    280.65, 280.55, 280.35, 279.95, 280.15, 280.15, 279.75, 279.75, 279.45, 
    279.35, 279.05, 279.05, 280.05, 280.25, 281.25, 280.85, 280.05, 280.75, 
    281.55, 281.05, 280.35, 280.45, 280.35, 279.85, 279.55, 279.25, 278.85, 
    278.75, 278.95, 278.85, 278.45, 277.95, 277.55, 278.95, 277.55, 277.95, 
    278.85, 279.35, 280.35, 280.25, 280.65, 280.25, 280.25, 280.15, 280.65, 
    280.45, 280.65, 281.15, 280.45, 280.65, 279.95, 279.85, 279.75, 279.65, 
    279.35, 279.35, 279.35, 279.25, 279.15, 279.05, 279.05, 279.15, 279.25, 
    279.05, 279.25, 279.95, 280.45, 280.35, 280.05, 279.45, 279.95, 279.75, 
    279.45, 279.35, 279.45, 279.35, 279.55, 280.15, 280.25, 279.85, 279.25, 
    279.35, 280.35, 280.55, 279.35, 280.35, 280.95, 281.65, 282.75, 283.35, 
    283.45, 282.85, 283.35, 284.75, 285.65, 283.95, 283.95, 283.95, 284.05, 
    283.95, 284.35, 283.55, 283.75, 283.15, 282.15, 281.95, 281.35, 281.65, 
    281.15, 282.55, 282.45, 282.65, 282.75, 282.35, 282.05, 281.95, 282.15, 
    281.75, 281.45, 281.75, 281.55, 281.45, 281.55, 281.85, 281.65, 281.45, 
    281.25, 281.25, 280.55, 280.75, 280.35, 280.85, 280.35, 280.35, 280.65, 
    282.15, 281.75, 282.05, 281.65, 281.85, 281.65, 281.55, 281.65, 281.85, 
    281.75, 281.85, 281.45, 281.35, 280.95, 280.45, 281.45, 282.15, 281.85, 
    281.75, 281.45, 280.45, 280.95, 281.15, 281.75, 282.35, 281.25, 281.75, 
    282.15, 281.95, 281.55, 281.25, 281.05, 280.25, 280.35, 279.05, 278.85, 
    278.55, 278.15, 278.35, 278.55, 278.35, 277.95, 278.45, 277.75, 277.55, 
    277.55, 278.65, 278.85, 278.75, 279.15, 279.75, 279.65, 279.35, 279.55, 
    279.55, 278.75, 279.15, 278.55, 278.15, 277.15, 276.45, 276.75, 276.55, 
    276.45, 276.45, 276.05, 276.35, 276.15, 276.15, 276.25, 277.05, 276.85, 
    276.95, 277.35, 277.15, 277.15, 277.35, 277.75, 278.05, 278.15, 277.95, 
    277.65, 277.35, 276.75, 275.85, 275.75, 274.35, 274.25, 273.85, 274.15, 
    274.45, 274.65, 274.75, 274.85, 275.05, 275.45, 276.05, 276.45, 276.75, 
    276.95, 276.95, 276.65, 276.75, 276.65, 276.65, 276.65, 276.45, 276.25, 
    276.15, 275.95, 275.65, 275.45, 275.35, 275.05, 274.75, 274.65, 274.75, 
    274.85, 274.65, 274.45, 274.75, 275.05, 275.25, 275.25, 275.15, 275.15, 
    275.25, 275.65, 275.65, 275.65, 275.55, 275.15, 275.05, 274.65, 274.55, 
    274.45, 274.85, 274.65, 274.05, 274.35, 274.65, 275.15, 275.55, 276.25, 
    277.05, 276.95, 277.65, 277.95, 277.45, 278.25, 278.35, 278.25, 278.25, 
    278.55, 278.05, 278.25, 278.15, 278.95, 279.45, 282.15, 282.15, 281.95, 
    281.35, 280.75, 280.85, 280.25, 279.75, 281.45, 280.75, 281.15, 281.45, 
    281.85, 283.25, 283.65, 282.35, 282.25, 282.05, 281.95, 281.45, 280.95, 
    280.25, 280.75, 279.85, 280.65, 279.95, 279.65, 279.35, 279.25, 279.95, 
    279.15, 278.65, 278.05, 278.15, 278.55, 278.65, 278.55, 278.45, 280.15, 
    279.75, 278.05, 278.15, 277.95, 278.05, 277.85, 277.75, 277.55, 277.35, 
    277.25, 277.05, 277.15, 277.25, 277.05, 276.95, 277.35, 278.15, 278.55, 
    278.75, 279.05, 278.95, 279.15, 279.25, 279.35, 279.25, 279.05, 278.95, 
    278.65, 278.05, 277.85, 277.95, 278.05, 278.35, 278.55, 278.35, 278.05, 
    277.75, 278.15, 277.75, 277.65, 278.45, 278.25, 278.25, 278.05, 278.15, 
    278.35, 277.65, 277.85, 278.25, 277.55, 277.35, 277.15, 277.05, 276.85, 
    277.25, 277.05, 276.75, 276.25, 276.05, 274.45, 275.15, 275.15, 275.45, 
    275.55, 276.15, 276.65, 276.75, 276.85, 277.05, 277.45, 277.95, 278.45, 
    279.25, 279.25, 279.05, 278.75, 278.45, 278.35, 277.85, 277.85, 277.65, 
    277.55, 277.65, 277.45, 277.05, 276.75, 276.55, 276.35, 276.35, 276.45, 
    276.45, 276.55, 276.75, 276.95, 277.85, 277.35, 278.05, 277.85, 278.25, 
    277.95, 277.55, 277.55, 277.45, 277.05, 276.95, 276.55, 276.25, 276.15, 
    276.05, 275.95, 275.25, 275.15, 275.35, 275.95, 276.25, 276.95, 276.85, 
    276.65, 276.55, 276.35, 276.05, 275.65, 275.55, 275.55, 275.15, 275.25, 
    274.75, 274.75, 273.75, 273.35, 273.35, 273.45, 273.55, 273.65, 273.85, 
    274.25, 273.95, 274.45, 274.85, 275.15, 275.95, 276.55, 276.15, 275.65, 
    276.15, 275.55, 275.65, 275.55, 275.25, 274.95, 274.95, 275.15, 274.95, 
    274.15, 274.65, 274.65, 273.95, 273.85, 273.95, 274.15, 274.35, 274.85, 
    275.45, 276.65, 277.25, 277.35, 276.95, 277.15, 277.05, 276.65, 276.65, 
    276.65, 276.55, 276.45, 276.45, 276.45, 276.75, 276.65, 277.05, 277.55, 
    277.35, 276.55, 279.65, 279.05, 279.15, 279.25, 279.45, 279.85, 279.75, 
    279.55, 280.55, 280.75, 281.05, 281.15, 280.45, 280.95, 279.95, 279.65, 
    279.85, 279.85, 278.75, 278.55, 278.25, 278.45, 277.95, 277.75, 278.25, 
    278.05, 279.45, 279.65, 280.15, 280.55, 280.05, 279.55, 279.75, 279.65, 
    279.05, 279.15, 278.05, 277.75, 277.85, 277.65, 277.75, 277.85, 277.25, 
    277.05, 276.35, 276.65, 277.05, 277.05, 277.15, 276.25, 276.35, 276.25, 
    276.65, 277.55, 277.75, 278.15, 277.55, 278.35, 277.35, 277.35, 277.15, 
    276.55, 275.85, 274.75, 274.85, 274.65, 275.05, 273.85, 275.45, 274.05, 
    274.15, 273.95, 274.35, 274.65, 275.25, 276.25, 276.35, 277.05, 276.35, 
    275.85, 276.55, 277.45, 277.55, 276.95, 276.05, 274.75, 275.45, 275.25, 
    275.95, 275.05, 275.15, 276.15, 275.85, 274.05, 274.35, 274.85, 275.35, 
    275.05, 275.35, 275.65, 275.75, 275.85, 275.95, 276.05, 276.85, 277.15, 
    276.15, 277.15, 277.45, 277.15, 276.85, 276.45, 278.45, 278.25, 277.45, 
    277.65, 277.75, 277.35, 276.85, 276.75, 276.35, 276.15, 277.35, 278.75, 
    279.15, 279.45, 279.85, 278.75, 278.95, 278.95, 280.05, 279.15, 279.55, 
    276.65, 277.15, 276.75, 277.45, 276.75, 275.95, 277.95, 275.85, 276.75, 
    276.25, 275.25, 275.45, 277.45, 276.35, 277.15, 278.35, 278.35, 278.45, 
    278.55, 277.95, 280.15, 280.45, 278.75, 277.55, 278.75, 277.95, 279.25, 
    279.45, 276.25, 276.65, 278.75, 277.55, 277.35, 277.35, 277.15, 278.05, 
    278.85, 281.35, 280.35, 281.45, 282.95, 283.65, 283.05, 281.85, 281.85, 
    282.75, 283.85, 281.55, 282.15, 282.15, 281.95, 281.95, 281.65, 281.95, 
    283.15, 280.65, 280.45, 280.45, 280.05, 279.75, 281.65, 279.05, 278.95, 
    279.15, 281.25, 280.85, 280.35, 280.75, 280.75, 280.75, 280.75, 279.75, 
    278.95, 277.95, 277.95, 278.15, 278.35, 277.95, 277.85, 277.75, 277.85, 
    277.45, 276.95, 276.75, 276.65, 276.75, 276.45, 276.75, 276.75, 277.35, 
    277.25, 276.95, 277.85, 278.05, 278.35, 278.55, 278.55, 278.55, 277.55, 
    277.55, 278.05, 277.85, 277.25, 276.65, 276.25, 276.65, 276.65, 276.85, 
    276.45, 276.65, 275.75, 275.95, 276.25, 276.55, 276.75, 276.45, 275.65, 
    275.45, 274.95, 275.25, 274.65, 273.65, 274.35, 272.95, 273.45, 273.05, 
    273.25, 272.85, 272.55, 271.85, 272.15, 271.95, 272.15, 272.25, 272.45, 
    272.75, 272.55, 273.45, 273.55, 273.35, 273.45, 273.35, 272.95, 272.55, 
    272.45, 272.65, 272.35, 272.15, 271.75, 271.45, 271.65, 271.75, 271.35, 
    270.95, 270.65, 270.65, 270.65, 271.25, 271.15, 270.95, 270.55, 270.65, 
    270.55, 270.85, 269.85, 270.15, 269.85, 269.95, 269.45, 268.95, 269.15, 
    268.45, 268.05, 267.85, 268.35, 267.95, 267.85, 267.85, 266.85, 266.85, 
    267.05, 267.15, 268.15, 269.05, 268.95, 269.65, 270.35, 269.65, 269.15, 
    269.65, 269.15, 269.15, 268.25, 268.95, 268.95, 268.55, 269.15, 269.05, 
    269.85, 268.95, 269.35, 269.95, 269.95, 269.15, 270.05, 271.15, 271.15, 
    271.25, 271.55, 273.05, 272.75, 271.95, 271.75, 272.55, 272.65, 272.55, 
    272.55, 272.35, 272.05, 272.55, 273.05, 272.65, 272.55, 272.95, 273.35, 
    273.35, 272.95, 272.45, 272.05, 271.75, 272.45, 273.95, 275.05, 275.75, 
    274.05, 274.05, 273.85, 273.95, 273.75, 273.85, 273.95, 271.75, 272.35, 
    272.95, 272.35, 271.95, 272.65, 273.35, 273.75, 274.15, 274.45, 274.55, 
    274.55, 274.05, 273.95, 274.05, 274.55, 274.95, 275.85, 276.15, 277.25, 
    275.35, 276.25, 276.35, 276.45, 277.35, 276.05, 276.25, 275.95, 275.45, 
    275.45, 275.95, 276.65, 276.85, 277.35, 275.55, 275.35, 275.95, 275.95, 
    276.25, 276.65, 276.75, 278.05, 278.15, 277.85, 277.55, 278.15, 276.35, 
    276.15, 277.65, 276.25, 276.35, 278.75, 278.55, 278.25, 277.75, 277.15, 
    276.65, 276.65, 276.25, 275.55, 276.25, 276.35, 275.65, 275.85, 275.75, 
    276.15, 275.65, 275.35, 274.75, 274.95, 275.15, 274.85, 274.55, 274.45, 
    274.65, 274.45, 274.35, 273.95, 274.35, 274.45, 273.95, 274.05, 273.35, 
    274.55, 273.85, 273.75, 273.65, 274.05, 273.85, 273.65, 273.65, 273.45, 
    273.35, 273.95, 272.05, 272.75, 272.55, 271.65, 271.65, 271.85, 271.85, 
    271.55, 271.05, 270.65, 270.95, 271.05, 271.75, 270.95, 271.05, 271.85, 
    271.55, 271.25, 271.55, 271.75, 272.25, 272.65, 272.05, 272.35, 272.75, 
    272.95, 273.35, 273.45, 273.45, 273.25, 271.15, 272.05, 270.25, 270.85, 
    270.05, 269.35, 270.85, 269.65, 268.75, 268.55, 268.75, 269.25, 268.95, 
    269.05, 269.75, 269.05, 270.15, 269.95, 269.75, 268.95, 269.25, 269.45, 
    269.05, 271.85, 267.75, 270.85, 269.85, 271.45, 271.05, 271.15, 271.45, 
    271.25, 270.65, 270.95, 271.35, 270.85, 271.75, 270.55, 270.75, 269.85, 
    269.25, 269.15, 267.75, 268.35, 269.05, 268.55, 271.25, 271.15, 272.75, 
    273.05, 273.15, 273.15, 272.75, 272.85, 272.95, 272.95, 272.95, 273.35, 
    273.05, 272.85, 272.95, 273.05, 272.25, 271.75, 271.45, 271.45, 271.55, 
    271.55, 271.55, 271.65, 271.75, 271.35, 271.55, 271.55, 271.25, 271.15, 
    271.15, 271.25, 270.95, 270.95, 271.05, 270.95, 270.85, 270.75, 271.55, 
    271.65, 271.35, 271.65, 271.35, 271.05, 271.25, 271.25, 271.25, 271.25, 
    271.45, 271.35, 271.15, 271.35, 272.05, 271.25, 271.45, 271.45, 271.75, 
    271.65, 271.55, 271.95, 271.95, 271.85, 272.25, 272.25, 271.65, 272.35, 
    272.45, 272.35, 272.75, 272.85, 272.75, 272.85, 272.95, 272.95, 273.15, 
    273.85, 273.45, 273.35, 273.55, 273.45, 273.55, 273.45, 273.85, 273.65, 
    273.05, 272.45, 272.75, 273.15, 273.15, 272.95, 273.15, 273.65, 273.75, 
    274.75, 274.95, 275.05, 275.25, 275.35, 275.55, 275.25, 275.05, 275.25, 
    275.15, 274.05, 272.95, 271.95, 270.95, 270.65, 270.75, 271.35, 271.85, 
    273.65, 272.95, 272.15, 271.35, 270.65, 269.95, 269.45, 269.35, 270.05, 
    270.35, 270.65, 268.85, 269.95, 270.85, 271.75, 272.65, 272.25, 271.55, 
    270.65, 270.45, 269.95, 268.95, 268.35, 267.75, 267.35, 266.95, 266.15, 
    265.55, 265.35, 264.75, 264.15, 264.55, 264.75, 264.45, 264.65, 263.65, 
    262.95, 262.85, 262.95, 262.25, 263.05, 262.55, 262.55, 262.85, 260.95, 
    260.75, 261.15, 262.05, 261.95, 262.55, 262.85, 263.55, 264.25, 264.45, 
    264.35, 266.45, 265.85, 265.75, 266.15, 265.75, 269.55, 268.15, 268.15, 
    267.45, 266.95, 267.55, 267.85, 267.95, 267.35, 266.85, 266.55, 268.15, 
    268.15, 268.55, 268.85, 268.85, 268.45, 269.15, 269.35, 269.45, 269.05, 
    269.05, 268.75, 268.65, 267.75, 267.25, 267.85, 267.25, 267.45, 268.75, 
    268.65, 270.35, 270.45, 271.95, 271.75, 271.45, 271.15, 270.85, 270.75, 
    270.95, 271.15, 271.15, 270.85, 270.65, 270.55, 270.05, 269.65, 270.25, 
    270.25, 269.95, 269.95, 270.05, 269.95, 269.65, 269.75, 269.75, 269.65, 
    268.45, 267.05, 265.85, 265.25, 266.05, 264.85, 265.25, 264.25, 263.95, 
    265.95, 265.45, 265.25, 265.25, 265.85, 266.65, 267.45, 266.85, 265.45, 
    264.05, 264.25, 265.25, 265.45, 264.95, 265.15, 264.15, 264.55, 264.85, 
    265.35, 265.35, 266.35, 266.05, 265.05, 265.55, 266.25, 266.85, 266.95, 
    265.15, 264.75, 264.85, 265.25, 264.45, 264.95, 264.75, 266.55, 266.55, 
    266.35, 266.25, 265.95, 265.75, 265.45, 265.45, 265.65, 265.75, 265.75, 
    265.85, 265.85, 265.25, 265.35, 265.55, 265.75, 265.75, 266.25, 266.55, 
    266.45, 266.55, 266.85, 266.85, 267.05, 267.05, 267.45, 267.45, 267.85, 
    267.85, 268.35, 268.05, 268.65, 267.75, 268.25, 267.15, 268.55, 268.55, 
    268.65, 267.05, 266.15, 265.15, 265.55, 264.65, 264.95, 264.25, 265.85, 
    265.95, 265.55, 265.35, 264.75, 264.05, 263.95, 264.55, 264.95, 264.25, 
    264.05, 265.05, 265.15, 265.65, 265.55, 265.85, 265.35, 265.45, 265.45, 
    266.35, 266.45, 266.25, 266.35, 266.55, 266.25, 266.25, 266.35, 265.25, 
    264.95, 264.95, 264.95, 265.15, 265.05, 265.05, 264.05, 263.05, 263.45, 
    263.25, 263.75, 262.95, 263.85, 264.15, 264.75, 264.95, 265.05, 265.25, 
    265.35, 265.45, 265.55, 265.75, 265.85, 266.05, 266.05, 264.95, 264.55, 
    264.75, 265.85, 266.85, 265.65, 265.95, 264.85, 264.95, 267.25, 266.85, 
    266.55, 265.45, 266.05, 265.75, 266.35, 265.05, 265.25, 265.65, 265.45, 
    265.55, 265.95, 265.85, 265.55, 265.25, 265.35, 265.35, 266.05, 264.35, 
    263.55, 265.65, 266.55, 264.95, 265.75, 264.65, 265.85, 263.15, 263.75, 
    265.05, 264.35, 264.75, 264.25, 264.35, 265.25, 265.85, 265.35, 265.45, 
    267.05, 267.35, 267.15, 266.95, 266.85, 266.75, 266.55, 266.25, 265.45, 
    264.45, 263.95, 261.65, 262.15, 261.45, 261.35, 262.35, 261.15, 260.95, 
    260.95, 261.95, 261.65, 261.25, 262.35, 262.25, 261.45, 262.05, 262.45, 
    261.75, 261.25, 261.55, 262.75, 261.95, 262.05, 263.95, 263.75, 263.05, 
    262.55, 262.45, 262.35, 262.35, 261.65, 262.15, 261.55, 261.45, 261.85, 
    261.95, 263.25, 262.85, 262.65, 262.55, 262.55, 260.95, 261.25, 260.35, 
    260.25, 260.55, 261.25, 261.05, 260.45, 260.05, 259.75, 259.65, 259.95, 
    259.95, 260.65, 260.85, 260.75, 261.25, 261.65, 261.35, 259.85, 259.85, 
    260.45, 259.95, 260.55, 260.65, 261.45, 261.35, 261.05, 261.65, 261.35, 
    262.65, 261.55, 262.05, 262.25, 262.75, 263.05, 263.15, 263.45, 263.95, 
    264.25, 264.25, 264.45, 264.65, 264.95, 264.85, 265.25, 265.25, 265.45, 
    265.55, 265.65, 266.05, 266.45, 266.25, 266.35, 266.95, 266.75, 267.25, 
    266.85, 267.15, 266.85, 267.45, 267.45, 267.15, 267.35, 267.35, 267.35, 
    267.35, 267.65, 267.75, 267.75, 267.75, 267.85, 267.85, 267.65, 268.05, 
    267.95, 268.45, 268.05, 268.55, 268.35, 268.45, 268.65, 268.65, 268.85, 
    269.15, 269.45, 269.45, 269.45, 269.65, 269.65, 269.85, 269.65, 269.85, 
    269.85, 269.65, 269.55, 269.65, 269.35, 269.15, 269.15, 269.05, 268.65, 
    268.35, 268.65, 268.55, 268.35, 268.45, 268.35, 268.15, 268.05, 267.95, 
    267.05, 266.35, 265.15, 266.35, 266.65, 265.85, 266.45, 266.45, 266.45, 
    266.45, 266.05, 265.15, 266.35, 266.75, 266.45, 264.45, 267.25, 266.45, 
    266.05, 265.05, 265.15, 265.15, 265.15, 265.05, 261.45, 263.25, 262.45, 
    260.95, 262.45, 261.55, 261.75, 261.95, 260.45, 261.25, 260.25, 260.25, 
    261.05, 261.35, 261.75, 261.95, 260.75, 260.65, 261.35, 261.15, 260.25, 
    261.65, 261.65, 261.15, 260.95, 260.85, 261.15, 261.75, 261.65, 261.65, 
    261.45, 260.85, 261.75, 262.05, 261.95, 261.15, 262.25, 261.15, 262.45, 
    262.35, 263.45, 261.95, 262.65, 263.85, 266.65, 265.75, 265.45, 265.95, 
    265.55, 265.65, 265.75, 262.95, 262.45, 262.35, 262.65, 264.35, 263.95, 
    264.35, 266.95, 267.95, 267.85, 268.15, 268.45, 267.95, 265.65, 266.05, 
    268.55, 266.95, 266.55, 267.05, 268.25, 269.65, 269.85, 265.95, 265.75, 
    264.55, 266.95, 267.85, 267.15, 266.55, 266.35, 266.55, 267.75, 267.75, 
    267.75, 268.05, 267.45, 267.45, 267.75, 267.55, 267.75, 267.75, 268.25, 
    267.45, 267.85, 267.95, 267.65, 269.05, 269.15, 267.05, 265.75, 265.15, 
    265.45, 266.15, 265.95, 266.35, 265.05, 266.75, 268.55, 268.55, 268.75, 
    268.75, 268.85, 269.45, 270.45, 270.95, 270.55, 270.75, 271.45, 271.55, 
    271.65, 272.35, 273.15, 273.95, 274.45, 274.55, 273.15, 273.55, 274.85, 
    274.75, 274.75, 273.65, 271.55, 270.95, 270.55, 270.95, 270.95, 269.85, 
    270.65, 270.15, 271.15, 269.25, 268.85, 268.35, 267.85, 267.15, 267.35, 
    267.15, 267.15, 267.25, 267.25, 267.05, 266.85, 266.85, 265.75, 265.55, 
    265.55, 264.85, 264.95, 264.85, 264.95, 264.85, 264.35, 264.45, 264.45, 
    264.05, 265.45, 265.55, 265.45, 265.55, 265.85, 265.35, 265.45, 265.55, 
    265.45, 265.55, 265.85, 265.85, 266.15, 265.75, 266.15, 265.75, 266.35, 
    264.85, 263.55, 263.05, 263.05, 263.95, 264.55, 265.35, 264.55, 264.45, 
    264.15, 263.55, 263.05, 261.55, 261.25, 261.65, 262.75, 262.05, 262.05, 
    262.75, 261.65, 262.55, 262.15, 260.95, 261.55, 260.05, 259.95, 260.05, 
    259.65, 259.35, 259.85, 259.15, 258.95, 259.05, 259.35, 259.85, 260.15, 
    260.55, 260.85, 261.35, 262.15, 262.75, 262.95, 263.05, 263.05, 263.05, 
    263.25, 263.75, 264.15, 263.65, 265.05, 264.55, 264.95, 265.45, 266.35, 
    266.75, 266.35, 268.05, 269.55, 268.65, 268.45, 268.05, 268.15, 268.45, 
    269.05, 268.45, 268.85, 268.55, 269.95, 269.15, 268.65, 267.35, 268.85, 
    268.95, 269.15, 269.65, 269.35, 269.55, 270.05, 270.35, 270.75, 270.85, 
    270.65, 270.45, 270.55, 270.55, 270.15, 269.75, 269.25, 269.25, 268.65, 
    268.65, 268.45, 268.05, 267.65, 267.25, 266.95, 266.05, 265.75, 265.05, 
    264.05, 264.15, 263.65, 263.15, 263.35, 262.15, 261.85, 260.25, 260.15, 
    258.95, 259.25, 259.15, 257.75, 259.05, 257.65, 259.15, 258.85, 257.65, 
    256.45, 255.65, 256.85, 255.85, 257.45, 257.15, 256.85, 258.35, 257.25, 
    258.95, 257.15, 258.15, 258.35, 259.95, 260.55, 261.25, 261.45, 264.45, 
    265.65, 265.65, 264.45, 265.55, 263.05, 265.35, 265.05, 264.65, 264.75, 
    262.55, 263.65, 261.75, 262.25, 261.55, 261.95, 262.25, 263.05, 263.35, 
    263.25, 262.65, 263.55, 262.35, 260.25, 260.65, 260.35, 260.25, 258.85, 
    260.05, 260.05, 260.75, 261.35, 261.45, 260.75, 261.15, 261.45, 261.55, 
    262.25, 263.35, 263.85, 264.25, 264.45, 264.55, 264.75, 265.15, 265.75, 
    266.15, 266.55, 266.95, 270.05, 270.25, 271.35, 272.35, 273.65, 275.25, 
    274.25, 272.55, 272.05, 271.55, 270.95, 271.95, 272.35, 272.85, 272.35, 
    272.95, 272.05, 271.05, 270.35, 269.95, 269.75, 269.25, 268.65, 268.25, 
    267.95, 267.65, 267.15, 266.55, 266.15, 265.75, 265.15, 264.95, 264.85, 
    264.65, 264.45, 264.15, 263.85, 262.75, 262.65, 262.15, 262.25, 261.85, 
    261.75, 261.65, 261.25, 260.95, 260.65, 260.45, 260.15, 259.85, 259.35, 
    259.65, 257.75, 257.45, 257.75, 256.95, 256.55, 257.15, 257.85, 258.35, 
    258.55, 258.15, 256.65, 257.75, 257.95, 257.95, 258.75, 258.65, 259.25, 
    259.95, 260.75, 261.45, 261.45, 261.65, 261.25, 261.15, 261.25, 261.85, 
    262.25, 262.15, 262.85, 262.75, 262.55, 261.55, 260.45, 260.05, 259.75, 
    259.55, 259.55, 260.45, 260.55, 260.25, 260.75, 260.85, 261.55, 261.75, 
    261.45, 260.75, 260.05, 262.45, 261.95, 266.25, 266.65, 267.15, 267.05, 
    266.85, 266.85, 266.85, 266.85, 266.75, 266.95, 267.65, 267.25, 267.25, 
    267.35, 267.45, 267.85, 268.05, 268.05, 268.35, 268.15, 267.55, 266.55, 
    265.85, 264.85, 264.35, 264.15, 264.55, 263.15, 262.85, 263.25, 262.95, 
    263.55, 262.65, 262.25, 262.65, 262.05, 262.55, 262.05, 261.65, 261.85, 
    261.95, 261.65, 261.55, 262.15, 263.85, 263.85, 264.25, 264.35, 263.85, 
    264.65, 264.15, 264.45, 264.25, 264.75, 265.25, 265.65, 266.15, 266.55, 
    266.85, 267.35, 267.65, 268.25, 267.75, 268.75, 269.05, 270.75, 270.45, 
    272.15, 273.65, 273.65, 273.75, 274.15, 273.45, 273.35, 272.95, 272.85, 
    272.95, 272.95, 272.95, 273.35, 273.65, 273.15, 273.35, 273.45, 273.55, 
    273.45, 273.35, 273.35, 273.55, 273.15, 272.65, 272.55, 272.55, 272.55, 
    272.45, 273.05, 272.75, 272.75, 273.45, 272.75, 272.05, 271.25, 270.75, 
    270.85, 270.85, 271.15, 269.45, 268.25, 268.35, 268.45, 268.55, 270.55, 
    269.65, 268.75, 272.75, 273.15, 272.75, 272.15, 272.25, 272.35, 271.85, 
    271.55, 270.95, 270.65, 270.45, 270.35, 270.05, 268.95, 268.55, 267.95, 
    267.65, 266.85, 266.65, 265.85, 265.75, 265.15, 264.85, 264.05, 263.45, 
    263.35, 262.95, 262.85, 262.65, 262.35, 262.15, 262.15, 262.05, 261.75, 
    261.25, 261.45, 261.05, 260.65, 260.25, 259.25, 259.75, 259.25, 258.15, 
    257.55, 257.35, 257.05, 256.35, 257.25, 256.75, 257.15, 257.15, 257.15, 
    257.25, 257.95, 257.95, 257.95, 257.75, 256.75, 257.15, 257.55, 257.65, 
    257.85, 257.05, 256.25, 256.45, 256.55, 256.35, 256.15, 256.15, 256.35, 
    254.65, 255.85, 256.25, 254.75, 254.85, 255.65, 255.65, 255.15, 256.25, 
    255.95, 255.65, 255.85, 256.15, 255.65, 256.45, 255.65, 256.05, 255.65, 
    255.95, 256.25, 256.25, 256.55, 256.35, 257.35, 256.05, 257.25, 256.55, 
    256.35, 256.15, 256.85, 256.45, 255.95, 255.55, 255.95, 256.85, 256.65, 
    256.55, 256.45, 255.85, 255.35, 255.55, 255.85, 253.85, 255.45, 255.05, 
    254.55, 255.25, 253.65, 255.05, 254.65, 254.55, 254.35, 253.25, 253.35, 
    253.95, 253.25, 253.25, 253.35, 252.95, 252.85, 253.35, 254.15, 254.15, 
    254.15, 254.95, 254.95, 255.15, 254.85, 255.45, 255.35, 254.75, 254.75, 
    254.35, 255.65, 256.25, 256.25, 255.75, 255.05, 254.75, 254.85, 255.75, 
    255.95, 255.65, 255.85, 256.05, 256.75, 256.55, 256.05, 257.75, 257.75, 
    257.95, 258.25, 258.25, 258.55, 258.35, 258.25, 258.25, 258.25, 257.65, 
    258.05, 257.85, 258.15, 258.55, 258.05, 256.55, 256.35, 255.85, 256.45, 
    256.45, 256.75, 255.75, 255.75, 256.05, 255.65, 255.65, 256.15, 255.95, 
    255.35, 253.95, 254.85, 254.85, 256.05, 255.45, 254.75, 256.35, 255.05, 
    255.85, 255.55, 254.55, 255.65, 255.35, 253.85, 255.65, 255.55, 254.95, 
    256.65, 256.55, 255.55, 256.55, 256.75, 256.35, 257.45, 256.75, 257.05, 
    258.45, 256.95, 257.75, 258.75, 257.45, 255.95, 257.85, 255.75, 256.35, 
    256.85, 257.15, 256.65, 256.55, 256.45, 256.35, 256.55, 257.25, 256.95, 
    257.75, 255.55, 255.75, 257.95, 259.05, 259.55, 259.65, 259.35, 259.25, 
    258.95, 258.85, 258.45, 258.15, 258.05, 257.65, 257.35, 257.35, 257.15, 
    256.75, 256.85, 256.35, 256.05, 255.55, 254.45, 253.65, 254.65, 254.85, 
    254.85, 255.05, 254.15, 255.15, 254.55, 255.15, 255.55, 255.05, 256.35, 
    257.35, 258.65, 258.85, 259.05, 259.85, 258.35, 259.85, 261.25, 261.55, 
    260.65, 259.75, 262.75, 262.95, 262.75, 262.25, 262.05, 260.25, 258.95, 
    260.15, 259.85, 258.25, 257.35, 257.05, 258.05, 257.25, 257.35, 257.35, 
    256.95, 256.15, 257.05, 257.25, 257.35, 256.95, 256.65, 256.45, 256.35, 
    256.35, 256.15, 254.65, 253.95, 253.75, 252.55, 252.85, 253.25, 254.25, 
    253.65, 254.65, 255.45, 255.05, 255.35, 255.75, 255.75, 255.55, 256.25, 
    257.25, 256.95, 257.55, 258.75, 260.05, 260.75, 260.45, 261.85, 262.15, 
    261.95, 260.95, 259.65, 260.05, 258.95, 259.45, 257.25, 256.85, 257.75, 
    257.55, 257.05, 256.85, 256.25, 256.25, 257.15, 256.25, 256.25, 254.25, 
    254.45, 255.55, 255.45, 255.05, 254.85, 255.25, 255.25, 256.55, 257.45, 
    258.45, 258.35, 258.45, 259.05, 258.75, 257.95, 258.65, 257.15, 259.15, 
    258.45, 260.45, 260.85, 261.15, 260.85, 261.95, 262.55, 262.75, 263.05, 
    263.75, 262.25, 262.45, 263.65, 262.85, 262.05, 262.55, 263.55, 261.15, 
    262.15, 261.45, 263.65, 263.75, 263.95, 262.25, 264.45, 264.65, 261.75, 
    263.05, 263.05, 262.95, 264.05, 262.95, 264.85, 267.55, 267.65, 267.05, 
    267.15, 266.65, 266.95, 267.15, 267.55, 267.55, 267.85, 267.85, 267.65, 
    267.15, 265.95, 265.75, 265.85, 266.65, 266.45, 265.45, 264.65, 263.95, 
    262.85, 262.95, 262.95, 263.15, 263.35, 263.75, 263.65, 263.75, 263.75, 
    263.75, 263.75, 263.45, 263.15, 262.95, 263.25, 263.45, 263.75, 263.75, 
    264.15, 264.45, 264.65, 264.95, 265.25, 265.65, 266.15, 266.35, 266.85, 
    267.35, 267.75, 267.85, 267.65, 267.05, 266.95, 267.05, 266.95, 266.75, 
    266.55, 266.05, 265.55, 265.05, 265.05, 264.75, 264.05, 262.35, 263.05, 
    261.85, 263.05, 261.75, 261.25, 262.55, 263.05, 262.75, 263.45, 263.95, 
    264.15, 264.35, 264.45, 265.25, 266.25, 266.25, 267.25, 266.75, 270.65, 
    271.25, 271.05, 270.45, 270.45, 270.75, 271.25, 271.75, 271.95, 272.45, 
    272.45, 272.25, 271.95, 271.85, 271.35, 271.65, 272.05, 272.15, 271.65, 
    271.95, 271.45, 270.35, 270.95, 270.05, 268.95, 268.05, 266.95, 266.65, 
    266.15, 267.05, 267.95, 270.15, 269.55, 269.95, 268.65, 269.95, 270.45, 
    271.95, 272.55, 273.15, 272.95, 273.55, 274.55, 273.95, 274.65, 274.85, 
    275.45, 275.75, 275.95, 275.65, 276.35, 275.95, 276.85, 277.75, 276.55, 
    276.15, 275.05, 275.85, 275.55, 275.25, 275.45, 275.75, 274.35, 275.65, 
    276.15, 275.95, 277.35, 277.05, 277.35, 277.45, 277.45, 276.95, 276.05, 
    276.95, 275.55, 275.25, 274.95, 274.55, 273.55, 273.15, 273.15, 272.35, 
    272.05, 272.05, 271.85, 271.55, 271.55, 271.75, 271.75, 270.95, 271.05, 
    271.25, 270.85, 270.85, 271.15, 271.25, 271.35, 271.25, 271.35, 271.45, 
    271.05, 270.55, 270.95, 270.55, 269.65, 269.55, 268.45, 269.15, 269.95, 
    268.85, 269.25, 268.45, 269.35, 269.15, 270.45, 269.55, 270.15, 271.05, 
    270.55, 269.85, 269.05, 268.65, 270.75, 271.05, 270.85, 270.95, 271.05, 
    271.35, 271.95, 272.45, 273.45, 271.05, 271.15, 272.05, 273.05, 272.55, 
    272.85, 272.45, 272.15, 272.35, 273.85, 272.15, 272.35, 272.35, 273.15, 
    273.15, 273.95, 275.25, 274.25, 272.85, 270.65, 272.25, 269.95, 271.35, 
    268.75, 267.15, 269.35, 270.55, 271.05, 269.65, 270.25, 268.25, 268.45, 
    268.55, 266.75, 267.65, 268.25, 265.95, 267.05, 267.45, 266.35, 267.75, 
    267.65, 269.35, 265.85, 266.85, 265.55, 268.35, 267.85, 267.75, 267.45, 
    267.05, 267.45, 266.75, 267.05, 268.85, 264.85, 267.35, 265.85, 264.75, 
    266.05, 266.35, 266.75, 268.95, 269.05, 268.75, 268.55, 267.95, 268.45, 
    267.65, 267.15, 266.25, 265.85, 264.75, 265.15, 265.95, 266.25, 266.95, 
    267.05, 266.85, 266.45, 266.75, 266.35, 266.15, 266.15, 266.25, 266.35, 
    266.05, 266.15, 266.35, 266.25, 266.35, 266.15, 266.15, 265.95, 266.25, 
    266.15, 265.95, 265.55, 265.65, 265.55, 265.35, 264.95, 264.85, 264.55, 
    264.35, 263.95, 263.75, 263.25, 262.95, 263.25, 262.85, 262.45, 262.05, 
    262.15, 261.65, 262.55, 262.45, 262.95, 262.55, 262.55, 262.25, 262.65, 
    263.05, 263.15, 263.45, 263.35, 263.05, 263.25, 263.45, 263.75, 263.55, 
    263.15, 263.45, 263.65, 263.55, 263.65, 263.75, 263.55, 264.25, 264.95, 
    265.15, 265.75, 265.85, 265.75, 265.95, 266.05, 266.05, 266.15, 265.95, 
    266.35, 266.35, 266.45, 266.45, 266.65, 266.55, 266.55, 266.55, 266.35, 
    266.35, 266.25, 266.15, 266.05, 265.75, 265.65, 266.05, 265.65, 265.65, 
    265.55, 265.35, 265.05, 265.15, 265.55, 265.55, 264.95, 265.25, 264.85, 
    264.15, 264.55, 264.15, 264.55, 264.65, 264.35, 264.75, 264.45, 261.95, 
    265.45, 265.35, 265.25, 264.55, 264.55, 264.75, 264.55, 264.95, 264.75, 
    264.85, 264.45, 264.65, 265.05, 265.05, 263.05, 262.55, 264.05, 263.75, 
    265.55, 265.45, 265.85, 265.85, 266.15, 266.35, 266.35, 266.75, 266.75, 
    266.95, 267.15, 266.95, 267.35, 267.35, 267.35, 267.45, 267.35, 267.25, 
    266.85, 266.55, 266.45, 266.45, 265.95, 265.65, 263.45, 263.95, 262.85, 
    263.95, 263.15, 261.95, 261.25, 261.85, 260.35, 261.05, 261.75, 260.45, 
    261.15, 260.75, 259.15, 259.55, 260.15, 260.95, 259.15, 259.75, 259.35, 
    258.85, 259.35, 259.65, 260.85, 258.75, 258.65, 258.35, 261.05, 259.85, 
    260.45, 260.25, 261.55, 261.35, 262.15, 261.45, 261.85, 261.75, 261.25, 
    260.75, 261.05, 261.55, 263.05, 262.25, 261.65, 262.65, 262.85, 263.15, 
    261.95, 263.15, 262.25, 262.85, 263.15, 262.45, 261.35, 260.25, 260.75, 
    261.35, 260.05, 260.95, 261.15, 260.85, 261.05, 261.55, 259.75, 261.15, 
    262.05, 262.45, 263.05, 263.05, 263.55, 263.75, 263.45, 263.45, 263.65, 
    263.65, 264.35, 264.95, 264.85, 265.15, 265.45, 268.75, 269.95, 269.85, 
    270.05, 269.65, 269.75, 269.85, 268.85, 268.75, 269.65, 269.25, 267.75, 
    268.65, 269.05, 268.55, 267.45, 269.05, 268.65, 268.05, 267.95, 268.15, 
    268.05, 268.05, 268.35, 267.65, 267.55, 267.15, 267.55, 266.85, 266.35, 
    266.75, 266.75, 267.55, 267.85, 267.55, 267.05, 267.35, 267.85, 269.55, 
    269.45, 268.15, 268.65, 268.45, 268.25, 267.55, 267.25, 266.45, 267.55, 
    266.85, 266.85, 266.85, 266.65, 267.25, 266.45, 266.65, 267.75, 269.75, 
    270.05, 269.95, 269.95, 269.65, 269.75, 270.15, 269.75, 269.55, 269.55, 
    268.95, 268.75, 268.55, 268.05, 267.35, 267.25, 266.55, 266.35, 266.15, 
    265.95, 265.45, 266.05, 264.55, 263.25, 263.55, 262.85, 260.05, 258.05, 
    261.25, 258.25, 258.25, 258.55, 257.75, 258.55, 256.45, 259.05, 260.35, 
    257.05, 260.65, 257.95, 257.75, 260.65, 260.15, 259.65, 258.55, 257.45, 
    257.45, 256.85, 257.25, 257.05, 257.45, 256.25, 255.85, 256.05, 255.75, 
    255.15, 255.65, 256.15, 255.65, 254.55, 255.85, 255.55, 255.35, 255.25, 
    254.85, 254.75, 254.45, 253.35, 254.05, 254.45, 254.15, 254.75, 252.75, 
    253.55, 252.85, 253.45, 254.05, 252.75, 254.15, 255.15, 253.55, 255.05, 
    256.75, 257.65, 255.95, 255.25, 257.05, 255.85, 254.85, 256.35, 255.75, 
    257.45, 255.75, 254.35, 256.25, 256.55, 256.65, 256.25, 255.35, 255.15, 
    254.85, 255.75, 254.35, 254.85, 253.85, 253.45, 254.45, 255.45, 253.95, 
    254.45, 254.45, 255.55, 254.45, 256.85, 254.75, 253.45, 255.65, 255.25, 
    254.35, 255.05, 255.55, 256.65, 256.95, 255.55, 258.45, 258.75, 258.45, 
    259.05, 259.45, 260.05, 260.25, 260.55, 260.75, 261.05, 261.05, 262.45, 
    263.55, 263.75, 263.85, 264.65, 264.55, 265.45, 269.05, 270.65, 270.75, 
    270.95, 271.25, 270.55, 272.05, 271.85, 271.75, 272.05, 272.05, 272.25, 
    271.55, 271.05, 271.15, 270.95, 270.45, 271.75, 271.95, 271.75, 271.05, 
    270.25, 271.25, 270.25, 270.15, 270.35, 270.65, 270.95, 270.45, 270.35, 
    270.25, 270.15, 269.55, 269.65, 269.25, 270.05, 269.45, 269.55, 269.85, 
    270.35, 270.75, 271.05, 271.35, 271.55, 271.45, 271.25, 271.15, 271.65, 
    271.55, 270.35, 269.75, 269.05, 268.45, 268.15, 269.05, 269.55, 268.65, 
    268.55, 268.25, 268.45, 268.05, 267.35, 268.45, 266.95, 267.55, 268.45, 
    269.55, 269.55, 266.65, 266.75, 266.85, 267.45, 266.05, 264.45, 264.75, 
    265.65, 265.35, 266.45, 263.65, 264.75, 265.25, 265.05, 264.45, 266.65, 
    266.85, 266.35, 266.45, 266.15, 267.35, 267.25, 266.95, 268.65, 270.95, 
    270.65, 270.45, 270.25, 269.45, 267.95, 266.65, 265.55, 267.55, 266.75, 
    263.45, 264.75, 262.25, 262.95, 263.95, 261.45, 263.55, 261.85, 262.05, 
    260.85, 261.15, 260.45, 261.25, 259.35, 261.65, 262.25, 263.35, 265.15, 
    263.75, 263.45, 263.35, 264.35, 264.15, 264.75, 265.35, 265.55, 266.15, 
    267.05, 267.95, 266.85, 267.25, 267.05, 268.25, 267.45, 268.65, 269.05, 
    269.05, 268.35, 268.05, 268.05, 268.45, 268.75, 268.55, 268.85, 269.35, 
    268.75, 269.45, 271.55, 274.45, 274.45, 274.35, 274.35, 273.65, 273.95, 
    274.15, 274.25, 274.35, 274.15, 274.15, 274.45, 274.15, 273.95, 273.85, 
    274.05, 273.45, 272.95, 274.05, 274.25, 274.35, 274.45, 274.45, 274.45, 
    274.35, 274.25, 273.15, 273.35, 273.55, 272.85, 272.45, 272.25, 272.15, 
    272.65, 272.35, 271.05, 271.95, 271.75, 271.95, 271.85, 271.95, 272.35, 
    272.55, 272.15, 273.65, 274.65, 275.05, 274.65, 275.05, 275.15, 274.65, 
    275.35, 275.15, 275.15, 274.95, 275.05, 275.15, 274.05, 272.05, 269.95, 
    269.25, 267.95, 267.15, 265.95, 266.85, 264.75, 264.05, 262.35, 261.45, 
    261.35, 262.15, 262.05, 260.95, 261.35, 258.85, 258.75, 259.25, 258.25, 
    259.35, 259.45, 260.15, 259.25, 259.25, 259.75, 259.25, 261.05, 258.15, 
    259.65, 260.25, 257.15, 256.05, 257.55, 260.15, 263.25, 259.75, 262.05, 
    261.55, 262.55, 262.95, 263.85, 263.75, 263.85, 264.65, 265.85, 265.55, 
    266.15, 266.45, 267.15, 266.65, 266.85, 267.35, 268.05, 269.05, 269.15, 
    269.95, 270.75, 270.95, 271.65, 271.05, 271.05, 271.95, 271.45, 269.95, 
    269.05, 269.35, 268.35, 267.95, 266.35, 266.45, 262.95, 263.35, 262.25, 
    264.55, 264.25, 263.55, 263.65, 262.65, 263.15, 264.05, 263.45, 265.85, 
    267.05, 267.05, 264.95, 266.85, 269.05, 269.25, 266.45, 268.45, 267.55, 
    269.55, 268.75, 269.35, 269.65, 268.95, 269.25, 269.85, 269.05, 270.05, 
    270.45, 270.75, 270.45, 271.45, 271.85, 275.45, 274.95, 274.95, 274.85, 
    275.25, 274.85, 273.75, 272.65, 272.75, 274.15, 273.55, 273.55, 274.55, 
    274.95, 273.45, 274.75, 273.65, 273.35, 272.85, 271.95, 269.45, 270.85, 
    271.75, 271.25, 270.65, 270.65, 270.95, 272.25, 272.15, 271.75, 271.15, 
    271.75, 271.75, 272.05, 272.45, 272.55, 272.55, 272.95, 273.05, 273.15, 
    271.65, 271.85, 271.65, 271.95, 273.05, 273.05, 272.55, 272.35, 272.35, 
    271.75, 271.95, 269.65, 269.25, 267.75, 269.05, 266.95, 268.05, 267.85, 
    267.15, 268.75, 266.85, 266.95, 264.75, 267.45, 265.45, 265.25, 266.65, 
    271.05, 270.35, 270.45, 270.85, 272.95, 272.75, 272.55, 271.85, 271.25, 
    272.75, 269.65, 270.95, 269.55, 270.15, 269.85, 269.35, 268.25, 269.05, 
    268.95, 266.15, 267.55, 268.85, 268.55, 268.05, 267.15, 269.45, 269.35, 
    270.05, 270.95, 269.55, 269.05, 269.15, 268.15, 267.35, 267.45, 267.05, 
    266.75, 267.15, 266.85, 267.25, 266.65, 266.25, 266.85, 267.05, 266.65, 
    265.45, 266.25, 266.95, 266.55, 265.05, 265.35, 265.85, 266.35, 267.35, 
    266.05, 266.75, 266.25, 266.25, 266.95, 266.85, 267.45, 266.95, 267.75, 
    269.15, 268.75, 268.25, 269.25, 269.15, 268.65, 268.85, 268.95, 268.75, 
    269.35, 269.45, 268.65, 269.45, 269.15, 269.15, 269.05, 269.55, 269.05, 
    269.15, 269.25, 269.15, 269.05, 269.15, 269.15, 266.75, 267.95, 267.35, 
    267.75, 268.05, 268.25, 268.15, 267.55, 267.65, 266.95, 266.85, 266.85, 
    267.45, 266.85, 267.75, 267.35, 267.25, 267.25, 268.75, 268.55, 268.05, 
    267.95, 267.75, 268.15, 267.85, 268.05, 268.95, 269.25, 271.35, 270.65, 
    270.65, 270.45, 269.55, 269.45, 268.75, 267.75, 267.95, 268.85, 269.65, 
    268.85, 268.85, 269.35, 269.05, 269.75, 269.55, 271.05, 271.85, 271.65, 
    272.25, 272.25, 272.35, 272.45, 273.95, 274.15, 274.05, 274.15, 274.35, 
    273.75, 273.65, 274.65, 274.15, 273.55, 273.65, 273.85, 273.25, 272.85, 
    271.95, 271.45, 270.95, 270.45, 269.85, 268.55, 266.45, 266.05, 264.95, 
    266.75, 264.75, 263.15, 264.15, 265.35, 264.35, 265.45, 265.85, 266.85, 
    266.55, 263.55, 263.35, 265.65, 266.05, 267.75, 269.55, 270.95, 270.35, 
    271.85, 271.55, 271.65, 271.05, 271.45, 271.15, 271.35, 271.35, 268.65, 
    269.95, 272.35, 272.35, 271.95, 271.65, 271.85, 271.35, 271.65, 271.75, 
    271.95, 271.95, 271.85, 272.15, 272.55, 272.55, 272.55, 272.75, 272.75, 
    273.05, 272.95, 273.15, 273.05, 272.85, 273.75, 272.45, 271.75, 272.75, 
    271.75, 272.25, 272.35, 272.35, 271.25, 270.05, 271.45, 271.65, 271.75, 
    270.45, 270.15, 270.75, 269.15, 268.95, 269.65, 268.95, 266.05, 267.25, 
    266.95, 269.15, 267.85, 267.55, 269.55, 267.95, 267.85, 269.45, 267.25, 
    266.95, 267.25, 266.35, 269.75, 270.05, 270.35, 270.85, 272.05, 272.95, 
    271.45, 271.05, 271.15, 270.65, 271.15, 271.15, 271.35, 270.55, 270.15, 
    269.55, 271.75, 269.35, 269.25, 270.55, 269.15, 270.75, 271.45, 271.95, 
    270.75, 272.25, 271.75, 271.15, 271.35, 271.65, 271.95, 272.05, 271.45, 
    271.55, 271.75, 271.85, 272.35, 272.65, 272.15, 272.45, 272.75, 272.95, 
    272.75, 272.15, 271.75, 272.75, 273.15, 272.55, 273.25, 273.45, 272.85, 
    272.15, 272.85, 272.85, 273.25, 272.75, 272.75, 273.25, 273.45, 272.85, 
    272.35, 271.95, 271.75, 270.85, 271.55, 271.85, 269.75, 270.15, 273.05, 
    272.25, 272.45, 272.85, 272.95, 273.05, 272.85, 272.45, 271.95, 271.85, 
    271.15, 271.45, 272.55, 272.05, 271.95, 272.55, 272.85, 272.65, 272.55, 
    271.45, 272.45, 272.95, 272.95, 272.25, 272.25, 272.05, 272.15, 272.45, 
    273.25, 273.15, 272.95, 272.85, 273.25, 273.25, 272.75, 273.45, 273.35, 
    272.65, 273.25, 272.35, 272.55, 273.15, 274.75, 273.85, 273.55, 273.75, 
    274.45, 273.75, 274.65, 275.35, 275.75, 275.75, 275.65, 275.65, 275.05, 
    274.15, 274.35, 275.25, 274.95, 273.75, 274.95, 273.95, 275.05, 274.05, 
    275.45, 275.45, 275.45, 274.45, 274.55, 274.75, 273.85, 272.65, 273.05, 
    273.15, 272.85, 273.85, 273.45, 273.35, 273.05, 272.75, 272.95, 272.95, 
    272.45, 272.55, 272.75, 272.25, 272.85, 272.05, 274.05, 274.75, 274.75, 
    274.85, 275.15, 276.15, 276.35, 277.95, 276.95, 277.15, 277.25, 277.15, 
    277.65, 277.85, 277.75, 276.55, 277.05, 277.55, 278.15, 277.95, 277.55, 
    278.05, 277.95, 278.05, 277.95, 277.55, 276.85, 276.35, 277.05, 276.25, 
    275.55, 275.85, 275.75, 275.75, 275.65, 275.75, 275.55, 274.85, 274.15, 
    274.35, 273.85, 274.25, 273.75, 273.15, 273.45, 273.25, 273.15, 272.55, 
    272.45, 272.45, 272.45, 272.95, 272.65, 272.65, 272.85, 272.85, 273.45, 
    272.85, 273.45, 273.65, 273.85, 274.15, 274.35, 274.55, 274.95, 274.15, 
    273.85, 273.45, 273.85, 273.15, 272.25, 271.75, 272.15, 271.95, 271.85, 
    272.05, 272.05, 272.15, 272.15, 272.15, 272.15, 272.65, 272.45, 272.65, 
    272.85, 272.65, 273.05, 273.25, 273.35, 273.75, 273.35, 273.65, 273.65, 
    273.95, 273.35, 273.25, 272.55, 271.85, 273.85, 273.05, 272.15, 272.35, 
    273.05, 274.25, 274.45, 274.05, 273.85, 273.85, 273.55, 273.75, 273.25, 
    269.95, 271.25, 271.65, 271.55, 271.35, 272.15, 270.75, 270.25, 270.15, 
    271.55, 271.45, 271.25, 271.75, 271.15, 271.55, 271.15, 271.15, 271.35, 
    269.95, 269.95, 270.75, 272.05, 273.25, 273.35, 273.55, 273.45, 273.45, 
    271.85, 272.35, 272.15, 273.15, 274.05, 274.35, 274.15, 274.35, 273.55, 
    273.15, 273.25, 272.85, 273.35, 273.05, 272.95, 272.85, 272.75, 271.95, 
    271.65, 271.35, 271.15, 270.35, 270.15, 270.25, 270.65, 270.55, 270.15, 
    270.95, 270.85, 270.75, 270.15, 269.75, 269.75, 269.75, 269.65, 269.75, 
    269.65, 269.25, 269.65, 269.15, 268.85, 268.85, 269.25, 267.75, 268.95, 
    268.85, 266.95, 265.95, 264.45, 264.05, 264.05, 264.75, 265.55, 264.65, 
    265.15, 265.25, 265.35, 265.85, 266.05, 266.35, 266.65, 266.95, 267.25, 
    267.25, 267.45, 267.65, 267.75, 267.65, 267.15, 266.95, 266.65, 266.75, 
    268.15, 269.85, 271.15, 271.15, 271.45, 271.75, 271.65, 271.95, 272.35, 
    272.75, 272.25, 272.05, 272.45, 271.65, 271.25, 271.25, 271.15, 271.25, 
    270.95, 270.85, 271.25, 271.05, 271.35, 271.95, 272.15, 272.05, 272.45, 
    271.95, 272.55, 271.55, 271.85, 272.55, 272.35, 272.05, 272.45, 271.95, 
    271.85, 272.05, 271.85, 271.75, 271.55, 271.45, 270.95, 270.15, 269.85, 
    269.95, 269.05, 269.85, 269.25, 269.65, 269.45, 269.65, 269.55, 269.15, 
    269.45, 269.75, 269.75, 269.15, 269.95, 268.75, 269.25, 268.55, 267.65, 
    267.45, 267.15, 268.25, 268.35, 266.15, 265.35, 265.75, 265.85, 267.25, 
    266.55, 268.15, 268.05, 268.45, 268.95, 268.95, 267.85, 269.05, 269.85, 
    269.45, 269.75, 270.05, 268.25, 269.75, 269.95, 270.05, 269.95, 269.85, 
    270.05, 269.85, 269.75, 269.85, 270.25, 270.65, 270.75, 270.05, 271.25, 
    270.65, 271.65, 271.55, 271.85, 272.05, 272.35, 272.55, 272.45, 272.95, 
    272.95, 272.65, 272.95, 273.05, 272.75, 272.45, 272.15, 272.55, 272.55, 
    272.35, 272.95, 273.15, 273.45, 273.55, 273.55, 273.65, 273.65, 273.45, 
    272.95, 272.35, 272.55, 271.95, 272.55, 269.95, 270.75, 270.45, 270.45, 
    270.15, 270.35, 270.15, 269.45, 269.55, 268.25, 266.85, 266.85, 266.95, 
    267.95, 267.35, 267.75, 268.55, 268.45, 269.25, 267.75, 267.15, 266.85, 
    265.35, 264.85, 264.65, 264.75, 264.75, 264.95, 265.25, 264.35, 264.15, 
    264.85, 265.45, 264.25, 264.45, 266.25, 264.85, 265.85, 265.35, 264.85, 
    264.25, 264.05, 263.75, 262.55, 262.05, 262.05, 259.85, 259.05, 259.15, 
    258.25, 259.25, 260.15, 258.95, 259.45, 258.85, 258.45, 257.75, 258.95, 
    260.75, 265.15, 263.85, 264.55, 264.05, 264.25, 263.85, 263.85, 264.75, 
    264.85, 264.75, 264.25, 262.65, 262.45, 262.45, 260.95, 261.95, 263.65, 
    261.15, 260.75, 260.25, 259.45, 260.85, 261.15, 260.85, 260.85, 260.05, 
    260.05, 259.15, 258.45, 257.95, 257.75, 257.65, 258.45, 257.35, 258.05, 
    256.75, 257.35, 258.05, 257.55, 258.45, 259.05, 258.95, 259.55, 259.85, 
    259.75, 259.65, 259.65, 259.95, 260.25, 260.25, 260.45, 261.25, 261.15, 
    261.75, 262.95, 263.25, 263.75, 264.15, 264.45, 264.45, 264.25, 265.15, 
    263.45, 264.45, 265.45, 265.95, 266.05, 266.45, 266.95, 268.95, 269.85, 
    270.15, 271.55, 272.05, 271.15, 272.25, 273.15, 272.05, 271.55, 271.15, 
    271.15, 271.15, 270.75, 270.35, 269.85, 269.45, 268.95, 268.55, 268.05, 
    267.65, 267.45, 267.05, 266.75, 266.55, 265.35, 265.55, 265.75, 265.55, 
    263.75, 262.45, 261.45, 260.95, 261.35, 261.35, 261.15, 260.25, 259.75, 
    260.85, 262.95, 262.05, 261.95, 261.25, 261.75, 262.25, 262.05, 263.75, 
    263.85, 264.35, 265.05, 265.75, 265.45, 266.15, 266.25, 266.25, 269.15, 
    268.85, 268.95, 268.35, 268.25, 268.15, 268.15, 268.25, 267.35, 266.65, 
    268.55, 268.45, 267.35, 265.15, 266.65, 265.15, 265.15, 265.65, 266.25, 
    267.25, 268.65, 271.25, 269.25, 271.85, 271.65, 272.25, 272.15, 272.75, 
    273.15, 273.25, 273.45, 273.65, 273.85, 274.05, 274.15, 274.75, 275.05, 
    275.85, 275.65, 275.25, 275.05, 274.25, 273.75, 274.35, 273.05, 272.45, 
    272.75, 273.95, 274.05, 274.65, 274.35, 273.65, 273.75, 274.05, 274.45, 
    274.55, 274.55, 274.55, 274.25, 273.85, 273.95, 273.35, 273.85, 274.05, 
    274.15, 274.65, 274.75, 274.75, 275.05, 274.55, 275.25, 274.65, 274.95, 
    274.75, 274.05, 274.65, 274.25, 273.75, 273.25, 274.45, 273.25, 273.25, 
    272.95, 273.05, 272.95, 272.35, 272.65, 272.45, 272.35, 272.15, 272.45, 
    272.45, 272.25, 271.45, 271.65, 272.05, 272.35, 272.55, 272.35, 272.65, 
    272.65, 272.15, 272.55, 272.25, 271.65, 271.15, 271.35, 271.05, 270.65, 
    270.35, 270.15, 270.95, 270.25, 270.15, 270.15, 268.85, 268.75, 269.55, 
    269.75, 269.45, 269.55, 269.55, 268.55, 268.55, 268.85, 268.85, 268.65, 
    268.75, 268.05, 268.25, 267.85, 267.85, 267.55, 267.85, 267.95, 267.55, 
    267.95, 267.65, 267.65, 268.25, 267.95, 268.05, 267.85, 268.05, 267.85, 
    267.95, 268.15, 268.25, 268.35, 268.25, 267.85, 267.25, 267.25, 266.45, 
    266.45, 266.25, 265.75, 266.25, 265.65, 265.55, 264.85, 264.35, 264.05, 
    264.35, 263.25, 264.75, 264.95, 264.55, 264.35, 263.95, 263.95, 263.05, 
    262.65, 260.55, 259.85, 260.25, 260.05, 258.55, 258.85, 259.45, 257.65, 
    258.05, 257.75, 258.25, 255.25, 256.25, 255.15, 256.55, 256.15, 256.75, 
    257.55, 256.35, 255.25, 257.85, 257.75, 259.15, 260.25, 258.45, 259.25, 
    259.05, 257.05, 258.75, 256.95, 259.45, 258.05, 257.35, 259.35, 256.45, 
    258.75, 258.95, 258.55, 258.25, 257.65, 257.65, 259.65, 259.05, 258.45, 
    258.45, 259.25, 260.75, 260.55, 259.15, 259.35, 259.35, 258.85, 259.25, 
    257.75, 259.05, 258.35, 257.85, 257.45, 257.15, 257.05, 257.75, 258.15, 
    257.35, 256.55, 257.55, 256.95, 258.35, 259.15, 258.15, 259.05, 258.95, 
    259.05, 259.65, 259.45, 260.15, 258.55, 259.25, 258.05, 257.95, 257.45, 
    258.15, 256.85, 257.75, 258.15, 258.05, 257.85, 255.95, 257.15, 257.95, 
    255.95, 255.75, 256.65, 257.55, 256.75, 259.05, 259.95, 259.35, 257.35, 
    258.65, 257.25, 256.85, 255.95, 259.65, 259.85, 259.95, 263.15, 260.95, 
    258.75, 259.05, 259.25, 261.65, 262.35, 260.75, 261.95, 262.75, 262.55, 
    262.55, 263.55, 263.55, 263.95, 264.05, 264.05, 264.05, 264.15, 264.65, 
    264.75, 264.75, 265.25, 264.75, 264.65, 264.35, 264.15, 263.85, 263.85, 
    264.15, 263.95, 264.35, 264.35, 264.25, 264.25, 264.15, 263.75, 263.65, 
    263.65, 263.65, 263.55, 263.75, 262.65, 263.25, 262.45, 261.65, 262.15, 
    263.25, 261.75, 262.65, 262.75, 263.35, 263.65, 261.85, 258.65, 259.85, 
    261.05, 260.95, 260.65, 258.65, 261.25, 260.85, 260.85, 259.25, 257.75, 
    258.55, 260.25, 259.05, 259.45, 257.45, 258.35, 256.55, 256.75, 256.15, 
    257.15, 256.85, 257.05, 255.75, 257.15, 255.85, 255.55, 254.65, 256.15, 
    256.25, 258.25, 258.55, 259.65, 260.75, 260.85, 260.45, 260.55, 260.95, 
    259.95, 260.75, 260.45, 260.55, 260.45, 260.55, 261.05, 260.55, 260.35, 
    260.15, 260.15, 259.75, 261.55, 261.55, 261.35, 260.55, 261.45, 261.15, 
    261.25, 261.75, 262.85, 263.25, 260.15, 260.35, 260.35, 258.75, 259.45, 
    259.05, 258.25, 258.15, 258.25, 257.55, 258.45, 258.05, 257.55, 258.85, 
    258.15, 257.35, 258.35, 257.15, 258.05, 259.75, 258.85, 260.05, 260.45, 
    259.45, 258.65, 259.45, 257.95, 256.75, 255.95, 257.75, 257.75, 256.35, 
    256.85, 256.85, 255.75, 254.95, 255.75, 256.25, 255.85, 258.75, 258.25, 
    258.45, 258.15, 258.05, 258.35, 258.75, 257.85, 257.15, 256.15, 255.45, 
    255.75, 255.85, 255.85, 256.65, 255.65, 256.75, 255.35, 255.05, 254.75, 
    255.25, 255.65, 252.65, 253.65, 252.65, 253.45, 254.45, 254.05, 256.65, 
    255.95, 255.95, 255.55, 256.15, 255.55, 254.15, 253.85, 255.15, 255.35, 
    254.65, 255.15, 255.95, 256.85, 256.45, 256.25, 260.35, 257.65, 259.15, 
    261.85, 262.75, 262.85, 263.35, 262.85, 262.25, 262.35, 262.75, 262.75, 
    264.05, 264.15, 264.05, 263.05, 263.55, 261.65, 262.15, 260.35, 259.25, 
    258.95, 258.75, 257.75, 257.45, 257.75, 257.95, 257.95, 259.35, 258.15, 
    260.25, 259.45, 260.15, 261.25, 262.35, 263.65, 262.95, 262.65, 262.45, 
    261.85, 259.75, 260.25, 258.65, 259.95, 259.35, 257.75, 259.95, 259.55, 
    258.55, 258.25, 261.05, 260.45, 260.85, 260.45, 260.35, 260.55, 264.15, 
    263.75, 264.75, 263.95, 263.75, 263.65, 263.35, 263.65, 265.25, 265.45, 
    266.25, 267.15, 268.15, 268.25, 267.45, 268.05, 268.25, 267.65, 270.65, 
    269.75, 269.65, 269.35, 269.05, 268.35, 267.45, 266.95, 266.75, 266.25, 
    265.25, 264.95, 265.15, 265.15, 264.95, 264.15, 263.45, 262.05, 262.45, 
    261.75, 262.65, 262.15, 262.55, 262.95, 261.85, 261.65, 261.45, 261.65, 
    260.75, 261.15, 261.65, 261.65, 261.25, 262.45, 261.95, 261.05, 260.65, 
    260.75, 257.95, 257.35, 257.55, 257.65, 257.55, 258.65, 255.55, 256.35, 
    257.15, 253.55, 257.35, 256.75, 257.55, 257.55, 258.05, 258.85, 258.95, 
    259.85, 258.65, 258.05, 259.05, 259.35, 258.85, 258.75, 257.25, 258.55, 
    257.75, 258.35, 258.05, 258.65, 256.85, 257.85, 258.15, 258.85, 259.15, 
    258.65, 259.85, 259.75, 260.65, 261.45, 262.05, 262.15, 261.85, 260.35, 
    260.75, 259.35, 259.05, 260.25, 259.75, 259.75, 259.15, 257.35, 257.15, 
    254.15, 254.65, 254.15, 257.25, 255.85, 255.45, 256.45, 256.75, 257.85, 
    258.05, 259.55, 259.55, 259.15, 259.05, 259.05, 259.35, 259.65, 258.95, 
    258.05, 257.05, 256.75, 259.05, 259.95, 259.95, 256.85, 257.35, 257.45, 
    256.55, 256.15, 256.35, 255.55, 256.75, 257.75, 260.35, 259.15, 259.65, 
    258.55, 259.45, 258.75, 258.05, 257.95, 257.15, 256.15, 255.95, 256.35, 
    256.25, 256.05, 255.35, 256.75, 256.95, 255.55, 255.95, 256.05, 254.85, 
    254.75, 254.55, 254.75, 257.45, 257.65, 256.95, 260.15, 257.55, 257.35, 
    259.95, 258.15, 257.75, 258.05, 256.85, 256.55, 256.45, 255.35, 254.05, 
    253.15, 255.05, 254.55, 254.65, 255.65, 254.55, 255.55, 254.85, 256.75, 
    256.35, 258.85, 258.55, 259.75, 260.05, 259.45, 257.35, 259.35, 258.95, 
    259.95, 259.35, 256.35, 257.25, 257.05, 255.25, 257.65, 256.35, 253.45, 
    257.25, 255.95, 256.65, 255.85, 256.95, 257.95, 259.05, 259.35, 258.65, 
    259.05, 259.25, 258.85, 258.75, 256.85, 258.15, 257.25, 256.55, 256.55, 
    255.45, 254.45, 254.85, 254.25, 253.25, 254.95, 258.25, 257.15, 255.05, 
    257.05, 256.35, 257.35, 258.85, 258.55, 261.65, 259.35, 259.55, 259.55, 
    259.95, 258.15, 257.95, 257.65, 256.15, 257.65, 257.35, 254.45, 257.15, 
    256.25, 254.95, 255.15, 256.15, 254.25, 254.15, 254.65, 256.75, 256.85, 
    257.75, 259.65, 259.75, 259.55, 260.95, 259.35, 260.15, 259.55, 258.25, 
    257.75, 256.75, 257.45, 256.65, 255.15, 255.45, 255.45, 255.75, 257.15, 
    257.25, 258.75, 258.25, 258.35, 258.65, 259.95, 261.05, 260.35, 261.95, 
    261.85, 262.85, 262.55, 263.15, 262.45, 262.05, 262.85, 262.55, 262.05, 
    263.55, 263.65, 263.15, 263.05, 263.25, 263.65, 263.65, 263.45, 263.45, 
    265.05, 265.35, 267.05, 267.95, 268.65, 269.55, 268.75, 269.55, 269.35, 
    269.05, 268.95, 269.35, 269.55, 269.65, 269.95, 269.95, 270.25, 270.15, 
    270.45, 270.05, 270.35, 270.85, 270.25, 270.85, 272.35, 272.25, 272.85, 
    272.75, 272.85, 273.05, 272.65, 272.85, 272.95, 272.75, 272.95, 272.35, 
    272.05, 271.65, 270.55, 270.35, 269.15, 266.95, 265.85, 264.95, 264.65, 
    265.05, 265.75, 265.95, 266.05, 266.85, 266.85, 266.75, 267.35, 267.45, 
    267.95, 266.85, 266.35, 265.75, 265.25, 264.15, 263.05, 263.15, 262.45, 
    261.85, 261.45, 261.45, 261.05, 260.75, 260.35, 258.45, 258.45, 257.65, 
    257.95, 257.35, 256.95, 257.65, 258.95, 259.25, 259.05, 259.35, 260.05, 
    259.25, 259.45, 258.25, 257.75, 256.55, 255.15, 255.45, 253.75, 255.05, 
    253.65, 254.35, 254.35, 254.15, 253.65, 253.45, 254.15, 254.35, 256.55, 
    255.95, 256.75, 257.45, 256.75, 259.65, 259.55, 258.75, 258.95, 257.65, 
    256.25, 257.45, 256.35, 254.45, 256.65, 255.05, 253.65, 255.85, 255.75, 
    253.35, 254.65, 254.65, 254.85, 255.55, 257.25, 258.75, 258.95, 259.75, 
    258.85, 261.15, 259.25, 260.75, 260.65, 257.45, 258.05, 258.05, 255.95, 
    255.05, 253.75, 254.85, 255.55, 255.85, 256.05, 256.35, 256.45, 257.25, 
    257.95, 258.35, 258.35, 260.55, 261.25, 262.75, 265.55, 262.35, 263.05, 
    263.05, 262.95, 263.55, 263.05, 262.85, 263.25, 263.45, 261.55, 261.55, 
    263.25, 264.25, 264.95, 264.65, 265.75, 265.55, 266.35, 267.25, 267.55, 
    269.35, 270.75, 269.95, 269.75, 269.95, 271.15, 271.35, 271.75, 271.75, 
    271.65, 270.75, 270.25, 270.25, 270.35, 270.05, 269.85, 270.35, 269.95, 
    269.55, 269.25, 269.05, 268.25, 267.85, 267.45, 265.85, 265.15, 264.85, 
    263.25, 263.65, 263.75, 263.45, 262.75, 261.85, 261.35, 262.25, 261.55, 
    260.55, 260.25, 260.55, 259.15, 259.15, 256.95, 257.75, 258.35, 255.05, 
    256.05, 258.55, 257.45, 258.45, 259.45, 259.65, 259.55, 260.15, 259.25, 
    259.75, 259.25, 260.35, 258.85, 256.75, 256.45, 255.25, 256.35, 255.15, 
    255.45, 254.05, 255.95, 254.85, 255.15, 255.05, 256.85, 257.65, 255.95, 
    256.95, 258.15, 259.55, 259.55, 260.05, 261.15, 261.05, 262.45, 261.05, 
    261.05, 260.65, 259.55, 257.35, 256.85, 258.45, 257.55, 257.95, 256.35, 
    257.55, 256.55, 256.95, 257.55, 257.65, 260.15, 260.75, 263.75, 262.05, 
    262.85, 263.95, 264.35, 264.75, 265.25, 265.35, 265.05, 265.05, 262.95, 
    262.65, 262.55, 262.75, 263.55, 262.65, 262.45, 263.05, 261.75, 263.35, 
    263.25, 263.35, 265.25, 265.95, 264.75, 266.05, 267.35, 266.25, 267.15, 
    266.55, 266.45, 266.45, 264.95, 264.55, 263.45, 262.25, 262.15, 261.35, 
    260.65, 260.05, 260.65, 259.75, 260.25, 260.45, 259.15, 260.35, 261.35, 
    261.95, 261.75, 261.65, 263.45, 263.25, 263.25, 262.95, 262.25, 261.45, 
    261.05, 260.35, 258.55, 258.35, 258.35, 257.95, 258.95, 258.55, 258.55, 
    257.95, 260.55, 259.65, 259.75, 261.95, 263.25, 262.95, 263.15, 264.05, 
    264.25, 265.35, 265.25, 266.75, 268.15, 265.85, 265.75, 264.25, 263.95, 
    263.95, 262.45, 262.25, 261.85, 260.15, 261.65, 261.25, 260.55, 260.45, 
    261.65, 262.65, 263.85, 264.35, 264.85, 266.05, 267.15, 266.15, 265.85, 
    265.45, 265.05, 264.75, 263.55, 262.45, 259.65, 258.45, 257.55, 257.95, 
    257.85, 258.45, 258.25, 258.85, 260.05, 260.65, 262.65, 262.55, 265.65, 
    264.45, 266.85, 265.75, 265.65, 266.35, 265.65, 264.75, 265.25, 264.95, 
    264.55, 263.55, 262.95, 262.15, 260.95, 259.65, 260.15, 259.35, 257.55, 
    258.85, 258.15, 260.55, 259.25, 261.95, 261.85, 261.35, 262.15, 264.05, 
    266.85, 267.45, 266.55, 265.85, 265.35, 264.85, 264.35, 263.65, 261.05, 
    261.25, 259.15, 259.25, 258.15, 257.65, 257.95, 259.25, 259.05, 259.85, 
    261.25, 261.15, 261.05, 261.25, 261.95, 262.05, 263.05, 262.95, 263.25, 
    263.35, 262.85, 262.55, 262.55, 261.95, 261.55, 261.85, 259.85, 258.75, 
    258.25, 258.25, 257.15, 257.75, 259.05, 259.95, 263.55, 264.25, 264.55, 
    264.95, 265.45, 266.55, 266.75, 267.95, 266.85, 266.75, 266.85, 265.95, 
    264.15, 264.85, 262.55, 261.45, 260.35, 260.15, 258.75, 260.45, 260.05, 
    260.65, 261.85, 261.35, 262.45, 263.75, 264.75, 264.75, 264.65, 264.55, 
    266.35, 267.05, 266.55, 267.35, 266.95, 266.05, 265.65, 264.55, 264.55, 
    262.05, 261.35, 261.35, 262.15, 262.05, 262.25, 262.95, 263.15, 264.95, 
    265.25, 265.95, 265.95, 265.75, 266.45, 266.05, 266.75, 267.25, 267.75, 
    267.65, 266.85, 265.95, 266.95, 266.55, 266.15, 266.05, 265.45, 265.45, 
    266.35, 266.35, 266.25, 266.75, 266.95, 267.15, 266.85, 267.15, 267.25, 
    267.75, 267.65, 268.05, 268.15, 268.25, 267.75, 267.55, 267.35, 266.95, 
    266.95, 266.95, 266.65, 266.45, 266.65, 266.35, 266.35, 265.95, 266.15, 
    266.05, 265.85, 265.25, 265.95, 266.85, 266.45, 266.25, 265.45, 266.45, 
    267.05, 266.45, 267.05, 266.85, 266.45, 265.55, 266.35, 264.95, 265.35, 
    263.25, 262.25, 261.05, 260.45, 259.35, 260.75, 261.15, 261.15, 261.75, 
    262.45, 263.15, 266.05, 264.75, 265.25, 265.35, 265.55, 265.55, 265.85, 
    265.35, 264.65, 264.65, 264.95, 264.35, 263.65, 262.05, 261.25, 260.65, 
    260.95, 261.55, 261.25, 260.15, 261.55, 262.95, 262.65, 264.15, 265.95, 
    267.75, 267.95, 270.55, 266.95, 269.95, 268.35, 267.75, 267.25, 266.85, 
    267.05, 266.65, 266.35, 263.75, 263.15, 264.45, 263.45, 263.45, 263.95, 
    265.85, 265.15, 265.35, 266.45, 267.75, 267.85, 270.35, 268.85, 270.15, 
    269.95, 271.25, 270.05, 270.15, 270.55, 269.75, 270.35, 270.35, 269.85, 
    269.45, 270.35, 273.35, 272.95, 272.95, 272.95, 272.95, 273.05, 273.05, 
    273.15, 273.25, 273.65, 273.45, 274.75, 274.15, 274.55, 273.75, 274.75, 
    275.15, 274.65, 274.45, 274.45, 274.55, 274.55, 274.35, 274.75, 274.65, 
    274.45, 274.05, 274.05, 274.15, 274.25, 274.05, 274.25, 274.45, 274.35, 
    274.65, 274.55, 275.05, 275.35, 275.25, 275.35, 275.35, 275.45, 275.45, 
    275.15, 275.15, 275.05, 275.15, 275.05, 274.65, 274.45, 274.45, 274.75, 
    274.35, 274.45, 274.55, 274.35, 274.25, 274.25, 274.35, 274.75, 274.75, 
    274.05, 272.85, 271.85, 272.45, 272.45, 271.65, 270.75, 270.05, 269.25, 
    268.85, 269.15, 268.65, 268.95, 268.75, 268.65, 268.55, 268.45, 269.25, 
    269.55, 268.75, 270.75, 270.05, 269.15, 270.75, 271.15, 270.95, 270.75, 
    271.65, 272.45, 272.35, 270.15, 269.85, 270.05, 269.35, 268.95, 269.05, 
    268.85, 268.65, 268.25, 267.55, 267.95, 268.55, 267.95, 267.75, 268.15, 
    268.05, 268.75, 269.15, 270.05, 268.85, 268.85, 269.05, 267.95, 267.75, 
    266.95, 266.25, 265.45, 265.25, 264.85, 264.65, 264.35, 263.95, 264.05, 
    263.75, 264.15, 263.95, 264.05, 264.15, 264.25, 264.45, 264.65, 265.25, 
    264.55, 265.05, 265.25, 264.65, 264.85, 264.55, 264.55, 264.45, 264.15, 
    263.55, 261.25, 261.15, 260.25, 258.85, 259.55, 259.85, 261.55, 260.55, 
    261.25, 262.55, 263.05, 263.45, 263.75, 265.05, 265.35, 265.75, 265.95, 
    266.65, 266.55, 265.55, 266.25, 265.85, 265.15, 264.55, 264.25, 263.95, 
    263.25, 262.45, 263.05, 262.75, 263.85, 263.45, 264.25, 265.35, 266.85, 
    266.25, 267.55, 267.35, 267.75, 267.35, 267.55, 267.05, 266.65, 266.55, 
    266.65, 266.05, 265.95, 265.75, 265.45, 265.45, 264.95, 264.75, 264.75, 
    264.75, 264.75, 264.75, 264.95, 265.15, 265.25, 265.05, 264.95, 265.05, 
    265.15, 265.35, 265.45, 265.55, 265.45, 265.45, 265.35, 265.25, 264.95, 
    264.75, 264.35, 263.35, 262.65, 261.75, 260.75, 261.75, 262.85, 262.35, 
    263.35, 263.95, 264.55, 265.25, 265.35, 266.05, 265.55, 266.35, 266.95, 
    266.75, 266.75, 265.85, 265.55, 264.85, 265.75, 265.65, 265.85, 266.55, 
    266.75, 265.95, 266.05, 266.05, 265.85, 266.65, 268.15, 267.95, 267.85, 
    269.25, 269.95, 270.25, 270.55, 271.25, 271.65, 271.35, 271.65, 272.35, 
    272.85, 273.45, 273.35, 273.95, 273.65, 274.45, 274.95, 276.15, 275.45, 
    275.75, 275.85, 274.95, 274.45, 273.65, 273.05, 272.45, 272.75, 272.75, 
    272.45, 272.35, 272.65, 272.55, 272.75, 273.15, 272.05, 271.35, 270.05, 
    269.35, 268.75, 268.15, 268.95, 268.75, 268.65, 268.35, 268.55, 268.85, 
    269.35, 269.65, 269.75, 270.55, 270.55, 270.65, 271.55, 270.35, 270.35, 
    271.05, 271.15, 270.25, 270.45, 270.75, 269.45, 267.95, 266.25, 266.85, 
    264.75, 265.15, 264.95, 266.65, 267.45, 268.15, 268.85, 269.85, 270.35, 
    270.45, 270.95, 271.05, 271.75, 271.95, 270.85, 270.65, 271.05, 270.85, 
    271.55, 270.85, 270.05, 269.75, 269.65, 269.65, 269.85, 269.85, 269.25, 
    268.65, 269.35, 269.55, 271.35, 271.45, 271.15, 272.15, 272.25, 271.35, 
    271.05, 271.15, 272.05, 271.25, 270.25, 270.15, 270.95, 268.65, 268.15, 
    267.65, 268.25, 266.85, 267.85, 267.25, 267.65, 269.95, 268.65, 269.45, 
    269.95, 271.15, 272.45, 272.45, 272.15, 272.45, 272.85, 272.15, 272.25, 
    272.35, 272.15, 271.75, 271.35, 271.25, 269.05, 269.25, 268.45, 267.85, 
    266.05, 265.55, 267.05, 265.95, 268.55, 267.05, 268.05, 268.15, 269.75, 
    270.05, 271.05, 271.55, 271.05, 271.55, 271.35, 271.25, 273.05, 272.35, 
    272.65, 271.65, 270.75, 270.35, 269.45, 269.85, 268.55, 267.75, 267.25, 
    268.55, 268.85, 269.75, 270.25, 270.95, 271.65, 272.25, 273.65, 274.25, 
    273.65, 273.15, 274.15, 274.85, 273.85, 273.35, 273.75, 273.55, 274.05, 
    274.05, 272.45, 272.05, 271.85, 270.45, 270.05, 268.85, 270.15, 271.05, 
    271.25, 271.85, 272.25, 272.45, 272.75, 274.25, 274.35, 274.15, 274.85, 
    274.55, 273.35, 272.65, 272.15, 272.55, 272.05, 271.45, 270.65, 269.95, 
    269.65, 267.05, 267.45, 267.65, 268.15, 270.65, 268.55, 270.65, 273.05, 
    271.55, 271.55, 272.45, 272.25, 272.85, 273.55, 273.05, 272.55, 271.85, 
    273.55, 273.45, 272.55, 270.75, 269.55, 270.05, 269.95, 267.85, 268.35, 
    269.35, 269.05, 270.95, 271.85, 271.85, 273.35, 273.15, 274.05, 274.25, 
    274.45, 273.95, 275.75, 273.75, 274.15, 274.45, 276.25, 274.45, 273.25, 
    273.25, 273.35, 273.05, 273.45, 275.15, 275.25, 275.15, 275.25, 275.25, 
    275.95, 275.75, 275.95, 275.85, 276.05, 276.35, 276.25, 275.75, 275.95, 
    275.75, 275.75, 275.65, 275.45, 275.75, 275.95, 275.95, 275.75, 275.65, 
    275.55, 275.45, 275.35, 275.35, 275.45, 275.85, 275.65, 275.45, 275.85, 
    276.05, 276.15, 276.25, 276.05, 276.15, 276.25, 276.15, 275.95, 275.75, 
    275.75, 275.95, 275.25, 274.95, 274.85, 274.05, 273.95, 273.75, 273.75, 
    273.85, 274.35, 274.65, 274.85, 276.05, 276.45, 276.45, 276.25, 276.75, 
    276.55, 276.65, 276.75, 276.55, 276.15, 275.95, 276.15, 275.85, 275.75, 
    275.65, 275.55, 276.15, 275.65, 275.75, 275.85, 275.75, 275.65, 275.55, 
    275.85, 276.05, 276.15, 275.85, 275.95, 275.75, 275.25, 275.45, 274.95, 
    273.85, 273.95, 274.55, 274.85, 274.45, 274.35, 274.15, 273.75, 273.85, 
    274.05, 274.15, 274.25, 274.45, 274.35, 274.05, 273.35, 273.75, 273.65, 
    273.95, 274.05, 274.15, 274.25, 274.25, 274.05, 273.75, 273.85, 273.35, 
    273.25, 273.05, 272.75, 272.55, 272.35, 272.25, 272.25, 272.25, 272.15, 
    272.15, 272.15, 272.25, 272.15, 272.05, 272.15, 272.45, 272.65, 272.75, 
    273.15, 273.05, 273.05, 273.25, 273.45, 273.15, 273.35, 273.35, 273.25, 
    273.25, 273.15, 272.85, 272.95, 272.05, 270.95, 271.25, 272.15, 272.35, 
    272.55, 273.45, 273.45, 273.35, 273.55, 274.05, 274.55, 274.65, 274.75, 
    274.95, 275.25, 275.45, 275.25, 275.05, 274.75, 274.85, 274.65, 274.75, 
    274.95, 274.95, 274.55, 274.75, 274.65, 275.05, 275.55, 274.25, 275.05, 
    274.95, 274.75, 273.95, 274.25, 274.55, 275.15, 275.15, 274.65, 274.65, 
    274.45, 273.95, 274.15, 273.35, 272.85, 272.95, 272.75, 271.85, 270.85, 
    272.25, 272.45, 272.25, 272.95, 273.65, 274.15, 273.95, 274.65, 275.15, 
    275.55, 275.85, 275.75, 276.15, 275.75, 275.85, 275.95, 275.95, 276.05, 
    275.95, 274.85, 274.05, 273.75, 273.35, 274.75, 274.35, 274.65, 275.35, 
    275.15, 275.35, 275.15, 275.75, 276.85, 276.05, 276.65, 277.05, 277.35, 
    276.95, 277.45, 277.65, 277.55, 277.15, 277.65, 277.75, 277.45, 276.55, 
    276.45, 276.05, 274.75, 276.15, 277.35, 277.05, 276.65, 277.75, 278.15, 
    278.45, 278.95, 278.35, 279.05, 279.55, 279.25, 278.75, 278.45, 278.55, 
    278.15, 277.95, 277.75, 277.45, 277.05, 277.05, 276.85, 276.35, 276.25, 
    276.35, 276.15, 276.15, 276.05, 276.15, 276.25, 276.45, 276.65, 276.75, 
    276.75, 277.15, 276.55, 276.85, 276.85, 276.85, 276.45, 276.55, 276.75, 
    276.35, 276.05, 275.95, 275.65, 275.75, 275.95, 276.55, 276.65, 276.55, 
    276.75, 276.75, 276.95, 277.75, 277.35, 276.85, 277.65, 277.75, 277.75, 
    278.35, 277.95, 277.35, 277.35, 277.95, 277.75, 277.45, 277.15, 277.05, 
    276.95, 276.85, 276.55, 276.75, 276.95, 276.05, 276.15, 276.35, 276.45, 
    276.15, 276.95, 277.25, 277.15, 277.15, 277.45, 277.25, 276.95, 277.05, 
    276.65, 276.35, 276.35, 275.55, 275.95, 275.75, 275.75, 276.05, 275.75, 
    275.95, 276.15, 276.35, 276.45, 276.65, 276.75, 277.05, 277.05, 277.25, 
    278.15, 277.85, 277.65, 277.55, 277.85, 277.65, 277.85, 277.75, 277.65, 
    277.55, 277.25, 277.05, 276.45, 276.75, 276.55, 276.15, 276.25, 277.05, 
    277.15, 276.75, 276.95, 276.95, 277.15, 276.65, 276.55, 277.25, 277.25, 
    277.25, 277.85, 277.25, 277.15, 277.15, 278.05, 276.85, 276.05, 275.65, 
    275.35, 275.15, 275.25, 275.95, 276.05, 275.95, 275.65, 275.75, 275.35, 
    275.55, 274.95, 275.85, 275.55, 275.75, 275.15, 275.05, 274.95, 274.55, 
    273.95, 274.35, 274.15, 274.75, 273.55, 274.15, 273.65, 273.45, 273.75, 
    274.25, 275.25, 274.55, 274.45, 275.15, 276.35, 276.85, 277.15, 277.15, 
    276.95, 276.65, 276.35, 276.45, 276.35, 276.25, 276.25, 276.15, 276.05, 
    276.05, 275.85, 275.75, 275.65, 275.75, 275.75, 276.25, 275.85, 275.35, 
    275.45, 275.65, 275.65, 276.15, 276.15, 276.35, 275.95, 275.35, 273.05, 
    272.45, 272.85, 273.85, 273.35, 274.05, 273.85, 273.85, 273.55, 271.75, 
    271.15, 270.95, 270.95, 270.85, 270.75, 270.95, 270.85, 271.65, 271.75, 
    271.75, 272.05, 271.85, 271.85, 272.35, 272.55, 272.05, 272.05, 272.25, 
    272.65, 272.95, 273.35, 273.45, 273.55, 273.55, 273.65, 272.65, 273.25, 
    273.55, 274.45, 274.35, 273.95, 274.85, 275.45, 275.85, 276.15, 276.55, 
    276.75, 277.45, 277.35, 278.05, 277.65, 277.45, 277.35, 277.25, 276.75, 
    275.35, 274.95, 274.55, 274.45, 273.85, 273.65, 273.75, 273.65, 273.95, 
    274.05, 274.25, 274.65, 275.25, 276.05, 276.25, 276.45, 276.65, 276.75, 
    276.95, 276.65, 276.65, 276.25, 276.25, 275.95, 275.65, 275.45, 275.25, 
    275.35, 274.95, 275.15, 275.05, 274.75, 274.25, 274.45, 274.75, 274.55, 
    274.85, 275.05, 275.45, 275.35, 274.35, 273.75, 273.25, 273.45, 273.35, 
    272.95, 273.05, 272.55, 272.85, 272.75, 273.15, 272.95, 273.25, 273.45, 
    273.45, 272.95, 273.25, 273.25, 273.95, 273.85, 274.35, 274.65, 274.85, 
    275.05, 275.15, 275.45, 275.45, 275.05, 275.35, 275.85, 275.65, 275.25, 
    275.25, 275.25, 274.95, 275.05, 274.65, 274.75, 274.85, 275.25, 275.35, 
    275.15, 275.85, 276.95, 276.95, 276.35, 276.55, 276.65, 277.65, 276.75, 
    277.55, 277.25, 277.05, 276.65, 276.75, 276.25, 276.05, 275.95, 275.85, 
    275.65, 275.25, 275.05, 275.15, 275.45, 275.85, 275.25, 275.85, 276.55, 
    277.05, 277.75, 278.65, 277.95, 277.65, 277.95, 278.35, 278.55, 278.25, 
    278.25, 278.25, 278.15, 278.05, 277.25, 276.95, 276.65, 276.55, 276.65, 
    277.05, 277.25, 277.35, 277.55, 278.05, 278.05, 278.65, 278.75, 278.85, 
    278.75, 278.95, 279.35, 279.35, 279.55, 279.75, 279.55, 278.95, 279.05, 
    278.95, 277.65, 277.75, 277.65, 277.55, 277.55, 277.45, 277.55, 277.55, 
    277.55, 278.05, 278.15, 277.85, 277.75, 278.15, 277.95, 277.95, 277.55, 
    278.05, 278.25, 278.55, 278.95, 278.95, 279.05, 278.95, 278.95, 278.75, 
    278.45, 278.25, 278.05, 277.75, 277.75, 278.15, 278.25, 278.15, 278.35, 
    278.55, 278.55, 278.45, 278.65, 278.95, 279.25, 279.35, 279.05, 279.55, 
    279.55, 279.75, 279.65, 279.55, 279.35, 279.15, 278.85, 278.45, 278.55, 
    278.05, 278.05, 278.35, 278.85, 279.05, 278.95, 279.35, 279.35, 279.65, 
    280.05, 279.95, 279.55, 279.45, 280.05, 279.85, 279.75, 278.95, 279.15, 
    278.85, 278.35, 278.15, 278.35, 278.15, 278.25, 278.55, 278.55, 278.95, 
    278.95, 279.05, 279.35, 279.45, 279.75, 280.05, 280.05, 280.15, 280.15, 
    279.85, 279.35, 279.05, 278.95, 279.15, 279.35, 278.75, 278.25, 278.45, 
    278.55, 278.65, 278.55, 277.85, 278.05, 277.85, 277.95, 278.15, 278.45, 
    278.95, 279.15, 280.35, 280.25, 280.45, 280.55, 280.65, 280.45, 280.75, 
    280.65, 280.05, 279.65, 279.05, 278.75, 278.75, 278.65, 278.65, 278.75, 
    279.05, 279.15, 279.15, 278.85, 279.05, 279.15, 279.35, 279.35, 279.95, 
    280.05, 280.25, 280.65, 281.05, 280.45, 280.65, 280.75, 280.95, 280.55, 
    280.35, 280.45, 280.85, 281.05, 280.55, 279.95, 280.35, 280.25, 280.25, 
    280.35, 280.05, 280.95, 280.75, 281.95, 282.75, 282.45, 283.35, 282.95, 
    282.05, 281.55, 281.35, 281.25, 281.15, 280.95, 280.95, 280.85, 280.85, 
    281.15, 280.95, 280.85, 281.15, 280.65, 281.05, 281.05, 280.75, 280.25, 
    280.35, 280.25, 280.45, 280.35, 279.55, 278.75, 278.35, 278.15, 278.55, 
    278.75, 278.85, 278.95, 278.75, 278.75, 278.65, 278.45, 278.45, 278.55, 
    278.55, 278.75, 278.95, 279.15, 279.35, 279.65, 280.45, 280.45, 280.75, 
    279.35, 280.25, 280.25, 281.25, 280.85, 280.55, 280.55, 279.95, 279.65, 
    279.55, 279.35, 279.15, 278.95, 278.45, 278.75, 278.65, 278.65, 278.85, 
    278.95, 278.95, 279.25, 280.35, 279.95, 280.65, 280.55, 280.35, 280.35, 
    280.45, 280.65, 280.55, 280.55, 280.55, 280.65, 280.35, 280.25, 280.05, 
    279.75, 279.35, 279.35, 279.35, 279.15, 278.95, 279.25, 279.35, 279.75, 
    279.85, 279.65, 279.75, 279.95, 279.95, 280.05, 280.05, 280.25, 279.75, 
    279.95, 279.45, 279.35, 279.55, 279.45, 279.35, 279.35, 279.45, 279.45, 
    279.95, 279.55, 279.35, 279.45, 279.65, 279.65, 279.95, 279.85, 280.15, 
    280.75, 280.85, 280.65, 280.65, 280.65, 280.65, 280.75, 280.85, 280.95, 
    280.55, 280.75, 280.55, 280.35, 279.85, 279.45, 279.25, 279.75, 279.85, 
    280.25, 280.25, 281.05, 282.05, 281.65, 281.95, 281.25, 281.95, 281.95, 
    281.65, 282.25, 281.75, 282.35, 282.25, 281.75, 281.55, 281.55, 280.75, 
    280.35, 279.95, 279.85, 279.45, 279.35, 279.55, 279.95, 280.25, 280.35, 
    280.15, 280.75, 280.55, 280.35, 280.15, 280.05, 280.05, 280.15, 280.25, 
    280.75, 280.45, 280.25, 280.45, 280.35, 280.45, 280.15, 280.05, 280.15, 
    280.05, 280.25, 280.55, 280.25, 280.25, 280.45, 280.25, 280.45, 280.55, 
    280.75, 281.35, 281.95, 281.45, 281.45, 281.65, 281.85, 281.95, 282.15, 
    281.85, 281.85, 281.85, 281.65, 281.35, 281.15, 281.35, 281.65, 282.35, 
    282.35, 283.25, 284.05, 283.45, 283.35, 283.45, 283.35, 283.65, 284.05, 
    284.05, 283.85, 284.35, 285.85, 285.25, 284.95, 282.65, 282.75, 281.25, 
    280.95, 280.75, 280.85, 280.85, 280.95, 281.15, 281.15, 281.65, 282.05, 
    281.65, 281.85, 281.75, 281.65, 281.45, 281.85, 281.55, 281.75, 281.75, 
    281.75, 281.45, 281.95, 281.95, 281.35, 281.35, 280.65, 280.85, 280.75, 
    280.75, 281.05, 280.95, 280.75, 280.75, 280.45, 280.75, 280.35, 280.25, 
    280.75, 280.35, 280.45, 280.35, 280.65, 280.65, 280.85, 281.25, 281.15, 
    281.05, 281.05, 280.95, 280.75, 280.75, 280.85, 280.85, 280.95, 281.05, 
    281.65, 281.45, 281.35, 281.65, 280.75, 280.55, 280.75, 280.85, 280.75, 
    280.85, 281.05, 280.75, 280.35, 280.45, 280.45, 280.35, 280.15, 280.15, 
    280.05, 279.95, 279.55, 279.35, 279.05, 278.25, 279.15, 278.35, 278.75, 
    278.75, 278.45, 278.65, 279.65, 279.95, 280.25, 280.05, 279.85, 279.85, 
    279.85, 279.65, 279.65, 279.45, 279.35, 279.45, 279.35, 279.25, 279.05, 
    278.95, 279.85, 280.15, 280.35, 280.35, 280.75, 281.75, 282.35, 283.05, 
    283.25, 282.65, 282.55, 283.65, 283.15, 283.05, 283.45, 283.15, 283.45, 
    283.05, 282.35, 281.55, 281.25, 280.75, 280.55, 280.55, 281.15, 280.75, 
    279.95, 280.15, 279.45, 279.45, 279.75, 279.35, 279.75, 280.15, 280.25, 
    280.25, 280.25, 280.35, 280.25, 280.15, 280.25, 280.05, 280.35, 280.55, 
    280.65, 279.45, 278.85, 278.85, 280.55, 281.35, 281.45, 281.55, 281.65, 
    281.85, 282.45, 282.85, 283.45, 283.55, 283.75, 284.05, 284.45, 283.95, 
    284.35, 284.05, 283.55, 283.15, 282.15, 281.95, 281.75, 281.35, 281.15, 
    280.95, 281.95, 281.95, 281.75, 282.25, 282.25, 283.25, 283.65, 284.05, 
    284.45, 285.05, 285.65, 286.35, 285.45, 285.55, 285.85, 284.65, 283.75, 
    283.85, 283.45, 283.25, 283.05, 282.55, 280.75, 280.65, 281.15, 281.05, 
    280.95, 280.95, 281.25, 281.45, 281.55, 281.55, 281.75, 281.95, 282.25, 
    282.15, 282.25, 281.95, 281.95, 282.05, 281.35, 281.25, 280.85, 281.05, 
    281.35, 281.45, 281.55, 281.65, 281.65, 281.55, 281.15, 281.55, 281.45, 
    281.55, 281.75, 281.35, 281.05, 281.35, 281.25, 281.25, 281.35, 281.55, 
    281.35, 281.15, 281.65, 281.55, 281.65, 281.55, 281.35, 281.15, 280.55, 
    280.45, 280.55, 280.45, 280.35, 280.65, 281.75, 281.35, 281.55, 281.15, 
    281.05, 280.95, 281.05, 281.25, 280.95, 280.75, 281.65, 281.25, 280.95, 
    280.65, 280.45, 280.85, 281.15, 280.75, 280.45, 280.45, 280.75, 281.15, 
    281.15, 281.05, 281.15, 281.35, 281.15, 282.45, 282.55, 283.15, 283.35, 
    284.25, 282.75, 283.45, 283.45, 282.35, 281.75, 280.85, 280.85, 280.65, 
    280.55, 280.65, 280.75, 280.25, 280.25, 280.75, 280.65, 280.65, 280.65, 
    280.85, 281.05, 281.25, 281.75, 282.05, 281.75, 280.75, 281.55, 281.55, 
    280.95, 281.05, 281.35, 281.15, 280.75, 280.65, 280.55, 280.45, 280.35, 
    279.85, 279.65, 279.85, 279.65, 279.85, 279.85, 279.75, 280.05, 280.45, 
    280.45, 280.85, 280.65, 281.15, 281.15, 281.65, 281.85, 282.15, 281.75, 
    281.35, 281.35, 281.15, 281.05, 280.85, 280.75, 280.65, 280.55, 280.55, 
    279.95, 279.85, 279.75, 280.05, 280.35, 280.35, 280.75, 280.75, 280.95, 
    281.05, 281.75, 281.55, 281.15, 281.85, 282.15, 282.35, 281.85, 281.95, 
    281.85, 281.55, 280.95, 280.95, 281.15, 281.05, 281.45, 282.25, 281.75, 
    281.85, 282.05, 282.65, 282.55, 282.45, 281.75, 282.15, 282.15, 282.35, 
    282.25, 281.95, 281.75, 281.25, 281.25, 280.75, 280.65, 280.65, 280.15, 
    279.35, 279.25, 279.55, 279.65, 279.55, 279.75, 280.05, 280.25, 280.35, 
    280.35, 280.65, 281.25, 281.75, 281.85, 282.15, 281.85, 282.35, 282.35, 
    281.85, 281.45, 281.25, 280.55, 280.05, 280.15, 279.85, 279.85, 279.95, 
    279.45, 280.05, 280.35, 280.75, 280.15, 280.75, 280.75, 280.55, 280.65, 
    280.65, 280.75, 281.35, 281.25, 281.05, 281.55, 281.55, 281.05, 280.75, 
    280.35, 279.85, 279.45, 279.55, 279.15, 279.55, 279.55, 279.45, 279.15, 
    279.05, 279.15, 279.35, 279.65, 279.35, 279.65, 279.85, 279.95, 279.75, 
    279.65, 279.25, 279.35, 279.35, 279.05, 279.05, 278.95, 279.25, 279.25, 
    279.25, 279.15, 278.65, 278.55, 278.85, 278.75, 278.35, 278.85, 279.95, 
    279.75, 279.55, 279.75, 280.05, 280.95, 281.15, 280.05, 279.85, 279.65, 
    279.75, 279.85, 279.95, 280.05, 279.95, 279.35, 279.15, 279.65, 279.45, 
    279.55, 280.65, 280.25, 280.15, 280.45, 281.55, 281.05, 280.85, 280.65, 
    280.85, 281.35, 280.85, 280.95, 280.45, 279.85, 279.95, 279.15, 278.75, 
    278.15, 277.85, 277.65, 277.55, 277.35, 277.65, 277.55, 278.25, 278.15, 
    278.35, 278.85, 279.65, 280.15, 280.35, 280.25, 280.15, 279.95, 279.85, 
    280.25, 280.05, 280.75, 279.75, 279.25, 278.15, 278.25, 277.15, 276.15, 
    276.55, 276.65, 276.75, 276.55, 277.05, 277.45, 278.15, 278.15, 278.15, 
    278.25, 278.35, 278.85, 278.65, 278.25, 277.95, 277.85, 277.85, 277.65, 
    277.45, 277.35, 277.25, 277.15, 276.95, 276.15, 275.95, 275.75, 276.45, 
    276.75, 277.25, 277.85, 278.05, 278.15, 278.75, 278.15, 278.15, 278.15, 
    278.55, 278.35, 278.45, 278.55, 278.25, 278.15, 278.05, 278.05, 277.45, 
    277.55, 277.45, 277.35, 277.25, 277.35, 277.65, 277.75, 278.25, 279.25, 
    278.55, 279.05, 279.25, 279.75, 279.95, 280.25, 280.45, 280.55, 280.35, 
    280.35, 279.95, 279.55, 278.85, 278.25, 277.45, 276.95, 276.65, 276.35, 
    276.35, 276.75, 277.15, 277.95, 278.05, 278.95, 279.75, 280.35, 280.95, 
    281.45, 281.95, 282.35, 282.75, 282.75, 282.55, 282.15, 281.45, 280.45, 
    279.45, 278.55, 277.65, 277.05, 277.15, 277.15, 277.05, 277.35, 277.65, 
    278.05, 279.85, 280.45, 282.85, 283.05, 281.45, 283.95, 284.25, 282.45, 
    282.45, 282.35, 282.05, 281.55, 280.75, 279.85, 279.05, 278.35, 277.55, 
    276.75, 276.05, 275.65, 275.25, 275.25, 275.45, 275.95, 277.25, 278.35, 
    282.45, 281.85, 281.65, 282.25, 282.15, 282.15, 282.15, 282.15, 282.05, 
    281.55, 281.55, 281.35, 281.05, 280.75, 280.65, 279.85, 279.75, 279.65, 
    279.65, 279.65, 279.85, 279.75, 279.85, 280.25, 279.75, 280.25, 280.25, 
    280.25, 280.85, 281.35, 281.15, 281.35, 282.25, 282.55, 282.25, 281.75, 
    281.25, 280.95, 280.85, 280.45, 280.45, 280.35, 280.35, 280.55, 280.45, 
    280.95, 281.15, 281.15, 281.05, 280.55, 280.75, 281.05, 280.85, 280.85, 
    280.75, 280.85, 281.05, 281.05, 281.25, 281.15, 280.75, 280.55, 280.25, 
    280.15, 279.95, 279.85, 279.65, 279.55, 279.35, 279.15, 279.65, 279.45, 
    279.65, 279.15, 279.25, 279.55, 280.05, 279.65, 279.65, 279.35, 279.55, 
    279.65, 279.55, 279.55, 279.55, 279.55, 279.55, 279.55, 279.55, 279.55, 
    279.75, 279.85, 279.95, 280.05, 280.05, 280.05, 280.05, 279.15, 279.35, 
    279.65, 279.85, 280.05, 280.05, 279.95, 280.05, 279.85, 280.35, 280.25, 
    280.55, 280.55, 280.45, 279.85, 279.65, 279.95, 279.65, 279.95, 280.05, 
    280.05, 280.15, 280.15, 280.15, 280.25, 280.35, 280.35, 280.55, 280.65, 
    280.75, 280.75, 281.15, 280.95, 280.75, 280.65, 280.55, 280.35, 280.25, 
    280.15, 279.95, 279.85, 279.65, 279.55, 280.15, 279.55, 279.85, 280.15, 
    280.25, 280.65, 281.75, 280.85, 280.75, 281.85, 281.55, 281.15, 280.85, 
    280.55, 280.15, 279.85, 279.85, 279.85, 279.85, 279.85, 279.55, 279.55, 
    279.65, 279.15, 279.25, 279.75, 279.85, 280.25, 280.75, 280.65, 280.55, 
    280.75, 281.35, 281.25, 281.95, 281.55, 281.35, 281.25, 281.25, 281.15, 
    280.95, 280.95, 280.75, 280.65, 280.65, 280.75, 280.75, 280.85, 280.85, 
    280.95, 280.95, 281.05, 281.05, 281.05, 281.15, 281.15, 281.65, 281.35, 
    281.55, 281.65, 281.55, 281.45, 280.85, 280.85, 280.75, 280.45, 280.15, 
    279.95, 279.35, 279.25, 279.05, 278.75, 279.35, 279.75, 280.05, 281.25, 
    281.75, 281.95, 282.65, 282.35, 282.65, 282.65, 282.25, 281.75, 281.25, 
    280.55, 279.75, 279.05, 278.85, 278.65, 278.15, 277.75, 277.75, 277.65, 
    277.45, 277.05, 277.45, 277.55, 277.95, 278.75, 280.15, 280.45, 279.75, 
    281.05, 280.95, 280.75, 280.65, 280.35, 279.95, 279.65, 279.55, 279.25, 
    278.35, 278.25, 278.15, 278.05, 277.85, 277.45, 277.75, 277.75, 277.75, 
    278.15, 278.05, 278.55, 279.75, 281.15, 280.25, 279.55, 279.65, 280.25, 
    280.35, 279.55, 280.25, 279.65, 279.45, 278.85, 278.25, 278.05, 277.35, 
    276.75, 276.35, 276.75, 276.25, 276.25, 276.75, 276.95, 277.15, 277.45, 
    278.95, 278.85, 279.35, 280.05, 280.25, 281.15, 281.05, 280.75, 280.35, 
    280.05, 279.85, 279.75, 279.55, 279.25, 278.75, 278.65, 278.15, 278.85, 
    278.45, 278.65, 278.95, 279.25, 279.45, 279.85, 280.25, 280.65, 280.95, 
    280.95, 280.95, 280.95, 281.15, 280.95, 280.65, 280.15, 279.75, 279.35, 
    278.95, 278.55, 278.15, 277.75, 277.35, 276.95, 276.55, 276.45, 277.35, 
    277.35, 278.05, 278.75, 278.15, 279.05, 279.05, 278.85, 278.95, 278.95, 
    278.55, 278.45, 278.05, 277.65, 277.25, 276.85, 276.65, 276.35, 276.05, 
    275.65, 275.35, 275.05, 274.75, 274.15, 274.65, 275.35, 276.15, 276.95, 
    277.75, 278.55, 279.25, 279.95, 280.85, 280.75, 280.45, 280.55, 280.75, 
    280.65, 280.95, 279.35, 278.25, 277.15, 276.45, 276.15, 275.45, 274.95, 
    274.55, 274.05, 274.75, 275.15, 275.85, 276.75, 277.05, 277.85, 277.75, 
    278.05, 278.55, 279.15, 279.25, 279.05, 279.05, 278.75, 279.05, 278.25, 
    277.55, 277.15, 276.75, 276.45, 276.25, 275.95, 275.85, 276.55, 276.35, 
    276.25, 276.55, 276.75, 277.35, 278.25, 279.35, 280.75, 280.15, 280.75, 
    280.35, 279.95, 279.55, 279.15, 278.65, 278.25, 277.85, 277.45, 277.05, 
    276.65, 276.65, 277.15, 277.05, 276.45, 276.55, 276.75, 277.05, 277.45, 
    277.85, 278.15, 278.55, 279.45, 279.75, 279.95, 279.95, 279.75, 279.05, 
    278.55, 278.15, 277.65, 277.15, 276.85, 276.25, 275.45, 275.25, 275.15, 
    274.45, 275.05, 274.95, 275.15, 275.95, 276.95, 278.15, 279.35, 280.45, 
    280.85, 280.85, 280.25, 280.15, 279.45, 278.85, 278.25, 278.85, 278.05, 
    277.05, 276.05, 274.85, 273.85, 273.65, 273.55, 274.45, 275.05, 275.55, 
    275.15, 276.25, 277.35, 277.35, 277.55, 277.85, 278.15, 278.35, 278.75, 
    279.35, 279.25, 279.45, 279.55, 279.25, 277.85, 276.75, 275.85, 275.35, 
    276.15, 276.15, 275.55, 275.85, 276.25, 276.55, 277.25, 277.15, 277.25, 
    277.35, 277.45, 278.35, 278.65, 279.25, 278.55, 278.65, 279.35, 278.75, 
    279.05, 279.05, 277.75, 276.95, 276.55, 276.05, 275.35, 274.75, 273.95, 
    273.55, 274.25, 274.25, 275.45, 275.75, 277.25, 277.05, 277.05, 277.35, 
    277.55, 277.55, 277.65, 277.95, 278.25, 278.25, 278.35, 278.55, 278.25, 
    277.35, 277.75, 277.55, 278.45, 278.15, 277.85, 277.95, 277.75, 277.65, 
    277.75, 277.95, 277.75, 277.75, 277.85, 277.95, 277.95, 278.25, 278.75, 
    279.25, 280.45, 280.35, 279.85, 279.65, 279.45, 278.95, 278.45, 278.65, 
    278.15, 278.65, 278.05, 277.55, 277.35, 277.25, 277.15, 277.25, 277.15, 
    277.05, 276.95, 276.95, 276.95, 277.05, 277.25, 276.75, 276.75, 276.75, 
    276.45, 276.55, 276.35, 276.15, 275.95, 276.15, 275.65, 275.45, 275.85, 
    275.45, 275.55, 275.35, 275.85, 276.45, 276.65, 277.15, 276.85, 277.05, 
    277.35, 277.55, 276.75, 277.35, 277.65, 277.55, 277.25, 276.95, 276.45, 
    276.75, 275.95, 275.95, 275.25, 274.75, 274.15, 275.45, 275.75, 276.05, 
    275.95, 276.95, 276.95, 277.05, 277.45, 278.05, 277.65, 277.55, 278.05, 
    277.25, 277.05, 276.75, 276.85, 276.45, 276.15, 276.05, 275.95, 275.75, 
    275.95, 275.55, 275.55, 275.65, 274.95, 274.45, 274.65, 275.05, 277.05, 
    276.75, 276.65, 275.95, 276.35, 276.65, 277.15, 276.65, 277.05, 276.85, 
    276.65, 276.35, 276.05, 275.75, 274.65, 273.65, 272.75, 273.45, 273.25, 
    273.65, 273.95, 273.95, 274.65, 274.75, 275.05, 276.15, 277.05, 277.25, 
    277.45, 277.55, 277.15, 277.35, 277.25, 276.95, 276.65, 276.65, 276.25, 
    275.65, 275.25, 275.15, 275.25, 275.15, 275.05, 274.65, 274.55, 275.25, 
    275.05, 275.45, 275.75, 276.15, 276.45, 276.35, 276.65, 277.05, 276.85, 
    277.05, 276.85, 276.75, 276.75, 276.75, 276.65, 276.55, 276.45, 276.45, 
    276.35, 276.45, 276.45, 276.55, 276.85, 276.75, 276.85, 276.75, 276.95, 
    277.45, 277.85, 277.85, 277.75, 277.75, 277.85, 277.75, 277.55, 277.45, 
    277.15, 277.05, 276.95, 276.85, 276.55, 276.55, 276.45, 276.25, 276.35, 
    276.35, 276.35, 276.45, 276.45, 276.65, 276.65, 276.95, 277.05, 277.15, 
    277.25, 277.35, 278.15, 278.05, 277.85, 277.75, 277.55, 277.45, 277.25, 
    277.15, 277.05, 276.55, 276.45, 276.05, 275.95, 275.95, 276.25, 276.45, 
    276.65, 276.95, 277.25, 277.45, 277.75, 278.35, 278.35, 278.15, 278.45, 
    278.35, 278.15, 277.65, 277.55, 277.35, 277.25, 277.05, 276.85, 276.85, 
    276.65, 276.55, 275.55, 275.35, 274.95, 273.95, 273.75, 273.85, 273.75, 
    273.65, 273.55, 273.45, 273.45, 273.45, 273.25, 273.65, 273.45, 273.55, 
    273.25, 272.05, 272.05, 271.75, 271.35, 271.05, 270.65, 270.05, 270.65, 
    270.35, 270.85, 270.75, 271.55, 271.75, 272.25, 272.65, 272.95, 273.25, 
    273.15, 272.65, 273.15, 273.25, 273.15, 273.15, 273.25, 273.45, 273.55, 
    273.35, 273.35, 273.45, 274.25, 273.35, 273.25, 273.35, 273.55, 273.85, 
    274.85, 274.85, 275.15, 275.25, 275.45, 275.45, 275.45, 275.45, 275.45, 
    275.35, 275.35, 275.15, 275.05, 274.75, 274.35, 274.25, 274.15, 274.05, 
    273.95, 273.75, 273.65, 273.55, 273.45, 273.35, 273.55, 273.75, 273.95, 
    274.35, 274.75, 275.15, 275.25, 275.15, 275.05, 274.95, 275.05, 274.85, 
    274.55, 274.25, 274.55, 274.45, 274.35, 274.25, 274.15, 274.15, 274.05, 
    273.95, 273.85, 273.75, 273.65, 273.65, 273.95, 274.15, 274.55, 274.75, 
    274.95, 274.95, 274.85, 274.85, 274.95, 274.85, 274.95, 275.05, 274.75, 
    274.85, 275.25, 275.15, 274.85, 274.85, 274.55, 274.25, 274.05, 273.65, 
    273.75, 274.55, 274.95, 275.15, 275.25, 275.65, 275.75, 275.75, 275.55, 
    275.25, 274.85, 274.85, 274.25, 274.35, 274.65, 274.75, 274.95, 275.05, 
    275.45, 275.65, 276.05, 278.45, 277.75, 277.15, 277.05, 277.65, 277.85, 
    278.05, 277.95, 278.45, 279.15, 278.45, 278.45, 279.05, 279.35, 278.95, 
    278.55, 278.15, 277.75, 277.15, 276.85, 276.75, 276.55, 276.45, 276.35, 
    275.45, 274.95, 274.85, 274.85, 274.45, 274.45, 274.15, 274.35, 273.95, 
    273.85, 274.35, 274.05, 273.55, 273.85, 273.65, 273.65, 273.65, 273.55, 
    273.55, 273.35, 272.95, 272.75, 272.75, 272.65, 272.15, 272.85, 272.45, 
    271.85, 272.35, 273.35, 273.95, 273.85, 274.55, 274.65, 274.45, 275.95, 
    275.15, 275.35, 274.55, 274.45, 274.55, 274.75, 274.85, 275.05, 275.15, 
    275.05, 275.25, 274.65, 274.75, 274.65, 274.65, 274.85, 275.15, 275.25, 
    275.35, 275.35, 275.35, 275.85, 275.65, 275.95, 277.55, 278.55, 280.75, 
    279.45, 279.15, 278.95, 279.05, 279.95, 278.85, 278.65, 278.55, 278.65, 
    278.35, 277.05, 275.75, 275.75, 275.25, 274.75, 274.15, 273.45, 272.95, 
    272.85, 273.05, 272.35, 272.65, 272.45, 271.95, 271.55, 271.35, 271.25, 
    271.55, 271.45, 271.75, 271.55, 271.55, 271.95, 271.95, 271.25, 271.45, 
    271.75, 271.95, 272.05, 272.25, 272.75, 272.35, 272.85, 272.35, 272.85, 
    272.75, 272.55, 272.35, 272.25, 272.05, 271.95, 271.75, 271.55, 271.45, 
    271.35, 271.35, 271.75, 271.65, 272.35, 271.95, 272.05, 272.25, 272.45, 
    272.55, 272.75, 272.75, 272.85, 272.55, 272.75, 272.15, 272.35, 272.05, 
    271.85, 271.85, 271.65, 271.55, 271.55, 271.35, 270.85, 270.35, 270.45, 
    270.55, 270.45, 270.35, 270.25, 270.15, 270.05, 270.05, 271.25, 272.05, 
    271.95, 271.75, 272.05, 272.35, 272.55, 272.55, 272.25, 271.95, 271.95, 
    271.95, 272.05, 271.65, 271.95, 271.95, 271.85, 271.75, 269.95, 270.75, 
    271.05, 270.75, 271.45, 271.75, 272.05, 272.35, 272.65, 272.85, 273.15, 
    273.45, 273.75, 274.05, 272.55, 272.25, 271.65, 271.55, 271.65, 271.75, 
    271.65, 271.35, 271.05, 270.85, 270.55, 270.45, 270.65, 271.15, 271.45, 
    271.75, 272.65, 272.85, 272.85, 272.95, 272.95, 273.05, 273.05, 273.05, 
    273.35, 273.25, 273.05, 272.95, 273.35, 273.15, 273.05, 272.85, 272.75, 
    272.65, 272.45, 273.35, 273.45, 274.05, 274.65, 275.15, 275.35, 275.55, 
    275.65, 275.65, 275.55, 275.65, 275.65, 275.75, 275.85, 275.95, 276.45, 
    276.55, 276.45, 276.35, 275.95, 276.05, 276.15, 276.15, 276.25, 276.25, 
    276.25, 276.55, 276.35, 276.95, 276.95, 276.95, 276.95, 276.95, 276.45, 
    276.45, 276.75, 276.55, 276.35, 275.55, 276.45, 276.55, 276.15, 276.05, 
    275.85, 275.95, 275.55, 274.75, 275.25, 275.75, 274.75, 275.15, 275.05, 
    275.05, 275.15, 275.35, 275.65, 275.85, 275.55, 274.95, 274.85, 274.95, 
    275.15, 275.35, 275.65, 275.85, 275.25, 274.95, 275.55, 275.65, 275.65, 
    275.75, 275.75, 275.55, 276.25, 276.85, 276.65, 276.35, 276.65, 276.85, 
    276.45, 276.35, 276.45, 275.95, 275.75, 275.55, 275.95, 275.45, 274.95, 
    274.65, 274.45, 274.35, 274.45, 275.05, 275.65, 276.05, 276.35, 276.55, 
    275.05, 275.45, 275.15, 275.65, 276.05, 276.15, 276.15, 275.95, 275.65, 
    275.25, 274.75, 274.25, 273.85, 273.85, 273.75, 273.25, 272.65, 272.05, 
    271.75, 271.65, 271.55, 270.65, 270.25, 270.05, 269.15, 270.75, 270.35, 
    270.65, 270.95, 271.15, 271.45, 271.75, 271.95, 271.75, 271.45, 271.55, 
    271.45, 271.25, 271.15, 270.95, 270.75, 270.55, 270.35, 270.05, 270.65, 
    270.75, 270.75, 270.65, 270.45, 270.85, 271.05, 271.25, 271.25, 271.45, 
    271.55, 271.65, 271.45, 271.15, 271.05, 270.75, 270.55, 270.35, 270.25, 
    270.25, 270.35, 270.65, 270.45, 270.15, 269.75, 269.55, 269.25, 268.95, 
    268.55, 268.35, 268.75, 268.95, 269.05, 269.25, 269.55, 269.65, 270.35, 
    270.05, 269.45, 268.95, 268.55, 268.45, 268.45, 268.65, 268.55, 268.45, 
    268.35, 268.15, 267.95, 267.65, 267.35, 267.15, 266.85, 266.55, 266.35, 
    266.05, 266.05, 267.55, 267.15, 266.75, 267.55, 267.75, 268.85, 269.55, 
    270.65, 270.35, 270.85, 272.45, 273.85, 274.25, 274.65, 275.05, 275.45, 
    275.95, 276.35, 275.05, 275.35, 275.65, 275.85, 275.45, 276.15, 275.95, 
    275.65, 275.75, 275.15, 275.05, 274.95, 274.95, 274.85, 274.75, 274.65, 
    274.85, 274.75, 274.95, 275.75, 276.35, 276.65, 276.25, 276.45, 276.15, 
    275.45, 276.05, 275.85, 275.55, 275.35, 275.45, 275.75, 276.05, 275.65, 
    275.45, 276.65, 277.15, 276.55, 277.45, 278.35, 278.35, 278.35, 278.45, 
    278.75, 279.05, 279.45, 279.85, 279.95, 279.85, 279.65, 279.15, 278.55, 
    278.05, 278.85, 278.25, 278.75, 278.95, 279.35, 277.75, 277.15, 277.05, 
    276.65, 276.05, 275.75, 276.05, 276.65, 277.15, 277.35, 277.25, 277.15, 
    277.95, 277.95, 277.35, 277.05, 276.75, 276.45, 276.05, 275.75, 275.45, 
    275.15, 275.05, 274.55, 273.85, 273.75, 274.85, 275.15, 275.45, 276.55, 
    275.65, 275.95, 275.65, 275.35, 275.45, 275.85, 276.25, 276.25, 276.05, 
    275.75, 275.45, 275.15, 274.85, 274.55, 274.25, 273.95, 273.65, 273.35, 
    273.15, 273.15, 272.95, 272.65, 272.45, 272.35, 272.75, 273.15, 272.95, 
    272.65, 272.15, 271.55, 271.15, 270.95, 270.85, 270.85, 270.65, 270.25, 
    270.15, 270.55, 271.15, 270.85, 270.35, 270.65, 269.45, 268.45, 270.25, 
    270.35, 270.65, 269.35, 268.95, 269.15, 269.05, 268.95, 269.05, 268.75, 
    267.65, 268.15, 268.55, 267.55, 267.65, 267.35, 267.35, 267.95, 267.85, 
    267.95, 268.25, 268.05, 267.35, 267.45, 266.75, 267.15, 267.65, 267.35, 
    268.05, 268.45, 268.75, 269.05, 268.95, 268.75, 269.05, 269.25, 269.25, 
    269.05, 269.05, 268.85, 268.55, 268.95, 269.25, 269.45, 269.55, 269.55, 
    269.55, 269.45, 269.65, 269.85, 270.05, 270.05, 270.25, 270.45, 270.45, 
    270.25, 270.15, 270.55, 270.45, 270.55, 270.45, 270.55, 270.95, 270.85, 
    270.55, 270.25, 270.15, 270.55, 270.85, 271.15, 271.55, 271.35, 270.95, 
    270.85, 270.75, 270.35, 270.75, 270.55, 270.45, 270.35, 270.45, 269.35, 
    269.05, 269.55, 270.15, 270.95, 271.15, 270.95, 271.05, 270.75, 270.75, 
    270.85, 270.05, 269.85, 269.65, 269.05, 268.25, 267.65, 267.45, 267.65, 
    268.05, 268.65, 269.15, 269.15, 269.05, 269.15, 268.35, 268.55, 268.15, 
    268.65, 268.65, 268.75, 268.35, 268.35, 268.55, 268.65, 268.45, 268.25, 
    268.55, 267.15, 268.05, 268.35, 268.55, 268.65, 268.75, 269.25, 268.15, 
    267.55, 266.85, 264.45, 264.95, 265.75, 265.05, 264.95, 264.95, 265.25, 
    265.95, 266.65, 266.85, 266.35, 266.45, 266.35, 266.35, 266.15, 265.85, 
    265.45, 264.75, 265.15, 265.05, 265.35, 264.55, 264.25, 263.85, 263.75, 
    263.85, 264.15, 264.25, 264.65, 265.75, 265.55, 265.15, 265.35, 265.55, 
    265.45, 263.35, 263.25, 264.05, 264.85, 265.55, 266.35, 266.75, 266.55, 
    266.35, 265.95, 265.55, 264.95, 264.85, 264.05, 263.25, 262.45, 261.75, 
    261.55, 260.05, 260.85, 260.05, 261.75, 261.05, 261.25, 261.35, 260.75, 
    260.95, 260.35, 260.55, 260.45, 260.05, 259.55, 259.15, 259.35, 260.95, 
    261.75, 262.85, 263.55, 263.55, 264.25, 264.75, 264.75, 265.35, 265.35, 
    265.25, 265.35, 265.65, 265.95, 265.75, 265.95, 266.75, 266.95, 266.85, 
    266.85, 266.65, 266.65, 266.65, 266.65, 266.65, 266.75, 267.15, 267.25, 
    267.25, 267.35, 267.05, 267.15, 266.85, 266.85, 266.75, 265.05, 264.75, 
    263.75, 262.75, 262.65, 262.85, 262.85, 262.85, 262.75, 262.75, 262.65, 
    262.65, 261.75, 261.45, 261.85, 262.15, 262.35, 262.15, 262.45, 262.65, 
    262.85, 263.05, 263.15, 262.55, 263.65, 264.25, 264.25, 264.15, 262.85, 
    262.05, 261.85, 262.15, 262.25, 262.25, 262.35, 262.45, 262.45, 262.55, 
    262.45, 262.65, 262.95, 263.95, 264.05, 264.25, 264.65, 264.65, 264.85, 
    265.05, 265.45, 265.55, 265.65, 265.85, 266.15, 266.35, 266.25, 266.25, 
    266.55, 266.75, 266.85, 267.05, 267.05, 267.35, 267.75, 268.15, 267.55, 
    268.05, 268.05, 268.15, 268.45, 268.45, 268.05, 267.55, 266.45, 267.55, 
    267.45, 267.45, 267.55, 266.85, 266.85, 267.15, 267.25, 267.15, 266.85, 
    266.85, 267.25, 265.95, 266.75, 266.45, 267.65, 268.25, 267.35, 266.85, 
    266.65, 267.55, 268.65, 266.55, 267.55, 268.35, 267.65, 266.05, 266.15, 
    266.55, 266.95, 267.45, 267.85, 268.35, 268.85, 269.35, 269.85, 270.35, 
    270.25, 270.85, 272.25, 271.85, 272.25, 272.75, 272.95, 273.05, 273.25, 
    273.75, 274.05, 274.55, 274.75, 274.45, 274.65, 274.25, 274.35, 273.85, 
    274.35, 273.35, 273.35, 273.35, 273.45, 273.45, 273.45, 273.45, 273.45, 
    273.55, 273.45, 273.55, 273.65, 273.05, 273.75, 276.55, 274.85, 277.45, 
    276.15, 277.15, 276.85, 276.55, 276.15, 275.65, 274.75, 275.25, 274.15, 
    274.25, 275.85, 272.45, 272.85, 273.85, 274.55, 275.75, 275.95, 275.75, 
    275.45, 275.15, 275.35, 274.85, 275.35, 275.25, 274.45, 274.85, 275.45, 
    276.05, 276.75, 277.35, 277.95, 278.35, 277.85, 277.95, 277.65, 277.35, 
    277.05, 276.75, 275.95, 275.45, 275.45, 275.65, 275.95, 275.75, 275.65, 
    276.55, 276.45, 275.95, 275.85, 276.95, 279.05, 279.75, 278.75, 278.65, 
    278.55, 276.95, 276.85, 277.45, 278.25, 278.65, 277.55, 277.65, 276.85, 
    277.15, 276.65, 277.05, 276.85, 276.85, 276.75, 276.65, 276.55, 276.85, 
    276.45, 276.75, 276.95, 276.65, 276.55, 276.55, 276.45, 276.35, 275.95, 
    276.05, 276.65, 277.15, 277.15, 277.45, 276.85, 276.85, 276.75, 276.65, 
    276.55, 276.45, 276.35, 276.65, 276.65, 276.75, 276.85, 276.25, 276.05, 
    275.85, 275.65, 275.65, 275.65, 275.55, 275.45, 275.35, 275.15, 275.15, 
    275.15, 274.95, 274.95, 274.85, 274.75, 274.75, 274.65, 274.45, 274.35, 
    274.05, 273.95, 273.65, 273.95, 273.85, 273.55, 273.45, 273.35, 273.15, 
    272.95, 272.85, 272.75, 272.65, 272.45, 272.25, 272.15, 271.95, 271.75, 
    271.65, 271.45, 271.25, 271.45, 271.55, 271.35, 271.55, 271.25, 271.25, 
    270.85, 270.55, 270.15, 270.15, 269.45, 269.55, 269.95, 270.05, 269.55, 
    269.45, 269.25, 269.25, 269.15, 269.05, 268.95, 268.75, 268.65, 268.65, 
    268.25, 267.95, 265.15, 265.15, 265.35, 265.25, 265.95, 266.15, 266.35, 
    266.85, 267.25, 267.15, 267.05, 267.25, 267.35, 267.35, 267.75, 267.75, 
    267.95, 267.75, 267.95, 268.75, 268.55, 267.95, 267.35, 266.25, 266.55, 
    267.05, 266.95, 267.25, 266.95, 267.25, 267.05, 267.25, 267.45, 267.75, 
    267.85, 268.05, 268.05, 268.35, 268.25, 268.25, 268.35, 267.95, 267.05, 
    267.75, 266.55, 265.45, 265.85, 265.45, 265.25, 265.25, 265.45, 265.45, 
    265.75, 265.85, 265.55, 265.25, 265.15, 265.15, 265.75, 265.65, 265.55, 
    265.45, 265.65, 265.35, 265.35, 265.25, 264.75, 264.75, 264.15, 263.55, 
    264.05, 264.25, 264.05, 264.45, 265.05, 264.95, 265.05, 264.95, 264.85, 
    264.55, 263.85, 263.55, 263.35, 263.15, 263.15, 262.95, 262.65, 262.65, 
    262.55, 261.75, 262.15, 261.95, 261.55, 261.25, 261.05, 260.25, 259.65, 
    259.35, 259.45, 259.35, 259.45, 259.55, 258.95, 259.35, 259.45, 259.95, 
    258.95, 259.35, 260.35, 258.35, 259.15, 257.05, 257.25, 256.65, 257.05, 
    257.55, 257.25, 257.15, 257.35, 256.95, 256.25, 258.15, 258.55, 259.25, 
    259.45, 259.75, 259.95, 259.65, 259.75, 259.95, 259.65, 259.75, 260.05, 
    260.25, 260.45, 260.75, 260.95, 261.05, 261.15, 261.25, 261.45, 261.25, 
    260.15, 260.75, 260.65, 260.65, 261.05, 261.85, 262.45, 263.45, 260.95, 
    261.75, 261.75, 262.25, 260.55, 259.45, 261.25, 259.55, 259.95, 259.05, 
    259.25, 259.75, 259.45, 258.95, 259.15, 258.85, 258.65, 258.15, 258.55, 
    258.45, 259.25, 259.45, 259.05, 258.95, 259.15, 259.25, 259.55, 259.85, 
    260.15, 260.55, 261.35, 261.25, 261.35, 262.05, 262.75, 264.25, 263.45, 
    264.85, 265.05, 265.25, 265.45, 265.95, 266.45, 266.35, 266.65, 267.05, 
    266.45, 266.15, 266.35, 266.45, 266.75, 268.05, 269.45, 269.85, 268.55, 
    268.55, 270.05, 269.25, 269.05, 268.95, 267.95, 267.55, 267.35, 266.55, 
    267.45, 267.85, 267.95, 267.25, 267.55, 266.85, 266.25, 265.55, 265.55, 
    265.35, 265.25, 265.25, 265.65, 265.65, 265.35, 265.45, 265.35, 265.05, 
    264.75, 264.55, 264.65, 264.35, 264.35, 264.35, 264.15, 263.85, 263.65, 
    263.65, 264.05, 263.75, 264.15, 263.55, 263.25, 263.25, 262.85, 262.55, 
    262.45, 262.05, 262.35, 261.65, 261.35, 261.25, 260.25, 260.85, 259.85, 
    257.95, 258.95, 258.95, 259.45, 259.05, 259.15, 258.85, 259.15, 257.85, 
    257.75, 258.65, 256.65, 258.55, 258.15, 258.65, 258.55, 257.75, 257.45, 
    257.55, 258.25, 257.25, 258.85, 258.95, 260.15, 258.75, 257.85, 259.65, 
    259.75, 259.25, 259.85, 259.65, 258.95, 256.95, 256.55, 257.05, 257.95, 
    257.15, 258.05, 258.55, 258.15, 258.35, 258.55, 258.75, 258.65, 258.45, 
    258.15, 257.25, 258.15, 257.45, 258.45, 258.45, 256.55, 257.95, 258.55, 
    257.15, 258.35, 258.05, 258.45, 258.25, 258.35, 258.45, 258.15, 258.75, 
    259.05, 258.95, 259.85, 259.55, 258.65, 257.65, 258.05, 259.05, 259.55, 
    258.05, 258.15, 258.45, 257.75, 257.65, 258.75, 257.75, 257.75, 257.05, 
    257.35, 257.65, 258.25, 257.45, 256.65, 257.85, 259.25, 257.85, 257.65, 
    257.85, 259.05, 258.65, 259.75, 259.95, 259.25, 258.65, 259.05, 257.35, 
    259.05, 258.75, 259.95, 260.05, 260.55, 260.75, 261.45, 261.05, 261.95, 
    261.35, 261.35, 262.35, 262.15, 262.65, 262.65, 262.45, 262.85, 263.25, 
    263.55, 264.15, 264.55, 266.85, 271.85, 272.75, 274.55, 273.65, 273.75, 
    275.25, 275.05, 274.85, 274.75, 273.45, 273.05, 271.95, 271.15, 270.35, 
    266.85, 266.45, 265.95, 264.95, 264.45, 263.85, 262.65, 262.75, 262.15, 
    261.85, 260.45, 259.75, 261.15, 260.65, 259.55, 258.45, 259.35, 260.05, 
    259.65, 259.15, 259.15, 259.35, 259.95, 259.25, 258.35, 260.15, 259.65, 
    259.85, 260.15, 261.05, 261.55, 262.65, 263.35, 263.85, 263.85, 263.45, 
    263.15, 263.95, 264.55, 264.45, 264.75, 265.25, 266.05, 266.05, 267.25, 
    267.05, 267.65, 267.95, 269.25, 269.45, 269.55, 268.85, 268.85, 268.55, 
    268.45, 268.45, 268.55, 268.55, 269.15, 268.35, 267.95, 268.05, 268.55, 
    267.95, 267.85, 268.65, 268.15, 267.75, 268.15, 267.95, 267.65, 267.25, 
    266.95, 266.75, 267.05, 266.85, 266.35, 266.75, 267.15, 266.75, 266.65, 
    266.55, 266.05, 266.05, 266.05, 265.45, 265.85, 265.55, 265.15, 264.75, 
    263.55, 262.65, 262.85, 261.85, 261.15, 259.95, 259.75, 258.95, 256.45, 
    255.15, 254.75, 254.55, 253.45, 255.65, 253.65, 254.25, 254.35, 254.45, 
    255.45, 256.75, 256.45, 257.15, 257.35, 257.55, 256.95, 256.65, 259.05, 
    260.35, 260.65, 260.75, 260.45, 262.35, 262.25, 262.65, 262.65, 262.85, 
    262.25, 262.35, 262.55, 262.65, 262.95, 263.55, 263.75, 264.05, 264.65, 
    265.45, 265.35, 265.45, 265.95, 266.65, 265.85, 265.95, 266.25, 266.45, 
    266.35, 266.45, 267.65, 267.45, 268.45, 269.15, 269.05, 269.55, 268.95, 
    268.95, 268.95, 269.25, 269.15, 269.55, 270.05, 270.65, 271.55, 272.75, 
    275.25, 275.75, 275.25, 275.65, 274.95, 274.85, 274.75, 274.75, 275.05, 
    275.35, 275.75, 275.55, 275.65, 275.75, 275.45, 275.25, 275.35, 275.25, 
    275.35, 275.45, 275.05, 275.45, 275.55, 276.15, 276.35, 275.55, 276.35, 
    275.75, 276.45, 276.05, 276.25, 276.45, 275.75, 275.65, 275.55, 274.65, 
    273.05, 271.05, 269.05, 268.15, 267.05, 266.65, 266.45, 265.05, 263.45, 
    262.85, 262.25, 262.05, 262.75, 263.55, 264.25, 264.15, 264.25, 264.45, 
    265.15, 265.65, 265.95, 266.35, 265.95, 266.25, 266.85, 267.45, 267.65, 
    267.55, 267.85, 268.25, 268.75, 268.95, 269.05, 269.15, 269.65, 269.25, 
    270.55, 270.45, 270.45, 270.75, 271.05, 271.15, 271.65, 271.75, 271.75, 
    271.65, 272.25, 272.25, 272.15, 272.15, 272.25, 271.85, 272.25, 272.35, 
    272.35, 273.65, 273.55, 273.55, 273.75, 273.25, 273.55, 271.95, 271.95, 
    271.95, 272.15, 272.35, 272.15, 272.45, 272.15, 272.45, 271.95, 271.75, 
    272.05, 271.85, 272.15, 272.45, 271.85, 272.15, 272.35, 272.45, 272.65, 
    272.95, 272.35, 273.95, 276.55, 276.25, 275.45, 275.05, 274.45, 273.85, 
    275.25, 274.55, 273.95, 272.75, 272.25, 269.85, 271.55, 269.85, 269.75, 
    269.95, 270.15, 270.55, 270.55, 270.25, 269.75, 269.15, 268.55, 270.35, 
    270.55, 270.15, 269.55, 268.45, 269.95, 270.45, 270.15, 268.45, 266.35, 
    266.45, 264.95, 263.95, 263.15, 262.25, 261.85, 262.05, 261.95, 261.85, 
    261.65, 261.45, 262.15, 261.85, 261.85, 262.75, 263.45, 263.95, 264.35, 
    264.65, 265.15, 265.75, 266.15, 266.55, 267.05, 267.35, 267.95, 268.25, 
    268.65, 268.75, 269.05, 269.35, 269.25, 269.95, 269.75, 270.15, 269.65, 
    269.55, 270.35, 270.35, 270.95, 271.15, 270.85, 270.75, 270.55, 270.65, 
    270.75, 271.05, 270.95, 271.15, 271.25, 271.05, 271.05, 271.05, 270.75, 
    270.75, 270.55, 270.45, 270.25, 269.95, 269.15, 268.55, 266.05, 265.95, 
    267.35, 267.45, 267.65, 272.05, 272.65, 272.55, 272.05, 272.45, 272.45, 
    272.35, 271.95, 272.25, 271.85, 272.25, 271.95, 271.65, 271.55, 271.35, 
    270.65, 270.55, 269.55, 269.45, 268.65, 268.15, 267.95, 267.75, 267.25, 
    266.85, 266.85, 266.85, 266.45, 266.25, 265.95, 264.95, 264.45, 263.75, 
    263.45, 263.75, 263.75, 263.55, 263.95, 263.05, 263.45, 263.85, 264.35, 
    263.75, 262.85, 262.15, 262.25, 261.85, 261.85, 261.55, 261.35, 261.65, 
    262.25, 262.65, 262.55, 262.45, 262.35, 262.65, 263.15, 263.65, 263.55, 
    263.45, 263.15, 262.85, 262.75, 262.85, 262.95, 262.65, 263.15, 263.25, 
    263.35, 263.25, 260.35, 259.75, 261.25, 260.15, 259.95, 260.75, 260.35, 
    260.65, 259.75, 260.95, 260.25, 259.95, 260.65, 260.15, 260.55, 260.75, 
    259.75, 260.35, 260.95, 260.95, 260.45, 265.55, 266.35, 266.65, 266.45, 
    266.25, 265.55, 265.65, 265.85, 266.15, 266.35, 266.55, 266.05, 265.75, 
    265.85, 265.55, 265.45, 265.45, 266.35, 266.05, 265.95, 265.95, 266.75, 
    267.65, 267.55, 267.85, 267.85, 268.95, 267.75, 268.05, 268.75, 267.65, 
    268.15, 267.45, 267.65, 267.25, 267.35, 267.35, 267.25, 267.55, 268.05, 
    268.75, 268.95, 269.15, 269.25, 269.45, 269.15, 269.35, 270.15, 270.15, 
    270.05, 270.15, 270.15, 269.75, 270.05, 270.05, 270.25, 270.25, 270.15, 
    270.05, 270.25, 269.95, 269.75, 269.45, 269.05, 269.45, 269.95, 269.55, 
    269.05, 269.25, 269.35, 269.35, 268.95, 268.75, 268.45, 268.15, 267.95, 
    267.65, 267.15, 266.95, 266.75, 266.55, 266.35, 266.05, 265.85, 265.45, 
    265.15, 264.85, 264.65, 264.65, 263.05, 262.35, 262.55, 262.25, 261.75, 
    260.75, 261.45, 260.45, 261.15, 260.45, 261.45, 260.85, 260.15, 260.35, 
    259.55, 259.65, 260.65, 260.85, 260.05, 259.55, 260.55, 260.95, 262.15, 
    262.55, 262.85, 263.25, 263.65, 264.15, 264.65, 265.05, 263.55, 261.95, 
    261.45, 261.05, 260.55, 261.65, 262.15, 261.55, 260.85, 261.05, 260.35, 
    261.05, 261.85, 262.45, 261.85, 263.45, 263.45, 264.85, 265.55, 265.55, 
    266.75, 267.05, 266.95, 267.05, 266.95, 268.15, 268.35, 268.45, 268.45, 
    268.35, 269.05, 268.85, 268.55, 268.35, 268.15, 267.85, 268.05, 268.35, 
    268.15, 268.05, 267.55, 268.05, 267.65, 268.05, 267.15, 267.05, 266.95, 
    267.05, 266.85, 266.65, 266.05, 266.95, 266.05, 266.15, 266.15, 266.15, 
    265.45, 265.15, 265.35, 265.45, 266.05, 267.55, 267.65, 267.45, 267.25, 
    266.95, 266.65, 267.05, 266.85, 266.05, 266.95, 266.35, 266.45, 264.85, 
    264.45, 264.25, 263.65, 263.35, 262.65, 263.05, 262.85, 262.25, 262.35, 
    261.85, 262.35, 261.65, 262.15, 262.25, 263.05, 264.25, 264.55, 264.55, 
    264.75, 265.35, 264.55, 264.95, 264.35, 263.75, 263.05, 262.55, 263.45, 
    264.25, 264.95, 265.05, 264.95, 264.85, 265.15, 265.35, 265.75, 265.85, 
    265.95, 266.35, 266.75, 266.75, 266.95, 267.05, 267.05, 266.75, 266.75, 
    266.85, 266.85, 267.05, 266.75, 266.45, 266.65, 266.65, 266.75, 266.85, 
    266.95, 266.95, 267.35, 267.05, 266.75, 266.45, 266.05, 265.55, 265.35, 
    264.55, 264.65, 264.35, 264.05, 263.95, 264.05, 263.55, 262.95, 264.05, 
    264.15, 264.65, 263.05, 260.75, 264.55, 262.35, 261.05, 262.65, 262.65, 
    262.15, 262.35, 264.95, 264.85, 264.95, 265.75, 266.45, 266.45, 266.45, 
    267.05, 266.45, 266.35, 266.45, 265.35, 264.65, 263.95, 263.55, 262.45, 
    263.25, 264.05, 263.25, 262.85, 262.35, 261.55, 263.35, 263.15, 261.65, 
    262.35, 260.75, 261.65, 260.85, 261.45, 261.35, 262.15, 261.25, 259.75, 
    261.95, 262.45, 262.35, 261.75, 261.45, 261.75, 259.55, 261.35, 260.95, 
    259.45, 260.05, 259.15, 261.25, 259.25, 258.65, 259.45, 260.35, 257.95, 
    258.75, 257.15, 258.85, 259.95, 259.45, 260.15, 259.75, 261.55, 261.25, 
    261.35, 261.95, 262.35, 262.05, 260.45, 260.15, 260.15, 263.35, 263.75, 
    264.65, 263.95, 264.65, 264.95, 265.15, 264.45, 265.25, 266.95, 267.35, 
    267.45, 267.35, 267.25, 266.85, 267.05, 266.45, 265.85, 265.15, 265.45, 
    265.95, 265.35, 265.45, 265.55, 265.45, 265.75, 264.95, 264.15, 264.45, 
    263.55, 262.75, 261.65, 261.15, 260.55, 259.75, 259.05, 258.05, 259.15, 
    257.15, 256.05, 257.05, 257.65, 257.65, 257.45, 255.65, 255.55, 256.05, 
    256.75, 255.85, 255.75, 256.25, 255.25, 255.75, 256.65, 255.65, 256.85, 
    258.05, 255.15, 255.05, 256.45, 256.05, 255.95, 257.65, 258.15, 257.25, 
    257.75, 255.65, 257.15, 255.15, 256.85, 256.55, 257.55, 257.75, 256.85, 
    256.95, 258.15, 257.65, 258.15, 258.55, 258.85, 257.95, 257.85, 259.25, 
    257.75, 259.65, 259.45, 258.85, 258.25, 257.65, 258.55, 258.05, 257.55, 
    256.55, 256.85, 256.65, 255.65, 255.65, 255.35, 256.75, 256.35, 255.65, 
    254.75, 254.55, 255.45, 254.35, 255.15, 255.45, 254.75, 256.75, 255.55, 
    255.95, 258.95, 253.75, 255.15, 256.35, 256.05, 257.35, 257.15, 256.65, 
    259.05, 257.65, 259.65, 257.45, 258.55, 256.85, 257.55, 255.95, 254.45, 
    255.65, 258.55, 256.65, 256.65, 259.05, 258.95, 258.85, 258.65, 258.75, 
    258.05, 256.55, 258.25, 254.65, 258.25, 258.65, 258.45, 257.35, 257.05, 
    255.45, 255.75, 255.75, 255.05, 255.75, 256.75, 257.45, 256.95, 256.65, 
    257.95, 258.35, 258.55, 258.55, 260.15, 258.75, 257.45, 258.15, 259.25, 
    257.65, 257.95, 258.85, 258.85, 259.35, 258.25, 258.75, 257.35, 256.05, 
    256.05, 255.95, 255.25, 254.55, 255.55, 254.85, 254.65, 256.35, 255.15, 
    255.85, 256.85, 254.45, 254.25, 254.05, 254.95, 255.45, 255.55, 254.85, 
    255.05, 255.15, 254.65, 254.05, 252.85, 254.65, 255.65, 256.35, 255.95, 
    256.65, 256.35, 256.55, 257.15, 257.75, 258.45, 257.35, 258.75, 258.15, 
    259.15, 258.95, 259.85, 259.75, 260.85, 261.05, 262.05, 261.45, 262.25, 
    262.85, 265.15, 264.95, 265.45, 265.85, 266.65, 266.75, 267.05, 267.35, 
    267.15, 267.75, 267.75, 267.55, 267.25, 266.85, 266.55, 265.75, 265.95, 
    266.35, 265.45, 265.75, 265.95, 266.65, 264.95, 264.75, 264.75, 264.85, 
    266.45, 264.85, 266.35, 264.75, 266.35, 265.95, 265.25, 266.05, 265.65, 
    267.95, 267.35, 267.95, 268.45, 269.45, 269.45, 268.45, 268.45, 268.65, 
    269.05, 269.25, 269.45, 270.35, 270.35, 271.05, 271.55, 271.85, 271.95, 
    272.55, 271.75, 272.15, 272.25, 272.85, 273.05, 272.45, 272.45, 272.55, 
    272.45, 272.55, 272.45, 272.75, 273.05, 272.95, 273.05, 272.95, 272.65, 
    271.15, 270.65, 270.35, 270.85, 271.15, 271.05, 270.75, 270.25, 270.25, 
    270.35, 269.75, 269.95, 270.25, 270.15, 270.05, 270.15, 269.95, 269.85, 
    269.65, 269.65, 269.55, 270.05, 269.95, 270.45, 269.15, 269.05, 269.05, 
    269.15, 269.85, 270.15, 269.25, 269.05, 269.45, 269.15, 270.35, 270.25, 
    269.75, 270.05, 270.05, 269.65, 269.05, 268.55, 270.55, 269.55, 270.05, 
    271.35, 274.25, 273.75, 272.95, 272.25, 271.35, 271.05, 271.05, 271.25, 
    271.35, 271.25, 271.55, 272.35, 272.55, 272.35, 273.95, 273.25, 273.65, 
    273.75, 273.25, 272.95, 272.65, 272.25, 271.95, 271.85, 271.15, 270.95, 
    271.25, 271.25, 271.25, 270.75, 270.35, 270.15, 269.55, 269.85, 269.85, 
    269.45, 268.55, 267.45, 268.25, 268.25, 267.75, 266.45, 266.05, 266.65, 
    266.75, 266.05, 266.45, 266.25, 266.75, 265.95, 266.25, 265.35, 265.05, 
    263.95, 263.95, 265.65, 264.85, 265.75, 265.85, 266.05, 263.95, 264.15, 
    264.65, 265.15, 265.75, 266.95, 266.25, 266.85, 266.15, 266.15, 265.45, 
    266.45, 265.65, 266.45, 265.95, 267.75, 267.45, 268.25, 268.65, 268.15, 
    267.25, 265.75, 265.25, 264.95, 265.25, 265.45, 266.05, 267.65, 266.25, 
    266.55, 266.85, 265.75, 267.45, 268.55, 267.55, 268.25, 269.65, 270.15, 
    269.65, 272.05, 272.95, 273.45, 273.25, 273.75, 273.75, 273.95, 273.95, 
    273.15, 273.65, 273.85, 273.85, 273.55, 273.15, 272.65, 272.45, 272.25, 
    272.85, 273.35, 272.25, 272.25, 272.25, 271.85, 271.45, 271.75, 270.35, 
    270.85, 270.15, 270.25, 270.45, 270.85, 270.95, 271.25, 270.95, 271.05, 
    270.75, 270.95, 270.85, 271.15, 270.75, 270.15, 269.55, 273.35, 272.25, 
    272.35, 272.65, 272.65, 272.85, 273.35, 272.95, 273.05, 273.15, 273.95, 
    274.05, 274.05, 274.15, 274.75, 274.35, 274.15, 273.75, 274.25, 274.35, 
    274.45, 274.35, 274.05, 274.15, 273.95, 273.85, 273.55, 273.75, 273.25, 
    273.15, 272.95, 273.05, 272.75, 272.95, 272.15, 271.05, 270.55, 271.35, 
    271.35, 270.75, 270.45, 270.15, 270.45, 270.25, 270.25, 270.15, 269.65, 
    269.75, 269.65, 268.65, 269.15, 269.55, 269.65, 269.15, 270.45, 270.65, 
    271.85, 271.25, 270.25, 269.95, 269.65, 269.45, 269.25, 269.55, 269.35, 
    269.75, 269.95, 269.85, 269.95, 270.15, 269.95, 270.15, 269.75, 268.55, 
    269.15, 267.95, 268.05, 268.45, 268.15, 265.95, 265.05, 264.85, 264.35, 
    263.55, 263.65, 263.75, 263.15, 263.55, 261.65, 261.45, 261.05, 261.95, 
    262.15, 260.25, 261.85, 262.15, 260.65, 261.05, 261.45, 260.85, 260.95, 
    261.05, 262.25, 262.15, 262.85, 262.55, 263.25, 263.35, 263.35, 263.45, 
    269.55, 269.85, 265.95, 267.25, 266.45, 265.05, 264.35, 264.25, 264.55, 
    264.65, 265.15, 264.95, 264.55, 264.25, 262.05, 261.85, 262.55, 263.65, 
    264.65, 264.75, 264.85, 264.55, 263.95, 263.45, 263.25, 263.45, 263.35, 
    262.35, 263.45, 262.95, 262.75, 262.15, 259.75, 258.85, 260.85, 261.25, 
    260.45, 260.55, 259.85, 260.95, 260.45, 260.35, 260.45, 260.35, 259.45, 
    259.15, 259.35, 258.35, 257.85, 257.85, 257.95, 258.45, 258.35, 257.85, 
    258.75, 258.35, 258.55, 258.15, 258.35, 257.75, 257.45, 259.15, 260.05, 
    259.35, 259.75, 259.65, 259.95, 259.25, 260.35, 259.95, 260.25, 260.15, 
    260.35, 260.15, 260.55, 260.25, 259.85, 258.85, 256.85, 254.85, 254.45, 
    254.35, 254.75, 255.55, 254.45, 254.85, 256.45, 255.85, 256.25, 255.35, 
    255.65, 256.35, 255.65, 255.55, 253.65, 255.85, 254.85, 255.05, 255.35, 
    255.65, 255.05, 254.85, 254.65, 254.65, 254.05, 254.75, 254.25, 254.35, 
    253.65, 253.65, 254.25, 253.65, 254.65, 253.15, 255.15, 254.35, 252.55, 
    253.95, 255.25, 253.35, 254.45, 254.75, 256.35, 257.15, 257.05, 258.35, 
    259.15, 259.05, 259.25, 259.65, 260.15, 259.95, 260.05, 263.25, 262.05, 
    262.05, 261.05, 260.45, 260.45, 260.35, 260.65, 260.35, 259.65, 259.25, 
    260.35, 260.85, 261.15, 261.45, 262.15, 262.25, 262.35, 262.35, 264.15, 
    267.15, 270.15, 270.55, 270.55, 270.45, 270.05, 270.75, 270.35, 269.65, 
    269.65, 269.65, 270.05, 270.25, 270.25, 269.95, 270.35, 269.55, 269.55, 
    268.75, 268.25, 267.95, 267.85, 268.55, 268.15, 265.85, 265.25, 265.85, 
    264.05, 264.05, 264.95, 264.75, 265.45, 265.85, 265.45, 265.55, 265.25, 
    265.55, 263.85, 263.35, 263.45, 262.85, 262.35, 262.65, 263.55, 263.85, 
    263.35, 263.05, 265.25, 264.05, 264.25, 267.35, 267.95, 266.65, 268.45, 
    267.55, 268.35, 269.15, 269.85, 270.15, 270.35, 269.95, 270.15, 270.45, 
    275.65, 275.95, 275.65, 275.35, 275.35, 275.55, 275.05, 274.65, 274.85, 
    275.25, 274.95, 275.75, 275.75, 275.65, 275.75, 275.95, 275.75, 276.05, 
    275.95, 275.55, 276.05, 274.95, 275.45, 276.55, 275.85, 276.35, 276.05, 
    275.65, 275.85, 276.05, 276.05, 275.35, 274.45, 274.35, 274.65, 274.25, 
    274.55, 274.45, 273.75, 273.15, 272.25, 271.55, 270.45, 271.25, 271.35, 
    270.45, 270.55, 268.95, 270.85, 267.85, 268.85, 270.25, 272.15, 271.05, 
    271.25, 271.55, 271.85, 271.75, 271.55, 272.65, 272.65, 272.15, 271.45, 
    272.25, 271.65, 271.55, 271.35, 271.25, 271.55, 271.65, 271.35, 270.65, 
    270.45, 270.25, 270.35, 270.05, 268.85, 268.75, 267.65, 267.75, 267.75, 
    267.85, 267.35, 268.55, 267.25, 268.35, 267.85, 267.55, 268.15, 267.75, 
    269.15, 268.55, 268.05, 267.35, 266.95, 266.65, 266.65, 267.05, 266.55, 
    267.25, 267.15, 267.25, 266.55, 265.65, 265.65, 265.35, 264.55, 264.15, 
    263.45, 264.05, 262.25, 262.25, 262.35, 262.45, 260.85, 260.85, 260.85, 
    260.55, 259.95, 259.45, 258.95, 258.45, 257.95, 257.55, 257.95, 258.75, 
    257.65, 257.45, 257.55, 257.45, 257.35, 257.05, 256.25, 256.65, 256.75, 
    256.65, 255.35, 255.55, 254.45, 254.45, 254.55, 254.45, 254.35, 255.15, 
    253.95, 254.45, 254.65, 253.95, 253.15, 252.25, 252.35, 252.65, 251.35, 
    251.15, 251.65, 251.75, 252.35, 252.05, 252.95, 251.55, 252.75, 252.65, 
    252.75, 254.05, 254.75, 254.25, 253.35, 253.95, 254.35, 254.65, 253.75, 
    254.95, 253.65, 253.15, 253.45, 253.75, 252.15, 253.55, 252.65, 252.95, 
    252.65, 252.05, 251.05, 251.85, 250.25, 249.95, 250.25, 248.75, 250.65, 
    250.05, 248.85, 249.05, 249.25, 249.05, 249.15, 247.15, 249.55, 250.25, 
    249.85, 248.45, 249.15, 248.35, 249.35, 247.75, 249.05, 249.35, 248.95, 
    248.85, 248.85, 249.05, 249.65, 249.35, 249.25, 249.15, 248.35, 249.45, 
    248.65, 248.55, 248.85, 248.75, 250.25, 249.25, 249.25, 249.45, 249.85, 
    250.15, 250.35, 250.85, 250.45, 250.75, 251.25, 251.75, 252.75, 251.65, 
    252.75, 254.25, 253.95, 254.95, 255.15, 255.35, 255.85, 255.95, 255.45, 
    255.65, 255.55, 255.35, 254.65, 254.85, 255.35, 253.15, 254.25, 254.65, 
    252.95, 253.35, 253.35, 251.25, 250.35, 253.25, 250.25, 252.55, 251.55, 
    250.55, 249.85, 249.35, 249.35, 249.25, 251.25, 251.95, 254.75, 254.25, 
    252.55, 253.75, 254.75, 254.55, 252.55, 252.65, 254.65, 253.95, 257.45, 
    254.45, 253.15, 254.05, 255.05, 254.75, 253.25, 254.05, 254.15, 254.25, 
    254.85, 254.75, 254.05, 254.45, 255.05, 255.75, 257.35, 259.05, 260.25, 
    260.85, 260.85, 260.65, 260.65, 260.95, 262.65, 268.45, 270.25, 270.55, 
    270.35, 270.65, 270.45, 270.55, 270.55, 270.35, 270.55, 270.55, 270.45, 
    270.55, 270.85, 270.75, 270.45, 270.15, 269.95, 270.05, 270.25, 271.05, 
    271.15, 271.35, 272.65, 272.15, 272.95, 273.45, 273.75, 273.75, 273.35, 
    273.85, 273.45, 273.75, 273.85, 273.95, 274.15, 274.35, 274.35, 272.85, 
    270.25, 270.65, 270.05, 269.75, 269.05, 267.75, 266.45, 265.15, 264.95, 
    263.25, 263.35, 262.45, 261.65, 259.65, 258.65, 258.55, 257.85, 257.35, 
    256.85, 255.55, 254.95, 254.45, 254.15, 253.95, 254.15, 254.15, 253.75, 
    253.85, 254.95, 254.85, 255.05, 255.05, 255.55, 255.35, 254.95, 255.15, 
    255.25, 255.75, 256.35, 256.45, 256.25, 256.05, 256.05, 256.15, 256.25, 
    256.25, 255.65, 255.25, 256.15, 256.55, 256.95, 257.35, 257.25, 256.95, 
    256.75, 256.65, 256.75, 256.85, 257.15, 257.25, 257.25, 257.35, 257.35, 
    257.15, 256.95, 256.55, 256.15, 256.15, 256.15, 252.65, 255.55, 254.35, 
    253.15, 252.05, 251.15, 252.95, 252.15, 252.05, 251.95, 251.85, 251.35, 
    252.65, 253.85, 252.35, 251.75, 251.05, 249.15, 249.85, 247.95, 247.35, 
    248.25, 247.35, 247.85, 249.65, 248.35, 248.05, 248.55, 247.45, 248.15, 
    248.95, 249.35, 247.85, 248.75, 247.85, 249.05, 249.35, 251.15, 249.65, 
    250.65, 249.35, 248.65, 248.75, 249.15, 248.65, 247.95, 248.95, 248.05, 
    246.95, 246.95, 247.95, 247.95, 247.35, 246.95, 246.35, 245.55, 247.25, 
    246.55, 247.55, 245.95, 246.65, 247.15, 246.45, 247.65, 246.55, 247.45, 
    247.25, 247.55, 246.15, 247.85, 247.95, 248.15, 250.35, 250.65, 251.35, 
    252.95, 253.15, 253.95, 253.85, 254.15, 254.35, 254.55, 254.25, 254.25, 
    254.75, 254.45, 254.95, 255.15, 255.25, 255.55, 255.25, 255.25, 255.25, 
    255.35, 255.65, 255.65, 255.35, 255.65, 255.85, 255.85, 255.65, 255.35, 
    255.15, 255.55, 255.35, 254.55, 254.25, 254.15, 253.85, 253.45, 251.45, 
    252.25, 250.75, 250.15, 251.55, 250.75, 251.75, 252.35, 251.45, 250.25, 
    250.85, 249.65, 249.75, 249.45, 250.25, 249.55, 249.95, 249.85, 250.95, 
    251.05, 251.25, 250.75, 250.25, 251.15, 251.05, 250.05, 250.55, 251.05, 
    251.35, 250.15, 250.85, 249.45, 248.95, 250.05, 248.85, 247.35, 250.35, 
    247.55, 248.95, 249.05, 250.95, 249.75, 250.15, 249.55, 250.05, 248.25, 
    248.25, 250.05, 249.55, 247.95, 250.65, 251.15, 252.95, 252.75, 253.05, 
    253.45, 255.25, 256.15, 254.55, 256.05, 260.85, 263.65, 263.25, 264.45, 
    264.35, 264.85, 264.55, 265.75, 266.25, 267.45, 269.55, 269.25, 268.95, 
    269.55, 269.85, 269.35, 269.45, 272.95, 273.65, 274.45, 274.85, 276.35, 
    275.05, 275.55, 276.25, 276.15, 275.55, 277.35, 277.65, 276.45, 275.05, 
    276.85, 276.95, 275.45, 276.35, 275.85, 274.65, 274.65, 273.75, 273.45, 
    273.35, 273.15, 272.95, 272.45, 272.65, 272.45, 271.95, 271.95, 271.55, 
    270.75, 271.45, 270.75, 270.45, 271.75, 270.65, 272.15, 269.45, 270.45, 
    270.05, 270.45, 269.15, 269.25, 269.55, 266.95, 267.15, 268.75, 268.55, 
    268.25, 267.85, 267.35, 266.55, 266.35, 265.75, 265.45, 264.55, 263.85, 
    263.05, 263.35, 262.85, 262.75, 262.15, 261.65, 261.45, 261.25, 261.35, 
    261.25, 261.05, 260.85, 260.55, 260.45, 260.25, 260.05, 259.95, 259.85, 
    259.75, 259.25, 259.15, 258.85, 257.85, 257.55, 256.95, 255.55, 254.35, 
    253.15, 252.75, 252.45, 252.15, 252.15, 251.75, 250.25, 251.55, 251.25, 
    251.75, 251.65, 251.75, 251.95, 254.25, 252.05, 252.65, 251.15, 252.45, 
    252.05, 250.65, 252.05, 251.55, 250.85, 249.75, 249.75, 249.95, 251.05, 
    248.35, 250.15, 249.55, 249.95, 249.95, 249.85, 250.25, 250.05, 250.35, 
    249.75, 249.15, 248.75, 248.65, 248.55, 248.15, 248.45, 247.85, 247.55, 
    247.55, 247.35, 248.35, 247.75, 246.75, 247.85, 247.85, 246.85, 246.25, 
    246.45, 246.65, 246.75, 247.15, 247.55, 247.35, 247.35, 247.75, 246.05, 
    247.55, 247.15, 247.25, 246.75, 246.65, 246.95, 247.35, 247.55, 247.45, 
    246.65, 246.45, 245.75, 245.75, 246.95, 246.85, 247.45, 247.45, 245.85, 
    245.85, 246.15, 247.75, 245.55, 246.45, 247.55, 246.15, 249.15, 246.25, 
    249.35, 249.75, 247.95, 249.45, 250.95, 251.15, 248.95, 248.55, 249.55, 
    249.55, 249.85, 249.95, 251.55, 252.75, 252.95, 254.75, 256.15, 255.85, 
    255.55, 255.25, 255.25, 254.55, 256.95, 255.55, 257.75, 260.05, 263.15, 
    264.25, 262.95, 263.75, 263.15, 261.95, 263.55, 263.65, 263.55, 263.45, 
    262.55, 263.15, 263.45, 263.45, 263.15, 264.15, 264.95, 264.45, 264.35, 
    267.35, 266.95, 267.85, 268.15, 268.15, 268.75, 269.15, 269.25, 269.75, 
    270.35, 269.65, 268.55, 268.35, 269.15, 268.45, 267.75, 268.05, 266.75, 
    266.55, 266.05, 265.65, 264.95, 266.05, 265.95, 265.05, 264.55, 264.15, 
    264.15, 262.85, 262.35, 261.05, 260.15, 259.35, 258.75, 257.45, 256.95, 
    256.75, 255.75, 254.65, 254.55, 255.75, 254.55, 254.15, 254.05, 254.45, 
    254.85, 253.35, 254.85, 254.65, 251.95, 252.05, 253.75, 253.05, 252.35, 
    251.15, 252.95, 251.85, 252.75, 254.15, 253.35, 254.95, 255.65, 254.45, 
    254.35, 255.55, 254.35, 252.85, 258.05, 254.75, 255.65, 253.75, 258.35, 
    257.15, 255.55, 255.55, 256.95, 257.65, 257.35, 256.55, 258.65, 257.05, 
    255.15, 255.55, 263.25, 263.45, 263.55, 262.95, 263.35, 263.65, 263.05, 
    262.75, 263.25, 263.85, 263.65, 263.85, 264.05, 264.05, 264.45, 264.55, 
    264.75, 264.55, 264.95, 264.95, 264.85, 265.05, 265.85, 266.15, 267.15, 
    266.45, 266.35, 266.65, 266.55, 267.05, 266.85, 268.05, 267.75, 267.85, 
    268.05, 268.45, 268.85, 268.95, 268.95, 268.95, 270.15, 267.85, 267.45, 
    267.75, 267.85, 267.25, 267.85, 267.55, 267.95, 268.75, 268.25, 268.85, 
    269.65, 269.95, 270.35, 271.15, 272.05, 272.45, 272.25, 271.45, 271.85, 
    272.95, 272.65, 273.65, 272.25, 272.65, 271.75, 270.85, 273.05, 272.75, 
    270.45, 271.95, 270.55, 270.75, 271.85, 270.55, 270.65, 270.35, 271.25, 
    270.45, 269.35, 268.45, 267.65, 267.85, 267.45, 267.05, 266.95, 266.85, 
    266.65, 266.55, 266.45, 266.35, 266.55, 267.05, 267.25, 263.35, 264.25, 
    265.35, 265.95, 265.95, 266.65, 267.05, 266.35, 266.25, 266.85, 267.45, 
    267.35, 267.05, 267.45, 267.75, 267.95, 268.25, 269.15, 269.35, 269.45, 
    269.85, 269.75, 269.55, 269.25, 269.15, 268.95, 268.75, 268.25, 268.05, 
    268.15, 268.25, 268.25, 267.85, 267.65, 268.25, 269.05, 269.55, 270.45, 
    270.75, 270.65, 270.75, 270.85, 271.05, 271.25, 271.25, 271.25, 271.25, 
    271.35, 271.35, 270.95, 270.25, 269.95, 270.15, 269.85, 269.35, 269.05, 
    268.75, 269.25, 269.35, 269.55, 269.75, 269.75, 269.95, 269.85, 269.45, 
    269.25, 270.25, 271.05, 271.55, 271.65, 271.75, 271.75, 271.45, 271.75, 
    271.75, 271.55, 271.65, 271.65, 271.85, 271.95, 271.85, 271.85, 271.75, 
    271.65, 271.75, 271.55, 271.15, 270.75, 271.05, 271.65, 272.15, 272.15, 
    272.05, 271.95, 271.85, 271.65, 270.15, 270.15, 269.15, 269.05, 269.05, 
    268.95, 268.55, 267.55, 266.95, 267.35, 267.75, 267.45, 265.65, 266.25, 
    266.75, 267.75, 268.55, 269.15, 269.25, 269.05, 268.95, 268.95, 268.85, 
    268.85, 268.65, 268.65, 268.55, 268.05, 267.75, 268.25, 268.75, 268.85, 
    268.75, 268.65, 268.65, 268.55, 267.05, 266.65, 266.85, 266.75, 266.85, 
    266.95, 266.65, 266.05, 265.85, 265.95, 265.75, 264.25, 263.95, 263.65, 
    263.55, 263.35, 263.15, 262.85, 262.65, 262.35, 262.25, 262.15, 262.15, 
    261.95, 261.95, 262.25, 262.45, 262.55, 262.65, 262.75, 262.75, 262.65, 
    262.45, 262.05, 261.45, 261.55, 261.05, 260.25, 259.35, 258.25, 257.25, 
    256.45, 256.05, 255.25, 254.95, 254.75, 254.35, 253.95, 254.95, 255.95, 
    257.65, 259.25, 261.35, 262.85, 263.75, 264.25, 264.45, 264.55, 264.85, 
    265.45, 265.75, 265.75, 265.45, 265.45, 265.75, 265.85, 265.65, 265.55, 
    264.45, 262.85, 261.65, 260.05, 259.35, 259.15, 260.65, 261.75, 262.65, 
    263.55, 264.05, 264.55, 264.75, 264.85, 264.65, 265.05, 264.75, 264.65, 
    264.75, 264.95, 264.65, 264.15, 263.55, 263.05, 262.85, 261.85, 261.25, 
    258.85, 257.95, 257.35, 257.45, 257.55, 258.35, 259.05, 259.35, 259.25, 
    259.45, 260.65, 265.85, 267.35, 267.45, 268.05, 268.55, 268.75, 269.15, 
    268.75, 268.55, 269.75, 276.45, 276.35, 276.25, 275.65, 275.65, 274.95, 
    274.95, 275.05, 275.15, 275.55, 275.55, 274.95, 274.55, 273.45, 273.65, 
    274.35, 271.85, 270.75, 270.65, 270.75, 271.35, 271.05, 270.85, 270.25, 
    268.35, 263.45, 261.85, 262.95, 260.75, 260.35, 260.35, 260.45, 260.65, 
    260.75, 260.85, 260.85, 260.75, 260.35, 259.95, 260.65, 260.25, 260.05, 
    259.65, 259.05, 258.45, 258.05, 257.85, 258.35, 258.45, 258.45, 258.45, 
    258.25, 258.05, 257.95, 258.05, 258.25, 258.35, 258.25, 258.15, 258.95, 
    257.55, 258.75, 259.05, 258.45, 256.75, 258.15, 257.25, 256.45, 258.25, 
    254.05, 258.95, 258.05, 256.95, 258.55, 257.45, 257.45, 258.55, 259.45, 
    259.45, 260.75, 261.05, 261.15, 261.05, 260.85, 261.75, 261.05, 261.15, 
    261.55, 261.45, 261.15, 261.15, 260.95, 260.85, 260.15, 260.25, 259.55, 
    259.05, 253.15, 252.95, 258.35, 258.35, 257.65, 257.35, 258.05, 257.95, 
    257.25, 257.25, 257.15, 257.05, 256.45, 257.05, 256.25, 256.95, 256.55, 
    256.35, 256.05, 256.35, 256.35, 253.15, 254.95, 255.95, 255.55, 254.85, 
    256.05, 255.75, 256.35, 255.05, 252.45, 254.35, 253.15, 252.85, 253.95, 
    254.35, 251.85, 251.95, 252.15, 252.05, 252.55, 250.15, 250.35, 249.25, 
    248.75, 252.75, 250.05, 251.95, 252.95, 250.55, 251.55, 252.15, 253.15, 
    253.45, 254.55, 254.55, 255.45, 251.95, 253.85, 252.75, 253.75, 252.45, 
    252.75, 252.25, 253.75, 246.25, 254.45, 245.65, 256.65, 250.65, 252.65, 
    253.85, 246.75, 246.35, 253.45, 254.55, 247.35, 247.85, 248.75, 257.65, 
    258.55, 257.95, 257.05, 257.55, 257.85, 261.05, 252.05, 260.75, 260.05, 
    252.55, 259.55, 258.45, 259.05, 250.95, 256.05, 255.85, 247.65, 255.75, 
    255.95, 245.85, 257.35, 246.75, 256.35, 254.55, 255.85, 256.55, 256.45, 
    253.95, 253.15, 254.55, 254.85, 249.65, 255.55, 254.55, 253.95, 249.15, 
    254.35, 255.65, 254.55, 256.75, 255.45, 254.95, 256.85, 257.15, 257.25, 
    258.15, 259.25, 259.25, 258.65, 256.15, 257.25, 256.45, 254.75, 255.35, 
    254.75, 253.65, 253.75, 253.55, 252.65, 253.95, 253.05, 250.85, 251.45, 
    252.75, 252.55, 253.55, 254.35, 254.95, 253.25, 254.15, 253.55, 254.05, 
    256.25, 255.25, 254.95, 255.75, 258.15, 258.25, 259.05, 262.95, 264.15, 
    260.35, 263.25, 263.95, 264.75, 265.25, 266.75, 267.65, 268.35, 267.55, 
    267.35, 268.65, 274.75, 275.15, 275.45, 275.35, 275.05, 275.15, 275.05, 
    275.25, 275.25, 275.35, 275.45, 272.95, 273.75, 272.65, 273.85, 274.15, 
    273.95, 273.65, 274.35, 273.85, 273.25, 274.15, 274.35, 274.15, 271.75, 
    274.25, 271.65, 273.25, 273.85, 273.35, 273.45, 272.15, 271.05, 271.55, 
    271.35, 271.05, 270.35, 270.65, 269.95, 269.85, 269.75, 268.35, 270.35, 
    270.95, 271.15, 271.45, 270.85, 270.35, 270.05, 270.05, 270.65, 270.75, 
    269.95, 268.65, 267.85, 264.95, 264.45, 263.55, 264.05, 263.85, 263.95, 
    259.65, 264.35, 263.05, 263.55, 264.05, 264.25, 264.25, 265.45, 259.15, 
    260.05, 261.45, 262.75, 263.75, 264.65, 265.25, 265.75, 265.65, 262.95, 
    262.85, 261.95, 261.85, 261.75, 261.95, 262.25, 262.65, 263.05, 263.35, 
    263.55, 263.95, 263.55, 264.05, 264.75, 265.15, 265.65, 269.35, 269.15, 
    268.25, 268.75, 267.45, 268.15, 267.65, 267.65, 268.05, 267.95, 268.05, 
    268.15, 264.15, 263.65, 263.25, 268.95, 268.35, 262.65, 263.05, 264.95, 
    269.85, 265.75, 269.45, 267.15, 270.15, 269.65, 270.05, 269.15, 269.25, 
    269.95, 269.55, 269.15, 269.35, 269.25, 269.55, 269.25, 269.65, 268.65, 
    263.75, 267.95, 267.85, 267.85, 267.45, 267.65, 266.45, 266.65, 266.95, 
    266.95, 266.75, 266.55, 266.85, 266.45, 265.25, 264.75, 264.25, 263.75, 
    263.85, 263.75, 263.65, 263.25, 260.35, 263.05, 263.15, 262.65, 262.15, 
    262.75, 262.05, 261.75, 262.05, 262.15, 261.85, 262.15, 262.05, 262.35, 
    261.65, 262.35, 261.55, 261.35, 260.55, 260.65, 261.15, 260.75, 260.55, 
    260.75, 258.55, 260.45, 260.25, 260.05, 260.05, 259.95, 258.05, 257.45, 
    260.65, 260.35, 260.25, 260.95, 261.65, 260.65, 260.15, 260.55, 259.55, 
    258.45, 256.85, 254.55, 254.85, 255.85, 255.65, 253.85, 254.95, 252.65, 
    250.55, 252.95, 253.75, 254.35, 255.35, 254.05, 255.15, 258.45, 256.65, 
    259.15, 259.35, 259.05, 259.95, 261.35, 260.85, 261.45, 261.45, 259.15, 
    259.35, 260.65, 260.25, 257.65, 262.45, 260.75, 256.45, 262.85, 261.75, 
    263.25, 262.45, 263.15, 264.65, 265.65, 271.65, 270.95, 271.05, 270.65, 
    269.95, 268.65, 268.25, 267.95, 267.45, 266.45, 266.15, 266.75, 265.95, 
    266.65, 263.05, 266.75, 267.45, 268.15, 268.75, 269.55, 268.85, 266.55, 
    270.65, 270.75, 270.65, 270.75, 270.35, 271.75, 271.35, 272.25, 271.15, 
    271.65, 271.05, 270.55, 271.45, 270.55, 270.95, 270.05, 268.65, 269.55, 
    266.05, 268.05, 266.65, 266.25, 265.45, 266.05, 265.15, 267.75, 268.55, 
    268.15, 269.75, 270.25, 269.75, 270.35, 269.95, 266.75, 267.65, 267.15, 
    263.95, 264.15, 265.85, 267.45, 264.65, 265.15, 267.15, 264.85, 264.95, 
    265.35, 265.85, 266.25, 267.05, 269.45, 269.65, 270.25, 270.25, 270.15, 
    270.55, 269.85, 268.85, 268.85, 268.35, 266.65, 266.15, 266.25, 266.35, 
    266.85, 259.05, 258.45, 266.15, 264.95, 267.15, 267.65, 268.55, 262.25, 
    269.35, 270.35, 270.65, 271.05, 270.95, 271.05, 270.05, 270.35, 269.65, 
    269.65, 268.85, 267.75, 268.35, 267.55, 265.45, 265.55, 265.65, 265.95, 
    266.45, 267.25, 267.95, 266.65, 268.45, 269.15, 269.55, 270.25, 270.65, 
    271.45, 272.05, 271.45, 272.65, 272.95, 272.55, 272.45, 272.55, 272.45, 
    272.55, 271.95, 270.55, 269.95, 270.25, 268.45, 267.65, 267.05, 267.95, 
    267.05, 268.45, 270.35, 271.05, 270.55, 272.05, 272.75, 270.95, 273.25, 
    270.65, 268.85, 267.75, 268.25, 267.45, 267.05, 267.25, 268.05, 267.15, 
    268.25, 267.95, 266.65, 268.15, 268.15, 270.35, 271.35, 271.35, 269.75, 
    270.05, 267.65, 267.65, 268.35, 269.75, 269.55, 269.25, 267.65, 267.75, 
    268.95, 269.75, 270.15, 270.45, 268.95, 269.75, 270.05, 270.75, 271.15, 
    271.05, 271.15, 272.15, 273.65, 274.05, 272.55, 272.35, 272.25, 272.45, 
    272.95, 273.35, 273.65, 272.95, 273.05, 274.05, 274.35, 272.45, 273.25, 
    273.15, 273.05, 273.25, 273.35, 273.25, 273.05, 273.25, 272.45, 272.55, 
    272.55, 271.45, 271.35, 271.05, 271.15, 271.25, 271.15, 271.95, 272.35, 
    270.05, 271.55, 271.45, 271.35, 274.05, 274.05, 276.85, 277.65, 275.75, 
    275.65, 275.55, 278.45, 277.85, 277.85, 276.85, 277.25, 277.25, 276.75, 
    276.25, 277.25, 276.65, 275.05, 274.75, 274.15, 274.85, 273.65, 274.15, 
    274.35, 273.75, 273.45, 271.75, 271.75, 272.15, 272.45, 271.95, 271.35, 
    271.15, 270.45, 269.65, 270.05, 269.15, 268.95, 268.45, 268.15, 267.45, 
    268.05, 268.35, 268.35, 268.25, 268.75, 270.05, 269.65, 270.15, 270.45, 
    270.25, 272.25, 270.95, 272.45, 272.35, 271.45, 270.25, 271.75, 268.45, 
    268.25, 270.65, 270.75, 270.75, 270.35, 271.55, 271.45, 269.85, 269.65, 
    268.65, 269.15, 270.75, 270.75, 271.15, 272.35, 269.45, 270.75, 269.95, 
    268.95, 267.95, 266.65, 266.35, 265.55, 265.05, 261.75, 261.95, 262.15, 
    260.65, 261.55, 263.05, 262.85, 265.05, 264.45, 263.55, 264.05, 265.95, 
    265.25, 267.55, 266.55, 267.25, 266.05, 267.65, 269.75, 266.95, 266.55, 
    265.75, 265.55, 262.25, 263.05, 262.45, 262.15, 263.05, 263.05, 263.65, 
    264.05, 264.15, 264.55, 263.95, 265.65, 264.45, 265.25, 264.75, 265.25, 
    265.55, 265.05, 265.35, 263.85, 263.95, 262.45, 262.95, 264.85, 265.15, 
    265.35, 266.25, 267.75, 266.85, 266.35, 266.75, 267.05, 266.35, 266.05, 
    265.75, 265.25, 264.65, 264.05, 263.25, 261.85, 261.45, 260.85, 260.75, 
    260.95, 260.85, 260.55, 260.85, 260.75, 261.45, 262.05, 262.45, 262.55, 
    262.95, 260.75, 260.45, 259.95, 259.55, 258.15, 257.45, 259.05, 258.85, 
    259.55, 262.05, 263.15, 262.95, 263.85, 264.95, 266.85, 270.35, 270.65, 
    269.45, 270.55, 270.35, 268.15, 266.15, 264.15, 266.35, 269.35, 269.15, 
    270.05, 269.65, 270.15, 269.75, 269.65, 269.25, 267.95, 267.65, 267.55, 
    268.15, 267.65, 267.15, 265.85, 266.15, 265.55, 267.45, 267.55, 267.75, 
    267.85, 267.75, 268.05, 269.15, 267.85, 267.75, 266.65, 265.85, 265.85, 
    265.75, 266.55, 265.55, 266.65, 266.75, 266.95, 266.15, 266.15, 266.85, 
    266.55, 266.35, 266.55, 266.35, 265.65, 265.85, 266.25, 265.95, 264.75, 
    266.05, 263.45, 265.85, 266.25, 266.45, 267.05, 266.75, 266.65, 266.65, 
    266.55, 266.55, 266.55, 265.65, 265.55, 265.05, 264.55, 262.95, 262.35, 
    264.35, 264.15, 265.15, 266.05, 265.45, 264.95, 266.45, 266.95, 265.65, 
    265.75, 264.45, 264.65, 263.55, 261.85, 263.45, 263.75, 263.85, 264.75, 
    265.85, 264.45, 264.95, 265.25, 265.15, 265.25, 264.55, 263.55, 261.85, 
    260.95, 261.45, 261.25, 262.85, 263.55, 265.95, 264.45, 265.35, 265.65, 
    267.05, 266.85, 265.05, 264.95, 265.25, 263.95, 263.75, 262.65, 260.85, 
    261.65, 264.45, 265.15, 266.65, 265.65, 266.05, 267.85, 266.65, 265.95, 
    265.25, 267.15, 266.55, 265.25, 263.65, 262.45, 262.45, 260.65, 258.85, 
    259.15, 260.85, 261.75, 260.25, 264.25, 265.85, 265.75, 266.75, 266.35, 
    267.95, 268.15, 266.55, 266.05, 266.75, 266.45, 265.05, 262.55, 267.05, 
    267.65, 268.15, 268.75, 268.35, 268.25, 268.85, 267.65, 267.65, 265.45, 
    265.95, 265.05, 265.35, 265.35, 265.55, 265.65, 265.35, 265.65, 265.45, 
    266.05, 266.45, 267.25, 266.75, 269.45, 269.35, 266.95, 267.75, 267.35, 
    267.55, 267.85, 269.25, 267.45, 267.15, 267.65, 267.55, 266.25, 264.75, 
    265.05, 265.85, 267.25, 267.15, 267.65, 269.05, 269.65, 271.05, 272.55, 
    270.75, 274.25, 270.75, 272.25, 273.65, 270.75, 271.15, 271.05, 271.55, 
    271.95, 272.15, 271.35, 271.55, 272.75, 270.65, 270.05, 270.45, 270.15, 
    269.95, 271.45, 271.65, 272.05, 272.65, 273.45, 274.05, 273.75, 272.85, 
    273.35, 273.35, 272.05, 273.05, 272.85, 271.35, 270.35, 269.75, 268.75, 
    270.65, 270.25, 269.75, 271.75, 272.25, 272.55, 272.75, 272.85, 273.25, 
    273.75, 272.85, 272.85, 272.65, 272.25, 272.95, 271.95, 271.75, 271.15, 
    270.45, 270.75, 269.55, 269.15, 267.65, 266.65, 266.15, 267.05, 267.25, 
    268.45, 270.45, 269.35, 270.35, 269.75, 269.75, 271.05, 273.05, 270.95, 
    271.95, 271.85, 270.35, 269.25, 270.05, 269.25, 268.65, 268.45, 267.85, 
    267.55, 267.95, 268.25, 267.65, 267.65, 267.75, 267.85, 267.65, 267.75, 
    268.15, 268.15, 269.05, 268.55, 270.05, 271.15, 268.65, 269.05, 268.25, 
    268.35, 268.85, 268.45, 268.15, 268.25, 268.35, 268.05, 268.55, 269.25, 
    269.25, 269.85, 269.95, 270.45, 269.85, 270.15, 271.95, 271.25, 271.75, 
    270.65, 270.25, 270.45, 269.85, 269.85, 269.55, 269.55, 269.35, 269.25, 
    269.05, 268.45, 268.15, 268.95, 268.85, 269.35, 269.15, 268.55, 270.55, 
    269.95, 268.65, 268.95, 268.45, 268.15, 268.35, 268.05, 267.55, 266.75, 
    266.15, 265.85, 265.55, 265.05, 265.05, 263.75, 263.55, 264.05, 265.05, 
    265.75, 266.85, 266.05, 266.15, 266.25, 266.85, 266.85, 267.65, 267.65, 
    267.45, 267.85, 267.45, 266.55, 266.45, 265.75, 265.65, 265.25, 265.25, 
    264.75, 264.75, 264.65, 264.65, 264.75, 265.25, 265.45, 266.15, 267.35, 
    268.55, 268.05, 268.55, 268.85, 269.45, 269.85, 268.05, 268.15, 268.45, 
    267.95, 268.15, 268.15, 268.25, 268.35, 268.45, 269.35, 269.85, 269.85, 
    269.95, 269.85, 271.15, 273.55, 270.55, 270.85, 272.95, 271.75, 270.95, 
    272.05, 271.35, 271.05, 271.35, 271.65, 271.55, 271.35, 272.45, 273.05, 
    272.55, 272.65, 272.65, 272.85, 272.95, 272.55, 273.55, 274.45, 274.05, 
    274.45, 274.45, 274.15, 275.55, 275.75, 276.65, 276.55, 275.65, 274.95, 
    275.15, 275.45, 275.35, 275.05, 274.45, 274.25, 273.55, 273.25, 273.25, 
    273.25, 272.85, 273.05, 273.75, 273.85, 273.55, 272.75, 272.45, 272.55, 
    272.85, 273.25, 272.45, 272.15, 271.85, 271.55, 271.25, 271.55, 271.55, 
    272.05, 271.95, 272.95, 272.55, 272.75, 273.05, 273.35, 273.65, 273.65, 
    273.95, 273.65, 273.75, 273.75, 273.35, 273.15, 273.65, 273.05, 272.35, 
    272.05, 272.25, 271.95, 272.35, 272.85, 273.15, 273.85, 274.25, 273.55, 
    273.85, 274.75, 275.75, 277.55, 277.05, 277.05, 277.15, 277.15, 274.15, 
    274.95, 273.85, 272.65, 271.95, 271.45, 271.15, 273.35, 272.35, 272.85, 
    272.35, 276.75, 275.25, 277.45, 275.65, 276.55, 275.25, 275.25, 278.45, 
    276.35, 276.45, 275.75, 275.15, 275.75, 275.15, 274.85, 274.95, 274.85, 
    274.75, 274.45, 274.75, 274.65, 274.75, 275.25, 276.15, 275.75, 276.55, 
    276.25, 276.95, 276.55, 276.25, 276.75, 276.15, 275.75, 275.35, 276.25, 
    276.55, 275.35, 274.95, 275.05, 275.05, 274.55, 274.05, 273.95, 273.85, 
    273.45, 272.95, 272.05, 271.65, 271.95, 271.25, 272.25, 271.45, 272.45, 
    271.95, 271.35, 271.25, 270.45, 270.55, 270.55, 270.45, 270.15, 270.15, 
    270.45, 270.25, 269.45, 269.95, 270.65, 270.45, 271.35, 270.75, 271.45, 
    271.75, 271.95, 271.45, 272.55, 272.85, 272.05, 270.15, 269.65, 269.15, 
    268.65, 270.25, 269.95, 273.55, 273.15, 274.25, 273.85, 274.05, 273.95, 
    273.95, 273.55, 271.55, 270.65, 269.25, 269.65, 270.75, 270.65, 272.45, 
    273.25, 274.85, 274.75, 274.55, 273.95, 274.05, 274.55, 274.05, 273.35, 
    273.35, 273.35, 272.95, 272.75, 272.85, 272.35, 272.85, 272.65, 272.85, 
    273.05, 273.55, 273.95, 274.75, 274.75, 274.05, 274.05, 274.25, 275.75, 
    274.95, 275.75, 274.05, 273.65, 272.35, 271.45, 270.65, 270.85, 272.05, 
    273.15, 272.35, 273.35, 274.95, 276.05, 274.25, 274.75, 274.85, 274.35, 
    275.15, 274.75, 274.55, 274.15, 274.85, 274.25, 273.65, 273.05, 272.45, 
    271.85, 271.35, 270.75, 270.15, 269.55, 270.65, 271.15, 271.85, 271.65, 
    272.55, 272.45, 273.15, 272.85, 273.55, 274.55, 276.05, 274.45, 275.35, 
    275.75, 276.25, 274.75, 274.55, 274.45, 274.55, 274.95, 275.25, 274.25, 
    274.25, 273.45, 273.65, 273.55, 274.55, 274.45, 273.35, 274.55, 274.45, 
    274.45, 274.75, 274.95, 274.65, 274.95, 274.95, 275.25, 274.95, 274.75, 
    274.55, 274.45, 274.35, 274.15, 274.55, 274.05, 274.25, 274.45, 274.65, 
    274.55, 275.35, 275.25, 275.15, 276.25, 275.25, 275.85, 276.55, 276.55, 
    277.25, 275.85, 275.95, 275.95, 275.55, 275.95, 275.45, 274.65, 273.85, 
    273.35, 273.05, 272.55, 273.35, 272.55, 274.25, 273.85, 274.55, 274.95, 
    275.35, 275.65, 275.95, 276.05, 276.05, 278.15, 277.55, 276.85, 276.55, 
    276.35, 276.05, 275.95, 275.65, 275.15, 274.45, 273.95, 273.35, 272.75, 
    272.25, 273.15, 274.35, 274.45, 274.35, 274.45, 274.65, 275.15, 275.85, 
    276.45, 275.85, 276.55, 275.55, 275.95, 276.35, 275.95, 276.15, 276.15, 
    276.15, 276.25, 276.25, 276.25, 276.05, 276.45, 276.95, 276.65, 276.45, 
    276.55, 275.95, 276.55, 275.85, 276.75, 276.95, 277.15, 277.55, 277.35, 
    276.65, 277.15, 277.15, 276.95, 276.55, 275.65, 275.25, 274.85, 274.65, 
    274.95, 274.85, 274.85, 274.95, 275.35, 274.75, 274.95, 275.25, 275.15, 
    276.35, 276.15, 275.55, 277.05, 276.45, 276.85, 276.35, 277.15, 276.65, 
    277.15, 276.45, 275.95, 275.55, 275.75, 275.45, 274.25, 274.55, 275.05, 
    274.95, 275.15, 275.15, 275.55, 275.55, 275.35, 275.55, 275.85, 275.85, 
    275.95, 275.55, 275.45, 275.55, 275.45, 276.75, 276.55, 275.85, 275.35, 
    275.55, 276.35, 276.75, 276.15, 276.35, 276.35, 276.15, 276.05, 275.95, 
    276.85, 276.35, 276.95, 276.95, 277.05, 276.75, 276.75, 277.75, 277.65, 
    277.05, 276.75, 276.35, 276.45, 276.45, 276.65, 276.45, 275.95, 275.95, 
    275.85, 275.55, 275.25, 275.75, 275.85, 275.75, 274.95, 276.15, 276.05, 
    275.95, 275.75, 275.75, 276.95, 277.05, 277.85, 277.25, 277.15, 277.05, 
    276.95, 277.25, 276.25, 275.85, 275.55, 275.35, 275.25, 275.45, 275.25, 
    275.25, 275.45, 275.35, 275.35, 275.45, 275.75, 276.15, 275.45, 276.35, 
    277.05, 276.65, 277.25, 275.85, 276.15, 276.65, 275.65, 276.15, 276.65, 
    276.55, 276.25, 275.75, 275.05, 274.95, 275.05, 274.25, 274.65, 275.05, 
    274.85, 275.25, 275.35, 275.35, 275.25, 275.75, 275.65, 276.25, 276.55, 
    276.45, 276.55, 276.75, 276.45, 276.15, 276.15, 276.15, 275.75, 275.85, 
    275.35, 275.55, 275.65, 275.95, 275.95, 275.45, 276.15, 277.25, 276.75, 
    277.25, 277.95, 277.75, 278.95, 277.45, 278.05, 278.55, 277.85, 277.75, 
    277.85, 277.35, 277.65, 277.95, 278.25, 278.45, 278.35, 277.65, 277.25, 
    277.45, 277.35, 277.25, 276.95, 277.05, 277.35, 277.75, 277.95, 278.85, 
    278.55, 278.95, 279.15, 278.55, 278.95, 278.75, 278.95, 278.55, 278.15, 
    278.45, 278.75, 278.85, 278.25, 278.05, 278.05, 277.75, 278.15, 278.55, 
    278.25, 278.05, 278.05, 279.25, 278.45, 279.05, 278.55, 277.75, 277.25, 
    276.35, 276.25, 276.25, 275.05, 274.15, 274.75, 274.85, 275.05, 275.75, 
    275.35, 275.25, 276.35, 276.15, 276.25, 276.95, 276.85, 276.65, 276.25, 
    276.85, 276.65, 276.45, 276.45, 276.85, 276.45, 276.55, 277.35, 277.05, 
    276.75, 275.15, 275.35, 275.35, 275.85, 276.65, 277.05, 276.65, 276.65, 
    276.65, 276.85, 276.75, 277.45, 278.05, 278.05, 278.25, 278.15, 278.05, 
    278.05, 278.05, 278.15, 278.05, 277.75, 277.25, 277.15, 277.55, 277.35, 
    277.65, 277.95, 277.55, 277.75, 277.55, 277.35, 276.85, 277.15, 277.45, 
    277.35, 277.55, 277.55, 277.85, 278.65, 277.55, 280.05, 278.45, 278.85, 
    279.15, 278.95, 279.35, 279.15, 278.85, 278.45, 278.45, 277.85, 277.85, 
    278.55, 278.25, 279.55, 279.15, 277.05, 278.35, 278.05, 277.55, 278.15, 
    277.55, 278.95, 279.85, 278.95, 281.15, 280.95, 280.95, 281.55, 280.05, 
    280.35, 279.95, 279.95, 279.25, 278.95, 278.75, 278.45, 277.95, 277.55, 
    277.35, 276.95, 276.95, 276.75, 277.85, 277.95, 278.55, 279.05, 279.05, 
    279.25, 279.25, 279.35, 279.45, 279.15, 277.65, 278.05, 277.15, 277.25, 
    277.05, 276.65, 277.35, 276.95, 276.75, 276.45, 276.55, 275.95, 276.25, 
    276.75, 277.05, 276.95, 276.65, 276.75, 276.95, 277.25, 277.25, 277.65, 
    277.45, 277.45, 277.95, 277.25, 276.95, 276.85, 277.35, 277.65, 277.65, 
    277.35, 277.15, 277.25, 277.15, 276.85, 277.15, 277.15, 277.35, 277.35, 
    277.15, 277.25, 277.95, 277.65, 278.25, 278.35, 278.45, 278.55, 278.55, 
    278.65, 278.65, 278.45, 278.25, 278.25, 278.35, 278.25, 277.95, 278.05, 
    278.05, 277.75, 277.85, 277.95, 278.05, 278.15, 278.35, 277.95, 277.55, 
    278.55, 278.35, 278.45, 279.15, 278.95, 278.65, 278.85, 278.75, 278.35, 
    279.15, 277.95, 277.95, 277.95, 277.65, 277.75, 278.25, 278.25, 277.55, 
    277.45, 277.35, 278.35, 279.35, 279.95, 280.65, 281.35, 280.65, 280.85, 
    280.35, 280.65, 280.45, 280.45, 280.55, 280.65, 280.45, 279.75, 278.85, 
    278.65, 279.05, 279.45, 278.75, 278.95, 279.35, 280.15, 280.15, 279.35, 
    279.15, 279.25, 279.55, 279.25, 279.25, 279.55, 280.25, 280.45, 280.15, 
    280.25, 280.25, 279.85, 279.55, 279.75, 279.85, 279.45, 279.25, 279.15, 
    278.85, 278.65, 278.85, 279.45, 280.05, 279.95, 280.35, 281.05, 281.25, 
    281.75, 281.95, 281.05, 281.35, 281.25, 281.55, 281.15, 281.45, 281.25, 
    281.65, 281.65, 280.95, 280.25, 280.05, 279.95, 279.95, 279.75, 279.75, 
    279.75, 279.95, 280.05, 280.05, 280.25, 279.45, 279.65, 279.55, 279.55, 
    279.85, 280.85, 280.15, 280.55, 280.75, 280.45, 280.45, 280.15, 279.75, 
    279.35, 278.95, 279.25, 279.05, 278.75, 278.85, 279.25, 279.15, 279.05, 
    278.85, 279.15, 279.15, 279.15, 279.85, 278.65, 279.75, 280.55, 280.25, 
    280.15, 279.45, 279.15, 279.05, 279.05, 278.85, 278.65, 278.45, 278.45, 
    278.25, 278.35, 278.35, 278.55, 278.75, 278.85, 279.05, 279.05, 279.55, 
    279.55, 279.65, 279.25, 279.95, 279.75, 279.75, 279.45, 279.65, 279.65, 
    279.55, 279.85, 279.65, 279.45, 279.05, 278.65, 278.35, 278.45, 278.45, 
    278.35, 278.45, 278.35, 278.55, 278.65, 278.45, 279.75, 279.85, 280.45, 
    280.25, 280.25, 279.65, 279.45, 279.35, 279.25, 278.95, 279.25, 279.05, 
    279.15, 278.95, 278.95, 278.95, 278.95, 278.95, 278.75, 278.65, 278.65, 
    278.55, 278.05, 278.35, 278.15, 278.35, 278.45, 278.45, 278.35, 278.15, 
    278.05, 278.15, 277.95, 277.75, 277.45, 277.85, 277.95, 277.95, 277.75, 
    277.45, 277.15, 277.35, 277.45, 277.45, 277.55, 277.15, 277.55, 277.55, 
    277.45, 277.15, 277.05, 277.15, 276.75, 276.65, 276.75, 276.75, 276.95, 
    277.05, 277.15, 276.55, 276.45, 276.25, 276.15, 275.75, 276.15, 276.25, 
    276.05, 275.95, 275.95, 276.25, 276.25, 276.75, 277.15, 277.15, 277.65, 
    277.45, 277.45, 277.85, 278.55, 278.15, 278.45, 278.65, 278.25, 278.05, 
    278.05, 277.75, 277.25, 277.15, 277.25, 277.55, 277.25, 277.15, 277.35, 
    277.95, 278.35, 278.65, 278.85, 279.35, 279.85, 280.55, 281.35, 282.15, 
    280.75, 280.45, 280.65, 280.85, 281.25, 281.05, 281.05, 280.45, 280.05, 
    279.65, 279.75, 279.55, 280.55, 280.25, 280.05, 278.85, 278.85, 279.05, 
    278.75, 278.85, 278.85, 279.15, 279.25, 279.55, 278.75, 278.85, 278.55, 
    278.45, 277.95, 278.05, 277.95, 278.25, 278.35, 278.35, 278.25, 278.05, 
    278.15, 278.15, 278.45, 278.65, 278.85, 278.85, 279.05, 278.95, 279.65, 
    279.65, 279.25, 279.25, 278.85, 279.15, 279.25, 278.95, 277.85, 277.35, 
    277.15, 277.25, 277.25, 277.55, 277.55, 277.55, 278.05, 277.75, 278.25, 
    278.35, 278.35, 278.35, 278.45, 278.25, 278.75, 279.35, 279.45, 279.55, 
    279.75, 280.05, 280.45, 279.75, 279.45, 279.75, 278.95, 278.55, 278.65, 
    278.55, 278.85, 279.25, 279.65, 279.95, 280.15, 280.45, 279.45, 279.75, 
    279.95, 280.15, 280.75, 281.15, 281.65, 281.05, 281.05, 280.85, 281.25, 
    281.25, 281.05, 280.25, 280.15, 280.05, 280.05, 279.75, 279.25, 279.55, 
    279.55, 279.15, 279.35, 279.45, 280.15, 280.05, 279.95, 280.25, 280.15, 
    280.65, 280.55, 280.85, 280.75, 281.35, 280.95, 281.05, 281.25, 280.55, 
    279.55, 279.35, 278.85, 278.55, 278.65, 278.65, 280.45, 279.95, 279.55, 
    280.15, 280.45, 281.15, 281.55, 282.05, 282.05, 282.75, 283.55, 283.35, 
    282.85, 282.55, 283.25, 282.25, 282.75, 281.85, 281.45, 280.95, 280.85, 
    279.75, 280.65, 280.25, 281.85, 281.05, 281.15, 281.95, 280.75, 281.95, 
    281.25, 281.25, 281.05, 281.05, 280.95, 280.65, 280.45, 280.65, 280.85, 
    280.55, 281.55, 280.45, 281.05, 281.25, 280.95, 281.65, 281.25, 281.15, 
    281.05, 280.65, 280.95, 281.25, 280.85, 281.65, 280.75, 279.95, 280.65, 
    280.75, 281.05, 280.55, 280.45, 280.65, 281.05, 281.35, 281.65, 281.95, 
    282.15, 281.95, 282.25, 282.55, 282.25, 282.25, 281.95, 281.75, 282.55, 
    283.95, 284.45, 285.45, 285.25, 285.75, 286.45, 286.45, 286.95, 286.45, 
    286.55, 285.65, 285.45, 285.35, 285.35, 285.25, 284.55, 284.55, 283.95, 
    283.15, 282.95, 282.95, 283.25, 283.65, 284.35, 284.55, 285.05, 285.15, 
    285.45, 284.75, 284.35, 284.55, 285.85, 285.95, 285.65, 287.15, 288.45, 
    287.25, 285.15, 285.65, 284.25, 283.35, 282.35, 281.65, 282.75, 283.35, 
    282.35, 281.05, 279.65, 279.65, 279.45, 279.55, 280.35, 280.85, 280.85, 
    281.15, 281.25, 281.25, 281.05, 280.75, 280.05, 279.35, 279.15, 278.85, 
    278.55, 278.25, 278.55, 278.15, 277.95, 277.85, 277.65, 277.55, 277.95, 
    278.15, 278.35, 278.35, 278.85, 279.35, 280.05, 281.05, 281.75, 281.15, 
    280.95, 280.65, 280.05, 279.65, 279.35, 279.05, 278.95, 278.65, 278.25, 
    278.25, 278.25, 278.25, 278.55, 278.15, 278.45, 278.15, 278.45, 279.15, 
    279.05, 279.65, 279.95, 280.25, 281.45, 281.75, 281.65, 281.65, 281.55, 
    281.75, 281.55, 281.25, 281.55, 281.75, 281.85, 281.95, 282.25, 282.15, 
    282.05, 282.15, 282.35, 283.45, 283.65, 284.75, 285.25, 285.85, 285.65, 
    285.45, 286.05, 286.65, 286.35, 285.95, 285.75, 285.85, 285.05, 283.75, 
    282.65, 282.15, 281.75, 281.35, 280.85, 280.55, 280.85, 281.15, 280.95, 
    281.45, 281.45, 281.75, 283.05, 283.65, 283.45, 282.45, 281.15, 284.65, 
    282.75, 281.55, 281.65, 280.45, 279.25, 279.55, 278.25, 277.35, 276.85, 
    277.05, 276.35, 275.95, 276.75, 277.25, 277.85, 277.85, 279.35, 279.95, 
    279.75, 279.35, 279.25, 279.15, 279.75, 280.45, 280.75, 280.95, 281.45, 
    281.25, 280.15, 279.85, 279.45, 280.45, 280.95, 281.05, 282.05, 281.75, 
    281.95, 281.75, 281.45, 281.25, 281.65, 281.45, 282.05, 282.15, 284.15, 
    283.15, 282.65, 282.35, 282.35, 282.15, 281.65, 281.05, 281.15, 281.15, 
    281.15, 281.15, 280.55, 279.75, 279.25, 279.55, 279.75, 280.55, 280.45, 
    281.15, 282.45, 283.15, 283.35, 282.65, 281.85, 281.15, 282.65, 281.75, 
    281.15, 280.85, 281.35, 280.85, 281.15, 281.75, 281.55, 281.25, 281.25, 
    280.85, 280.55, 279.85, 279.35, 278.85, 279.45, 279.85, 280.15, 279.45, 
    279.65, 279.95, 279.35, 279.85, 279.95, 280.75, 281.15, 280.25, 280.15, 
    280.25, 280.35, 280.25, 280.75, 279.55, 280.45, 279.25, 278.65, 279.05, 
    278.85, 279.95, 278.65, 280.95, 281.55, 283.35, 282.55, 283.15, 282.95, 
    283.65, 283.75, 283.75, 283.75, 283.15, 283.95, 283.65, 282.85, 281.75, 
    280.75, 281.05, 280.05, 279.95, 280.15, 280.75, 279.85, 280.25, 281.15, 
    281.15, 282.45, 284.35, 283.95, 284.25, 284.45, 284.65, 284.35, 283.75, 
    283.35, 283.15, 282.95, 282.95, 282.95, 282.55, 282.05, 282.05, 281.55, 
    281.25, 280.65, 280.85, 281.05, 281.25, 281.55, 281.65, 281.85, 281.95, 
    282.15, 281.55, 282.65, 282.45, 282.55, 282.25, 282.15, 282.05, 282.05, 
    282.95, 280.55, 280.55, 280.85, 280.35, 280.15, 280.75, 279.35, 279.15, 
    279.15, 279.45, 279.85, 280.45, 280.05, 279.05, 279.35, 278.95, 279.05, 
    278.95, 279.55, 280.15, 279.75, 279.65, 279.35, 279.35, 279.05, 278.45, 
    278.75, 278.85, 278.75, 278.45, 278.15, 278.35, 278.25, 278.25, 278.65, 
    278.15, 278.35, 278.75, 279.05, 279.15, 279.15, 279.65, 279.25, 279.15, 
    278.75, 278.95, 279.05, 278.95, 278.75, 278.85, 278.25, 277.95, 278.05, 
    277.95, 277.75, 277.45, 277.25, 277.85, 278.05, 278.35, 278.15, 278.55, 
    278.65, 278.75, 279.55, 279.35, 279.15, 280.75, 281.25, 279.65, 280.95, 
    280.55, 280.35, 280.05, 279.45, 279.85, 279.65, 279.35, 278.75, 279.05, 
    279.05, 279.25, 278.95, 279.15, 279.75, 279.95, 280.45, 279.45, 280.05, 
    279.45, 279.85, 280.25, 280.05, 280.45, 280.15, 279.75, 279.75, 278.85, 
    279.25, 279.25, 279.15, 278.75, 278.95, 278.95, 278.85, 279.35, 279.35, 
    278.95, 279.25, 279.35, 279.65, 279.95, 280.25, 280.45, 280.65, 281.45, 
    281.45, 281.35, 281.65, 281.55, 281.35, 281.65, 281.25, 281.75, 281.65, 
    281.05, 280.75, 280.55, 281.25, 280.75, 280.45, 280.05, 280.45, 280.45, 
    280.55, 280.85, 280.75, 280.55, 280.55, 279.65, 278.85, 279.65, 279.85, 
    279.65, 280.25, 280.55, 280.65, 281.25, 281.15, 281.75, 281.15, 281.45, 
    281.75, 282.55, 281.75, 282.35, 283.25, 283.95, 283.85, 283.75, 285.35, 
    284.45, 284.65, 285.15, 286.75, 283.85, 283.15, 283.15, 283.75, 283.95, 
    284.15, 282.85, 283.65, 283.25, 283.25, 283.75, 282.95, 282.75, 282.15, 
    283.95, 286.35, 286.25, 285.95, 286.85, 287.95, 286.75, 287.15, 288.15, 
    288.55, 288.35, 288.65, 288.55, 288.05, 287.25, 285.75, 284.85, 285.35, 
    284.35, 285.35, 284.55, 284.25, 285.55, 285.25, 286.25, 288.15, 288.65, 
    288.45, 288.45, 289.05, 289.85, 288.25, 288.65, 288.75, 288.65, 288.35, 
    286.65, 287.55, 286.15, 285.45, 285.75, 284.45, 284.75, 284.75, 285.25, 
    285.35, 286.65, 286.55, 287.45, 286.15, 286.15, 288.25, 288.25, 287.75, 
    286.85, 286.65, 286.75, 286.95, 287.45, 286.45, 286.35, 286.05, 285.15, 
    285.25, 284.55, 283.95, 284.05, 284.55, 283.95, 283.85, 284.05, 284.65, 
    283.65, 285.15, 286.35, 285.75, 286.35, 285.55, 286.05, 285.35, 286.35, 
    286.45, 286.05, 286.65, 285.85, 285.75, 285.05, 283.85, 283.95, 283.85, 
    282.95, 283.85, 282.25, 282.55, 282.95, 282.35, 284.15, 284.05, 283.75, 
    284.05, 284.55, 286.95, 285.15, 285.05, 285.35, 285.05, 284.45, 283.45, 
    281.95, 281.35, 281.75, 281.65, 281.35, 281.35, 281.05, 281.25, 280.75, 
    281.15, 280.85, 280.85, 281.15, 280.85, 280.85, 281.55, 281.05, 281.45, 
    282.05, 282.15, 282.25, 282.35, 281.75, 281.95, 282.15, 281.85, 281.75, 
    282.35, 282.95, 281.75, 281.25, 280.65, 281.25, 280.25, 281.15, 281.45, 
    281.35, 280.75, 282.35, 282.65, 282.25, 283.45, 283.85, 285.35, 284.25, 
    285.85, 285.65, 285.75, 284.75, 283.85, 283.05, 282.85, 282.85, 282.85, 
    282.45, 282.15, 281.55, 281.15, 281.45, 281.25, 281.05, 280.85, 281.25, 
    281.15, 281.35, 281.25, 281.45, 281.35, 281.05, 280.95, 280.85, 280.75, 
    280.65, 280.85, 281.05, 280.75, 280.75, 280.65, 280.35, 280.35, 280.15, 
    280.25, 280.25, 280.25, 280.85, 281.15, 280.95, 281.35, 280.95, 281.45, 
    282.05, 281.95, 281.65, 282.05, 281.25, 281.25, 281.35, 281.05, 280.95, 
    280.75, 280.65, 280.55, 280.45, 280.45, 280.45, 279.65, 279.65, 279.85, 
    280.15, 280.85, 280.95, 281.05, 281.35, 281.95, 282.25, 282.35, 281.85, 
    281.95, 281.95, 281.95, 281.85, 281.65, 281.45, 281.55, 281.25, 281.05, 
    280.75, 280.55, 280.35, 280.45, 280.45, 280.05, 280.15, 280.15, 280.15, 
    280.95, 280.95, 281.05, 280.95, 280.95, 281.25, 281.45, 281.55, 281.55, 
    280.85, 280.75, 280.85, 280.75, 280.65, 280.45, 280.15, 280.15, 280.15, 
    280.25, 280.25, 280.05, 280.45, 280.65, 280.95, 280.75, 281.15, 281.05, 
    281.15, 281.65, 281.55, 281.45, 281.55, 281.65, 281.35, 281.25, 281.25, 
    281.75, 281.35, 281.35, 280.85, 280.85, 280.95, 280.85, 281.45, 281.45, 
    282.25, 282.15, 281.75, 282.05, 282.55, 283.25, 283.45, 282.55, 283.55, 
    282.65, 282.45, 281.85, 282.05, 281.85, 281.55, 281.25, 281.05, 280.75, 
    280.75, 280.45, 280.75, 280.85, 280.75, 281.55, 280.85, 282.55, 282.95, 
    282.55, 283.25, 283.55, 283.45, 283.35, 283.75, 284.35, 285.05, 285.65, 
    285.85, 285.85, 285.55, 285.15, 284.45, 284.25, 284.25, 283.55, 283.45, 
    283.55, 283.35, 283.45, 283.55, 283.85, 284.55, 285.75, 285.65, 286.35, 
    286.65, 286.55, 286.35, 286.15, 285.95, 285.95, 285.15, 284.35, 283.05, 
    282.55, 282.15, 281.65, 280.65, 280.45, 280.35, 279.65, 281.05, 281.85, 
    282.85, 284.35, 284.55, 281.55, 281.45, 281.25, 281.25, 281.75, 281.55, 
    281.85, 281.45, 281.05, 280.85, 280.65, 280.25, 280.05, 280.25, 280.05, 
    279.95, 279.75, 279.75, 279.95, 279.95, 279.85, 280.15, 279.95, 280.55, 
    279.85, 279.85, 279.65, 279.75, 279.95, 279.85, 279.85, 279.95, 280.35, 
    279.95, 279.65, 279.65, 279.25, 279.45, 279.55, 279.35, 279.45, 279.35, 
    279.75, 279.75, 279.75, 280.05, 279.85, 280.45, 280.55, 280.55, 280.65, 
    281.45, 280.25, 281.65, 283.15, 281.45, 283.55, 283.65, 281.75, 280.95, 
    280.85, 280.75, 281.05, 280.55, 280.55, 280.55, 280.65, 280.65, 281.15, 
    280.85, 281.25, 280.55, 281.05, 280.85, 281.75, 281.45, 281.65, 281.15, 
    281.05, 281.15, 281.25, 280.95, 280.05, 280.05, 280.05, 280.65, 281.35, 
    281.15, 280.45, 280.25, 279.95, 279.55, 279.55, 280.75, 281.25, 281.15, 
    281.95, 282.15, 282.25, 282.25, 281.55, 281.25, 281.25, 280.95, 280.75, 
    280.45, 280.65, 280.25, 280.05, 280.25, 279.55, 279.35, 279.65, 279.85, 
    279.25, 280.35, 280.85, 280.35, 280.25, 280.55, 280.45, 280.25, 280.35, 
    280.25, 280.25, 280.35, 280.35, 280.05, 279.95, 279.65, 279.35, 279.15, 
    278.85, 278.85, 278.85, 278.85, 278.75, 278.65, 278.55, 279.05, 279.25, 
    278.95, 278.65, 279.15, 279.15, 279.45, 279.75, 279.95, 280.65, 280.45, 
    280.15, 280.15, 280.85, 280.95, 280.45, 279.45, 278.85, 278.95, 279.05, 
    278.95, 279.05, 278.85, 278.95, 278.85, 278.85, 278.65, 279.25, 279.95, 
    280.55, 280.65, 280.95, 280.95, 281.55, 280.95, 280.65, 280.55, 280.35, 
    280.55, 280.35, 280.05, 279.55, 279.35, 279.05, 278.75, 278.55, 278.65, 
    278.65, 278.65, 278.85, 279.25, 279.65, 279.95, 280.35, 281.55, 282.15, 
    281.95, 281.55, 281.15, 280.75, 280.25, 280.15, 280.15, 280.45, 280.25, 
    279.35, 279.55, 280.05, 280.15, 279.65, 280.05, 280.05, 280.25, 280.45, 
    280.45, 280.25, 280.15, 280.05, 279.95, 280.25, 280.65, 280.75, 280.25, 
    280.05, 279.95, 279.75, 279.65, 279.75, 279.55, 279.15, 278.55, 278.55, 
    278.65, 278.65, 278.65, 278.55, 278.45, 278.55, 278.55, 278.75, 278.65, 
    278.65, 278.85, 278.85, 279.05, 278.95, 279.05, 279.25, 279.35, 279.65, 
    279.65, 279.75, 279.65, 279.45, 279.35, 279.05, 278.55, 278.35, 278.05, 
    277.85, 277.85, 277.85, 278.05, 278.15, 278.25, 278.65, 278.95, 279.05, 
    279.35, 279.55, 279.25, 279.25, 279.15, 279.85, 278.85, 278.65, 278.55, 
    278.05, 276.95, 275.95, 275.85, 276.45, 275.25, 275.95, 275.75, 276.35, 
    277.55, 278.45, 278.95, 278.05, 278.15, 278.95, 279.25, 279.25, 279.45, 
    279.35, 279.45, 279.35, 278.95, 278.65, 278.25, 278.05, 277.75, 277.05, 
    277.75, 277.95, 277.65, 277.55, 277.65, 277.65, 277.65, 277.85, 277.95, 
    278.15, 278.35, 278.25, 278.35, 278.15, 277.95, 278.25, 278.25, 278.65, 
    277.95, 277.75, 277.55, 277.55, 276.25, 276.45, 275.95, 276.05, 275.15, 
    275.25, 274.95, 275.55, 276.05, 277.15, 276.95, 277.65, 277.75, 277.95, 
    277.95, 277.95, 277.65, 277.25, 277.25, 277.15, 277.15, 276.95, 276.75, 
    276.65, 276.35, 276.35, 276.05, 275.35, 275.45, 275.45, 275.75, 275.65, 
    273.75, 273.55, 273.45, 273.65, 273.65, 273.95, 274.65, 275.95, 276.75, 
    277.65, 278.65, 278.45, 278.85, 278.75, 278.45, 278.05, 278.75, 278.45, 
    278.45, 277.85, 277.65, 277.55, 278.05, 278.25, 277.85, 278.05, 278.35, 
    278.15, 277.85, 278.15, 278.15, 278.15, 278.15, 278.05, 278.15, 278.15, 
    277.65, 277.15, 276.95, 276.15, 276.65, 276.75, 277.35, 277.35, 277.15, 
    276.65, 276.55, 276.55, 276.75, 276.15, 276.55, 277.05, 276.55, 276.65, 
    276.55, 276.55, 276.75, 277.25, 277.35, 276.95, 276.35, 276.15, 275.95, 
    276.05, 275.65, 275.35, 275.65, 274.85, 274.75, 274.55, 274.45, 274.45, 
    274.85, 275.15, 275.15, 275.15, 275.85, 275.35, 275.35, 275.15, 275.25, 
    275.05, 274.95, 274.85, 274.75, 274.65, 274.35, 274.25, 274.15, 273.75, 
    273.75, 273.35, 272.75, 272.35, 272.75, 273.45, 274.35, 274.65, 275.05, 
    274.75, 274.55, 274.65, 274.45, 274.55, 274.35, 274.15, 274.15, 274.05, 
    274.05, 274.05, 274.25, 274.05, 274.05, 274.15, 273.35, 273.45, 274.45, 
    274.25, 273.95, 274.65, 274.65, 274.65, 274.95, 275.45, 275.85, 275.85, 
    276.05, 275.95, 276.05, 276.25, 276.35, 276.35, 276.35, 276.35, 276.25, 
    276.45, 276.35, 275.45, 275.45, 275.15, 275.15, 275.15, 274.95, 274.95, 
    275.05, 274.75, 275.45, 275.65, 276.25, 276.35, 276.35, 276.25, 276.25, 
    276.35, 275.85, 275.55, 275.75, 275.35, 274.95, 274.65, 274.65, 274.45, 
    274.25, 274.15, 273.65, 273.85, 273.65, 273.15, 273.35, 273.75, 274.15, 
    274.75, 274.95, 275.45, 275.65, 275.35, 275.15, 275.05, 275.05, 275.05, 
    274.75, 274.65, 274.45, 274.35, 274.25, 274.05, 273.95, 274.05, 274.25, 
    273.85, 273.95, 274.25, 274.55, 274.65, 275.05, 275.45, 275.35, 275.55, 
    275.75, 275.95, 276.35, 276.45, 276.45, 276.35, 275.95, 275.55, 275.45, 
    275.05, 274.05, 274.05, 273.85, 274.05, 273.65, 274.15, 273.75, 274.25, 
    274.45, 275.05, 276.05, 277.45, 277.15, 276.65, 277.05, 277.85, 278.45, 
    277.45, 277.75, 277.65, 277.55, 277.05, 276.75, 276.25, 276.15, 275.45, 
    274.95, 274.85, 275.15, 275.45, 275.45, 275.95, 276.05, 276.05, 276.35, 
    276.75, 276.75, 276.65, 276.75, 276.85, 276.75, 276.45, 276.75, 275.75, 
    274.75, 274.25, 273.65, 273.65, 273.25, 272.85, 273.35, 273.45, 273.15, 
    272.65, 273.05, 273.15, 272.95, 273.55, 273.85, 274.15, 274.35, 274.65, 
    274.95, 275.15, 275.15, 274.65, 274.55, 274.15, 273.45, 272.15, 271.55, 
    271.45, 272.35, 271.95, 272.35, 272.25, 272.65, 272.75, 273.15, 273.45, 
    273.75, 274.15, 274.45, 274.75, 274.75, 274.65, 274.65, 274.65, 274.75, 
    275.05, 275.45, 276.35, 276.45, 276.25, 276.25, 276.25, 275.55, 275.85, 
    275.65, 275.25, 273.65, 273.45, 273.35, 273.35, 273.45, 273.65, 273.75, 
    274.15, 274.25, 274.45, 274.85, 275.15, 276.55, 278.15, 278.45, 278.65, 
    278.15, 278.65, 278.55, 278.45, 278.85, 278.95, 278.75, 278.45, 277.95, 
    278.05, 277.25, 276.85, 276.55, 275.95, 276.35, 276.75, 277.05, 276.95, 
    276.45, 275.65, 275.45, 275.65, 275.85, 275.95, 275.85, 275.85, 275.85, 
    275.95, 276.65, 276.65, 277.45, 279.55, 279.25, 278.75, 278.55, 278.35, 
    278.35, 278.45, 278.55, 278.55, 278.55, 278.55, 278.65, 279.05, 278.55, 
    278.75, 278.55, 278.35, 277.95, 278.15, 277.95, 277.65, 277.15, 276.85, 
    276.95, 277.35, 277.65, 277.15, 277.45, 277.35, 277.55, 278.15, 278.15, 
    277.55, 277.55, 278.55, 279.55, 279.35, 279.25, 278.05, 278.15, 278.25, 
    278.75, 278.55, 278.25, 278.15, 278.35, 278.85, 278.95, 278.65, 278.35, 
    278.15, 277.45, 277.45, 277.15, 277.25, 277.45, 277.65, 277.25, 277.45, 
    277.25, 276.95, 275.85, 275.95, 276.05, 275.85, 275.85, 275.45, 275.55, 
    275.05, 275.15, 275.15, 274.35, 274.65, 273.35, 273.35, 273.15, 273.25, 
    273.65, 274.25, 274.05, 274.45, 274.55, 274.65, 274.85, 275.05, 275.25, 
    275.55, 275.45, 275.25, 275.55, 275.45, 275.35, 274.85, 275.05, 275.95, 
    275.65, 276.65, 276.55, 276.75, 276.35, 276.75, 276.05, 276.25, 276.35, 
    276.25, 276.55, 276.85, 277.05, 277.15, 277.15, 276.95, 276.45, 276.15, 
    275.65, 275.05, 275.15, 275.05, 274.75, 274.35, 274.05, 273.65, 273.45, 
    273.25, 273.05, 272.75, 272.65, 272.55, 272.35, 272.15, 272.25, 272.15, 
    271.95, 272.05, 272.05, 272.65, 273.35, 272.65, 272.85, 272.85, 272.65, 
    272.95, 273.35, 274.15, 273.85, 273.05, 272.85, 274.05, 273.15, 273.25, 
    273.65, 274.55, 274.85, 274.65, 274.85, 275.05, 274.95, 274.95, 274.95, 
    274.95, 275.15, 275.15, 274.75, 274.75, 274.05, 274.35, 274.15, 274.25, 
    274.25, 274.25, 274.05, 274.15, 273.75, 273.75, 273.85, 274.25, 274.25, 
    274.85, 274.85, 274.75, 274.85, 275.05, 274.45, 274.75, 274.35, 274.95, 
    275.25, 275.05, 275.05, 275.05, 274.65, 274.05, 274.45, 274.55, 274.75, 
    273.85, 274.85, 274.15, 274.55, 274.35, 274.55, 274.85, 274.75, 274.05, 
    273.95, 274.05, 274.05, 274.15, 274.45, 274.45, 274.45, 274.65, 274.55, 
    274.45, 274.35, 274.55, 274.65, 275.75, 275.45, 276.55, 276.05, 275.85, 
    275.65, 275.85, 276.15, 276.05, 277.25, 276.95, 276.85, 277.05, 277.25, 
    277.25, 277.25, 277.35, 277.25, 277.25, 277.55, 277.15, 277.35, 277.05, 
    276.75, 277.75, 277.25, 277.05, 277.05, 276.85, 276.95, 277.05, 277.65, 
    278.45, 277.75, 277.45, 277.45, 277.65, 277.95, 277.85, 277.65, 277.95, 
    277.85, 277.45, 277.25, 277.15, 276.95, 277.05, 276.95, 276.75, 276.35, 
    276.15, 276.05, 275.65, 275.45, 275.35, 275.25, 275.05, 275.25, 275.95, 
    276.15, 276.15, 275.85, 275.85, 275.85, 275.45, 274.95, 275.25, 275.15, 
    274.55, 274.85, 274.65, 274.65, 274.35, 274.75, 274.45, 274.65, 274.45, 
    274.25, 274.35, 274.65, 275.25, 275.85, 275.85, 276.15, 276.15, 276.15, 
    276.15, 276.35, 275.65, 275.85, 275.45, 274.55, 273.85, 274.05, 273.85, 
    274.25, 273.95, 274.25, 273.95, 274.55, 274.55, 274.25, 274.85, 274.75, 
    275.15, 275.45, 275.65, 275.55, 275.25, 274.95, 274.65, 274.35, 274.25, 
    273.65, 274.15, 273.85, 273.75, 273.25, 273.95, 273.75, 273.85, 273.85, 
    273.85, 273.75, 273.55, 273.65, 273.45, 273.45, 273.55, 273.75, 273.85, 
    273.75, 273.65, 273.65, 273.65, 273.85, 273.95, 273.95, 273.95, 273.95, 
    274.05, 274.25, 273.85, 273.95, 274.05, 274.55, 274.75, 274.95, 275.45, 
    275.95, 275.25, 275.25, 275.65, 275.45, 275.45, 275.95, 276.75, 276.45, 
    276.45, 276.95, 276.55, 275.95, 276.25, 276.45, 276.15, 275.65, 275.05, 
    274.95, 275.25, 275.25, 274.75, 274.85, 277.85, 276.25, 277.65, 276.05, 
    276.55, 276.35, 276.15, 276.65, 278.95, 278.75, 277.95, 278.65, 278.45, 
    277.45, 277.85, 277.95, 277.95, 277.65, 277.65, 277.95, 277.35, 277.75, 
    277.75, 276.55, 276.35, 276.75, 276.65, 276.55, 276.45, 276.35, 276.05, 
    275.35, 274.05, 272.55, 272.15, 271.55, 271.15, 270.95, 270.85, 270.85, 
    270.65, 270.65, 270.35, 270.65, 270.75, 271.05, 270.55, 270.35, 270.05, 
    269.75, 269.55, 269.65, 269.95, 269.65, 269.55, 269.45, 269.65, 269.85, 
    270.05, 270.05, 270.05, 270.15, 270.15, 269.85, 269.35, 269.75, 270.25, 
    269.85, 270.45, 269.65, 270.05, 270.05, 269.55, 269.55, 269.55, 270.15, 
    269.95, 270.15, 270.35, 269.55, 270.05, 269.95, 269.45, 268.65, 268.85, 
    268.55, 268.05, 268.25, 268.55, 268.65, 268.75, 268.65, 268.45, 268.55, 
    268.85, 268.45, 269.05, 268.95, 269.15, 269.35, 269.65, 269.85, 270.25, 
    270.35, 270.75, 270.75, 270.55, 270.45, 270.35, 269.95, 269.95, 269.35, 
    269.15, 269.45, 269.75, 270.05, 269.65, 269.75, 269.85, 269.85, 270.55, 
    270.55, 271.05, 270.45, 270.85, 271.85, 271.05, 270.95, 269.55, 269.35, 
    269.15, 268.65, 268.25, 267.75, 267.55, 267.55, 267.55, 266.85, 267.25, 
    267.35, 267.55, 267.25, 266.85, 267.25, 266.85, 267.15, 266.85, 267.95, 
    268.25, 268.75, 269.25, 268.25, 269.25, 268.65, 268.15, 267.35, 267.35, 
    266.65, 267.65, 266.95, 267.45, 266.75, 267.75, 268.25, 269.05, 269.55, 
    269.55, 269.85, 270.35, 270.75, 271.05, 271.45, 271.85, 272.25, 272.55, 
    272.25, 272.15, 272.05, 272.05, 271.85, 272.05, 272.45, 272.85, 272.65, 
    272.95, 272.65, 273.35, 273.65, 274.25, 274.05, 274.05, 273.55, 273.85, 
    273.75, 273.85, 274.35, 274.45, 274.85, 274.65, 274.85, 275.05, 275.05, 
    274.85, 274.35, 274.65, 274.35, 274.65, 275.15, 275.05, 274.45, 273.95, 
    273.75, 273.85, 274.35, 274.25, 274.05, 274.35, 273.65, 273.85, 273.75, 
    274.35, 274.25, 274.05, 274.45, 274.05, 273.35, 273.75, 272.25, 272.45, 
    271.65, 271.85, 271.25, 270.65, 271.75, 271.05, 270.45, 270.75, 270.55, 
    269.85, 270.25, 271.05, 271.05, 270.65, 270.85, 271.15, 271.45, 271.45, 
    270.65, 270.45, 269.45, 270.95, 269.25, 269.75, 271.25, 271.95, 272.15, 
    272.95, 273.55, 273.95, 272.95, 273.05, 274.55, 275.65, 275.25, 275.55, 
    275.15, 275.65, 275.85, 276.35, 276.45, 275.75, 275.15, 275.65, 275.25, 
    274.95, 275.85, 275.65, 276.25, 277.25, 277.05, 275.85, 275.75, 275.45, 
    276.05, 276.85, 277.35, 275.65, 275.85, 275.75, 275.05, 275.45, 274.65, 
    274.35, 274.65, 275.05, 275.75, 275.05, 275.35, 275.85, 275.05, 275.55, 
    275.55, 275.55, 274.95, 273.45, 273.15, 273.55, 272.95, 273.75, 272.85, 
    272.95, 272.95, 273.75, 272.75, 272.55, 272.65, 272.75, 272.85, 272.95, 
    273.05, 272.95, 272.45, 272.25, 272.15, 272.65, 272.55, 272.75, 272.75, 
    272.65, 272.65, 272.85, 272.35, 272.55, 271.85, 272.15, 272.35, 271.95, 
    271.95, 272.65, 271.95, 272.05, 272.15, 272.15, 271.85, 272.25, 272.05, 
    272.55, 272.35, 272.45, 271.65, 270.35, 269.85, 271.95, 270.55, 270.15, 
    270.25, 271.45, 270.65, 270.75, 270.05, 269.45, 269.15, 268.55, 269.05, 
    270.35, 272.55, 273.15, 273.45, 273.75, 273.85, 273.75, 272.55, 272.15, 
    272.35, 272.65, 273.55, 273.45, 272.85, 272.65, 273.95, 273.45, 273.35, 
    272.45, 270.65, 271.95, 271.85, 270.35, 270.55, 270.85, 271.25, 271.75, 
    271.55, 271.85, 271.75, 271.65, 271.65, 272.05, 272.45, 272.75, 272.95, 
    272.95, 273.05, 273.85, 275.05, 274.85, 274.35, 274.35, 274.25, 273.55, 
    273.35, 273.55, 273.45, 273.05, 273.45, 273.45, 273.65, 274.05, 273.65, 
    273.45, 273.25, 273.35, 273.65, 273.05, 273.05, 273.25, 273.15, 273.15, 
    273.45, 272.65, 273.25, 272.45, 271.15, 270.35, 270.25, 272.15, 272.25, 
    272.35, 271.65, 271.35, 270.55, 269.65, 267.75, 269.85, 269.85, 270.55, 
    270.65, 270.05, 270.05, 270.15, 269.75, 270.35, 270.75, 270.55, 270.25, 
    271.55, 270.35, 270.25, 270.65, 270.85, 271.05, 271.35, 271.55, 271.65, 
    271.55, 271.55, 271.45, 271.75, 271.85, 272.55, 272.75, 273.05, 272.45, 
    272.55, 272.55, 272.65, 273.55, 273.25, 273.25, 273.75, 273.45, 273.95, 
    275.35, 275.95, 275.45, 275.45, 276.05, 276.55, 276.45, 276.05, 276.15, 
    276.05, 275.15, 275.15, 275.05, 273.75, 272.55, 271.15, 270.65, 270.65, 
    270.25, 269.65, 268.75, 268.45, 268.05, 267.75, 267.45, 267.45, 267.45, 
    267.45, 267.15, 267.25, 267.35, 267.25, 266.95, 266.95, 266.85, 267.05, 
    267.05, 267.25, 267.45, 267.55, 267.65, 267.75, 267.75, 267.85, 267.85, 
    267.85, 267.75, 267.75, 267.95, 267.75, 268.05, 268.05, 268.05, 268.45, 
    269.15, 269.35, 269.45, 269.65, 269.85, 269.85, 270.05, 270.35, 270.55, 
    270.75, 270.95, 271.05, 271.45, 271.45, 271.55, 271.65, 271.65, 271.85, 
    272.15, 272.35, 272.35, 272.25, 271.75, 271.55, 271.65, 271.75, 271.45, 
    271.65, 271.35, 271.65, 271.25, 271.65, 271.55, 271.55, 271.35, 271.55, 
    271.65, 271.65, 271.35, 271.65, 271.45, 271.35, 271.65, 271.85, 272.05, 
    272.25, 272.45, 272.55, 272.55, 272.75, 272.55, 272.85, 273.35, 273.45, 
    273.45, 273.45, 273.15, 272.25, 273.35, 273.75, 273.95, 274.25, 274.75, 
    275.05, 274.15, 274.15, 274.55, 272.55, 270.55, 269.05, 268.45, 268.65, 
    269.95, 270.25, 271.85, 274.05, 274.15, 274.25, 274.05, 274.55, 274.05, 
    274.85, 274.45, 274.25, 274.65, 274.75, 274.65, 274.55, 274.75, 274.65, 
    274.75, 274.85, 274.55, 274.75, 274.45, 275.05, 274.65, 273.75, 273.55, 
    272.55, 272.25, 271.55, 271.05, 270.85, 270.85, 270.75, 270.15, 269.85, 
    269.75, 268.95, 269.15, 269.15, 269.25, 269.55, 269.45, 269.55, 269.35, 
    269.15, 269.05, 269.15, 268.75, 268.55, 268.25, 268.15, 267.85, 267.25, 
    265.95, 266.85, 265.55, 265.05, 265.85, 262.25, 264.25, 264.05, 262.65, 
    262.85, 263.55, 263.45, 263.95, 264.15, 263.95, 262.95, 261.85, 262.35, 
    261.55, 261.85, 261.15, 260.85, 260.15, 260.65, 260.65, 260.65, 260.05, 
    260.05, 259.55, 259.15, 260.45, 259.35, 259.85, 258.85, 260.15, 258.65, 
    259.45, 259.85, 261.25, 260.75, 261.65, 260.95, 261.05, 261.25, 261.55, 
    261.25, 260.35, 260.45, 260.35, 260.55, 261.05, 261.65, 262.25, 261.95, 
    262.55, 262.45, 262.65, 262.55, 262.65, 262.75, 263.55, 263.45, 263.45, 
    263.75, 264.45, 265.05, 264.95, 264.95, 265.25, 265.25, 265.35, 265.45, 
    266.25, 266.45, 266.55, 266.95, 267.65, 268.15, 268.55, 268.75, 269.15, 
    269.75, 269.65, 270.05, 270.25, 270.45, 272.05, 273.75, 275.35, 276.35, 
    276.45, 276.45, 276.55, 276.45, 276.05, 275.75, 276.05, 275.65, 276.25, 
    275.95, 276.25, 276.25, 276.35, 276.05, 275.55, 276.05, 276.55, 276.45, 
    276.15, 276.15, 275.75, 275.25, 275.25, 275.55, 275.45, 275.85, 275.55, 
    275.35, 275.25, 274.45, 273.85, 274.05, 273.85, 273.05, 272.95, 272.15, 
    272.75, 272.75, 272.55, 273.35, 273.75, 273.35, 273.45, 275.05, 275.85, 
    275.35, 275.35, 275.65, 275.55, 274.55, 275.05, 275.15, 275.45, 275.55, 
    275.35, 275.95, 275.05, 275.05, 274.35, 274.65, 274.45, 275.15, 273.85, 
    274.55, 273.85, 274.25, 273.85, 274.65, 274.35, 274.45, 273.85, 273.95, 
    274.35, 274.35, 274.25, 274.75, 274.75, 274.05, 273.85, 272.85, 272.75, 
    272.35, 271.65, 271.45, 270.75, 270.75, 270.55, 270.05, 269.85, 269.65, 
    269.45, 269.55, 269.35, 269.15, 269.05, 268.65, 268.55, 268.65, 268.45, 
    268.45, 268.35, 267.85, 267.65, 267.75, 267.75, 267.35, 267.35, 266.75, 
    266.85, 267.05, 266.75, 266.95, 267.05, 266.45, 265.85, 265.75, 265.65, 
    265.45, 265.35, 265.45, 265.75, 265.55, 265.25, 264.75, 266.15, 265.85, 
    265.65, 265.55, 265.25, 265.05, 264.85, 264.65, 264.25, 263.85, 263.55, 
    263.15, 262.85, 262.55, 262.15, 261.95, 261.65, 261.15, 260.55, 259.95, 
    259.25, 258.95, 258.65, 258.75, 258.45, 258.45, 257.95, 258.55, 259.05, 
    258.35, 258.25, 259.35, 258.15, 258.35, 258.85, 257.65, 258.25, 258.45, 
    258.75, 259.45, 258.75, 260.05, 260.35, 260.95, 259.95, 261.35, 260.55, 
    259.65, 260.35, 261.05, 260.15, 260.55, 260.65, 259.95, 260.95, 262.25, 
    261.25, 263.15, 263.55, 263.65, 264.15, 264.75, 265.25, 265.35, 266.05, 
    265.95, 266.05, 266.15, 266.85, 267.15, 267.95, 268.05, 268.95, 268.35, 
    268.35, 268.75, 268.25, 268.85, 268.85, 268.95, 268.95, 269.05, 268.85, 
    269.35, 269.85, 269.25, 269.75, 271.45, 271.55, 272.25, 272.25, 272.45, 
    273.95, 274.95, 275.75, 274.85, 274.75, 275.25, 275.35, 274.65, 274.45, 
    274.65, 274.25, 274.95, 274.35, 273.55, 276.85, 273.25, 273.35, 275.75, 
    275.35, 276.35, 276.05, 276.25, 277.45, 276.35, 275.85, 276.05, 275.25, 
    275.25, 275.55, 275.45, 274.95, 275.55, 272.75, 272.65, 273.15, 274.35, 
    275.35, 275.95, 277.15, 276.95, 276.95, 276.45, 276.35, 276.35, 276.45, 
    276.15, 276.35, 275.95, 276.25, 276.25, 276.45, 276.45, 277.15, 277.15, 
    276.75, 277.05, 276.85, 277.35, 277.25, 276.85, 276.65, 276.75, 276.65, 
    277.15, 277.55, 277.15, 276.85, 276.85, 276.75, 276.95, 276.95, 276.85, 
    277.55, 276.65, 276.25, 276.15, 275.95, 275.85, 275.45, 275.35, 275.15, 
    275.55, 275.25, 274.85, 273.55, 273.65, 274.85, 274.95, 275.15, 275.05, 
    275.35, 275.25, 275.45, 275.65, 275.65, 275.65, 275.35, 274.85, 274.95, 
    274.65, 274.85, 274.65, 274.45, 273.95, 274.15, 273.95, 274.25, 274.05, 
    273.65, 273.65, 273.85, 273.65, 273.65, 272.85, 272.75, 272.95, 272.55, 
    272.55, 272.25, 272.15, 272.65, 272.35, 272.35, 272.45, 272.95, 272.25, 
    272.45, 272.85, 272.65, 272.25, 272.15, 272.05, 271.95, 271.65, 271.95, 
    271.85, 271.75, 271.65, 272.15, 271.75, 271.25, 271.65, 271.65, 271.55, 
    271.15, 271.35, 271.15, 271.25, 271.25, 271.45, 271.45, 271.45, 270.95, 
    271.65, 271.95, 272.15, 272.35, 272.95, 272.95, 272.75, 272.95, 273.55, 
    273.65, 273.95, 274.35, 274.75, 275.15, 275.65, 275.65, 276.05, 275.95, 
    275.75, 275.15, 275.95, 275.85, 275.95, 275.65, 275.65, 275.65, 275.15, 
    275.65, 275.15, 275.35, 275.05, 275.35, 274.85, 273.75, 272.95, 274.05, 
    274.35, 274.55, 274.45, 274.25, 273.85, 271.75, 270.15, 270.65, 270.95, 
    268.95, 269.15, 268.65, 268.55, 267.15, 267.75, 266.45, 267.35, 266.95, 
    266.85, 266.85, 267.05, 267.95, 267.15, 267.15, 266.45, 266.75, 267.25, 
    267.85, 268.05, 268.65, 269.05, 268.75, 269.25, 269.25, 269.85, 269.85, 
    269.15, 268.75, 268.45, 267.85, 267.15, 267.35, 266.35, 266.25, 265.55, 
    265.15, 265.25, 265.15, 264.85, 263.95, 263.95, 264.05, 263.65, 263.55, 
    263.15, 262.95, 262.55, 262.65, 262.95, 262.95, 262.75, 262.95, 262.85, 
    262.65, 262.65, 262.75, 262.45, 262.35, 262.15, 262.05, 262.25, 262.05, 
    261.65, 261.65, 261.25, 260.45, 260.35, 260.55, 260.55, 260.25, 260.25, 
    260.25, 260.25, 260.05, 260.15, 260.45, 260.15, 260.75, 261.15, 261.15, 
    261.15, 261.25, 261.35, 260.75, 261.25, 262.05, 261.35, 260.95, 261.15, 
    261.25, 261.45, 261.65, 261.75, 262.25, 261.85, 263.05, 263.55, 264.05, 
    264.25, 264.35, 264.05, 263.85, 263.75, 263.95, 263.45, 263.15, 262.65, 
    262.75, 262.95, 263.05, 262.95, 262.35, 261.85, 261.75, 260.95, 260.95, 
    260.45, 260.35, 260.05, 261.05, 260.85, 261.65, 262.25, 262.95, 262.35, 
    262.95, 262.55, 263.15, 263.05, 263.15, 263.75, 264.35, 264.95, 264.95, 
    265.65, 265.85, 267.35, 267.65, 267.95, 265.95, 265.65, 263.95, 263.65, 
    263.55, 263.25, 262.35, 261.95, 262.15, 262.05, 263.15, 262.55, 262.65, 
    262.55, 262.35, 262.15, 262.25, 261.45, 262.15, 261.25, 261.35, 260.25, 
    263.25, 262.45, 263.25, 263.75, 263.05, 262.05, 261.45, 263.05, 261.95, 
    263.55, 262.85, 262.85, 264.45, 265.95, 265.35, 265.35, 264.45, 263.45, 
    266.75, 265.75, 265.25, 264.85, 264.85, 265.35, 266.35, 266.75, 265.35, 
    264.95, 265.15, 265.35, 265.45, 265.55, 264.75, 264.75, 264.15, 263.75, 
    264.25, 266.35, 265.85, 265.25, 265.75, 266.35, 266.35, 266.75, 266.55, 
    266.95, 266.75, 267.75, 268.05, 270.35, 270.45, 270.45, 270.55, 270.55, 
    270.15, 270.35, 270.35, 270.45, 270.15, 270.05, 269.95, 269.85, 268.75, 
    268.15, 267.75, 267.65, 268.05, 270.25, 270.75, 270.85, 271.05, 271.15, 
    270.95, 270.75, 270.55, 270.85, 270.45, 270.65, 271.05, 270.75, 270.65, 
    270.35, 269.75, 270.45, 270.45, 270.45, 270.65, 271.05, 271.15, 270.25, 
    270.95, 270.85, 271.05, 271.65, 272.25, 272.55, 272.25, 272.15, 271.85, 
    271.05, 270.75, 270.35, 270.25, 269.85, 270.15, 269.85, 270.55, 270.15, 
    270.35, 269.85, 269.65, 269.85, 269.25, 269.25, 269.35, 269.35, 269.15, 
    268.95, 268.85, 268.75, 268.75, 268.65, 268.75, 268.55, 268.45, 268.65, 
    268.55, 268.45, 268.55, 268.35, 268.45, 268.55, 268.75, 268.55, 268.85, 
    269.05, 269.15, 269.35, 269.55, 269.95, 270.05, 270.25, 269.95, 270.45, 
    269.95, 269.45, 269.65, 270.05, 269.45, 269.65, 270.25, 270.45, 270.85, 
    270.95, 270.95, 270.85, 271.25, 271.75, 271.85, 271.65, 271.75, 272.35, 
    272.55, 273.05, 272.15, 272.85, 273.45, 273.15, 273.45, 273.75, 274.15, 
    273.95, 273.55, 273.05, 272.95, 272.55, 272.55, 272.65, 272.35, 272.65, 
    272.55, 273.05, 272.95, 273.65, 274.15, 274.65, 274.85, 274.95, 274.55, 
    274.65, 274.95, 274.65, 274.65, 274.55, 275.15, 273.65, 275.05, 275.45, 
    275.75, 274.45, 273.75, 273.55, 273.75, 273.45, 273.75, 273.45, 273.65, 
    273.85, 273.95, 274.15, 274.35, 274.15, 273.35, 272.85, 272.95, 272.75, 
    272.05, 272.95, 272.85, 272.55, 272.55, 272.55, 272.65, 272.65, 272.55, 
    272.65, 272.95, 273.85, 274.35, 274.45, 274.25, 273.95, 271.75, 273.85, 
    274.05, 273.95, 273.25, 272.85, 272.35, 271.25, 271.05, 270.55, 270.15, 
    270.35, 271.55, 271.85, 271.65, 271.55, 271.75, 271.65, 272.45, 272.35, 
    272.25, 272.15, 271.85, 271.75, 271.55, 271.15, 271.25, 272.05, 272.65, 
    272.55, 272.35, 272.15, 271.95, 271.55, 271.75, 271.35, 270.15, 268.65, 
    269.05, 269.85, 270.15, 269.85, 269.05, 269.05, 268.85, 268.25, 268.65, 
    268.65, 268.65, 268.65, 268.95, 268.65, 269.75, 270.75, 272.55, 272.75, 
    272.45, 271.65, 271.75, 271.55, 274.45, 273.85, 272.95, 272.85, 272.85, 
    273.05, 273.55, 273.15, 273.05, 272.95, 272.15, 271.85, 271.65, 271.45, 
    271.15, 270.55, 270.55, 270.45, 270.35, 270.25, 270.45, 271.05, 271.25, 
    271.15, 271.55, 271.85, 271.65, 271.45, 271.15, 271.15, 271.25, 271.15, 
    271.05, 270.65, 270.15, 269.85, 269.75, 269.85, 268.45, 268.25, 268.05, 
    268.25, 268.05, 269.05, 268.25, 268.25, 267.85, 266.85, 267.85, 268.65, 
    267.65, 265.95, 266.25, 265.55, 264.45, 263.95, 264.55, 263.35, 265.15, 
    264.95, 264.75, 264.45, 264.05, 263.85, 263.35, 263.55, 263.45, 263.65, 
    263.25, 264.65, 263.85, 263.25, 262.65, 262.65, 262.75, 262.45, 262.65, 
    262.75, 263.55, 264.15, 262.75, 264.15, 264.65, 264.45, 263.55, 265.05, 
    264.75, 264.75, 263.95, 263.75, 262.75, 262.75, 262.55, 261.55, 262.15, 
    261.65, 261.85, 261.85, 261.35, 261.55, 261.35, 260.95, 260.75, 261.35, 
    260.45, 261.35, 262.25, 261.95, 262.65, 262.95, 263.05, 263.15, 263.25, 
    263.45, 263.15, 263.55, 264.05, 265.35, 265.65, 266.15, 265.95, 264.95, 
    263.35, 261.55, 262.15, 261.65, 260.45, 260.95, 260.65, 260.55, 261.35, 
    261.15, 260.45, 260.25, 261.45, 261.25, 262.85, 262.35, 262.55, 262.25, 
    261.95, 261.75, 261.55, 260.95, 260.65, 260.55, 260.05, 260.05, 259.75, 
    259.55, 259.55, 259.25, 259.15, 258.85, 256.75, 256.95, 257.05, 256.95, 
    256.95, 255.65, 255.55, 256.15, 255.95, 256.15, 254.85, 254.95, 255.65, 
    254.55, 255.05, 256.85, 254.65, 254.55, 254.25, 254.05, 254.15, 253.35, 
    253.55, 253.25, 253.15, 252.85, 253.65, 253.45, 253.95, 253.35, 253.35, 
    252.95, 253.25, 253.55, 253.75, 253.55, 253.65, 254.45, 253.95, 255.15, 
    255.35, 254.95, 254.95, 255.35, 254.95, 254.75, 255.65, 256.65, 256.25, 
    256.55, 256.85, 257.25, 257.75, 258.25, 258.25, 257.65, 258.15, 259.05, 
    259.15, 259.35, 260.55, 260.35, 260.55, 260.55, 260.15, 260.55, 261.05, 
    261.05, 261.45, 261.35, 261.25, 260.55, 260.35, 259.95, 260.35, 258.85, 
    259.75, 259.85, 260.15, 260.85, 262.15, 261.85, 262.05, 262.95, 263.15, 
    262.95, 262.65, 262.65, 262.25, 262.65, 264.15, 263.35, 263.15, 263.65, 
    264.25, 264.15, 263.85, 263.55, 263.05, 261.05, 260.75, 260.15, 261.75, 
    258.15, 258.55, 259.95, 259.15, 258.25, 257.65, 257.95, 257.85, 257.95, 
    257.85, 256.65, 257.35, 257.05, 256.25, 257.25, 257.45, 257.75, 257.85, 
    257.85, 258.25, 259.15, 260.65, 260.65, 260.95, 260.15, 258.65, 258.05, 
    258.75, 261.05, 262.65, 262.35, 262.25, 261.95, 262.45, 262.75, 263.25, 
    263.45, 262.75, 263.55, 263.65, 264.25, 264.05, 264.65, 264.95, 265.55, 
    265.95, 266.75, 267.45, 268.15, 268.55, 268.65, 269.05, 269.35, 269.95, 
    269.45, 269.35, 269.55, 269.95, 269.95, 269.85, 269.95, 269.95, 269.85, 
    270.15, 270.25, 270.55, 271.05, 271.25, 271.45, 271.25, 271.25, 271.35, 
    271.55, 272.05, 271.45, 271.55, 271.45, 270.85, 270.85, 271.25, 271.55, 
    271.25, 271.85, 272.45, 272.55, 272.95, 272.95, 272.05, 271.75, 272.25, 
    272.25, 272.45, 272.75, 273.05, 273.15, 272.85, 273.55, 273.85, 272.95, 
    273.55, 272.95, 273.25, 273.35, 272.65, 272.95, 272.55, 272.25, 272.25, 
    272.35, 272.95, 272.05, 271.75, 272.25, 271.95, 271.65, 271.05, 268.15, 
    268.25, 268.25, 267.25, 267.05, 267.55, 267.35, 266.35, 267.85, 267.45, 
    267.45, 266.55, 267.35, 267.45, 269.25, 270.35, 267.45, 268.85, 267.25, 
    267.25, 266.75, 267.05, 267.35, 267.45, 268.85, 268.95, 268.55, 267.45, 
    265.35, 264.05, 264.45, 263.75, 263.75, 263.55, 263.45, 264.55, 263.85, 
    264.35, 265.05, 263.75, 263.35, 263.55, 264.05, 264.15, 263.95, 265.65, 
    265.55, 265.25, 264.95, 264.85, 265.45, 265.85, 265.85, 265.85, 265.95, 
    266.25, 265.75, 265.95, 266.05, 266.65, 267.15, 268.15, 268.45, 269.45, 
    270.15, 270.15, 270.45, 269.95, 269.35, 269.95, 268.65, 269.05, 268.85, 
    268.75, 268.85, 268.75, 269.35, 269.05, 269.05, 268.95, 268.85, 269.35, 
    269.05, 268.55, 268.95, 268.65, 268.75, 268.75, 269.05, 269.25, 268.55, 
    268.15, 267.45, 266.85, 266.55, 266.15, 265.75, 265.75, 265.35, 264.85, 
    264.65, 264.65, 264.15, 263.95, 263.55, 263.05, 262.65, 262.15, 261.95, 
    261.65, 261.65, 261.35, 260.95, 260.55, 260.35, 260.15, 259.75, 259.55, 
    259.35, 259.15, 258.95, 259.05, 259.05, 258.95, 258.75, 258.45, 258.45, 
    257.35, 257.95, 257.45, 257.05, 256.95, 256.75, 256.85, 257.25, 256.95, 
    256.85, 256.75, 256.75, 256.75, 256.85, 257.05, 255.35, 255.55, 255.45, 
    255.25, 254.65, 255.95, 255.95, 255.55, 255.25, 254.75, 255.45, 254.35, 
    252.95, 254.95, 255.55, 255.35, 256.15, 256.35, 256.55, 257.35, 258.55, 
    259.65, 260.65, 261.55, 261.55, 262.45, 262.05, 262.25, 263.25, 263.65, 
    265.95, 267.35, 268.25, 268.75, 268.85, 269.15, 269.25, 269.85, 269.65, 
    269.45, 269.25, 268.55, 271.75, 272.85, 273.75, 274.35, 274.95, 275.45, 
    275.25, 274.55, 274.45, 274.65, 275.85, 274.35, 274.45, 273.85, 274.35, 
    274.05, 274.15, 274.55, 274.65, 275.25, 274.35, 273.85, 275.45, 280.35, 
    280.85, 280.85, 279.75, 280.15, 280.45, 279.95, 279.75, 277.85, 278.15, 
    277.85, 277.95, 277.15, 275.95, 276.95, 275.65, 275.65, 275.35, 274.45, 
    275.25, 275.15, 275.25, 275.35, 276.15, 274.85, 274.05, 275.25, 273.95, 
    277.65, 275.15, 276.35, 278.55, 278.35, 278.95, 278.15, 279.25, 278.65, 
    278.45, 278.15, 277.15, 277.65, 277.45, 277.55, 275.85, 276.45, 276.35, 
    277.05, 276.75, 276.65, 276.45, 277.05, 277.85, 277.25, 278.15, 276.75, 
    276.65, 276.15, 276.15, 276.15, 275.55, 276.45, 276.25, 275.45, 276.75, 
    276.15, 275.95, 276.05, 274.85, 275.45, 275.85, 275.85, 275.55, 276.05, 
    276.25, 276.25, 276.45, 277.55, 278.45, 276.85, 276.55, 275.95, 275.75, 
    276.15, 276.25, 275.65, 275.25, 276.35, 275.65, 274.75, 273.65, 273.55, 
    274.95, 275.15, 275.15, 275.45, 276.15, 275.65, 275.85, 276.05, 275.45, 
    274.45, 274.45, 275.25, 276.05, 276.75, 277.45, 277.35, 277.15, 277.65, 
    278.25, 277.65, 277.35, 278.15, 277.75, 277.15, 277.95, 276.95, 276.05, 
    276.75, 276.35, 276.05, 275.15, 274.25, 273.55, 273.15, 272.85, 272.15, 
    272.35, 272.25, 272.25, 272.35, 272.35, 272.55, 272.45, 272.45, 272.35, 
    271.95, 272.05, 271.95, 272.15, 272.35, 272.25, 272.45, 272.15, 271.95, 
    271.85, 271.75, 270.55, 270.05, 269.95, 268.95, 268.15, 267.75, 267.95, 
    267.85, 268.75, 268.75, 268.15, 268.25, 268.05, 267.85, 267.45, 267.15, 
    267.15, 266.65, 266.75, 265.95, 266.15, 265.95, 265.35, 265.15, 264.75, 
    264.15, 263.75, 263.65, 263.15, 263.25, 263.15, 263.15, 263.55, 263.65, 
    263.65, 263.95, 263.65, 263.65, 263.55, 263.25, 263.15, 263.35, 262.65, 
    263.15, 262.95, 263.25, 263.05, 263.45, 263.85, 264.05, 265.15, 265.35, 
    264.95, 266.25, 266.95, 267.15, 266.55, 266.75, 266.65, 266.85, 266.85, 
    266.45, 266.15, 266.15, 265.85, 265.45, 264.75, 264.15, 263.15, 262.65, 
    262.55, 262.25, 262.35, 262.15, 260.75, 260.15, 260.05, 260.55, 262.05, 
    263.15, 263.75, 264.25, 264.35, 264.55, 264.95, 265.25, 265.75, 265.95, 
    265.95, 265.95, 265.85, 265.95, 266.05, 266.15, 266.25, 266.05, 266.15, 
    266.15, 266.05, 265.95, 265.95, 265.85, 265.65, 265.35, 263.55, 263.75, 
    263.55, 264.25, 264.55, 266.35, 265.95, 266.25, 266.05, 266.15, 264.45, 
    266.25, 266.35, 266.15, 265.75, 265.55, 265.35, 262.35, 263.55, 263.65, 
    263.65, 262.45, 262.15, 262.45, 262.75, 263.15, 263.25, 265.25, 265.35, 
    265.65, 265.05, 264.75, 266.05, 265.55, 263.65, 265.05, 266.25, 266.65, 
    266.35, 266.55, 266.55, 266.65, 266.75, 267.05, 267.05, 266.95, 266.65, 
    266.55, 266.65, 266.35, 266.15, 266.25, 266.55, 266.35, 266.25, 266.25, 
    266.15, 266.35, 266.35, 266.25, 264.75, 264.65, 264.15, 263.35, 265.05, 
    264.75, 263.75, 263.75, 263.65, 262.45, 263.75, 263.75, 263.75, 261.95, 
    263.25, 261.95, 262.65, 262.15, 261.65, 262.05, 261.75, 261.15, 261.35, 
    261.95, 261.65, 261.65, 260.75, 261.95, 261.45, 261.25, 261.65, 261.65, 
    261.25, 260.75, 261.35, 260.55, 261.55, 260.65, 260.95, 261.65, 261.75, 
    261.45, 260.95, 261.55, 262.15, 262.45, 262.15, 262.45, 262.35, 263.25, 
    262.75, 262.85, 263.55, 263.85, 264.75, 264.35, 266.45, 265.45, 266.25, 
    265.95, 267.75, 267.05, 266.45, 267.45, 267.35, 267.45, 267.35, 267.15, 
    266.65, 266.35, 266.25, 265.75, 265.55, 265.25, 264.45, 264.95, 264.75, 
    264.15, 264.15, 264.05, 263.65, 263.75, 263.75, 264.05, 264.45, 264.65, 
    264.55, 264.85, 265.15, 265.35, 265.45, 266.05, 266.05, 266.75, 266.15, 
    266.75, 266.75, 266.95, 266.05, 269.15, 267.45, 267.65, 267.75, 267.85, 
    268.15, 268.45, 269.75, 270.15, 270.75, 271.25, 271.15, 270.55, 271.45, 
    271.25, 270.45, 270.55, 270.75, 271.65, 272.15, 271.75, 271.65, 271.65, 
    271.85, 271.55, 271.15, 271.35, 271.25, 268.55, 270.65, 267.95, 267.65, 
    267.65, 269.25, 268.85, 265.75, 265.85, 267.15, 264.95, 265.95, 266.65, 
    267.05, 268.05, 269.05, 269.35, 269.55, 269.05, 269.45, 269.95, 269.35, 
    269.45, 270.15, 271.85, 271.95, 271.85, 271.65, 271.35, 271.05, 271.05, 
    271.25, 270.85, 270.65, 270.35, 270.05, 269.85, 269.75, 269.45, 267.95, 
    267.85, 267.95, 269.15, 268.45, 268.05, 269.45, 270.85, 271.95, 271.35, 
    271.45, 270.35, 269.55, 271.55, 271.55, 271.35, 270.95, 270.95, 270.75, 
    270.15, 269.35, 269.25, 268.25, 268.35, 267.25, 267.25, 266.75, 266.25, 
    265.95, 266.75, 265.15, 266.85, 266.45, 265.85, 266.85, 267.15, 266.85, 
    266.05, 266.45, 265.05, 265.95, 266.95, 266.25, 266.45, 266.75, 266.45, 
    267.15, 267.55, 267.35, 266.85, 265.75, 264.05, 264.45, 263.85, 263.65, 
    261.75, 260.75, 261.55, 259.65, 260.45, 260.55, 260.55, 260.15, 260.25, 
    260.05, 261.95, 261.55, 262.25, 263.05, 263.35, 264.05, 264.25, 264.45, 
    264.85, 265.25, 265.95, 266.35, 266.65, 266.85, 266.95, 266.95, 268.25, 
    268.45, 268.15, 269.25, 268.75, 268.95, 269.15, 268.85, 269.25, 269.15, 
    269.25, 269.55, 269.05, 270.05, 270.15, 270.45, 269.65, 270.35, 270.45, 
    270.55, 270.95, 270.85, 271.25, 271.45, 270.95, 270.75, 270.75, 270.85, 
    270.45, 271.05, 270.65, 270.95, 271.45, 271.35, 271.45, 271.65, 271.55, 
    272.05, 271.45, 271.45, 270.85, 270.95, 270.95, 271.95, 272.45, 272.15, 
    271.75, 271.65, 271.85, 272.25, 272.65, 272.85, 272.85, 273.35, 273.55, 
    273.15, 272.55, 272.35, 274.85, 272.75, 274.65, 276.35, 276.05, 275.95, 
    275.75, 275.15, 274.85, 275.45, 275.05, 274.45, 273.85, 273.65, 273.95, 
    273.75, 274.05, 273.95, 273.95, 273.85, 273.55, 273.65, 273.35, 273.35, 
    272.85, 273.05, 273.15, 273.05, 272.95, 272.45, 272.55, 272.45, 272.45, 
    272.55, 272.05, 271.65, 271.45, 271.45, 270.45, 270.45, 270.55, 270.55, 
    270.55, 270.55, 270.45, 270.25, 270.25, 270.15, 269.65, 269.75, 269.65, 
    269.85, 269.75, 269.65, 269.75, 269.85, 269.75, 269.85, 269.65, 269.55, 
    269.25, 269.55, 269.25, 269.05, 269.05, 268.85, 269.15, 269.15, 268.75, 
    268.75, 268.65, 268.25, 268.65, 268.55, 268.75, 268.45, 268.15, 268.05, 
    268.35, 268.25, 268.55, 268.35, 268.45, 268.45, 268.45, 268.25, 267.75, 
    267.45, 268.25, 267.75, 267.85, 267.45, 266.95, 267.35, 268.15, 268.25, 
    268.85, 269.35, 268.65, 268.35, 268.65, 268.25, 268.35, 268.15, 268.05, 
    268.45, 268.45, 268.55, 268.25, 268.25, 267.95, 267.65, 267.55, 267.55, 
    267.65, 266.95, 265.55, 265.75, 264.15, 263.05, 262.95, 264.05, 263.05, 
    263.35, 263.45, 262.75, 263.25, 263.45, 264.95, 266.25, 266.35, 266.65, 
    267.55, 269.05, 271.65, 273.75, 274.25, 273.25, 274.85, 275.05, 274.85, 
    274.25, 274.25, 273.85, 273.65, 273.65, 274.25, 273.95, 273.85, 273.35, 
    272.65, 272.55, 272.05, 271.95, 270.95, 270.95, 271.05, 270.85, 271.25, 
    271.15, 270.65, 270.15, 270.45, 270.25, 269.95, 269.95, 270.05, 270.15, 
    270.45, 270.65, 270.65, 270.55, 270.85, 271.05, 271.35, 271.15, 271.15, 
    271.25, 271.05, 270.95, 271.45, 272.15, 272.25, 272.85, 272.05, 272.45, 
    272.25, 271.85, 272.05, 271.75, 271.65, 271.65, 271.55, 271.75, 271.65, 
    271.65, 271.65, 271.75, 271.85, 271.65, 271.35, 271.65, 271.15, 271.15, 
    270.65, 270.25, 270.45, 270.75, 270.25, 270.25, 270.25, 269.45, 270.15, 
    270.05, 269.95, 269.45, 268.55, 267.75, 267.25, 267.15, 267.05, 267.35, 
    267.45, 267.45, 266.55, 267.25, 267.05, 267.05, 267.15, 267.25, 267.45, 
    267.55, 267.55, 267.45, 267.05, 266.75, 266.45, 266.55, 266.15, 266.35, 
    266.05, 265.45, 265.75, 266.15, 266.85, 267.55, 268.25, 268.55, 268.75, 
    269.35, 269.65, 269.75, 269.75, 269.25, 269.45, 268.45, 268.35, 268.25, 
    267.85, 268.05, 268.05, 267.75, 267.35, 267.25, 266.65, 266.55, 265.85, 
    265.55, 263.25, 263.25, 263.45, 262.75, 263.65, 263.25, 262.75, 263.45, 
    262.65, 262.95, 263.25, 263.65, 262.95, 262.85, 263.45, 263.25, 262.95, 
    262.85, 262.75, 262.75, 262.45, 263.05, 263.25, 262.95, 263.35, 263.15, 
    263.35, 263.35, 263.35, 263.55, 263.55, 263.65, 263.75, 263.75, 263.35, 
    262.65, 260.65, 260.75, 260.75, 259.35, 260.35, 260.35, 260.95, 260.95, 
    261.45, 260.05, 260.25, 260.65, 260.05, 259.95, 259.95, 259.45, 259.35, 
    258.85, 260.05, 259.05, 258.15, 258.65, 258.85, 259.35, 258.95, 258.45, 
    258.85, 258.65, 260.75, 259.05, 260.55, 260.45, 258.85, 260.05, 259.85, 
    260.75, 262.15, 261.55, 260.75, 260.05, 261.15, 261.65, 261.85, 262.15, 
    263.85, 264.35, 263.55, 262.75, 262.25, 263.95, 264.35, 263.95, 263.75, 
    263.65, 263.65, 263.85, 263.55, 261.05, 262.05, 260.55, 262.25, 262.55, 
    262.65, 260.75, 262.55, 262.25, 262.65, 262.95, 263.45, 263.75, 263.95, 
    264.05, 264.65, 264.15, 265.25, 266.05, 267.05, 267.45, 267.55, 268.05, 
    268.55, 268.65, 269.15, 269.15, 269.45, 269.35, 269.25, 269.25, 269.15, 
    268.95, 268.75, 267.95, 267.25, 266.95, 266.25, 265.85, 265.35, 264.85, 
    264.45, 264.05, 263.65, 262.75, 263.15, 261.55, 261.45, 260.55, 259.65, 
    261.05, 260.45, 260.25, 260.05, 259.85, 259.25, 259.75, 259.45, 259.35, 
    259.15, 258.85, 259.05, 259.35, 259.55, 258.95, 259.05, 258.65, 258.65, 
    259.35, 259.25, 259.15, 259.45, 259.85, 259.35, 259.55, 259.85, 260.05, 
    260.95, 259.55, 260.85, 261.25, 261.75, 262.05, 262.85, 262.95, 262.75, 
    262.55, 261.75, 261.45, 261.35, 261.55, 261.05, 260.85, 260.75, 261.15, 
    261.65, 259.95, 260.95, 260.35, 260.75, 260.25, 260.05, 260.35, 260.75, 
    260.95, 260.95, 260.85, 261.45, 260.75, 261.95, 261.25, 260.65, 261.75, 
    261.15, 261.35, 259.15, 258.65, 257.85, 258.55, 258.35, 258.55, 259.15, 
    259.85, 258.75, 260.45, 260.75, 261.05, 261.95, 262.05, 263.75, 264.35, 
    264.55, 264.15, 265.15, 264.55, 264.85, 267.15, 268.55, 267.45, 266.45, 
    268.25, 271.15, 270.55, 270.35, 271.05, 271.05, 270.95, 270.85, 271.35, 
    270.95, 270.95, 270.85, 270.75, 270.75, 271.05, 271.45, 271.85, 271.95, 
    271.65, 271.95, 272.25, 272.15, 272.05, 272.35, 272.45, 272.65, 272.15, 
    271.65, 271.35, 272.55, 272.65, 272.65, 273.65, 272.25, 272.15, 272.15, 
    271.25, 271.35, 270.95, 271.15, 270.85, 270.45, 271.45, 269.35, 269.95, 
    270.15, 270.85, 270.65, 270.75, 271.55, 271.35, 271.45, 270.85, 270.95, 
    271.15, 270.65, 270.35, 270.45, 270.65, 270.15, 269.95, 270.15, 269.35, 
    269.55, 268.95, 268.75, 268.95, 269.45, 269.65, 269.95, 269.95, 269.85, 
    270.35, 270.55, 270.65, 270.45, 271.15, 270.15, 270.55, 270.15, 270.75, 
    270.65, 270.75, 270.75, 270.85, 270.75, 270.75, 270.85, 271.05, 270.05, 
    269.75, 269.85, 269.15, 269.15, 269.55, 269.75, 270.15, 270.35, 270.05, 
    269.85, 270.85, 270.55, 270.75, 270.25, 269.75, 270.55, 272.15, 274.45, 
    272.85, 272.05, 272.35, 272.15, 272.95, 272.95, 272.05, 270.55, 270.15, 
    269.65, 267.45, 266.65, 267.65, 267.75, 267.05, 267.45, 266.95, 266.65, 
    267.25, 266.55, 266.05, 267.35, 268.65, 267.65, 269.35, 269.05, 268.85, 
    267.85, 269.35, 269.45, 270.85, 269.75, 270.65, 271.65, 271.25, 271.05, 
    270.85, 270.45, 270.15, 270.45, 268.75, 268.55, 269.45, 268.45, 270.25, 
    269.65, 269.55, 269.65, 269.85, 269.45, 269.45, 269.55, 269.45, 269.75, 
    269.45, 270.05, 269.85, 269.35, 268.75, 268.25, 267.75, 267.85, 268.55, 
    270.35, 270.85, 271.45, 271.75, 271.75, 271.75, 273.15, 272.85, 272.45, 
    272.45, 272.45, 272.45, 272.15, 271.95, 272.35, 272.65, 272.85, 272.95, 
    273.05, 273.35, 273.05, 272.95, 272.75, 273.25, 273.35, 273.15, 273.35, 
    274.05, 274.25, 273.75, 273.15, 273.25, 273.85, 273.15, 272.75, 273.75, 
    273.45, 273.45, 273.75, 274.15, 272.65, 273.35, 273.95, 273.35, 273.95, 
    273.65, 273.85, 273.55, 274.65, 273.85, 274.05, 273.65, 273.75, 272.75, 
    273.45, 273.35, 273.25, 273.85, 273.65, 273.55, 273.15, 272.75, 272.55, 
    272.55, 272.55, 272.55, 272.85, 272.35, 272.05, 271.35, 271.25, 271.25, 
    270.65, 270.05, 270.35, 270.05, 267.25, 267.85, 268.25, 267.85, 266.95, 
    267.45, 266.95, 267.25, 266.85, 266.05, 266.45, 266.55, 265.35, 264.25, 
    264.35, 264.65, 263.75, 265.15, 265.25, 264.75, 264.85, 265.65, 265.45, 
    267.05, 265.95, 265.25, 265.75, 266.05, 265.85, 265.35, 266.45, 264.65, 
    264.85, 263.85, 264.85, 264.95, 264.05, 264.65, 263.05, 265.05, 263.25, 
    263.95, 264.05, 264.45, 264.15, 264.55, 265.05, 263.75, 263.55, 262.35, 
    263.55, 262.75, 263.85, 262.75, 262.65, 262.95, 262.85, 263.65, 261.95, 
    263.25, 262.35, 262.65, 262.95, 263.35, 263.25, 264.35, 262.95, 263.05, 
    263.25, 262.75, 262.75, 263.05, 263.55, 263.65, 263.25, 263.55, 263.75, 
    263.55, 263.55, 263.35, 263.35, 262.75, 262.65, 262.95, 263.05, 263.55, 
    264.05, 265.15, 265.05, 264.15, 264.75, 263.85, 263.55, 263.35, 263.85, 
    262.85, 260.95, 261.25, 261.65, 262.35, 262.45, 262.85, 262.95, 262.85, 
    262.75, 263.45, 263.95, 263.65, 263.65, 263.55, 264.25, 264.35, 264.85, 
    265.55, 265.25, 265.75, 265.05, 263.95, 263.35, 264.35, 263.25, 263.95, 
    263.35, 263.25, 264.95, 264.95, 265.35, 266.05, 265.85, 265.75, 267.35, 
    266.75, 266.25, 266.75, 266.35, 266.25, 266.55, 266.55, 266.45, 266.85, 
    266.15, 265.45, 264.75, 264.65, 264.45, 263.35, 263.25, 264.35, 264.55, 
    265.25, 264.75, 266.05, 269.55, 270.25, 271.05, 271.45, 272.45, 271.55, 
    272.45, 270.95, 270.35, 271.35, 270.85, 271.75, 271.45, 271.35, 272.55, 
    271.95, 273.05, 273.35, 274.45, 275.25, 275.85, 275.05, 274.65, 274.65, 
    274.15, 273.45, 273.45, 273.55, 273.55, 274.05, 273.05, 273.15, 273.45, 
    273.75, 273.85, 273.75, 273.15, 272.45, 272.55, 272.35, 272.35, 272.75, 
    273.15, 273.35, 272.85, 273.35, 274.65, 272.55, 272.85, 271.85, 272.55, 
    272.85, 272.55, 271.95, 271.95, 270.45, 272.45, 274.95, 275.45, 275.55, 
    274.25, 273.95, 274.55, 274.35, 273.85, 272.85, 272.35, 272.15, 272.35, 
    271.35, 271.65, 271.35, 271.25, 271.25, 271.25, 271.15, 270.25, 270.15, 
    269.45, 268.45, 268.65, 267.75, 267.95, 268.35, 269.35, 269.35, 270.45, 
    270.05, 270.35, 270.85, 271.25, 271.45, 271.55, 271.45, 271.55, 271.65, 
    271.55, 271.35, 271.25, 271.25, 270.85, 270.85, 271.05, 270.65, 270.55, 
    270.45, 270.25, 270.15, 269.45, 269.75, 269.05, 269.35, 268.25, 267.35, 
    267.95, 268.35, 268.45, 268.65, 268.45, 268.25, 268.45, 268.45, 268.35, 
    268.45, 268.45, 268.55, 268.95, 269.15, 268.95, 269.25, 268.45, 268.25, 
    267.25, 267.85, 268.15, 268.15, 267.85, 268.25, 267.05, 267.45, 267.25, 
    268.15, 268.75, 269.05, 268.45, 268.05, 267.15, 267.55, 265.95, 267.45, 
    265.65, 265.75, 266.35, 267.35, 265.95, 267.85, 267.55, 267.95, 268.35, 
    267.35, 267.25, 265.95, 265.35, 264.85, 265.65, 264.35, 266.15, 265.65, 
    266.15, 266.45, 265.85, 265.05, 265.25, 266.75, 268.65, 269.05, 268.65, 
    268.35, 268.05, 268.95, 269.85, 269.55, 269.05, 269.15, 266.85, 267.15, 
    265.75, 265.25, 265.25, 265.75, 264.95, 264.55, 264.35, 264.05, 264.75, 
    265.85, 266.55, 266.65, 266.75, 266.35, 266.65, 266.55, 266.65, 266.25, 
    266.15, 265.55, 265.55, 265.55, 266.35, 267.75, 268.05, 267.95, 267.85, 
    267.85, 268.75, 267.55, 268.55, 269.25, 269.45, 269.25, 269.75, 270.55, 
    270.55, 270.05, 270.35, 271.65, 272.45, 271.15, 271.05, 269.95, 269.55, 
    270.85, 271.65, 271.15, 272.05, 273.05, 272.75, 272.65, 273.15, 273.75, 
    273.65, 273.85, 273.15, 272.95, 272.55, 272.75, 273.95, 273.75, 272.95, 
    274.25, 274.35, 275.25, 275.35, 275.75, 275.25, 275.45, 276.35, 276.35, 
    276.45, 275.45, 275.55, 275.05, 275.35, 276.05, 275.55, 276.55, 276.05, 
    276.35, 275.55, 274.65, 275.25, 275.15, 275.05, 275.35, 277.15, 276.05, 
    276.15, 275.95, 275.35, 275.25, 275.05, 274.85, 275.05, 274.65, 274.65, 
    274.35, 273.95, 272.15, 270.35, 269.95, 269.35, 269.35, 267.05, 266.55, 
    266.35, 265.55, 265.05, 265.05, 264.75, 265.55, 266.15, 266.15, 266.55, 
    266.95, 267.15, 266.45, 266.15, 266.25, 267.25, 267.75, 268.75, 269.15, 
    269.85, 269.55, 269.65, 269.75, 269.15, 271.15, 271.45, 271.45, 271.65, 
    271.35, 271.15, 270.85, 268.95, 268.15, 267.35, 267.05, 266.15, 265.65, 
    265.45, 265.25, 264.85, 264.35, 262.75, 260.85, 261.85, 261.35, 262.95, 
    262.35, 261.65, 260.75, 259.45, 258.95, 258.55, 258.45, 258.35, 258.55, 
    258.15, 257.35, 257.35, 257.65, 257.45, 257.05, 257.15, 257.05, 257.25, 
    256.95, 256.65, 256.05, 256.05, 256.05, 255.75, 255.95, 255.95, 255.85, 
    256.25, 256.25, 256.65, 257.15, 257.55, 257.85, 258.05, 257.85, 257.85, 
    258.35, 258.25, 258.15, 257.85, 257.95, 257.75, 258.15, 257.75, 257.55, 
    257.55, 257.65, 257.95, 257.95, 258.15, 257.65, 256.85, 256.45, 257.15, 
    258.75, 259.15, 258.25, 260.75, 256.95, 258.85, 259.05, 261.35, 259.05, 
    258.75, 259.45, 259.15, 258.25, 261.35, 261.45, 258.65, 259.95, 258.35, 
    259.15, 257.05, 259.65, 258.85, 257.55, 259.65, 260.15, 259.05, 260.95, 
    262.05, 259.05, 259.75, 259.45, 261.45, 259.25, 257.95, 257.75, 258.65, 
    259.05, 258.65, 257.95, 258.55, 259.25, 257.65, 258.25, 256.75, 256.65, 
    257.15, 258.65, 258.15, 258.05, 258.45, 259.35, 258.45, 257.65, 257.85, 
    257.65, 257.65, 257.45, 256.95, 256.95, 257.85, 256.95, 257.25, 257.25, 
    257.45, 257.75, 257.75, 257.85, 257.85, 258.45, 258.75, 257.95, 257.55, 
    257.25, 258.45, 258.85, 259.35, 258.05, 259.55, 258.55, 258.15, 257.05, 
    257.05, 256.65, 255.75, 255.55, 254.65, 255.35, 254.65, 255.25, 255.05, 
    254.45, 255.15, 254.05, 255.15, 256.05, 255.35, 256.95, 257.35, 256.45, 
    256.35, 257.25, 257.15, 256.65, 256.45, 256.05, 254.55, 256.85, 255.65, 
    255.05, 255.75, 256.05, 255.95, 255.35, 256.35, 256.85, 257.05, 257.75, 
    258.85, 261.05, 260.65, 260.75, 260.65, 262.35, 261.25, 260.65, 260.25, 
    260.95, 260.95, 260.05, 260.15, 260.65, 260.15, 260.25, 258.35, 258.45, 
    257.65, 257.75, 257.85, 257.25, 256.65, 258.05, 257.95, 259.25, 259.05, 
    259.45, 260.05, 260.15, 259.95, 259.85, 260.85, 259.25, 258.45, 258.45, 
    257.95, 257.45, 256.45, 257.35, 255.85, 256.65, 256.95, 255.95, 256.05, 
    256.95, 257.45, 257.35, 256.85, 257.55, 258.75, 259.95, 259.45, 261.95, 
    260.15, 261.65, 260.45, 260.25, 259.95, 257.65, 258.15, 257.55, 258.85, 
    258.35, 259.15, 257.85, 258.35, 258.75, 258.95, 258.25, 259.25, 258.95, 
    260.15, 260.65, 261.55, 263.05, 263.65, 264.15, 265.05, 264.65, 264.35, 
    264.75, 263.75, 263.35, 263.15, 262.15, 262.75, 262.15, 262.85, 263.65, 
    263.85, 264.95, 265.05, 265.75, 266.65, 269.15, 269.65, 269.65, 270.35, 
    270.35, 270.35, 270.05, 270.55, 271.35, 270.85, 271.75, 272.15, 272.55, 
    272.65, 272.75, 273.35, 273.15, 273.75, 272.75, 273.15, 272.85, 271.95, 
    274.25, 274.55, 273.35, 273.35, 273.75, 273.55, 274.75, 274.65, 273.35, 
    273.85, 274.15, 273.75, 273.35, 272.75, 272.65, 272.25, 272.05, 272.15, 
    271.35, 270.65, 269.95, 269.15, 268.85, 268.55, 268.35, 268.55, 268.25, 
    268.25, 268.45, 268.95, 267.75, 266.75, 268.15, 267.45, 268.15, 268.15, 
    267.95, 265.05, 266.55, 265.05, 265.65, 265.95, 265.35, 265.75, 266.15, 
    266.25, 267.15, 266.85, 265.85, 267.25, 267.75, 267.95, 267.05, 265.75, 
    264.95, 267.45, 269.55, 269.75, 269.35, 269.55, 270.05, 270.55, 270.25, 
    270.25, 270.35, 270.15, 270.35, 270.35, 270.25, 270.15, 269.95, 269.85, 
    269.65, 269.55, 269.75, 269.85, 269.85, 269.85, 270.05, 269.85, 269.75, 
    269.55, 269.05, 268.65, 268.35, 267.85, 267.55, 267.65, 266.55, 266.65, 
    266.65, 264.45, 264.15, 263.15, 264.15, 261.95, 261.55, 260.25, 261.35, 
    262.15, 262.55, 263.75, 263.25, 263.55, 264.05, 264.95, 266.45, 263.45, 
    263.65, 263.55, 262.75, 261.25, 260.95, 260.75, 261.35, 262.45, 261.45, 
    263.35, 262.95, 263.15, 263.35, 263.35, 264.25, 264.05, 264.85, 265.25, 
    266.25, 265.85, 265.75, 266.55, 266.55, 266.95, 266.45, 266.85, 266.55, 
    266.75, 266.45, 267.05, 267.05, 266.95, 266.65, 267.65, 267.65, 267.35, 
    266.75, 267.65, 268.25, 268.65, 268.55, 269.05, 269.65, 268.85, 271.25, 
    271.15, 271.45, 271.45, 271.35, 271.55, 271.25, 271.35, 270.75, 270.55, 
    270.45, 270.45, 269.05, 268.35, 269.65, 270.65, 271.45, 271.55, 271.55, 
    271.55, 271.25, 271.75, 271.75, 272.15, 271.45, 271.15, 270.65, 269.55, 
    269.15, 269.35, 269.35, 268.95, 268.75, 268.95, 268.65, 268.65, 268.45, 
    268.45, 267.95, 267.85, 267.85, 267.75, 267.85, 267.65, 267.55, 267.75, 
    267.75, 267.65, 267.95, 268.05, 267.75, 267.85, 267.35, 267.05, 267.45, 
    267.05, 266.85, 266.35, 266.35, 266.05, 265.95, 265.95, 265.65, 261.95, 
    261.65, 262.65, 261.75, 263.35, 265.05, 265.55, 266.95, 265.65, 267.15, 
    267.35, 268.35, 267.55, 267.15, 266.45, 267.95, 267.95, 267.25, 267.45, 
    268.25, 267.65, 267.95, 268.15, 267.85, 268.25, 268.25, 268.45, 268.45, 
    268.95, 268.75, 270.35, 269.55, 270.45, 270.45, 270.65, 270.65, 270.15, 
    271.45, 270.55, 270.45, 269.55, 269.55, 269.35, 269.35, 269.05, 268.85, 
    269.25, 268.95, 268.95, 268.65, 268.85, 268.95, 268.75, 268.95, 269.45, 
    269.55, 270.15, 270.15, 270.35, 271.05, 270.45, 270.15, 269.95, 269.15, 
    268.85, 268.55, 268.25, 268.35, 268.45, 268.75, 268.35, 267.75, 268.45, 
    268.25, 268.05, 268.75, 268.65, 268.35, 269.65, 269.15, 269.25, 268.85, 
    269.15, 269.85, 269.45, 269.55, 269.35, 269.25, 268.55, 268.35, 268.05, 
    267.65, 267.35, 266.75, 266.95, 266.45, 266.15, 265.75, 265.35, 265.35, 
    264.95, 264.75, 264.45, 264.35, 264.45, 263.95, 264.45, 263.75, 262.75, 
    261.95, 262.75, 261.55, 261.25, 256.55, 256.55, 256.65, 259.05, 256.55, 
    257.85, 255.95, 255.15, 254.75, 257.05, 257.25, 257.55, 258.05, 257.95, 
    257.65, 257.85, 258.35, 258.85, 258.85, 258.35, 258.55, 258.45, 259.15, 
    259.75, 259.85, 259.35, 259.15, 257.65, 257.15, 256.25, 257.35, 257.05, 
    257.15, 258.65, 259.65, 259.65, 260.75, 261.05, 261.45, 261.35, 262.05, 
    262.05, 262.25, 262.55, 262.95, 262.55, 261.95, 261.75, 259.65, 258.25, 
    258.75, 259.15, 259.35, 258.65, 258.85, 259.15, 258.45, 257.95, 258.65, 
    259.25, 259.95, 260.35, 260.45, 260.95, 262.65, 261.75, 262.05, 261.55, 
    262.15, 261.85, 261.45, 259.65, 258.25, 257.55, 257.45, 259.15, 259.05, 
    258.75, 258.95, 259.85, 258.65, 260.75, 260.95, 264.25, 264.65, 264.65, 
    266.05, 266.05, 266.05, 265.75, 265.35, 265.35, 265.95, 265.85, 265.95, 
    266.45, 265.85, 265.15, 264.85, 265.05, 263.55, 263.85, 262.65, 262.55, 
    263.45, 263.05, 264.55, 264.85, 264.55, 264.55, 265.05, 264.45, 264.15, 
    264.35, 264.65, 264.45, 264.65, 264.85, 264.65, 264.75, 264.25, 264.35, 
    263.65, 264.05, 263.95, 263.25, 262.25, 261.75, 262.15, 261.85, 263.05, 
    263.25, 263.75, 265.55, 265.85, 265.95, 265.75, 265.25, 265.65, 266.15, 
    265.75, 264.95, 264.35, 264.65, 263.65, 262.35, 262.65, 262.55, 262.75, 
    262.95, 262.25, 261.65, 262.55, 262.15, 263.05, 264.75, 265.25, 265.25, 
    266.15, 266.15, 266.55, 266.75, 266.75, 266.65, 266.15, 266.05, 266.05, 
    265.65, 265.65, 265.05, 265.05, 264.85, 264.95, 265.05, 264.65, 264.75, 
    263.45, 263.15, 264.55, 264.45, 262.95, 263.05, 264.85, 264.85, 265.15, 
    265.05, 264.65, 265.15, 265.65, 264.65, 263.65, 262.95, 262.35, 261.35, 
    260.95, 260.65, 259.85, 260.05, 259.05, 259.45, 259.25, 258.75, 260.55, 
    260.95, 263.65, 262.95, 264.25, 263.25, 263.45, 263.15, 263.05, 263.25, 
    263.05, 263.15, 261.35, 261.35, 260.75, 259.75, 259.25, 260.25, 259.05, 
    259.95, 259.45, 259.45, 260.05, 259.85, 260.75, 261.05, 262.25, 263.45, 
    264.25, 265.55, 264.45, 264.75, 264.95, 265.45, 264.95, 264.35, 264.55, 
    263.55, 261.55, 260.45, 260.95, 261.55, 259.95, 260.15, 259.25, 258.75, 
    260.25, 261.45, 261.25, 262.65, 264.25, 264.35, 263.35, 263.75, 264.25, 
    264.45, 264.25, 265.55, 266.15, 264.65, 265.25, 265.15, 264.85, 264.75, 
    264.95, 264.85, 265.55, 265.25, 265.75, 266.25, 267.05, 268.55, 268.65, 
    268.95, 269.25, 268.65, 269.95, 270.85, 271.15, 270.75, 270.75, 271.35, 
    271.25, 270.25, 269.95, 270.05, 269.55, 269.85, 269.25, 268.85, 269.45, 
    269.45, 269.35, 269.25, 269.45, 269.45, 270.65, 272.35, 272.15, 271.15, 
    273.45, 273.85, 272.85, 274.55, 271.85, 271.55, 271.15, 270.15, 268.65, 
    268.45, 267.35, 266.25, 265.95, 265.45, 266.05, 266.55, 267.25, 266.95, 
    266.25, 266.15, 266.75, 266.85, 266.15, 267.15, 267.55, 268.05, 268.55, 
    268.35, 267.65, 267.95, 266.85, 266.45, 265.65, 265.45, 264.25, 263.15, 
    263.85, 263.15, 262.15, 263.25, 263.55, 263.05, 262.75, 263.15, 262.45, 
    264.05, 265.05, 264.85, 265.45, 265.75, 266.05, 267.15, 265.95, 266.75, 
    267.45, 263.95, 265.75, 266.05, 265.65, 265.35, 265.15, 264.85, 264.65, 
    264.85, 265.15, 265.25, 264.55, 264.55, 264.85, 265.95, 268.05, 266.75, 
    267.85, 269.45, 268.15, 268.55, 268.15, 269.15, 268.15, 268.05, 268.35, 
    268.75, 267.85, 267.25, 267.85, 267.65, 267.85, 268.25, 267.85, 268.05, 
    267.75, 267.55, 267.55, 268.25, 268.65, 271.55, 272.35, 271.05, 271.55, 
    271.75, 273.15, 273.25, 273.05, 272.55, 272.75, 271.75, 270.05, 267.95, 
    268.15, 266.25, 266.75, 266.55, 267.25, 267.35, 265.75, 268.05, 266.85, 
    268.85, 270.95, 273.15, 271.95, 270.95, 271.15, 270.75, 270.25, 270.75, 
    271.25, 271.05, 271.25, 271.25, 269.05, 269.15, 269.25, 268.85, 268.55, 
    268.05, 267.25, 268.05, 267.45, 268.55, 268.75, 269.85, 270.65, 271.05, 
    271.65, 272.35, 273.45, 272.95, 274.75, 273.25, 272.65, 272.55, 272.15, 
    272.45, 271.35, 269.95, 270.05, 268.45, 268.75, 267.45, 267.95, 267.95, 
    266.85, 270.55, 269.05, 270.65, 271.95, 273.85, 274.15, 273.65, 273.45, 
    274.05, 272.85, 274.25, 274.85, 272.95, 272.85, 272.65, 272.25, 270.25, 
    270.45, 270.95, 271.15, 271.45, 271.15, 271.35, 271.85, 271.85, 271.55, 
    272.35, 272.25, 273.15, 272.35, 272.35, 272.55, 273.25, 273.55, 274.35, 
    274.85, 274.85, 275.05, 274.85, 274.95, 274.45, 274.75, 275.35, 275.35, 
    273.35, 273.25, 273.05, 272.85, 272.95, 273.35, 274.45, 275.15, 277.05, 
    277.65, 275.15, 276.05, 275.95, 275.15, 275.05, 274.15, 273.75, 273.85, 
    274.15, 273.65, 273.35, 273.35, 272.95, 272.95, 272.95, 272.85, 272.75, 
    272.85, 272.95, 273.45, 272.95, 272.95, 272.65, 272.75, 272.55, 272.85, 
    272.85, 272.45, 272.55, 272.85, 272.85, 272.55, 272.45, 272.35, 272.05, 
    271.95, 271.55, 271.55, 271.45, 271.45, 271.15, 271.45, 271.15, 271.25, 
    271.25, 271.35, 271.45, 271.55, 271.65, 272.25, 271.65, 271.65, 271.85, 
    271.85, 272.05, 271.95, 271.65, 271.35, 271.35, 270.85, 270.95, 270.95, 
    271.25, 271.55, 271.65, 271.85, 272.25, 272.55, 272.75, 272.65, 272.95, 
    272.75, 272.85, 273.05, 272.15, 271.75, 271.15, 271.05, 270.85, 270.35, 
    269.95, 269.95, 269.85, 269.85, 269.95, 270.35, 270.35, 270.45, 270.65, 
    269.55, 270.05, 270.45, 271.25, 271.85, 272.05, 273.05, 273.35, 274.15, 
    274.35, 273.55, 273.05, 272.85, 273.55, 273.75, 273.65, 273.35, 273.35, 
    273.25, 273.25, 273.25, 273.25, 273.15, 273.15, 273.25, 273.05, 273.05, 
    273.05, 273.35, 273.25, 273.75, 273.55, 273.55, 273.25, 273.75, 273.75, 
    273.35, 273.75, 273.75, 273.45, 273.25, 273.35, 273.15, 273.65, 273.35, 
    274.05, 274.15, 274.25, 273.65, 273.85, 274.25, 274.55, 275.35, 275.55, 
    276.15, 275.55, 275.45, 275.25, 276.05, 276.45, 276.35, 276.85, 277.05, 
    275.25, 275.55, 273.65, 274.05, 273.45, 273.25, 273.35, 272.95, 273.45, 
    273.05, 273.25, 273.25, 273.35, 273.95, 273.35, 273.85, 274.15, 274.55, 
    273.45, 273.95, 273.55, 273.85, 273.55, 273.95, 273.45, 273.25, 273.15, 
    272.95, 273.65, 273.65, 273.45, 273.65, 273.45, 273.35, 273.25, 273.45, 
    273.75, 274.05, 273.25, 273.25, 272.65, 273.05, 274.35, 273.65, 273.35, 
    274.15, 274.35, 274.45, 273.75, 273.55, 273.75, 273.35, 273.25, 273.45, 
    273.15, 273.15, 272.95, 274.15, 274.75, 274.25, 274.35, 274.45, 274.55, 
    274.75, 274.15, 274.65, 275.25, 275.15, 275.25, 275.35, 275.05, 274.65, 
    274.45, 274.25, 273.85, 273.75, 273.35, 273.45, 273.95, 274.35, 274.95, 
    275.45, 275.85, 275.85, 276.75, 276.55, 277.35, 277.35, 277.15, 276.95, 
    277.15, 276.85, 276.75, 276.85, 276.75, 276.95, 276.45, 276.45, 275.95, 
    275.65, 275.75, 275.65, 275.35, 275.05, 274.75, 274.65, 274.75, 274.55, 
    274.45, 274.45, 274.55, 274.55, 274.75, 274.75, 275.35, 274.95, 274.95, 
    274.85, 274.85, 274.55, 274.65, 274.75, 274.65, 273.95, 273.65, 273.35, 
    273.15, 273.25, 273.55, 273.95, 274.55, 274.45, 274.95, 275.05, 275.55, 
    275.55, 275.85, 275.65, 275.55, 275.65, 274.95, 273.55, 274.25, 275.15, 
    274.85, 275.05, 275.25, 275.15, 275.75, 275.75, 276.25, 275.95, 276.45, 
    276.15, 276.05, 274.75, 274.75, 274.75, 275.05, 274.75, 274.65, 274.35, 
    274.15, 274.15, 274.35, 274.65, 275.05, 274.95, 274.65, 274.25, 274.35, 
    275.25, 274.95, 274.95, 275.05, 274.85, 274.85, 274.85, 275.45, 275.45, 
    275.65, 275.65, 275.85, 276.05, 275.65, 274.95, 275.45, 275.25, 275.35, 
    275.05, 275.85, 275.05, 274.85, 275.25, 275.05, 274.35, 273.95, 274.15, 
    273.65, 273.85, 273.95, 274.15, 274.35, 274.55, 274.35, 273.95, 273.85, 
    273.95, 273.85, 274.15, 273.85, 274.35, 274.95, 274.65, 275.05, 274.45, 
    273.55, 273.75, 273.85, 273.15, 272.55, 272.85, 272.75, 272.85, 272.85, 
    272.85, 272.95, 273.25, 273.55, 273.65, 273.75, 274.15, 273.35, 273.25, 
    273.45, 272.75, 272.55, 272.75, 272.75, 272.45, 272.25, 271.95, 271.85, 
    271.55, 271.55, 271.25, 271.15, 271.05, 270.95, 271.05, 270.75, 270.85, 
    270.75, 271.15, 271.15, 271.25, 271.45, 270.95, 270.75, 270.75, 270.75, 
    270.75, 271.15, 271.35, 271.65, 271.25, 271.35, 271.35, 271.25, 271.35, 
    271.35, 270.95, 271.15, 271.35, 271.15, 271.05, 271.35, 271.45, 271.95, 
    272.35, 272.95, 273.25, 273.45, 273.75, 273.65, 273.35, 273.15, 273.55, 
    273.95, 274.45, 273.05, 271.55, 271.75, 270.95, 270.45, 270.85, 271.45, 
    272.15, 271.95, 272.05, 272.35, 272.65, 272.55, 273.65, 275.25, 275.15, 
    275.15, 275.35, 275.15, 275.45, 275.45, 275.15, 275.15, 274.95, 274.75, 
    274.45, 274.45, 274.65, 274.45, 274.55, 274.65, 274.65, 274.75, 274.95, 
    275.35, 275.55, 275.25, 275.55, 275.35, 276.05, 276.15, 275.65, 276.45, 
    276.65, 276.25, 276.65, 275.95, 275.35, 274.85, 274.45, 273.75, 273.45, 
    274.75, 275.45, 275.55, 275.85, 276.05, 275.65, 276.05, 276.35, 276.25, 
    275.85, 276.05, 275.95, 276.05, 276.45, 277.05, 277.25, 276.75, 276.65, 
    276.65, 276.15, 276.15, 276.25, 276.45, 275.95, 275.95, 275.75, 276.15, 
    276.05, 276.15, 276.25, 276.35, 276.85, 277.15, 277.35, 277.55, 277.75, 
    277.85, 277.65, 277.95, 278.25, 276.65, 276.25, 276.35, 276.15, 275.55, 
    275.45, 274.95, 275.05, 275.05, 275.05, 275.05, 275.05, 274.75, 275.05, 
    274.95, 274.95, 275.15, 275.45, 275.45, 275.75, 274.95, 274.55, 274.65, 
    274.65, 274.45, 274.75, 274.55, 274.85, 274.95, 274.35, 274.35, 274.35, 
    274.35, 274.15, 273.95, 274.35, 274.35, 274.65, 275.05, 275.05, 275.15, 
    275.45, 275.75, 275.85, 276.15, 276.05, 276.25, 275.25, 276.05, 276.75, 
    277.35, 277.35, 277.75, 277.35, 276.45, 276.05, 277.15, 277.05, 277.25, 
    277.15, 277.65, 278.35, 278.15, 278.05, 278.95, 279.95, 280.45, 279.85, 
    279.35, 278.35, 278.05, 277.35, 277.35, 275.25, 276.15, 276.05, 276.45, 
    276.65, 276.15, 276.15, 275.65, 274.95, 274.95, 275.45, 275.45, 275.65, 
    276.15, 276.95, 277.35, 277.05, 276.75, 276.85, 277.05, 277.05, 276.85, 
    276.85, 276.95, 277.05, 276.95, 276.25, 276.45, 276.05, 275.35, 274.95, 
    274.75, 274.95, 274.65, 275.35, 275.05, 275.85, 275.55, 275.95, 276.85, 
    277.15, 276.25, 277.35, 277.55, 278.15, 278.25, 278.75, 278.65, 278.75, 
    278.15, 277.95, 276.95, 277.25, 277.05, 276.95, 277.45, 277.65, 277.55, 
    277.95, 277.95, 277.15, 277.45, 278.75, 278.55, 279.25, 278.75, 279.05, 
    278.75, 278.85, 277.55, 277.95, 277.25, 278.05, 277.35, 277.05, 277.35, 
    277.55, 277.45, 277.25, 277.05, 276.65, 276.65, 277.15, 276.85, 276.85, 
    277.25, 277.35, 277.25, 277.45, 277.45, 277.45, 277.35, 277.15, 277.05, 
    276.75, 276.75, 276.85, 276.95, 276.95, 276.85, 276.65, 276.75, 276.55, 
    276.45, 276.25, 276.05, 275.85, 275.95, 276.45, 276.65, 276.85, 277.05, 
    276.75, 277.85, 278.55, 278.35, 278.55, 278.85, 278.75, 278.65, 278.45, 
    278.25, 277.95, 277.75, 277.25, 277.05, 277.05, 276.75, 276.45, 276.75, 
    276.35, 276.55, 276.55, 276.55, 276.25, 276.45, 276.55, 276.85, 276.75, 
    277.45, 277.55, 277.05, 276.65, 276.45, 276.15, 276.05, 275.45, 275.25, 
    275.05, 274.65, 274.75, 273.95, 274.05, 273.95, 274.05, 275.05, 274.65, 
    275.45, 275.55, 275.35, 275.25, 275.05, 276.15, 276.05, 276.15, 277.05, 
    276.25, 276.05, 275.65, 274.85, 274.65, 274.35, 273.35, 272.95, 272.65, 
    272.55, 272.25, 272.25, 272.65, 272.75, 272.65, 273.35, 274.05, 273.95, 
    274.35, 274.45, 274.25, 274.05, 274.05, 274.45, 274.35, 274.75, 274.15, 
    274.15, 273.75, 273.35, 272.85, 272.75, 272.65, 272.55, 272.65, 272.95, 
    273.25, 273.75, 273.55, 273.55, 273.65, 273.85, 273.85, 273.95, 274.05, 
    274.25, 274.35, 274.15, 274.25, 274.15, 274.35, 274.15, 274.15, 273.95, 
    273.85, 273.95, 273.75, 274.05, 274.05, 273.95, 273.95, 273.75, 273.65, 
    273.85, 273.75, 273.75, 274.05, 274.55, 274.75, 275.05, 275.05, 274.75, 
    274.85, 274.85, 274.75, 274.85, 274.75, 274.65, 274.55, 274.45, 274.45, 
    274.35, 274.35, 274.35, 274.75, 275.05, 275.15, 275.05, 275.15, 275.15, 
    275.25, 275.55, 275.85, 275.95, 276.35, 276.35, 276.65, 276.65, 276.85, 
    276.75, 276.45, 276.65, 276.35, 276.15, 275.85, 275.05, 275.05, 275.25, 
    275.65, 276.45, 276.45, 276.35, 276.65, 277.15, 276.95, 276.45, 276.75, 
    277.65, 278.35, 278.65, 277.55, 277.45, 277.15, 276.65, 276.55, 276.55, 
    276.75, 276.35, 276.45, 276.25, 276.15, 276.65, 276.85, 276.75, 277.15, 
    277.75, 278.05, 277.95, 278.35, 278.75, 279.25, 279.75, 280.05, 280.35, 
    280.55, 280.55, 280.55, 280.35, 280.25, 279.75, 279.05, 278.75, 278.25, 
    277.35, 277.75, 277.35, 277.35, 277.75, 277.55, 277.65, 277.95, 277.05, 
    278.25, 278.95, 279.45, 279.85, 278.85, 278.25, 277.65, 277.65, 277.35, 
    277.85, 277.95, 277.65, 277.65, 277.75, 277.25, 276.65, 276.45, 276.35, 
    276.15, 277.75, 276.55, 276.85, 276.95, 277.25, 277.35, 277.25, 277.05, 
    277.45, 276.95, 276.95, 276.55, 276.55, 276.55, 276.35, 275.95, 276.45, 
    275.85, 275.85, 275.85, 275.35, 275.45, 275.55, 275.55, 275.95, 275.95, 
    275.95, 276.25, 276.55, 276.35, 276.55, 277.05, 276.55, 276.55, 276.65, 
    277.05, 277.05, 277.15, 277.05, 277.05, 277.15, 276.85, 276.75, 276.95, 
    277.05, 277.15, 277.05, 277.15, 277.15, 277.35, 277.85, 277.75, 277.95, 
    278.35, 278.05, 278.25, 278.55, 279.25, 279.15, 278.75, 278.45, 278.35, 
    278.95, 279.25, 279.15, 279.25, 278.75, 278.45, 278.35, 278.25, 278.05, 
    278.35, 278.45, 278.55, 278.75, 278.75, 278.85, 279.35, 279.75, 280.05, 
    280.35, 280.65, 280.55, 280.55, 280.85, 280.05, 280.35, 280.35, 280.55, 
    279.25, 279.85, 279.65, 279.15, 278.55, 279.65, 279.65, 279.25, 279.25, 
    278.25, 278.25, 279.95, 280.15, 278.65, 279.35, 279.85, 280.55, 280.55, 
    280.25, 279.95, 279.55, 279.85, 279.25, 279.15, 278.95, 278.95, 279.35, 
    279.15, 278.65, 278.75, 279.05, 279.55, 278.95, 279.65, 279.45, 279.25, 
    278.95, 279.35, 278.75, 279.85, 279.45, 279.25, 279.25, 279.65, 279.05, 
    278.95, 278.85, 279.05, 279.05, 278.85, 278.85, 278.85, 279.05, 278.65, 
    278.75, 278.75, 278.55, 279.05, 278.35, 279.25, 279.25, 278.75, 279.45, 
    279.95, 279.25, 279.05, 278.95, 278.55, 278.55, 278.65, 278.85, 276.75, 
    277.15, 277.25, 277.35, 277.45, 277.65, 277.75, 277.75, 278.05, 277.75, 
    278.35, 278.85, 278.55, 277.95, 277.95, 278.45, 278.65, 278.45, 278.65, 
    278.45, 278.75, 278.75, 279.25, 279.15, 278.85, 277.85, 277.65, 277.35, 
    277.15, 277.15, 277.55, 277.65, 277.85, 277.95, 278.25, 278.65, 279.25, 
    279.45, 279.55, 279.85, 279.65, 279.65, 279.95, 279.65, 279.65, 279.65, 
    279.65, 279.15, 278.95, 278.45, 278.15, 277.95, 277.95, 277.85, 277.75, 
    277.35, 277.45, 277.95, 277.45, 277.95, 278.05, 278.05, 278.65, 278.75, 
    278.85, 279.15, 279.05, 279.15, 278.65, 279.05, 278.65, 278.35, 278.35, 
    278.05, 278.05, 277.85, 277.85, 277.85, 278.15, 278.35, 278.55, 278.55, 
    278.25, 278.65, 278.75, 278.75, 279.05, 279.25, 279.55, 279.55, 279.65, 
    279.65, 279.55, 279.35, 279.35, 279.45, 278.85, 278.75, 278.85, 278.75, 
    278.45, 278.35, 278.55, 278.65, 278.85, 278.85, 278.75, 278.95, 279.45, 
    279.75, 279.85, 279.75, 280.65, 281.05, 281.25, 280.55, 280.15, 280.25, 
    279.75, 279.85, 279.55, 279.35, 279.45, 279.25, 279.65, 279.65, 279.05, 
    278.75, 278.05, 278.05, 278.45, 278.35, 278.55, 278.05, 278.05, 278.25, 
    278.05, 278.05, 277.75, 278.75, 278.25, 277.65, 277.45, 277.35, 277.55, 
    277.85, 278.05, 278.05, 277.85, 278.15, 278.45, 278.75, 278.35, 278.85, 
    278.65, 279.65, 279.65, 279.75, 279.65, 279.45, 279.65, 280.45, 280.75, 
    280.05, 280.15, 280.15, 279.85, 279.65, 279.45, 279.45, 279.55, 278.95, 
    279.05, 278.85, 279.45, 279.95, 279.55, 279.35, 279.95, 280.45, 279.65, 
    280.15, 280.25, 280.45, 280.25, 279.95, 279.85, 280.15, 280.15, 280.65, 
    280.45, 280.75, 280.75, 280.55, 280.85, 280.75, 279.85, 279.95, 280.25, 
    280.45, 280.55, 280.55, 280.55, 280.05, 280.15, 280.65, 280.65, 280.45, 
    280.85, 280.95, 281.35, 281.25, 281.05, 280.85, 280.45, 280.75, 280.75, 
    280.65, 279.95, 279.65, 279.85, 279.45, 279.25, 279.35, 279.35, 279.45, 
    279.65, 279.35, 280.25, 280.45, 279.85, 280.05, 280.85, 280.45, 280.65, 
    280.65, 280.45, 280.35, 280.05, 280.85, 280.05, 280.05, 280.05, 279.85, 
    279.25, 278.85, 279.65, 280.55, 281.25, 280.35, 280.85, 282.35, 282.05, 
    282.45, 282.95, 283.05, 283.45, 283.95, 284.65, 284.85, 284.25, 283.75, 
    283.85, 283.35, 283.15, 283.35, 282.75, 282.45, 282.25, 282.15, 281.65, 
    281.55, 281.55, 281.45, 281.25, 280.85, 281.45, 280.95, 281.05, 281.85, 
    282.15, 282.85, 282.75, 282.15, 282.35, 282.05, 282.05, 282.35, 281.25, 
    281.35, 281.75, 281.45, 281.25, 281.25, 281.05, 280.15, 279.95, 280.35, 
    280.65, 280.75, 280.65, 280.65, 280.85, 281.35, 281.65, 281.65, 281.55, 
    281.75, 281.65, 281.65, 281.25, 281.15, 281.45, 281.25, 281.35, 281.35, 
    281.15, 280.95, 281.35, 281.15, 281.55, 281.75, 282.35, 283.05, 283.35, 
    283.45, 283.35, 283.25, 283.45, 283.45, 283.85, 284.25, 284.25, 284.25, 
    284.35, 284.05, 283.95, 282.75, 282.25, 281.85, 281.15, 281.15, 281.65, 
    283.65, 283.45, 283.15, 283.75, 284.15, 285.25, 285.95, 286.45, 286.95, 
    287.75, 288.15, 288.45, 288.45, 288.55, 288.45, 287.75, 286.15, 285.65, 
    284.25, 283.95, 283.55, 282.85, 282.45, 282.55, 285.25, 285.65, 284.25, 
    284.75, 286.15, 287.45, 289.25, 289.35, 288.65, 288.35, 287.75, 287.55, 
    286.55, 286.95, 286.65, 285.75, 285.95, 286.15, 284.25, 284.45, 283.75, 
    282.65, 283.35, 282.35, 281.15, 280.85, 281.05, 281.25, 280.65, 279.65, 
    279.35, 279.25, 278.75, 279.35, 279.65, 279.55, 279.35, 278.85, 279.35, 
    279.55, 279.75, 279.55, 279.35, 278.55, 277.75, 278.05, 278.45, 278.75, 
    278.95, 278.95, 278.95, 280.25, 279.75, 279.65, 280.05, 280.15, 279.65, 
    280.55, 280.95, 280.75, 280.85, 281.45, 281.55, 281.95, 282.15, 281.65, 
    280.45, 280.35, 280.05, 279.75, 279.35, 279.45, 281.15, 280.55, 280.85, 
    281.75, 280.85, 280.95, 281.35, 281.65, 282.45, 282.45, 282.45, 282.75, 
    282.85, 283.55, 283.35, 283.85, 282.85, 282.85, 281.95, 281.85, 282.15, 
    281.85, 280.85, 280.85, 280.85, 280.95, 281.65, 282.05, 282.05, 282.75, 
    282.45, 282.15, 281.65, 281.95, 282.05, 282.25, 282.15, 282.65, 283.25, 
    282.55, 283.25, 282.85, 282.15, 282.25, 282.45, 282.65, 282.75, 283.05, 
    283.55, 283.35, 282.75, 282.95, 284.15, 284.15, 284.15, 284.05, 284.75, 
    285.15, 284.25, 284.65, 284.85, 285.25, 284.05, 283.95, 283.65, 283.95, 
    283.35, 283.25, 282.25, 282.25, 282.05, 282.15, 283.35, 283.35, 283.45, 
    283.25, 284.55, 284.15, 284.85, 284.45, 284.35, 284.75, 284.25, 284.45, 
    284.45, 284.45, 284.35, 284.55, 284.45, 283.65, 282.55, 282.25, 281.75, 
    281.35, 281.75, 283.05, 282.55, 283.15, 283.25, 283.35, 284.15, 285.05, 
    284.95, 284.65, 285.15, 285.35, 285.05, 285.95, 286.15, 286.25, 286.15, 
    285.55, 285.15, 285.25, 283.65, 283.05, 282.75, 282.75, 281.95, 281.35, 
    280.55, 280.35, 280.75, 280.55, 281.15, 282.05, 282.15, 283.75, 283.75, 
    283.95, 284.65, 285.85, 284.75, 284.85, 284.55, 284.85, 283.25, 283.05, 
    282.35, 283.45, 283.45, 282.85, 284.35, 283.95, 283.45, 283.85, 285.05, 
    284.05, 284.35, 283.95, 284.15, 284.05, 285.25, 283.85, 283.55, 283.45, 
    282.55, 282.85, 282.75, 282.05, 282.35, 281.95, 281.65, 282.65, 281.65, 
    282.05, 281.85, 281.75, 281.65, 281.95, 280.95, 280.95, 281.15, 281.05, 
    281.05, 280.65, 281.25, 281.85, 281.45, 282.05, 281.15, 282.05, 282.05, 
    282.75, 282.75, 282.25, 281.55, 281.75, 282.05, 282.15, 281.55, 282.95, 
    283.45, 284.15, 282.45, 283.65, 284.85, 285.05, 286.15, 287.05, 287.35, 
    288.25, 288.75, 288.75, 288.45, 288.55, 287.85, 286.35, 284.65, 284.45, 
    284.55, 283.25, 283.35, 283.35, 283.85, 283.75, 284.35, 283.45, 283.25, 
    284.35, 283.45, 284.35, 285.95, 284.45, 284.65, 284.65, 283.45, 284.45, 
    285.45, 284.45, 283.85, 283.75, 283.35, 282.85, 283.05, 282.95, 283.35, 
    282.95, 282.95, 283.15, 282.95, 282.85, 283.05, 282.65, 283.15, 282.35, 
    282.05, 283.05, 282.85, 282.95, 283.05, 282.55, 282.55, 282.05, 282.15, 
    282.25, 282.15, 281.45, 281.25, 280.65, 280.55, 280.55, 280.55, 280.75, 
    280.75, 280.95, 280.75, 280.95, 281.15, 281.55, 282.15, 282.15, 282.45, 
    283.15, 282.85, 283.25, 283.25, 283.25, 283.75, 283.35, 284.55, 284.35, 
    284.15, 283.55, 283.35, 283.55, 284.25, 283.95, 284.15, 284.15, 283.55, 
    284.35, 283.75, 283.95, 284.05, 284.05, 283.25, 283.65, 284.25, 283.95, 
    284.75, 285.45, 285.55, 285.75, 285.95, 285.35, 286.15, 285.95, 285.15, 
    284.25, 284.55, 283.55, 284.35, 285.25, 285.85, 285.65, 285.65, 285.75, 
    284.85, 284.15, 282.95, 282.35, 282.85, 283.05, 282.85, 282.55, 283.05, 
    282.65, 282.25, 282.15, 281.95, 282.05, 281.35, 281.25, 281.15, 281.35, 
    281.65, 281.15, 281.05, 281.05, 281.35, 281.45, 281.65, 281.15, 280.75, 
    280.45, 280.05, 280.35, 280.85, 280.85, 280.85, 281.35, 281.35, 281.35, 
    281.15, 281.35, 281.05, 281.55, 281.35, 280.85, 280.45, 280.55, 280.85, 
    281.25, 281.55, 282.25, 282.55, 283.05, 282.85, 283.25, 282.55, 281.95, 
    282.55, 282.25, 282.65, 282.55, 282.65, 282.35, 282.25, 281.95, 281.65, 
    281.25, 280.85, 280.55, 280.45, 280.25, 279.95, 280.45, 280.35, 280.45, 
    280.85, 281.05, 281.25, 281.45, 281.55, 281.65, 281.85, 281.85, 281.85, 
    281.85, 280.95, 280.85, 280.85, 280.85, 280.95, 280.45, 280.25, 279.65, 
    279.55, 280.35, 280.05, 280.25, 281.15, 281.35, 280.95, 281.35, 281.25, 
    281.65, 281.75, 281.95, 281.85, 282.05, 281.95, 281.95, 282.35, 281.95, 
    281.65, 281.55, 281.45, 280.15, 279.95, 279.85, 279.85, 279.45, 280.05, 
    279.75, 280.05, 280.25, 280.75, 280.35, 280.75, 281.25, 281.15, 281.45, 
    281.45, 281.45, 281.75, 281.75, 281.65, 281.55, 280.65, 281.15, 281.45, 
    281.55, 281.45, 279.95, 281.55, 281.25, 281.75, 282.55, 282.05, 281.75, 
    283.05, 282.25, 282.75, 282.45, 282.95, 283.15, 283.55, 282.35, 281.35, 
    282.15, 282.05, 281.75, 281.75, 281.75, 281.55, 281.25, 281.15, 281.35, 
    281.15, 281.25, 281.55, 281.35, 282.05, 282.45, 281.55, 281.65, 282.35, 
    282.65, 283.15, 282.95, 283.15, 283.05, 283.15, 282.55, 282.55, 281.95, 
    281.25, 281.25, 280.35, 280.45, 280.25, 280.75, 280.95, 281.35, 281.35, 
    281.45, 282.15, 281.85, 282.35, 282.25, 282.35, 282.65, 282.15, 282.65, 
    282.45, 282.75, 282.65, 282.75, 283.15, 282.65, 282.05, 281.35, 280.95, 
    280.75, 280.05, 280.25, 279.65, 279.85, 281.35, 281.45, 281.65, 281.35, 
    281.45, 281.55, 281.55, 281.55, 281.25, 281.75, 281.85, 281.85, 281.65, 
    281.35, 280.85, 280.45, 280.45, 279.95, 279.95, 280.05, 280.05, 279.85, 
    279.75, 279.55, 279.45, 279.25, 279.15, 279.45, 279.65, 280.45, 280.55, 
    280.25, 281.05, 280.15, 279.55, 279.45, 279.35, 279.25, 279.65, 279.45, 
    279.35, 279.25, 278.65, 278.45, 278.25, 278.15, 278.35, 278.75, 278.35, 
    279.05, 278.65, 279.05, 279.75, 280.95, 280.75, 280.45, 280.45, 280.75, 
    281.45, 280.35, 280.65, 280.85, 281.45, 281.35, 281.65, 280.65, 279.65, 
    279.85, 279.15, 278.55, 278.35, 278.55, 278.65, 278.95, 279.35, 279.55, 
    280.25, 280.05, 280.15, 280.35, 280.45, 280.05, 280.45, 280.25, 279.45, 
    280.25, 280.55, 280.45, 280.65, 280.05, 279.35, 279.15, 278.75, 279.85, 
    279.25, 279.65, 280.05, 280.15, 281.05, 280.85, 280.85, 281.55, 281.45, 
    282.85, 282.15, 282.35, 282.45, 282.25, 282.25, 282.15, 281.75, 281.55, 
    281.25, 281.05, 281.25, 281.15, 281.25, 281.15, 281.45, 281.55, 282.05, 
    283.35, 282.55, 282.15, 283.45, 284.05, 284.95, 283.95, 284.45, 284.55, 
    284.85, 286.25, 286.65, 285.95, 284.95, 282.15, 281.25, 280.75, 280.75, 
    280.55, 279.95, 279.55, 279.65, 280.15, 279.65, 279.85, 279.95, 280.15, 
    280.65, 280.95, 280.85, 280.45, 280.85, 282.15, 282.45, 281.85, 281.45, 
    280.35, 279.95, 279.85, 279.65, 279.35, 279.25, 279.05, 278.85, 278.95, 
    278.95, 278.85, 279.05, 279.25, 279.65, 279.95, 279.95, 280.75, 281.35, 
    280.95, 281.35, 281.05, 281.25, 281.25, 281.15, 280.85, 280.25, 280.05, 
    279.65, 279.15, 278.75, 278.55, 278.45, 278.35, 278.35, 278.45, 278.55, 
    278.35, 278.65, 278.75, 278.75, 278.75, 278.65, 278.85, 278.95, 278.95, 
    279.25, 279.05, 279.25, 279.15, 279.25, 279.25, 279.05, 278.95, 278.85, 
    278.65, 278.75, 278.55, 278.15, 278.75, 278.45, 278.55, 279.25, 279.25, 
    279.65, 280.05, 279.95, 280.35, 280.15, 280.65, 280.15, 280.35, 280.25, 
    280.15, 279.75, 279.25, 279.25, 279.15, 278.75, 278.45, 278.55, 278.65, 
    278.55, 278.55, 278.45, 278.65, 278.85, 278.95, 278.95, 278.95, 278.95, 
    279.25, 278.85, 279.15, 279.05, 279.15, 279.25, 279.15, 279.45, 279.25, 
    279.15, 278.95, 278.65, 278.35, 278.35, 278.15, 277.95, 277.75, 277.65, 
    278.45, 279.15, 279.35, 279.15, 279.55, 280.05, 279.85, 279.95, 280.15, 
    280.15, 279.75, 280.05, 279.75, 279.95, 279.85, 280.05, 279.45, 278.95, 
    278.65, 278.35, 278.45, 278.65, 278.35, 278.45, 278.55, 279.25, 279.35, 
    279.75, 280.05, 280.95, 280.85, 281.05, 280.85, 281.25, 280.45, 280.25, 
    279.65, 279.65, 278.95, 278.25, 277.65, 277.15, 276.75, 276.65, 276.75, 
    276.85, 276.85, 277.65, 278.25, 279.05, 279.35, 279.45, 278.85, 278.95, 
    279.35, 279.65, 279.25, 279.35, 279.45, 279.35, 278.75, 278.15, 277.75, 
    277.25, 277.15, 277.15, 277.15, 277.25, 277.25, 277.35, 277.55, 278.05, 
    278.45, 278.75, 278.45, 278.35, 278.85, 279.35, 279.35, 279.05, 279.75, 
    279.55, 279.45, 279.05, 278.75, 278.75, 278.75, 278.35, 277.65, 277.65, 
    277.75, 277.65, 277.75, 278.65, 278.05, 277.95, 278.55, 278.95, 278.65, 
    278.65, 278.75, 279.05, 279.15, 279.35, 279.15, 278.85, 279.15, 279.25, 
    278.55, 278.75, 278.55, 278.05, 277.45, 277.45, 277.45, 277.65, 278.05, 
    278.15, 278.35, 278.75, 280.25, 278.95, 279.75, 279.85, 279.85, 280.35, 
    279.55, 279.65, 279.85, 280.35, 280.55, 280.25, 279.75, 279.15, 279.25, 
    279.15, 278.75, 278.35, 277.85, 277.95, 277.95, 278.05, 278.85, 279.45, 
    279.75, 279.45, 280.55, 280.05, 280.25, 280.65, 280.15, 279.75, 279.55, 
    279.35, 279.25, 278.95, 278.85, 279.15, 279.15, 278.75, 278.35, 277.75, 
    277.15, 277.15, 277.15, 277.45, 277.25, 277.55, 278.25, 278.45, 278.55, 
    278.45, 279.25, 279.05, 279.15, 279.25, 279.35, 279.25, 279.15, 279.05, 
    279.05, 278.95, 278.65, 278.65, 278.55, 278.35, 277.95, 277.85, 277.85, 
    277.95, 278.05, 278.25, 278.55, 278.65, 280.15, 279.85, 280.05, 280.85, 
    281.25, 281.55, 281.25, 281.15, 281.35, 280.65, 280.95, 280.55, 280.45, 
    280.15, 280.05, 279.85, 279.25, 278.75, 279.05, 278.65, 279.35, 279.85, 
    280.45, 280.95, 281.65, 280.35, 280.55, 280.85, 280.15, 280.15, 279.85, 
    279.65, 279.75, 280.95, 280.95, 280.85, 280.95, 280.95, 281.15, 281.05, 
    281.15, 280.85, 280.85, 281.75, 281.55, 281.45, 281.05, 280.75, 281.15, 
    281.45, 280.85, 280.25, 280.15, 280.15, 280.25, 279.75, 280.25, 282.05, 
    281.95, 281.75, 281.95, 282.15, 281.85, 282.05, 281.95, 282.15, 282.15, 
    281.85, 281.65, 281.35, 281.65, 281.55, 281.45, 281.95, 281.95, 282.15, 
    281.65, 282.05, 282.05, 281.95, 282.15, 281.95, 281.55, 280.95, 280.95, 
    281.35, 281.25, 281.15, 280.95, 280.85, 281.05, 280.45, 280.15, 279.95, 
    279.85, 280.05, 279.85, 279.95, 280.25, 280.25, 279.95, 280.05, 279.65, 
    279.85, 280.05, 280.85, 280.25, 280.95, 279.75, 279.75, 280.15, 279.75, 
    279.85, 279.45, 279.05, 278.75, 278.75, 278.55, 278.55, 278.75, 278.85, 
    279.05, 279.55, 280.35, 280.75, 281.15, 281.15, 281.85, 281.65, 281.25, 
    279.85, 279.25, 278.35, 278.05, 278.05, 277.85, 277.85, 277.85, 277.65, 
    277.75, 278.25, 278.25, 278.15, 278.35, 278.75, 277.95, 279.05, 279.35, 
    279.65, 279.85, 280.25, 280.75, 280.85, 279.65, 279.65, 279.15, 278.65, 
    277.85, 277.75, 277.55, 276.65, 276.75, 276.75, 276.65, 276.35, 277.15, 
    277.75, 277.05, 276.65, 276.45, 276.65, 276.55, 277.45, 278.05, 277.55, 
    277.35, 277.65, 277.05, 276.25, 275.95, 275.15, 274.75, 274.95, 274.65, 
    274.25, 273.85, 273.65, 274.45, 275.75, 276.25, 276.25, 276.15, 276.05, 
    276.65, 276.75, 276.95, 277.65, 277.35, 277.55, 277.95, 277.75, 277.65, 
    277.65, 277.45, 276.85, 276.35, 276.45, 276.35, 276.35, 276.35, 277.55, 
    277.65, 277.85, 277.65, 277.75, 277.85, 277.55, 277.95, 278.15, 277.85, 
    277.75, 275.95, 275.75, 275.25, 274.85, 274.85, 274.45, 274.15, 274.05, 
    273.95, 273.15, 273.45, 273.25, 273.35, 273.45, 273.75, 273.85, 274.55, 
    275.05, 274.65, 274.95, 275.05, 275.45, 275.85, 275.45, 274.95, 275.45, 
    275.55, 275.25, 275.25, 274.65, 274.65, 274.25, 274.05, 274.25, 274.15, 
    273.95, 273.65, 274.15, 274.25, 274.75, 275.15, 275.85, 276.25, 277.05, 
    277.55, 277.15, 277.15, 277.25, 277.65, 277.35, 277.05, 276.95, 276.85, 
    276.65, 276.25, 275.85, 275.45, 276.55, 277.65, 277.35, 277.15, 276.65, 
    276.55, 276.75, 276.35, 276.85, 276.85, 277.55, 278.15, 278.25, 278.45, 
    278.35, 278.25, 278.25, 278.45, 278.45, 278.55, 278.55, 277.55, 277.15, 
    277.15, 277.05, 277.05, 276.55, 276.45, 276.65, 276.35, 275.75, 276.35, 
    276.65, 277.05, 277.45, 276.45, 277.45, 277.75, 277.55, 277.55, 277.55, 
    276.95, 276.45, 276.65, 276.75, 276.95, 276.45, 276.35, 276.05, 275.85, 
    275.85, 275.65, 275.25, 274.95, 275.15, 274.65, 274.75, 275.65, 275.75, 
    275.35, 275.45, 275.25, 275.35, 275.65, 276.05, 276.05, 276.15, 275.95, 
    275.85, 275.75, 275.55, 275.85, 275.75, 275.45, 275.05, 275.35, 275.35, 
    275.55, 275.55, 275.85, 275.85, 275.25, 275.45, 275.65, 276.05, 276.55, 
    276.55, 276.65, 276.65, 276.55, 276.35, 277.15, 276.65, 276.25, 275.85, 
    275.45, 275.25, 274.85, 273.95, 273.35, 273.35, 273.15, 273.45, 274.55, 
    275.65, 276.05, 276.75, 276.65, 276.85, 277.05, 277.15, 276.85, 276.95, 
    276.65, 276.15, 275.85, 275.85, 275.55, 275.15, 274.85, 274.55, 273.75, 
    273.35, 274.05, 274.05, 274.05, 274.35, 274.65, 274.65, 275.45, 275.85, 
    275.85, 276.75, 276.65, 276.25, 276.55, 276.35, 276.05, 275.55, 275.55, 
    275.35, 274.85, 274.55, 274.55, 274.65, 273.95, 273.65, 273.85, 274.55, 
    274.35, 274.65, 275.05, 275.65, 275.85, 276.35, 276.65, 276.85, 276.75, 
    277.15, 277.35, 277.55, 276.95, 277.05, 276.85, 276.85, 277.15, 277.15, 
    276.25, 276.55, 276.35, 276.45, 276.25, 275.95, 276.25, 275.95, 276.85, 
    277.55, 278.15, 278.45, 278.05, 278.55, 278.75, 278.25, 278.35, 277.85, 
    278.05, 277.65, 276.75, 276.25, 275.45, 275.45, 276.15, 275.05, 273.65, 
    274.45, 274.35, 273.75, 273.85, 274.05, 276.05, 276.15, 276.95, 277.25, 
    277.45, 277.55, 277.25, 277.15, 277.15, 277.35, 277.15, 277.35, 277.25, 
    276.75, 276.35, 276.25, 276.55, 275.85, 276.45, 275.75, 276.15, 276.25, 
    275.75, 276.05, 276.15, 276.45, 276.85, 277.25, 277.75, 277.75, 277.55, 
    277.95, 278.05, 277.65, 277.85, 277.35, 277.25, 276.55, 276.05, 276.55, 
    276.05, 276.05, 276.25, 275.45, 275.45, 275.75, 275.65, 276.15, 276.65, 
    276.65, 276.75, 277.25, 277.35, 277.15, 277.45, 277.25, 277.25, 277.15, 
    277.15, 277.35, 277.25, 277.15, 276.95, 276.75, 276.55, 276.55, 276.35, 
    276.25, 276.15, 276.25, 276.45, 276.35, 276.65, 276.95, 277.35, 278.55, 
    277.85, 277.85, 278.05, 278.05, 278.05, 277.85, 277.95, 277.75, 277.65, 
    277.45, 277.15, 277.15, 276.65, 276.85, 276.95, 276.75, 276.35, 276.35, 
    276.45, 276.45, 276.35, 277.65, 277.85, 277.75, 277.55, 277.55, 277.25, 
    277.15, 277.65, 277.35, 276.65, 276.95, 276.15, 276.35, 275.85, 275.45, 
    275.65, 274.75, 274.25, 273.55, 273.15, 273.65, 273.65, 273.75, 275.05, 
    275.15, 275.75, 276.15, 276.25, 276.45, 276.45, 276.45, 276.75, 277.05, 
    276.45, 275.55, 275.05, 274.65, 273.95, 273.85, 272.95, 272.95, 273.25, 
    273.15, 273.25, 272.65, 272.75, 274.05, 274.05, 276.05, 275.35, 275.75, 
    276.35, 276.75, 277.65, 276.85, 276.25, 275.45, 275.25, 275.05, 275.15, 
    274.55, 274.35, 274.85, 274.85, 274.55, 274.05, 274.45, 274.85, 274.05, 
    274.25, 274.35, 276.35, 276.25, 277.15, 277.55, 277.45, 277.85, 277.45, 
    277.65, 277.75, 277.55, 277.35, 276.95, 275.05, 275.85, 274.65, 275.05, 
    274.85, 274.65, 274.95, 275.75, 275.15, 274.45, 274.35, 273.35, 274.55, 
    275.35, 275.65, 275.45, 276.65, 276.15, 276.05, 276.35, 276.25, 275.35, 
    276.05, 276.25, 275.95, 278.05, 278.05, 280.15, 278.95, 278.35, 277.85, 
    277.65, 276.95, 277.35, 277.25, 277.45, 278.25, 278.15, 278.85, 280.25, 
    281.15, 279.25, 280.65, 279.85, 279.65, 280.35, 279.95, 279.65, 279.45, 
    279.05, 279.35, 279.45, 279.65, 279.15, 278.75, 278.35, 278.45, 278.25, 
    277.25, 277.45, 277.55, 277.85, 277.95, 278.25, 278.55, 278.45, 279.75, 
    278.55, 279.75, 278.85, 279.05, 278.05, 277.65, 277.25, 277.15, 276.85, 
    276.85, 276.75, 275.95, 276.05, 275.95, 275.35, 275.55, 276.45, 275.95, 
    276.05, 276.75, 276.45, 276.45, 277.05, 277.15, 277.55, 277.45, 277.35, 
    277.25, 277.15, 276.85, 276.55, 276.05, 276.25, 276.45, 276.75, 277.05, 
    277.25, 277.45, 276.75, 276.35, 276.55, 276.85, 278.45, 279.25, 280.05, 
    280.65, 278.35, 280.25, 280.95, 280.45, 281.05, 281.95, 281.55, 281.75, 
    281.25, 281.35, 282.25, 281.85, 281.65, 281.25, 280.75, 280.25, 280.05, 
    278.95, 279.55, 279.35, 279.55, 279.95, 279.35, 279.35, 280.25, 282.65, 
    282.75, 281.45, 283.75, 283.35, 282.75, 282.75, 282.25, 282.25, 281.05, 
    280.25, 279.75, 279.05, 278.75, 278.65, 278.25, 278.15, 277.75, 277.25, 
    277.15, 277.05, 277.15, 277.05, 277.45, 277.55, 277.15, 277.15, 277.25, 
    277.25, 277.15, 276.95, 276.95, 277.05, 277.05, 276.65, 275.45, 275.65, 
    275.45, 275.75, 275.45, 275.65, 275.55, 275.85, 275.85, 276.05, 276.25, 
    276.15, 276.15, 276.35, 276.05, 275.85, 275.75, 275.35, 275.15, 275.15, 
    275.25, 275.45, 275.45, 275.45, 275.65, 276.25, 276.65, 276.65, 277.55, 
    278.25, 278.95, 277.95, 278.05, 280.15, 279.75, 279.65, 279.55, 279.85, 
    279.45, 278.95, 278.95, 278.85, 278.35, 278.45, 278.15, 278.15, 278.25, 
    277.85, 277.55, 277.95, 277.45, 277.35, 276.95, 276.75, 276.85, 276.55, 
    277.05, 276.85, 277.15, 278.25, 278.65, 278.35, 277.85, 277.35, 276.55, 
    275.25, 275.05, 274.65, 274.95, 274.65, 274.65, 274.65, 274.45, 274.35, 
    274.15, 273.85, 273.35, 273.45, 273.95, 274.05, 274.45, 274.55, 275.05, 
    275.85, 275.45, 274.85, 274.95, 275.15, 274.75, 274.85, 274.75, 274.95, 
    275.05, 275.25, 275.25, 275.55, 276.25, 276.95, 277.35, 277.45, 276.95, 
    276.65, 276.45, 276.85, 276.55, 276.65, 276.75, 276.75, 276.85, 276.95, 
    276.95, 276.95, 277.25, 277.15, 276.85, 276.95, 276.95, 276.85, 276.95, 
    277.05, 276.75, 276.55, 276.85, 276.75, 276.95, 276.75, 276.65, 277.05, 
    276.85, 277.15, 276.95, 277.55, 277.25, 277.35, 277.45, 277.35, 277.25, 
    277.45, 277.35, 277.15, 277.55, 276.95, 276.85, 276.35, 275.25, 275.65, 
    276.35, 275.45, 274.85, 274.75, 274.45, 274.55, 273.65, 273.95, 274.55, 
    274.75, 275.45, 276.25, 276.35, 276.55, 276.25, 276.85, 278.25, 279.65, 
    280.15, 280.05, 279.95, 280.25, 279.65, 278.95, 278.95, 278.85, 279.35, 
    279.45, 279.25, 279.55, 279.05, 278.45, 278.65, 278.45, 278.75, 279.25, 
    278.75, 278.15, 278.45, 279.15, 279.15, 279.85, 279.35, 278.75, 278.25, 
    278.25, 278.15, 278.05, 278.25, 277.95, 277.45, 278.05, 277.85, 277.95, 
    277.75, 278.05, 277.95, 278.25, 277.35, 278.15, 278.75, 277.95, 278.35, 
    278.15, 277.65, 277.25, 277.35, 276.35, 275.25, 275.55, 275.05, 275.45, 
    275.45, 276.25, 277.85, 277.85, 278.55, 277.75, 278.85, 277.65, 277.85, 
    278.05, 277.95, 277.85, 277.75, 277.95, 277.95, 277.75, 277.55, 277.15, 
    277.15, 276.95, 276.95, 276.85, 276.65, 276.45, 276.25, 276.05, 276.05, 
    275.65, 275.15, 275.35, 275.25, 275.95, 275.75, 275.95, 275.85, 275.95, 
    275.25, 275.25, 275.85, 275.85, 275.55, 275.65, 275.65, 275.85, 276.05, 
    275.75, 275.65, 275.45, 275.15, 275.25, 275.05, 275.65, 275.85, 275.65, 
    275.85, 276.35, 276.75, 276.95, 277.25, 278.05, 278.25, 277.35, 277.25, 
    277.95, 277.45, 276.95, 276.75, 276.55, 276.65, 277.15, 276.45, 276.35, 
    276.35, 276.35, 276.45, 276.45, 276.05, 275.65, 275.65, 275.75, 276.15, 
    276.45, 276.55, 276.55, 276.65, 276.65, 276.35, 275.95, 275.45, 275.45, 
    275.55, 275.45, 275.25, 275.05, 274.75, 274.25, 273.95, 273.75, 273.55, 
    273.05, 272.95, 272.45, 272.35, 272.15, 272.15, 271.95, 272.15, 272.15, 
    272.25, 270.85, 271.45, 271.45, 270.95, 271.05, 271.15, 271.25, 270.75, 
    270.45, 269.95, 269.65, 269.45, 269.75, 270.55, 269.85, 270.35, 270.65, 
    270.75, 270.75, 270.95, 271.05, 271.15, 271.45, 272.05, 272.65, 272.55, 
    272.75, 273.95, 275.65, 276.35, 278.05, 278.25, 277.75, 277.65, 277.45, 
    276.85, 276.25, 276.75, 276.75, 276.75, 277.95, 276.65, 276.75, 277.15, 
    277.85, 277.95, 277.95, 277.85, 277.85, 277.55, 277.25, 277.55, 277.75, 
    277.25, 276.75, 275.65, 276.75, 276.05, 275.85, 275.65, 275.85, 275.75, 
    275.35, 275.05, 274.35, 273.85, 273.25, 273.95, 274.55, 274.75, 274.45, 
    274.55, 274.25, 274.65, 274.25, 274.05, 273.55, 273.55, 273.55, 273.15, 
    274.05, 274.35, 274.75, 274.45, 274.75, 279.05, 279.35, 280.25, 280.55, 
    280.15, 280.05, 279.75, 279.65, 279.35, 279.25, 278.95, 278.55, 277.85, 
    277.45, 277.55, 277.55, 278.35, 277.45, 276.35, 276.55, 275.75, 274.95, 
    274.75, 274.65, 274.35, 273.95, 273.65, 274.05, 273.95, 273.15, 272.95, 
    273.95, 273.25, 273.35, 273.95, 273.95, 274.15, 274.25, 274.35, 273.95, 
    274.35, 274.45, 273.35, 273.95, 275.25, 275.55, 274.65, 275.45, 275.45, 
    276.05, 275.85, 276.05, 276.15, 275.75, 274.75, 274.35, 276.35, 276.55, 
    276.65, 276.05, 276.05, 277.35, 277.35, 277.55, 277.55, 277.95, 278.55, 
    278.45, 278.25, 278.05, 278.35, 279.35, 278.95, 278.55, 279.55, 279.35, 
    279.75, 279.65, 279.05, 279.15, 279.25, 279.15, 279.35, 279.45, 279.55, 
    279.65, 279.35, 279.15, 279.15, 278.85, 278.65, 278.45, 278.55, 278.55, 
    278.75, 278.95, 278.95, 278.85, 278.85, 278.65, 278.45, 277.85, 277.55, 
    277.25, 277.15, 277.55, 277.75, 276.95, 276.85, 277.15, 276.65, 276.25, 
    276.45, 276.55, 276.15, 275.95, 276.05, 275.75, 275.75, 275.95, 276.15, 
    276.05, 275.95, 276.45, 276.95, 276.75, 276.55, 276.25, 276.05, 275.95, 
    275.85, 275.85, 275.95, 275.35, 275.45, 274.65, 274.75, 274.65, 274.75, 
    274.55, 274.45, 274.25, 274.25, 273.75, 273.85, 273.85, 273.85, 273.55, 
    273.35, 273.35, 273.25, 273.35, 273.35, 273.35, 273.05, 273.35, 273.45, 
    273.25, 272.75, 272.95, 273.15, 273.65, 273.15, 272.55, 272.75, 272.85, 
    273.05, 273.15, 273.15, 273.35, 273.35, 273.45, 273.55, 273.95, 273.85, 
    273.65, 273.65, 273.95, 278.05, 278.45, 278.45, 279.55, 279.45, 279.45, 
    279.45, 278.35, 278.65, 278.65, 278.45, 277.65, 277.45, 277.35, 277.65, 
    278.25, 277.85, 277.75, 276.85, 275.65, 274.65, 274.15, 273.35, 272.35, 
    271.25, 269.65, 269.55, 269.55, 269.65, 269.55, 269.75, 270.05, 270.15, 
    270.45, 270.85, 271.05, 270.75, 270.55, 270.35, 270.15, 269.95, 269.55, 
    269.45, 269.15, 269.45, 269.35, 269.55, 269.95, 269.85, 270.35, 270.45, 
    270.75, 271.05, 271.45, 270.95, 271.05, 271.05, 271.45, 271.45, 271.15, 
    271.35, 271.55, 271.95, 272.15, 272.15, 272.05, 272.05, 272.55, 272.95, 
    272.95, 273.15, 272.95, 273.05, 272.65, 273.65, 273.85, 273.45, 273.45, 
    273.75, 275.05, 274.95, 274.95, 274.65, 275.45, 275.65, 275.85, 275.15, 
    275.05, 274.65, 274.55, 274.75, 274.45, 274.75, 274.65, 274.75, 275.05, 
    275.25, 275.05, 275.05, 275.05, 274.95, 274.55, 274.85, 274.85, 275.85, 
    277.15, 277.35, 277.65, 277.85, 276.35, 277.25, 276.35, 276.65, 276.65, 
    276.95, 276.05, 276.25, 276.45, 275.55, 276.05, 275.65, 276.35, 275.75, 
    275.65, 275.65, 275.55, 275.55, 274.85, 275.15, 275.85, 276.25, 276.75, 
    278.15, 278.35, 278.15, 278.45, 278.75, 278.75, 279.15, 278.95, 278.75, 
    278.85, 278.65, 278.75, 278.65, 279.15, 279.45, 279.75, 279.45, 279.55, 
    279.45, 279.95, 280.05, 280.75, 281.05, 280.85, 280.75, 280.75, 280.65, 
    280.45, 280.65, 280.45, 280.15, 280.25, 279.85, 279.85, 280.25, 280.15, 
    279.85, 279.65, 279.45, 279.35, 279.15, 279.15, 278.95, 278.75, 278.25, 
    278.15, 278.25, 278.25, 278.45, 278.45, 278.75, 278.85, 279.65, 279.05, 
    279.05, 279.05, 277.65, 276.75, 275.85, 275.55, 275.45, 275.15, 274.65, 
    274.75, 274.25, 274.25, 274.35, 274.55, 274.25, 274.65, 274.05, 274.35, 
    273.95, 274.25, 274.35, 274.65, 275.15, 275.05, 275.05, 277.75, 278.65, 
    278.55, 278.85, 278.85, 279.05, 279.15, 279.05, 279.35, 279.05, 278.95, 
    278.45, 278.05, 278.05, 277.85, 278.25, 277.65, 277.55, 277.45, 277.75, 
    276.45, 276.75, 276.05, 275.95, 275.75, 275.75, 275.75, 275.65, 275.65, 
    275.55, 276.35, 276.35, 276.65, 276.55, 275.65, 275.65, 277.05, 275.65, 
    275.55, 274.95, 274.35, 275.35, 275.45, 275.15, 276.45, 276.35, 276.05, 
    276.15, 276.65, 276.65, 276.65, 275.75, 275.75, 275.05, 275.75, 275.05, 
    274.45, 274.25, 274.55, 274.35, 274.35, 274.15, 273.75, 273.85, 274.15, 
    274.65, 274.45, 274.85, 274.25, 274.85, 274.25, 274.05, 274.05, 275.45, 
    274.85, 274.75, 274.95, 274.75, 277.15, 276.75, 276.55, 279.55, 279.15, 
    278.55, 278.55, 277.25, 277.45, 277.65, 278.45, 280.05, 279.45, 278.75, 
    278.75, 278.35, 278.55, 278.95, 278.75, 278.55, 277.75, 277.55, 277.65, 
    277.25, 276.95, 277.05, 276.45, 276.95, 276.75, 276.75, 276.35, 276.25, 
    276.65, 276.25, 276.15, 276.45, 275.95, 275.95, 276.25, 276.55, 276.55, 
    276.85, 276.75, 276.55, 277.15, 277.15, 277.85, 277.95, 277.95, 277.35, 
    277.55, 277.35, 277.45, 277.75, 277.75, 277.05, 276.65, 276.55, 276.15, 
    276.15, 275.35, 275.15, 275.45, 275.65, 275.95, 276.15, 275.75, 275.55, 
    274.75, 274.65, 274.55, 274.25, 273.95, 273.85, 273.85, 273.35, 273.15, 
    272.65, 272.95, 273.25, 273.75, 273.65, 273.65, 273.45, 273.45, 273.45, 
    273.55, 273.55, 273.55, 273.55, 273.65, 273.55, 273.65, 273.55, 273.55, 
    273.45, 273.45, 272.25, 272.55, 272.75, 272.65, 272.65, 272.55, 272.05, 
    271.45, 271.45, 271.75, 271.75, 271.45, 270.95, 271.55, 271.75, 271.85, 
    271.75, 271.95, 271.75, 271.75, 271.55, 271.25, 271.55, 271.75, 271.25, 
    271.85, 271.65, 271.45, 271.45, 271.65, 271.35, 270.95, 270.35, 270.25, 
    270.35, 270.35, 270.65, 270.85, 270.45, 270.35, 270.05, 270.35, 270.35, 
    270.05, 270.25, 270.35, 270.35, 270.65, 270.85, 271.15, 271.15, 271.15, 
    271.05, 270.75, 270.35, 269.95, 269.65, 268.75, 268.95, 269.25, 269.45, 
    268.85, 269.55, 269.05, 269.15, 268.75, 268.15, 268.55, 269.25, 269.15, 
    268.95, 268.95, 269.15, 269.45, 269.95, 269.45, 269.85, 269.25, 269.45, 
    269.15, 269.35, 269.55, 269.55, 269.25, 269.25, 269.15, 269.15, 268.55, 
    269.25, 269.65, 269.85, 270.35, 270.45, 270.55, 270.55, 270.75, 270.85, 
    271.05, 271.25, 271.05, 271.05, 270.95, 270.85, 271.35, 271.15, 270.95, 
    270.25, 271.25, 271.25, 271.35, 270.95, 271.25, 271.35, 271.65, 271.65, 
    271.75, 272.25, 272.25, 272.45, 272.45, 272.25, 272.15, 272.35, 271.95, 
    272.45, 272.65, 272.45, 272.95, 272.95, 272.55, 272.05, 272.05, 271.95, 
    271.25, 271.05, 270.95, 270.85, 270.75, 269.95, 270.25, 269.75, 269.75, 
    269.85, 269.35, 269.35, 269.25, 267.75, 267.95, 268.35, 268.25, 268.65, 
    268.75, 269.05, 269.15, 269.05, 269.25, 269.25, 269.55, 270.15, 269.95, 
    271.15, 273.25, 273.65, 273.75, 273.45, 273.65, 274.15, 274.05, 274.25, 
    274.75, 275.35, 275.65, 275.25, 275.25, 274.85, 275.05, 276.35, 276.45, 
    277.05, 276.95, 276.95, 276.85, 276.35, 276.65, 276.75, 277.25, 277.25, 
    277.05, 275.85, 275.85, 276.35, 276.55, 276.35, 276.45, 277.05, 276.45, 
    276.25, 277.55, 278.05, 278.15, 278.65, 278.95, 278.95, 278.55, 278.05, 
    277.55, 276.35, 275.65, 275.35, 274.75, 274.55, 274.35, 274.25, 273.65, 
    273.55, 272.85, 272.45, 272.45, 271.95, 272.05, 272.25, 272.25, 272.15, 
    272.25, 271.85, 271.75, 271.85, 271.95, 272.05, 272.35, 272.65, 272.85, 
    273.05, 273.45, 274.35, 275.15, 276.75, 277.35, 277.75, 277.45, 277.35, 
    277.75, 277.55, 277.15, 276.95, 276.95, 276.85, 276.85, 277.05, 276.95, 
    276.65, 277.15, 276.45, 276.65, 276.35, 276.15, 276.05, 276.15, 276.05, 
    275.75, 276.35, 275.45, 275.55, 274.65, 274.75, 274.65, 274.85, 274.75, 
    274.65, 273.85, 273.45, 273.25, 273.15, 273.15, 273.95, 273.25, 274.25, 
    273.75, 274.15, 273.25, 274.35, 273.75, 273.85, 273.95, 273.65, 273.45, 
    274.55, 274.25, 274.15, 274.15, 274.65, 275.95, 273.75, 274.25, 274.35, 
    274.75, 274.55, 274.75, 274.45, 274.55, 274.45, 273.25, 273.05, 273.25, 
    273.45, 273.45, 273.55, 273.35, 273.65, 273.15, 273.45, 272.85, 273.45, 
    272.65, 272.65, 272.25, 272.95, 274.25, 274.05, 273.45, 273.65, 273.65, 
    273.55, 273.05, 273.25, 273.45, 271.85, 272.15, 272.05, 271.15, 271.75, 
    271.85, 272.55, 272.85, 272.95, 272.35, 273.45, 272.85, 272.95, 272.95, 
    272.35, 271.95, 271.85, 272.35, 272.85, 272.95, 272.65, 272.55, 272.55, 
    273.05, 273.65, 273.45, 273.35, 275.35, 277.45, 277.75, 278.85, 278.35, 
    278.55, 278.95, 278.65, 278.95, 278.25, 278.05, 278.35, 278.25, 277.45, 
    277.35, 276.75, 275.95, 275.25, 275.45, 275.65, 275.15, 275.85, 275.85, 
    275.95, 275.65, 275.85, 275.65, 275.15, 275.15, 274.55, 275.05, 275.35, 
    274.65, 274.75, 274.65, 274.65, 274.75, 274.75, 274.35, 274.55, 274.25, 
    274.45, 274.75, 277.85, 278.25, 278.15, 277.25, 277.15, 276.95, 277.15, 
    276.85, 277.75, 277.55, 278.45, 278.65, 278.55, 278.55, 278.35, 278.35, 
    277.95, 277.65, 277.95, 276.85, 276.15, 275.45, 274.45, 273.25, 273.55, 
    273.35, 274.05, 274.35, 274.05, 274.05, 274.15, 274.25, 274.15, 275.05, 
    274.75, 275.05, 275.25, 275.55, 275.25, 275.25, 275.45, 274.05, 273.85, 
    274.65, 273.65, 273.05, 273.85, 273.05, 272.75, 272.45, 273.35, 273.55, 
    273.75, 274.15, 274.65, 276.25, 276.25, 276.15, 275.95, 275.35, 275.35, 
    275.15, 274.55, 274.95, 274.65, 274.65, 275.75, 274.95, 274.65, 274.15, 
    273.45, 273.75, 274.15, 273.75, 273.65, 273.75, 274.05, 274.75, 275.45, 
    274.65, 274.25, 274.15, 273.95, 273.75, 273.45, 274.05, 274.35, 274.45, 
    274.85, 275.25, 275.15, 275.25, 275.55, 275.75, 275.75, 275.65, 275.35, 
    275.35, 275.05, 274.85, 275.05, 275.05, 274.65, 274.75, 275.25, 275.05, 
    275.25, 275.45, 275.75, 276.05, 275.55, 274.55, 274.75, 274.45, 274.25, 
    273.65, 274.25, 274.55, 274.05, 274.05, 273.95, 273.55, 273.85, 274.05, 
    273.55, 273.35, 273.35, 272.85, 272.65, 272.45, 272.45, 271.75, 271.45, 
    271.25, 269.35, 269.85, 269.65, 269.95, 269.95, 270.05, 270.25, 270.35, 
    270.55, 270.55, 270.55, 270.95, 270.85, 270.75, 270.75, 270.55, 270.65, 
    270.95, 270.75, 270.65, 270.75, 270.75, 270.75, 270.85, 270.95, 271.25, 
    271.65, 271.55, 271.25, 271.45, 271.35, 271.55, 271.35, 271.25, 271.25, 
    271.35, 271.25, 271.25, 271.25, 271.45, 271.25, 271.35, 271.45, 271.35, 
    271.55, 271.45, 271.45, 270.45, 269.95, 269.95, 270.45, 270.55, 270.75, 
    270.55, 271.05, 271.45, 271.65, 271.75, 271.65, 271.45, 271.45, 271.35, 
    271.25, 271.05, 270.85, 270.05, 269.55, 269.05, 269.05, 268.85, 268.75, 
    268.85, 268.95, 268.65, 268.55, 268.45, 268.35, 268.55, 268.65, 268.65, 
    268.65, 268.45, 268.45, 268.45, 268.45, 268.25, 268.05, 268.45, 268.85, 
    268.65, 269.45, 269.45, 269.25, 268.85, 268.95, 267.85, 267.95, 267.25, 
    266.15, 265.45, 265.35, 265.25, 265.15, 265.35, 265.05, 265.05, 264.85, 
    264.55, 264.85, 265.05, 265.35, 265.65, 265.75, 266.15, 266.15, 266.35, 
    266.15, 265.75, 265.05, 264.55, 264.85, 264.85, 264.65, 264.45, 264.95, 
    265.75, 265.75, 265.75, 266.15, 266.45, 266.55, 265.45, 266.15, 265.95, 
    264.75, 263.75, 264.85, 264.85, 263.95, 263.85, 264.15, 264.15, 265.15, 
    264.35, 262.95, 264.25, 263.65, 263.85, 263.75, 263.45, 263.75, 263.15, 
    264.05, 263.05, 264.15, 263.95, 264.25, 264.45, 264.05, 264.15, 264.85, 
    265.05, 264.65, 265.45, 267.75, 268.15, 269.15, 270.05, 270.65, 270.85, 
    270.65, 270.55, 270.55, 269.95, 269.95, 269.35, 269.75, 269.95, 270.25, 
    270.35, 270.55, 270.25, 270.35, 271.05, 271.25, 270.75, 270.35, 270.45, 
    270.25, 270.05, 270.25, 269.95, 269.75, 269.75, 269.25, 268.95, 269.15, 
    269.45, 269.35, 269.65, 269.75, 269.55, 268.75, 269.05, 268.65, 267.85, 
    268.25, 268.55, 268.75, 269.15, 269.05, 268.55, 268.45, 268.25, 267.45, 
    267.25, 267.15, 267.35, 267.35, 267.35, 267.55, 267.25, 266.65, 266.85, 
    266.65, 266.55, 266.15, 264.45, 265.05, 265.85, 266.25, 266.35, 266.55, 
    265.05, 263.95, 263.15, 263.05, 263.95, 262.75, 263.05, 262.85, 262.35, 
    262.65, 262.85, 263.75, 263.15, 263.45, 264.15, 263.75, 264.25, 264.25, 
    263.95, 263.95, 264.05, 264.05, 264.35, 264.25, 264.05, 264.45, 264.45, 
    264.75, 264.45, 264.75, 264.85, 265.05, 265.15, 265.45, 265.35, 265.25, 
    266.15, 267.25, 268.65, 269.15, 269.05, 269.55, 269.55, 269.55, 269.15, 
    269.85, 268.65, 268.05, 266.85, 264.45, 268.05, 266.55, 268.55, 268.25, 
    268.65, 268.65, 267.25, 266.65, 265.85, 266.25, 265.35, 264.25, 265.85, 
    265.95, 268.85, 269.75, 269.05, 268.85, 268.25, 267.85, 267.95, 267.95, 
    267.95, 268.35, 268.05, 268.15, 268.35, 268.05, 267.75, 267.65, 267.75, 
    267.55, 267.15, 266.75, 266.35, 265.85, 266.15, 264.95, 264.05, 263.95, 
    262.95, 263.85, 263.75, 264.05, 264.35, 263.35, 262.35, 262.15, 261.15, 
    260.25, 259.45, 258.75, 257.75, 257.05, 256.65, 256.65, 256.45, 256.95, 
    255.95, 255.35, 255.45, 255.65, 254.95, 254.35, 253.35, 253.15, 253.65, 
    253.25, 253.75, 254.25, 254.05, 253.85, 255.75, 256.25, 257.05, 257.95, 
    258.35, 258.25, 258.15, 258.15, 258.05, 258.05, 258.05, 257.65, 258.15, 
    258.05, 257.95, 258.05, 257.75, 257.65, 257.65, 257.85, 257.55, 257.15, 
    255.15, 254.45, 254.65, 254.25, 255.15, 255.15, 254.35, 254.65, 254.65, 
    254.55, 255.15, 254.85, 254.75, 254.85, 254.95, 254.75, 254.85, 254.95, 
    254.25, 254.85, 254.65, 254.85, 254.75, 254.75, 253.85, 253.75, 254.45, 
    255.55, 254.85, 255.05, 255.15, 257.35, 257.95, 258.15, 259.15, 260.05, 
    260.85, 262.35, 263.35, 264.25, 263.75, 263.25, 263.15, 262.85, 265.25, 
    264.45, 263.95, 263.15, 263.75, 263.15, 263.55, 262.85, 262.25, 261.95, 
    264.25, 263.95, 263.55, 262.45, 261.55, 263.25, 261.45, 261.95, 261.65, 
    261.05, 259.75, 260.15, 261.05, 261.85, 261.95, 261.45, 260.55, 260.15, 
    260.85, 260.65, 260.15, 260.25, 259.95, 260.65, 259.25, 259.55, 259.05, 
    258.25, 259.15, 259.05, 259.35, 259.35, 259.75, 259.45, 260.15, 260.95, 
    260.85, 261.25, 262.05, 261.15, 261.35, 262.05, 261.75, 261.65, 262.35, 
    261.55, 261.65, 261.65, 261.95, 261.85, 260.85, 262.35, 262.75, 262.15, 
    263.25, 263.75, 263.45, 262.15, 261.35, 261.95, 261.45, 261.85, 261.25, 
    261.55, 259.75, 261.35, 260.85, 260.75, 261.25, 261.05, 259.95, 260.25, 
    259.85, 259.85, 259.85, 259.95, 260.35, 260.35, 260.85, 259.75, 259.75, 
    260.05, 259.75, 259.85, 259.55, 259.55, 260.05, 260.85, 260.05, 260.55, 
    261.05, 260.55, 261.35, 260.85, 260.95, 260.85, 260.85, 261.25, 261.05, 
    261.65, 262.05, 262.65, 263.95, 264.85, 264.85, 265.05, 266.25, 266.15, 
    266.15, 266.45, 266.85, 267.55, 267.85, 268.75, 269.15, 269.25, 269.05, 
    268.35, 269.55, 269.85, 270.25, 269.35, 269.75, 269.35, 269.45, 269.75, 
    270.35, 270.75, 270.85, 271.35, 271.25, 271.35, 270.65, 271.65, 272.35, 
    271.65, 271.45, 271.55, 272.85, 272.65, 270.55, 272.05, 270.95, 270.65, 
    270.85, 270.65, 271.35, 271.85, 271.65, 271.35, 271.65, 271.75, 271.95, 
    272.25, 272.45, 272.65, 272.85, 272.25, 273.55, 271.85, 270.15, 270.15, 
    270.75, 270.55, 268.25, 267.85, 267.75, 269.45, 270.45, 270.65, 270.35, 
    268.45, 268.55, 268.35, 268.15, 269.15, 269.35, 268.65, 268.55, 269.15, 
    269.15, 269.45, 269.95, 269.95, 269.45, 270.05, 270.25, 270.95, 271.05, 
    271.75, 272.45, 272.75, 272.85, 273.05, 273.25, 273.75, 273.35, 273.45, 
    272.65, 273.55, 273.45, 273.05, 273.05, 272.95, 272.85, 272.75, 272.85, 
    272.65, 272.65, 272.75, 272.85, 274.55, 274.65, 273.85, 274.35, 274.15, 
    273.55, 272.85, 272.45, 272.15, 271.25, 270.95, 270.35, 270.15, 269.65, 
    269.45, 269.35, 269.25, 268.95, 268.55, 267.85, 267.25, 267.75, 268.35, 
    268.65, 269.75, 273.15, 274.05, 274.45, 273.55, 272.95, 272.15, 272.25, 
    273.15, 272.55, 272.75, 273.05, 273.25, 273.15, 272.45, 271.75, 272.05, 
    271.85, 272.35, 272.05, 271.85, 270.75, 269.75, 269.95, 270.05, 269.25, 
    269.65, 269.25, 269.45, 269.95, 270.15, 268.65, 268.45, 268.75, 269.35, 
    270.95, 271.65, 271.45, 270.45, 273.75, 274.05, 274.65, 274.75, 274.85, 
    274.25, 275.15, 273.65, 273.55, 273.55, 273.85, 276.55, 276.85, 277.15, 
    276.35, 276.65, 275.35, 275.55, 275.55, 274.75, 275.45, 273.95, 273.55, 
    273.55, 274.15, 273.85, 273.15, 273.45, 273.15, 273.45, 273.95, 273.55, 
    272.65, 273.45, 274.15, 274.35, 274.35, 273.95, 273.35, 274.95, 274.95, 
    274.75, 275.15, 274.55, 274.65, 274.65, 274.65, 274.05, 274.15, 273.85, 
    273.55, 273.75, 273.35, 273.15, 271.85, 271.05, 270.45, 269.95, 268.15, 
    267.85, 269.45, 267.85, 268.05, 267.75, 268.25, 267.55, 268.25, 267.95, 
    268.05, 268.15, 268.15, 267.95, 268.25, 268.45, 269.35, 269.05, 269.25, 
    269.25, 268.85, 268.55, 268.45, 270.25, 270.05, 270.25, 268.55, 268.25, 
    267.95, 268.15, 267.45, 266.35, 266.85, 266.45, 266.45, 267.05, 266.15, 
    266.35, 266.85, 266.85, 266.85, 267.55, 268.05, 267.65, 267.95, 267.35, 
    266.85, 267.45, 267.75, 267.95, 267.25, 265.85, 266.85, 267.15, 267.05, 
    266.85, 266.25, 265.35, 264.75, 264.95, 264.75, 264.25, 264.85, 265.15, 
    264.65, 265.35, 266.75, 265.55, 266.05, 268.45, 266.35, 267.45, 271.25, 
    270.55, 269.75, 269.95, 270.25, 271.15, 271.65, 272.75, 272.75, 272.45, 
    272.15, 272.05, 272.35, 272.25, 271.35, 271.35, 270.75, 270.25, 270.65, 
    269.75, 268.95, 268.15, 268.95, 267.45, 266.65, 267.55, 267.65, 267.35, 
    267.05, 267.25, 266.85, 267.05, 266.95, 266.45, 266.75, 266.95, 266.45, 
    263.25, 263.75, 265.15, 263.45, 264.05, 262.75, 264.55, 265.75, 268.55, 
    269.35, 269.65, 268.85, 269.75, 269.85, 270.15, 269.45, 268.85, 268.15, 
    267.85, 267.95, 268.45, 268.25, 267.95, 267.85, 268.15, 268.45, 268.75, 
    268.85, 268.95, 269.15, 269.45, 269.75, 269.85, 269.95, 269.75, 269.85, 
    269.75, 269.65, 269.55, 269.15, 268.75, 268.45, 268.35, 268.25, 267.85, 
    267.85, 267.55, 268.05, 268.35, 268.75, 268.55, 268.05, 268.15, 267.85, 
    267.85, 267.65, 267.45, 267.25, 266.45, 266.95, 266.85, 266.95, 267.05, 
    266.15, 266.35, 265.85, 265.65, 265.05, 265.05, 265.05, 264.75, 264.85, 
    264.85, 264.85, 265.05, 265.05, 264.85, 264.95, 264.85, 264.75, 265.05, 
    265.25, 265.15, 265.65, 265.45, 265.25, 264.55, 264.55, 264.85, 264.75, 
    264.55, 264.55, 264.75, 264.45, 264.45, 264.35, 264.35, 264.75, 264.05, 
    264.15, 264.05, 264.15, 264.15, 264.55, 264.25, 264.55, 264.55, 264.55, 
    264.35, 265.15, 265.45, 265.15, 264.35, 263.45, 262.05, 262.95, 263.35, 
    263.35, 266.35, 264.25, 266.75, 265.05, 266.55, 264.95, 266.55, 264.15, 
    266.05, 267.35, 267.25, 266.55, 266.75, 266.65, 265.75, 266.45, 266.65, 
    266.05, 266.15, 268.45, 268.25, 268.65, 268.55, 269.15, 269.15, 269.05, 
    269.55, 269.65, 269.05, 267.95, 267.55, 266.75, 267.75, 265.55, 265.35, 
    265.45, 264.25, 264.35, 264.85, 264.85, 264.95, 264.95, 264.85, 265.05, 
    265.05, 263.55, 263.35, 264.65, 263.45, 263.35, 263.55, 263.35, 263.55, 
    263.25, 263.15, 263.15, 262.95, 261.95, 264.15, 264.35, 265.05, 266.05, 
    265.55, 265.45, 266.05, 266.35, 267.05, 266.65, 266.55, 265.75, 267.15, 
    266.15, 264.45, 263.85, 264.65, 265.55, 264.85, 266.05, 267.15, 268.05, 
    270.25, 270.85, 271.35, 272.15, 272.55, 272.25, 271.75, 270.75, 269.75, 
    267.45, 266.65, 266.25, 265.85, 265.85, 265.15, 265.35, 264.65, 263.75, 
    263.15, 264.65, 262.25, 263.65, 261.15, 261.35, 261.15, 261.15, 262.65, 
    263.85, 264.05, 265.35, 268.75, 271.25, 271.15, 271.55, 271.25, 270.65, 
    270.35, 270.25, 270.25, 270.05, 269.95, 269.25, 268.55, 267.95, 267.65, 
    266.95, 266.45, 265.95, 265.35, 265.05, 264.45, 264.25, 264.35, 264.45, 
    264.15, 264.05, 263.75, 263.95, 263.45, 263.15, 262.95, 262.65, 262.15, 
    262.25, 260.85, 260.15, 259.75, 260.35, 260.05, 260.55, 260.85, 260.85, 
    261.45, 261.55, 261.45, 261.05, 260.95, 260.55, 260.65, 260.85, 260.65, 
    260.85, 260.55, 261.15, 261.05, 260.85, 260.85, 261.05, 260.95, 260.85, 
    260.45, 260.15, 260.65, 260.55, 260.15, 259.65, 259.45, 259.55, 259.25, 
    259.25, 259.15, 259.25, 259.55, 259.65, 259.25, 259.05, 258.85, 258.35, 
    258.85, 258.45, 258.55, 258.95, 258.65, 258.65, 257.85, 257.85, 257.65, 
    256.85, 256.15, 255.95, 256.15, 255.75, 255.95, 256.25, 256.55, 256.15, 
    255.45, 255.45, 255.25, 255.45, 255.55, 255.85, 256.05, 256.35, 256.35, 
    256.85, 256.35, 257.25, 256.55, 254.45, 257.05, 256.25, 254.55, 254.35, 
    255.35, 255.95, 257.45, 256.85, 257.25, 257.95, 256.35, 256.75, 257.45, 
    258.55, 257.95, 257.55, 258.65, 259.05, 259.65, 260.05, 259.85, 260.15, 
    260.85, 260.55, 260.55, 260.15, 259.05, 260.05, 261.05, 261.15, 260.05, 
    258.65, 259.45, 259.85, 259.85, 259.15, 260.85, 259.95, 259.65, 259.35, 
    259.65, 260.45, 260.75, 261.55, 259.35, 260.05, 259.35, 260.55, 260.05, 
    262.15, 262.25, 262.25, 261.35, 262.65, 262.35, 262.25, 262.15, 262.05, 
    262.05, 260.65, 261.15, 261.25, 260.15, 259.15, 260.45, 261.55, 260.15, 
    260.85, 262.35, 261.75, 262.25, 263.05, 262.65, 263.45, 263.65, 264.15, 
    264.65, 264.75, 264.75, 264.85, 265.15, 264.45, 264.85, 264.85, 265.05, 
    265.55, 265.05, 266.15, 265.95, 264.75, 265.65, 265.05, 265.25, 266.15, 
    264.85, 263.75, 262.95, 263.65, 264.35, 265.15, 263.15, 262.85, 263.65, 
    263.65, 264.15, 263.05, 263.25, 262.95, 262.65, 262.25, 263.35, 264.95, 
    263.85, 264.25, 264.65, 264.95, 265.25, 265.05, 264.85, 265.25, 265.25, 
    265.85, 265.95, 266.55, 267.15, 266.55, 267.25, 267.55, 270.65, 273.35, 
    274.05, 274.45, 274.45, 274.45, 274.05, 273.55, 275.05, 272.15, 273.55, 
    274.25, 274.25, 273.45, 273.15, 273.05, 272.25, 271.55, 271.85, 271.25, 
    269.85, 269.35, 268.35, 267.75, 267.15, 265.85, 265.25, 264.25, 263.55, 
    262.15, 262.15, 261.55, 260.05, 258.05, 257.25, 256.35, 256.15, 256.05, 
    256.25, 255.95, 255.85, 256.65, 256.35, 255.45, 257.35, 255.25, 256.45, 
    256.35, 256.15, 257.25, 257.35, 257.85, 258.65, 258.45, 256.25, 255.35, 
    257.45, 254.25, 254.95, 253.65, 255.75, 255.65, 255.55, 256.55, 256.85, 
    256.35, 256.25, 254.85, 255.65, 255.55, 256.15, 256.55, 255.45, 256.75, 
    257.45, 256.95, 256.15, 256.05, 257.45, 258.35, 256.85, 257.95, 258.15, 
    258.05, 258.45, 258.75, 259.05, 259.25, 260.25, 259.85, 260.45, 262.15, 
    261.85, 261.15, 262.75, 262.05, 262.25, 261.75, 261.55, 260.95, 261.75, 
    261.45, 261.55, 261.55, 261.15, 260.65, 259.75, 259.85, 259.95, 260.05, 
    261.35, 261.75, 262.05, 262.35, 262.75, 262.35, 262.85, 262.75, 264.05, 
    264.65, 265.35, 266.85, 267.25, 267.45, 266.95, 267.05, 267.05, 266.75, 
    266.55, 266.45, 265.85, 266.15, 265.55, 262.05, 260.85, 260.55, 261.75, 
    260.55, 262.45, 262.15, 262.25, 261.65, 259.45, 262.15, 262.05, 261.85, 
    261.65, 262.55, 262.05, 261.95, 260.65, 259.25, 258.85, 259.35, 258.65, 
    257.45, 258.85, 258.35, 258.55, 259.65, 258.45, 256.85, 257.65, 258.85, 
    259.25, 259.05, 257.85, 258.35, 259.35, 258.25, 258.45, 259.75, 260.25, 
    259.55, 261.55, 260.65, 262.95, 263.15, 262.45, 263.95, 262.15, 263.55, 
    264.25, 264.75, 265.25, 265.75, 265.75, 265.45, 266.35, 266.75, 266.85, 
    267.45, 269.05, 269.65, 270.85, 271.75, 271.75, 271.75, 271.15, 269.15, 
    267.65, 266.45, 265.45, 264.65, 263.95, 263.45, 263.25, 262.65, 262.75, 
    262.95, 263.75, 263.55, 263.05, 263.15, 262.75, 262.55, 262.45, 262.25, 
    262.35, 261.95, 262.05, 262.05, 261.85, 261.95, 261.65, 261.65, 261.35, 
    261.15, 260.45, 259.75, 259.15, 258.65, 258.05, 257.45, 257.15, 257.15, 
    257.15, 256.65, 256.75, 256.15, 254.35, 256.65, 254.35, 251.85, 253.75, 
    253.65, 253.95, 254.25, 251.85, 252.65, 252.85, 253.45, 253.85, 252.45, 
    252.15, 253.85, 253.55, 253.55, 253.95, 253.95, 253.55, 254.15, 254.05, 
    253.95, 252.75, 254.75, 255.25, 255.75, 256.55, 256.55, 256.45, 256.35, 
    256.45, 256.05, 254.65, 253.15, 253.45, 253.85, 253.35, 253.95, 253.15, 
    252.65, 253.15, 251.85, 252.85, 252.05, 252.55, 252.95, 251.45, 251.85, 
    252.75, 251.75, 254.25, 252.85, 251.55, 253.65, 253.65, 251.85, 251.45, 
    252.65, 252.75, 252.65, 251.05, 251.75, 250.35, 252.25, 252.35, 253.05, 
    252.85, 252.65, 253.35, 253.55, 253.85, 253.85, 254.65, 255.45, 255.55, 
    255.35, 255.35, 255.35, 253.55, 251.45, 251.75, 250.95, 251.15, 253.35, 
    253.85, 251.75, 252.45, 251.85, 250.65, 249.95, 252.45, 252.95, 248.45, 
    250.75, 250.95, 252.95, 252.95, 252.85, 253.15, 253.35, 253.15, 253.35, 
    253.85, 253.55, 254.15, 252.75, 255.35, 255.95, 256.35, 257.05, 256.75, 
    256.55, 256.85, 257.15, 257.05, 256.05, 255.75, 256.95, 257.15, 256.35, 
    256.45, 252.55, 252.45, 255.45, 255.85, 254.75, 254.75, 254.55, 253.55, 
    254.25, 253.75, 253.35, 252.85, 252.85, 252.05, 253.55, 253.45, 253.45, 
    254.25, 254.45, 254.75, 255.25, 256.25, 256.55, 256.75, 256.65, 257.05, 
    257.65, 259.05, 259.15, 259.85, 260.65, 261.55, 262.35, 263.15, 263.65, 
    263.65, 263.15, 264.15, 262.35, 263.75, 264.45, 263.55, 263.65, 264.25, 
    263.75, 262.75, 263.55, 263.45, 263.35, 264.25, 264.55, 265.05, 265.85, 
    266.25, 267.25, 267.35, 268.05, 268.15, 268.45, 268.35, 267.95, 268.85, 
    268.15, 269.35, 269.35, 269.55, 270.25, 270.55, 270.55, 270.55, 271.35, 
    270.85, 270.75, 271.15, 271.35, 271.05, 271.95, 272.05, 272.25, 272.85, 
    272.95, 272.55, 272.25, 272.85, 272.35, 272.15, 272.85, 273.45, 272.25, 
    271.55, 270.75, 270.45, 270.15, 269.75, 269.55, 269.15, 269.25, 269.35, 
    270.25, 270.15, 270.35, 270.55, 270.45, 270.55, 270.75, 270.65, 270.45, 
    270.35, 270.15, 270.45, 270.55, 272.45, 273.45, 275.45, 275.75, 275.65, 
    276.55, 276.25, 276.95, 276.55, 276.55, 276.15, 276.75, 276.25, 277.05, 
    276.85, 276.65, 276.45, 276.65, 276.65, 276.85, 276.65, 276.75, 276.15, 
    276.25, 276.55, 275.75, 275.15, 276.95, 276.15, 275.85, 275.65, 275.85, 
    276.05, 275.75, 275.65, 276.45, 275.65, 275.75, 276.05, 276.75, 276.55, 
    275.85, 277.05, 277.15, 276.95, 277.15, 276.85, 276.55, 276.75, 277.15, 
    276.35, 276.45, 275.95, 275.95, 275.95, 275.65, 276.05, 276.65, 276.85, 
    276.75, 276.75, 276.45, 276.35, 276.45, 276.35, 276.05, 276.75, 276.05, 
    276.05, 276.15, 275.95, 275.85, 275.95, 276.65, 276.15, 275.85, 276.05, 
    276.05, 276.15, 276.15, 276.45, 276.05, 276.45, 276.65, 276.15, 276.05, 
    276.25, 276.35, 275.95, 275.95, 275.65, 276.25, 275.75, 275.75, 275.75, 
    275.65, 275.65, 275.95, 276.15, 275.35, 276.05, 275.95, 276.15, 275.95, 
    275.85, 275.85, 276.15, 276.05, 275.85, 275.55, 275.15, 275.35, 274.95, 
    274.75, 274.95, 274.25, 274.65, 274.75, 275.15, 275.05, 275.55, 275.05, 
    274.65, 275.05, 276.05, 275.95, 275.35, 275.95, 275.05, 275.55, 276.25, 
    275.65, 275.45, 275.45, 275.95, 276.35, 276.05, 276.55, 276.45, 276.15, 
    275.65, 274.95, 274.85, 275.05, 275.05, 274.85, 274.75, 274.75, 274.85, 
    274.85, 274.65, 274.85, 274.65, 273.95, 274.55, 273.95, 274.65, 274.55, 
    274.75, 274.35, 274.05, 273.65, 273.55, 273.55, 273.85, 273.55, 272.45, 
    272.35, 272.15, 271.85, 274.15, 274.65, 274.25, 274.35, 274.55, 274.85, 
    274.45, 273.35, 271.95, 271.05, 271.55, 271.35, 269.45, 268.25, 267.95, 
    268.35, 267.05, 266.25, 266.15, 266.55, 266.25, 266.05, 265.25, 265.25, 
    265.15, 264.85, 264.75, 264.75, 264.15, 263.75, 263.45, 263.15, 262.75, 
    263.15, 263.25, 262.75, 262.15, 262.25, 261.65, 261.25, 260.15, 261.05, 
    260.65, 259.45, 259.25, 258.15, 259.15, 258.95, 258.15, 258.55, 258.45, 
    257.55, 257.65, 258.05, 259.35, 258.55, 259.05, 258.95, 258.85, 258.75, 
    258.95, 259.15, 259.75, 260.55, 260.95, 261.75, 262.45, 262.35, 262.85, 
    262.95, 263.45, 263.55, 263.75, 264.15, 265.25, 264.85, 263.65, 262.95, 
    262.15, 261.45, 261.05, 260.35, 259.55, 258.75, 258.15, 257.95, 257.45, 
    256.85, 256.65, 256.35, 256.05, 256.45, 256.05, 255.75, 255.55, 255.55, 
    255.35, 255.85, 256.05, 255.05, 255.75, 255.75, 256.15, 254.75, 254.75, 
    254.75, 254.55, 254.45, 254.35, 253.95, 254.05, 253.35, 253.35, 253.75, 
    253.55, 253.35, 253.45, 253.05, 252.95, 253.05, 253.15, 253.45, 253.35, 
    254.75, 252.95, 254.65, 253.55, 252.75, 253.45, 253.05, 253.15, 252.25, 
    252.45, 251.55, 252.75, 251.95, 252.15, 252.25, 252.25, 252.05, 252.15, 
    251.95, 252.15, 252.85, 253.55, 253.65, 252.95, 252.75, 252.85, 253.45, 
    253.55, 253.95, 253.75, 254.25, 254.05, 254.05, 254.85, 255.35, 256.05, 
    256.15, 256.75, 257.15, 257.65, 258.05, 258.65, 259.05, 259.55, 262.15, 
    262.45, 262.25, 262.15, 262.35, 262.05, 261.95, 261.65, 261.45, 261.45, 
    260.75, 261.55, 261.45, 260.55, 260.05, 259.55, 258.95, 259.45, 258.85, 
    259.05, 258.85, 258.35, 258.35, 258.45, 258.45, 259.05, 260.05, 261.05, 
    263.65, 265.75, 266.15, 266.65, 267.55, 268.15, 268.75, 269.05, 269.45, 
    269.65, 269.15, 269.05, 268.85, 269.55, 270.05, 269.95, 269.15, 268.85, 
    268.45, 268.25, 267.45, 266.65, 266.55, 266.25, 266.15, 266.15, 265.35, 
    264.75, 263.25, 262.25, 261.65, 260.95, 260.85, 260.55, 260.25, 260.55, 
    260.75, 260.95, 261.35, 261.85, 261.95, 262.35, 261.75, 262.25, 262.15, 
    262.15, 261.95, 262.05, 261.75, 261.05, 260.75, 260.85, 260.55, 260.45, 
    260.35, 260.55, 260.75, 260.65, 260.85, 261.25, 261.45, 261.35, 261.25, 
    261.15, 260.85, 260.65, 260.55, 260.15, 260.05, 260.15, 260.15, 260.05, 
    260.35, 260.45, 260.55, 260.85, 261.25, 261.65, 262.25, 262.75, 263.15, 
    263.65, 264.35, 264.65, 264.95, 265.25, 265.45, 265.25, 265.35, 265.45, 
    265.75, 265.35, 265.55, 264.45, 264.05, 263.85, 263.85, 263.35, 263.65, 
    263.25, 263.55, 262.25, 261.95, 261.55, 260.25, 260.35, 260.35, 259.05, 
    258.55, 257.75, 258.45, 257.55, 258.45, 258.75, 259.15, 257.55, 258.25, 
    258.55, 258.25, 257.25, 258.15, 258.25, 257.45, 258.75, 257.35, 258.05, 
    256.95, 256.85, 256.65, 256.65, 257.45, 256.45, 257.15, 258.05, 258.15, 
    258.05, 259.35, 258.25, 257.95, 259.55, 260.45, 258.95, 260.35, 260.55, 
    260.45, 260.45, 260.05, 259.75, 259.95, 260.05, 259.75, 259.35, 259.05, 
    258.85, 259.25, 260.65, 260.45, 259.75, 260.45, 260.65, 259.65, 259.95, 
    259.25, 260.15, 260.55, 261.05, 262.55, 261.55, 260.55, 261.45, 262.35, 
    262.65, 262.75, 261.85, 261.15, 261.55, 262.25, 261.95, 261.75, 261.55, 
    260.85, 261.75, 262.95, 260.45, 260.45, 261.35, 261.25, 261.65, 260.75, 
    259.35, 260.55, 260.35, 261.75, 261.65, 259.45, 259.05, 260.05, 258.25, 
    258.95, 259.35, 259.35, 257.45, 258.65, 259.95, 258.15, 258.55, 258.05, 
    257.95, 259.55, 258.85, 259.35, 259.25, 257.65, 258.55, 258.45, 258.35, 
    260.55, 260.45, 259.75, 258.55, 259.05, 259.85, 258.95, 259.05, 258.95, 
    259.05, 258.55, 257.55, 259.75, 259.15, 259.15, 259.95, 260.35, 259.05, 
    260.45, 261.05, 260.85, 261.35, 262.15, 261.35, 262.65, 262.65, 262.35, 
    262.15, 259.95, 261.45, 260.55, 260.65, 260.85, 259.85, 261.25, 261.55, 
    260.55, 259.85, 260.15, 260.25, 260.75, 260.75, 260.85, 261.25, 261.25, 
    260.85, 260.65, 261.55, 261.85, 262.25, 262.15, 262.05, 261.55, 261.55, 
    261.15, 262.75, 279.15, 262.35, 263.15, 263.05, 264.45, 263.95, 263.15, 
    263.85, 264.55, 265.15, 264.95, 265.15, 265.45, 265.05, 265.45, 265.55, 
    265.75, 265.95, 266.25, 266.45, 266.55, 266.75, 266.75, 266.95, 267.05, 
    266.85, 267.25, 267.25, 267.35, 267.25, 267.25, 267.55, 267.65, 267.45, 
    268.45, 268.15, 267.75, 267.45, 267.95, 267.95, 268.05, 267.95, 267.15, 
    266.65, 266.15, 264.65, 264.15, 263.45, 261.85, 260.85, 260.15, 260.15, 
    259.35, 258.65, 258.65, 258.55, 258.55, 258.05, 258.55, 258.45, 258.35, 
    258.55, 258.65, 258.85, 259.05, 259.25, 259.65, 259.65, 260.35, 260.45, 
    260.55, 261.15, 261.55, 261.45, 261.55, 262.65, 263.05, 262.65, 262.55, 
    262.25, 263.55, 263.95, 264.15, 264.75, 265.35, 265.75, 266.35, 266.75, 
    266.95, 267.25, 267.35, 266.65, 267.05, 266.65, 266.55, 266.55, 266.85, 
    267.05, 267.05, 267.05, 267.45, 267.25, 267.55, 267.45, 267.75, 268.05, 
    268.95, 268.65, 268.75, 268.35, 267.85, 265.95, 266.15, 265.85, 265.95, 
    266.15, 265.55, 264.85, 264.85, 264.75, 264.35, 263.55, 262.45, 263.05, 
    264.75, 264.65, 264.45, 264.35, 263.95, 263.85, 263.75, 263.55, 263.35, 
    263.25, 263.05, 262.75, 262.75, 262.85, 262.65, 261.65, 261.05, 259.55, 
    260.55, 260.85, 260.55, 260.55, 260.35, 260.75, 260.75, 260.75, 260.55, 
    260.95, 260.85, 260.85, 261.25, 261.75, 261.95, 261.85, 261.25, 261.35, 
    260.85, 258.35, 255.15, 254.55, 253.55, 252.55, 252.55, 252.15, 252.15, 
    251.85, 251.75, 251.75, 251.05, 250.65, 249.95, 249.65, 249.65, 248.85, 
    248.75, 248.25, 248.35, 248.45, 249.05, 249.95, 248.85, 248.55, 248.65, 
    248.55, 249.15, 249.55, 250.25, 250.75, 250.75, 251.35, 251.65, 252.25, 
    254.15, 253.95, 255.35, 254.45, 255.55, 256.75, 255.85, 254.65, 254.85, 
    253.65, 254.25, 254.85, 254.65, 254.05, 254.15, 253.55, 253.05, 252.65, 
    254.05, 254.65, 254.75, 256.05, 256.55, 257.45, 258.05, 258.45, 259.15, 
    259.65, 259.65, 260.65, 261.05, 261.15, 261.65, 262.25, 263.05, 263.75, 
    264.95, 265.05, 266.35, 267.45, 267.85, 267.45, 267.25, 267.15, 267.95, 
    267.95, 268.35, 268.05, 268.85, 269.55, 269.75, 269.95, 270.55, 270.45, 
    271.15, 271.85, 271.75, 271.85, 273.05, 272.85, 272.95, 273.65, 272.85, 
    272.85, 272.45, 271.95, 271.55, 273.35, 273.45, 273.65, 273.85, 273.75, 
    273.35, 272.95, 272.65, 272.35, 271.75, 271.45, 270.85, 270.25, 270.05, 
    269.85, 268.95, 268.75, 268.35, 268.35, 267.75, 267.15, 266.55, 265.75, 
    265.25, 264.65, 264.05, 263.65, 263.15, 262.45, 261.85, 261.45, 260.85, 
    260.25, 259.65, 258.85, 258.55, 258.05, 257.65, 258.55, 258.25, 257.75, 
    257.15, 257.25, 256.75, 256.65, 256.55, 256.35, 256.15, 255.95, 255.85, 
    255.75, 254.75, 254.45, 254.65, 253.95, 253.65, 254.15, 254.25, 252.95, 
    254.25, 254.45, 254.45, 253.95, 253.45, 253.55, 253.05, 252.95, 252.55, 
    252.25, 252.85, 252.45, 251.65, 251.65, 251.25, 251.05, 250.65, 250.75, 
    250.75, 250.05, 250.45, 249.85, 249.35, 249.05, 248.95, 248.55, 248.55, 
    249.05, 249.55, 250.15, 250.35, 249.45, 249.95, 247.75, 247.75, 247.35, 
    248.45, 247.75, 246.85, 248.15, 247.25, 248.35, 248.75, 249.15, 249.35, 
    250.25, 251.35, 251.65, 251.75, 251.85, 251.55, 252.75, 253.15, 253.05, 
    253.95, 253.05, 253.95, 254.15, 255.05, 256.15, 255.85, 256.45, 256.65, 
    256.45, 257.15, 256.35, 255.65, 255.45, 255.35, 255.15, 254.95, 254.55, 
    253.95, 253.55, 253.85, 253.95, 254.05, 253.65, 254.65, 254.75, 255.25, 
    255.45, 254.35, 254.35, 255.45, 253.75, 254.05, 254.95, 255.75, 254.05, 
    255.25, 254.75, 254.05, 254.85, 254.85, 254.75, 254.65, 255.95, 256.95, 
    256.75, 257.05, 257.45, 259.45, 258.95, 259.25, 259.35, 258.35, 257.05, 
    258.85, 255.55, 256.45, 257.35, 258.05, 257.05, 256.85, 258.15, 256.35, 
    257.35, 258.85, 258.95, 259.95, 258.85, 258.85, 259.95, 259.65, 260.45, 
    261.15, 262.25, 262.25, 261.45, 262.25, 262.65, 261.65, 265.15, 264.65, 
    265.15, 265.55, 265.45, 265.35, 264.95, 264.85, 264.65, 264.55, 263.55, 
    264.65, 263.75, 263.55, 263.95, 264.55, 264.95, 264.85, 264.85, 264.95, 
    264.85, 265.65, 265.35, 263.55, 262.35, 261.55, 260.55, 260.25, 260.65, 
    259.75, 259.35, 260.55, 258.75, 258.75, 258.65, 258.85, 258.95, 259.45, 
    258.35, 259.85, 258.55, 258.15, 258.55, 259.45, 259.85, 260.35, 259.55, 
    259.35, 258.15, 257.65, 257.75, 257.25, 256.95, 256.55, 255.35, 254.45, 
    255.05, 254.45, 255.75, 256.05, 256.15, 258.15, 258.65, 259.85, 260.45, 
    261.45, 261.85, 262.05, 261.65, 262.05, 263.75, 263.05, 263.05, 263.35, 
    263.65, 263.55, 262.75, 263.15, 263.05, 262.65, 262.65, 262.25, 262.55, 
    262.45, 262.65, 262.55, 262.35, 261.75, 260.35, 260.65, 259.85, 258.25, 
    257.55, 256.15, 255.95, 255.55, 255.05, 254.15, 254.15, 253.95, 253.45, 
    251.15, 252.85, 253.75, 253.75, 253.45, 252.85, 252.45, 251.95, 252.25, 
    252.65, 252.55, 251.75, 251.85, 252.05, 252.25, 254.05, 254.05, 254.85, 
    254.55, 254.85, 254.35, 253.95, 254.25, 255.95, 256.25, 253.25, 252.75, 
    253.95, 256.15, 254.15, 254.05, 252.85, 254.25, 252.45, 252.95, 254.15, 
    252.95, 253.55, 252.55, 253.75, 252.75, 254.25, 255.05, 254.65, 254.25, 
    253.65, 253.05, 253.25, 252.95, 253.05, 252.35, 251.55, 251.45, 251.35, 
    251.45, 252.25, 252.85, 252.95, 253.45, 253.65, 254.85, 254.45, 255.35, 
    254.75, 255.25, 255.15, 255.25, 253.55, 253.95, 253.65, 253.75, 253.45, 
    252.85, 253.35, 253.15, 253.35, 253.55, 253.25, 253.75, 254.35, 254.15, 
    253.65, 254.25, 255.05, 255.85, 256.75, 257.75, 257.85, 257.25, 256.95, 
    257.35, 255.95, 256.05, 254.15, 255.75, 255.35, 255.35, 254.65, 254.35, 
    254.95, 254.35, 255.55, 254.15, 255.05, 254.45, 254.45, 255.85, 258.05, 
    257.65, 257.25, 255.15, 256.15, 255.25, 255.55, 254.75, 253.45, 252.95, 
    252.85, 252.65, 252.35, 252.65, 252.35, 251.45, 251.45, 250.75, 249.45, 
    249.05, 249.05, 249.85, 250.75, 250.95, 251.95, 253.65, 253.25, 253.95, 
    253.55, 253.95, 254.75, 255.35, 254.25, 253.25, 254.25, 253.35, 253.75, 
    253.25, 252.25, 253.25, 254.35, 253.95, 252.95, 253.85, 254.05, 254.15, 
    255.75, 256.15, 258.55, 258.75, 258.25, 259.95, 259.35, 258.25, 256.75, 
    258.95, 258.45, 258.85, 258.85, 258.05, 258.75, 260.15, 260.35, 260.15, 
    259.85, 260.05, 260.15, 259.65, 260.55, 260.15, 260.65, 260.35, 260.55, 
    260.95, 260.95, 261.05, 260.85, 262.05, 260.95, 261.45, 261.05, 260.15, 
    259.75, 259.15, 257.95, 257.85, 257.05, 256.15, 254.95, 254.95, 254.45, 
    254.15, 254.25, 254.45, 254.75, 255.15, 255.65, 256.05, 256.95, 255.55, 
    255.15, 255.55, 255.95, 255.35, 254.55, 253.75, 253.35, 253.55, 253.25, 
    252.95, 253.15, 253.35, 253.45, 254.55, 255.75, 256.75, 258.15, 259.45, 
    262.65, 263.55, 262.55, 264.45, 264.25, 264.35, 263.95, 264.55, 264.35, 
    262.85, 263.45, 264.05, 264.75, 264.85, 263.05, 261.75, 262.75, 261.35, 
    263.25, 262.35, 261.65, 261.25, 262.65, 262.85, 262.95, 262.85, 264.25, 
    264.55, 265.75, 264.85, 265.15, 264.45, 264.35, 264.05, 263.75, 260.55, 
    261.25, 260.35, 261.35, 262.15, 259.85, 261.35, 260.55, 259.25, 259.85, 
    260.35, 261.35, 261.65, 262.95, 263.35, 264.75, 265.85, 265.85, 266.55, 
    263.85, 266.95, 264.65, 265.75, 264.65, 263.45, 261.65, 262.65, 260.85, 
    262.05, 262.85, 260.55, 262.65, 260.25, 260.55, 259.95, 260.75, 263.45, 
    264.35, 263.85, 263.45, 264.55, 264.75, 264.45, 265.25, 266.55, 267.85, 
    267.15, 268.75, 268.05, 267.85, 268.45, 268.75, 268.65, 268.35, 269.25, 
    269.15, 270.15, 269.75, 269.35, 269.15, 269.05, 269.55, 269.95, 269.75, 
    270.85, 269.95, 272.05, 271.65, 271.55, 271.35, 271.65, 271.25, 270.85, 
    271.25, 270.95, 270.55, 270.75, 270.75, 270.75, 270.05, 270.25, 270.75, 
    270.35, 269.95, 269.85, 269.85, 269.95, 270.65, 270.55, 270.75, 270.65, 
    270.25, 268.35, 268.65, 267.55, 267.65, 266.65, 264.85, 265.15, 263.95, 
    263.25, 262.75, 262.15, 261.85, 262.55, 260.75, 260.75, 260.65, 263.65, 
    264.65, 264.15, 264.05, 264.95, 266.55, 267.25, 267.05, 265.65, 265.15, 
    264.85, 263.45, 261.05, 260.95, 260.95, 261.55, 261.55, 262.65, 260.45, 
    260.75, 262.45, 262.75, 263.05, 264.05, 263.55, 263.55, 265.35, 265.75, 
    267.95, 266.85, 267.95, 267.05, 267.45, 268.15, 265.55, 265.55, 265.55, 
    262.75, 262.05, 263.15, 262.25, 260.45, 261.05, 261.35, 261.75, 263.75, 
    264.05, 262.25, 263.35, 264.55, 265.65, 268.05, 266.75, 267.25, 264.95, 
    268.55, 267.75, 265.75, 264.55, 265.25, 264.15, 262.25, 263.45, 265.05, 
    264.45, 265.25, 266.05, 265.75, 265.55, 265.95, 264.25, 263.25, 262.85, 
    261.05, 261.05, 260.45, 260.55, 261.35, 260.65, 260.55, 260.35, 259.95, 
    258.55, 257.35, 256.75, 255.65, 253.85, 254.05, 253.85, 253.35, 251.65, 
    253.45, 253.95, 253.75, 254.25, 254.15, 254.55, 255.15, 256.45, 255.65, 
    256.15, 256.45, 256.45, 257.05, 256.55, 256.55, 256.35, 256.05, 255.55, 
    254.25, 254.15, 254.95, 255.15, 255.65, 255.95, 254.65, 254.35, 255.35, 
    255.05, 254.55, 254.85, 255.05, 255.65, 256.25, 257.35, 259.15, 257.75, 
    259.55, 256.85, 258.15, 258.15, 256.75, 255.65, 254.35, 253.75, 253.25, 
    253.85, 253.45, 254.45, 252.55, 254.65, 254.45, 255.25, 256.15, 257.45, 
    257.45, 259.75, 260.15, 261.25, 259.75, 261.75, 261.55, 262.85, 263.15, 
    263.45, 262.65, 262.65, 261.85, 261.45, 261.15, 263.15, 263.35, 262.65, 
    262.15, 262.35, 262.05, 262.55, 262.45, 261.85, 263.65, 265.05, 265.75, 
    265.25, 264.75, 263.45, 263.75, 263.85, 262.35, 263.15, 263.25, 261.45, 
    260.05, 258.85, 258.35, 258.55, 257.35, 255.95, 257.05, 257.35, 256.55, 
    257.15, 257.85, 261.95, 262.75, 263.15, 261.95, 262.35, 262.75, 262.85, 
    262.85, 263.55, 263.15, 262.75, 262.65, 262.45, 260.75, 260.25, 260.65, 
    259.65, 259.65, 259.85, 259.65, 261.65, 261.55, 261.75, 261.65, 262.35, 
    264.75, 266.25, 267.35, 267.95, 267.85, 267.95, 269.25, 269.65, 269.65, 
    270.75, 270.15, 270.35, 269.85, 269.35, 268.25, 268.25, 267.55, 267.55, 
    267.35, 267.15, 267.85, 268.85, 268.95, 268.75, 268.65, 268.85, 269.35, 
    269.35, 269.65, 269.65, 269.75, 269.55, 269.65, 269.35, 269.25, 269.05, 
    269.15, 269.15, 270.05, 269.05, 270.05, 269.55, 269.35, 268.05, 267.05, 
    266.75, 267.15, 266.95, 267.95, 268.65, 268.65, 268.95, 269.05, 268.75, 
    269.05, 269.05, 268.75, 267.35, 267.15, 266.55, 264.85, 263.85, 263.25, 
    263.25, 263.05, 262.95, 260.85, 261.55, 262.55, 263.45, 263.75, 263.55, 
    263.85, 264.55, 263.75, 263.75, 264.25, 264.75, 265.35, 264.85, 265.25, 
    264.55, 264.95, 263.85, 263.15, 262.25, 261.45, 260.85, 259.35, 260.15, 
    260.65, 260.35, 259.55, 258.95, 259.35, 261.55, 262.45, 263.45, 263.05, 
    265.85, 264.35, 264.05, 264.85, 264.35, 264.05, 263.15, 263.35, 262.85, 
    260.95, 260.25, 259.25, 258.55, 257.95, 258.25, 258.75, 258.55, 258.05, 
    258.95, 260.15, 260.75, 262.05, 264.15, 264.85, 264.95, 264.65, 265.45, 
    264.25, 264.25, 263.75, 263.45, 263.35, 262.75, 261.65, 261.05, 259.95, 
    260.15, 260.35, 260.15, 259.35, 259.25, 259.35, 261.35, 262.35, 263.35, 
    263.35, 263.05, 263.55, 263.85, 264.15, 264.85, 265.15, 265.35, 265.65, 
    265.55, 265.55, 265.05, 264.95, 264.85, 264.55, 264.45, 264.45, 264.35, 
    267.45, 268.05, 268.35, 268.75, 269.45, 269.75, 270.45, 269.75, 269.45, 
    269.45, 268.15, 268.85, 268.45, 269.15, 268.65, 267.75, 267.85, 267.85, 
    267.75, 268.45, 267.95, 268.35, 269.45, 269.95, 270.55, 273.15, 273.65, 
    273.45, 273.55, 273.45, 274.25, 274.95, 275.95, 275.05, 274.75, 274.65, 
    274.05, 273.85, 274.35, 274.95, 274.35, 273.95, 273.75, 274.35, 274.85, 
    275.05, 275.15, 274.85, 274.75, 274.75, 275.15, 274.75, 275.25, 275.35, 
    275.45, 275.45, 275.55, 275.85, 276.15, 275.75, 275.35, 274.65, 274.15, 
    271.65, 268.85, 268.35, 267.15, 266.05, 265.25, 264.25, 263.15, 263.25, 
    263.75, 264.85, 265.15, 265.55, 267.15, 267.15, 267.15, 267.05, 268.25, 
    268.25, 268.25, 268.65, 268.75, 269.55, 268.85, 268.95, 269.55, 269.45, 
    269.45, 269.45, 269.55, 269.45, 269.25, 269.45, 269.55, 269.45, 269.45, 
    269.15, 269.65, 270.05, 270.65, 270.85, 270.85, 271.55, 271.05, 271.45, 
    271.25, 271.55, 271.15, 271.05, 271.15, 269.95, 270.15, 269.95, 270.05, 
    270.05, 269.65, 269.55, 269.55, 269.35, 269.05, 268.75, 268.45, 268.55, 
    268.55, 268.75, 268.95, 268.75, 269.35, 269.15, 268.85, 268.45, 268.05, 
    267.55, 267.45, 266.95, 266.25, 266.65, 266.85, 267.05, 267.05, 267.55, 
    268.05, 267.65, 268.05, 268.85, 268.75, 269.25, 269.15, 269.55, 269.15, 
    268.95, 268.95, 269.45, 269.75, 269.95, 270.45, 273.65, 275.05, 274.95, 
    274.85, 275.05, 274.75, 274.75, 273.45, 273.25, 273.25, 273.55, 273.35, 
    273.35, 273.85, 274.75, 274.25, 274.05, 273.75, 273.05, 272.95, 272.55, 
    271.75, 271.55, 270.85, 270.85, 270.65, 269.15, 269.15, 269.35, 268.55, 
    268.15, 267.55, 267.25, 266.55, 265.75, 265.35, 265.45, 265.25, 265.15, 
    265.15, 264.95, 265.15, 265.25, 265.05, 265.25, 264.85, 264.55, 263.45, 
    266.25, 263.95, 263.35, 263.55, 262.35, 262.05, 261.65, 261.45, 260.95, 
    260.75, 258.85, 259.85, 260.85, 261.25, 262.05, 262.95, 262.85, 263.05, 
    261.45, 263.35, 261.75, 263.15, 264.45, 263.35, 263.15, 262.85, 262.95, 
    261.95, 262.05, 262.15, 262.65, 262.25, 262.55, 262.55, 263.15, 262.25, 
    263.05, 263.05, 263.25, 264.25, 264.25, 264.65, 264.45, 264.95, 265.15, 
    264.35, 264.45, 265.05, 264.35, 264.05, 263.05, 262.65, 261.85, 261.75, 
    261.65, 261.35, 261.05, 260.85, 260.35, 260.25, 260.55, 261.05, 261.55, 
    261.65, 262.05, 262.75, 262.45, 262.85, 262.35, 262.35, 261.85, 262.85, 
    262.35, 261.05, 261.85, 260.95, 260.15, 260.15, 259.95, 259.65, 259.25, 
    259.25, 259.05, 259.15, 259.45, 259.95, 260.55, 261.25, 261.05, 261.95, 
    261.85, 263.15, 262.65, 263.15, 263.25, 263.25, 263.75, 263.95, 262.95, 
    262.35, 261.95, 261.95, 262.05, 261.85, 261.85, 261.85, 261.65, 261.75, 
    262.05, 262.65, 263.05, 262.55, 262.85, 263.45, 264.05, 264.35, 265.55, 
    264.65, 264.35, 264.65, 264.35, 264.05, 264.15, 263.25, 262.65, 262.25, 
    262.05, 261.95, 261.65, 261.85, 260.75, 262.45, 263.05, 263.95, 264.65, 
    264.95, 265.45, 265.95, 266.35, 266.45, 266.15, 266.45, 266.25, 266.15, 
    265.95, 265.35, 264.95, 264.55, 263.85, 263.55, 263.15, 263.05, 262.35, 
    261.95, 261.25, 262.15, 262.55, 262.65, 263.65, 264.55, 265.05, 265.65, 
    265.65, 266.05, 266.25, 266.95, 267.15, 266.85, 266.45, 266.75, 265.75, 
    265.55, 264.45, 264.15, 263.85, 263.55, 263.85, 263.15, 262.85, 264.05, 
    263.55, 265.25, 265.35, 266.15, 267.75, 267.55, 267.25, 268.25, 268.05, 
    268.45, 268.25, 268.65, 269.55, 269.45, 269.25, 268.55, 267.85, 267.45, 
    267.05, 266.45, 266.55, 266.15, 265.85, 266.75, 266.95, 267.45, 268.25, 
    269.35, 269.55, 269.75, 270.65, 270.75, 271.45, 271.75, 272.05, 272.05, 
    271.25, 271.65, 271.25, 271.65, 271.65, 271.25, 270.15, 270.35, 269.75, 
    270.85, 272.95, 272.65, 272.55, 271.95, 272.15, 271.65, 271.65, 271.45, 
    270.55, 269.85, 270.05, 270.25, 270.25, 269.95, 269.55, 268.75, 267.15, 
    266.85, 265.55, 264.95, 263.75, 262.75, 262.25, 261.75, 261.85, 263.25, 
    264.25, 264.15, 265.75, 266.65, 266.15, 267.15, 268.05, 268.35, 269.05, 
    269.25, 268.85, 268.75, 268.65, 267.85, 267.75, 267.35, 265.75, 263.75, 
    264.45, 263.25, 263.35, 263.25, 262.85, 262.95, 263.75, 264.75, 266.05, 
    266.95, 266.35, 266.65, 267.45, 267.05, 267.65, 267.65, 267.15, 267.05, 
    267.35, 266.95, 266.85, 266.85, 266.65, 266.95, 266.95, 266.65, 266.65, 
    266.65, 266.75, 266.75, 266.95, 267.15, 267.45, 267.75, 268.05, 268.25, 
    268.85, 269.15, 269.65, 271.25, 270.85, 270.25, 269.35, 269.45, 269.15, 
    269.05, 268.75, 268.25, 268.45, 268.35, 268.55, 268.55, 268.25, 267.85, 
    267.65, 268.25, 268.85, 269.15, 269.95, 270.75, 270.65, 270.65, 270.75, 
    270.55, 270.35, 271.15, 271.55, 270.85, 270.75, 269.65, 269.95, 269.65, 
    269.65, 269.55, 269.45, 269.45, 269.55, 269.55, 270.35, 270.95, 270.95, 
    271.35, 272.75, 272.75, 272.85, 273.05, 273.05, 273.55, 273.25, 273.65, 
    273.55, 273.55, 273.25, 273.15, 272.95, 272.85, 272.55, 271.95, 272.45, 
    272.55, 272.55, 272.75, 273.15, 273.35, 274.25, 273.45, 274.75, 274.35, 
    275.55, 274.75, 275.05, 275.85, 275.85, 274.85, 274.15, 273.85, 273.75, 
    273.35, 272.65, 272.15, 270.95, 270.15, 269.65, 269.85, 269.95, 269.55, 
    269.05, 268.75, 269.45, 267.65, 269.05, 268.85, 268.75, 267.35, 267.05, 
    266.25, 268.75, 267.25, 266.85, 268.25, 266.55, 267.05, 266.75, 267.05, 
    266.55, 266.35, 266.15, 266.65, 266.95, 267.25, 267.45, 267.65, 267.15, 
    267.55, 267.05, 267.25, 267.55, 268.25, 267.65, 268.05, 268.55, 268.15, 
    267.45, 267.55, 267.65, 267.65, 266.85, 266.45, 266.15, 265.55, 265.45, 
    265.25, 264.75, 265.25, 265.85, 266.35, 267.95, 267.85, 268.35, 268.25, 
    269.25, 268.75, 269.25, 269.75, 269.05, 269.35, 268.95, 268.55, 268.55, 
    267.65, 267.45, 267.35, 267.45, 267.05, 266.95, 266.75, 266.55, 266.85, 
    266.25, 266.05, 267.45, 267.65, 267.05, 267.15, 267.45, 268.35, 267.75, 
    267.45, 268.05, 268.35, 267.95, 267.65, 267.75, 267.25, 266.95, 266.65, 
    266.65, 266.35, 266.15, 265.85, 266.15, 266.75, 267.35, 267.95, 268.75, 
    268.65, 269.05, 269.15, 269.55, 270.15, 270.55, 270.55, 270.15, 270.35, 
    269.95, 269.95, 268.85, 268.15, 268.35, 267.75, 267.35, 267.15, 266.55, 
    266.75, 266.45, 266.25, 266.95, 266.85, 267.75, 268.35, 268.55, 268.95, 
    269.35, 270.05, 270.15, 269.55, 270.25, 269.65, 269.85, 269.95, 269.65, 
    269.55, 268.75, 269.15, 268.75, 268.55, 268.35, 268.35, 267.75, 268.05, 
    269.05, 269.45, 269.65, 269.75, 269.75, 269.85, 270.65, 270.75, 269.95, 
    269.85, 269.65, 270.35, 270.25, 269.65, 269.45, 268.75, 268.85, 268.55, 
    268.45, 267.85, 267.55, 267.75, 267.75, 268.05, 268.35, 268.35, 268.85, 
    268.65, 269.05, 270.25, 270.35, 270.85, 270.85, 270.95, 272.25, 270.85, 
    271.55, 271.75, 272.95, 271.35, 270.45, 272.35, 271.85, 272.05, 272.55, 
    272.75, 273.25, 273.25, 273.35, 273.95, 273.95, 274.55, 274.55, 274.95, 
    276.15, 277.05, 278.45, 279.05, 280.65, 279.35, 279.25, 279.75, 279.35, 
    278.05, 277.45, 278.45, 278.05, 278.15, 278.75, 278.75, 278.75, 278.35, 
    277.95, 277.25, 277.55, 278.75, 278.65, 278.65, 280.35, 280.15, 279.85, 
    280.55, 278.35, 280.35, 278.55, 277.55, 278.05, 279.25, 278.05, 277.25, 
    275.95, 273.55, 273.75, 273.15, 273.65, 274.25, 274.45, 274.35, 274.75, 
    275.55, 274.45, 275.15, 275.85, 275.05, 275.45, 275.25, 275.35, 275.35, 
    275.25, 275.35, 275.75, 275.95, 275.15, 273.75, 272.95, 272.85, 272.65, 
    272.55, 272.55, 274.25, 274.45, 273.85, 274.75, 274.55, 274.45, 275.05, 
    274.65, 274.65, 274.65, 274.75, 274.75, 274.55, 274.55, 274.65, 274.45, 
    274.25, 274.05, 274.15, 274.25, 274.25, 274.15, 274.25, 273.95, 273.75, 
    273.95, 274.15, 274.35, 274.25, 274.35, 274.25, 274.75, 275.15, 275.05, 
    275.35, 275.35, 275.05, 274.95, 274.75, 274.85, 274.65, 274.65, 274.55, 
    274.35, 274.65, 274.25, 274.35, 274.15, 274.25, 274.25, 274.35, 274.65, 
    274.55, 274.75, 274.85, 274.95, 275.25, 275.45, 275.55, 275.95, 275.55, 
    275.45, 276.05, 275.85, 275.85, 275.75, 274.55, 274.35, 274.15, 273.85, 
    274.05, 274.45, 274.55, 274.15, 273.85, 274.05, 273.65, 274.85, 274.95, 
    275.65, 276.85, 276.65, 278.15, 279.75, 279.05, 279.35, 278.15, 278.75, 
    279.45, 279.75, 277.35, 277.75, 277.25, 276.45, 276.35, 278.15, 279.95, 
    280.45, 280.35, 281.05, 281.65, 279.45, 279.25, 279.45, 278.75, 278.95, 
    279.85, 279.55, 279.25, 277.75, 277.15, 277.95, 277.75, 276.95, 277.05, 
    275.35, 275.75, 275.75, 276.25, 275.45, 275.55, 275.95, 276.15, 276.65, 
    277.45, 278.35, 277.95, 278.55, 278.25, 278.35, 277.85, 278.05, 276.95, 
    276.55, 275.95, 275.65, 275.85, 275.85, 275.55, 275.75, 275.75, 275.45, 
    275.85, 276.15, 275.95, 275.25, 276.35, 276.55, 276.55, 277.05, 277.95, 
    278.15, 278.25, 279.15, 278.85, 279.05, 279.55, 279.95, 279.85, 280.05, 
    280.45, 280.65, 278.15, 277.55, 277.45, 277.35, 276.55, 278.25, 279.25, 
    278.75, 277.35, 277.85, 278.05, 278.45, 278.45, 278.35, 278.75, 278.55, 
    279.15, 278.45, 278.55, 278.15, 278.15, 278.05, 277.95, 277.55, 277.75, 
    277.55, 277.75, 277.25, 277.25, 277.15, 277.55, 277.65, 277.15, 277.55, 
    277.35, 277.45, 277.75, 277.95, 278.25, 278.65, 278.25, 278.35, 279.45, 
    278.65, 280.45, 278.65, 278.55, 278.35, 278.35, 278.55, 278.05, 277.95, 
    277.75, 277.55, 278.05, 277.95, 278.95, 279.75, 280.05, 279.75, 279.75, 
    278.95, 279.25, 280.05, 280.45, 281.15, 280.75, 281.35, 281.25, 280.65, 
    280.75, 280.35, 279.65, 278.95, 278.65, 278.15, 277.75, 278.65, 279.75, 
    279.85, 279.25, 279.25, 277.85, 277.75, 277.15, 277.45, 277.75, 277.75, 
    277.65, 277.75, 278.55, 278.35, 277.85, 277.85, 277.55, 277.45, 277.35, 
    276.75, 276.75, 276.55, 276.95, 276.85, 276.95, 277.45, 277.55, 277.95, 
    277.35, 277.75, 277.55, 277.45, 277.55, 277.25, 277.25, 277.45, 277.35, 
    277.35, 277.05, 277.25, 277.15, 277.15, 277.15, 276.85, 276.75, 276.55, 
    276.75, 276.75, 276.75, 276.75, 277.15, 277.45, 277.95, 278.75, 279.55, 
    278.95, 279.75, 279.75, 279.75, 279.65, 279.15, 278.65, 278.35, 278.15, 
    277.55, 277.45, 277.25, 277.35, 276.85, 276.55, 276.45, 276.25, 276.25, 
    276.55, 276.65, 277.35, 277.55, 277.95, 277.85, 277.75, 277.65, 277.25, 
    277.35, 277.55, 277.65, 277.45, 277.85, 277.65, 277.35, 277.55, 277.35, 
    277.15, 276.85, 276.75, 276.15, 275.65, 275.85, 275.75, 275.55, 275.85, 
    276.15, 276.05, 276.35, 276.45, 276.75, 276.95, 276.95, 277.25, 277.55, 
    277.25, 277.05, 276.85, 276.85, 276.55, 276.45, 276.25, 275.95, 275.75, 
    275.45, 275.15, 275.35, 275.85, 275.95, 276.25, 276.95, 277.45, 278.05, 
    277.55, 277.25, 277.35, 276.95, 277.45, 277.95, 278.35, 277.95, 277.25, 
    277.45, 276.95, 276.75, 276.85, 276.35, 276.55, 276.45, 276.45, 276.75, 
    276.95, 277.15, 277.35, 277.15, 277.35, 277.55, 278.15, 278.15, 278.45, 
    278.45, 278.95, 278.85, 279.75, 279.75, 279.25, 278.75, 279.05, 278.75, 
    278.05, 277.65, 277.85, 278.35, 278.85, 278.65, 278.85, 279.25, 279.05, 
    279.15, 279.15, 279.15, 279.45, 279.75, 280.25, 279.95, 279.55, 279.25, 
    279.25, 279.25, 278.65, 278.85, 278.45, 278.75, 278.85, 278.75, 278.45, 
    277.95, 277.75, 277.65, 277.15, 277.35, 276.95, 276.55, 276.45, 277.15, 
    277.15, 277.75, 278.55, 278.45, 278.35, 278.35, 277.95, 278.35, 278.65, 
    278.25, 278.25, 278.15, 278.15, 278.25, 278.25, 278.15, 278.45, 278.25, 
    277.65, 277.95, 278.75, 279.45, 279.35, 279.05, 279.75, 280.45, 280.15, 
    280.35, 280.85, 280.55, 281.05, 280.55, 280.75, 280.85, 280.35, 279.35, 
    279.85, 279.05, 278.45, 278.35, 278.35, 278.35, 278.15, 278.15, 277.75, 
    277.65, 278.45, 278.15, 277.65, 278.15, 278.55, 278.55, 278.25, 277.95, 
    277.85, 277.85, 277.75, 277.45, 277.45, 277.45, 277.35, 277.05, 276.95, 
    276.75, 276.75, 276.85, 277.15, 277.55, 277.45, 277.75, 278.75, 278.45, 
    278.45, 278.95, 279.25, 280.05, 279.35, 279.45, 279.45, 278.75, 278.85, 
    278.95, 279.05, 279.25, 278.05, 277.25, 277.75, 277.65, 277.15, 277.45, 
    277.75, 277.25, 277.35, 277.95, 278.65, 279.15, 279.35, 279.15, 279.55, 
    279.65, 279.75, 279.85, 279.65, 279.45, 279.65, 279.75, 279.45, 279.25, 
    279.55, 279.15, 278.65, 278.65, 278.65, 278.95, 280.15, 279.25, 279.35, 
    279.65, 280.45, 280.15, 280.35, 281.05, 279.75, 280.25, 280.15, 279.65, 
    278.95, 278.75, 278.35, 278.65, 278.55, 278.55, 278.75, 278.85, 278.75, 
    278.65, 278.55, 278.55, 278.65, 278.65, 279.35, 278.85, 279.15, 278.65, 
    278.45, 278.95, 279.35, 279.55, 279.45, 279.35, 279.25, 278.85, 278.95, 
    278.85, 278.15, 277.95, 277.95, 277.95, 277.65, 277.75, 277.45, 277.55, 
    277.35, 277.75, 277.45, 277.65, 277.85, 278.45, 279.35, 279.65, 279.95, 
    279.75, 279.75, 279.75, 279.15, 278.65, 278.35, 278.25, 278.25, 277.85, 
    277.55, 277.45, 277.35, 277.15, 277.05, 277.35, 277.95, 278.25, 278.95, 
    279.05, 279.25, 279.55, 279.55, 279.45, 279.55, 279.05, 279.65, 280.35, 
    279.85, 280.15, 279.55, 279.45, 279.45, 279.55, 279.35, 279.25, 278.95, 
    278.65, 278.35, 278.25, 278.15, 278.05, 278.55, 278.25, 278.45, 278.85, 
    279.85, 280.65, 280.55, 280.25, 279.65, 280.55, 279.55, 279.35, 278.45, 
    278.05, 277.75, 277.25, 276.95, 276.75, 276.55, 276.65, 276.65, 276.95, 
    276.85, 276.85, 276.95, 277.35, 277.35, 278.15, 278.65, 278.85, 278.75, 
    278.65, 278.35, 278.35, 278.05, 278.35, 277.15, 277.05, 276.75, 276.55, 
    276.65, 276.55, 276.75, 276.95, 277.15, 277.05, 277.35, 277.35, 277.55, 
    278.25, 278.25, 278.45, 278.55, 278.45, 278.75, 279.05, 279.45, 279.45, 
    279.85, 279.45, 279.25, 279.05, 279.05, 278.95, 278.45, 278.05, 277.65, 
    277.75, 277.75, 277.95, 277.95, 278.35, 278.85, 278.65, 278.45, 279.05, 
    279.35, 279.25, 279.25, 279.25, 279.35, 279.05, 278.65, 279.25, 278.65, 
    278.15, 277.85, 277.55, 277.05, 276.85, 276.65, 276.45, 276.45, 277.35, 
    277.25, 277.65, 278.05, 277.85, 278.45, 277.55, 278.15, 277.95, 277.85, 
    278.35, 278.55, 278.35, 278.65, 278.45, 277.95, 277.75, 277.95, 278.05, 
    278.25, 277.95, 277.75, 277.85, 277.75, 278.05, 277.95, 277.95, 278.35, 
    278.55, 278.95, 279.25, 278.95, 279.15, 279.55, 279.35, 279.35, 279.35, 
    278.75, 278.65, 278.55, 278.25, 277.85, 277.85, 277.85, 277.75, 277.55, 
    277.55, 277.65, 277.85, 278.15, 278.35, 278.65, 279.15, 279.45, 279.85, 
    280.45, 280.55, 280.65, 280.65, 281.05, 280.45, 280.55, 280.15, 279.55, 
    279.45, 278.95, 278.55, 278.75, 278.75, 278.85, 278.75, 278.55, 278.95, 
    278.95, 279.35, 279.95, 279.85, 280.05, 279.85, 280.15, 279.95, 278.95, 
    279.45, 279.45, 279.25, 278.95, 278.85, 278.75, 278.65, 278.65, 278.45, 
    278.45, 278.05, 278.45, 278.25, 278.45, 278.35, 278.35, 278.35, 278.55, 
    278.55, 279.45, 279.75, 279.35, 279.25, 279.45, 279.85, 279.75, 279.55, 
    279.55, 279.55, 279.45, 279.45, 279.35, 279.25, 279.25, 279.25, 279.05, 
    279.15, 278.85, 278.75, 278.85, 278.95, 279.45, 279.85, 279.85, 279.65, 
    279.55, 279.55, 279.65, 280.05, 279.95, 280.15, 279.85, 279.55, 279.65, 
    279.55, 279.25, 279.05, 278.25, 278.05, 277.55, 277.25, 277.55, 277.55, 
    277.45, 277.55, 277.55, 278.65, 278.15, 278.65, 278.85, 279.05, 279.55, 
    279.45, 279.75, 279.85, 280.15, 279.95, 280.25, 280.05, 280.05, 279.85, 
    279.55, 279.55, 279.45, 279.65, 279.45, 279.75, 279.55, 279.55, 280.45, 
    280.95, 280.95, 281.25, 281.45, 281.45, 281.85, 282.05, 282.15, 282.25, 
    282.55, 282.45, 281.85, 281.75, 281.65, 280.65, 279.95, 280.05, 280.85, 
    280.45, 280.25, 280.25, 280.55, 280.25, 281.25, 281.25, 281.85, 281.45, 
    281.75, 282.15, 281.95, 281.65, 281.25, 281.25, 281.55, 281.35, 281.05, 
    281.05, 280.75, 280.65, 280.65, 280.25, 280.25, 279.65, 279.45, 280.55, 
    280.15, 280.05, 280.25, 281.05, 282.05, 281.75, 281.85, 282.45, 282.85, 
    282.95, 282.65, 282.35, 281.85, 282.25, 281.65, 281.45, 281.65, 281.55, 
    281.15, 280.75, 280.95, 280.75, 280.45, 280.35, 280.15, 279.85, 279.75, 
    279.65, 279.35, 279.35, 279.35, 279.45, 279.75, 279.85, 280.15, 280.15, 
    279.95, 280.15, 280.45, 280.85, 280.85, 281.35, 281.15, 280.85, 280.55, 
    280.45, 280.35, 280.45, 280.65, 280.85, 281.35, 281.05, 280.75, 280.45, 
    279.95, 279.75, 279.65, 279.75, 279.85, 279.95, 278.95, 279.05, 279.05, 
    279.25, 279.55, 279.55, 279.85, 279.85, 279.75, 279.75, 279.95, 280.15, 
    280.15, 280.25, 280.55, 280.15, 280.95, 280.95, 281.05, 281.05, 281.25, 
    281.15, 281.25, 281.45, 281.65, 281.35, 281.65, 281.55, 281.65, 281.15, 
    281.85, 281.65, 282.55, 282.65, 282.25, 282.65, 282.85, 283.15, 283.35, 
    283.05, 282.65, 282.15, 281.05, 281.05, 280.75, 281.55, 282.95, 281.35, 
    281.85, 281.45, 281.55, 281.55, 281.35, 281.55, 281.65, 281.35, 281.35, 
    281.55, 281.45, 282.35, 283.25, 283.25, 282.65, 282.95, 283.55, 285.65, 
    284.45, 285.35, 284.45, 284.15, 284.05, 284.65, 284.35, 284.55, 284.25, 
    284.95, 284.55, 283.95, 283.65, 283.35, 282.85, 283.15, 282.25, 283.15, 
    282.75, 283.35, 283.05, 283.55, 282.05, 282.55, 282.85, 282.45, 281.85, 
    282.35, 282.45, 282.75, 284.15, 282.75, 282.15, 283.25, 282.95, 282.55, 
    282.05, 281.95, 280.85, 281.25, 281.45, 281.25, 281.25, 280.95, 281.15, 
    281.05, 281.45, 280.65, 281.15, 281.35, 281.05, 280.95, 280.85, 280.85, 
    280.95, 280.95, 281.15, 280.85, 280.05, 279.75, 279.35, 279.15, 279.15, 
    279.45, 279.25, 278.55, 278.85, 278.95, 278.85, 278.75, 279.05, 279.45, 
    280.15, 279.65, 280.15, 279.45, 279.75, 280.25, 280.05, 279.65, 279.95, 
    280.45, 280.75, 280.65, 280.85, 280.85, 280.25, 280.35, 280.45, 280.35, 
    280.15, 280.25, 280.65, 281.25, 281.05, 281.05, 280.95, 280.75, 280.65, 
    280.75, 281.05, 281.05, 281.15, 280.75, 280.85, 280.35, 280.25, 280.15, 
    279.85, 280.05, 280.25, 280.25, 280.15, 280.15, 280.65, 280.35, 280.25, 
    280.05, 280.35, 280.45, 280.65, 281.25, 281.15, 281.15, 281.35, 281.55, 
    281.65, 281.65, 281.95, 281.85, 281.35, 281.45, 281.75, 281.35, 281.25, 
    281.05, 281.15, 281.55, 280.85, 280.45, 280.35, 280.05, 280.35, 280.45, 
    281.65, 281.25, 280.85, 280.55, 281.85, 282.15, 282.85, 282.15, 280.95, 
    280.55, 280.05, 279.65, 279.25, 279.25, 279.05, 278.65, 278.85, 278.85, 
    279.55, 279.95, 279.75, 279.95, 279.75, 280.15, 280.65, 280.75, 281.05, 
    280.85, 281.15, 281.45, 281.15, 281.15, 280.55, 280.65, 280.35, 280.45, 
    280.45, 280.35, 280.15, 280.25, 280.45, 280.45, 279.95, 280.25, 280.15, 
    280.25, 280.35, 280.15, 280.55, 280.65, 280.65, 281.25, 281.25, 281.95, 
    281.95, 282.25, 282.45, 282.75, 281.85, 280.95, 281.65, 281.25, 281.35, 
    280.95, 280.85, 280.55, 280.75, 280.75, 280.95, 281.05, 281.55, 281.75, 
    282.45, 282.55, 282.35, 282.05, 281.85, 281.15, 282.05, 281.55, 281.55, 
    281.15, 280.75, 280.25, 279.95, 279.65, 279.75, 279.55, 279.45, 279.25, 
    279.65, 279.45, 279.35, 279.25, 279.55, 279.75, 279.15, 280.45, 281.05, 
    280.45, 280.55, 281.05, 281.25, 281.35, 281.45, 281.15, 280.75, 280.45, 
    280.05, 280.25, 279.95, 279.85, 279.85, 280.15, 279.85, 279.95, 280.15, 
    279.85, 279.85, 280.55, 280.35, 279.55, 279.95, 279.05, 279.35, 279.45, 
    279.15, 279.55, 279.05, 278.05, 277.95, 278.95, 278.45, 278.35, 278.25, 
    278.05, 277.85, 278.35, 279.15, 278.85, 279.35, 279.15, 279.35, 279.15, 
    279.75, 279.65, 279.65, 280.45, 280.85, 281.05, 281.55, 280.85, 281.25, 
    280.75, 280.55, 280.25, 280.05, 279.75, 279.35, 279.25, 279.15, 279.45, 
    279.55, 279.75, 279.55, 279.35, 280.15, 280.45, 281.05, 280.55, 280.85, 
    281.05, 281.55, 281.75, 281.75, 282.35, 282.15, 281.85, 281.15, 281.35, 
    280.95, 280.45, 280.65, 280.25, 279.65, 279.75, 280.55, 280.15, 280.95, 
    280.95, 280.45, 280.65, 281.25, 281.55, 282.25, 281.95, 281.85, 281.65, 
    281.65, 281.35, 281.45, 281.25, 280.65, 280.35, 280.15, 280.45, 280.45, 
    280.25, 280.15, 280.35, 280.05, 280.05, 279.85, 279.95, 280.15, 279.95, 
    280.05, 280.35, 280.45, 280.65, 280.75, 281.25, 281.05, 281.05, 280.95, 
    281.15, 281.25, 280.65, 279.85, 280.25, 280.15, 280.05, 280.15, 280.65, 
    281.55, 281.15, 282.25, 283.05, 282.95, 282.85, 282.75, 282.35, 282.85, 
    284.05, 283.65, 283.35, 284.65, 284.35, 284.35, 284.15, 283.25, 282.55, 
    282.15, 280.95, 281.05, 280.45, 280.75, 280.65, 281.15, 281.45, 281.55, 
    281.75, 281.95, 282.15, 282.45, 282.45, 282.25, 282.75, 282.85, 282.95, 
    283.45, 283.25, 282.75, 282.05, 282.65, 282.15, 281.25, 281.15, 281.05, 
    280.65, 280.45, 280.55, 280.65, 280.45, 280.45, 280.85, 280.95, 281.05, 
    281.35, 281.35, 281.55, 281.75, 281.35, 281.45, 281.55, 281.75, 281.35, 
    281.05, 281.15, 280.85, 280.55, 280.25, 279.85, 279.65, 279.25, 278.95, 
    279.25, 279.15, 279.35, 279.65, 279.95, 279.75, 279.95, 280.15, 280.15, 
    280.25, 280.45, 280.85, 280.65, 280.55, 280.75, 281.05, 280.95, 281.05, 
    280.95, 280.85, 280.55, 280.45, 280.55, 280.35, 280.15, 280.35, 280.95, 
    280.85, 281.35, 281.45, 281.25, 281.15, 281.45, 281.55, 281.85, 281.85, 
    282.25, 281.85, 281.65, 281.55, 281.45, 281.25, 281.15, 280.95, 280.85, 
    280.65, 280.55, 280.55, 280.75, 280.65, 281.25, 281.05, 280.85, 280.85, 
    280.85, 280.45, 280.75, 281.25, 281.65, 281.75, 281.85, 281.25, 281.35, 
    281.25, 281.05, 280.95, 280.45, 280.25, 280.25, 280.25, 280.25, 280.05, 
    280.05, 280.55, 280.55, 280.75, 281.15, 281.55, 281.55, 281.55, 281.65, 
    281.95, 282.15, 281.85, 282.05, 282.15, 281.95, 281.35, 281.05, 280.65, 
    280.25, 280.05, 279.85, 279.65, 279.55, 279.25, 279.25, 279.25, 279.35, 
    279.45, 279.65, 279.95, 279.75, 279.75, 280.05, 280.05, 280.25, 280.35, 
    280.25, 280.35, 280.55, 280.25, 280.25, 279.55, 279.45, 279.05, 279.75, 
    279.95, 279.55, 279.85, 279.95, 280.25, 280.25, 280.15, 280.05, 280.25, 
    279.95, 279.95, 279.95, 279.95, 280.15, 280.15, 280.05, 280.65, 280.25, 
    280.35, 279.65, 279.95, 280.25, 280.15, 280.55, 280.75, 280.55, 280.75, 
    280.55, 281.05, 281.65, 281.25, 281.75, 281.45, 281.75, 281.55, 281.25, 
    281.65, 281.25, 281.15, 281.15, 280.95, 280.55, 280.25, 279.95, 279.95, 
    280.55, 280.45, 280.05, 279.95, 279.85, 280.05, 280.55, 280.55, 280.85, 
    281.65, 281.45, 281.05, 282.15, 282.05, 281.65, 281.15, 281.85, 280.45, 
    280.75, 281.05, 281.15, 281.35, 281.55, 281.55, 281.15, 280.85, 280.85, 
    281.15, 279.95, 279.95, 280.45, 280.45, 280.45, 280.05, 279.65, 280.15, 
    281.05, 281.55, 281.75, 281.95, 281.45, 281.35, 281.15, 281.55, 281.15, 
    281.25, 281.05, 280.75, 281.35, 280.65, 280.25, 279.95, 279.45, 279.75, 
    279.95, 280.05, 280.35, 280.85, 280.75, 281.05, 280.35, 280.65, 279.95, 
    280.45, 280.55, 280.45, 280.45, 280.35, 280.15, 279.75, 280.15, 280.15, 
    280.05, 279.85, 279.75, 279.35, 279.15, 279.15, 279.05, 278.55, 278.25, 
    278.35, 278.55, 278.45, 278.65, 278.45, 278.35, 278.55, 278.75, 278.95, 
    279.55, 279.55, 279.55, 279.35, 279.35, 279.05, 279.05, 278.95, 278.85, 
    278.75, 278.75, 278.85, 278.85, 278.35, 278.05, 277.85, 278.15, 278.85, 
    279.75, 280.45, 281.25, 280.65, 280.25, 279.55, 279.25, 278.95, 277.95, 
    277.55, 277.35, 276.85, 276.15, 275.75, 275.25, 275.25, 275.15, 275.05, 
    275.65, 275.95, 276.25, 276.45, 276.85, 277.45, 277.65, 277.55, 277.65, 
    278.05, 278.05, 277.65, 277.15, 276.95, 276.65, 276.45, 276.25, 276.15, 
    276.05, 275.85, 275.75, 275.75, 275.95, 276.05, 276.25, 276.35, 276.45, 
    276.65, 276.55, 276.85, 277.75, 278.15, 277.55, 278.45, 278.15, 277.95, 
    278.45, 278.85, 278.75, 278.45, 278.05, 277.55, 277.15, 276.75, 276.05, 
    276.05, 275.75, 274.95, 274.45, 275.65, 276.45, 277.15, 277.35, 277.25, 
    277.65, 277.85, 277.75, 278.05, 278.25, 278.95, 278.65, 278.55, 278.45, 
    278.25, 278.05, 277.65, 277.55, 277.25, 276.55, 276.75, 276.65, 276.55, 
    276.55, 276.75, 277.35, 277.65, 277.95, 278.65, 278.25, 278.15, 278.45, 
    279.25, 278.65, 278.55, 278.85, 279.05, 278.55, 278.45, 277.75, 277.65, 
    277.45, 276.75, 276.45, 275.65, 275.45, 275.65, 276.35, 277.05, 277.25, 
    277.45, 278.65, 278.25, 278.55, 278.75, 279.25, 279.95, 279.85, 280.15, 
    280.55, 280.35, 280.75, 280.85, 280.15, 279.75, 279.25, 279.45, 279.05, 
    278.95, 278.65, 278.25, 278.25, 278.55, 278.25, 278.05, 277.85, 278.45, 
    278.05, 278.45, 278.65, 278.85, 278.85, 279.15, 279.15, 279.55, 279.35, 
    278.75, 278.25, 277.45, 276.75, 276.55, 276.15, 276.35, 276.95, 277.15, 
    277.35, 277.55, 277.95, 278.35, 278.55, 278.95, 278.95, 278.75, 278.95, 
    279.05, 279.15, 279.55, 279.35, 279.25, 278.95, 278.65, 278.65, 278.35, 
    278.15, 278.05, 277.95, 277.85, 277.95, 277.85, 278.15, 277.45, 277.85, 
    277.85, 278.05, 278.05, 278.65, 278.85, 278.75, 279.15, 279.75, 279.45, 
    278.75, 279.15, 279.05, 279.45, 279.45, 278.85, 278.85, 279.05, 279.85, 
    279.55, 279.65, 279.25, 279.25, 279.45, 279.65, 279.65, 280.05, 280.65, 
    280.05, 279.95, 280.05, 279.95, 279.95, 280.85, 280.35, 280.55, 279.75, 
    279.25, 279.25, 279.15, 278.75, 278.35, 278.05, 277.95, 277.75, 277.75, 
    277.25, 277.65, 277.65, 277.75, 278.15, 278.25, 278.55, 279.15, 278.85, 
    278.45, 278.45, 278.05, 277.75, 277.25, 277.05, 276.55, 276.35, 276.15, 
    275.05, 274.95, 274.25, 274.65, 274.35, 274.25, 274.55, 274.85, 275.35, 
    275.45, 275.45, 275.15, 276.05, 276.85, 277.35, 276.85, 276.85, 277.55, 
    277.45, 277.25, 277.25, 277.25, 277.05, 276.35, 275.95, 276.15, 275.85, 
    275.45, 275.35, 275.55, 275.35, 275.25, 276.15, 276.55, 276.85, 277.25, 
    277.65, 278.45, 278.75, 278.85, 278.75, 278.55, 278.35, 278.55, 278.55, 
    278.45, 278.55, 278.15, 278.15, 278.05, 277.95, 277.35, 277.45, 277.75, 
    277.95, 277.85, 278.15, 278.85, 279.25, 279.55, 279.35, 279.85, 280.25, 
    281.25, 281.75, 281.65, 281.35, 281.05, 281.45, 281.65, 281.55, 281.65, 
    280.45, 280.65, 279.65, 279.75, 279.25, 279.05, 278.65, 278.65, 278.35, 
    278.45, 278.15, 278.15, 277.85, 277.85, 277.45, 276.65, 276.75, 276.55, 
    276.45, 276.35, 276.05, 275.65, 275.65, 275.45, 274.65, 274.45, 273.95, 
    273.85, 273.45, 273.15, 273.15, 272.95, 272.95, 273.35, 273.55, 273.95, 
    274.45, 274.05, 273.85, 274.25, 274.45, 274.15, 274.25, 273.95, 273.95, 
    272.95, 272.95, 272.35, 271.85, 271.65, 271.35, 271.25, 271.45, 272.15, 
    272.55, 272.95, 273.75, 274.45, 274.25, 274.65, 274.85, 275.15, 275.45, 
    275.85, 275.95, 276.15, 276.05, 276.05, 275.85, 275.85, 275.85, 275.85, 
    275.85, 275.65, 275.85, 275.85, 275.85, 275.95, 276.35, 276.85, 277.15, 
    277.25, 278.05, 278.15, 278.85, 279.45, 279.35, 278.35, 278.85, 279.15, 
    279.45, 279.75, 279.35, 279.75, 280.15, 279.95, 279.85, 279.85, 279.55, 
    279.45, 279.45, 279.95, 279.85, 278.75, 279.25, 279.75, 280.05, 280.25, 
    280.25, 280.85, 281.35, 282.05, 282.15, 282.55, 281.55, 281.05, 281.45, 
    280.55, 279.85, 279.55, 279.15, 278.25, 277.75, 277.75, 277.55, 277.45, 
    277.35, 277.25, 277.15, 277.45, 277.45, 277.55, 277.55, 277.75, 278.15, 
    278.65, 278.05, 278.35, 278.55, 278.25, 277.75, 277.15, 276.35, 276.35, 
    275.65, 275.05, 275.25, 275.05, 275.55, 275.25, 274.95, 276.15, 276.15, 
    276.45, 276.85, 276.95, 276.95, 277.45, 277.65, 279.25, 279.85, 281.05, 
    278.45, 278.85, 279.25, 277.55, 277.35, 277.15, 277.05, 276.55, 277.05, 
    276.25, 276.65, 276.45, 276.55, 276.65, 277.05, 277.35, 277.55, 277.55, 
    279.15, 279.25, 279.85, 280.65, 281.55, 281.55, 281.05, 280.25, 280.45, 
    280.05, 280.25, 279.45, 278.95, 279.25, 279.65, 278.75, 278.15, 278.45, 
    280.35, 279.25, 280.05, 280.05, 279.45, 279.85, 279.65, 280.35, 280.45, 
    279.85, 279.85, 279.75, 280.45, 280.55, 280.25, 280.15, 280.15, 280.05, 
    279.75, 279.45, 278.75, 278.55, 278.55, 278.65, 278.75, 278.55, 278.65, 
    278.75, 278.85, 279.15, 280.15, 279.45, 279.55, 279.95, 279.95, 280.35, 
    280.45, 280.45, 279.15, 279.25, 280.05, 279.15, 279.35, 278.45, 277.85, 
    278.25, 277.85, 277.95, 277.85, 277.75, 277.05, 277.85, 278.15, 278.25, 
    277.95, 277.75, 277.85, 277.75, 278.05, 278.15, 278.05, 277.95, 277.45, 
    276.55, 275.75, 275.75, 275.35, 275.55, 275.45, 275.35, 275.35, 275.35, 
    276.55, 275.45, 276.75, 277.35, 277.35, 278.55, 278.55, 279.65, 280.15, 
    280.75, 280.25, 280.55, 279.95, 279.45, 278.95, 278.55, 278.95, 278.45, 
    279.05, 278.85, 279.45, 279.25, 279.15, 279.25, 279.05, 279.05, 279.45, 
    280.15, 279.85, 279.85, 279.95, 280.85, 280.95, 281.05, 280.75, 280.15, 
    279.65, 279.25, 279.15, 278.85, 278.75, 278.95, 278.75, 278.45, 278.65, 
    278.55, 278.75, 278.65, 278.75, 278.85, 278.75, 279.05, 278.95, 279.25, 
    279.45, 279.15, 279.15, 279.05, 278.65, 278.35, 278.75, 278.55, 278.55, 
    278.25, 278.25, 277.75, 277.55, 277.65, 277.35, 277.05, 277.15, 276.85, 
    276.75, 276.75, 277.05, 276.95, 277.65, 277.55, 277.85, 278.35, 277.95, 
    278.35, 278.05, 278.05, 277.95, 277.65, 277.55, 277.15, 277.55, 277.95, 
    277.85, 277.45, 277.25, 277.45, 277.35, 277.05, 276.95, 277.35, 277.25, 
    277.55, 277.75, 277.65, 277.65, 278.15, 278.05, 277.65, 278.15, 277.75, 
    277.35, 276.15, 274.85, 274.45, 273.85, 274.85, 274.35, 274.45, 273.85, 
    274.85, 273.55, 273.85, 274.35, 273.55, 273.95, 274.75, 274.65, 274.95, 
    276.35, 276.25, 276.35, 276.75, 276.95, 276.45, 275.45, 274.85, 274.15, 
    273.75, 273.15, 272.85, 272.85, 272.45, 272.45, 272.75, 273.25, 273.45, 
    273.45, 273.55, 273.75, 273.75, 273.95, 274.25, 274.65, 274.15, 274.15, 
    274.15, 274.15, 274.15, 273.55, 273.25, 273.15, 273.15, 273.25, 273.35, 
    273.75, 273.95, 273.95, 274.65, 274.85, 274.65, 274.95, 275.65, 275.45, 
    275.35, 275.95, 276.55, 276.55, 277.55, 277.65, 277.75, 277.25, 277.25, 
    276.55, 275.55, 274.45, 274.95, 274.95, 274.75, 275.15, 274.65, 274.15, 
    274.75, 274.85, 275.05, 275.05, 275.25, 275.55, 275.75, 275.95, 276.45, 
    279.35, 279.25, 278.25, 279.75, 278.25, 278.15, 280.55, 282.55, 282.65, 
    282.35, 282.35, 281.85, 281.05, 281.35, 281.25, 281.35, 281.35, 281.55, 
    281.05, 280.85, 280.55, 280.95, 280.65, 279.65, 278.65, 277.15, 276.65, 
    276.25, 275.85, 275.45, 274.95, 274.95, 274.95, 274.45, 274.35, 274.25, 
    274.15, 273.95, 273.75, 273.35, 273.65, 273.35, 273.15, 273.05, 273.25, 
    273.45, 273.45, 273.85, 273.75, 273.95, 273.95, 274.05, 274.05, 274.05, 
    274.05, 274.05, 274.05, 273.85, 273.85, 273.75, 273.65, 273.75, 273.45, 
    273.35, 273.35, 273.35, 273.55, 273.35, 273.55, 273.85, 274.25, 274.65, 
    274.85, 274.95, 275.05, 275.15, 275.05, 275.05, 275.15, 275.05, 274.95, 
    275.05, 274.85, 274.85, 274.65, 274.75, 274.85, 274.55, 274.75, 274.45, 
    274.55, 274.65, 274.25, 274.55, 274.45, 274.85, 275.15, 275.05, 275.25, 
    275.15, 275.05, 275.35, 275.05, 275.15, 275.25, 275.25, 275.25, 275.15, 
    275.25, 275.05, 275.35, 275.15, 275.25, 275.35, 275.45, 275.95, 275.75, 
    275.55, 276.55, 276.05, 276.45, 279.85, 279.75, 280.25, 280.05, 279.55, 
    279.65, 279.55, 279.45, 279.25, 278.75, 278.45, 278.65, 278.65, 278.25, 
    277.55, 277.55, 277.85, 277.45, 277.25, 276.65, 276.75, 276.75, 276.85, 
    276.75, 277.35, 277.25, 277.05, 276.95, 276.85, 276.75, 276.25, 275.75, 
    276.05, 276.05, 276.05, 276.55, 276.55, 276.75, 276.45, 276.65, 277.05, 
    276.85, 276.75, 276.35, 276.65, 276.75, 277.05, 277.65, 277.75, 279.85, 
    280.75, 280.85, 279.45, 279.65, 279.85, 279.25, 282.35, 282.35, 282.25, 
    281.95, 281.25, 280.85, 280.15, 280.45, 280.35, 279.95, 279.85, 279.85, 
    279.85, 280.05, 279.95, 280.05, 280.05, 279.85, 279.75, 279.25, 279.25, 
    279.15, 279.15, 278.85, 278.85, 278.95, 278.75, 278.35, 278.25, 278.15, 
    278.15, 277.95, 278.25, 278.45, 278.15, 278.15, 278.15, 278.25, 278.45, 
    278.65, 278.55, 278.75, 279.95, 279.65, 279.25, 278.65, 278.75, 278.45, 
    277.85, 277.85, 278.45, 279.25, 280.25, 279.95, 280.05, 280.45, 280.35, 
    280.45, 281.05, 281.05, 281.05, 279.65, 279.85, 280.85, 281.35, 280.65, 
    280.65, 280.75, 281.25, 281.65, 280.95, 281.55, 280.45, 280.45, 280.25, 
    280.65, 279.65, 279.35, 279.75, 280.75, 280.35, 280.15, 278.75, 278.65, 
    279.25, 278.85, 278.35, 278.45, 278.85, 279.05, 277.85, 278.05, 277.75, 
    277.75, 278.05, 277.95, 277.75, 277.95, 278.35, 278.65, 277.65, 277.85, 
    277.85, 277.55, 277.45, 277.85, 277.75, 277.55, 277.65, 277.55, 277.85, 
    278.55, 277.95, 278.55, 279.25, 278.35, 278.45, 278.45, 279.35, 279.05, 
    278.85, 279.95, 278.05, 278.85, 277.95, 278.55, 277.25, 277.35, 277.75, 
    276.15, 277.05, 277.45, 275.25, 275.95, 276.85, 276.45, 276.05, 276.45, 
    276.65, 276.55, 273.65, 276.05, 273.65, 275.65, 276.25, 275.65, 275.25, 
    275.35, 275.95, 275.25, 274.65, 274.35, 274.25, 273.55, 273.95, 274.05, 
    274.05, 275.25, 274.65, 274.55, 274.25, 274.65, 275.25, 275.45, 274.65, 
    273.85, 273.95, 273.85, 273.85, 274.25, 273.85, 273.65, 273.05, 274.25, 
    273.35, 274.35, 273.25, 273.05, 272.85, 273.35, 273.95, 275.05, 274.15, 
    274.45, 275.25, 274.95, 274.45, 274.55, 274.55, 274.15, 274.25, 275.05, 
    274.85, 275.85, 275.05, 274.75, 274.45, 273.95, 273.75, 273.75, 273.55, 
    273.35, 273.05, 272.75, 273.35, 273.45, 274.15, 274.55, 275.15, 274.95, 
    274.85, 274.75, 274.75, 274.35, 275.05, 275.15, 274.85, 274.75, 274.65, 
    274.85, 274.65, 274.55, 274.65, 273.85, 273.55, 273.35, 273.45, 274.15, 
    274.25, 274.25, 274.15, 274.15, 274.25, 274.35, 274.45, 274.25, 274.45, 
    274.25, 273.95, 274.15, 273.95, 273.65, 273.65, 273.55, 273.35, 273.25, 
    273.45, 273.55, 272.85, 272.55, 272.55, 272.55, 273.35, 273.45, 274.15, 
    274.55, 275.15, 273.35, 273.85, 273.85, 273.85, 272.85, 273.05, 272.85, 
    271.75, 271.45, 271.45, 270.85, 269.65, 270.05, 269.45, 269.95, 269.95, 
    269.35, 270.15, 269.75, 268.75, 269.55, 269.85, 270.45, 270.85, 270.85, 
    270.95, 270.95, 270.45, 270.75, 269.75, 269.75, 270.15, 270.55, 270.85, 
    270.65, 270.75, 270.95, 270.75, 270.65, 270.75, 270.45, 270.65, 270.35, 
    270.35, 270.25, 270.25, 270.35, 270.45, 270.65, 270.65, 270.55, 270.95, 
    270.95, 271.05, 271.25, 271.55, 271.75, 271.95, 272.05, 272.25, 272.55, 
    272.55, 272.65, 272.85, 273.05, 273.05, 273.15, 273.35, 273.65, 273.45, 
    273.65, 274.15, 274.35, 274.55, 274.15, 274.45, 273.95, 273.95, 274.05, 
    273.95, 273.55, 273.65, 273.65, 273.85, 274.05, 274.05, 273.65, 273.25, 
    273.85, 273.45, 273.95, 274.25, 275.05, 274.65, 274.65, 274.05, 273.85, 
    274.25, 274.15, 274.15, 274.55, 274.45, 274.25, 274.45, 274.45, 274.45, 
    274.75, 274.45, 273.95, 274.15, 273.95, 272.75, 272.65, 273.55, 273.65, 
    273.75, 273.75, 273.15, 273.25, 272.95, 272.45, 272.25, 270.65, 270.65, 
    269.55, 269.55, 270.05, 270.35, 270.35, 270.25, 270.35, 270.45, 270.55, 
    269.25, 269.95, 271.75, 270.95, 272.25, 270.55, 270.65, 271.05, 272.75, 
    270.75, 272.15, 273.75, 271.95, 271.55, 271.65, 271.65, 273.45, 272.35, 
    275.05, 275.45, 276.65, 276.95, 277.35, 277.85, 276.95, 277.05, 277.05, 
    277.55, 277.75, 277.65, 277.45, 277.45, 277.15, 277.15, 277.35, 277.55, 
    277.75, 277.65, 278.05, 278.65, 278.45, 278.65, 278.55, 278.45, 278.85, 
    278.65, 278.75, 278.75, 278.55, 278.85, 278.65, 278.55, 278.25, 278.55, 
    278.75, 278.05, 278.25, 277.65, 277.15, 277.15, 276.95, 277.35, 277.45, 
    277.55, 277.35, 277.25, 277.65, 277.75, 277.75, 278.05, 278.05, 277.95, 
    278.25, 277.85, 277.85, 277.95, 277.85, 277.85, 277.95, 277.95, 277.85, 
    277.45, 277.55, 277.95, 277.75, 277.75, 277.65, 277.65, 278.05, 277.65, 
    277.95, 277.85, 277.65, 277.65, 277.75, 277.45, 277.85, 277.25, 277.65, 
    277.25, 277.25, 277.55, 277.35, 277.35, 277.05, 277.35, 277.55, 277.05, 
    277.55, 277.65, 277.35, 277.15, 276.95, 277.05, 277.15, 277.35, 276.95, 
    277.65, 278.25, 277.45, 277.45, 276.85, 276.75, 276.55, 276.85, 276.35, 
    275.95, 275.15, 274.85, 275.25, 275.15, 275.25, 275.55, 275.25, 275.35, 
    275.25, 275.75, 275.65, 274.85, 274.45, 274.35, 273.85, 275.15, 275.05, 
    274.85, 274.55, 274.25, 274.25, 274.15, 273.65, 273.65, 273.45, 273.35, 
    273.15, 273.15, 273.15, 273.15, 272.85, 272.75, 272.35, 272.35, 272.45, 
    272.65, 272.55, 272.15, 271.75, 272.15, 271.85, 271.75, 271.25, 271.25, 
    270.75, 270.85, 270.65, 271.05, 271.35, 271.65, 271.75, 272.05, 272.15, 
    272.15, 272.15, 272.35, 272.55, 272.55, 272.55, 272.75, 272.65, 272.95, 
    273.35, 273.05, 273.35, 273.55, 273.15, 273.15, 273.25, 273.05, 273.75, 
    273.65, 273.75, 273.75, 273.75, 273.85, 274.35, 274.25, 273.65, 273.75, 
    274.05, 273.75, 273.75, 273.55, 273.35, 273.85, 274.15, 273.35, 273.25, 
    273.75, 273.65, 273.45, 273.15, 272.85, 272.65, 272.95, 273.15, 273.05, 
    273.35, 272.95, 273.25, 273.25, 273.35, 273.05, 272.85, 272.95, 272.85, 
    272.95, 272.95, 272.65, 272.95, 273.35, 272.85, 272.85, 272.15, 271.65, 
    272.45, 272.95, 272.95, 272.85, 272.95, 273.25, 273.05, 273.35, 273.35, 
    273.55, 273.85, 274.75, 275.45, 275.65, 276.55, 277.15, 277.75, 277.85, 
    277.65, 277.45, 277.65, 278.65, 278.45, 278.55, 278.65, 278.75, 278.45, 
    278.45, 278.75, 279.35, 279.25, 278.55, 278.25, 278.25, 277.95, 277.15, 
    275.75, 274.45, 274.15, 273.65, 272.95, 272.45, 272.05, 272.05, 271.55, 
    271.15, 270.95, 270.65, 270.35, 270.25, 270.25, 269.95, 269.65, 269.35, 
    269.15, 269.05, 269.25, 269.15, 268.75, 268.45, 268.55, 268.75, 268.65, 
    268.55, 268.45, 268.25, 267.65, 267.45, 267.65, 267.45, 267.55, 267.45, 
    267.05, 266.75, 266.55, 266.25, 266.15, 266.35, 266.35, 266.15, 266.55, 
    266.65, 266.85, 266.95, 267.25, 267.25, 267.05, 266.95, 267.25, 267.65, 
    267.75, 267.85, 268.05, 268.25, 268.35, 268.45, 268.55, 268.65, 268.75, 
    268.95, 269.15, 269.45, 269.55, 269.75, 270.15, 270.15, 269.95, 270.05, 
    270.35, 270.65, 270.75, 272.65, 272.55, 272.55, 272.85, 273.05, 273.25, 
    273.55, 273.95, 274.25, 273.75, 273.55, 272.85, 272.95, 272.95, 272.45, 
    272.15, 271.85, 271.95, 271.95, 271.75, 271.55, 271.15, 270.95, 270.85, 
    270.45, 270.05, 269.55, 269.35, 269.75, 269.75, 269.45, 269.35, 269.05, 
    268.85, 268.65, 268.35, 268.25, 267.95, 268.25, 269.55, 269.15, 268.75, 
    268.05, 267.65, 267.75, 268.05, 268.25, 268.25, 268.35, 268.35, 268.65, 
    268.65, 268.55, 268.05, 268.45, 268.05, 267.75, 267.45, 267.35, 267.45, 
    267.35, 267.25, 267.45, 267.55, 267.85, 268.45, 268.65, 268.75, 268.75, 
    268.65, 268.45, 269.05, 268.65, 269.05, 268.75, 269.15, 269.45, 269.65, 
    269.85, 270.05, 270.55, 270.65, 271.05, 271.35, 271.45, 271.55, 271.45, 
    271.35, 271.25, 271.75, 271.35, 271.85, 272.05, 271.75, 271.25, 271.25, 
    271.35, 271.05, 270.85, 271.15, 271.25, 271.05, 271.45, 271.25, 270.75, 
    270.85, 270.65, 269.85, 270.25, 268.95, 268.65, 268.05, 268.25, 268.15, 
    268.15, 268.25, 268.45, 268.45, 267.15, 267.45, 268.15, 268.25, 268.15, 
    267.85, 267.75, 268.15, 267.85, 267.65, 268.25, 267.65, 267.75, 267.95, 
    268.15, 268.35, 268.45, 268.25, 268.35, 267.85, 267.45, 267.85, 268.05, 
    267.75, 267.25, 267.65, 267.65, 267.85, 267.95, 268.75, 268.95, 269.45, 
    271.05, 271.45, 270.95, 271.25, 271.55, 271.35, 271.25, 271.45, 271.65, 
    271.65, 271.65, 271.65, 272.05, 272.05, 271.65, 271.55, 271.75, 272.35, 
    271.65, 271.95, 272.25, 271.65, 271.95, 272.05, 272.45, 272.25, 272.45, 
    272.95, 272.85, 273.15, 272.95, 272.85, 272.45, 272.25, 271.95, 271.75, 
    272.15, 272.35, 272.55, 272.75, 272.95, 272.85, 273.15, 273.05, 273.25, 
    273.65, 273.45, 273.35, 273.95, 274.15, 274.45, 274.45, 274.95, 275.85, 
    274.65, 274.25, 274.25, 273.85, 273.25, 273.05, 272.45, 271.95, 271.95, 
    271.45, 271.35, 271.15, 271.15, 271.35, 271.35, 270.85, 270.95, 271.05, 
    271.25, 271.55, 271.65, 271.85, 272.25, 272.05, 272.55, 272.15, 271.95, 
    272.05, 272.05, 272.25, 271.85, 272.05, 272.15, 271.95, 271.85, 271.65, 
    271.35, 270.95, 271.05, 270.65, 270.75, 270.35, 270.45, 271.15, 270.75, 
    270.25, 270.45, 270.15, 270.35, 269.65, 269.15, 268.25, 269.85, 269.95, 
    270.05, 269.45, 269.75, 269.55, 270.25, 269.95, 269.95, 269.95, 269.45, 
    267.65, 266.95, 266.15, 266.05, 266.75, 266.45, 266.55, 265.75, 265.65, 
    265.45, 265.65, 265.75, 265.65, 265.35, 265.25, 265.65, 265.55, 266.25, 
    266.35, 266.75, 266.55, 266.55, 269.15, 269.45, 269.85, 270.05, 269.75, 
    270.25, 270.65, 271.15, 271.55, 271.45, 271.25, 271.65, 271.35, 271.55, 
    272.25, 272.05, 272.05, 272.25, 272.25, 272.25, 272.65, 272.45, 272.05, 
    272.05, 271.35, 270.45, 270.45, 270.35, 269.75, 269.65, 269.75, 269.95, 
    270.05, 270.65, 271.15, 271.45, 271.75, 272.15, 272.35, 272.95, 273.35, 
    273.45, 273.25, 273.75, 273.45, 273.65, 273.75, 274.05, 273.95, 274.15, 
    274.05, 274.35, 274.65, 275.25, 274.55, 273.55, 272.55, 272.05, 271.65, 
    271.95, 272.65, 272.75, 273.05, 272.75, 272.05, 271.95, 272.35, 272.25, 
    272.25, 272.35, 272.35, 272.25, 272.25, 272.25, 271.95, 271.85, 271.95, 
    271.45, 271.85, 271.95, 272.05, 271.75, 271.85, 272.35, 272.85, 272.85, 
    273.05, 273.35, 273.15, 273.35, 273.45, 273.45, 273.75, 274.15, 274.15, 
    274.25, 274.35, 274.45, 274.35, 274.25, 274.15, 274.25, 274.55, 274.65, 
    274.75, 274.85, 275.05, 275.05, 275.25, 274.95, 274.85, 273.95, 274.85, 
    274.55, 273.55, 273.05, 272.55, 272.55, 272.85, 273.15, 273.45, 273.45, 
    272.65, 273.25, 272.55, 272.95, 273.15, 272.65, 272.05, 272.25, 272.85, 
    273.05, 273.35, 273.35, 272.85, 272.55, 272.65, 272.35, 271.95, 272.35, 
    272.85, 273.25, 273.05, 272.95, 272.95, 272.65, 272.65, 272.95, 273.15, 
    272.85, 273.15, 272.35, 272.95, 273.25, 272.75, 272.95, 273.25, 272.85, 
    272.45, 272.35, 273.05, 272.95, 272.55, 273.55, 273.55, 273.55, 273.55, 
    273.75, 274.15, 273.65, 274.25, 275.85, 275.65, 275.95, 275.65, 275.35, 
    275.65, 275.75, 275.65, 275.25, 275.35, 275.25, 274.85, 274.95, 274.85, 
    274.65, 273.75, 274.15, 274.65, 274.85, 274.75, 274.35, 274.15, 273.95, 
    274.15, 274.05, 273.75, 273.55, 272.65, 272.35, 272.45, 272.25, 271.75, 
    271.35, 270.85, 270.95, 270.95, 271.05, 271.35, 271.45, 271.25, 270.95, 
    270.75, 270.65, 270.45, 270.05, 270.05, 270.05, 269.85, 269.95, 269.55, 
    269.55, 269.15, 269.25, 269.05, 268.75, 268.85, 269.25, 269.65, 269.85, 
    270.05, 269.95, 270.35, 270.65, 270.75, 271.15, 271.05, 271.25, 270.85, 
    271.25, 271.15, 271.05, 271.25, 271.15, 271.65, 271.65, 271.85, 272.35, 
    271.65, 271.55, 271.25, 271.15, 270.95, 270.85, 270.45, 270.25, 269.95, 
    269.65, 269.15, 269.35, 269.55, 269.55, 269.65, 269.55, 269.55, 269.15, 
    269.05, 268.75, 268.45, 268.15, 268.35, 268.25, 268.35, 268.15, 268.35, 
    268.25, 268.25, 268.35, 268.25, 268.25, 268.25, 268.25, 267.95, 268.15, 
    268.35, 268.35, 269.05, 269.05, 269.05, 268.95, 269.25, 269.35, 269.55, 
    269.25, 269.15, 269.35, 269.65, 269.45, 269.75, 269.55, 269.95, 270.05, 
    270.25, 270.25, 270.15, 270.15, 269.75, 269.65, 269.55, 269.35, 269.25, 
    269.35, 269.05, 268.85, 268.55, 268.55, 268.75, 269.05, 269.25, 269.45, 
    269.25, 268.75, 268.35, 268.45, 268.25, 268.35, 267.75, 267.35, 267.45, 
    267.85, 267.95, 268.55, 268.55, 268.75, 268.75, 268.85, 268.95, 268.55, 
    268.85, 268.65, 268.65, 268.75, 268.75, 269.15, 269.05, 269.25, 269.25, 
    269.15, 269.25, 269.35, 269.15, 269.35, 269.35, 269.15, 268.65, 268.55, 
    269.05, 269.25, 268.85, 268.75, 268.75, 268.55, 268.75, 269.15, 268.95, 
    268.95, 268.95, 269.25, 269.15, 269.35, 269.15, 269.05, 269.05, 269.15, 
    268.95, 269.25, 269.15, 268.75, 268.85, 268.85, 268.75, 268.85, 268.75, 
    268.65, 268.55, 268.45, 268.75, 268.65, 267.95, 268.05, 267.85, 267.85, 
    267.95, 267.55, 267.45, 267.15, 267.15, 266.95, 267.15, 266.95, 266.75, 
    266.85, 266.85, 266.95, 266.85, 266.95, 263.95, 264.45, 264.25, 264.55, 
    264.85, 263.95, 263.85, 264.45, 264.45, 264.05, 263.35, 263.65, 264.05, 
    263.85, 262.75, 263.95, 263.65, 263.45, 264.15, 264.35, 262.65, 263.45, 
    263.55, 264.25, 264.25, 264.05, 263.95, 263.55, 263.35, 262.65, 263.05, 
    263.45, 264.05, 264.15, 264.75, 264.15, 264.95, 265.45, 264.45, 264.65, 
    264.85, 264.65, 264.65, 264.45, 264.45, 264.75, 264.35, 264.85, 264.65, 
    265.05, 265.25, 265.35, 265.75, 265.75, 265.65, 265.65, 266.65, 266.95, 
    268.65, 267.55, 267.25, 266.95, 266.65, 266.05, 265.65, 265.25, 265.05, 
    265.05, 264.55, 264.25, 263.65, 263.55, 262.95, 262.75, 262.75, 262.65, 
    262.35, 263.65, 263.95, 264.15, 264.05, 263.15, 262.35, 260.85, 261.25, 
    261.15, 261.85, 261.45, 262.35, 262.05, 262.15, 262.15, 264.15, 264.05, 
    265.25, 268.65, 268.25, 267.75, 267.65, 267.15, 264.25, 262.75, 263.75, 
    265.55, 265.75, 265.45, 265.35, 263.65, 264.55, 264.25, 262.45, 262.35, 
    261.95, 261.75, 261.55, 261.45, 261.25, 261.35, 261.65, 261.75, 262.15, 
    262.55, 262.45, 262.65, 262.75, 263.35, 263.05, 262.95, 263.15, 263.25, 
    263.65, 264.15, 263.65, 263.55, 264.65, 266.05, 266.25, 266.55, 267.85, 
    268.75, 268.85, 269.35, 269.65, 269.55, 268.65, 268.45, 268.05, 269.75, 
    270.15, 271.05, 271.35, 271.95, 271.85, 272.05, 272.15, 270.65, 269.95, 
    269.65, 269.35, 268.85, 268.35, 267.85, 266.55, 266.25, 265.25, 264.55, 
    265.35, 265.55, 266.35, 265.75, 266.05, 266.15, 265.95, 267.55, 268.65, 
    269.75, 269.65, 269.85, 269.55, 269.55, 269.95, 269.85, 269.45, 269.35, 
    269.15, 269.95, 269.35, 269.05, 269.25, 268.85, 268.75, 268.85, 268.85, 
    269.25, 268.35, 266.95, 265.25, 265.65, 266.25, 266.55, 266.95, 267.45, 
    268.05, 268.95, 271.05, 273.05, 273.45, 273.85, 273.65, 273.65, 273.95, 
    273.85, 274.25, 274.35, 274.35, 273.65, 273.45, 273.55, 273.45, 273.35, 
    273.55, 273.25, 272.75, 273.05, 273.05, 272.85, 272.65, 272.55, 272.55, 
    272.55, 272.55, 272.65, 273.15, 272.85, 273.15, 272.85, 272.95, 272.65, 
    272.25, 271.95, 271.95, 271.85, 271.85, 271.85, 271.25, 270.65, 269.75, 
    268.85, 267.35, 267.65, 268.85, 268.85, 266.45, 266.85, 267.85, 267.85, 
    267.85, 268.45, 268.65, 269.05, 269.15, 269.65, 269.25, 269.15, 268.65, 
    268.95, 269.05, 268.75, 268.25, 268.35, 269.15, 269.45, 269.95, 270.05, 
    270.15, 270.25, 270.45, 270.55, 271.15, 271.05, 271.25, 271.25, 271.05, 
    270.85, 270.65, 270.45, 270.35, 270.35, 270.15, 270.25, 269.95, 270.25, 
    270.55, 269.95, 269.65, 269.55, 269.05, 269.15, 269.05, 268.85, 268.95, 
    268.85, 268.95, 268.85, 268.95, 268.95, 268.85, 269.55, 269.75, 270.45, 
    270.75, 271.15, 271.55, 272.25, 271.85, 271.55, 271.05, 270.85, 270.55, 
    270.35, 270.35, 270.35, 270.15, 270.15, 270.45, 270.55, 271.05, 271.55, 
    271.95, 271.95, 272.55, 272.85, 273.15, 272.65, 272.35, 272.25, 271.55, 
    271.65, 271.55, 271.25, 271.05, 271.95, 272.35, 272.25, 272.45, 272.15, 
    272.35, 271.75, 271.55, 270.95, 270.85, 270.25, 269.85, 269.65, 269.25, 
    269.05, 269.25, 269.15, 268.95, 267.05, 267.05, 267.95, 267.45, 267.35, 
    267.05, 266.85, 267.85, 267.95, 267.95, 268.25, 268.65, 268.25, 268.25, 
    268.45, 268.35, 268.45, 268.75, 269.15, 268.75, 270.85, 270.75, 270.85, 
    270.95, 271.45, 271.75, 271.45, 271.75, 271.45, 271.55, 271.15, 270.55, 
    270.45, 270.15, 269.85, 270.05, 270.25, 270.35, 270.95, 270.85, 270.45, 
    270.95, 271.75, 272.05, 272.55, 272.85, 272.35, 272.85, 272.95, 272.95, 
    272.95, 273.45, 274.15, 274.25, 273.85, 273.25, 272.95, 272.75, 273.05, 
    272.95, 272.55, 272.85, 272.65, 272.75, 272.65, 272.35, 272.35, 272.25, 
    272.15, 271.95, 271.55, 271.75, 271.05, 271.45, 271.15, 270.75, 270.35, 
    269.85, 269.65, 269.35, 266.15, 264.65, 265.85, 265.35, 265.45, 267.15, 
    267.85, 268.65, 268.95, 267.45, 268.85, 271.15, 273.15, 272.25, 271.05, 
    269.55, 271.75, 270.35, 273.55, 273.35, 273.15, 273.25, 272.65, 272.95, 
    272.05, 272.25, 271.95, 272.05, 271.95, 272.05, 272.05, 272.25, 271.65, 
    271.35, 270.75, 269.95, 269.75, 269.55, 269.25, 269.05, 268.95, 268.25, 
    267.65, 267.45, 267.25, 267.15, 266.95, 265.45, 266.65, 266.65, 265.05, 
    264.55, 264.85, 264.55, 263.35, 264.45, 264.95, 264.95, 263.75, 264.15, 
    265.05, 265.45, 265.75, 265.75, 266.05, 265.85, 265.85, 265.75, 265.75, 
    265.85, 265.65, 265.85, 266.15, 266.35, 265.75, 266.15, 265.75, 265.35, 
    265.75, 266.05, 265.95, 266.55, 266.85, 267.35, 267.05, 267.35, 267.25, 
    267.65, 267.75, 267.55, 267.55, 268.65, 268.65, 269.05, 269.15, 269.15, 
    269.05, 268.85, 268.85, 268.95, 269.05, 270.15, 270.55, 269.65, 269.35, 
    269.85, 269.55, 269.05, 269.65, 270.05, 269.65, 269.05, 268.85, 268.65, 
    268.45, 268.45, 268.45, 268.45, 268.05, 268.25, 267.35, 268.05, 267.15, 
    265.45, 265.35, 264.65, 265.25, 265.05, 263.65, 263.15, 264.25, 263.75, 
    262.75, 263.45, 263.65, 263.55, 265.05, 265.85, 266.35, 266.55, 267.25, 
    267.65, 267.15, 266.75, 266.75, 267.55, 267.85, 267.65, 268.45, 269.05, 
    268.75, 270.45, 272.05, 272.95, 273.15, 273.75, 273.55, 273.55, 272.35, 
    272.15, 272.85, 272.95, 273.15, 273.35, 273.35, 273.25, 272.95, 273.35, 
    273.15, 272.85, 272.75, 273.05, 272.85, 273.85, 273.75, 272.85, 271.85, 
    272.05, 270.25, 269.15, 271.05, 270.95, 271.25, 271.45, 271.35, 272.45, 
    272.35, 271.75, 271.55, 271.05, 270.15, 270.75, 270.95, 271.25, 271.15, 
    271.35, 271.95, 272.05, 272.35, 272.35, 272.55, 272.05, 270.75, 271.65, 
    271.25, 271.45, 273.55, 273.15, 271.65, 271.85, 271.65, 272.45, 273.75, 
    273.35, 273.35, 273.75, 273.75, 273.85, 273.45, 273.45, 274.05, 274.15, 
    274.25, 274.25, 274.25, 274.15, 274.25, 274.15, 273.45, 273.05, 272.15, 
    270.05, 270.55, 270.25, 267.45, 269.35, 273.25, 273.55, 273.35, 273.55, 
    273.55, 273.65, 273.85, 273.75, 273.55, 273.45, 273.25, 273.55, 273.55, 
    273.85, 274.15, 274.35, 274.55, 273.75, 274.25, 273.95, 274.05, 273.25, 
    273.45, 273.35, 272.65, 272.25, 271.95, 271.35, 271.45, 271.15, 270.35, 
    270.05, 267.75, 267.05, 267.15, 268.55, 266.95, 264.45, 268.05, 270.25, 
    269.85, 269.25, 268.95, 269.55, 268.85, 268.15, 269.75, 269.75, 270.05, 
    270.05, 269.95, 270.25, 269.85, 270.15, 270.45, 270.35, 270.45, 270.75, 
    270.65, 270.85, 270.45, 271.05, 270.85, 270.75, 270.15, 270.35, 270.45, 
    267.75, 265.65, 267.05, 266.35, 266.85, 270.75, 269.15, 269.15, 269.05, 
    269.15, 269.35, 269.15, 269.05, 269.05, 269.25, 268.85, 269.15, 269.25, 
    269.35, 268.85, 269.05, 268.25, 268.75, 269.05, 268.55, 268.45, 268.65, 
    268.95, 268.75, 267.95, 267.75, 267.85, 267.75, 266.95, 266.35, 266.05, 
    265.55, 264.95, 264.25, 263.55, 263.55, 263.45, 263.25, 263.55, 263.85, 
    262.75, 263.15, 261.05, 262.55, 261.95, 263.05, 262.65, 262.75, 263.25, 
    263.85, 264.75, 264.95, 265.05, 266.85, 264.15, 261.25, 261.15, 260.35, 
    260.65, 261.25, 261.35, 261.35, 261.25, 261.65, 260.95, 260.55, 262.35, 
    261.55, 261.85, 260.75, 260.45, 259.55, 259.15, 258.85, 258.55, 257.85, 
    255.95, 256.05, 257.05, 256.95, 256.65, 255.65, 256.25, 255.85, 255.35, 
    255.65, 256.05, 256.15, 256.15, 255.65, 255.65, 255.85, 256.35, 255.55, 
    256.15, 256.25, 255.35, 254.95, 256.25, 256.85, 257.25, 256.65, 255.85, 
    255.15, 255.05, 254.65, 254.65, 254.35, 255.65, 255.25, 255.65, 254.85, 
    253.95, 255.95, 254.15, 255.25, 254.95, 254.75, 256.05, 254.95, 256.35, 
    255.25, 255.95, 255.75, 256.25, 256.25, 256.05, 255.95, 255.75, 256.05, 
    255.65, 256.15, 256.05, 256.15, 256.75, 257.55, 256.05, 257.45, 256.65, 
    256.15, 257.15, 257.05, 256.65, 257.65, 257.65, 255.95, 257.35, 257.65, 
    257.05, 257.55, 256.85, 257.15, 257.35, 257.75, 258.15, 258.05, 258.35, 
    258.85, 258.35, 258.05, 258.15, 257.15, 258.15, 258.25, 257.75, 257.75, 
    257.65, 257.95, 258.85, 257.75, 258.95, 257.85, 257.65, 258.05, 257.35, 
    258.05, 257.45, 258.95, 259.65, 257.95, 259.15, 259.75, 260.45, 259.95, 
    262.15, 263.05, 262.25, 260.35, 259.15, 259.15, 259.55, 259.45, 259.15, 
    257.15, 256.55, 257.65, 257.35, 258.45, 258.85, 258.95, 258.05, 257.65, 
    256.25, 256.65, 256.35, 256.55, 257.25, 257.05, 256.25, 257.55, 255.45, 
    256.75, 257.15, 256.95, 255.35, 256.25, 257.45, 255.15, 256.65, 254.65, 
    255.95, 256.75, 257.45, 256.35, 257.05, 256.25, 257.75, 257.55, 257.15, 
    258.65, 258.45, 258.95, 259.95, 260.05, 259.95, 260.85, 261.05, 260.95, 
    261.65, 261.35, 260.85, 261.05, 262.25, 261.95, 261.65, 260.55, 260.85, 
    262.05, 261.75, 262.85, 262.15, 263.15, 262.45, 263.45, 263.35, 264.15, 
    265.55, 265.75, 265.85, 266.25, 266.15, 266.15, 266.25, 267.05, 266.65, 
    267.05, 267.35, 267.15, 267.15, 267.55, 267.85, 267.85, 268.15, 268.15, 
    267.35, 267.25, 266.15, 265.85, 265.95, 265.75, 264.55, 264.75, 264.75, 
    262.95, 261.75, 262.35, 261.95, 262.45, 261.95, 261.55, 261.15, 261.15, 
    263.15, 263.05, 263.75, 264.65, 265.55, 267.45, 268.05, 267.55, 268.35, 
    268.15, 268.85, 268.95, 269.45, 269.25, 269.85, 269.45, 269.95, 270.45, 
    271.25, 269.45, 270.25, 270.85, 270.85, 271.35, 271.05, 271.05, 270.75, 
    270.15, 269.85, 268.65, 267.95, 267.95, 268.05, 268.75, 268.45, 266.95, 
    267.65, 267.85, 269.15, 269.15, 269.25, 269.75, 269.15, 268.75, 268.85, 
    268.75, 269.55, 269.25, 268.85, 268.95, 269.75, 269.75, 269.65, 269.65, 
    268.75, 270.05, 270.25, 270.05, 270.15, 270.45, 270.35, 269.85, 269.25, 
    269.15, 268.75, 266.15, 266.95, 266.65, 267.45, 267.55, 267.25, 266.45, 
    267.65, 268.05, 268.25, 268.65, 268.95, 269.05, 269.05, 269.55, 269.45, 
    269.85, 270.45, 269.95, 269.95, 269.85, 270.25, 270.35, 270.15, 270.35, 
    269.95, 270.15, 270.15, 270.05, 270.75, 271.55, 270.85, 270.35, 270.55, 
    270.75, 271.15, 271.05, 271.55, 271.15, 271.25, 271.25, 271.35, 270.05, 
    270.05, 270.35, 270.25, 270.35, 269.75, 270.05, 270.35, 270.45, 270.65, 
    271.25, 271.35, 271.65, 271.35, 271.25, 271.95, 271.95, 271.95, 271.55, 
    271.15, 272.15, 272.25, 272.15, 271.65, 271.65, 272.45, 273.75, 273.55, 
    273.45, 273.25, 273.45, 273.15, 272.85, 272.55, 272.25, 272.35, 271.85, 
    272.05, 272.25, 272.85, 272.05, 272.05, 272.95, 273.65, 275.95, 277.75, 
    277.15, 277.05, 275.95, 277.05, 277.35, 277.55, 277.05, 277.45, 277.35, 
    277.25, 277.35, 277.15, 276.85, 276.65, 276.35, 275.85, 275.45, 275.05, 
    274.05, 273.35, 272.85, 272.35, 272.15, 271.55, 271.55, 271.65, 271.25, 
    271.25, 271.25, 271.05, 270.85, 270.85, 270.85, 270.95, 270.85, 270.95, 
    270.85, 271.45, 271.35, 272.35, 272.85, 272.15, 272.75, 272.95, 272.15, 
    272.15, 272.45, 273.35, 272.75, 273.25, 274.85, 274.15, 274.65, 274.85, 
    274.55, 274.15, 273.65, 273.05, 272.35, 273.45, 273.85, 273.55, 273.55, 
    273.65, 272.65, 272.75, 274.15, 274.15, 273.95, 273.25, 273.15, 272.65, 
    272.45, 271.75, 271.25, 270.65, 270.15, 271.05, 271.15, 271.35, 271.15, 
    271.05, 271.15, 271.35, 271.35, 271.15, 271.25, 271.65, 271.45, 271.75, 
    271.75, 271.25, 271.75, 271.45, 270.75, 270.75, 270.65, 270.85, 270.65, 
    270.35, 269.95, 270.25, 269.95, 269.75, 270.75, 270.55, 270.75, 271.25, 
    271.05, 271.35, 271.25, 271.05, 271.35, 270.95, 271.05, 271.15, 270.15, 
    270.35, 270.95, 271.15, 271.15, 271.25, 270.75, 270.75, 270.75, 270.05, 
    270.65, 272.05, 272.25, 272.25, 272.05, 271.75, 269.55, 268.55, 267.65, 
    268.45, 268.05, 268.05, 268.05, 268.05, 269.15, 269.05, 268.85, 269.45, 
    268.75, 268.65, 268.95, 269.25, 270.25, 270.25, 270.35, 269.85, 270.75, 
    270.55, 270.45, 269.85, 269.55, 269.05, 268.75, 268.75, 268.65, 268.65, 
    268.55, 268.25, 267.85, 267.75, 267.65, 268.15, 268.15, 268.75, 269.05, 
    268.65, 269.45, 268.75, 268.65, 268.35, 267.85, 266.65, 265.95, 265.45, 
    265.15, 264.95, 264.65, 264.25, 263.85, 263.55, 263.35, 263.25, 265.85, 
    264.85, 264.25, 263.55, 263.45, 263.25, 263.05, 262.85, 265.35, 265.85, 
    264.95, 264.15, 265.65, 266.05, 266.35, 266.55, 265.65, 265.65, 268.25, 
    267.35, 266.85, 266.95, 267.35, 269.05, 267.95, 268.05, 268.35, 268.15, 
    267.75, 267.75, 267.65, 267.15, 266.95, 267.45, 267.75, 268.45, 267.75, 
    266.25, 267.65, 268.85, 268.95, 268.55, 268.25, 267.75, 267.35, 268.35, 
    268.65, 268.15, 268.15, 268.15, 268.05, 268.05, 268.05, 267.85, 267.95, 
    267.95, 267.75, 269.15, 269.55, 269.55, 268.45, 268.45, 268.75, 268.75, 
    268.45, 269.45, 268.75, 268.45, 267.65, 267.85, 267.95, 268.25, 267.95, 
    267.95, 267.75, 267.05, 265.95, 264.85, 266.35, 266.45, 266.25, 266.45, 
    266.85, 266.95, 264.95, 264.45, 265.75, 266.05, 265.95, 264.95, 265.25, 
    264.95, 263.25, 263.15, 262.65, 261.75, 263.35, 263.95, 264.15, 264.15, 
    264.35, 264.35, 262.65, 263.45, 263.25, 263.45, 263.55, 263.65, 263.85, 
    263.85, 264.35, 264.75, 263.85, 264.15, 263.35, 263.05, 263.25, 263.35, 
    263.25, 263.45, 263.15, 262.85, 262.85, 262.65, 261.35, 260.55, 261.65, 
    261.55, 261.15, 261.05, 261.25, 260.85, 260.95, 261.05, 261.35, 261.85, 
    261.65, 261.25, 259.85, 259.15, 259.15, 259.35, 259.15, 259.15, 258.05, 
    258.15, 257.65, 257.75, 257.95, 258.25, 258.65, 259.45, 260.35, 261.35, 
    263.55, 264.75, 264.65, 264.65, 264.15, 263.45, 262.65, 264.45, 264.35, 
    264.45, 264.95, 265.75, 266.75, 265.55, 264.65, 264.05, 263.35, 263.05, 
    262.95, 262.95, 262.75, 262.35, 260.75, 261.55, 262.25, 262.55, 260.05, 
    261.25, 259.15, 258.55, 258.75, 258.55, 258.15, 257.85, 257.55, 257.45, 
    257.65, 257.65, 259.15, 258.05, 257.65, 257.55, 257.45, 257.35, 257.25, 
    257.15, 257.15, 257.05, 256.55, 256.05, 258.55, 257.95, 259.05, 259.45, 
    259.25, 259.05, 258.95, 258.85, 258.85, 258.85, 258.65, 259.05, 259.25, 
    259.15, 258.95, 258.95, 258.85, 258.85, 258.75, 258.95, 258.75, 258.55, 
    257.95, 258.45, 258.15, 258.75, 258.35, 257.45, 257.35, 256.95, 256.65, 
    256.55, 256.45, 256.45, 256.55, 256.85, 257.45, 257.15, 256.65, 256.25, 
    256.05, 256.15, 256.05, 256.25, 256.55, 256.15, 256.05, 255.85, 256.85, 
    256.55, 255.75, 255.35, 255.15, 255.05, 255.45, 255.95, 255.85, 257.55, 
    258.45, 258.75, 256.45, 255.85, 255.25, 254.55, 256.65, 257.85, 258.45, 
    257.75, 256.45, 255.85, 255.45, 255.05, 256.55, 256.35, 255.85, 255.45, 
    255.15, 255.15, 255.05, 254.85, 254.75, 254.75, 258.65, 258.75, 255.45, 
    256.05, 258.55, 258.65, 259.25, 260.25, 260.95, 260.55, 259.95, 259.35, 
    259.05, 258.95, 259.05, 259.05, 259.95, 260.65, 260.95, 261.25, 263.75, 
    265.75, 266.95, 267.55, 267.45, 267.35, 267.15, 266.45, 267.45, 267.95, 
    266.85, 266.25, 265.25, 265.75, 267.85, 267.25, 267.85, 267.95, 267.45, 
    270.35, 271.35, 272.15, 272.45, 272.65, 272.35, 272.65, 272.85, 273.25, 
    272.65, 272.15, 272.15, 272.05, 272.55, 273.45, 273.35, 272.75, 272.35, 
    272.35, 272.05, 271.35, 271.05, 270.75, 270.55, 271.45, 272.05, 271.75, 
    271.75, 272.15, 273.15, 273.45, 274.25, 275.25, 274.45, 274.05, 273.95, 
    273.65, 272.95, 273.15, 272.45, 271.65, 271.45, 271.25, 270.85, 270.55, 
    270.25, 270.55, 270.05, 270.35, 269.65, 269.45, 270.45, 271.05, 270.95, 
    270.45, 269.65, 268.75, 268.05, 267.65, 267.55, 266.95, 265.85, 265.15, 
    264.35, 266.15, 267.05, 268.05, 268.35, 268.45, 269.35, 268.25, 266.65, 
    265.65, 265.25, 265.05, 264.85, 264.85, 265.35, 265.25, 265.35, 266.05, 
    266.85, 267.35, 266.85, 268.25, 268.45, 268.65, 269.15, 269.35, 268.75, 
    268.75, 268.35, 268.95, 268.65, 267.75, 265.45, 264.15, 263.45, 262.45, 
    261.85, 264.45, 266.35, 266.85, 267.05, 267.35, 268.55, 268.25, 268.55, 
    268.95, 269.25, 268.65, 268.05, 267.75, 266.85, 266.95, 264.75, 263.35, 
    263.35, 263.95, 262.45, 262.05, 261.55, 260.95, 260.45, 260.15, 260.25, 
    262.75, 264.25, 264.95, 265.35, 265.75, 266.05, 267.45, 265.25, 264.65, 
    264.05, 263.15, 267.15, 267.35, 266.55, 265.85, 267.95, 267.95, 270.05, 
    270.05, 269.95, 270.35, 271.45, 271.55, 272.25, 273.15, 273.05, 273.05, 
    273.05, 273.15, 271.65, 269.35, 269.15, 270.25, 271.05, 271.95, 271.85, 
    272.05, 271.85, 271.95, 271.75, 271.55, 272.55, 272.25, 271.45, 271.75, 
    272.55, 272.15, 270.75, 270.05, 270.25, 270.35, 270.75, 271.05, 271.25, 
    271.25, 270.35, 271.85, 271.75, 271.35, 270.75, 269.85, 269.05, 268.35, 
    267.45, 266.75, 266.15, 265.85, 265.35, 264.95, 264.85, 264.85, 264.25, 
    263.45, 261.95, 260.55, 259.85, 259.45, 260.25, 260.05, 260.05, 259.55, 
    259.15, 258.75, 258.95, 259.05, 258.95, 258.95, 258.75, 259.05, 262.95, 
    263.75, 264.15, 264.45, 264.85, 265.05, 265.25, 265.25, 265.35, 265.45, 
    265.45, 265.45, 265.65, 265.25, 264.85, 264.45, 264.75, 264.95, 264.95, 
    264.85, 265.05, 265.75, 265.75, 265.15, 265.65, 265.05, 262.75, 261.15, 
    261.15, 261.25, 260.95, 260.85, 260.85, 260.65, 260.55, 260.35, 260.35, 
    260.35, 260.05, 259.75, 259.55, 259.55, 259.55, 259.25, 259.15, 259.25, 
    259.25, 259.25, 260.55, 260.35, 260.15, 260.05, 259.85, 259.65, 259.55, 
    259.55, 259.45, 259.35, 259.25, 258.95, 257.65, 257.55, 257.35, 260.55, 
    261.45, 260.95, 261.55, 261.25, 260.15, 256.55, 256.55, 256.55, 258.45, 
    258.35, 257.95, 257.85, 257.85, 257.75, 257.55, 257.35, 257.15, 257.05, 
    256.85, 256.75, 256.45, 256.35, 256.15, 255.95, 255.85, 255.85, 255.85, 
    255.75, 255.75, 255.75, 255.75, 255.55, 255.55, 255.85, 256.15, 256.25, 
    256.05, 255.85, 255.65, 255.65, 255.55, 255.55, 255.45, 255.45, 255.15, 
    255.15, 255.25, 255.05, 254.85, 254.65, 254.65, 254.55, 254.45, 254.25, 
    253.75, 253.55, 252.15, 252.45, 252.65, 252.75, 252.35, 252.05, 251.75, 
    251.55, 251.65, 251.85, 252.05, 252.35, 254.05, 254.05, 254.05, 253.65, 
    253.35, 253.35, 253.35, 253.35, 253.45, 253.85, 254.35, 254.75, 257.65, 
    257.55, 257.55, 257.65, 257.75, 257.65, 257.65, 257.75, 257.85, 257.85, 
    257.85, 257.85, 259.05, 258.95, 259.05, 259.35, 259.35, 259.15, 259.05, 
    259.05, 259.05, 259.15, 259.65, 259.75, 261.05, 260.75, 260.55, 261.45, 
    262.65, 263.35, 262.85, 262.55, 261.95, 261.75, 261.85, 261.55, 259.55, 
    259.95, 260.35, 260.25, 260.35, 260.25, 259.35, 259.05, 258.75, 258.75, 
    258.65, 258.65, 258.55, 258.25, 258.45, 257.35, 257.35, 257.35, 256.25, 
    259.75, 259.65, 257.55, 256.75, 256.35, 257.55, 256.95, 256.25, 255.45, 
    254.75, 254.25, 254.05, 253.65, 253.35, 253.55, 253.65, 253.65, 254.05, 
    253.95, 253.45, 252.65, 252.55, 253.05, 253.15, 253.35, 253.55, 253.75, 
    253.75, 253.45, 253.65, 253.35, 252.95, 253.45, 253.45, 253.65, 254.05, 
    254.45, 255.25, 255.45, 255.45, 254.65, 256.55, 256.75, 256.95, 256.95, 
    261.05, 263.55, 264.75, 264.85, 264.95, 265.15, 265.45, 265.85, 266.85, 
    267.15, 267.25, 267.25, 267.35, 267.45, 267.55, 267.45, 267.45, 267.65, 
    267.65, 267.35, 266.65, 266.85, 267.45, 268.45, 269.95, 270.35, 270.05, 
    269.85, 269.95, 269.95, 269.95, 269.85, 270.55, 269.85, 269.55, 269.25, 
    269.55, 272.15, 271.55, 270.65, 270.35, 269.75, 269.55, 269.95, 269.95, 
    269.95, 262.85, 262.65, 262.25, 261.95, 261.95, 261.45, 261.15, 260.75, 
    260.65, 260.65, 264.65, 264.45, 264.55, 264.45, 264.55, 264.45, 264.65, 
    265.65, 267.35, 268.55, 268.45, 272.85, 271.05, 273.05, 273.65, 274.05, 
    274.35, 274.75, 275.05, 275.25, 275.15, 274.95, 274.95, 274.85, 274.55, 
    274.55, 274.55, 274.75, 274.75, 274.85, 275.35, 275.35, 275.55, 275.55, 
    275.25, 275.25, 275.05, 274.65, 274.75, 274.75, 274.75, 274.75, 274.65, 
    274.55, 274.55, 274.45, 274.45, 274.45, 274.25, 274.15, 274.15, 274.25, 
    274.35, 274.35, 274.35, 274.05, 273.85, 274.05, 274.25, 273.65, 267.65, 
    266.65, 266.15, 265.95, 265.75, 265.15, 263.95, 263.35, 263.45, 262.95, 
    262.75, 262.15, 261.85, 261.55, 261.15, 260.55, 263.05, 262.95, 262.55, 
    262.45, 261.55, 260.95, 261.05, 260.55, 260.15, 259.85, 259.95, 260.25, 
    260.05, 259.65, 259.45, 259.45, 258.75, 259.35, 258.95, 258.85, 258.85, 
    257.35, 257.25, 257.85, 258.65, 257.85, 257.55, 257.55, 257.05, 257.35, 
    256.95, 257.25, 256.75, 257.55, 259.25, 260.15, 260.65, 261.05, 260.95, 
    260.75, 261.85, 262.05, 262.35, 261.85, 262.25, 262.45, 262.15, 262.15, 
    262.25, 262.45, 261.95, 261.95, 262.45, 262.45, 261.95, 261.75, 262.15, 
    262.45, 262.35, 263.25, 261.35, 260.45, 259.55, 259.05, 259.05, 258.65, 
    258.75, 258.85, 258.85, 261.15, 261.35, 261.35, 262.05, 262.75, 261.45, 
    260.35, 261.15, 262.15, 262.75, 262.35, 262.55, 261.75, 263.45, 263.75, 
    263.05, 262.95, 262.35, 263.55, 263.35, 263.15, 263.55, 262.85, 261.25, 
    260.75, 260.35, 261.45, 260.85, 260.55, 258.95, 260.05, 260.25, 260.45, 
    260.15, 260.05, 259.95, 259.75, 261.05, 260.55, 261.25, 259.95, 262.25, 
    262.45, 261.75, 260.65, 259.35, 260.15, 258.55, 261.25, 258.65, 259.95, 
    260.05, 260.75, 259.25, 258.65, 258.45, 257.45, 257.25, 257.95, 258.25, 
    258.05, 257.45, 257.95, 258.25, 258.05, 257.95, 258.15, 257.45, 257.75, 
    257.65, 258.15, 257.65, 257.45, 256.75, 257.25, 256.75, 257.95, 256.15, 
    256.55, 256.85, 256.15, 256.35, 254.75, 255.05, 254.55, 256.25, 254.45, 
    256.45, 255.15, 254.65, 254.25, 255.25, 253.95, 254.75, 253.95, 254.25, 
    254.85, 253.25, 254.95, 255.55, 256.15, 254.15, 254.65, 255.05, 253.75, 
    254.05, 253.75, 253.55, 252.35, 254.25, 253.15, 252.55, 252.95, 253.55, 
    252.75, 252.65, 252.05, 252.65, 253.35, 252.25, 253.45, 251.75, 252.65, 
    254.85, 254.65, 252.75, 252.85, 253.25, 252.55, 253.15, 251.65, 252.65, 
    252.85, 252.05, 251.55, 252.45, 251.35, 251.95, 251.45, 251.95, 252.25, 
    251.15, 252.35, 251.25, 251.55, 251.45, 254.05, 253.15, 255.05, 252.25, 
    252.55, 252.95, 252.85, 251.45, 251.95, 252.25, 251.45, 251.55, 253.65, 
    252.15, 251.75, 251.65, 251.85, 252.55, 252.75, 252.45, 252.95, 252.35, 
    252.45, 254.85, 254.95, 255.55, 255.55, 253.85, 254.25, 253.95, 254.85, 
    254.45, 254.35, 254.85, 256.45, 256.05, 254.65, 254.55, 254.65, 255.55, 
    257.55, 256.85, 254.05, 256.35, 254.15, 255.05, 254.95, 255.95, 255.75, 
    258.65, 257.35, 256.05, 257.55, 254.75, 257.45, 256.05, 254.95, 255.75, 
    255.05, 254.45, 255.05, 254.15, 254.45, 253.75, 254.05, 254.35, 254.15, 
    253.65, 253.75, 253.75, 255.85, 254.25, 254.75, 256.65, 258.15, 256.15, 
    255.35, 254.55, 255.65, 256.05, 254.15, 255.75, 254.25, 255.15, 255.25, 
    255.65, 255.55, 254.65, 253.85, 256.85, 256.25, 253.75, 256.65, 254.15, 
    255.55, 256.65, 256.65, 257.95, 257.35, 256.25, 256.05, 256.95, 254.45, 
    253.55, 255.25, 256.75, 254.55, 254.35, 254.75, 255.75, 255.75, 255.65, 
    255.85, 254.75, 256.35, 256.75, 255.05, 255.15, 256.25, 257.15, 257.25, 
    259.45, 257.85, 258.75, 258.95, 258.25, 257.95, 258.55, 257.05, 257.75, 
    257.35, 256.55, 257.05, 257.05, 259.45, 256.35, 256.45, 258.75, 256.25, 
    257.75, 256.55, 255.35, 257.05, 257.75, 257.65, 258.45, 258.35, 258.95, 
    258.55, 257.65, 259.65, 258.65, 260.65, 260.35, 261.25, 262.05, 260.85, 
    260.85, 261.25, 261.25, 261.65, 261.35, 261.85, 263.05, 263.25, 263.05, 
    263.25, 263.15, 264.05, 264.65, 264.45, 264.75, 263.95, 264.35, 265.05, 
    264.15, 264.95, 267.25, 264.85, 264.95, 265.25, 266.05, 266.95, 268.75, 
    268.95, 267.15, 269.55, 271.85, 271.55, 272.45, 271.85, 272.75, 272.55, 
    272.95, 273.35, 273.35, 273.25, 273.45, 273.45, 273.35, 272.65, 272.25, 
    272.15, 271.65, 271.65, 271.05, 270.55, 270.65, 270.85, 269.35, 268.35, 
    267.75, 267.45, 267.15, 266.95, 267.05, 266.85, 266.55, 266.55, 266.35, 
    265.95, 265.05, 264.35, 263.35, 262.65, 261.85, 261.05, 260.35, 259.55, 
    259.25, 259.05, 258.45, 257.05, 256.25, 256.05, 255.95, 255.15, 254.75, 
    254.85, 256.55, 257.25, 256.45, 256.35, 257.05, 255.75, 255.15, 254.45, 
    255.25, 254.45, 253.45, 253.15, 252.95, 253.15, 251.95, 253.35, 252.25, 
    252.95, 251.85, 252.05, 251.45, 251.55, 252.55, 252.55, 252.95, 253.95, 
    254.65, 255.25, 254.55, 254.55, 254.55, 255.25, 254.35, 255.55, 254.45, 
    255.05, 254.25, 255.25, 254.95, 255.55, 254.85, 254.45, 255.15, 255.85, 
    255.25, 255.05, 255.85, 256.25, 255.45, 255.65, 256.35, 256.05, 258.25, 
    255.75, 256.25, 256.15, 255.55, 255.65, 255.85, 254.45, 253.85, 252.45, 
    253.15, 252.05, 251.95, 251.85, 252.65, 252.15, 253.15, 254.05, 253.15, 
    253.45, 254.25, 254.15, 255.35, 260.55, 261.15, 261.05, 261.95, 261.15, 
    263.25, 263.35, 263.35, 262.45, 262.65, 262.75, 262.25, 260.55, 261.95, 
    263.15, 263.15, 261.65, 260.35, 263.15, 263.45, 263.05, 263.15, 263.25, 
    264.45, 264.25, 264.25, 264.25, 264.45, 263.65, 262.95, 262.45, 260.85, 
    260.35, 259.25, 260.35, 256.25, 258.05, 257.75, 260.85, 261.25, 262.05, 
    261.25, 261.45, 260.15, 260.35, 259.05, 258.35, 259.65, 259.25, 260.05, 
    263.35, 261.75, 262.75, 263.45, 262.95, 262.55, 261.85, 261.55, 260.35, 
    259.35, 260.25, 258.45, 258.95, 258.15, 257.35, 258.75, 258.35, 258.55, 
    259.15, 259.65, 258.45, 260.55, 262.15, 263.15, 261.35, 260.95, 260.65, 
    259.75, 259.35, 259.95, 259.05, 258.95, 258.55, 259.05, 259.15, 259.25, 
    263.45, 262.85, 263.05, 264.35, 262.95, 264.65, 263.95, 265.15, 265.65, 
    266.15, 266.05, 264.75, 264.95, 265.05, 265.25, 265.15, 265.55, 264.75, 
    264.05, 263.85, 263.45, 261.85, 260.95, 260.85, 260.75, 260.05, 258.85, 
    259.45, 259.45, 260.15, 259.35, 261.05, 261.35, 261.55, 261.65, 262.65, 
    261.15, 260.55, 259.45, 260.35, 260.45, 260.55, 259.75, 259.55, 259.45, 
    259.15, 259.45, 259.95, 260.75, 260.95, 261.35, 260.85, 261.85, 261.05, 
    261.15, 261.25, 262.35, 264.35, 264.45, 264.45, 263.75, 263.45, 262.55, 
    262.45, 262.15, 260.45, 258.85, 258.65, 258.35, 257.85, 258.85, 258.45, 
    256.95, 256.55, 257.25, 256.95, 255.15, 257.35, 257.35, 257.65, 257.55, 
    260.45, 260.45, 260.35, 260.05, 260.55, 260.65, 258.85, 258.15, 255.65, 
    256.05, 256.85, 256.55, 254.85, 255.75, 255.55, 254.95, 255.25, 255.05, 
    256.25, 256.75, 255.55, 256.75, 258.25, 258.75, 259.85, 259.15, 258.55, 
    259.95, 258.65, 258.65, 257.75, 256.55, 256.55, 255.65, 255.45, 255.25, 
    254.65, 254.85, 255.65, 254.05, 253.85, 253.15, 253.65, 254.15, 255.35, 
    255.65, 257.65, 256.85, 257.45, 257.05, 257.45, 257.85, 258.15, 257.95, 
    256.55, 256.15, 254.95, 253.55, 253.25, 254.85, 253.95, 255.25, 255.55, 
    256.35, 257.15, 258.05, 259.05, 259.35, 259.45, 259.45, 260.55, 260.15, 
    260.15, 259.95, 259.85, 259.35, 260.45, 260.25, 258.75, 258.25, 255.85, 
    256.45, 256.75, 256.25, 255.05, 256.65, 255.95, 254.95, 255.15, 256.05, 
    255.25, 256.65, 257.25, 255.55, 257.15, 259.95, 259.45, 260.35, 260.35, 
    259.75, 260.05, 258.45, 259.65, 258.65, 257.85, 257.35, 258.35, 257.85, 
    258.65, 257.25, 257.75, 257.55, 257.25, 258.05, 257.35, 257.25, 258.45, 
    258.85, 260.05, 261.35, 260.35, 260.55, 261.05, 261.65, 259.95, 260.65, 
    260.15, 259.75, 258.15, 257.65, 256.75, 257.25, 257.25, 257.55, 256.75, 
    256.15, 255.65, 255.75, 255.85, 257.05, 256.85, 258.05, 257.95, 260.25, 
    260.55, 261.05, 259.55, 259.55, 259.95, 259.35, 258.85, 257.85, 256.75, 
    256.95, 256.65, 257.05, 255.45, 256.25, 255.05, 255.35, 255.25, 252.95, 
    254.65, 254.25, 255.65, 257.15, 257.05, 258.55, 258.05, 259.55, 259.15, 
    259.05, 260.15, 259.25, 259.05, 257.45, 256.65, 255.85, 256.45, 254.95, 
    256.25, 256.85, 254.75, 254.35, 255.35, 255.65, 256.95, 257.45, 257.05, 
    257.15, 258.65, 259.05, 261.05, 259.05, 259.65, 259.25, 260.95, 261.55, 
    260.75, 259.85, 258.85, 257.85, 258.85, 257.45, 257.35, 256.55, 256.35, 
    256.45, 256.05, 256.95, 256.55, 255.55, 256.15, 258.25, 258.55, 260.65, 
    259.45, 259.95, 260.15, 260.05, 259.05, 260.55, 258.25, 258.95, 258.55, 
    257.65, 256.25, 256.65, 257.45, 256.25, 256.05, 257.05, 255.65, 255.85, 
    257.25, 257.25, 257.15, 258.55, 261.05, 261.25, 261.95, 263.45, 262.15, 
    263.55, 263.05, 263.85, 261.05, 261.55, 261.15, 258.65, 260.75, 260.25, 
    259.65, 259.85, 261.75, 260.85, 260.65, 261.55, 259.15, 261.05, 262.05, 
    262.45, 262.25, 262.75, 262.85, 265.45, 264.85, 264.85, 266.05, 265.35, 
    265.25, 265.55, 265.55, 264.15, 264.35, 261.45, 260.95, 260.25, 260.35, 
    260.05, 257.85, 255.25, 256.15, 258.05, 258.75, 258.45, 257.65, 258.65, 
    259.65, 260.55, 262.35, 258.85, 261.25, 259.95, 259.65, 258.75, 259.45, 
    257.25, 257.85, 256.25, 259.25, 258.35, 258.95, 260.55, 260.35, 259.95, 
    261.15, 261.55, 262.35, 262.45, 263.25, 263.55, 263.35, 264.05, 264.65, 
    265.05, 265.95, 265.75, 266.55, 265.85, 265.25, 265.15, 264.75, 265.05, 
    265.85, 265.95, 265.85, 266.35, 265.35, 266.15, 265.55, 265.65, 265.85, 
    266.15, 266.65, 267.35, 267.15, 267.85, 267.85, 268.15, 268.65, 269.15, 
    268.85, 268.55, 270.95, 273.85, 274.15, 274.25, 273.85, 273.35, 272.65, 
    272.65, 272.75, 271.95, 270.85, 270.95, 271.05, 270.85, 270.15, 268.55, 
    269.05, 269.35, 269.75, 268.55, 267.75, 267.95, 267.05, 265.85, 264.25, 
    262.95, 263.05, 261.15, 262.15, 260.15, 261.95, 258.05, 259.45, 258.45, 
    260.45, 259.25, 261.05, 260.95, 262.05, 263.05, 260.25, 259.65, 264.15, 
    265.25, 264.55, 264.35, 264.45, 265.15, 264.85, 264.45, 264.05, 265.65, 
    266.55, 266.65, 261.65, 263.25, 262.05, 262.35, 261.95, 260.65, 263.05, 
    264.25, 264.25, 263.95, 267.65, 263.45, 263.85, 266.55, 265.25, 264.85, 
    265.65, 265.55, 265.35, 266.35, 265.05, 265.75, 266.15, 266.05, 266.75, 
    266.85, 267.05, 266.85, 268.35, 268.55, 268.55, 271.65, 270.85, 270.05, 
    270.95, 271.75, 271.95, 272.25, 270.95, 271.05, 271.25, 271.45, 270.95, 
    270.65, 270.15, 270.05, 269.85, 269.65, 269.65, 269.65, 270.05, 270.95, 
    271.25, 270.25, 270.45, 269.75, 268.25, 267.85, 269.45, 268.05, 267.45, 
    269.15, 266.15, 264.95, 264.95, 263.75, 263.95, 263.75, 263.15, 262.45, 
    258.45, 259.45, 262.15, 262.65, 262.15, 261.05, 260.25, 260.35, 261.45, 
    263.55, 263.85, 263.95, 263.95, 263.35, 263.55, 264.55, 262.75, 263.05, 
    263.75, 262.85, 262.65, 260.45, 259.85, 260.15, 260.15, 258.85, 258.95, 
    258.85, 259.35, 258.45, 260.45, 259.65, 260.05, 263.25, 263.35, 264.55, 
    262.95, 264.05, 266.25, 263.35, 264.15, 263.15, 263.45, 262.65, 261.15, 
    261.05, 258.35, 259.55, 259.25, 258.15, 256.75, 258.85, 255.35, 259.65, 
    258.85, 258.85, 260.85, 259.95, 262.55, 262.45, 263.55, 265.65, 262.05, 
    263.05, 263.75, 264.35, 264.65, 265.15, 264.55, 264.15, 263.95, 263.35, 
    263.25, 263.35, 263.65, 263.95, 264.15, 264.35, 264.85, 265.45, 267.45, 
    266.85, 267.45, 268.25, 268.95, 268.35, 268.35, 271.95, 271.65, 270.95, 
    269.35, 268.65, 268.45, 268.85, 268.75, 268.05, 267.45, 268.05, 268.35, 
    264.45, 265.95, 266.45, 263.05, 265.55, 266.25, 266.05, 267.05, 268.05, 
    268.65, 270.95, 270.25, 268.85, 269.25, 267.75, 267.25, 266.65, 265.05, 
    264.45, 263.75, 262.75, 260.95, 261.05, 261.15, 256.85, 259.05, 260.35, 
    259.75, 262.45, 261.85, 263.25, 264.65, 266.05, 265.65, 265.25, 266.55, 
    267.95, 265.15, 265.45, 264.35, 263.95, 263.85, 263.85, 263.75, 263.75, 
    263.65, 263.35, 262.85, 260.25, 259.25, 259.45, 260.05, 259.05, 261.25, 
    261.25, 261.95, 263.05, 262.85, 262.55, 263.35, 262.55, 262.05, 262.35, 
    263.95, 263.75, 260.65, 259.15, 257.55, 258.75, 258.55, 257.55, 255.95, 
    257.45, 256.35, 257.75, 258.05, 255.95, 257.95, 259.65, 261.35, 262.25, 
    262.55, 260.95, 261.25, 263.45, 262.45, 262.55, 261.95, 261.75, 261.55, 
    258.95, 258.05, 258.35, 257.25, 256.75, 257.05, 255.35, 256.25, 257.95, 
    256.75, 256.85, 259.65, 260.65, 262.75, 263.05, 264.55, 262.35, 263.45, 
    265.45, 261.55, 261.95, 261.65, 262.35, 261.75, 259.35, 258.15, 257.25, 
    256.45, 257.35, 257.25, 255.05, 256.55, 255.35, 257.95, 257.15, 260.15, 
    259.05, 262.35, 264.25, 262.65, 264.05, 264.25, 263.35, 265.55, 263.45, 
    262.15, 261.35, 261.35, 261.05, 260.25, 259.15, 260.15, 260.45, 258.75, 
    261.15, 261.05, 261.55, 262.15, 263.05, 265.65, 264.65, 265.15, 266.65, 
    264.95, 266.55, 267.05, 266.55, 266.75, 267.45, 266.95, 266.25, 265.45, 
    265.15, 263.35, 263.55, 263.95, 265.35, 264.85, 266.05, 265.05, 264.85, 
    265.55, 266.35, 266.65, 267.45, 267.35, 268.65, 270.25, 273.15, 270.55, 
    272.75, 268.45, 269.15, 268.95, 267.45, 266.25, 266.55, 266.25, 266.45, 
    265.85, 266.05, 265.55, 266.75, 267.15, 268.25, 267.25, 267.85, 268.85, 
    269.45, 270.85, 270.05, 270.25, 270.75, 270.65, 270.55, 270.35, 270.95, 
    270.95, 269.55, 270.45, 269.55, 269.55, 268.75, 268.55, 269.05, 269.35, 
    269.25, 268.65, 268.95, 270.25, 270.65, 270.65, 272.15, 270.65, 272.45, 
    272.55, 273.75, 273.45, 274.25, 275.15, 272.95, 274.35, 271.75, 272.35, 
    271.85, 271.65, 271.35, 271.25, 270.25, 271.05, 270.05, 270.85, 271.65, 
    270.55, 270.75, 271.55, 272.75, 272.95, 274.35, 273.45, 274.05, 273.65, 
    275.15, 273.25, 273.75, 274.75, 275.35, 275.35, 273.05, 270.05, 267.45, 
    268.95, 265.75, 267.75, 268.15, 267.85, 270.05, 269.85, 269.55, 271.85, 
    270.75, 272.85, 272.75, 274.15, 274.25, 274.25, 276.15, 277.45, 276.15, 
    275.95, 276.25, 276.55, 276.85, 276.45, 276.85, 277.35, 276.65, 276.65, 
    276.45, 276.35, 276.35, 277.55, 276.25, 276.75, 277.25, 277.15, 277.95, 
    277.95, 279.45, 277.55, 278.15, 277.95, 278.35, 278.35, 277.85, 275.65, 
    275.35, 274.75, 275.25, 274.85, 274.15, 271.55, 272.15, 272.45, 275.35, 
    275.45, 276.15, 276.65, 278.45, 278.55, 279.35, 279.65, 279.55, 279.65, 
    278.35, 280.25, 279.05, 278.45, 277.75, 277.35, 275.05, 275.45, 276.15, 
    276.15, 275.25, 275.15, 275.25, 274.85, 275.15, 275.65, 274.75, 273.85, 
    275.45, 276.25, 276.25, 275.85, 275.75, 274.85, 275.75, 276.05, 274.25, 
    274.35, 274.25, 274.35, 273.55, 273.15, 273.35, 273.45, 274.55, 274.65, 
    274.85, 274.55, 274.95, 274.45, 275.25, 274.85, 274.45, 274.15, 275.45, 
    275.35, 275.65, 275.75, 275.65, 275.75, 275.55, 275.05, 273.95, 274.05, 
    273.95, 274.55, 275.05, 275.45, 275.85, 275.45, 275.05, 275.25, 275.05, 
    274.95, 275.35, 276.55, 277.55, 275.15, 275.15, 274.95, 274.55, 274.45, 
    274.95, 275.05, 274.45, 274.05, 274.75, 273.75, 273.95, 274.05, 274.15, 
    274.25, 274.05, 273.45, 273.65, 273.65, 272.85, 273.65, 273.45, 273.65, 
    274.75, 273.95, 274.75, 274.55, 275.35, 275.15, 274.65, 273.95, 273.85, 
    273.45, 273.85, 275.05, 274.65, 275.05, 275.45, 275.15, 275.75, 275.65, 
    275.25, 275.25, 274.45, 273.95, 274.65, 275.15, 274.75, 275.95, 277.05, 
    277.65, 276.75, 276.95, 277.25, 276.55, 277.25, 276.15, 274.55, 274.15, 
    274.15, 273.95, 273.25, 273.35, 273.65, 273.85, 273.45, 273.75, 273.95, 
    274.35, 275.35, 275.05, 275.55, 275.55, 276.45, 277.45, 276.65, 276.75, 
    275.85, 275.05, 274.25, 273.95, 273.75, 273.55, 273.55, 273.35, 273.15, 
    273.05, 273.05, 272.75, 273.15, 273.45, 273.75, 274.05, 274.25, 274.75, 
    275.55, 275.65, 275.45, 275.55, 275.05, 275.35, 275.45, 275.75, 274.95, 
    275.15, 274.65, 274.55, 274.25, 273.75, 272.25, 271.85, 271.25, 272.75, 
    273.15, 273.55, 272.95, 273.45, 273.55, 274.15, 273.95, 273.95, 273.45, 
    273.65, 273.55, 273.65, 277.15, 276.25, 276.05, 275.05, 275.25, 274.75, 
    273.55, 273.45, 273.45, 272.65, 272.35, 273.15, 273.35, 272.25, 272.65, 
    272.65, 272.85, 273.85, 274.05, 274.75, 274.25, 275.45, 274.85, 274.85, 
    275.95, 275.65, 274.65, 274.95, 274.35, 274.15, 273.85, 273.55, 273.25, 
    272.55, 272.75, 271.85, 272.35, 271.55, 272.25, 272.25, 272.55, 272.25, 
    272.85, 273.85, 273.65, 273.75, 273.55, 274.35, 274.75, 273.65, 274.65, 
    274.25, 274.25, 274.65, 274.25, 273.85, 274.65, 274.65, 273.85, 273.85, 
    274.35, 275.15, 274.25, 274.65, 274.35, 275.95, 274.75, 274.85, 274.75, 
    274.55, 275.15, 275.25, 274.85, 274.65, 274.95, 274.65, 275.05, 275.05, 
    274.85, 275.05, 276.95, 277.45, 277.45, 277.55, 277.25, 277.75, 277.65, 
    277.05, 277.75, 278.05, 277.35, 277.25, 277.15, 277.55, 276.75, 276.85, 
    276.85, 276.95, 277.15, 275.95, 275.95, 276.35, 276.15, 276.45, 276.45, 
    275.85, 275.95, 276.05, 275.85, 276.35, 276.55, 276.45, 276.55, 276.15, 
    276.45, 276.45, 276.35, 276.45, 276.25, 276.25, 276.85, 277.55, 276.85, 
    276.25, 275.65, 276.35, 276.15, 276.05, 275.55, 275.15, 275.15, 275.15, 
    275.25, 275.65, 275.75, 275.85, 275.45, 275.35, 275.45, 275.65, 276.35, 
    276.45, 276.25, 276.45, 276.15, 276.05, 276.45, 276.05, 275.05, 274.85, 
    274.85, 275.05, 275.25, 274.55, 274.45, 274.75, 273.95, 274.45, 274.25, 
    274.95, 274.25, 274.95, 274.05, 274.35, 274.75, 275.25, 275.15, 275.85, 
    275.45, 275.15, 276.05, 275.75, 275.95, 275.65, 275.65, 274.25, 273.95, 
    273.55, 272.85, 272.85, 272.45, 272.55, 272.15, 272.65, 272.75, 273.25, 
    273.45, 274.25, 274.45, 274.45, 274.05, 274.45, 274.45, 274.45, 274.15, 
    273.65, 273.35, 273.35, 273.05, 272.75, 272.55, 272.45, 272.15, 272.05, 
    272.05, 271.95, 272.05, 272.25, 272.35, 272.35, 272.65, 272.45, 272.65, 
    273.15, 272.85, 272.95, 273.25, 273.35, 273.55, 273.45, 273.35, 273.45, 
    273.35, 273.15, 273.05, 273.15, 273.35, 273.15, 273.15, 273.35, 273.35, 
    273.55, 273.95, 274.25, 273.95, 274.35, 274.35, 275.05, 274.95, 274.65, 
    274.45, 274.15, 274.05, 274.25, 274.45, 273.75, 273.05, 272.95, 273.15, 
    273.65, 274.05, 274.55, 274.25, 274.25, 273.95, 274.45, 274.45, 274.25, 
    274.95, 275.85, 276.95, 277.95, 277.25, 277.85, 276.35, 277.25, 277.55, 
    277.55, 276.65, 276.15, 275.65, 275.05, 274.45, 274.65, 274.85, 274.75, 
    274.35, 274.65, 273.75, 273.55, 273.75, 273.75, 273.75, 273.75, 273.15, 
    273.45, 273.85, 274.15, 274.15, 274.05, 274.35, 273.45, 273.25, 273.35, 
    273.55, 273.45, 273.35, 272.85, 272.95, 272.65, 272.55, 272.45, 272.15, 
    272.15, 272.15, 272.15, 272.05, 272.25, 272.65, 272.65, 273.45, 273.85, 
    274.35, 273.95, 274.25, 274.35, 273.85, 273.95, 273.45, 273.05, 273.05, 
    272.95, 273.05, 272.95, 272.95, 272.85, 273.05, 273.35, 273.95, 274.15, 
    275.05, 275.25, 275.55, 275.45, 274.55, 274.65, 275.05, 274.65, 274.65, 
    274.35, 274.65, 274.55, 274.75, 274.25, 274.35, 274.15, 274.55, 274.35, 
    274.15, 274.35, 273.75, 274.15, 274.55, 274.15, 274.65, 274.95, 275.15, 
    275.75, 276.25, 276.25, 276.75, 276.95, 276.65, 276.85, 276.35, 276.75, 
    277.05, 276.55, 276.45, 275.95, 275.95, 276.35, 275.25, 274.75, 274.35, 
    274.05, 273.85, 273.75, 274.15, 274.05, 274.55, 273.95, 274.15, 274.35, 
    274.75, 274.75, 274.65, 275.05, 274.95, 274.75, 274.65, 274.95, 274.95, 
    274.75, 274.45, 274.35, 273.95, 274.05, 274.15, 274.35, 274.45, 274.15, 
    274.35, 274.45, 274.75, 275.05, 274.85, 275.05, 275.55, 276.45, 276.45, 
    275.85, 276.65, 276.45, 276.15, 275.85, 274.95, 275.05, 275.15, 274.95, 
    274.85, 274.85, 275.35, 275.75, 276.25, 276.25, 276.75, 277.25, 276.95, 
    276.75, 276.35, 277.15, 276.45, 276.25, 276.55, 276.65, 276.85, 277.15, 
    277.55, 277.35, 277.15, 276.75, 276.35, 276.45, 276.35, 276.45, 276.35, 
    276.85, 276.15, 276.95, 277.05, 278.45, 277.85, 278.05, 278.25, 277.65, 
    278.45, 278.25, 278.45, 278.35, 277.95, 277.65, 277.35, 277.15, 277.15, 
    276.35, 276.65, 276.45, 276.15, 275.95, 276.15, 275.95, 275.75, 275.85, 
    275.85, 275.95, 275.95, 276.25, 276.45, 276.85, 277.05, 276.05, 276.55, 
    276.15, 275.45, 275.05, 274.55, 274.75, 274.65, 274.65, 274.45, 274.25, 
    274.35, 273.95, 274.15, 274.15, 274.05, 274.15, 274.35, 274.85, 275.35, 
    275.45, 275.85, 275.75, 275.95, 276.05, 276.15, 276.25, 276.05, 275.75, 
    275.75, 275.75, 275.55, 275.65, 275.75, 275.55, 275.75, 275.75, 275.75, 
    276.05, 275.75, 276.15, 276.05, 276.05, 276.55, 276.75, 277.15, 277.15, 
    277.25, 277.05, 276.75, 277.15, 277.25, 276.55, 276.95, 276.05, 275.65, 
    275.45, 275.05, 274.95, 275.05, 274.95, 274.85, 274.85, 275.25, 275.45, 
    275.95, 275.95, 275.65, 275.45, 275.75, 275.25, 275.45, 275.35, 275.45, 
    274.65, 274.25, 274.35, 273.95, 273.75, 273.75, 273.65, 273.55, 273.55, 
    273.55, 273.45, 273.55, 273.75, 274.15, 274.25, 274.05, 274.45, 274.25, 
    274.65, 274.85, 275.25, 275.55, 275.35, 275.45, 275.55, 275.85, 276.15, 
    276.15, 276.35, 276.25, 275.95, 276.25, 276.05, 275.95, 276.55, 276.05, 
    276.75, 276.65, 276.45, 276.45, 278.25, 276.35, 276.35, 276.55, 276.15, 
    275.75, 275.75, 275.55, 275.25, 275.95, 275.45, 275.25, 275.45, 275.65, 
    275.85, 275.95, 276.05, 275.55, 275.75, 275.15, 275.35, 275.85, 275.85, 
    275.95, 277.15, 277.75, 277.65, 277.45, 276.75, 276.65, 276.55, 277.05, 
    277.45, 277.55, 277.35, 276.35, 275.75, 275.65, 275.65, 275.45, 275.25, 
    275.05, 275.05, 274.95, 274.95, 274.85, 274.75, 274.95, 275.05, 275.65, 
    275.65, 275.85, 275.85, 275.95, 275.85, 275.65, 275.75, 275.65, 275.35, 
    275.05, 274.75, 274.65, 274.55, 274.45, 274.25, 273.85, 273.55, 273.65, 
    273.55, 273.85, 273.95, 274.35, 274.45, 274.75, 274.95, 275.35, 275.65, 
    275.55, 275.35, 274.75, 274.95, 274.95, 274.85, 274.95, 274.85, 274.95, 
    274.95, 274.95, 274.85, 274.85, 274.85, 274.85, 275.15, 275.05, 275.25, 
    275.05, 275.25, 275.15, 275.35, 275.45, 275.15, 275.15, 275.15, 275.05, 
    275.05, 274.45, 273.85, 274.15, 273.55, 273.75, 273.45, 273.65, 273.75, 
    273.25, 272.35, 272.15, 272.85, 273.35, 273.35, 273.15, 273.45, 274.55, 
    274.75, 274.35, 274.75, 274.85, 274.85, 274.85, 275.35, 275.15, 275.15, 
    275.05, 274.45, 274.45, 274.65, 273.85, 273.55, 273.45, 273.65, 273.35, 
    273.55, 273.75, 274.05, 274.35, 274.65, 274.45, 274.65, 274.45, 274.45, 
    274.55, 274.35, 274.15, 274.25, 274.05, 274.15, 274.25, 274.25, 274.05, 
    274.75, 274.25, 274.25, 274.05, 274.25, 273.85, 273.85, 274.45, 274.75, 
    274.55, 275.15, 275.05, 275.45, 275.25, 275.85, 276.15, 275.85, 276.15, 
    276.35, 276.25, 276.15, 276.25, 275.75, 275.95, 275.75, 275.65, 275.85, 
    275.75, 275.85, 276.05, 276.35, 276.85, 277.65, 278.75, 278.15, 278.45, 
    277.85, 278.35, 278.15, 278.65, 278.05, 277.35, 279.05, 280.95, 280.65, 
    280.25, 279.25, 279.05, 279.65, 279.05, 278.15, 277.15, 276.75, 276.35, 
    277.05, 276.65, 277.35, 278.85, 279.95, 280.25, 281.55, 281.15, 280.85, 
    281.25, 281.45, 281.65, 282.75, 282.75, 282.45, 281.95, 280.75, 281.35, 
    281.35, 281.05, 280.75, 280.85, 280.45, 280.45, 280.35, 279.75, 280.15, 
    279.25, 279.35, 279.45, 278.85, 277.35, 277.75, 277.55, 277.25, 277.35, 
    277.15, 276.65, 276.55, 276.65, 276.25, 276.25, 276.25, 276.55, 276.45, 
    276.45, 276.55, 276.75, 276.65, 276.55, 276.75, 277.35, 277.55, 278.05, 
    278.15, 278.75, 279.15, 279.15, 279.35, 278.25, 278.75, 278.85, 278.35, 
    278.15, 278.25, 277.15, 276.85, 277.25, 277.25, 277.05, 278.55, 279.45, 
    280.95, 280.15, 279.55, 280.25, 279.05, 278.65, 280.05, 281.55, 281.75, 
    281.35, 281.15, 281.15, 280.05, 279.25, 278.65, 277.85, 277.75, 277.55, 
    277.75, 278.05, 277.85, 278.35, 277.55, 277.35, 276.85, 277.35, 277.85, 
    277.55, 277.55, 277.55, 278.45, 277.95, 277.55, 277.55, 278.05, 278.15, 
    278.35, 279.05, 279.05, 278.85, 278.85, 278.65, 278.65, 278.65, 278.45, 
    278.25, 278.25, 278.55, 279.15, 279.75, 279.85, 280.15, 280.45, 279.75, 
    280.15, 280.25, 279.95, 280.25, 279.75, 279.75, 279.55, 280.75, 280.85, 
    280.25, 280.05, 279.25, 279.05, 278.35, 278.15, 277.45, 277.25, 277.15, 
    277.75, 277.75, 278.55, 278.55, 278.45, 279.15, 278.85, 279.45, 278.65, 
    279.15, 278.35, 277.65, 279.65, 280.55, 280.55, 280.15, 281.35, 279.95, 
    279.05, 279.25, 279.35, 278.75, 279.65, 280.55, 280.15, 279.45, 279.65, 
    280.15, 280.75, 280.35, 278.95, 279.15, 279.75, 280.25, 279.55, 280.85, 
    282.35, 282.45, 283.05, 282.95, 283.75, 281.15, 281.95, 281.45, 282.05, 
    281.75, 281.35, 282.85, 280.85, 281.25, 280.45, 280.25, 279.85, 279.45, 
    279.45, 278.95, 279.35, 279.05, 279.15, 279.65, 279.75, 279.35, 279.85, 
    279.55, 279.55, 279.55, 279.35, 279.15, 279.15, 278.45, 278.45, 278.15, 
    277.95, 277.85, 278.15, 278.05, 277.75, 277.95, 277.95, 277.85, 278.55, 
    278.15, 278.25, 278.45, 278.15, 278.35, 278.95, 278.35, 278.25, 277.95, 
    278.35, 277.55, 277.55, 277.75, 278.05, 277.95, 277.95, 278.05, 278.05, 
    278.35, 278.55, 279.25, 279.35, 279.65, 279.85, 280.15, 279.95, 280.05, 
    280.45, 280.75, 280.75, 280.95, 280.95, 280.75, 280.65, 280.25, 279.85, 
    279.55, 279.25, 279.35, 279.75, 280.35, 280.45, 279.95, 279.25, 279.25, 
    279.95, 279.75, 279.65, 278.95, 279.55, 280.05, 279.75, 279.95, 279.95, 
    279.75, 279.75, 279.55, 279.45, 278.95, 278.75, 278.65, 278.35, 278.35, 
    278.25, 278.25, 278.45, 278.05, 278.75, 278.25, 278.05, 277.95, 278.95, 
    279.25, 278.45, 278.95, 278.95, 279.25, 279.15, 279.25, 278.55, 277.85, 
    277.85, 278.05, 278.15, 278.15, 278.25, 278.45, 278.25, 278.05, 277.75, 
    278.25, 278.35, 278.55, 278.95, 279.15, 279.75, 279.15, 280.15, 279.65, 
    279.75, 279.45, 279.25, 279.55, 278.75, 278.25, 278.05, 277.75, 277.85, 
    277.85, 277.85, 278.55, 278.65, 278.35, 279.15, 279.85, 279.55, 278.95, 
    279.65, 280.25, 279.65, 280.15, 280.65, 280.65, 279.65, 279.55, 278.25, 
    277.95, 277.55, 277.05, 277.25, 276.95, 276.65, 276.65, 276.45, 276.65, 
    276.95, 276.75, 277.15, 277.75, 278.25, 278.05, 277.65, 277.95, 278.35, 
    278.45, 278.45, 277.75, 277.45, 277.15, 276.85, 276.85, 276.85, 276.65, 
    276.75, 276.85, 277.25, 277.35, 277.75, 277.85, 278.15, 278.65, 278.75, 
    279.55, 279.65, 279.45, 279.25, 278.65, 278.65, 278.75, 278.55, 278.65, 
    278.75, 278.65, 278.45, 278.35, 278.15, 278.35, 278.35, 278.25, 278.35, 
    278.25, 278.05, 278.35, 278.35, 278.35, 278.65, 279.85, 280.75, 281.15, 
    280.95, 282.15, 281.05, 281.35, 282.15, 282.45, 281.55, 282.05, 283.55, 
    283.75, 284.15, 282.75, 282.05, 281.75, 282.55, 282.45, 281.45, 280.95, 
    280.05, 280.25, 280.65, 280.15, 280.45, 280.75, 280.95, 281.25, 279.85, 
    279.55, 279.65, 280.35, 280.15, 279.85, 279.65, 279.55, 279.15, 279.15, 
    279.95, 279.35, 279.55, 279.55, 279.25, 279.45, 279.25, 279.95, 279.55, 
    279.45, 279.55, 279.15, 279.05, 279.25, 279.45, 279.75, 280.35, 281.15, 
    281.05, 281.25, 281.75, 281.25, 280.15, 280.45, 280.25, 280.35, 280.15, 
    279.25, 279.05, 278.95, 278.85, 279.05, 279.65, 279.55, 279.35, 279.85, 
    280.25, 280.15, 280.55, 281.25, 281.75, 281.75, 282.05, 282.65, 282.95, 
    281.95, 281.75, 281.15, 280.95, 280.85, 280.95, 281.55, 282.15, 282.85, 
    283.15, 282.35, 281.95, 282.05, 282.65, 282.25, 282.55, 282.25, 282.95, 
    283.35, 281.95, 282.15, 282.05, 281.65, 281.15, 281.55, 281.65, 281.35, 
    281.25, 280.75, 282.45, 282.15, 282.05, 281.85, 282.15, 282.05, 282.65, 
    282.25, 282.45, 282.65, 283.15, 282.05, 281.75, 281.75, 280.85, 281.15, 
    280.55, 280.25, 280.05, 280.15, 279.55, 279.65, 279.65, 279.25, 279.15, 
    279.55, 279.35, 279.55, 279.25, 279.35, 279.35, 279.45, 279.85, 280.05, 
    279.65, 279.05, 279.25, 279.25, 279.45, 279.25, 279.35, 279.25, 279.45, 
    279.15, 279.25, 279.15, 279.25, 279.55, 278.85, 278.85, 278.75, 278.85, 
    279.05, 279.25, 279.25, 278.85, 279.45, 279.25, 279.15, 279.45, 279.55, 
    280.25, 280.55, 280.05, 279.95, 279.75, 279.65, 279.35, 279.15, 278.55, 
    278.55, 278.65, 278.25, 278.15, 277.95, 277.85, 277.85, 277.65, 278.05, 
    279.05, 278.75, 278.95, 279.25, 279.35, 278.95, 279.35, 279.45, 279.25, 
    279.35, 279.35, 279.15, 279.05, 278.85, 278.55, 278.35, 278.45, 278.15, 
    278.05, 278.25, 278.55, 278.35, 279.05, 278.75, 278.75, 279.05, 278.95, 
    279.45, 279.45, 278.75, 279.45, 280.05, 280.05, 279.45, 279.35, 279.25, 
    279.15, 278.95, 278.75, 278.55, 278.35, 278.35, 277.65, 277.65, 277.65, 
    277.75, 278.25, 278.75, 278.85, 278.75, 278.45, 278.55, 278.65, 279.35, 
    278.95, 278.15, 278.35, 278.45, 277.95, 278.65, 278.45, 278.35, 278.45, 
    278.45, 278.35, 278.35, 278.15, 278.35, 278.15, 278.05, 278.35, 278.35, 
    278.35, 278.55, 278.65, 278.65, 278.95, 279.05, 279.05, 279.45, 279.15, 
    279.45, 278.65, 279.05, 279.65, 279.65, 279.55, 279.25, 279.15, 279.15, 
    278.85, 278.85, 278.85, 278.95, 279.35, 279.65, 280.75, 280.85, 281.05, 
    281.65, 281.95, 282.35, 282.55, 282.55, 282.15, 282.25, 281.85, 281.85, 
    281.65, 281.45, 281.35, 280.85, 279.85, 279.35, 279.25, 279.25, 279.35, 
    279.75, 280.05, 281.15, 281.25, 281.55, 281.85, 282.15, 282.05, 282.25, 
    282.05, 281.75, 282.45, 281.25, 281.55, 281.35, 281.25, 281.25, 281.15, 
    280.85, 280.15, 279.75, 279.55, 279.55, 279.55, 279.35, 279.55, 279.65, 
    280.05, 279.95, 280.25, 280.45, 280.25, 280.25, 280.15, 280.25, 280.65, 
    280.65, 280.55, 280.35, 279.95, 279.45, 279.25, 279.35, 279.55, 279.25, 
    279.15, 279.15, 279.55, 279.85, 280.45, 280.45, 280.95, 281.55, 282.15, 
    281.85, 282.95, 282.15, 282.05, 282.45, 282.45, 282.45, 282.15, 281.95, 
    281.65, 281.25, 280.55, 280.65, 280.55, 280.45, 280.15, 280.15, 280.25, 
    280.35, 280.75, 281.65, 282.65, 281.65, 282.25, 283.25, 283.25, 283.05, 
    282.95, 283.65, 283.75, 282.45, 282.85, 281.75, 282.55, 282.05, 282.45, 
    282.05, 282.45, 282.25, 282.25, 282.05, 281.85, 282.05, 281.85, 282.35, 
    281.25, 281.05, 282.35, 281.75, 281.95, 282.85, 282.15, 281.35, 281.05, 
    281.65, 280.75, 280.95, 280.65, 280.65, 280.55, 280.05, 279.65, 280.05, 
    279.95, 279.85, 279.45, 279.35, 278.95, 279.05, 279.05, 279.25, 279.05, 
    279.35, 279.65, 279.55, 279.45, 279.25, 279.35, 279.05, 279.25, 279.35, 
    279.55, 279.55, 279.55, 279.45, 279.35, 279.15, 279.45, 279.65, 279.65, 
    279.55, 279.55, 279.75, 280.35, 280.75, 280.85, 282.15, 282.05, 282.15, 
    281.95, 282.05, 281.85, 282.25, 281.85, 282.25, 281.75, 281.55, 281.65, 
    281.35, 281.45, 280.85, 281.05, 281.05, 280.65, 280.95, 281.25, 280.65, 
    281.25, 281.65, 281.85, 282.05, 282.15, 282.25, 282.55, 282.55, 282.55, 
    282.25, 282.65, 283.35, 282.95, 282.95, 282.85, 282.45, 282.65, 282.55, 
    282.95, 282.45, 282.35, 282.05, 282.15, 281.45, 281.35, 281.85, 281.55, 
    281.35, 281.25, 280.45, 280.25, 280.15, 280.25, 280.15, 279.85, 279.45, 
    278.95, 279.05, 278.95, 278.95, 278.75, 278.35, 278.45, 278.45, 278.55, 
    278.85, 279.25, 279.15, 279.25, 279.45, 280.05, 279.45, 280.25, 280.45, 
    280.95, 280.95, 281.55, 281.45, 281.95, 282.55, 282.55, 282.25, 281.85, 
    282.35, 281.05, 280.85, 280.45, 280.55, 280.15, 280.25, 279.85, 280.85, 
    280.75, 279.65, 279.75, 279.45, 279.25, 280.45, 280.15, 280.05, 279.55, 
    279.45, 279.35, 278.95, 278.85, 278.95, 278.95, 278.85, 278.75, 279.05, 
    279.25, 279.25, 278.85, 278.85, 279.45, 279.35, 279.85, 280.35, 280.05, 
    280.35, 281.15, 280.45, 281.45, 281.35, 280.75, 280.35, 280.55, 280.05, 
    280.05, 280.25, 279.95, 279.65, 279.15, 279.15, 279.35, 278.55, 278.95, 
    278.75, 278.75, 279.25, 280.85, 280.95, 281.15, 281.25, 281.25, 281.65, 
    281.25, 281.35, 281.35, 281.05, 281.15, 281.05, 281.15, 280.85, 280.95, 
    281.85, 281.85, 281.05, 280.45, 280.15, 280.05, 280.15, 279.85, 280.05, 
    280.15, 280.45, 280.55, 280.75, 281.25, 281.55, 280.95, 282.05, 281.95, 
    281.45, 281.25, 280.75, 280.55, 280.45, 280.85, 280.25, 280.15, 280.25, 
    280.35, 280.15, 281.05, 279.55, 280.05, 280.95, 281.45, 281.15, 281.75, 
    282.15, 282.85, 283.25, 283.55, 283.35, 283.25, 283.35, 283.75, 284.05, 
    283.75, 282.15, 281.25, 281.35, 281.85, 281.65, 281.85, 281.65, 282.05, 
    282.45, 282.35, 282.15, 282.05, 282.45, 283.15, 283.65, 284.35, 284.15, 
    285.75, 285.55, 285.25, 285.55, 285.35, 285.25, 283.85, 284.15, 284.35, 
    283.35, 283.45, 283.05, 283.15, 283.35, 282.95, 282.45, 282.55, 282.05, 
    282.55, 283.95, 284.15, 284.05, 285.25, 285.25, 285.55, 286.25, 286.25, 
    285.55, 286.55, 286.45, 287.25, 285.15, 284.25, 285.25, 285.15, 285.45, 
    284.95, 284.75, 284.95, 284.95, 285.65, 286.15, 285.95, 286.15, 286.35, 
    286.15, 286.65, 285.85, 286.75, 286.85, 285.35, 284.45, 284.55, 283.85, 
    283.55, 283.45, 283.35, 283.35, 283.95, 282.95, 282.65, 282.75, 282.55, 
    281.75, 281.55, 281.75, 282.15, 282.15, 282.05, 282.15, 282.35, 281.85, 
    281.75, 281.85, 281.75, 281.45, 281.65, 281.85, 281.65, 281.45, 281.45, 
    280.85, 280.75, 280.75, 280.85, 280.55, 280.35, 280.35, 280.65, 281.35, 
    281.05, 281.05, 281.65, 281.45, 282.05, 281.85, 282.15, 282.75, 282.45, 
    282.15, 282.55, 282.15, 282.05, 281.75, 281.65, 282.05, 282.05, 281.65, 
    281.95, 281.25, 282.05, 281.95, 281.85, 282.15, 282.45, 282.35, 282.65, 
    282.85, 283.15, 283.45, 284.15, 282.75, 283.05, 283.65, 283.25, 282.75, 
    282.35, 282.05, 281.65, 281.15, 280.65, 280.55, 280.35, 281.05, 281.65, 
    282.45, 283.05, 283.95, 283.95, 283.85, 284.25, 283.75, 283.75, 282.95, 
    282.15, 282.65, 283.25, 282.85, 282.35, 281.85, 281.45, 282.05, 282.15, 
    281.05, 281.65, 280.95, 280.65, 282.05, 281.85, 281.25, 280.75, 281.45, 
    281.05, 282.25, 280.75, 282.45, 282.65, 282.75, 281.15, 280.35, 280.75, 
    281.05, 280.55, 280.25, 279.45, 280.85, 280.85, 280.45, 279.35, 279.75, 
    280.15, 279.75, 280.15, 279.75, 280.25, 281.15, 280.75, 280.85, 280.75, 
    280.75, 280.65, 281.05, 281.45, 281.75, 281.85, 282.35, 282.05, 279.85, 
    280.15, 279.85, 279.45, 279.35, 279.25, 279.45, 279.85, 279.55, 279.25, 
    279.15, 278.95, 279.05, 279.15, 279.25, 279.45, 279.65, 279.55, 279.95, 
    279.95, 280.25, 280.65, 280.45, 280.25, 280.45, 280.25, 280.05, 279.85, 
    279.95, 279.75, 279.65, 278.85, 278.65, 278.25, 278.35, 278.65, 278.65, 
    278.85, 279.25, 279.65, 279.65, 280.05, 279.65, 279.95, 280.25, 280.15, 
    280.05, 280.15, 280.25, 280.05, 280.25, 279.95, 279.65, 279.25, 278.95, 
    279.05, 279.05, 279.55, 279.15, 279.05, 278.95, 278.95, 279.25, 279.35, 
    279.45, 279.55, 279.85, 279.85, 279.65, 279.85, 279.95, 280.25, 279.75, 
    280.35, 280.45, 280.45, 280.45, 280.25, 280.15, 279.95, 279.75, 279.65, 
    279.65, 279.55, 279.55, 279.85, 280.05, 280.25, 280.45, 280.65, 280.75, 
    281.25, 281.85, 281.65, 281.15, 280.85, 280.75, 280.45, 279.85, 279.65, 
    279.25, 278.95, 278.75, 278.85, 279.05, 278.75, 279.05, 279.55, 280.25, 
    281.05, 281.55, 281.45, 281.85, 281.95, 281.95, 281.75, 282.15, 281.95, 
    281.95, 281.85, 281.55, 281.35, 280.45, 279.85, 279.35, 278.15, 277.95, 
    277.95, 277.65, 277.25, 277.95, 278.55, 278.85, 278.55, 278.45, 278.75, 
    278.85, 278.75, 278.95, 279.15, 278.95, 278.95, 278.95, 278.95, 278.75, 
    278.65, 278.55, 278.25, 278.05, 277.95, 277.75, 277.75, 277.65, 277.65, 
    277.55, 277.55, 277.95, 277.65, 277.75, 277.75, 277.95, 278.25, 278.65, 
    279.35, 279.25, 279.05, 279.55, 279.95, 279.95, 279.85, 279.75, 279.65, 
    279.65, 279.45, 279.15, 278.65, 278.65, 279.05, 279.25, 279.05, 279.15, 
    279.15, 279.25, 279.65, 279.75, 279.75, 279.95, 280.55, 280.45, 280.15, 
    280.35, 280.65, 280.35, 280.15, 279.85, 279.55, 279.15, 279.15, 279.35, 
    279.85, 279.95, 279.95, 279.75, 280.05, 280.25, 280.95, 281.05, 280.55, 
    280.35, 280.65, 280.65, 280.85, 280.75, 280.05, 280.05, 280.05, 280.05, 
    279.65, 279.65, 281.05, 281.85, 282.55, 283.35, 282.75, 283.35, 283.55, 
    283.25, 283.45, 283.35, 282.55, 279.75, 279.05, 278.85, 278.65, 278.55, 
    278.45, 278.45, 278.95, 278.35, 277.85, 277.65, 277.55, 277.45, 277.35, 
    277.15, 276.95, 276.95, 276.95, 276.75, 276.75, 276.95, 277.15, 277.45, 
    277.55, 277.75, 277.95, 278.45, 279.35, 279.95, 279.35, 278.65, 278.65, 
    278.75, 279.15, 279.25, 279.15, 279.05, 278.85, 278.95, 278.75, 278.55, 
    278.45, 278.35, 278.55, 278.55, 278.65, 279.15, 280.35, 280.25, 280.45, 
    281.25, 281.15, 281.25, 281.25, 281.25, 280.65, 280.45, 280.35, 280.35, 
    280.35, 279.75, 279.25, 278.85, 278.65, 280.55, 279.75, 279.35, 280.15, 
    280.35, 280.75, 280.55, 280.55, 280.85, 280.15, 281.15, 281.95, 281.45, 
    280.85, 280.25, 279.45, 279.05, 278.45, 278.95, 278.55, 278.25, 278.25, 
    277.95, 278.25, 277.95, 277.85, 277.95, 277.95, 277.95, 277.95, 278.15, 
    278.55, 279.45, 279.45, 279.05, 279.45, 279.95, 279.95, 279.75, 279.75, 
    279.35, 279.25, 279.15, 278.65, 278.55, 278.65, 278.35, 277.95, 277.75, 
    278.25, 278.25, 277.95, 278.45, 278.25, 278.75, 278.45, 278.75, 278.65, 
    279.05, 279.45, 279.45, 279.25, 279.55, 280.15, 280.15, 280.35, 280.25, 
    279.45, 279.45, 279.55, 279.95, 279.65, 278.85, 279.15, 278.85, 278.35, 
    278.25, 278.85, 278.55, 278.85, 279.05, 279.45, 279.65, 279.65, 279.55, 
    279.45, 279.25, 279.25, 279.25, 278.85, 278.75, 278.45, 278.45, 277.75, 
    277.55, 277.45, 277.35, 276.75, 277.25, 276.95, 277.05, 277.55, 278.05, 
    278.05, 278.15, 278.85, 278.55, 278.65, 278.35, 277.65, 277.35, 277.35, 
    277.25, 277.05, 276.95, 277.15, 277.15, 277.15, 277.15, 277.25, 276.35, 
    276.35, 277.05, 276.35, 277.15, 277.05, 277.15, 277.55, 277.95, 278.05, 
    277.75, 277.95, 277.95, 278.05, 277.95, 277.85, 277.85, 277.75, 277.65, 
    277.25, 276.95, 276.25, 275.65, 276.05, 275.55, 275.55, 275.35, 275.75, 
    276.05, 276.25, 276.85, 277.05, 277.45, 277.95, 277.95, 277.85, 278.05, 
    278.05, 277.95, 277.85, 277.85, 277.75, 277.55, 277.35, 277.15, 276.35, 
    276.35, 276.15, 275.75, 276.05, 275.55, 275.05, 276.55, 276.55, 277.95, 
    276.95, 277.35, 277.65, 277.45, 277.95, 278.65, 279.05, 279.55, 279.15, 
    278.65, 278.05, 278.15, 277.75, 277.55, 277.25, 276.95, 276.75, 276.65, 
    276.45, 276.25, 276.65, 277.05, 276.75, 277.45, 277.55, 277.65, 277.45, 
    277.15, 277.15, 277.15, 277.85, 277.75, 277.95, 278.35, 278.85, 278.85, 
    278.55, 278.55, 278.85, 278.95, 279.25, 279.45, 278.95, 278.95, 278.85, 
    279.15, 279.25, 280.05, 279.65, 281.15, 280.45, 281.25, 282.05, 283.15, 
    283.55, 282.95, 283.35, 283.75, 280.65, 279.75, 280.05, 279.95, 279.95, 
    280.25, 280.55, 279.85, 278.65, 278.75, 278.45, 278.25, 278.25, 278.45, 
    278.65, 278.75, 278.45, 279.05, 278.85, 278.75, 279.35, 278.65, 278.55, 
    278.25, 278.15, 277.25, 277.35, 276.55, 276.95, 275.85, 275.75, 276.55, 
    276.05, 275.65, 274.55, 274.45, 274.85, 274.95, 275.55, 276.35, 277.15, 
    277.55, 278.15, 278.05, 277.95, 277.65, 278.45, 278.75, 278.75, 278.95, 
    278.75, 279.05, 278.65, 279.15, 278.85, 278.85, 279.65, 279.85, 280.05, 
    279.15, 280.45, 280.05, 280.05, 280.95, 280.55, 280.05, 280.45, 280.35, 
    280.55, 279.75, 279.75, 279.25, 279.05, 279.15, 279.85, 279.05, 278.75, 
    278.85, 278.45, 278.15, 278.15, 278.35, 278.05, 277.25, 277.75, 278.55, 
    278.25, 279.75, 280.75, 281.25, 281.15, 282.15, 281.55, 281.35, 281.15, 
    280.85, 280.05, 279.85, 279.85, 279.05, 278.55, 278.45, 278.35, 277.35, 
    277.55, 276.85, 277.05, 277.55, 277.55, 277.55, 277.95, 278.25, 278.95, 
    279.25, 278.85, 278.85, 279.25, 278.75, 278.55, 279.15, 279.65, 278.95, 
    278.55, 278.55, 278.35, 278.35, 278.35, 278.45, 278.05, 278.15, 278.25, 
    277.55, 277.45, 277.65, 277.85, 277.75, 277.55, 278.45, 279.05, 279.35, 
    278.85, 279.15, 279.35, 279.05, 278.85, 278.75, 279.15, 278.55, 278.25, 
    277.75, 277.55, 277.55, 276.65, 275.95, 275.75, 275.55, 275.85, 276.25, 
    276.45, 276.65, 277.55, 276.85, 277.25, 276.75, 276.35, 276.75, 276.05, 
    276.65, 276.85, 276.35, 275.85, 275.45, 274.95, 274.65, 275.25, 275.05, 
    274.45, 274.05, 274.15, 274.15, 274.25, 274.15, 274.95, 274.95, 274.65, 
    275.75, 276.95, 277.05, 277.45, 277.75, 277.55, 277.35, 277.35, 277.15, 
    276.95, 276.85, 276.45, 276.65, 276.85, 276.75, 276.65, 276.25, 275.95, 
    275.65, 275.65, 276.05, 276.65, 276.65, 276.55, 276.45, 276.25, 276.25, 
    276.55, 276.35, 276.45, 277.35, 278.05, 277.65, 277.35, 276.75, 277.05, 
    277.15, 277.55, 277.25, 276.95, 277.35, 276.85, 277.95, 278.05, 278.25, 
    278.15, 278.75, 278.65, 278.65, 278.95, 279.05, 278.95, 279.25, 279.15, 
    279.05, 278.95, 278.85, 278.75, 278.65, 278.55, 277.95, 277.95, 277.75, 
    277.55, 277.65, 278.35, 277.55, 277.65, 278.45, 278.15, 278.35, 278.75, 
    278.55, 278.65, 278.75, 278.75, 278.25, 278.25, 278.25, 278.15, 278.05, 
    277.65, 277.55, 276.95, 276.65, 276.25, 275.55, 275.35, 275.55, 275.45, 
    276.55, 278.05, 278.85, 279.25, 279.75, 279.45, 279.95, 279.95, 279.95, 
    279.55, 279.55, 279.15, 278.65, 278.35, 277.75, 277.35, 277.25, 277.05, 
    276.85, 276.65, 276.45, 276.55, 276.35, 275.85, 276.25, 276.75, 276.85, 
    276.65, 278.15, 277.75, 278.15, 277.65, 278.65, 278.05, 277.95, 277.55, 
    277.05, 276.35, 276.35, 276.15, 275.65, 275.15, 274.95, 274.55, 274.15, 
    274.15, 273.05, 272.15, 272.05, 272.95, 273.05, 273.85, 274.65, 274.95, 
    274.75, 274.65, 274.65, 274.65, 274.75, 274.65, 274.35, 274.55, 274.35, 
    274.25, 273.75, 273.85, 273.65, 272.85, 272.85, 273.25, 273.15, 273.75, 
    274.35, 274.25, 274.05, 273.95, 273.95, 274.05, 274.25, 274.35, 274.25, 
    274.65, 274.65, 274.75, 274.55, 274.25, 274.35, 274.35, 274.25, 273.95, 
    273.95, 273.55, 273.35, 273.15, 273.35, 272.95, 272.95, 273.15, 273.15, 
    272.95, 272.95, 273.25, 273.55, 274.05, 273.75, 273.95, 274.65, 274.05, 
    273.75, 272.55, 271.35, 271.55, 271.25, 271.65, 271.65, 271.25, 270.95, 
    269.85, 270.85, 270.55, 270.95, 271.25, 272.05, 272.85, 273.95, 274.35, 
    274.25, 275.05, 275.05, 275.55, 275.35, 275.05, 273.15, 274.95, 273.35, 
    273.55, 273.75, 272.55, 273.15, 273.45, 272.55, 273.25, 273.05, 272.35, 
    272.75, 274.15, 271.95, 273.55, 275.05, 275.45, 276.25, 276.15, 276.25, 
    276.35, 275.85, 275.85, 275.65, 275.05, 275.45, 275.15, 275.05, 274.55, 
    272.55, 272.55, 271.15, 272.05, 271.75, 271.15, 272.25, 271.85, 271.85, 
    272.35, 271.85, 273.05, 273.15, 273.65, 275.15, 273.75, 273.65, 273.55, 
    273.15, 272.45, 272.05, 271.25, 270.65, 270.25, 270.15, 270.55, 270.65, 
    269.95, 269.95, 269.95, 269.85, 269.75, 270.05, 271.15, 271.75, 272.25, 
    272.95, 273.45, 274.15, 273.75, 273.85, 273.75, 273.45, 273.05, 273.35, 
    271.25, 271.75, 270.65, 270.55, 273.75, 273.65, 273.75, 274.05, 273.85, 
    273.75, 274.15, 274.65, 274.65, 274.55, 274.55, 274.75, 274.45, 274.25, 
    274.25, 274.25, 273.85, 273.25, 273.25, 273.25, 273.25, 273.05, 272.95, 
    273.25, 272.95, 273.05, 273.15, 273.25, 273.35, 273.75, 273.25, 273.15, 
    273.65, 273.75, 273.95, 274.45, 274.55, 274.65, 274.65, 274.45, 274.25, 
    274.45, 274.05, 273.85, 273.45, 273.75, 272.05, 270.85, 271.45, 270.65, 
    270.25, 270.55, 271.45, 271.35, 272.65, 273.65, 274.35, 275.05, 275.05, 
    274.85, 275.05, 275.05, 275.25, 275.75, 275.45, 275.35, 274.95, 274.35, 
    274.65, 274.05, 273.95, 274.65, 275.05, 274.95, 274.35, 274.55, 274.95, 
    275.05, 275.95, 275.75, 276.25, 276.75, 277.25, 277.05, 276.75, 277.05, 
    277.05, 277.05, 277.35, 277.65, 277.85, 277.55, 278.35, 278.35, 278.65, 
    278.45, 279.15, 279.25, 279.75, 278.75, 279.05, 278.65, 278.95, 278.05, 
    277.85, 277.65, 276.95, 277.25, 277.45, 277.95, 277.85, 277.95, 277.35, 
    277.25, 276.55, 276.35, 276.05, 275.45, 275.65, 275.55, 275.45, 275.35, 
    275.45, 275.15, 275.45, 275.55, 275.55, 275.45, 275.45, 275.15, 275.15, 
    275.35, 275.25, 275.15, 274.95, 274.75, 273.75, 273.65, 273.45, 273.05, 
    272.95, 272.75, 272.45, 272.15, 272.05, 271.95, 271.65, 271.55, 271.05, 
    271.05, 270.95, 270.85, 270.75, 270.75, 270.85, 271.05, 270.45, 270.55, 
    270.45, 270.35, 270.25, 270.05, 269.75, 268.15, 267.85, 268.15, 267.45, 
    267.05, 267.25, 266.75, 266.85, 266.85, 267.25, 267.35, 266.65, 267.35, 
    266.95, 267.75, 268.45, 268.65, 268.85, 268.85, 268.75, 269.05, 269.15, 
    269.35, 268.65, 268.55, 268.35, 268.95, 268.45, 268.75, 268.65, 268.65, 
    269.05, 268.65, 268.35, 268.65, 268.35, 268.15, 268.05, 268.35, 268.85, 
    269.55, 269.55, 268.85, 268.55, 268.55, 268.75, 267.85, 268.45, 268.45, 
    268.85, 268.75, 268.85, 269.35, 269.25, 269.55, 269.95, 269.85, 269.45, 
    269.05, 268.35, 267.45, 267.35, 267.55, 268.15, 269.15, 269.75, 268.75, 
    268.75, 267.45, 267.85, 267.85, 267.45, 266.85, 266.65, 265.95, 265.65, 
    265.45, 266.95, 266.05, 265.75, 265.65, 266.15, 266.25, 266.15, 265.85, 
    266.05, 266.45, 266.55, 266.25, 266.75, 265.65, 266.45, 266.35, 265.25, 
    265.75, 265.35, 264.95, 264.95, 264.85, 264.05, 264.15, 264.45, 264.55, 
    263.65, 265.15, 264.55, 265.05, 265.75, 266.15, 268.25, 267.75, 268.85, 
    269.55, 270.25, 269.85, 270.25, 270.95, 270.55, 271.35, 272.15, 272.25, 
    272.55, 272.85, 272.55, 272.95, 273.15, 273.25, 273.05, 273.15, 272.75, 
    272.75, 272.85, 273.05, 272.25, 272.05, 272.55, 272.15, 272.35, 272.65, 
    273.55, 273.85, 273.35, 273.35, 273.55, 273.35, 273.25, 273.05, 273.25, 
    273.35, 273.45, 273.45, 273.35, 273.25, 271.45, 270.45, 270.75, 270.45, 
    270.95, 271.05, 273.95, 272.25, 272.55, 273.25, 273.55, 272.65, 273.05, 
    272.35, 272.95, 271.95, 273.85, 271.05, 271.35, 272.55, 272.55, 272.15, 
    272.55, 272.55, 271.85, 270.95, 270.75, 271.45, 271.75, 270.55, 269.65, 
    269.35, 270.45, 268.45, 268.75, 267.85, 267.45, 267.75, 267.05, 267.05, 
    267.45, 268.45, 268.85, 268.65, 268.45, 268.25, 268.05, 268.05, 267.95, 
    267.75, 267.65, 267.45, 267.25, 267.45, 267.45, 267.55, 267.85, 267.95, 
    267.85, 267.95, 267.65, 267.05, 267.35, 267.65, 267.65, 267.65, 267.75, 
    267.85, 267.95, 268.05, 268.15, 267.05, 267.55, 267.75, 268.25, 268.55, 
    268.45, 268.65, 269.15, 267.75, 266.95, 268.35, 266.05, 265.75, 265.85, 
    266.65, 265.75, 266.95, 267.55, 267.75, 268.05, 268.25, 268.25, 268.25, 
    268.45, 268.25, 268.25, 266.15, 268.05, 267.35, 266.55, 265.55, 267.15, 
    267.35, 267.95, 267.85, 267.95, 269.15, 267.25, 268.45, 268.15, 268.05, 
    267.25, 265.75, 267.05, 266.05, 267.65, 267.75, 267.55, 267.35, 266.45, 
    267.85, 267.25, 265.15, 265.55, 266.85, 266.05, 265.05, 265.75, 266.45, 
    266.25, 265.75, 265.05, 265.85, 265.55, 264.25, 264.55, 264.95, 264.75, 
    264.85, 265.15, 265.35, 264.25, 264.45, 263.55, 264.85, 266.55, 266.75, 
    266.95, 266.85, 267.25, 267.75, 267.85, 267.55, 267.05, 266.05, 265.45, 
    266.15, 265.65, 265.45, 266.35, 266.95, 266.45, 265.15, 265.45, 265.35, 
    265.45, 266.95, 267.15, 265.45, 265.65, 264.45, 265.25, 265.85, 265.45, 
    267.15, 266.75, 264.35, 262.85, 265.05, 264.65, 264.95, 265.45, 263.05, 
    264.85, 264.85, 264.55, 264.15, 264.85, 265.55, 265.85, 266.95, 266.55, 
    266.75, 266.55, 267.15, 267.55, 267.25, 266.25, 267.85, 267.75, 268.65, 
    269.15, 269.15, 269.15, 269.75, 269.35, 269.25, 269.75, 270.35, 270.55, 
    270.75, 270.75, 271.05, 271.55, 272.05, 271.65, 271.65, 271.25, 271.25, 
    271.55, 271.35, 271.65, 271.75, 272.05, 272.85, 272.65, 272.45, 272.35, 
    272.55, 272.55, 272.85, 273.35, 274.05, 274.35, 274.35, 274.45, 274.65, 
    275.55, 274.35, 274.05, 274.55, 275.65, 275.15, 275.55, 276.25, 276.75, 
    276.35, 276.35, 277.05, 277.55, 277.75, 277.35, 277.25, 276.55, 276.35, 
    276.95, 276.15, 276.45, 277.35, 276.55, 276.55, 276.75, 276.95, 276.95, 
    277.15, 276.85, 277.05, 277.35, 279.35, 279.45, 280.75, 280.05, 279.05, 
    278.35, 278.55, 277.55, 278.25, 277.75, 276.75, 275.75, 275.25, 275.45, 
    275.25, 276.05, 274.85, 274.95, 274.75, 275.05, 275.25, 275.25, 275.15, 
    275.55, 275.55, 275.65, 275.25, 276.05, 275.95, 275.45, 275.15, 274.75, 
    274.75, 274.45, 274.55, 274.65, 274.75, 274.55, 274.05, 274.65, 275.65, 
    274.65, 274.75, 274.25, 275.25, 276.55, 275.25, 275.45, 274.75, 274.85, 
    275.15, 275.25, 275.25, 275.05, 274.25, 274.45, 274.25, 274.45, 274.05, 
    273.75, 273.65, 273.75, 273.55, 273.25, 273.05, 273.25, 273.05, 273.15, 
    272.85, 273.05, 272.55, 272.75, 272.85, 272.75, 272.85, 272.45, 272.45, 
    272.35, 271.05, 271.65, 271.25, 270.85, 270.85, 270.45, 270.75, 270.85, 
    270.45, 270.45, 269.65, 269.95, 269.75, 269.55, 270.25, 270.25, 270.55, 
    270.45, 270.45, 271.15, 271.35, 270.45, 271.05, 270.35, 270.55, 270.15, 
    269.45, 269.45, 268.85, 269.55, 268.25, 269.05, 268.35, 268.45, 268.15, 
    268.65, 268.25, 267.85, 267.35, 268.35, 267.75, 266.95, 267.35, 267.85, 
    267.55, 267.05, 267.75, 267.85, 266.95, 267.05, 267.35, 266.45, 266.45, 
    265.95, 266.55, 265.95, 266.25, 266.15, 266.85, 266.65, 266.25, 266.05, 
    267.45, 266.35, 267.05, 267.35, 267.25, 268.25, 268.35, 268.45, 269.05, 
    269.45, 269.55, 269.55, 270.55, 274.65, 275.15, 275.45, 275.75, 276.45, 
    276.95, 277.05, 276.85, 276.55, 276.75, 276.95, 277.15, 276.65, 277.05, 
    277.05, 277.15, 277.05, 277.25, 277.25, 276.85, 276.85, 277.05, 276.75, 
    277.25, 277.05, 277.15, 277.15, 276.75, 276.95, 277.25, 277.75, 277.85, 
    277.65, 277.55, 278.35, 278.75, 277.65, 278.55, 277.65, 277.35, 277.55, 
    277.55, 277.55, 277.55, 277.55, 277.55, 277.85, 277.55, 277.35, 277.05, 
    277.15, 277.05, 277.25, 277.25, 276.65, 276.25, 276.15, 276.15, 276.15, 
    276.25, 276.05, 275.85, 275.65, 275.55, 275.35, 274.85, 274.25, 274.75, 
    273.75, 273.75, 273.25, 273.35, 273.15, 273.45, 273.45, 273.45, 273.25, 
    272.85, 272.85, 272.75, 272.85, 273.05, 272.65, 272.65, 272.55, 272.15, 
    272.15, 272.15, 272.25, 272.65, 272.65, 272.75, 272.65, 272.55, 272.75, 
    272.55, 272.45, 272.75, 272.35, 272.25, 272.05, 272.05, 271.95, 272.15, 
    272.15, 272.15, 272.25, 272.15, 272.05, 271.85, 271.95, 272.15, 272.15, 
    272.05, 271.65, 270.85, 270.85, 270.75, 269.95, 269.95, 268.45, 271.25, 
    271.05, 271.65, 271.65, 271.65, 271.55, 271.55, 271.85, 271.75, 271.55, 
    271.35, 270.85, 270.85, 270.45, 270.15, 269.75, 269.85, 269.65, 269.65, 
    269.25, 269.25, 268.95, 268.75, 267.35, 267.35, 266.85, 267.35, 266.35, 
    268.75, 268.65, 268.05, 267.65, 267.15, 267.55, 267.45, 267.45, 266.85, 
    267.75, 267.35, 266.65, 266.05, 266.95, 266.55, 265.85, 265.45, 265.05, 
    264.85, 264.95, 264.85, 264.95, 264.65, 264.95, 265.25, 265.45, 265.65, 
    265.55, 265.75, 265.85, 265.25, 264.55, 264.05, 263.75, 263.65, 263.75, 
    263.15, 263.65, 264.65, 265.35, 266.15, 266.45, 267.45, 267.85, 267.45, 
    268.05, 268.75, 268.65, 268.35, 268.45, 269.55, 269.65, 270.65, 271.25, 
    271.45, 271.15, 272.45, 272.05, 272.95, 271.95, 272.35, 272.25, 272.05, 
    272.25, 272.15, 272.95, 272.15, 274.75, 274.25, 271.75, 271.15, 270.85, 
    270.35, 270.55, 269.85, 268.85, 267.85, 268.05, 267.95, 267.85, 265.85, 
    266.15, 265.55, 265.75, 265.45, 266.05, 266.35, 265.65, 266.45, 267.65, 
    268.25, 269.45, 270.05, 271.45, 271.45, 271.35, 271.35, 270.85, 271.25, 
    271.05, 270.95, 270.85, 270.75, 270.85, 270.85, 271.05, 271.35, 271.15, 
    271.35, 271.25, 271.25, 271.25, 272.15, 272.05, 271.95, 271.85, 272.05, 
    272.05, 272.05, 271.95, 272.15, 272.25, 271.95, 272.05, 271.95, 272.65, 
    272.85, 273.15, 272.95, 272.75, 272.55, 272.65, 272.25, 272.25, 272.05, 
    271.85, 271.65, 271.55, 271.55, 271.75, 271.45, 271.65, 271.45, 271.45, 
    271.25, 271.15, 271.25, 271.15, 271.15, 270.65, 270.45, 270.25, 270.15, 
    269.95, 269.65, 269.45, 269.15, 268.75, 268.95, 268.85, 268.65, 268.65, 
    268.35, 268.15, 267.65, 267.25, 266.95, 266.65, 266.75, 266.75, 266.45, 
    267.05, 267.15, 267.45, 267.55, 267.35, 267.65, 267.55, 267.75, 267.35, 
    267.85, 266.85, 265.95, 266.25, 266.05, 266.35, 268.55, 268.85, 267.85, 
    267.35, 265.65, 267.35, 268.95, 267.35, 267.75, 270.75, 271.25, 271.95, 
    272.65, 273.25, 273.85, 274.25, 274.05, 274.25, 274.55, 274.25, 274.05, 
    274.15, 274.35, 274.55, 275.05, 275.35, 275.45, 275.55, 275.85, 275.35, 
    276.45, 275.85, 276.05, 276.55, 276.35, 276.45, 275.55, 275.45, 275.05, 
    274.65, 274.05, 274.05, 273.75, 273.75, 273.85, 273.45, 273.25, 272.85, 
    272.75, 272.55, 272.15, 271.95, 272.15, 271.95, 271.75, 271.85, 271.85, 
    271.75, 271.55, 271.05, 271.35, 270.95, 271.55, 271.25, 271.05, 270.85, 
    270.65, 270.65, 270.45, 270.55, 270.95, 270.55, 270.75, 270.55, 270.55, 
    270.25, 269.85, 269.85, 269.65, 269.65, 269.75, 269.85, 269.85, 269.55, 
    270.85, 271.25, 271.75, 272.35, 272.85, 272.35, 271.85, 271.85, 271.95, 
    271.95, 270.75, 270.45, 270.65, 270.65, 270.65, 270.45, 270.35, 270.35, 
    270.75, 270.95, 271.35, 270.95, 270.95, 271.45, 271.35, 270.75, 270.15, 
    270.35, 269.95, 269.75, 269.85, 268.45, 268.25, 268.65, 268.65, 269.15, 
    269.25, 268.95, 269.75, 269.65, 269.05, 269.45, 269.25, 269.75, 270.15, 
    270.55, 270.85, 270.85, 270.45, 270.55, 271.05, 271.35, 271.95, 271.85, 
    271.65, 272.05, 272.05, 272.05, 272.45, 272.05, 272.45, 272.85, 272.45, 
    273.15, 272.85, 272.85, 273.05, 273.15, 272.75, 272.25, 272.55, 272.85, 
    272.95, 273.45, 273.25, 273.05, 273.15, 274.25, 273.75, 273.25, 273.65, 
    273.45, 273.85, 273.25, 273.15, 273.25, 273.95, 274.65, 274.35, 274.25, 
    274.45, 274.55, 275.75, 275.65, 275.45, 275.15, 274.95, 274.75, 274.45, 
    274.65, 274.35, 273.85, 274.85, 274.25, 273.85, 273.15, 272.45, 270.95, 
    270.35, 269.45, 268.15, 267.65, 267.05, 267.75, 266.15, 266.75, 266.15, 
    265.45, 265.55, 265.65, 265.55, 265.15, 264.35, 264.75, 263.85, 265.15, 
    264.85, 265.25, 264.55, 264.85, 264.45, 264.75, 265.35, 264.75, 264.35, 
    264.75, 264.85, 264.65, 264.85, 265.05, 265.15, 265.05, 265.45, 266.55, 
    264.15, 264.35, 264.65, 264.75, 264.75, 264.05, 264.55, 264.95, 264.85, 
    263.65, 264.15, 264.85, 264.45, 264.45, 264.85, 265.15, 265.35, 265.55, 
    265.45, 265.45, 265.45, 265.45, 265.75, 265.75, 265.75, 265.75, 265.85, 
    265.75, 265.65, 265.85, 266.15, 266.15, 266.45, 266.55, 266.95, 267.35, 
    267.85, 267.75, 267.85, 267.35, 266.45, 267.45, 267.85, 267.65, 268.05, 
    268.55, 268.65, 269.15, 268.45, 268.75, 269.05, 268.85, 268.55, 267.85, 
    267.35, 266.65, 265.85, 265.75, 264.95, 264.65, 264.05, 263.65, 263.25, 
    263.45, 263.25, 263.15, 263.15, 263.15, 262.95, 262.85, 262.65, 262.95, 
    262.65, 262.45, 263.15, 263.05, 262.95, 262.65, 261.55, 260.55, 259.65, 
    259.55, 259.35, 259.95, 261.05, 262.15, 261.75, 262.25, 262.95, 263.25, 
    263.75, 263.25, 264.05, 263.55, 263.95, 264.05, 264.65, 264.85, 265.55, 
    265.75, 266.35, 266.45, 267.05, 266.95, 266.85, 268.85, 268.55, 269.05, 
    269.15, 269.35, 270.35, 271.75, 272.25, 272.95, 274.05, 275.85, 275.55, 
    275.25, 276.05, 275.25, 275.35, 275.55, 275.45, 274.65, 276.05, 276.15, 
    276.65, 277.05, 276.65, 276.65, 276.35, 276.25, 276.45, 276.45, 276.65, 
    275.85, 277.05, 276.05, 277.55, 276.95, 276.35, 276.35, 276.85, 277.95, 
    276.65, 276.65, 275.85, 275.45, 275.35, 274.75, 273.75, 272.95, 272.55, 
    271.95, 271.25, 271.25, 269.75, 270.45, 270.25, 270.65, 270.15, 268.05, 
    267.25, 267.05, 266.45, 266.15, 266.05, 265.15, 264.65, 264.75, 263.85, 
    263.85, 263.65, 262.75, 262.75, 262.15, 261.45, 261.15, 261.05, 261.35, 
    262.15, 262.55, 262.95, 262.95, 262.95, 262.95, 262.75, 262.65, 263.05, 
    263.25, 264.15, 264.45, 264.15, 262.65, 262.15, 263.65, 264.35, 264.55, 
    264.45, 263.75, 264.05, 262.95, 264.15, 263.45, 262.75, 262.85, 262.15, 
    262.05, 262.15, 261.55, 262.25, 262.35, 262.05, 261.95, 262.55, 262.15, 
    263.05, 263.35, 264.75, 265.25, 265.75, 266.15, 266.95, 267.25, 266.75, 
    267.05, 267.15, 267.35, 268.65, 269.35, 269.65, 272.05, 271.95, 272.25, 
    272.45, 272.75, 272.55, 272.65, 272.75, 272.95, 272.95, 272.15, 272.15, 
    271.85, 271.65, 271.55, 270.95, 271.05, 270.45, 270.75, 270.45, 269.95, 
    269.95, 269.75, 269.75, 269.65, 269.05, 267.95, 267.75, 268.35, 267.95, 
    268.35, 267.85, 267.95, 266.55, 267.35, 267.15, 267.35, 267.25, 266.95, 
    266.75, 266.45, 266.15, 266.25, 264.75, 266.15, 265.95, 265.25, 265.55, 
    264.55, 265.75, 265.55, 265.55, 265.15, 264.85, 263.75, 263.25, 263.25, 
    263.45, 262.75, 263.45, 262.95, 263.25, 263.25, 264.85, 263.15, 262.95, 
    262.75, 261.95, 262.95, 262.25, 261.95, 261.75, 262.05, 261.45, 261.35, 
    260.85, 260.95, 260.65, 262.55, 262.15, 260.95, 261.65, 261.95, 261.45, 
    261.25, 261.15, 261.35, 261.25, 261.25, 260.45, 260.55, 260.85, 260.45, 
    261.05, 261.65, 260.75, 262.05, 262.55, 261.95, 263.35, 263.55, 263.55, 
    263.75, 264.25, 265.25, 264.65, 267.95, 269.45, 270.05, 270.55, 269.85, 
    271.05, 272.15, 269.35, 266.85, 265.95, 265.45, 265.15, 265.05, 264.65, 
    264.55, 264.65, 264.85, 265.05, 264.25, 264.75, 263.65, 261.35, 261.75, 
    261.35, 260.75, 260.85, 262.05, 257.85, 261.95, 261.65, 266.25, 266.95, 
    267.55, 267.05, 267.75, 269.55, 269.05, 268.95, 269.25, 269.25, 268.55, 
    266.85, 267.75, 267.55, 268.05, 270.75, 270.65, 270.45, 270.75, 271.05, 
    271.05, 270.85, 270.55, 270.45, 270.25, 270.05, 270.15, 269.55, 270.15, 
    269.85, 269.65, 269.55, 269.75, 269.55, 270.15, 270.05, 270.25, 270.25, 
    270.45, 270.15, 270.35, 270.55, 270.65, 270.75, 270.95, 271.05, 271.15, 
    270.85, 270.95, 270.05, 270.45, 271.05, 270.35, 270.65, 270.85, 271.25, 
    271.15, 270.55, 270.95, 270.55, 270.15, 269.95, 269.85, 269.15, 269.75, 
    269.35, 269.25, 269.55, 269.15, 269.45, 269.75, 269.75, 269.85, 269.85, 
    270.05, 269.95, 269.85, 269.65, 269.35, 269.15, 268.65, 268.55, 268.25, 
    268.65, 268.25, 268.15, 268.65, 269.55, 269.95, 269.95, 270.45, 270.85, 
    271.05, 271.55, 271.55, 271.15, 271.15, 270.85, 270.65, 270.45, 270.35, 
    270.25, 270.15, 270.75, 270.85, 270.85, 270.95, 270.55, 270.55, 270.45, 
    270.65, 270.75, 270.75, 270.85, 271.45, 271.75, 272.15, 272.35, 272.05, 
    272.25, 273.15, 273.35, 273.45, 273.85, 274.45, 275.25, 275.25, 275.15, 
    275.05, 274.85, 275.15, 275.25, 275.35, 275.15, 274.75, 275.35, 275.15, 
    275.55, 275.15, 275.45, 275.75, 275.85, 275.65, 275.45, 276.25, 276.15, 
    275.15, 274.95, 275.05, 273.45, 274.35, 275.05, 274.65, 274.35, 274.75, 
    274.65, 275.25, 275.75, 275.55, 275.45, 274.85, 274.55, 275.25, 274.55, 
    274.65, 274.25, 272.85, 272.75, 272.95, 274.25, 273.85, 272.95, 273.45, 
    272.65, 272.25, 272.35, 273.05, 272.65, 272.25, 272.35, 272.25, 272.55, 
    272.15, 272.25, 272.35, 271.45, 271.75, 271.65, 271.65, 272.35, 273.45, 
    273.65, 272.95, 272.75, 272.55, 272.35, 272.15, 272.15, 272.05, 271.95, 
    272.15, 272.05, 271.75, 272.15, 273.05, 272.65, 272.95, 272.95, 272.55, 
    272.45, 272.55, 272.95, 272.75, 273.15, 273.25, 273.45, 274.65, 274.45, 
    274.45, 274.65, 274.35, 274.35, 273.75, 274.25, 274.25, 273.95, 273.85, 
    273.95, 273.55, 273.85, 273.75, 273.95, 273.75, 273.45, 273.15, 272.85, 
    272.75, 272.65, 272.85, 271.85, 271.55, 270.95, 271.75, 271.35, 270.65, 
    269.85, 269.95, 269.65, 270.65, 270.65, 270.45, 270.55, 270.15, 270.25, 
    270.15, 269.95, 269.75, 269.75, 269.65, 269.75, 267.25, 266.75, 267.45, 
    267.05, 267.55, 268.05, 267.45, 267.15, 266.95, 266.15, 266.65, 266.85, 
    267.35, 264.65, 264.55, 264.65, 265.75, 265.45, 265.25, 264.55, 264.45, 
    264.25, 263.45, 262.15, 261.55, 261.45, 260.25, 261.05, 260.35, 261.55, 
    260.65, 261.45, 260.35, 262.05, 262.35, 262.25, 263.05, 263.65, 263.25, 
    263.15, 263.45, 263.75, 262.95, 262.15, 262.65, 264.75, 265.25, 264.75, 
    265.05, 265.45, 265.65, 265.35, 265.95, 265.75, 265.55, 264.55, 263.75, 
    263.35, 263.05, 262.65, 262.75, 262.45, 262.05, 261.95, 261.25, 260.85, 
    261.25, 261.15, 262.45, 263.15, 263.15, 263.55, 264.05, 264.85, 265.05, 
    266.05, 265.75, 266.05, 265.55, 266.25, 266.25, 266.95, 267.65, 269.25, 
    269.05, 268.85, 269.15, 269.55, 269.95, 269.95, 271.75, 272.35, 271.85, 
    272.95, 274.35, 275.25, 274.95, 274.25, 274.15, 273.85, 273.65, 273.85, 
    273.55, 273.35, 274.05, 273.65, 274.25, 273.45, 272.45, 271.35, 271.35, 
    270.75, 271.25, 269.95, 269.05, 267.95, 268.75, 266.45, 266.15, 268.25, 
    265.85, 268.05, 267.15, 267.55, 269.35, 269.15, 268.85, 270.55, 271.95, 
    271.35, 271.95, 272.35, 272.15, 271.95, 271.05, 270.95, 270.85, 271.05, 
    271.05, 270.85, 270.95, 270.95, 270.85, 271.45, 272.05, 273.25, 272.45, 
    272.75, 272.65, 275.25, 275.55, 275.45, 275.35, 275.75, 275.95, 275.95, 
    276.25, 275.25, 273.85, 273.25, 271.65, 269.25, 266.95, 264.65, 264.25, 
    262.75, 262.35, 260.65, 259.75, 258.95, 258.45, 258.15, 258.65, 257.85, 
    257.15, 258.05, 258.15, 258.25, 256.55, 259.45, 258.05, 258.85, 257.95, 
    259.25, 260.75, 258.85, 260.15, 260.45, 259.35, 259.35, 259.95, 258.95, 
    259.05, 260.35, 260.95, 260.15, 259.65, 258.75, 259.85, 258.75, 260.45, 
    257.65, 258.65, 258.45, 258.75, 257.75, 258.85, 257.85, 259.05, 258.75, 
    259.15, 259.45, 260.05, 260.15, 260.75, 261.05, 261.35, 261.45, 261.85, 
    262.25, 262.65, 263.75, 264.75, 266.05, 266.35, 266.05, 266.15, 266.55, 
    267.05, 268.55, 269.05, 270.55, 272.55, 274.55, 276.25, 276.35, 276.45, 
    276.75, 276.35, 275.65, 275.55, 276.25, 276.35, 276.55, 276.75, 276.05, 
    275.65, 275.75, 275.35, 275.35, 274.35, 273.95, 273.35, 273.25, 273.15, 
    272.85, 273.05, 272.65, 272.65, 272.85, 272.75, 272.45, 273.15, 272.95, 
    272.75, 272.65, 272.95, 272.35, 271.85, 271.95, 273.35, 272.75, 273.15, 
    273.45, 273.45, 273.85, 273.65, 272.75, 272.65, 272.05, 272.45, 272.65, 
    273.75, 274.05, 273.75, 273.85, 273.75, 273.85, 274.25, 274.05, 273.75, 
    274.15, 273.45, 273.25, 273.55, 273.45, 273.75, 273.65, 273.45, 273.25, 
    272.95, 272.95, 272.55, 272.45, 272.85, 272.65, 272.15, 272.85, 271.75, 
    272.15, 275.15, 274.45, 274.05, 273.85, 273.25, 273.85, 274.15, 273.15, 
    271.85, 272.45, 271.75, 271.25, 270.95, 270.15, 269.05, 268.05, 267.25, 
    266.85, 266.25, 265.55, 264.65, 264.35, 263.75, 263.15, 262.35, 262.05, 
    261.85, 261.45, 261.25, 260.75, 260.45, 259.85, 259.65, 259.75, 259.05, 
    258.75, 257.45, 256.35, 256.35, 255.75, 255.35, 256.25, 255.45, 255.15, 
    255.05, 254.75, 255.25, 255.65, 256.45, 256.15, 256.15, 255.85, 256.65, 
    257.75, 258.15, 258.85, 259.35, 260.15, 260.55, 261.75, 261.85, 262.35, 
    262.75, 262.95, 263.35, 263.55, 265.25, 264.95, 264.65, 264.85, 264.45, 
    264.25, 264.05, 264.05, 263.85, 263.65, 263.95, 263.75, 263.55, 263.25, 
    263.25, 263.45, 263.35, 262.85, 262.65, 262.65, 262.95, 262.85, 262.45, 
    262.05, 261.85, 261.85, 261.65, 261.55, 261.45, 261.45, 261.35, 261.25, 
    260.95, 260.45, 259.95, 259.35, 258.95, 258.85, 258.55, 258.35, 257.95, 
    257.65, 257.45, 256.95, 256.75, 256.55, 256.45, 255.95, 255.95, 255.75, 
    255.65, 255.95, 254.05, 254.25, 253.65, 253.45, 253.35, 253.55, 253.15, 
    253.75, 253.15, 253.15, 252.25, 252.55, 252.05, 252.35, 251.95, 252.55, 
    251.65, 251.75, 252.15, 252.45, 252.85, 253.75, 253.95, 254.35, 254.95, 
    255.55, 255.85, 255.35, 253.45, 253.95, 252.35, 252.15, 250.95, 251.15, 
    250.45, 250.25, 251.25, 250.75, 250.85, 251.15, 251.55, 252.65, 253.75, 
    254.15, 254.45, 254.15, 254.75, 254.05, 253.35, 253.55, 254.95, 254.25, 
    254.25, 254.65, 254.85, 254.45, 254.45, 254.25, 254.55, 254.65, 254.15, 
    254.95, 256.65, 259.05, 258.75, 258.05, 257.65, 258.35, 257.65, 257.25, 
    259.15, 257.75, 256.95, 256.15, 256.05, 256.05, 255.85, 255.35, 255.75, 
    255.85, 255.25, 255.65, 254.45, 254.95, 255.95, 254.95, 255.35, 254.75, 
    256.55, 256.15, 256.35, 255.65, 254.25, 255.45, 255.55, 254.75, 253.35, 
    253.95, 253.85, 254.25, 255.25, 253.15, 253.75, 254.25, 255.05, 253.95, 
    252.55, 253.35, 253.25, 252.65, 252.85, 253.15, 253.45, 252.75, 253.75, 
    255.15, 255.65, 254.65, 254.95, 255.05, 254.95, 255.15, 255.75, 254.95, 
    254.15, 255.25, 255.35, 257.45, 255.25, 255.05, 254.35, 255.75, 255.45, 
    256.85, 256.65, 256.55, 256.45, 256.75, 256.45, 256.05, 256.75, 255.45, 
    255.75, 255.45, 255.65, 255.55, 255.95, 256.45, 255.45, 255.15, 255.75, 
    255.55, 255.15, 254.75, 254.65, 255.05, 253.55, 255.55, 256.45, 257.05, 
    257.65, 258.55, 259.45, 260.25, 260.55, 260.55, 260.75, 261.95, 262.05, 
    262.95, 262.95, 263.55, 264.15, 264.75, 265.35, 265.85, 266.45, 267.25, 
    265.65, 264.65, 265.55, 265.35, 265.05, 265.85, 264.25, 263.75, 262.95, 
    264.05, 264.05, 262.25, 263.05, 263.05, 262.45, 263.45, 263.25, 262.35, 
    264.15, 263.85, 264.05, 263.75, 261.65, 263.65, 264.35, 265.35, 266.05, 
    266.35, 266.65, 266.85, 267.35, 267.85, 268.05, 268.55, 268.95, 269.85, 
    269.55, 269.35, 268.85, 268.15, 268.25, 267.95, 267.85, 267.25, 267.75, 
    268.15, 267.85, 268.65, 268.35, 268.25, 268.05, 268.05, 268.35, 268.25, 
    268.35, 268.55, 267.95, 268.25, 268.25, 268.55, 268.75, 268.85, 268.85, 
    268.75, 268.85, 269.05, 269.05, 268.75, 268.35, 268.45, 268.25, 267.85, 
    267.45, 266.85, 266.95, 266.75, 266.45, 266.25, 266.25, 266.55, 266.55, 
    266.35, 266.05, 265.95, 265.95, 265.95, 265.85, 266.05, 265.75, 265.45, 
    265.05, 265.45, 265.45, 266.15, 266.95, 267.55, 267.75, 267.85, 268.95, 
    269.55, 269.45, 269.35, 269.35, 268.85, 268.65, 268.15, 268.05, 267.75, 
    267.65, 267.55, 267.05, 267.05, 266.95, 266.65, 266.55, 266.15, 265.95, 
    265.85, 265.75, 265.35, 265.55, 265.55, 265.85, 265.45, 265.25, 264.85, 
    263.65, 264.45, 264.65, 264.35, 264.75, 265.05, 265.05, 265.05, 264.75, 
    265.45, 265.85, 266.25, 266.35, 267.15, 267.45, 267.45, 266.45, 265.55, 
    264.75, 264.55, 263.75, 264.15, 263.55, 263.35, 262.45, 262.75, 263.25, 
    262.85, 262.35, 262.95, 262.85, 263.15, 263.95, 269.25, 268.75, 268.65, 
    267.95, 269.15, 269.75, 269.35, 268.95, 270.15, 269.05, 268.25, 267.15, 
    267.15, 266.25, 266.05, 266.05, 266.05, 266.05, 264.95, 264.65, 264.35, 
    263.95, 263.45, 262.85, 262.65, 262.85, 262.45, 262.45, 262.65, 262.65, 
    262.65, 262.55, 262.55, 262.45, 262.35, 262.65, 262.45, 262.45, 262.25, 
    261.85, 261.85, 261.65, 261.35, 261.25, 260.05, 261.65, 261.35, 260.55, 
    259.95, 259.55, 259.35, 260.15, 261.05, 261.25, 260.85, 258.85, 257.85, 
    257.75, 258.55, 258.55, 257.25, 258.05, 256.85, 258.15, 258.25, 259.55, 
    260.75, 261.05, 261.25, 260.65, 259.75, 259.95, 259.15, 259.35, 260.15, 
    260.65, 260.75, 263.35, 264.15, 264.55, 265.05, 265.15, 265.15, 265.25, 
    265.45, 265.25, 265.05, 264.35, 263.45, 262.85, 263.45, 263.35, 263.55, 
    261.65, 259.15, 260.85, 259.85, 260.75, 259.75, 260.35, 259.95, 260.85, 
    259.85, 260.55, 259.95, 260.05, 259.05, 259.75, 260.25, 258.95, 259.15, 
    260.75, 259.75, 259.35, 258.75, 258.85, 258.15, 258.85, 258.75, 258.35, 
    257.85, 258.65, 257.95, 257.55, 257.45, 257.65, 257.65, 256.35, 257.75, 
    257.55, 257.65, 257.65, 256.75, 257.05, 256.75, 256.85, 256.45, 256.85, 
    256.45, 255.45, 255.85, 257.45, 256.85, 256.65, 256.85, 256.95, 255.75, 
    255.75, 257.65, 257.85, 257.15, 256.95, 257.35, 257.95, 258.55, 258.55, 
    258.85, 258.65, 258.85, 259.05, 259.15, 259.15, 259.75, 260.25, 261.15, 
    261.25, 261.25, 262.45, 261.85, 262.65, 262.35, 261.75, 259.65, 259.85, 
    260.45, 260.25, 261.25, 260.85, 260.35, 260.75, 261.25, 259.75, 259.35, 
    258.15, 257.35, 256.55, 255.45, 257.45, 256.75, 256.65, 257.85, 259.45, 
    259.25, 256.75, 256.55, 256.55, 256.75, 259.55, 258.25, 259.25, 259.35, 
    259.55, 259.25, 259.15, 259.05, 258.85, 258.75, 258.35, 258.15, 258.05, 
    258.05, 257.75, 258.15, 257.85, 257.55, 257.45, 257.35, 257.55, 257.05, 
    257.15, 256.55, 255.25, 255.25, 255.35, 254.75, 254.35, 254.45, 253.75, 
    253.15, 253.95, 254.15, 252.85, 253.25, 253.15, 253.75, 253.85, 253.95, 
    254.15, 254.45, 253.55, 254.15, 253.55, 254.05, 254.25, 253.85, 253.65, 
    253.75, 254.05, 253.45, 253.85, 253.05, 253.15, 253.15, 253.25, 252.45, 
    252.65, 252.85, 252.05, 252.15, 252.35, 253.25, 253.05, 251.95, 252.85, 
    251.95, 251.25, 252.05, 251.95, 251.05, 251.45, 252.25, 252.25, 251.55, 
    253.15, 251.85, 252.85, 252.95, 251.65, 252.25, 252.95, 250.75, 253.45, 
    253.45, 253.55, 251.95, 253.65, 254.05, 254.15, 254.65, 253.85, 254.85, 
    253.55, 253.95, 254.25, 254.75, 253.55, 252.95, 254.75, 253.55, 254.05, 
    253.55, 254.35, 253.85, 252.75, 254.15, 253.75, 255.15, 254.35, 254.65, 
    254.85, 255.55, 253.95, 254.15, 254.65, 254.75, 255.95, 255.95, 254.85, 
    255.15, 255.95, 255.65, 256.65, 255.75, 256.55, 257.05, 256.95, 256.75, 
    256.25, 258.75, 257.75, 256.25, 256.95, 255.75, 258.45, 255.85, 257.35, 
    257.15, 258.45, 258.15, 256.85, 256.85, 257.45, 257.45, 257.95, 256.75, 
    258.35, 257.95, 260.65, 259.15, 260.05, 260.15, 260.85, 260.55, 261.75, 
    261.55, 262.35, 262.35, 262.45, 263.15, 262.95, 263.65, 263.35, 264.15, 
    263.85, 263.05, 263.55, 263.45, 263.75, 262.95, 263.75, 263.75, 263.15, 
    261.85, 262.25, 261.95, 260.85, 262.65, 263.05, 262.05, 261.05, 262.35, 
    263.25, 261.45, 260.65, 261.65, 262.25, 263.35, 260.65, 262.25, 261.95, 
    265.05, 262.15, 262.55, 265.35, 263.45, 265.35, 265.85, 264.45, 264.95, 
    264.85, 265.75, 264.45, 266.05, 264.25, 263.85, 265.25, 266.85, 264.85, 
    265.35, 265.95, 265.45, 267.35, 266.55, 266.75, 266.15, 266.25, 265.75, 
    265.45, 265.65, 264.35, 265.65, 265.85, 265.35, 266.05, 266.45, 266.95, 
    268.05, 267.45, 266.45, 265.95, 264.95, 266.65, 264.55, 264.25, 263.45, 
    262.65, 261.65, 263.05, 264.15, 262.05, 262.45, 263.05, 262.95, 263.45, 
    265.55, 267.05, 267.75, 268.45, 268.25, 268.95, 269.05, 269.35, 268.85, 
    268.55, 267.95, 268.65, 268.95, 268.85, 269.25, 269.25, 269.25, 269.25, 
    268.95, 269.15, 269.05, 269.05, 269.55, 269.55, 269.55, 269.85, 270.35, 
    270.25, 270.95, 270.85, 270.45, 269.75, 269.25, 271.25, 271.75, 271.65, 
    271.65, 271.75, 271.65, 271.65, 271.95, 271.95, 271.35, 271.85, 272.45, 
    272.25, 272.05, 272.05, 271.85, 272.05, 271.95, 272.55, 272.95, 272.85, 
    271.85, 271.45, 271.45, 270.05, 269.15, 268.85, 267.45, 266.45, 269.05, 
    268.75, 269.85, 271.35, 269.95, 270.55, 271.05, 271.55, 272.05, 270.65, 
    272.95, 271.85, 272.55, 272.45, 272.95, 272.75, 272.55, 272.25, 272.35, 
    272.35, 272.05, 271.95, 271.45, 271.55, 270.75, 270.15, 269.55, 269.15, 
    269.75, 269.65, 269.65, 269.15, 269.75, 269.05, 269.35, 269.55, 267.85, 
    267.45, 267.45, 268.25, 267.95, 268.15, 267.95, 268.85, 268.45, 268.55, 
    270.05, 270.15, 270.35, 270.25, 270.25, 270.15, 270.25, 270.45, 270.45, 
    270.15, 270.45, 270.55, 270.25, 270.75, 271.05, 271.05, 270.95, 270.75, 
    271.15, 271.45, 271.95, 271.15, 271.25, 271.45, 271.35, 271.05, 270.85, 
    271.15, 271.05, 271.45, 271.15, 271.35, 271.05, 271.15, 271.05, 271.35, 
    270.65, 269.25, 269.95, 269.65, 269.95, 270.25, 270.75, 270.65, 271.15, 
    269.95, 271.25, 270.75, 270.75, 270.15, 270.85, 269.65, 270.45, 270.75, 
    270.45, 269.75, 270.75, 269.45, 269.65, 270.45, 270.55, 270.05, 269.55, 
    269.65, 270.15, 269.65, 269.65, 269.85, 269.85, 269.75, 269.65, 268.95, 
    269.15, 267.95, 268.35, 268.35, 268.05, 267.85, 267.55, 267.15, 267.25, 
    267.35, 267.55, 266.75, 266.35, 264.95, 265.55, 264.65, 264.65, 264.95, 
    264.25, 264.55, 263.95, 264.25, 264.55, 264.25, 263.85, 264.15, 264.05, 
    263.35, 263.35, 264.55, 264.45, 264.95, 264.35, 264.85, 265.15, 265.15, 
    264.55, 262.95, 264.75, 264.55, 268.25, 268.75, 269.15, 268.95, 269.15, 
    269.15, 268.95, 268.75, 268.75, 268.85, 268.65, 268.35, 268.65, 268.35, 
    268.25, 268.05, 268.15, 267.75, 267.05, 267.05, 266.85, 267.15, 267.65, 
    267.25, 266.95, 266.75, 267.15, 267.25, 267.25, 267.25, 266.15, 266.85, 
    266.55, 265.55, 265.15, 263.45, 266.45, 265.85, 264.05, 265.75, 265.95, 
    266.15, 265.35, 265.35, 265.35, 263.85, 264.45, 263.25, 262.65, 263.05, 
    263.65, 264.05, 264.55, 265.95, 265.55, 264.95, 264.85, 264.55, 262.55, 
    261.25, 261.85, 260.05, 260.95, 260.75, 260.65, 262.45, 261.25, 260.15, 
    259.75, 260.15, 259.95, 260.75, 260.05, 260.35, 260.15, 261.35, 261.35, 
    262.35, 264.15, 263.45, 262.75, 262.55, 262.15, 262.25, 262.05, 262.25, 
    261.55, 261.05, 260.95, 260.35, 260.45, 259.85, 259.05, 259.35, 258.75, 
    259.25, 259.05, 260.55, 259.35, 259.45, 260.15, 260.55, 261.35, 262.15, 
    263.95, 264.75, 265.05, 265.15, 265.25, 265.35, 265.55, 265.35, 264.95, 
    264.35, 264.15, 263.65, 263.35, 263.15, 263.35, 262.75, 262.25, 262.45, 
    262.45, 262.05, 261.95, 262.25, 261.75, 261.85, 261.55, 261.75, 261.45, 
    261.15, 261.05, 261.05, 260.55, 260.15, 259.85, 259.45, 258.85, 258.25, 
    256.15, 256.55, 255.95, 255.85, 255.65, 255.15, 255.35, 254.95, 254.45, 
    254.85, 253.95, 254.15, 254.05, 253.55, 253.05, 255.25, 254.15, 253.55, 
    254.35, 253.65, 253.15, 253.55, 253.35, 254.85, 253.75, 254.45, 254.35, 
    254.95, 256.55, 255.05, 257.25, 256.55, 257.85, 257.35, 257.65, 259.35, 
    257.55, 261.25, 259.35, 259.55, 258.95, 259.55, 258.25, 260.25, 257.95, 
    258.35, 259.85, 258.65, 257.35, 257.65, 258.15, 258.95, 258.65, 258.65, 
    259.35, 259.65, 259.85, 260.45, 261.05, 259.65, 258.95, 257.95, 258.55, 
    258.45, 257.95, 257.05, 256.45, 257.05, 257.65, 255.85, 255.85, 257.75, 
    256.15, 256.55, 256.85, 260.15, 259.35, 258.95, 258.15, 257.75, 257.15, 
    257.25, 257.75, 257.65, 257.35, 257.05, 256.65, 256.05, 255.35, 254.95, 
    254.95, 254.45, 253.85, 253.25, 252.85, 251.85, 251.15, 250.35, 250.75, 
    249.45, 248.55, 247.15, 247.45, 247.95, 248.15, 248.15, 248.55, 248.35, 
    248.55, 248.75, 248.85, 248.75, 249.05, 248.75, 249.05, 249.15, 249.25, 
    248.55, 248.55, 248.25, 248.25, 249.05, 248.15, 248.65, 249.05, 248.35, 
    248.35, 248.35, 247.95, 248.55, 248.85, 250.65, 248.15, 248.15, 248.25, 
    246.95, 247.95, 247.45, 248.35, 249.15, 249.65, 250.05, 249.15, 249.15, 
    249.65, 249.45, 249.05, 249.15, 249.25, 248.85, 248.55, 248.85, 248.75, 
    248.45, 248.25, 248.75, 248.05, 247.35, 246.95, 247.65, 248.85, 247.15, 
    247.95, 247.85, 247.95, 248.05, 247.45, 249.35, 249.35, 248.55, 250.05, 
    249.55, 250.25, 250.85, 250.45, 251.15, 251.05, 251.65, 251.85, 251.75, 
    252.35, 252.85, 253.05, 252.75, 252.65, 252.15, 252.05, 253.65, 252.95, 
    253.35, 252.45, 253.55, 255.05, 255.85, 256.25, 257.05, 257.85, 257.75, 
    258.15, 259.65, 258.95, 259.15, 259.05, 259.55, 258.85, 258.85, 258.55, 
    258.35, 258.35, 258.45, 258.95, 259.65, 260.55, 259.85, 260.15, 260.55, 
    260.35, 261.05, 261.75, 272.25, 272.55, 271.85, 272.15, 272.85, 273.05, 
    273.45, 273.35, 273.35, 273.25, 273.05, 273.95, 274.45, 274.25, 273.35, 
    273.25, 273.35, 272.95, 272.55, 271.95, 271.85, 271.85, 271.05, 271.95, 
    271.05, 270.55, 270.65, 271.85, 273.55, 272.95, 272.15, 269.85, 269.95, 
    268.45, 268.55, 267.75, 267.55, 267.15, 267.45, 265.05, 264.45, 264.55, 
    264.05, 262.45, 262.75, 263.15, 263.05, 263.65, 263.45, 263.05, 263.05, 
    263.15, 263.85, 263.35, 262.85, 262.95, 263.15, 263.15, 264.75, 264.65, 
    264.95, 264.85, 264.15, 264.05, 263.75, 263.35, 262.95, 261.55, 260.35, 
    259.55, 258.85, 257.25, 257.05, 256.95, 255.95, 254.95, 254.35, 253.95, 
    253.95, 253.85, 253.35, 253.45, 253.25, 253.15, 252.75, 251.05, 250.45, 
    251.35, 250.65, 249.75, 249.25, 249.15, 249.25, 249.35, 250.25, 251.15, 
    251.15, 250.75, 250.75, 250.25, 250.75, 250.35, 250.85, 251.35, 250.05, 
    250.05, 251.05, 251.15, 252.05, 250.95, 250.75, 251.45, 253.15, 253.45, 
    255.05, 253.85, 255.35, 255.75, 256.65, 256.15, 258.65, 257.45, 258.35, 
    257.75, 258.25, 258.75, 258.15, 258.15, 258.85, 256.95, 258.95, 259.75, 
    258.45, 258.25, 257.45, 259.45, 258.55, 258.65, 258.15, 257.85, 257.15, 
    256.25, 256.45, 257.85, 258.35, 258.05, 257.55, 257.35, 258.05, 258.05, 
    257.55, 258.05, 257.95, 257.85, 258.55, 257.65, 257.45, 256.75, 256.95, 
    256.95, 257.45, 256.85, 256.75, 257.45, 256.25, 256.75, 257.35, 256.95, 
    256.45, 256.45, 257.15, 257.35, 256.95, 256.45, 256.25, 255.75, 255.55, 
    255.45, 254.75, 255.05, 255.05, 254.95, 256.25, 255.85, 255.75, 256.15, 
    256.25, 256.35, 257.35, 256.35, 256.35, 255.25, 255.65, 255.45, 255.25, 
    254.85, 254.55, 255.15, 254.85, 254.65, 254.15, 255.45, 255.25, 254.95, 
    254.45, 254.45, 255.05, 253.15, 252.95, 252.15, 251.45, 252.35, 252.95, 
    253.05, 252.05, 252.85, 251.65, 253.15, 252.65, 252.25, 253.25, 254.05, 
    256.45, 254.65, 255.75, 255.55, 255.85, 254.55, 254.65, 254.25, 254.35, 
    253.85, 254.15, 253.85, 254.05, 253.65, 253.35, 252.85, 252.65, 252.35, 
    251.95, 251.95, 251.55, 252.05, 251.65, 252.15, 251.65, 250.85, 250.85, 
    249.15, 250.55, 253.05, 251.85, 251.65, 252.95, 254.05, 254.45, 254.15, 
    254.35, 253.45, 252.45, 252.45, 252.85, 251.25, 250.75, 251.55, 250.75, 
    251.25, 251.15, 251.95, 252.35, 252.75, 252.35, 252.55, 253.65, 253.65, 
    253.55, 252.45, 253.75, 254.35, 253.85, 253.15, 252.45, 252.45, 251.85, 
    253.05, 252.05, 251.75, 254.25, 253.25, 252.85, 252.45, 250.85, 250.95, 
    250.55, 252.65, 252.05, 253.05, 254.35, 256.25, 258.55, 261.85, 259.45, 
    262.25, 262.25, 262.35, 262.55, 262.65, 261.65, 261.25, 261.85, 262.05, 
    258.95, 258.55, 259.55, 259.45, 259.65, 259.35, 257.45, 260.05, 259.55, 
    257.35, 255.65, 256.15, 255.35, 255.35, 258.25, 255.05, 257.55, 255.95, 
    254.25, 256.05, 254.75, 254.65, 254.95, 255.25, 255.75, 255.35, 255.95, 
    255.35, 255.55, 255.95, 254.85, 254.15, 254.25, 254.45, 254.45, 255.75, 
    254.95, 254.85, 254.35, 254.75, 254.45, 253.85, 253.75, 254.15, 254.15, 
    252.35, 252.95, 254.85, 255.45, 254.25, 252.55, 253.55, 254.85, 253.35, 
    252.75, 253.95, 254.25, 254.15, 255.35, 253.85, 253.75, 254.45, 253.35, 
    253.85, 254.35, 253.75, 255.95, 255.05, 255.05, 256.05, 255.35, 256.55, 
    257.95, 256.25, 256.85, 256.35, 256.05, 255.95, 254.95, 254.65, 255.85, 
    255.05, 254.55, 253.85, 255.15, 255.25, 255.45, 256.35, 254.65, 255.55, 
    254.05, 253.25, 254.35, 254.05, 253.05, 253.35, 253.25, 252.55, 253.85, 
    254.85, 252.25, 252.65, 251.65, 252.95, 251.65, 251.15, 251.35, 252.65, 
    251.35, 252.85, 254.25, 254.05, 253.75, 253.15, 251.65, 252.25, 252.75, 
    252.65, 252.35, 251.85, 252.25, 252.95, 253.55, 253.25, 252.35, 252.45, 
    253.65, 252.85, 252.35, 253.25, 252.85, 251.55, 253.15, 252.15, 252.95, 
    252.85, 253.55, 253.55, 254.05, 253.75, 253.55, 253.55, 254.55, 254.85, 
    255.45, 255.55, 255.25, 254.25, 254.85, 254.75, 254.65, 255.05, 254.35, 
    255.35, 256.45, 255.55, 255.25, 254.05, 253.75, 254.15, 254.95, 254.65, 
    254.25, 253.65, 252.85, 254.65, 253.85, 252.45, 253.65, 251.75, 251.35, 
    253.75, 252.65, 252.95, 252.65, 252.15, 252.55, 252.95, 251.55, 251.95, 
    251.45, 253.55, 252.05, 254.65, 255.55, 254.05, 252.45, 252.45, 252.75, 
    253.05, 253.25, 252.35, 251.85, 252.45, 252.15, 251.75, 253.65, 251.65, 
    253.15, 251.85, 253.05, 254.55, 254.75, 255.05, 254.55, 255.35, 255.75, 
    256.05, 255.85, 256.65, 256.55, 256.15, 255.75, 255.85, 256.25, 255.75, 
    255.55, 255.45, 255.15, 254.25, 254.15, 253.85, 253.05, 252.85, 253.15, 
    251.55, 251.15, 251.75, 251.85, 253.15, 254.05, 253.35, 255.25, 254.65, 
    253.35, 254.15, 252.65, 253.05, 253.75, 251.55, 249.65, 251.15, 251.85, 
    249.95, 249.65, 251.55, 249.55, 251.85, 249.65, 251.05, 251.75, 250.25, 
    250.45, 251.95, 255.25, 253.45, 253.25, 254.75, 254.95, 254.05, 253.35, 
    254.65, 256.05, 257.05, 256.55, 256.45, 257.05, 257.05, 257.55, 257.45, 
    260.65, 262.05, 262.65, 261.15, 260.55, 260.75, 263.65, 264.75, 269.45, 
    270.15, 269.95, 270.45, 270.25, 270.55, 269.95, 268.45, 267.45, 265.45, 
    263.95, 263.55, 262.15, 262.75, 261.85, 261.35, 260.95, 260.25, 260.15, 
    260.25, 260.65, 260.45, 260.95, 261.35, 262.05, 262.05, 261.95, 262.55, 
    261.65, 261.75, 261.55, 261.15, 261.95, 261.25, 263.15, 265.15, 263.65, 
    267.45, 268.45, 268.75, 269.15, 269.15, 270.25, 271.25, 271.45, 272.45, 
    272.85, 275.25, 275.25, 276.05, 275.15, 275.35, 275.75, 274.85, 273.85, 
    273.55, 273.15, 272.75, 272.55, 272.05, 271.55, 271.75, 271.45, 271.35, 
    270.05, 269.45, 269.85, 267.85, 268.15, 267.35, 266.15, 267.95, 266.15, 
    267.15, 266.95, 266.55, 265.55, 264.15, 263.75, 263.55, 264.65, 266.65, 
    265.35, 264.45, 264.05, 263.15, 265.05, 262.15, 265.65, 267.15, 266.35, 
    268.35, 267.65, 271.15, 269.25, 270.45, 270.45, 270.05, 270.25, 269.75, 
    269.45, 268.95, 268.55, 268.25, 265.75, 265.45, 264.45, 263.95, 262.85, 
    263.35, 263.45, 262.85, 264.05, 264.05, 264.15, 264.15, 265.65, 265.15, 
    265.75, 266.25, 266.55, 266.65, 268.15, 268.35, 267.75, 267.25, 266.85, 
    266.95, 266.85, 265.35, 265.45, 262.95, 262.85, 262.95, 263.25, 261.05, 
    261.75, 264.15, 263.65, 265.15, 266.65, 265.95, 265.95, 265.85, 265.75, 
    266.35, 265.75, 264.35, 263.85, 262.65, 261.75, 260.85, 259.35, 258.25, 
    257.55, 255.85, 255.55, 256.45, 255.85, 257.25, 258.45, 259.75, 262.65, 
    263.55, 263.45, 262.85, 262.45, 263.15, 262.45, 262.25, 262.85, 262.75, 
    262.05, 260.95, 262.25, 261.65, 261.05, 260.35, 260.15, 259.95, 259.35, 
    258.65, 258.45, 257.85, 256.75, 255.05, 254.55, 255.05, 256.15, 255.65, 
    256.15, 256.75, 257.45, 258.65, 258.95, 258.75, 260.05, 260.45, 260.85, 
    261.15, 261.55, 260.25, 260.25, 261.15, 260.85, 261.05, 261.15, 261.85, 
    262.85, 264.65, 264.55, 264.45, 265.85, 265.75, 265.05, 265.15, 264.95, 
    266.35, 267.05, 267.85, 267.15, 267.85, 267.05, 267.05, 267.05, 266.35, 
    266.95, 266.95, 267.05, 265.25, 265.75, 265.35, 267.65, 267.95, 268.05, 
    267.45, 267.35, 267.05, 266.15, 266.75, 267.35, 267.25, 267.65, 267.85, 
    268.25, 267.75, 267.85, 267.45, 268.25, 268.85, 268.25, 269.95, 270.25, 
    270.25, 270.35, 270.45, 270.55, 269.75, 269.45, 269.25, 269.75, 269.35, 
    269.65, 270.05, 270.05, 270.15, 270.25, 269.75, 269.65, 270.05, 269.55, 
    269.15, 269.95, 269.65, 267.85, 267.65, 267.45, 267.05, 266.35, 266.75, 
    265.45, 266.15, 267.25, 266.65, 267.25, 267.05, 267.65, 267.95, 267.55, 
    268.05, 266.95, 265.85, 266.45, 266.85, 266.85, 265.15, 264.65, 264.55, 
    263.45, 262.75, 260.95, 260.55, 260.55, 260.75, 260.75, 260.35, 261.05, 
    259.65, 259.05, 259.95, 260.85, 260.35, 260.85, 260.65, 261.55, 261.25, 
    260.75, 260.75, 261.05, 260.85, 260.55, 260.25, 259.65, 260.15, 259.55, 
    259.65, 259.15, 257.85, 259.35, 257.85, 258.35, 257.15, 257.35, 257.25, 
    258.05, 258.45, 259.15, 260.15, 259.55, 259.65, 260.25, 260.65, 260.25, 
    259.05, 259.45, 258.45, 258.85, 258.65, 258.45, 257.75, 258.15, 257.75, 
    256.15, 257.85, 256.15, 256.55, 256.85, 256.75, 256.95, 257.15, 257.65, 
    258.05, 257.95, 257.85, 257.75, 257.95, 258.45, 257.35, 256.05, 254.75, 
    255.45, 254.45, 255.75, 254.65, 254.95, 254.25, 254.85, 255.35, 255.75, 
    255.55, 256.15, 256.85, 257.05, 258.05, 258.55, 260.35, 260.55, 260.15, 
    260.75, 260.65, 260.35, 259.45, 258.75, 258.75, 257.75, 257.75, 257.85, 
    257.25, 256.95, 258.05, 257.45, 256.85, 256.75, 256.55, 257.95, 258.15, 
    259.75, 260.75, 261.65, 261.45, 261.65, 263.35, 263.45, 263.35, 263.15, 
    263.55, 263.45, 264.35, 263.25, 264.95, 266.05, 266.05, 267.85, 266.75, 
    265.55, 271.55, 270.25, 270.05, 269.15, 269.35, 269.55, 269.25, 269.45, 
    268.75, 268.55, 267.65, 266.35, 265.75, 265.25, 264.15, 263.85, 263.75, 
    264.05, 264.55, 262.55, 262.35, 263.25, 262.55, 263.25, 264.15, 263.45, 
    263.05, 262.85, 263.55, 263.65, 264.45, 264.95, 265.45, 265.35, 264.95, 
    266.65, 266.15, 266.35, 266.65, 266.45, 265.85, 265.55, 264.15, 264.35, 
    263.85, 263.65, 263.35, 264.05, 263.75, 262.75, 262.55, 262.35, 261.15, 
    261.55, 262.65, 261.35, 262.15, 262.95, 262.15, 264.35, 262.05, 264.15, 
    261.25, 260.45, 260.85, 258.95, 258.05, 258.95, 257.15, 258.35, 258.85, 
    258.45, 257.05, 257.85, 259.35, 258.95, 259.85, 258.95, 261.75, 261.95, 
    260.15, 261.25, 262.15, 262.95, 264.55, 262.35, 261.45, 260.15, 259.05, 
    258.85, 259.15, 260.15, 261.55, 260.75, 261.25, 261.95, 261.75, 263.05, 
    263.35, 262.75, 264.75, 265.45, 266.65, 266.95, 266.45, 266.25, 266.75, 
    267.05, 267.15, 267.15, 267.35, 268.15, 268.35, 268.85, 268.35, 267.85, 
    268.85, 268.75, 268.45, 268.25, 268.45, 268.75, 269.85, 270.05, 269.25, 
    270.15, 270.55, 271.65, 271.85, 271.95, 271.85, 273.05, 273.05, 272.85, 
    271.65, 271.65, 271.05, 270.55, 270.25, 269.55, 268.85, 268.35, 268.15, 
    267.65, 267.25, 266.65, 266.75, 266.55, 266.55, 266.05, 266.85, 265.75, 
    266.35, 266.35, 266.85, 266.15, 264.55, 263.55, 263.95, 264.15, 264.25, 
    264.15, 264.45, 264.25, 263.95, 263.75, 263.85, 263.85, 263.95, 264.15, 
    265.35, 265.85, 266.05, 266.45, 266.65, 268.45, 268.25, 268.15, 267.45, 
    268.35, 268.35, 268.35, 267.85, 268.55, 267.15, 267.15, 267.15, 267.65, 
    267.45, 267.55, 267.75, 267.45, 267.15, 268.15, 268.55, 268.55, 269.35, 
    269.85, 270.65, 269.55, 270.15, 269.85, 269.95, 269.55, 269.85, 270.05, 
    270.05, 270.65, 269.35, 268.45, 268.25, 268.25, 268.15, 268.65, 268.25, 
    268.15, 267.45, 267.55, 267.65, 268.05, 268.45, 268.25, 269.25, 269.35, 
    269.45, 269.85, 270.45, 270.95, 271.25, 272.05, 272.95, 272.35, 272.05, 
    271.85, 270.95, 270.35, 270.15, 270.15, 270.15, 269.65, 268.75, 268.35, 
    267.75, 267.85, 268.65, 268.55, 268.65, 269.05, 269.15, 269.15, 269.15, 
    269.15, 269.05, 268.75, 268.95, 269.35, 269.15, 269.05, 269.05, 269.85, 
    275.35, 275.65, 275.85, 275.45, 275.55, 274.85, 275.15, 275.15, 275.35, 
    275.35, 275.35, 275.45, 275.45, 275.65, 275.65, 275.45, 275.35, 275.65, 
    275.35, 275.55, 275.45, 275.15, 274.95, 274.95, 274.25, 275.05, 274.25, 
    273.75, 274.05, 274.75, 274.75, 274.25, 274.15, 273.95, 274.25, 274.55, 
    274.65, 274.65, 274.45, 274.25, 274.05, 274.85, 273.95, 273.95, 273.35, 
    273.35, 273.75, 274.45, 275.45, 275.65, 275.55, 275.35, 275.65, 275.65, 
    275.45, 275.15, 275.45, 275.25, 275.15, 275.45, 275.45, 275.55, 275.75, 
    275.45, 275.25, 275.15, 275.15, 274.75, 275.75, 276.35, 275.85, 276.05, 
    275.75, 275.45, 276.65, 276.75, 275.65, 275.45, 275.45, 275.75, 275.75, 
    275.65, 276.25, 276.75, 276.35, 275.85, 276.35, 275.45, 275.25, 275.15, 
    274.75, 274.05, 273.55, 273.35, 273.25, 272.55, 272.25, 272.15, 271.55, 
    270.05, 268.85, 268.25, 267.85, 268.45, 268.15, 268.45, 269.35, 269.55, 
    271.65, 270.45, 270.55, 270.45, 270.75, 271.55, 271.75, 270.45, 270.05, 
    270.35, 269.55, 268.35, 267.95, 268.35, 268.25, 267.85, 267.55, 267.05, 
    267.25, 267.35, 266.95, 267.05, 267.25, 267.65, 267.45, 268.05, 267.85, 
    267.95, 267.95, 266.55, 265.35, 265.45, 264.55, 263.65, 263.15, 262.15, 
    261.25, 261.25, 260.65, 260.05, 259.75, 259.05, 260.15, 260.45, 261.05, 
    260.65, 261.55, 262.75, 262.65, 262.75, 263.75, 265.35, 265.95, 264.35, 
    264.35, 263.55, 263.15, 263.95, 262.35, 261.95, 262.25, 261.85, 261.95, 
    262.95, 262.55, 262.85, 263.05, 264.05, 263.25, 264.65, 265.25, 267.05, 
    266.75, 267.95, 269.15, 267.25, 268.35, 267.55, 267.55, 267.15, 266.65, 
    266.85, 266.65, 266.45, 266.25, 265.55, 264.15, 264.35, 264.35, 264.35, 
    265.05, 265.55, 265.85, 266.25, 267.85, 268.35, 268.35, 268.75, 269.25, 
    270.45, 270.65, 269.05, 269.05, 269.25, 268.75, 268.75, 268.45, 268.55, 
    268.45, 268.85, 269.35, 269.35, 269.85, 270.35, 271.35, 271.25, 271.75, 
    271.85, 272.25, 272.75, 272.85, 271.95, 271.25, 270.85, 271.05, 271.05, 
    270.95, 271.25, 270.95, 270.95, 270.55, 270.65, 270.75, 270.35, 270.35, 
    270.35, 270.45, 270.65, 270.85, 270.75, 271.85, 272.55, 273.05, 273.35, 
    273.85, 274.65, 272.55, 272.55, 273.55, 271.85, 271.55, 271.65, 272.15, 
    271.55, 271.35, 271.25, 271.15, 270.95, 271.15, 270.85, 271.25, 271.45, 
    271.65, 271.05, 271.75, 272.55, 272.35, 272.35, 272.35, 273.55, 275.25, 
    273.45, 273.15, 273.95, 272.85, 272.95, 272.35, 272.15, 272.35, 272.35, 
    272.45, 272.35, 272.25, 272.05, 272.05, 271.95, 271.95, 272.75, 273.15, 
    273.65, 273.85, 274.85, 274.65, 275.15, 276.65, 275.15, 276.45, 275.75, 
    274.45, 274.85, 273.95, 273.85, 273.45, 273.45, 273.45, 273.55, 273.65, 
    273.45, 273.15, 272.95, 273.05, 272.75, 273.25, 273.25, 273.35, 273.45, 
    273.85, 273.85, 274.05, 273.95, 273.05, 273.25, 273.25, 270.95, 270.55, 
    268.95, 266.95, 268.55, 266.75, 267.25, 266.75, 265.85, 266.15, 265.05, 
    265.05, 264.35, 264.45, 264.75, 265.35, 265.05, 265.75, 265.95, 266.05, 
    265.25, 264.45, 265.55, 265.85, 263.95, 264.75, 265.65, 265.65, 264.35, 
    264.45, 263.95, 262.55, 263.15, 263.05, 263.65, 263.55, 262.75, 263.65, 
    263.55, 263.55, 263.35, 263.85, 263.85, 262.45, 262.35, 262.65, 262.45, 
    262.15, 261.15, 261.05, 260.95, 260.55, 260.45, 260.05, 260.15, 260.55, 
    261.55, 262.45, 263.75, 263.25, 264.15, 265.25, 265.85, 266.95, 268.15, 
    267.95, 266.85, 268.05, 268.15, 266.15, 266.35, 266.15, 268.05, 269.05, 
    268.35, 268.65, 269.05, 270.05, 269.05, 269.05, 269.85, 270.65, 269.15, 
    268.15, 269.05, 269.55, 268.75, 268.55, 270.15, 269.15, 269.15, 269.55, 
    268.55, 269.45, 270.15, 269.35, 269.05, 267.85, 267.35, 267.25, 266.25, 
    266.05, 265.05, 266.05, 264.45, 264.95, 265.05, 266.15, 265.85, 266.45, 
    266.75, 267.35, 267.45, 267.45, 267.75, 268.05, 268.55, 268.35, 268.55, 
    268.55, 268.55, 267.85, 267.05, 265.95, 265.95, 264.85, 264.35, 263.35, 
    263.35, 263.25, 264.05, 264.05, 264.85, 265.15, 266.15, 266.15, 266.35, 
    266.55, 266.55, 266.95, 266.85, 266.75, 266.65, 267.15, 266.05, 265.85, 
    265.25, 265.45, 265.45, 264.85, 264.95, 265.15, 265.65, 265.45, 265.85, 
    266.65, 267.45, 266.85, 267.05, 267.95, 267.95, 269.85, 270.25, 270.55, 
    271.55, 271.35, 270.75, 271.35, 270.75, 269.45, 269.95, 268.25, 267.95, 
    268.05, 267.25, 266.45, 266.25, 266.55, 266.45, 267.25, 267.65, 268.05, 
    268.65, 268.55, 268.55, 268.35, 268.25, 269.25, 269.65, 270.15, 269.45, 
    268.95, 268.75, 269.05, 268.75, 268.15, 267.75, 267.45, 267.45, 266.95, 
    266.95, 266.95, 267.15, 266.95, 267.05, 266.45, 267.15, 267.35, 267.35, 
    267.25, 267.45, 267.55, 267.55, 267.85, 267.25, 266.65, 266.95, 266.45, 
    266.15, 265.55, 265.55, 265.75, 265.55, 265.45, 265.35, 265.65, 266.25, 
    266.85, 267.15, 267.25, 267.75, 267.75, 267.95, 267.45, 267.95, 268.25, 
    268.55, 268.25, 268.25, 267.85, 268.45, 268.25, 267.85, 267.05, 267.05, 
    266.95, 265.95, 264.85, 265.45, 265.15, 265.55, 265.25, 266.35, 266.75, 
    267.65, 267.85, 268.15, 268.85, 269.25, 269.55, 269.55, 269.25, 269.55, 
    268.95, 269.15, 268.65, 268.25, 266.95, 266.75, 266.15, 265.95, 265.65, 
    265.25, 265.05, 266.25, 267.05, 267.05, 268.15, 268.45, 268.65, 268.95, 
    269.95, 270.85, 271.55, 271.15, 270.95, 271.25, 271.15, 271.45, 272.15, 
    271.75, 271.55, 271.35, 271.15, 271.25, 271.25, 271.75, 271.35, 271.95, 
    271.95, 272.05, 272.55, 272.75, 272.75, 272.85, 272.95, 272.35, 272.65, 
    273.85, 274.45, 273.15, 273.15, 273.35, 272.85, 272.55, 272.75, 272.65, 
    273.05, 273.15, 273.35, 273.65, 274.05, 274.35, 274.35, 274.65, 274.65, 
    274.55, 274.35, 273.25, 273.35, 273.55, 273.65, 275.25, 274.75, 273.15, 
    272.45, 272.65, 272.85, 273.05, 273.95, 273.55, 273.75, 273.55, 273.55, 
    273.55, 273.75, 273.75, 274.25, 274.35, 274.45, 274.25, 274.15, 273.95, 
    274.15, 275.15, 274.15, 273.15, 273.45, 273.05, 273.15, 273.15, 272.95, 
    273.05, 272.75, 272.65, 272.55, 272.55, 271.95, 272.15, 272.55, 272.85, 
    273.25, 273.65, 273.95, 273.85, 273.55, 273.65, 274.15, 273.95, 274.45, 
    274.15, 274.05, 273.95, 274.55, 273.95, 274.15, 273.85, 273.75, 273.85, 
    273.55, 273.65, 273.55, 273.75, 273.45, 273.45, 273.55, 273.95, 276.25, 
    274.65, 274.75, 274.65, 275.45, 275.55, 275.45, 275.65, 276.65, 274.55, 
    275.15, 275.25, 275.05, 274.35, 274.35, 273.75, 273.55, 273.25, 273.15, 
    272.95, 272.95, 272.75, 272.75, 272.95, 272.85, 273.35, 273.45, 273.95, 
    274.15, 274.25, 274.25, 274.25, 274.25, 274.05, 274.25, 274.25, 274.15, 
    274.15, 274.05, 273.85, 273.75, 273.65, 273.35, 273.45, 273.35, 273.35, 
    273.25, 273.65, 273.55, 273.55, 273.75, 274.05, 273.95, 274.25, 274.25, 
    274.15, 274.65, 274.35, 274.35, 274.45, 274.15, 273.95, 273.75, 273.15, 
    272.85, 272.95, 272.75, 272.95, 272.75, 272.75, 272.45, 272.35, 272.05, 
    271.95, 271.95, 272.05, 271.95, 271.85, 271.75, 272.15, 271.75, 271.45, 
    271.55, 271.75, 271.25, 271.35, 271.35, 271.15, 271.25, 271.15, 271.25, 
    271.15, 271.05, 271.25, 271.15, 271.15, 270.95, 270.95, 271.25, 271.15, 
    271.15, 270.95, 270.45, 269.85, 269.55, 269.35, 269.25, 269.15, 268.95, 
    268.85, 268.75, 268.75, 268.65, 268.35, 268.35, 268.05, 267.85, 267.85, 
    268.15, 267.85, 267.95, 268.65, 268.55, 269.45, 270.25, 270.85, 270.55, 
    270.65, 270.85, 271.55, 271.55, 271.45, 271.55, 271.25, 271.05, 270.75, 
    270.65, 270.65, 269.95, 269.95, 269.75, 270.25, 270.15, 269.95, 271.25, 
    271.15, 271.35, 271.65, 272.75, 272.65, 272.25, 272.55, 272.35, 271.95, 
    271.75, 272.35, 272.45, 272.25, 272.15, 271.95, 271.05, 271.05, 270.75, 
    270.65, 270.95, 270.75, 271.05, 270.35, 271.05, 271.95, 272.05, 271.75, 
    271.25, 271.15, 272.05, 272.05, 271.85, 271.65, 271.35, 270.75, 271.05, 
    271.85, 271.45, 270.65, 270.65, 270.75, 271.05, 270.45, 269.85, 269.95, 
    269.55, 269.15, 269.65, 269.95, 270.45, 269.95, 270.15, 270.35, 270.25, 
    270.25, 270.15, 270.05, 270.05, 270.15, 269.35, 268.65, 267.75, 267.25, 
    266.75, 266.45, 265.75, 265.65, 265.95, 265.75, 266.15, 266.95, 267.15, 
    267.05, 267.15, 267.45, 267.15, 267.55, 267.05, 267.15, 267.25, 267.45, 
    267.45, 267.15, 267.65, 267.65, 267.85, 268.15, 268.75, 268.95, 269.15, 
    269.15, 269.15, 270.15, 270.15, 270.15, 270.45, 270.65, 270.95, 271.45, 
    271.55, 271.65, 271.35, 272.25, 272.45, 272.15, 272.45, 272.25, 271.45, 
    270.85, 270.55, 270.55, 269.15, 268.45, 268.25, 267.85, 268.15, 269.35, 
    269.65, 270.25, 270.95, 271.25, 271.25, 271.45, 271.65, 272.25, 272.15, 
    272.55, 272.95, 272.75, 272.85, 273.15, 272.85, 272.55, 272.95, 272.55, 
    272.15, 271.35, 271.65, 271.65, 271.25, 271.35, 271.35, 271.35, 272.05, 
    272.75, 272.65, 272.35, 273.45, 273.25, 274.05, 273.55, 273.05, 272.45, 
    272.25, 272.55, 272.55, 272.35, 272.35, 271.95, 271.55, 271.55, 271.45, 
    271.85, 271.85, 272.15, 272.65, 272.75, 272.95, 273.35, 274.05, 274.55, 
    275.45, 275.85, 276.45, 276.65, 276.65, 276.95, 276.05, 276.25, 275.55, 
    275.45, 274.95, 274.95, 274.15, 274.05, 273.55, 273.45, 273.25, 273.75, 
    274.25, 273.85, 274.85, 274.85, 274.85, 275.35, 276.25, 277.55, 276.45, 
    275.45, 275.45, 275.35, 276.05, 275.65, 275.05, 274.85, 275.65, 275.55, 
    276.05, 276.05, 276.35, 277.15, 277.25, 277.05, 275.15, 275.05, 275.35, 
    275.45, 275.35, 276.15, 279.25, 277.75, 278.35, 278.75, 278.95, 278.35, 
    277.75, 277.15, 277.55, 278.15, 276.35, 276.75, 277.55, 276.75, 276.25, 
    275.95, 275.65, 275.55, 274.75, 274.65, 274.65, 274.85, 275.05, 275.15, 
    275.15, 275.05, 275.55, 275.55, 275.75, 275.75, 276.55, 276.65, 276.45, 
    276.25, 275.15, 274.75, 274.35, 273.75, 273.05, 273.05, 273.95, 274.95, 
    274.85, 274.75, 275.55, 275.95, 275.65, 276.05, 275.75, 274.65, 274.55, 
    275.35, 275.15, 275.35, 274.45, 274.25, 273.85, 273.55, 273.15, 273.15, 
    271.85, 271.15, 271.35, 271.25, 271.25, 271.15, 271.35, 271.65, 273.25, 
    272.45, 274.15, 274.75, 274.25, 274.95, 275.45, 276.55, 274.85, 275.05, 
    275.45, 275.05, 275.25, 275.25, 274.85, 275.45, 275.45, 275.05, 274.65, 
    274.35, 274.05, 273.95, 273.55, 274.05, 274.65, 275.15, 274.95, 274.55, 
    275.25, 275.75, 276.25, 275.85, 276.05, 275.75, 275.75, 275.15, 275.25, 
    275.55, 275.35, 275.45, 275.05, 274.95, 274.85, 274.95, 274.95, 274.85, 
    275.15, 275.15, 275.15, 275.45, 274.95, 275.05, 274.75, 275.05, 275.35, 
    275.05, 275.05, 276.15, 275.75, 275.85, 276.25, 275.35, 274.55, 274.65, 
    274.85, 274.95, 274.95, 275.25, 275.05, 275.05, 275.35, 275.55, 275.65, 
    275.75, 275.85, 275.95, 276.05, 276.45, 276.85, 276.85, 276.65, 276.05, 
    276.15, 275.55, 275.55, 275.35, 275.65, 275.55, 275.35, 275.45, 275.25, 
    274.85, 274.65, 275.25, 275.25, 275.55, 276.05, 276.85, 276.55, 276.55, 
    276.35, 276.45, 276.55, 276.55, 276.45, 276.55, 276.25, 276.65, 276.45, 
    276.45, 276.25, 275.95, 275.85, 275.65, 275.65, 275.55, 275.55, 275.85, 
    276.05, 276.15, 276.35, 276.65, 276.75, 276.75, 276.95, 277.05, 277.05, 
    277.05, 276.35, 276.75, 276.05, 276.25, 276.25, 276.05, 275.75, 275.65, 
    275.15, 275.05, 275.25, 275.15, 275.65, 275.75, 275.65, 275.55, 276.15, 
    276.35, 276.45, 277.05, 277.85, 277.95, 277.15, 277.45, 277.65, 278.25, 
    278.35, 278.15, 278.15, 278.15, 277.55, 277.15, 276.15, 275.85, 275.85, 
    275.95, 276.05, 277.25, 277.35, 278.05, 278.65, 279.45, 279.25, 279.55, 
    279.55, 279.55, 280.75, 279.05, 279.15, 279.55, 279.65, 279.25, 279.55, 
    279.15, 278.65, 277.55, 277.75, 277.35, 277.05, 276.75, 277.45, 279.45, 
    277.85, 278.45, 278.65, 279.45, 279.55, 279.55, 280.35, 280.15, 280.35, 
    278.75, 278.45, 277.95, 278.25, 278.15, 277.55, 276.95, 276.75, 277.95, 
    277.85, 277.25, 276.85, 277.15, 277.45, 277.75, 277.95, 278.05, 278.25, 
    277.65, 277.55, 277.85, 277.95, 277.95, 277.95, 278.65, 278.55, 277.85, 
    278.35, 277.65, 277.65, 277.45, 276.95, 276.85, 276.95, 276.85, 276.85, 
    275.85, 276.45, 276.15, 276.15, 275.75, 276.25, 276.85, 277.25, 277.35, 
    277.65, 277.95, 278.15, 278.65, 278.55, 278.55, 277.95, 278.05, 277.35, 
    277.45, 276.95, 276.85, 276.75, 276.35, 276.85, 276.85, 276.75, 276.35, 
    276.25, 276.25, 276.65, 276.75, 277.25, 277.65, 277.95, 278.35, 278.55, 
    278.65, 278.85, 279.05, 279.15, 277.85, 277.85, 278.15, 279.65, 278.75, 
    278.25, 278.35, 277.85, 278.05, 278.55, 279.65, 277.85, 278.05, 277.95, 
    277.45, 278.15, 277.15, 277.15, 279.05, 279.25, 280.35, 279.75, 280.65, 
    280.45, 279.85, 279.15, 279.65, 278.15, 278.25, 277.95, 277.55, 276.95, 
    277.45, 277.85, 277.55, 278.05, 278.05, 277.95, 278.75, 278.05, 279.05, 
    279.55, 279.05, 278.75, 278.45, 279.85, 279.15, 278.65, 277.95, 277.95, 
    277.35, 276.85, 277.15, 276.25, 276.45, 276.75, 276.75, 276.35, 276.05, 
    276.15, 276.05, 276.25, 276.95, 276.95, 276.75, 276.35, 276.15, 276.75, 
    275.95, 276.75, 277.95, 278.15, 277.95, 277.35, 277.35, 277.55, 277.15, 
    277.25, 277.55, 277.85, 276.95, 276.95, 277.25, 278.25, 278.15, 279.15, 
    280.05, 279.05, 280.55, 279.25, 279.45, 279.05, 279.05, 277.95, 278.95, 
    279.25, 279.15, 277.45, 277.85, 278.05, 278.25, 278.35, 278.15, 277.85, 
    277.85, 278.15, 278.55, 278.85, 279.45, 280.05, 280.15, 279.15, 279.55, 
    280.55, 280.35, 281.25, 281.35, 281.05, 281.75, 282.05, 282.35, 281.85, 
    281.55, 280.75, 280.75, 280.65, 280.25, 278.95, 278.65, 279.95, 279.45, 
    280.05, 279.95, 280.05, 280.35, 280.75, 281.05, 281.05, 281.75, 281.45, 
    282.45, 282.65, 281.65, 282.05, 281.75, 281.45, 280.75, 279.95, 279.65, 
    279.55, 279.45, 279.15, 278.85, 279.65, 279.95, 279.65, 279.95, 280.55, 
    280.45, 280.95, 281.15, 281.45, 281.35, 282.15, 280.95, 280.95, 282.45, 
    281.25, 281.15, 280.05, 280.45, 280.35, 279.85, 279.45, 279.85, 279.25, 
    278.65, 279.05, 279.25, 279.25, 279.55, 279.85, 280.75, 281.05, 281.85, 
    282.05, 282.35, 281.75, 281.85, 281.75, 282.65, 282.45, 282.25, 282.55, 
    282.05, 282.55, 282.85, 281.95, 282.15, 282.05, 282.05, 281.65, 281.85, 
    281.95, 281.95, 281.95, 281.95, 282.55, 283.05, 283.25, 283.45, 283.35, 
    283.25, 282.95, 283.35, 282.25, 282.65, 282.45, 281.55, 281.35, 281.25, 
    281.85, 281.75, 281.95, 281.95, 281.55, 281.05, 281.45, 281.15, 281.95, 
    282.25, 282.45, 282.65, 283.25, 284.45, 284.55, 284.05, 283.95, 283.75, 
    283.55, 283.35, 283.05, 281.95, 281.95, 281.65, 281.55, 281.15, 280.85, 
    280.95, 281.05, 280.85, 280.55, 280.55, 281.05, 281.35, 280.95, 280.95, 
    281.35, 281.65, 281.65, 282.05, 281.75, 281.65, 280.75, 280.85, 280.65, 
    280.35, 279.85, 279.55, 279.35, 279.15, 279.05, 279.05, 279.45, 279.25, 
    279.75, 279.65, 279.45, 279.75, 280.05, 280.45, 279.85, 279.25, 279.35, 
    279.25, 279.25, 279.25, 279.15, 278.95, 279.25, 279.25, 279.15, 279.15, 
    278.85, 279.15, 279.05, 278.55, 278.35, 278.55, 278.65, 278.55, 278.45, 
    278.05, 277.85, 277.75, 277.75, 277.85, 277.75, 277.55, 277.15, 277.55, 
    277.55, 276.95, 276.95, 275.95, 276.05, 275.45, 274.25, 273.15, 273.55, 
    273.35, 274.05, 274.65, 275.25, 275.25, 275.75, 276.65, 276.45, 276.55, 
    276.65, 276.75, 276.95, 277.55, 277.85, 278.05, 277.95, 277.95, 277.95, 
    278.25, 277.75, 277.85, 277.35, 276.85, 278.05, 277.45, 277.25, 276.75, 
    277.45, 276.25, 275.45, 276.35, 277.25, 277.85, 277.85, 278.15, 278.35, 
    278.35, 278.95, 279.05, 279.15, 279.45, 279.45, 279.05, 278.65, 277.55, 
    277.85, 278.65, 278.65, 279.05, 279.55, 279.85, 280.15, 280.75, 280.85, 
    280.85, 280.75, 280.35, 280.55, 281.55, 281.95, 282.55, 280.65, 280.75, 
    280.65, 280.15, 279.85, 281.35, 281.35, 281.05, 281.55, 281.75, 281.85, 
    282.55, 282.35, 281.85, 282.95, 283.95, 284.05, 284.35, 284.65, 284.15, 
    284.45, 285.15, 285.35, 285.85, 285.85, 285.15, 283.65, 284.85, 285.75, 
    286.55, 285.85, 285.85, 285.65, 285.55, 285.75, 285.75, 285.45, 284.65, 
    284.85, 283.75, 284.05, 283.65, 283.45, 284.15, 283.65, 282.95, 282.65, 
    284.35, 284.05, 283.45, 283.85, 284.65, 284.05, 282.55, 282.15, 282.15, 
    281.05, 281.25, 281.25, 282.25, 280.45, 279.75, 279.65, 279.25, 279.45, 
    279.05, 278.95, 278.95, 279.15, 279.25, 279.55, 279.45, 279.35, 279.65, 
    279.85, 279.45, 279.05, 278.65, 279.05, 278.75, 278.65, 278.15, 277.55, 
    277.25, 278.45, 278.85, 279.25, 278.75, 279.25, 280.65, 281.35, 281.65, 
    281.95, 282.55, 282.45, 283.25, 284.05, 283.95, 284.35, 284.35, 284.75, 
    283.35, 282.85, 281.75, 281.75, 282.35, 283.55, 284.65, 283.85, 282.95, 
    284.25, 284.85, 284.85, 284.25, 284.65, 285.35, 283.15, 282.95, 283.15, 
    283.85, 284.35, 283.05, 284.35, 283.25, 283.35, 283.35, 282.55, 282.75, 
    283.65, 281.25, 280.65, 281.55, 281.15, 282.35, 282.85, 282.85, 283.25, 
    283.45, 283.85, 283.25, 284.85, 282.85, 283.35, 283.15, 284.15, 286.55, 
    285.35, 283.85, 287.15, 286.65, 285.25, 284.35, 283.95, 283.85, 282.95, 
    282.25, 282.75, 282.55, 282.25, 283.35, 283.55, 284.75, 285.75, 286.25, 
    286.35, 285.45, 285.45, 284.15, 285.15, 283.85, 282.35, 282.65, 282.75, 
    283.65, 283.05, 282.95, 282.75, 282.95, 283.15, 283.05, 283.25, 283.45, 
    283.45, 284.95, 285.75, 286.25, 286.35, 286.85, 286.85, 286.95, 286.85, 
    287.45, 288.15, 287.85, 287.65, 283.35, 283.55, 284.25, 283.95, 282.85, 
    282.25, 282.85, 283.05, 281.95, 281.65, 281.95, 282.15, 282.55, 283.65, 
    281.85, 281.85, 281.75, 282.25, 282.05, 282.25, 282.15, 283.05, 283.05, 
    282.85, 282.65, 283.85, 282.95, 283.35, 282.65, 282.05, 281.55, 280.95, 
    281.05, 281.15, 281.55, 281.25, 281.35, 281.15, 280.95, 280.85, 280.65, 
    280.85, 281.05, 281.05, 281.45, 281.35, 281.45, 281.35, 281.15, 280.95, 
    280.85, 280.85, 280.75, 280.85, 280.65, 280.75, 280.55, 280.65, 280.75, 
    280.75, 280.75, 280.75, 280.85, 280.85, 280.85, 280.95, 281.05, 281.05, 
    281.55, 281.85, 281.55, 281.25, 281.35, 281.25, 280.75, 281.35, 280.95, 
    280.15, 279.75, 279.55, 279.25, 279.25, 279.35, 279.95, 280.05, 280.65, 
    280.85, 280.75, 280.25, 280.45, 280.75, 280.85, 280.55, 280.65, 280.85, 
    280.75, 280.65, 280.45, 280.25, 280.15, 279.85, 279.55, 279.65, 279.85, 
    279.55, 279.65, 279.65, 279.85, 279.55, 279.05, 278.55, 278.25, 278.75, 
    278.95, 278.95, 278.85, 279.35, 280.15, 280.25, 279.45, 278.65, 279.15, 
    278.95, 278.85, 278.55, 278.65, 278.55, 278.75, 278.75, 278.75, 279.05, 
    279.25, 279.85, 280.05, 279.95, 280.05, 280.15, 280.15, 280.75, 280.35, 
    280.55, 281.15, 281.35, 281.05, 280.65, 280.15, 280.05, 279.95, 280.05, 
    279.85, 279.75, 279.75, 279.75, 279.75, 279.65, 279.65, 280.15, 280.05, 
    280.25, 280.35, 280.55, 280.65, 280.85, 280.75, 281.05, 280.75, 280.85, 
    280.75, 280.75, 280.65, 280.35, 280.35, 280.35, 280.25, 280.15, 280.15, 
    280.05, 280.15, 280.15, 280.35, 280.25, 280.45, 280.85, 280.85, 280.45, 
    280.65, 280.65, 280.75, 280.95, 281.15, 281.35, 280.85, 280.55, 280.05, 
    280.15, 279.75, 279.75, 279.65, 279.75, 279.55, 279.55, 279.65, 279.85, 
    279.95, 279.95, 280.05, 280.55, 280.95, 281.15, 281.35, 281.25, 281.05, 
    281.55, 281.15, 281.25, 281.55, 281.15, 281.35, 280.85, 280.35, 280.15, 
    280.05, 279.85, 279.75, 279.85, 279.95, 280.45, 280.35, 280.25, 280.25, 
    280.55, 280.55, 280.35, 280.25, 280.55, 280.75, 280.55, 282.45, 281.35, 
    280.55, 280.05, 280.15, 280.15, 280.35, 280.05, 278.85, 278.75, 278.65, 
    278.85, 278.95, 279.15, 279.35, 279.45, 279.25, 280.15, 279.95, 280.65, 
    280.75, 281.35, 280.95, 281.35, 281.25, 281.25, 281.15, 280.85, 280.85, 
    280.95, 280.95, 280.65, 280.95, 280.95, 281.05, 281.05, 280.55, 280.75, 
    280.65, 280.85, 281.05, 281.65, 281.75, 281.45, 281.55, 281.65, 281.65, 
    281.65, 281.65, 281.55, 280.95, 281.55, 281.55, 282.05, 281.45, 281.25, 
    281.15, 280.95, 280.65, 280.15, 280.05, 279.75, 279.55, 279.75, 280.25, 
    279.85, 279.95, 280.55, 280.35, 280.25, 279.75, 279.35, 280.35, 280.65, 
    280.45, 280.55, 280.35, 280.55, 280.55, 280.25, 280.15, 279.85, 279.85, 
    279.95, 280.05, 280.15, 280.15, 280.75, 280.95, 281.65, 281.75, 281.75, 
    280.95, 281.75, 281.15, 281.35, 281.35, 280.85, 280.85, 280.85, 280.75, 
    280.55, 280.55, 280.75, 280.65, 280.75, 280.45, 280.05, 280.05, 280.45, 
    281.15, 281.35, 281.65, 282.45, 282.35, 282.35, 282.35, 282.25, 281.95, 
    281.65, 281.55, 281.95, 282.05, 281.85, 281.45, 281.45, 281.55, 281.45, 
    281.15, 281.25, 281.25, 281.15, 281.05, 281.05, 281.35, 281.85, 281.85, 
    281.85, 282.15, 282.05, 281.55, 283.05, 283.05, 283.85, 283.85, 283.85, 
    282.65, 282.55, 282.25, 281.85, 281.75, 280.95, 280.85, 280.75, 279.95, 
    279.45, 279.85, 280.45, 280.85, 280.25, 281.15, 281.35, 282.15, 282.55, 
    282.85, 283.25, 283.05, 283.25, 283.25, 282.95, 282.25, 282.25, 282.35, 
    281.95, 281.35, 281.15, 281.25, 280.85, 280.75, 280.55, 280.45, 280.85, 
    280.85, 280.95, 281.95, 281.85, 282.55, 282.65, 282.85, 283.25, 283.65, 
    284.15, 284.05, 284.65, 284.75, 284.95, 283.75, 282.75, 282.05, 281.95, 
    281.85, 281.35, 281.05, 280.45, 281.25, 281.85, 282.05, 282.25, 282.85, 
    283.85, 283.45, 283.35, 284.95, 285.05, 284.95, 284.95, 285.35, 285.05, 
    285.15, 285.05, 284.65, 284.55, 282.35, 282.05, 281.75, 281.25, 281.15, 
    281.45, 281.55, 281.65, 282.25, 282.55, 283.45, 284.75, 284.95, 285.75, 
    285.95, 286.85, 287.15, 287.45, 287.35, 287.65, 287.25, 287.75, 287.65, 
    286.45, 285.75, 285.45, 284.85, 284.15, 282.75, 283.05, 281.65, 282.05, 
    282.75, 282.95, 283.05, 283.45, 283.45, 283.35, 283.15, 283.65, 283.45, 
    283.45, 283.45, 282.75, 282.45, 282.55, 282.55, 282.65, 281.75, 282.25, 
    282.25, 282.15, 282.05, 282.15, 282.15, 281.75, 281.85, 282.15, 282.15, 
    282.45, 282.05, 281.55, 282.15, 281.65, 281.85, 281.65, 281.85, 282.05, 
    282.15, 282.65, 282.05, 281.95, 281.95, 281.35, 281.35, 281.25, 280.95, 
    281.25, 281.45, 280.35, 280.65, 280.55, 280.75, 281.05, 281.15, 281.45, 
    281.75, 282.25, 282.45, 283.75, 285.85, 286.35, 286.55, 286.45, 285.85, 
    286.05, 284.15, 283.45, 282.45, 281.95, 281.45, 281.05, 280.55, 281.85, 
    281.75, 281.55, 280.15, 279.95, 279.85, 280.25, 280.35, 280.55, 280.65, 
    280.95, 281.25, 281.65, 281.65, 281.85, 281.95, 281.85, 282.25, 281.85, 
    281.75, 281.65, 281.55, 281.45, 281.25, 280.75, 280.55, 281.05, 281.25, 
    281.35, 281.65, 282.55, 282.55, 282.55, 283.15, 283.35, 283.45, 284.35, 
    284.15, 284.35, 283.75, 282.85, 282.55, 282.05, 281.75, 281.15, 280.75, 
    280.55, 280.85, 281.25, 281.05, 280.95, 281.55, 281.25, 282.15, 282.15, 
    282.95, 283.45, 283.95, 284.35, 283.95, 283.85, 282.95, 282.75, 281.75, 
    281.65, 281.45, 281.15, 280.85, 280.55, 280.55, 280.45, 279.85, 280.05, 
    280.05, 280.05, 279.95, 279.95, 279.75, 280.05, 280.25, 280.35, 280.55, 
    280.95, 280.95, 281.25, 281.55, 281.75, 282.05, 281.95, 281.85, 281.65, 
    281.95, 281.55, 281.25, 280.85, 280.65, 280.95, 280.75, 281.25, 281.95, 
    282.35, 282.35, 282.85, 283.45, 283.25, 283.65, 283.95, 283.95, 284.85, 
    285.15, 284.65, 283.95, 283.55, 282.55, 282.25, 281.15, 280.95, 279.65, 
    280.25, 279.65, 280.45, 281.85, 281.25, 282.35, 282.85, 282.65, 282.25, 
    282.95, 283.75, 283.15, 284.35, 284.35, 283.75, 282.65, 281.95, 281.55, 
    280.45, 279.75, 279.15, 279.35, 278.75, 278.65, 278.45, 278.45, 278.75, 
    278.95, 279.65, 279.95, 280.45, 280.45, 280.85, 280.95, 280.65, 280.75, 
    281.55, 280.95, 281.55, 281.55, 281.35, 281.55, 281.45, 281.15, 281.15, 
    281.15, 280.85, 281.35, 281.05, 281.05, 281.25, 281.05, 280.95, 280.95, 
    280.95, 282.15, 282.75, 282.05, 282.65, 282.45, 282.55, 282.55, 283.05, 
    282.65, 282.15, 281.75, 281.85, 281.65, 280.95, 280.45, 279.85, 279.85, 
    279.85, 279.95, 280.05, 280.45, 280.55, 280.65, 280.85, 280.45, 280.35, 
    280.25, 280.35, 279.95, 280.15, 280.25, 280.35, 280.65, 280.75, 280.65, 
    280.25, 280.05, 279.65, 279.45, 278.95, 278.35, 277.85, 277.25, 277.35, 
    277.95, 278.05, 278.75, 278.75, 278.35, 279.15, 279.15, 279.25, 279.25, 
    279.65, 279.25, 279.85, 279.75, 279.45, 278.45, 279.25, 277.85, 277.45, 
    277.55, 277.65, 277.65, 277.55, 277.35, 276.85, 277.35, 277.45, 278.05, 
    278.05, 278.75, 278.55, 278.75, 279.55, 279.65, 279.85, 280.05, 279.75, 
    280.05, 278.85, 278.75, 279.35, 278.75, 278.55, 277.75, 277.45, 277.45, 
    277.25, 278.15, 277.75, 277.75, 277.85, 277.95, 278.85, 279.05, 278.95, 
    279.05, 279.65, 278.95, 279.35, 278.85, 278.55, 278.45, 278.55, 278.35, 
    278.25, 277.85, 277.45, 277.65, 277.75, 277.75, 277.55, 277.25, 277.65, 
    277.35, 277.65, 277.95, 277.75, 278.45, 278.45, 278.45, 279.35, 280.05, 
    280.65, 280.55, 280.15, 280.35, 279.95, 279.65, 280.65, 280.05, 279.45, 
    279.25, 279.35, 279.05, 278.85, 279.05, 278.85, 278.35, 278.05, 278.05, 
    277.95, 277.95, 278.15, 278.65, 278.95, 279.45, 279.65, 279.35, 279.05, 
    278.85, 278.55, 278.45, 278.05, 278.05, 277.55, 277.55, 277.45, 276.95, 
    276.95, 276.95, 276.95, 276.95, 277.15, 277.05, 276.95, 276.85, 276.45, 
    276.45, 276.65, 276.85, 276.95, 276.75, 276.45, 276.15, 275.95, 275.75, 
    275.25, 275.05, 274.55, 274.35, 274.45, 274.45, 273.95, 274.25, 274.95, 
    276.05, 276.25, 276.35, 276.85, 276.65, 277.15, 277.75, 277.65, 277.55, 
    277.45, 278.25, 278.15, 278.15, 278.15, 277.45, 276.95, 276.75, 276.85, 
    276.75, 276.75, 276.75, 276.45, 276.55, 276.35, 276.75, 276.95, 277.05, 
    277.15, 277.25, 277.65, 278.65, 278.95, 278.75, 278.85, 278.85, 278.75, 
    278.35, 279.05, 278.05, 277.95, 277.85, 277.75, 277.45, 277.25, 276.85, 
    276.55, 276.65, 276.95, 277.15, 277.35, 277.55, 277.85, 278.15, 278.55, 
    279.05, 279.05, 278.85, 278.75, 278.65, 278.35, 278.15, 278.35, 278.35, 
    278.15, 277.95, 277.75, 277.45, 277.15, 277.25, 276.85, 276.85, 276.85, 
    276.85, 277.55, 277.65, 278.05, 278.75, 278.75, 279.05, 278.35, 279.05, 
    278.95, 278.65, 278.05, 277.95, 278.15, 278.25, 278.35, 278.45, 278.45, 
    278.25, 278.05, 278.15, 277.85, 277.25, 277.75, 277.55, 278.15, 278.35, 
    278.75, 279.05, 279.65, 280.05, 279.85, 280.45, 279.95, 279.65, 279.45, 
    279.55, 279.15, 279.25, 278.85, 278.85, 278.55, 278.45, 278.25, 278.05, 
    277.85, 278.75, 277.95, 277.05, 276.65, 277.05, 277.15, 276.75, 277.05, 
    277.75, 278.15, 277.75, 277.45, 277.55, 278.15, 277.35, 276.75, 276.05, 
    275.35, 274.95, 274.95, 274.65, 273.85, 273.65, 273.65, 273.65, 273.55, 
    273.85, 273.95, 274.85, 275.25, 275.45, 275.85, 276.25, 276.45, 276.85, 
    277.75, 278.35, 277.85, 277.65, 277.55, 277.55, 277.35, 276.95, 276.45, 
    276.55, 276.05, 275.95, 276.25, 275.55, 276.15, 276.75, 276.05, 276.45, 
    276.85, 276.95, 277.15, 277.55, 277.65, 277.95, 278.15, 277.85, 277.65, 
    277.55, 277.15, 276.95, 275.95, 275.75, 275.75, 275.85, 275.75, 275.95, 
    276.15, 276.25, 277.45, 277.65, 276.75, 276.15, 276.45, 276.75, 277.05, 
    276.85, 276.95, 276.95, 276.95, 277.35, 277.75, 278.15, 277.85, 277.95, 
    277.85, 277.35, 276.95, 276.75, 276.35, 276.15, 275.95, 275.85, 275.85, 
    276.05, 276.35, 278.05, 276.65, 277.05, 277.15, 277.65, 278.35, 278.55, 
    278.45, 278.55, 278.65, 278.65, 278.45, 278.35, 278.35, 278.25, 278.05, 
    277.95, 277.65, 277.65, 277.65, 277.75, 278.05, 278.45, 277.45, 278.25, 
    278.55, 278.75, 279.25, 279.35, 279.95, 280.55, 280.35, 279.75, 279.75, 
    278.75, 278.35, 276.45, 275.85, 275.85, 276.35, 276.75, 277.15, 277.55, 
    279.15, 279.65, 279.25, 276.15, 275.85, 277.95, 277.95, 278.25, 278.25, 
    279.05, 278.75, 278.35, 278.35, 278.35, 278.65, 278.75, 279.15, 279.35, 
    279.05, 278.65, 279.45, 279.95, 279.45, 279.65, 279.75, 279.75, 279.65, 
    279.55, 277.95, 278.75, 280.05, 280.25, 280.25, 280.55, 280.45, 280.05, 
    279.65, 279.65, 279.45, 279.55, 279.15, 279.55, 279.85, 279.35, 279.05, 
    278.65, 278.85, 279.25, 279.15, 278.95, 279.45, 280.05, 279.55, 279.45, 
    279.45, 280.35, 280.35, 280.85, 281.05, 280.95, 281.25, 281.25, 281.15, 
    281.05, 280.95, 281.25, 281.95, 282.15, 282.25, 282.65, 282.05, 282.75, 
    282.25, 281.15, 280.85, 280.95, 280.75, 281.25, 280.95, 281.45, 281.35, 
    282.75, 282.45, 281.25, 283.75, 282.15, 282.65, 282.45, 282.65, 281.95, 
    282.35, 281.75, 282.35, 281.75, 281.55, 281.65, 281.05, 280.65, 280.55, 
    280.45, 280.35, 279.95, 279.75, 279.75, 279.65, 279.25, 279.75, 279.85, 
    280.45, 280.35, 280.25, 280.25, 280.25, 279.45, 279.25, 279.25, 279.15, 
    278.85, 278.65, 278.45, 278.25, 278.15, 277.95, 277.95, 278.05, 278.55, 
    278.15, 278.85, 279.35, 278.95, 279.55, 279.65, 280.15, 280.25, 280.05, 
    279.85, 280.25, 280.05, 279.75, 279.45, 279.05, 278.25, 278.15, 277.85, 
    278.05, 277.85, 277.35, 277.05, 277.85, 278.75, 279.15, 279.75, 281.15, 
    281.15, 281.25, 280.85, 281.55, 279.95, 280.15, 279.55, 279.25, 279.05, 
    278.65, 278.55, 278.05, 277.55, 277.25, 276.95, 277.35, 277.25, 277.25, 
    277.55, 277.55, 277.55, 277.55, 278.05, 278.05, 278.35 ;

 air_pressure_at_sea_level = 100710, 100720, 100680, 100680, 100690, 100690, 
    100680, 100670, 100730, 100720, 100740, 100760, 100760, 100760, 100760, 
    100760, 100760, 100770, 100790, 100800, 100700, 100710, 100690, 100690, 
    100670, 100670, 100660, 100650, 100650, 100640, 100640, 100630, 100670, 
    100670, 100660, 100660, 100660, 100650, 100620, 100600, 100590, 100570, 
    100540, 100530, 100480, 100480, 100470, 100460, 100460, 100460, 100430, 
    100400, 100370, 100340, 100320, 100330, 100350, 100340, 100330, 100340, 
    100340, 100340, 100330, 100330, 100310, 100320, 100340, 100350, 100360, 
    100380, 100400, 100270, 100280, 100470, 100470, 100370, 100400, 100400, 
    100440, 100450, 100500, 100540, 100560, 100600, 100610, 100640, 100640, 
    100650, 100670, 100700, 100690, 100670, 100690, 100690, 100710, 100740, 
    100750, 100730, 100750, 100770, 100770, 100770, 100800, 100800, 100840, 
    100880, 100910, 100940, 100970, 100980, 100990, 101010, 101030, 101030, 
    101040, 101030, 101030, 101030, 101060, 101060, 101070, 101070, 101080, 
    101060, 101040, 101030, 101020, 100990, 101010, 101010, 101000, 101030, 
    101020, 101010, 101030, 101020, 101040, 101060, 101100, 101130, 101180, 
    101240, 101290, 101360, 101420, 101480, 101530, 101590, 101650, 101710, 
    101750, 101790, 101850, 101890, 101900, 101970, 101990, 102010, 102040, 
    102070, 102080, 102060, 102080, 102090, _, 102230, 102260, 102310, 
    102340, 102370, 102410, 102440, 102450, 102460, 102460, 102500, 102530, 
    102550, 102590, 102640, 102620, 102620, 102630, 102660, 102650, 102610, 
    102590, 102580, 102540, 102590, 102580, 102560, 102610, 102600, 102580, 
    102560, 102560, 102560, 102470, 102450, 102430, 102410, 102410, 102410, 
    102420, 102430, 102430, 102410, 102410, 102380, 102370, 102370, 102390, 
    102440, 102460, 102510, 102520, 102540, 102570, 102590, 102570, 102590, 
    102600, 102640, 102660, 102700, 102730, 102780, 102820, 102860, 102870, 
    102900, 102930, 102960, 102950, 102990, 103030, 103050, 103090, 103160, 
    103180, 103220, 103250, 103270, 103290, 103310, 103350, 103360, 103390, 
    103400, 103450, 103470, 103480, 103500, 103480, 103500, 103510, 103510, 
    103510, 103510, 103490, 103500, 103480, 103470, 103460, 103430, 103410, 
    103430, 103440, 103410, 103400, 103390, 103400, 103420, 103410, 103400, 
    103420, 103420, 103400, 103390, 103390, 103360, 103360, 103370, 103360, 
    103370, 103370, 103400, 103440, 103440, 103440, 103440, 103450, 103450, 
    103460, 103440, 103440, 103460, 103490, 103510, 103510, 103490, 103500, 
    103530, 103530, 103540, 103510, 103510, 103500, 103480, 103500, 103500, 
    103500, 103490, 103490, 103470, 103480, 103480, 103480, 103500, 103510, 
    103520, 103540, 103550, 103590, 103580, 103580, 103610, 103610, 103630, 
    103640, 103650, 103650, 103640, 103680, 103710, 103730, 103740, 103750, 
    103740, 103700, 103690, 103630, 103600, 103590, 103570, 103550, 103510, 
    103480, 103440, 103380, 103340, 103310, 103260, 103230, 103190, 103120, 
    103080, 103050, 103030, 102990, 102970, 102920, 102870, 102810, 102770, 
    102720, 102670, 102620, 102580, 102530, 102500, 102450, 102420, 102370, 
    102360, 102350, 102340, 102320, 102310, 102340, 102370, 102380, 102410, 
    102450, 102470, 102460, 102480, 102480, 102490, 102470, 102460, 102460, 
    102470, 102460, 102480, 102490, 102470, 102480, 102460, 102450, 102450, 
    102440, 102430, 102430, 102400, 102400, 102400, 102410, 102400, 102380, 
    102360, 102340, 102330, 102330, 102320, 102320, 102320, 102320, 102320, 
    102310, 102290, 102290, 102270, 102250, 102220, 102200, 102150, 102140, 
    102110, 102120, 102130, 102130, 102090, 102060, 102040, 102020, 101990, 
    101960, 101950, 101930, 101910, 101890, 101860, 101850, 101830, 101790, 
    101750, 101710, 101700, 101690, 101650, 101620, 101620, 101620, 101610, 
    101590, 101570, 101570, 101530, 101510, 101500, 101460, 101450, 101450, 
    101410, 101380, 101340, 101320, 101260, 101210, 101160, 101140, 101110, 
    101080, 101050, 101030, 101010, 101000, 101010, 101000, 100980, 100980, 
    100970, 100950, 100950, 100940, 100930, 100890, 100930, 100980, 100960, 
    101010, 101030, 101080, 101130, 101180, 101240, 101300, 101350, 101370, 
    101460, 101550, 101620, 101670, 101720, 101740, 101780, 101830, 101900, 
    101970, 102030, 102070, 102150, 102230, 102290, 102340, 102400, 102460, 
    102520, 102580, 102650, 102710, 102770, 102820, 102890, 102970, 103040, 
    103090, 103120, 103160, 103180, 103210, 103200, 103160, 103150, 103130, 
    103060, 103040, 103010, 102950, 102900, 102790, 102670, 102580, 102490, 
    102340, 102210, 102120, 102020, 101980, 101950, 101930, 101920, 101920, 
    101900, 101910, 101910, 101920, 101920, 101910, 101920, 101920, 101950, 
    101990, 102020, 102050, 102090, 102130, 102160, 102170, 102190, 102210, 
    102240, 102230, 102230, 102260, 102270, 102260, 102270, 102270, 102300, 
    102330, 102360, 102340, 102380, 102410, 102470, 102520, 102560, 102580, 
    102600, 102630, 102660, 102680, 102710, 102740, 102770, 102820, 102890, 
    102930, 102950, 102990, 103030, 103070, 103080, 103100, 103130, 103170, 
    103190, 103200, 103220, 103220, 103190, 103180, 103130, 103080, 103050, 
    103010, 102940, 102900, 102870, 102830, 102790, 102750, 102730, 102670, 
    102620, 102570, 102520, 102470, 102430, 102390, 102330, 102310, 102300, 
    102270, 102250, 102210, 102180, 102140, 102120, 102120, 102080, 102060, 
    102050, 102070, 102070, 102040, 102020, 102010, 102010, 102010, 102000, 
    101970, 101960, 101950, 101990, 102030, 102030, 102030, 102040, 102050, 
    102080, 102100, 102100, 102130, 102150, 102160, 102180, 102200, 102220, 
    102220, 102180, 102120, 102070, 102010, 101940, 101810, 101690, 101570, 
    101450, 101320, 101240, 101140, 101060, 100970, 100910, 100850, 100770, 
    100660, 100580, 100520, 100500, 100530, 100540, 100550, 100550, 100570, 
    100580, 100600, 100600, 100600, 100610, 100610, 100600, 100580, 100550, 
    100530, 100510, 100480, 100460, 100470, 100450, 100430, 100470, 100530, 
    100610, 100710, 100810, 100900, 101010, 101120, 101240, 101360, 101460, 
    101560, 101660, 101720, 101830, 101910, 101980, 102060, 102080, 102160, 
    102220, 102270, 102310, 102360, 102420, 102470, 102530, 102610, 102680, 
    102740, 102800, 102850, 102910, 102960, 103010, 103050, 103100, 103130, 
    103150, 103200, 103200, 103220, 103220, 103200, 103170, 103150, 103110, 
    103020, 102950, 102850, 102740, 102600, 102460, 102350, 102250, 102100, 
    101950, 101840, 101760, 101670, 101660, 101720, 101820, 101940, 101980, 
    102060, 102160, 102180, 102300, 102350, 102430, 102510, 102520, 102580, 
    102660, 102730, 102800, 102850, 102870, 102900, 102920, 102940, 102990, 
    103000, 103020, 103040, 103050, 103030, 103040, 103040, 103030, 103010, 
    102980, 102960, 102920, 102890, 102860, 102830, 102800, 102770, 102740, 
    102700, 102610, 102500, 102380, 102290, 102160, 102040, 101850, 101730, 
    101610, 101500, 101410, 101290, 101190, 101090, 101000, 100990, 100940, 
    100910, 100840, 100800, 100740, 100740, 100740, 100670, 100670, 100610, 
    100500, 100420, 100390, 100380, 100400, 100460, 100470, 100530, 100610, 
    100610, 100600, 100690, 100870, 100980, 101090, 101210, 101320, 101440, 
    101550, 101650, 101790, 101930, 102030, 102120, 102200, 102270, 102330, 
    102380, 102430, 102420, 102460, 102500, 102480, 102490, 102450, 102410, 
    102340, 102270, 102210, 102140, 102050, 101980, 101910, 101850, 101790, 
    101710, 101660, 101560, 101490, 101420, 101330, 101270, 101200, 101090, 
    101020, 100960, 100890, 100790, 100730, 100660, 100630, 100580, 100540, 
    100490, 100450, 100380, 100340, 100290, 100240, 100160, 100110, 100020, 
    99950, 99890, 99870, 99850, 99840, 99840, 99850, 99870, 99900, 99890, 
    99900, 99900, 99890, 99900, 99890, 99890, 99860, 99860, 99870, 99870, 
    99860, 99850, 99810, 99760, 99700, 99660, 99550, 99520, 99510, 99470, 
    99390, 99300, 99280, 99260, 99240, 99180, 99120, 99080, 99050, 99020, 
    98970, 98930, 98880, 98840, 98840, 98810, 98770, 98710, 98670, 98660, 
    98660, 98670, 98680, 98690, 98710, 98740, 98790, 98840, 98860, 98870, 
    98900, 98950, 99000, 99060, 99120, 99150, 99190, 99260, 99340, 99400, 
    99460, 99510, 99580, 99660, 99750, 99840, 99910, 100000, 100050, 100110, 
    100170, 100230, 100290, 100340, 100360, 100420, 100450, 100460, 100470, 
    100490, 100520, 100520, 100540, 100530, 100520, 100510, 100440, 100410, 
    100320, 100190, 100090, 100040, 100000, 99970, 99950, 99910, 99890, 
    99880, 99930, 99970, 100020, 100040, 100050, 100060, 100150, 100190, 
    100290, 100360, 100430, 100460, 100490, 100540, 100530, 100570, 100600, 
    100610, 100650, 100660, 100700, 100720, 100710, 100700, 100690, 100610, 
    100520, 100430, 100380, 100350, 100310, 100300, 100320, 100320, 100310, 
    100300, 100230, 100180, 100130, 100110, 100110, 100110, 100090, 100080, 
    100060, 100070, 100060, 100020, 99960, 99950, 99870, 99810, 99780, 99740, 
    99710, 99670, 99630, 99620, 99560, 99530, 99560, 99510, 99490, 99500, 
    99490, 99460, 99430, 99360, 99450, 99400, 99400, 99440, 99460, 99470, 
    99460, 99490, 99530, 99530, 99570, 99590, 99620, 99600, 99570, 99550, 
    99570, 99560, 99560, 99520, 99540, 99530, 99530, 99520, 99550, 99550, 
    99540, 99530, 99500, 99490, 99470, 99420, 99440, 99460, 99480, 99500, 
    99490, 99520, 99500, 99490, 99470, 99440, 99390, 99360, 99310, 99260, 
    99250, 99220, 99210, 99160, 99140, 99100, 99070, 99050, 99040, 99030, 
    99010, 99030, 99060, 99070, 99120, 99190, 99230, 99260, 99320, 99360, 
    99410, 99460, 99520, 99550, 99610, 99660, 99710, 99780, 99860, 99920, 
    99990, 100050, 100120, 100180, 100250, 100310, 100370, 100450, 100530, 
    100600, 100670, 100710, 100760, 100810, 100860, 100930, 100980, 101020, 
    101080, 101140, 101200, 101260, 101300, 101330, 101380, 101430, 101480, 
    101500, 101520, 101540, 101570, 101580, 101580, 101610, 101620, 101620, 
    101600, 101590, 101530, 101490, 101430, 101360, 101290, 101200, 101070, 
    100950, 100840, 100720, 100590, 100430, 100210, 100030, 99820, 99720, 
    99660, 99610, 99570, 99530, 99500, 99480, 99480, 99420, 99370, 99320, 
    99270, 99210, 99180, 99140, 99120, 99090, 99110, 99130, 99180, 99210, 
    99250, 99280, 99290, 99330, 99350, 99360, 99380, 99380, 99360, 99340, 
    99330, 99400, 99440, 99550, 99630, 99670, 99710, 99790, 99840, 99900, 
    99910, 99930, 99930, 99970, 100000, 100010, 100050, 100070, 100130, 
    100170, 100210, 100290, 100330, 100390, 100460, 100520, 100590, 100680, 
    100760, 100810, 100880, 100980, 101010, 101080, 101180, 101200, 101260, 
    101300, 101320, 101330, 101400, 101440, 101480, 101510, 101540, 101550, 
    101540, 101540, 101530, 101460, 101430, 101400, 101350, 101280, 101260, 
    101220, 101200, 101220, 101210, 101190, 101130, 101190, 101200, 101190, 
    101170, 101180, 101120, 101070, 101010, 100910, 100810, 100710, 100590, 
    100490, 100430, 100310, 100250, 100210, 100090, 99990, 99870, 99750, 
    99590, 99400, 99330, 99310, 99310, 99320, 99300, 99300, 99370, 99400, 
    99490, 99570, 99640, 99720, 99750, 99810, 99850, 99880, 99950, 100020, 
    100070, 100160, 100280, 100380, 100490, 100570, 100690, 100770, 100890, 
    100990, 101060, 101140, 101220, 101300, 101370, 101430, 101480, 101530, 
    101580, 101600, 101620, 101650, 101680, 101680, 101720, 101740, 101770, 
    101790, 101800, 101820, 101830, 101850, 101860, 101900, 101910, 101910, 
    101920, 101940, 101960, 101990, 102030, 102040, 102080, 102080, 102110, 
    102130, 102120, 102100, 102120, 102140, 102150, 102160, 102200, 102210, 
    102230, 102210, 102220, 102220, 102220, 102250, 102240, 102280, 102330, 
    102350, 102370, 102380, 102410, 102420, 102430, 102420, 102430, 102430, 
    102400, 102390, 102380, 102350, 102340, 102320, 102310, 102280, 102250, 
    102200, 102170, 102120, 102080, 102060, 102040, 102010, 101970, 101930, 
    101880, 101830, 101740, 101680, 101630, 101560, 101460, 101370, 101290, 
    101190, 101090, 100940, 100880, 100770, 100690, 100580, 100500, 100420, 
    100370, 100310, 100290, 100290, 100300, 100310, 100310, 100310, 100310, 
    100310, 100300, 100310, 100330, 100350, 100360, 100360, 100360, 100360, 
    100340, 100320, 100300, 100260, 100230, 100230, 100230, 100220, 100230, 
    100210, 100230, 100220, 100180, 100140, 100110, 100120, 100110, 100110, 
    100100, 100070, 100060, 99990, 99980, 100020, 100040, 100140, 100200, 
    100300, 100360, 100410, 100460, 100510, 100580, 100630, 100670, 100750, 
    100770, 100820, 100900, 100950, 101020, 101080, 101130, 101190, 101270, 
    101350, 101420, 101450, 101460, 101500, 101510, 101540, 101560, 101580, 
    101580, 101610, 101640, 101660, 101650, 101640, 101610, 101600, 101580, 
    101570, 101520, 101460, 101400, 101360, 101330, 101260, 101180, 101110, 
    101040, 100950, 100840, 100750, 100670, 100560, 100450, 100330, 100260, 
    100130, 99990, 99930, 99820, 99700, 99620, 99560, 99520, 99490, 99480, 
    99500, 99540, 99580, 99620, 99680, 99730, 99800, 99860, 99940, 100070, 
    100190, 100280, 100370, 100490, 100610, 100710, 100800, 100900, 101050, 
    101140, 101170, 101230, 101300, 101360, 101410, 101480, 101520, 101510, 
    101520, 101540, 101550, 101570, 101530, 101530, 101510, 101500, 101500, 
    101490, 101490, 101470, 101450, 101430, 101420, 101420, 101400, 101410, 
    101470, 101490, 101540, 101570, 101590, 101610, 101630, 101700, 101730, 
    101770, 101740, 101750, 101760, 101780, 101850, 101910, 101990, 102040, 
    102090, 102130, 102130, 102150, 102140, 102160, 102170, 102210, 102210, 
    102220, 102230, 102230, 102240, 102210, 102180, 102170, 102180, 102160, 
    102110, 102090, 102060, 102000, 101950, 101930, 101880, 101800, 101780, 
    101710, 101630, 101580, 101530, 101460, 101410, 101380, 101340, 101320, 
    101300, 101270, 101240, 101210, 101200, 101200, 101200, 101190, 101190, 
    101180, 101150, 101120, 101120, 101090, 101050, 101040, 101040, 101030, 
    101010, 100990, 100980, 100950, 100910, 100910, 100910, 100890, 100890, 
    100920, 100930, 100920, 100900, 100890, 100890, 100890, 100880, 100880, 
    100870, 100860, 100870, 100890, 100870, 100850, 100830, 100820, 100810, 
    100800, 100800, 100780, 100770, 100760, 100770, 100740, 100720, 100700, 
    100690, 100700, 100710, 100700, 100710, 100720, 100720, 100720, 100690, 
    100670, 100660, 100650, 100640, 100630, 100650, 100640, 100640, 100640, 
    100620, 100610, 100620, 100620, 100610, 100600, 100610, 100610, 100610, 
    100610, 100630, 100630, 100640, 100630, 100630, 100630, 100630, 100620, 
    100600, 100590, 100600, 100590, 100600, 100590, 100590, 100590, 100580, 
    100580, 100580, 100580, 100580, 100580, 100610, 100640, 100650, 100660, 
    100650, 100630, 100650, 100640, 100610, 100630, 100620, 100610, 100600, 
    100580, 100560, 100540, 100530, 100510, 100490, 100460, 100420, 100380, 
    100350, 100340, 100330, 100320, 100310, 100290, 100250, 100230, 100220, 
    100200, 100190, 100170, 100170, 100170, 100180, 100190, 100180, 100180, 
    100180, 100180, 100180, 100210, 100200, 100160, 100100, 100080, 100090, 
    100090, 100100, 100110, 100120, 100120, 100140, 100170, 100180, 100180, 
    100180, 100210, 100240, 100280, 100310, 100340, 100340, 100330, 100340, 
    100350, 100350, 100330, 100320, 100340, 100360, 100390, 100420, 100450, 
    100480, 100470, 100510, 100490, 100480, 100480, 100470, 100460, 100460, 
    100460, 100460, 100450, 100450, 100470, 100480, 100470, 100450, 100460, 
    100450, 100440, 100420, 100420, 100370, 100350, 100340, 100320, 100290, 
    100280, 100270, 100260, 100250, 100220, 100230, 100230, 100230, 100210, 
    100180, 100200, 100220, 100220, 100180, 100180, 100190, 100200, 100230, 
    100250, 100250, 100270, 100280, 100280, 100300, 100310, 100310, 100290, 
    100310, 100300, 100310, 100330, 100350, 100340, 100330, 100320, 100320, 
    100310, 100290, 100280, 100290, 100280, 100280, 100260, 100250, 100250, 
    100230, 100220, 100220, 100220, 100230, 100220, 100230, 100240, 100230, 
    100260, 100320, 100360, 100390, 100420, 100460, 100510, 100550, 100590, 
    100630, 100680, 100730, 100780, 100830, 100860, 100890, 100930, 100950, 
    101000, 101060, 101110, 101170, 101200, 101260, 101300, 101350, 101370, 
    101410, 101440, 101460, 101510, 101540, 101560, 101580, 101590, 101630, 
    101630, 101640, 101630, 101630, 101600, 101580, 101600, 101590, 101600, 
    101590, 101570, 101560, 101560, 101540, 101530, 101510, 101500, 101480, 
    101450, 101430, 101410, 101390, 101400, 101400, 101400, 101400, 101410, 
    101410, 101420, 101420, 101430, 101420, 101400, 101380, 101360, 101350, 
    101350, 101350, 101360, 101380, 101380, 101350, 101330, 101300, 101300, 
    101300, 101250, 101250, 101260, 101240, 101260, 101260, 101240, 101230, 
    101230, 101210, 101210, 101200, 101190, 101180, 101180, 101170, 101160, 
    101160, 101130, 101110, 101080, 101040, 101010, 101000, 101010, 101000, 
    100990, 100970, 100940, 100920, 100930, 100940, 100980, 101030, 101080, 
    101110, 101150, 101190, 101250, 101300, 101340, 101390, 101470, 101540, 
    101590, 101620, 101640, 101640, 101660, 101660, 101640, 101660, 101590, 
    101530, 101440, 101350, 101210, 101130, 101090, 101130, 101160, 101170, 
    101270, 101350, 101440, 101500, 101600, 101680, 101750, 101820, 101880, 
    101920, 101960, 102000, 102020, 102060, 102060, 102070, 102070, 102050, 
    102070, 102060, 102060, 102050, 102070, 102080, 102120, 102140, 102160, 
    102170, 102220, 102290, 102340, 102360, 102360, 102380, 102430, 102460, 
    102530, 102580, 102600, 102630, 102640, 102650, 102640, 102640, 102630, 
    102640, 102640, 102610, 102610, 102570, 102520, 102470, 102410, 102340, 
    102310, 102280, 102260, 102250, 102230, 102200, 102230, 102240, 102240, 
    102230, 102190, 102160, 102140, 102100, 102050, 102010, 101970, 101900, 
    101850, 101790, 101750, 101660, 101570, 101510, 101420, 101340, 101270, 
    101210, 101170, 101130, 101090, 101040, 100990, 100950, 100910, 100870, 
    100840, 100810, 100800, 100790, 100790, 100820, 100850, 100890, 100920, 
    100940, 100940, 100940, 100950, 100950, 100960, 101010, 101060, 101140, 
    101260, 101360, 101500, 101570, 101650, 101710, 101780, 101840, 101860, 
    101910, 101960, 102030, 102080, 102110, 102140, 102120, 102130, 102160, 
    102180, 102200, 102210, 102210, 102200, 102210, 102240, 102260, 102270, 
    102250, 102220, 102160, 102070, 102000, 101980, 101990, 101990, 101970, 
    101940, 101920, 101880, 101820, 101780, 101750, 101750, 101720, 101690, 
    101670, 101670, 101660, 101660, 101660, 101620, 101600, 101610, 101590, 
    101590, 101610, 101630, 101650, 101680, 101750, 101780, 101840, 101890, 
    101930, 101970, 101980, 101980, 102030, 102070, 102120, 102170, 102230, 
    102280, 102330, 102370, 102380, 102400, 102430, 102430, 102440, 102430, 
    102410, 102400, 102380, 102350, 102330, 102310, 102250, 102260, 102240, 
    102220, 102240, 102240, 102270, 102280, 102300, 102330, 102340, 102330, 
    102330, 102340, 102340, 102280, 102260, 102210, 102200, 102190, 102160, 
    102130, 102080, 102050, 101980, 101900, 101870, 101820, 101750, 101670, 
    101580, 101500, 101460, 101390, 101330, 101260, 101210, 101200, 101190, 
    101230, 101280, 101360, 101440, 101520, 101600, 101700, 101780, 101860, 
    101940, 101970, 102020, 102080, 102130, 102170, 102240, 102300, 102360, 
    102410, 102460, 102510, 102540, 102580, 102620, 102660, 102680, 102670, 
    102710, 102720, 102720, 102700, 102710, 102650, 102560, 102490, 102450, 
    102440, 102380, 102300, 102190, 102100, 102020, 101930, 101890, 101850, 
    101830, 101850, 101820, 101820, 101830, 101850, 101870, 101890, 101910, 
    101930, 101980, 102000, 102010, 102060, 102100, 102120, 102140, 102140, 
    102160, 102170, 102170, 102170, 102180, 102180, 102180, 102150, 102100, 
    102100, 102070, 102020, 101960, 101930, 101920, 101910, 101870, 101850, 
    101820, 101810, 101810, 101790, 101810, 101820, 101830, 101850, 101900, 
    101950, 101990, 102030, 102050, 102080, 102090, 102080, 102080, 102070, 
    102050, 102030, 102010, 101960, 101920, 101860, 101810, 101730, 101640, 
    101550, 101450, 101330, 101230, 101120, 101000, 100940, 100910, 100830, 
    100750, 100680, 100660, 100640, 100650, 100660, 100640, 100650, 100670, 
    100710, 100800, 100870, 100930, 100980, 101020, 101080, 101170, 101260, 
    101350, 101440, 101540, 101640, 101720, 101810, 101890, 101970, 102060, 
    102110, 102160, 102210, 102220, 102260, 102280, 102280, 102280, 102270, 
    102250, 102220, 102140, 102080, 102010, 101950, 101910, 101880, 101830, 
    101830, 101870, 101850, 101850, 101830, 101810, 101830, 101840, 101860, 
    101880, 101930, 101970, 102000, 102030, 102030, 102050, 102030, 102030, 
    102040, 102060, 102040, 102030, 102040, 102060, 102090, 102130, 102130, 
    102130, 102140, 102150, 102170, 102160, 102130, 102100, 102070, 102090, 
    102090, 102040, 102020, 102030, 102000, 101970, 101950, 101920, 101900, 
    101880, 101880, 101850, 101850, 101830, 101810, 101790, 101810, 101780, 
    101760, 101760, 101730, 101680, 101640, 101610, 101600, 101590, 101570, 
    101550, 101520, 101510, 101500, 101490, 101490, 101490, 101480, 101490, 
    101530, 101560, 101560, 101590, 101590, 101590, 101590, 101600, 101610, 
    101620, 101630, 101650, 101670, 101680, 101710, 101720, 101710, 101720, 
    101730, 101730, 101710, 101690, 101690, 101690, 101710, 101750, 101750, 
    101790, 101810, 101850, 101870, 101890, 101900, 101930, 101950, 101950, 
    101980, 101980, 101970, 101970, 101950, 101930, 101900, 101900, 101880, 
    101880, 101890, 101920, 101940, 101970, 101980, 101980, 101970, 101970, 
    101980, 101980, 101990, 101970, 101950, 101920, 101870, 101840, 101820, 
    101830, 101840, 101800, 101880, 101910, 102050, 102160, 102140, 102200, 
    102250, 102330, 102330, 102350, 102430, 102520, 102590, 102620, 102660, 
    102740, 102820, 102840, 102880, 102940, 102920, 102950, 102930, 102970, 
    102960, 102920, 102880, 102850, 102860, 102870, 102910, 102910, 102900, 
    102870, 102840, 102800, 102790, 102760, 102740, 102720, 102710, 102680, 
    102670, 102650, 102620, 102580, 102540, 102510, 102480, 102460, 102440, 
    102420, 102440, 102460, 102470, 102480, 102510, 102540, 102560, 102580, 
    102600, 102640, 102670, 102710, 102750, 102790, 102820, 102860, 102910, 
    102950, 102960, 102990, 103020, 103040, 103050, 103050, 103090, 103090, 
    103110, 103130, 103110, 103090, 103060, 103030, 102970, 102940, 102860, 
    102810, 102770, 102730, 102700, 102650, 102630, 102630, 102590, 102580, 
    102560, 102520, 102480, 102480, 102410, 102390, 102400, 102370, 102330, 
    102360, 102330, 102320, 102270, 102250, 102240, 102300, 102300, 102310, 
    102280, 102260, 102230, 102220, 102200, 102180, 102150, 102110, 102100, 
    102070, 102090, 102110, 102110, 102100, 102130, 102190, 102250, 102300, 
    102360, 102380, 102400, 102400, 102420, 102460, 102490, 102510, 102520, 
    102530, 102540, 102560, 102570, 102580, 102580, 102590, 102750, 102750, 
    102750, 102610, 102620, 102620, 102610, 102580, 102550, 102530, 102520, 
    102490, 102430, 102410, 102370, 102360, 102330, 102250, 102240, 102260, 
    102290, 102250, 102240, 102230, 102220, 102230, 102230, 102270, 102270, 
    102290, 102250, 102240, 102230, 102230, 102190, 102190, 102150, 102110, 
    102110, 102080, 102040, 101990, 101950, 101910, 101860, 101820, 101750, 
    101690, 101630, 101600, 101540, 101490, 101460, 101410, 101350, 101300, 
    101260, 101230, 101170, 101140, 101080, 101060, 101040, 101010, 100970, 
    100930, 100890, 100860, 100820, 100770, 100720, 100680, 100630, 100610, 
    100580, 100530, 100480, 100450, 100410, 100380, 100350, 100340, 100350, 
    100360, 100390, 100400, 100390, 100380, 100420, 100500, 100540, 100560, 
    100570, 100600, 100600, 100630, 100690, 100760, 100810, 100870, 100910, 
    100940, 100950, 100960, 100960, 100970, 100980, 101010, 101030, 101080, 
    101110, 101130, 101130, 101120, 101120, 101120, 101150, 101210, 101250, 
    101280, 101330, 101360, 101420, 101470, 101530, 101600, 101660, 101740, 
    101790, 101860, 101910, 101980, 102110, 102220, 102320, 102430, 102480, 
    102550, 102620, 102680, 102720, 102770, 102830, 102890, 102950, 103020, 
    103070, 103100, 103120, 103160, 103200, 103230, 103270, 103280, 103310, 
    103340, 103390, 103450, 103540, 103590, 103660, 103720, 103770, 103820, 
    103900, 103940, 104040, 104120, 104200, 104270, 104330, 104420, 104440, 
    104500, 104590, 104630, 104650, 104680, 104710, 104740, 104750, 104780, 
    104820, 104890, 104920, 104990, 105100, 105120, 105150, 105200, 105230, 
    105260, 105280, 105300, 105310, 105300, 105290, 105270, 105280, 105300, 
    105320, 105310, 105320, 105330, 105370, 105430, 105460, 105480, 105500, 
    105520, 105520, 105560, 105570, 105590, 105590, 105590, 105610, 105640, 
    105690, 105720, 105730, 105730, 105740, 105730, 105740, 105710, 105700, 
    105700, 105690, 105680, 105660, 105660, 105640, 105610, 105780, 105560, 
    105540, 105510, 105460, 105460, 105430, 105410, 105380, 105340, 105300, 
    105260, 105220, 105170, 105110, 105070, 105020, 104950, 104890, 104880, 
    104830, 104800, 104750, 104680, 104750, 104700, 104460, 104390, 104330, 
    104270, 104200, 104150, 104100, 104030, 103980, 103890, 103830, 103780, 
    103760, 103710, 103700, 103630, 103600, 103600, 103580, 103540, 103500, 
    103460, 103450, 103430, 103370, 103380, 103350, 103300, 103320, 103340, 
    103380, 103380, 103400, 103380, 103350, 103330, 103300, 103300, 103280, 
    103250, 103210, 103130, 103100, 103080, 103030, 102990, 102940, 102890, 
    102890, 102860, 102860, 102870, 102880, 102900, 102930, 102950, 102970, 
    102970, 102960, 102980, 103000, 103020, 103030, 103020, 103050, 103070, 
    103090, 103100, 103070, 103060, 103200, 103030, 103020, 103010, 102990, 
    102960, 102960, 102950, 102940, 102930, 102900, 102880, 102850, 102810, 
    102780, 102740, 102710, 102670, 102640, 102630, 102630, 102600, 102580, 
    102520, 102490, 102490, 102440, 102430, 102400, 102360, 102330, 102310, 
    102260, 102240, 102200, 102160, 102110, 102060, 102000, 101950, 101900, 
    101870, 101810, 101750, 101710, 101630, 101560, 101470, 101390, 101310, 
    101210, 101180, 101120, 101120, 101140, 101200, 101150, 101190, 101230, 
    101280, 101280, 101290, 101240, 101330, 101350, 101320, 101300, 101310, 
    101260, 101200, 101200, 101180, 101200, 101220, 101250, 101300, 101350, 
    101390, 101440, 101510, 101560, 101610, 101650, 101690, 101730, 101750, 
    101780, 101800, 101820, 101830, 101840, 101860, 101850, 101850, 101820, 
    101800, 101800, 101790, 101750, 101750, 101750, 101730, 101700, 101690, 
    101680, 101670, 101650, 101620, 101590, 101550, 101540, 101510, 101470, 
    101450, 101430, 101400, 101380, 101360, 101350, 101340, 101310, 101260, 
    101230, 101200, 101160, 101130, 101090, 101070, 101040, 100990, 101000, 
    100970, 100920, 100880, 100850, 100820, 100780, 100750, 100690, 100650, 
    100610, 100590, 100560, 100520, 100480, 100440, 100390, 100360, 100340, 
    100280, 100250, 100250, 100240, 100220, 100200, 100190, 100180, 100180, 
    100180, 100190, 100200, 100180, 100180, 100180, 100180, 100190, 100200, 
    100210, 100210, 100220, 100220, 100210, 100230, 100230, 100260, 100300, 
    100320, 100350, 100380, 100420, 100440, 100460, 100490, 100500, 100540, 
    100590, 100640, 100670, 100720, 100780, 100820, 100860, 101090, 100920, 
    100950, 101010, 101030, 101070, 101120, 101160, 101220, 101250, 101280, 
    101310, 101360, 101370, 101380, 101400, 101420, 101420, 101440, 101470, 
    101500, 101490, 101500, 101580, 101540, 101550, 101540, 101550, 101550, 
    101550, 101580, 101590, 101610, 101650, 101660, 101680, 101690, 101700, 
    101710, 101730, 101770, 101780, 101820, 101850, 101910, 101950, 101960, 
    101990, 102000, 102020, 102040, 102070, 102110, 102140, 102150, 102170, 
    102200, 102200, 102210, 102270, 102280, 102290, 102280, 102270, 102220, 
    102280, 102340, 102340, 102390, 102420, 102450, 102440, 102480, 102520, 
    102540, 102530, 102540, 102540, 102540, 102520, 102570, 102560, 102550, 
    102510, 102480, 102460, 102450, 102460, 102590, 102680, 102750, 102800, 
    102810, 102830, 102830, 102810, 102790, 102760, 102720, 102640, 102610, 
    102570, 102550, 102490, 102440, 102380, 102320, 102230, 102150, 102080, 
    101990, 101900, 101830, 101790, 101740, 101710, 101730, 101710, 101700, 
    101700, 101710, 101720, 101710, 101710, 101740, 101780, 101830, 101860, 
    101880, 101880, 101890, 101880, 101840, 101830, 101790, 101780, 101720, 
    101680, 101670, 101670, 101630, 101580, 101560, 101520, 101510, 101490, 
    101450, 101390, 101340, 101290, 101260, 101240, 101200, 101170, 101140, 
    101110, 101080, 101070, 101050, 101030, 101030, 100990, 101000, 101010, 
    101020, 101050, 101060, 101060, 101070, 101070, 101070, 101080, 101080, 
    101090, 101100, 101110, 101120, 101120, 101110, 101110, 101120, 101110, 
    101090, 101080, 101080, 101090, 101090, 101100, 101120, 101100, 101090, 
    101080, 101050, 101050, 101040, 101060, 101050, 101050, 101040, 101050, 
    101060, 101050, 101050, 101050, 101060, 101070, 101050, 101030, 101040, 
    101060, 101090, 101130, 101160, 101150, 101140, 101170, 101170, 101190, 
    101160, 101200, 101230, 101250, 101280, 101300, 101340, 101390, 101410, 
    101430, 101450, 101490, 101510, 101520, 101530, 101580, 101610, 101650, 
    101660, 101660, 101650, 101650, 101650, 101670, 101680, 101660, 101630, 
    101610, 101620, 101610, 101600, 101580, 101550, 101530, 101510, 101510, 
    101490, 101450, 101450, 101440, 101440, 101440, 101450, 101450, 101450, 
    101440, 101430, 101430, 101410, 101410, 101400, 101390, 101410, 101430, 
    101430, 101410, 101410, 101380, 101350, 101360, 101340, 101330, 101320, 
    101300, 101270, 101270, 101260, 101240, 101220, 101210, 101190, 101180, 
    101160, 101150, 101130, 101110, 101100, 101090, 101080, 101080, 101070, 
    101060, 101050, 101040, 101040, 101010, 101000, 100990, 100990, 100990, 
    100980, 100980, 100960, 100960, 100950, 100940, 100960, 100950, 100940, 
    100940, 100940, 100940, 100950, 100960, 100960, 100970, 100980, 101000, 
    101030, 101040, 101070, 101070, 101090, 101110, 101120, 101140, 101170, 
    101190, 101180, 101180, 101200, 101180, 101170, 101190, 101190, 101200, 
    101170, 101160, 101140, 101120, 101100, 101070, 101010, 100970, 100930, 
    100880, 100840, 100800, 100770, 100720, 100670, 100630, 100590, 100550, 
    100490, 100440, 100410, 100370, 100360, 100340, 100320, 100320, 100300, 
    100310, 100310, 100300, 100300, 100330, 100310, 100350, 100360, 100390, 
    100390, 100420, 100440, 100470, 100490, 100490, 100500, 100480, 100460, 
    100480, 100490, 100490, 100470, 100470, 100480, 100510, 100480, 100490, 
    100470, 100460, 100460, 100470, 100470, 100480, 100470, 100450, 100440, 
    100440, 100440, 100410, 100390, 100380, 100390, 100400, 100420, 100460, 
    100470, 100480, 100510, 100530, 100560, 100580, 100630, 100680, 100700, 
    100740, 100890, 100840, 100880, 100910, 100940, 100990, 101040, 101080, 
    101110, 101160, 101220, 101250, 101290, 101350, 101400, 101440, 101480, 
    101510, 101540, 101590, 101590, 101610, 101650, 101670, 101670, 101700, 
    101740, 101760, 101750, 101760, 101760, 101750, 101740, 101740, 101720, 
    101700, 101690, 101680, 101630, 101580, 101550, 101510, 101480, 101440, 
    101350, 101250, 101160, 101080, 100960, 100810, 100670, 100460, 100300, 
    100150, 100000, 99820, 99720, 99640, 99600, 99590, 99580, 99590, 99610, 
    99650, 99660, 99650, 99620, 99600, 99560, 99520, 99490, 99450, 99400, 
    99350, 99300, 99270, 99230, 99180, 99150, 99140, 99130, 99120, 99120, 
    99120, 99190, 99140, 99160, 99200, 99220, 99240, 99260, 99280, 99270, 
    99280, 99290, 99300, 99330, 99330, 99320, 99320, 99310, 99270, 99250, 
    99200, 99210, 99170, 99140, 99120, 99070, 99060, 99030, 99010, 99000, 
    99020, 99020, 99040, 99060, 99070, 99100, 99140, 99170, 99200, 99240, 
    99280, 99310, 99340, 99360, 99400, 99430, 99460, 99510, 99540, 99570, 
    99590, 99610, 99630, 99660, 99690, 99720, 99730, 99760, 99790, 99840, 
    99870, 99910, 99950, 99970, 100000, 100030, 100050, 100070, 100070, 
    100080, 100100, 100110, 100140, 100150, 100140, 100140, 100130, 100110, 
    100090, 100090, 100090, 100090, 100090, 100120, 100140, 100170, 100190, 
    100220, 100260, 100280, 100320, 100350, 100370, 100390, 100420, 100460, 
    100500, 100550, 100590, 100630, 100680, 100740, 100790, 100840, 100880, 
    100910, 100950, 100970, 101020, 101060, 101100, 101130, 101140, 101170, 
    101190, 101200, 101200, 101180, 101160, 101150, 101130, 101120, 101120, 
    101110, 101080, 101080, 101050, 101060, 101030, 100980, 100950, 100910, 
    100870, 100820, 100770, 100750, 100710, 100650, 100640, 100620, 100590, 
    100570, 100560, 100540, 100540, 100550, 100570, 100560, 100590, 100630, 
    100640, 100680, 100690, 100720, 100720, 100740, 100760, 100770, 100790, 
    100820, 100840, 100860, 100860, 100850, 100860, 100880, 100890, 100880, 
    100870, 100900, 100930, 100950, 100970, 100990, 101020, 101040, 101050, 
    101040, 101040, 101070, 101090, 101110, 101140, 101170, 101190, 101190, 
    101190, 101190, 101210, 101220, 101220, 101220, 101240, 101240, 101260, 
    101280, 101280, 101280, 101260, 101230, 101230, 101210, 101200, 101180, 
    101160, 101140, 101130, 101110, 101080, 101070, 101050, 101010, 101000, 
    100960, 100950, 100940, 100960, 100960, 100950, 100940, 100920, 100900, 
    100890, 100880, 100860, 100840, 100800, 100770, 100720, 100710, 100680, 
    100640, 100630, 100600, 100560, 100530, 100510, 100460, 100450, 100470, 
    100480, 100470, 100490, 100520, 100530, 100540, 100560, 100580, 100610, 
    100620, 100630, 100650, 100660, 100670, 100710, 100760, 100790, 100830, 
    100860, 100890, 100920, 100940, 100970, 101010, 101020, 101050, 101100, 
    101150, 101160, 101180, 101200, 101210, 101230, 101260, 101260, 101250, 
    101300, 101320, 101330, 101370, 101400, 101420, 101430, 101430, 101420, 
    101410, 101420, 101420, 101430, 101440, 101470, 101470, 101480, 101510, 
    101520, 101560, 101580, 101580, 101580, 101590, 101600, 101610, 101620, 
    101640, 101670, 101640, 101640, 101590, 101570, 101560, 101540, 101520, 
    101490, 101470, 101450, 101430, 101420, 101400, 101370, 101330, 101290, 
    101240, 101190, 101170, 101130, 101100, 101090, 101050, 101010, 100970, 
    100950, 100920, 100900, 100870, 100830, 100770, 100730, 100680, 100660, 
    100610, 100590, 100560, 100560, 100540, 100520, 100510, 100520, 100520, 
    100550, 100580, 100610, 100640, 100660, 100700, 100720, 100750, 100770, 
    100800, 100840, 100870, 100930, 100970, 101020, 101060, 101110, 101160, 
    101190, 101230, 101250, 101270, 101300, 101310, 101360, 101400, 101440, 
    101480, 101530, 101540, 101570, 101600, 101610, 101600, 101620, 101620, 
    101640, 101640, 101640, 101630, 101620, 101620, 101610, 101590, 101560, 
    101550, 101530, 101500, 101490, 101470, 101460, 101450, 101430, 101400, 
    101380, 101340, 101290, 101250, 101150, 101120, 101060, 101020, 100990, 
    100980, 100980, 100970, 100980, 100990, 100970, 100960, 100950, 100950, 
    100950, 100980, 101000, 101020, 101060, 101090, 101110, 101120, 101140, 
    101160, 101190, 101230, 101280, 101300, 101340, 101380, 101430, 101470, 
    101500, 101560, 101600, 101640, 101670, 101710, 101750, 101810, 101870, 
    101910, 101930, 101940, 101990, 102010, 102030, 102040, 102060, 102090, 
    102120, 102150, 102170, 102190, 102210, 102250, 102280, 102310, 102330, 
    102340, 102390, 102410, 102430, 102480, 102530, 102580, 102620, 102660, 
    102680, 102720, 102750, 102790, 102810, 102830, 102850, 102880, 102910, 
    102930, 102960, 102970, 102970, 102980, 102980, 102970, 102960, 102950, 
    102970, 102960, 102970, 102970, 102960, 102930, 102930, 102900, 102860, 
    102840, 102820, 102820, 102800, 102780, 102780, 102770, 102750, 102740, 
    102730, 102710, 102690, 102680, 102640, 102630, 102610, 102600, 102600, 
    102600, 102590, 102550, 102530, 102500, 102480, 102460, 102440, 102430, 
    102450, 102460, 102450, 102430, 102430, 102430, 102440, 102430, 102440, 
    102440, 102440, 102450, 102480, 102520, 102550, 102580, 102590, 102620, 
    102640, 102680, 102720, 102760, 102790, 102830, 102870, 102910, 102950, 
    102970, 103020, 103050, 103070, 103060, 103080, 103090, 103120, 103120, 
    103130, 103120, 103110, 103110, 103130, 103110, 103050, 103050, 103030, 
    102950, 102890, 102860, 102810, 102770, 102730, 102660, 102580, 102540, 
    102430, 102280, 102190, 102070, 101940, 101810, 101720, 101600, 101510, 
    101430, 101350, 101270, 101200, 101150, 101070, 101010, 100980, 100960, 
    100970, 100990, 101000, 101060, 101110, 101170, 101200, 101280, 101340, 
    101390, 101450, 101490, 101540, 101600, 101680, 101750, 101830, 101920, 
    102000, 102070, 102130, 102200, 102260, 102310, 102340, 102360, 102430, 
    102500, 102530, 102570, 102560, 102580, 102600, 102590, 102580, 102580, 
    102560, 102570, 102550, 102530, 102530, 102520, 102500, 102490, 102460, 
    102420, 102390, 102350, 102330, 102330, 102340, 102350, 102350, 102340, 
    102340, 102320, 102300, 102270, 102240, 102220, 102190, 102160, 102150, 
    102150, 102140, 102110, 102080, 102040, 102010, 101990, 101970, 101950, 
    101930, 101940, 101940, 101960, 101960, 101960, 101950, 101940, 101930, 
    101950, 101960, 102000, 102010, 102040, 102110, 102130, 102160, 102160, 
    102180, 102180, 102200, 102210, 102210, 102210, 102230, 102230, 102270, 
    102290, 102310, 102320, 102300, 102310, 102330, 102340, 102350, 102330, 
    102330, 102360, 102390, 102390, 102370, 102350, 102320, 102260, 102230, 
    102160, 102140, 102080, 102050, 102020, 101970, 101920, 101880, 101840, 
    101770, 101690, 101600, 101500, 101410, 101310, 101230, 101150, 101080, 
    101010, 100950, 100900, 100810, 100770, 100680, 100580, 100490, 100420, 
    100350, 100270, 100220, 100200, 100180, 100130, 100100, 100060, 100090, 
    100100, 100120, 100150, 100160, 100230, 100300, 100370, 100440, 100570, 
    100650, 100740, 100830, 100900, 100950, 101030, 101130, 101220, 101320, 
    101410, 101500, 101580, 101650, 101740, 101800, 101870, 101930, 101990, 
    102050, 102110, 102140, 102150, 102180, 102210, 102230, 102210, 102220, 
    102200, 102190, 102170, 102190, 102170, 102170, 102170, 102170, 102150, 
    102150, 102150, 102110, 102090, 102080, 102060, 102040, 102020, 102010, 
    102000, 102000, 101980, 101960, 101920, 101910, 101870, 101840, 101820, 
    101800, 101790, 101780, 101780, 101790, 101810, 101800, 101790, 101760, 
    101740, 101740, 101740, 101740, 101780, 101820, 101860, 101920, 101990, 
    102060, 102090, 102140, 102170, 102200, 102260, 102300, 102340, 102380, 
    102420, 102460, 102510, 102510, 102520, 102530, 102540, 102560, 102540, 
    102530, 102550, 102520, 102470, 102410, 102350, 102230, 102160, 102140, 
    102090, 102040, 102050, 102110, 102140, 102190, 102240, 102280, 102310, 
    102330, 102380, 102400, 102380, 102340, 102320, 102310, 102300, 102300, 
    102290, 102260, 102240, 102190, 102150, 102090, 102060, 102010, 101960, 
    101900, 101860, 101810, 101780, 101760, 101730, 101710, 101650, 101630, 
    101600, 101580, 101550, 101570, 101550, 101550, 101560, 101570, 101580, 
    101610, 101590, 101620, 101630, 101660, 101670, 101700, 101750, 101800, 
    101830, 101880, 101900, 101930, 101960, 101990, 102010, 102040, 102090, 
    102100, 102150, 102190, 102220, 102260, 102270, 102300, 102340, 102370, 
    102380, 102400, 102420, 102460, 102480, 102510, 102540, 102570, 102580, 
    102580, 102570, 102560, 102550, 102550, 102560, 102550, 102540, 102550, 
    102560, 102560, 102560, 102540, 102510, 102510, 102470, 102420, 102380, 
    102340, 102330, 102360, 102360, 102300, 102270, 102240, 102200, 102140, 
    102130, 102080, 102030, 102010, 101970, 101960, 101920, 101850, 101790, 
    101710, 101650, 101620, 101530, 101460, 101440, 101400, 101430, 101430, 
    101440, 101440, 101430, 101390, 101340, 101230, 101150, 101070, 101040, 
    101020, 100990, 101020, 101070, 101130, 101150, 101190, 101190, 101280, 
    101300, 101390, 101450, 101470, 101550, 101590, 101660, 101700, 101720, 
    101720, 101740, 101790, 101840, 101850, 101910, 101940, 101950, 101970, 
    101980, 101970, 101920, 101850, 101770, 101700, 101650, 101590, 101560, 
    101540, 101470, 101430, 101440, 101450, 101410, 101400, 101350, 101310, 
    101290, 101280, 101270, 101270, 101270, 101280, 101310, 101300, 101300, 
    101280, 101280, 101290, 101300, 101310, 101320, 101340, 101400, 101410, 
    101420, 101430, 101410, 101450, 101420, 101410, 101430, 101400, 101370, 
    101330, 101280, 101280, 101210, 101140, 101080, 100990, 100910, 100810, 
    100760, 100730, 100680, 100730, 100770, 100820, 100890, 101020, 101130, 
    101210, 101300, 101360, 101450, 101470, 101500, 101520, 101550, 101580, 
    101610, 101640, 101650, 101660, 101670, 101670, 101670, 101660, 101660, 
    101670, 101660, 101650, 101680, 101660, 101650, 101620, 101580, 101560, 
    101530, 101480, 101430, 101380, 101330, 101300, 101270, 101200, 101140, 
    101090, 101020, 100960, 100890, 100830, 100770, 100760, 100750, 100740, 
    100730, 100730, 100750, 100780, 100790, 100800, 100810, 100830, 100840, 
    100850, 100910, 100950, 101000, 101050, 101090, 101100, 101100, 101130, 
    101140, 101120, 101140, 101150, 101160, 101140, 101160, 101160, 101140, 
    101140, 101150, 101170, 101190, 101210, 101200, 101240, 101260, 101300, 
    101320, 101350, 101370, 101390, 101410, 101420, 101430, 101440, 101430, 
    101430, 101440, 101450, 101460, 101470, 101460, 101450, 101420, 101380, 
    101330, 101280, 101230, 101200, 101180, 101160, 101140, 101100, 101070, 
    101010, 100970, 100910, 100880, 100840, 100800, 100800, 100790, 100790, 
    100800, 100800, 100800, 100780, 100770, 100780, 100810, 100820, 100850, 
    100860, 100880, 100910, 100920, 100930, 100950, 100940, 100930, 100900, 
    100880, 100860, 100830, 100810, 100790, 100780, 100740, 100730, 100660, 
    100620, 100600, 100590, 100550, 100520, 100480, 100410, 100360, 100370, 
    100350, 100320, 100270, 100240, 100230, 100190, 100150, 100100, 100080, 
    100060, 100060, 100090, 100100, 100110, 100130, 100130, 100130, 100140, 
    100140, 100150, 100140, 100120, 100110, 100120, 100110, 100120, 100140, 
    100160, 100190, 100200, 100220, 100220, 100220, 100260, 100290, 100330, 
    100350, 100390, 100420, 100450, 100470, 100490, 100500, 100520, 100540, 
    100530, 100540, 100550, 100570, 100590, 100580, 100590, 100590, 100590, 
    100570, 100570, 100560, 100560, 100550, 100550, 100530, 100530, 100540, 
    100550, 100550, 100530, 100490, 100450, 100410, 100390, 100380, 100390, 
    100380, 100380, 100370, 100360, 100330, 100290, 100250, 100240, 100210, 
    100170, 100160, 100170, 100190, 100210, 100240, 100240, 100270, 100290, 
    100280, 100260, 100280, 100300, 100320, 100340, 100350, 100360, 100390, 
    100420, 100440, 100480, 100500, 100500, 100510, 100530, 100580, 100590, 
    100620, 100610, 100630, 100650, 100680, 100710, 100700, 100740, 100740, 
    100750, 100750, 100760, 100790, 100830, 100870, 100930, 100950, 100980, 
    101000, 101010, 101020, 101030, 101050, 101060, 101080, 101110, 101100, 
    101120, 101110, 101100, 101060, 101070, 101020, 100980, 100970, 100950, 
    100970, 100980, 100970, 100960, 100940, 100930, 100930, 100930, 100920, 
    100930, 100920, 100920, 100930, 100910, 100900, 100860, 100850, 100830, 
    100820, 100800, 100790, 100780, 100780, 100790, 100800, 100780, 100770, 
    100770, 100780, 100800, 100780, 100790, 100810, 100810, 100800, 100820, 
    100840, 100870, 100880, 100890, 100890, 100900, 100930, 100930, 100960, 
    100990, 101040, 101080, 101110, 101130, 101140, 101130, 101120, 101100, 
    101100, 101090, 101060, 101000, 100970, 100970, 100950, 100930, 100880, 
    100840, 100830, 100770, 100720, 100670, 100600, 100530, 100490, 100450, 
    100360, 100320, 100260, 100230, 100170, 100130, 100080, 100040, 100020, 
    100010, 99980, 99990, 99980, 99970, 99960, 99960, 99960, 99960, 99960, 
    100000, 100010, 100030, 100070, 100120, 100180, 100250, 100260, 100290, 
    100370, 100420, 100480, 100520, 100540, 100610, 100720, 100800, 100890, 
    100970, 101050, 101110, 101190, 101250, 101290, 101350, 101400, 101330, 
    101380, 101420, 101540, 101560, 101570, 101590, 101580, 101590, 101590, 
    101590, 101600, 101590, 101580, 101570, 101550, 101550, 101550, 101540, 
    101530, 101500, 101490, 101460, 101420, 101380, 101370, 101360, 101350, 
    101340, 101330, 101310, 101300, 101290, 101280, 101250, 101230, 101230, 
    101230, 101260, 101280, 101260, 101240, 101220, 101210, 101160, 101130, 
    101110, 101130, 101150, 101170, 101200, 101230, 101260, 101280, 101290, 
    101320, 101340, 101320, 101320, 101340, 101340, 101350, 101380, 101410, 
    101440, 101470, 101490, 101520, 101530, 101520, 101510, 101490, 101500, 
    101490, 101480, 101460, 101430, 101390, 101390, 101390, 101380, 101340, 
    101300, 101320, 101310, 101330, 101380, 101440, 101500, 101560, 101590, 
    101600, 101600, 101580, 101560, 101540, 101500, 101500, 101460, 101430, 
    101420, 101370, 101330, 101280, 101200, 101130, 101060, 101000, 100950, 
    100910, 100850, 100810, 100790, 100760, 100760, 100760, 100760, 100750, 
    100780, 100800, 100830, 100900, 100950, 101010, 101030, 101050, 101090, 
    101060, 101030, 101010, 101010, 100940, 100910, 100830, 100780, 100780, 
    100720, 100630, 100620, 100570, 100560, 100530, 100500, 100480, 100480, 
    100560, 100630, 100700, 100720, 100740, 100760, 100730, 100730, 100730, 
    100730, 100710, 100700, 100700, 100720, 100730, 100730, 100710, 100700, 
    100700, 100710, 100700, 100660, 100610, 100590, 100590, 100620, 100690, 
    100740, 100780, 100830, 100850, 100870, 100910, 100930, 100980, 101000, 
    101000, 101040, 101060, 101080, 101080, 101080, 101080, 101080, 101070, 
    101080, 101110, 101100, 101140, 101180, 101220, 101220, 101190, 101180, 
    101190, 101170, 101150, 101140, 101130, 101120, 101100, 101110, 101110, 
    101070, 101020, 101000, 100950, 100940, 100910, 100870, 100820, 100780, 
    100750, 100730, 100730, 100700, 100670, 100650, 100590, 100550, 100540, 
    100500, 100460, 100420, 100390, 100390, 100360, 100340, 100340, 100320, 
    100330, 100340, 100330, 100320, 100320, 100320, 100320, 100320, 100340, 
    100340, 100340, 100330, 100340, 100350, 100360, 100370, 100380, 100410, 
    100450, 100490, 100530, 100560, 100590, 100640, 100650, 100660, 100670, 
    100680, 100700, 100720, 100710, 100690, 100670, 100660, 100650, 100610, 
    100580, 100570, 100550, 100520, 100510, 100510, 100550, 100600, 100630, 
    100670, 100690, 100680, 100650, 100620, 100590, 100580, 100580, 100580, 
    100580, 100590, 100620, 100620, 100610, 100610, 100590, 100550, 100520, 
    100460, 100420, 100380, 100330, 100310, 100290, 100260, 100240, 100200, 
    100180, 100130, 100060, 99990, 99980, 100010, 100060, 100130, 100170, 
    100190, 100220, 100230, 100190, 100170, 100140, 100120, 100100, 100080, 
    100070, 100040, 100030, 100050, 100030, 100000, 99980, 99960, 99960, 
    99940, 99930, 99920, 99900, 99910, 99910, 99910, 99910, 99900, 99890, 
    99900, 99890, 99890, 99880, 99870, 99880, 99900, 99910, 99910, 99900, 
    99880, 99850, 99820, 99790, 99770, 99780, 99760, 99730, 99720, 99720, 
    99720, 99680, 99660, 99650, 99640, 99620, 99610, 99600, 99600, 99600, 
    99610, 99620, 99640, 99670, 99680, 99690, 99700, 99710, 99740, 99750, 
    99780, 99810, 99850, 99910, 99920, 99960, 99990, 100040, 100070, 100110, 
    100140, 100180, 100210, 100260, 100290, 100330, 100380, 100420, 100460, 
    100500, 100540, 100580, 100610, 100620, 100660, 100710, 100770, 100820, 
    100880, 100930, 100980, 101030, 101070, 101120, 101150, 101190, 101230, 
    101280, 101320, 101380, 101420, 101470, 101500, 101530, 101550, 101570, 
    101590, 101610, 101610, 101600, 101630, 101630, 101630, 101620, 101620, 
    101620, 101600, 101590, 101570, 101550, 101540, 101520, 101470, 101440, 
    101410, 101400, 101360, 101320, 101290, 101250, 101200, 101170, 101160, 
    101130, 101100, 101110, 101080, 101040, 101020, 100970, 100960, 100930, 
    100890, 100840, 100800, 100750, 100720, 100700, 100670, 100640, 100620, 
    100610, 100530, 100510, 100480, 100450, 100420, 100390, 100340, 100310, 
    100260, 100240, 100270, 100210, 100170, 100140, 100100, 100090, 100020, 
    100000, 99980, 99940, 99920, 99920, 99880, 99850, 99800, 99780, 99760, 
    99730, 99690, 99710, 99680, 99690, 99710, 99700, 99730, 99770, 99790, 
    99790, 99820, 99830, 99820, 99830, 99860, 99890, 99930, 99970, 100010, 
    100040, 100080, 100110, 100140, 100160, 100230, 100290, 100340, 100370, 
    100430, 100460, 100510, 100550, 100570, 100600, 100630, 100640, 100690, 
    100720, 100780, 100800, 100850, 100890, 100930, 100970, 101000, 101020, 
    101040, 101070, 101080, 101100, 101110, 101150, 101170, 101190, 101200, 
    101210, 101220, 101220, 101220, 101250, 101270, 101300, 101320, 101330, 
    101350, 101370, 101390, 101410, 101420, 101430, 101440, 101480, 101500, 
    101540, 101570, 101600, 101630, 101670, 101700, 101700, 101730, 101730, 
    101720, 101720, 101750, 101770, 101790, 101770, 101800, 101790, 101790, 
    101790, 101790, 101780, 101770, 101740, 101680, 101640, 101610, 101550, 
    101520, 101440, 101360, 101310, 101250, 101150, 101050, 100940, 100900, 
    100770, 100700, 100650, 100610, 100520, 100470, 100420, 100320, 100240, 
    100170, 100120, 100050, 99990, 99960, 99940, 99930, 99930, 99940, 99940, 
    99960, 99980, 99990, 100010, 100020, 100090, 100160, 100270, 100320, 
    100380, 100430, 100500, 100550, 100610, 100670, 100730, 100760, 100760, 
    100800, 100850, 100880, 100900, 100920, 100940, 100970, 100980, 101010, 
    101060, 101100, 101130, 101120, 101130, 101150, 101160, 101160, 101170, 
    101180, 101190, 101200, 101230, 101270, 101310, 101330, 101360, 101390, 
    101430, 101440, 101450, 101470, 101480, 101500, 101510, 101500, 101510, 
    101530, 101560, 101570, 101560, 101580, 101590, 101600, 101580, 101610, 
    101630, 101640, 101650, 101680, 101700, 101710, 101730, 101740, 101750, 
    101730, 101730, 101750, 101760, 101750, 101750, 101720, 101720, 101710, 
    101710, 101730, 101750, 101720, 101690, 101670, 101670, 101670, 101670, 
    101650, 101650, 101640, 101640, 101640, 101630, 101620, 101600, 101570, 
    101560, 101560, 101540, 101520, 101510, 101490, 101490, 101490, 101490, 
    101480, 101480, 101470, 101480, 101470, 101470, 101480, 101480, 101470, 
    101470, 101470, 101460, 101440, 101410, 101370, 101340, 101310, 101280, 
    101250, 101230, 101220, 101210, 101190, 101140, 101100, 101060, 101050, 
    101020, 100970, 100960, 100950, 100940, 100930, 100900, 100900, 100890, 
    100900, 100880, 100870, 100880, 100880, 100900, 100910, 100910, 100910, 
    100940, 100970, 100970, 100990, 100980, 100980, 101000, 101030, 101070, 
    101120, 101160, 101180, 101220, 101260, 101290, 101330, 101350, 101380, 
    101380, 101400, 101440, 101460, 101470, 101470, 101480, 101470, 101460, 
    101440, 101440, 101430, 101430, 101420, 101440, 101430, 101450, 101450, 
    101460, 101450, 101450, 101460, 101460, 101440, 101430, 101450, 101460, 
    101470, 101500, 101510, 101510, 101500, 101490, 101490, 101490, 101480, 
    101490, 101490, 101520, 101520, 101520, 101520, 101520, 101500, 101500, 
    101490, 101450, 101430, 101440, 101440, 101410, 101400, 101410, 101400, 
    101360, 101340, 101320, 101310, 101280, 101260, 101270, 101250, 101230, 
    101220, 101230, 101240, 101250, 101250, 101250, 101210, 101200, 101180, 
    101170, 101140, 101160, 101140, 101150, 101150, 101150, 101160, 101170, 
    101170, 101160, 101130, 101110, 101090, 101090, 101040, 101020, 101030, 
    101010, 100970, 100930, 100880, 100840, 100800, 100760, 100690, 100650, 
    100580, 100550, 100470, 100350, 100250, 100190, 100140, 100110, 100080, 
    100090, 100050, 100050, 100060, 100140, 100170, 100190, 100210, 100270, 
    100320, 100380, 100440, 100490, 100550, 100620, 100680, 100740, 100790, 
    100850, 100890, 100940, 100980, 101030, 101070, 101110, 101160, 101200, 
    101260, 101300, 101370, 101420, 101470, 101500, 101530, 101530, 101560, 
    101570, 101590, 101600, 101610, 101630, 101640, 101650, 101650, 101650, 
    101640, 101640, 101630, 101620, 101630, 101620, 101620, 101660, 101680, 
    101680, 101660, 101650, 101590, 101600, 101590, 101590, 101630, 101630, 
    101610, 101640, 101620, 101620, 101620, 101590, 101570, 101570, 101540, 
    101530, 101520, 101520, 101470, 101450, 101430, 101430, 101440, 101400, 
    101380, 101350, 101350, 101350, 101340, 101360, 101370, 101370, 101370, 
    101370, 101380, 101370, 101380, 101410, 101430, 101440, 101440, 101470, 
    101490, 101500, 101520, 101530, 101530, 101540, 101530, 101510, 101520, 
    101500, 101510, 101520, 101500, 101500, 101510, 101490, 101450, 101420, 
    101390, 101360, 101330, 101320, 101300, 101270, 101240, 101230, 101210, 
    101210, 101150, 101100, 101060, 101020, 100970, 100910, 100840, 100810, 
    100770, 100750, 100680, 100620, 100570, 100550, 100510, 100500, 100490, 
    100470, 100480, 100500, 100520, 100540, 100570, 100580, 100620, 100630, 
    100650, 100690, 100690, 100710, 100730, 100750, 100780, 100800, 100810, 
    100800, 100820, 100800, 100800, 100800, 100800, 100790, 100810, 100800, 
    100800, 100800, 100800, 100800, 100790, 100780, 100780, 100760, 100780, 
    100780, 100790, 100780, 100800, 100810, 100810, 100810, 100800, 100800, 
    100800, 100790, 100770, 100770, 100720, 100680, 100650, 100630, 100600, 
    100570, 100520, 100490, 100430, 100320, 100270, 100180, 100140, 100090, 
    100070, 100060, 100100, 100120, 100120, 100150, 100180, 100210, 100260, 
    100310, 100380, 100420, 100470, 100480, 100520, 100550, 100540, 100540, 
    100510, 100470, 100440, 100400, 100350, 100330, 100300, 100280, 100230, 
    100180, 100140, 100110, 100040, 99970, 99900, 99860, 99810, 99770, 99730, 
    99700, 99690, 99640, 99570, 99500, 99450, 99420, 99410, 99390, 99370, 
    99390, 99400, 99410, 99420, 99440, 99460, 99490, 99510, 99510, 99550, 
    99580, 99630, 99660, 99670, 99680, 99700, 99710, 99720, 99710, 99700, 
    99680, 99660, 99620, 99610, 99620, 99610, 99620, 99630, 99640, 99660, 
    99700, 99740, 99770, 99850, 99930, 100000, 100060, 100140, 100190, 
    100250, 100290, 100360, 100400, 100440, 100470, 100500, 100520, 100540, 
    100540, 100540, 100520, 100440, 100370, 100270, 100170, 100060, 100000, 
    99920, 99840, 99780, 99770, 99750, 99760, 99790, 99850, 99940, 99980, 
    100040, 100100, 100140, 100160, 100190, 100220, 100270, 100300, 100320, 
    100340, 100340, 100330, 100340, 100340, 100340, 100330, 100320, 100310, 
    100300, 100290, 100310, 100300, 100320, 100300, 100280, 100260, 100250, 
    100250, 100280, 100300, 100320, 100330, 100350, 100360, 100380, 100410, 
    100440, 100450, 100480, 100490, 100510, 100540, 100560, 100580, 100610, 
    100620, 100650, 100640, 100640, 100610, 100600, 100620, 100640, 100640, 
    100680, 100660, 100630, 100620, 100580, 100580, 100560, 100530, 100500, 
    100520, 100500, 100540, 100560, 100540, 100570, 100600, 100620, 100590, 
    100570, 100580, 100550, 100510, 100520, 100540, 100490, 100480, 100470, 
    100430, 100410, 100390, 100400, 100390, 100400, 100400, 100380, 100390, 
    100420, 100410, 100400, 100370, 100390, 100410, 100450, 100450, 100410, 
    100380, 100400, 100420, 100420, 100400, 100370, 100330, 100290, 100240, 
    100200, 100210, 100200, 100180, 100170, 100180, 100210, 100210, 100180, 
    100160, 100150, 100100, 100060, 100010, 99990, 99960, 99940, 99910, 
    99890, 99880, 99880, 99860, 99860, 99860, 99860, 99870, 99870, 99880, 
    99870, 99880, 99890, 99920, 99930, 99940, 99980, 99980, 99980, 99990, 
    100000, 100000, 100010, 100010, 100020, 100040, 100070, 100100, 100110, 
    100120, 100140, 100150, 100160, 100170, 100180, 100190, 100220, 100240, 
    100260, 100270, 100300, 100340, 100360, 100370, 100380, 100360, 100390, 
    100430, 100460, 100480, 100510, 100550, 100570, 100590, 100620, 100650, 
    100660, 100670, 100700, 100710, 100730, 100760, 100770, 100780, 100800, 
    100800, 100790, 100780, 100750, 100720, 100680, 100660, 100650, 100610, 
    100570, 100530, 100470, 100390, 100320, 100260, 100200, 100150, 100130, 
    100130, 100140, 100170, 100220, 100320, 100450, 100570, 100680, 100790, 
    100890, 100990, 101060, 101150, 101240, 101330, 101400, 101440, 101490, 
    101550, 101580, 101610, 101650, 101670, 101710, 101730, 101780, 101800, 
    101830, 101850, 101850, 101850, 101850, 101860, 101830, 101830, 101820, 
    101810, 101790, 101770, 101740, 101670, 101620, 101580, 101530, 101450, 
    101380, 101300, 101220, 101170, 101090, 101000, 100930, 100870, 100850, 
    100810, 100720, 100590, 100500, 100440, 100390, 100360, 100310, 100270, 
    100220, 100140, 100040, 99940, 99790, 99670, 99630, 99570, 99480, 99400, 
    99360, 99330, 99270, 99250, 99240, 99220, 99240, 99260, 99260, 99280, 
    99270, 99320, 99350, 99380, 99400, 99430, 99440, 99480, 99500, 99510, 
    99500, 99520, 99530, 99530, 99540, 99530, 99540, 99550, 99560, 99550, 
    99540, 99530, 99530, 99550, 99540, 99530, 99520, 99530, 99510, 99470, 
    99470, 99440, 99420, 99390, 99390, 99360, 99320, 99310, 99280, 99260, 
    99240, 99190, 99190, 99170, 99140, 99110, 99090, 99120, 99110, 99080, 
    99050, 99050, 99030, 99020, 99050, 99070, 99090, 99110, 99130, 99190, 
    99230, 99280, 99320, 99330, 99380, 99470, 99500, 99590, 99640, 99710, 
    99730, 99810, 99900, 99970, 100050, 100110, 100160, 100230, 100290, 
    100360, 100410, 100460, 100500, 100570, 100630, 100680, 100730, 100790, 
    100840, 100900, 100940, 100960, 101010, 101050, 101070, 101100, 101120, 
    101150, 101160, 101200, 101250, 101280, 101310, 101340, 101350, 101390, 
    101390, 101410, 101440, 101460, 101480, 101510, 101540, 101560, 101560, 
    101570, 101570, 101580, 101590, 101590, 101590, 101580, 101610, 101620, 
    101630, 101630, 101620, 101610, 101600, 101590, 101580, 101570, 101570, 
    101560, 101560, 101560, 101570, 101560, 101540, 101530, 101520, 101520, 
    101510, 101500, 101500, 101500, 101500, 101520, 101510, 101500, 101510, 
    101500, 101500, 101500, 101510, 101500, 101480, 101470, 101490, 101490, 
    101490, 101500, 101490, 101450, 101410, 101390, 101370, 101350, 101320, 
    101300, 101300, 101310, 101320, 101320, 101310, 101260, 101220, 101180, 
    101120, 101090, 101030, 100980, 100980, 100950, 100930, 100870, 100830, 
    100800, 100770, 100770, 100760, 100750, 100750, 100730, 100720, 100740, 
    100730, 100720, 100700, 100650, 100610, 100550, 100530, 100510, 100500, 
    100500, 100500, 100460, 100470, 100450, 100410, 100370, 100320, 100260, 
    100230, 100250, 100280, 100280, 100290, 100270, 100260, 100230, 100190, 
    100140, 100130, 100100, 100080, 100070, 100070, 100050, 100020, 99980, 
    100000, 100000, 100010, 100040, 100050, 100060, 100070, 100080, 100090, 
    100080, 100110, 100130, 100150, 100130, 100140, 100160, 100180, 100190, 
    100180, 100160, 100140, 100130, 100110, 100090, 100060, 100040, 100000, 
    99940, 99900, 99860, 99850, 99860, 99880, 99940, 99970, 100010, 100080, 
    100150, 100220, 100250, 100290, 100320, 100330, 100370, 100380, 100370, 
    100340, 100290, 100190, 100100, 100050, 100020, 99930, 99910, 99890, 
    99870, 99920, 99970, 100020, 100090, 100190, 100290, 100370, 100430, 
    100470, 100520, 100570, 100620, 100640, 100690, 100700, 100720, 100730, 
    100700, 100690, 100670, 100620, 100610, 100610, 100600, 100620, 100630, 
    100700, 100750, 100820, 100890, 100920, 101000, 101030, 101120, 101130, 
    101240, 101310, 101360, 101400, 101460, 101490, 101510, 101560, 101570, 
    101570, 101570, 101600, 101570, 101610, 101580, 101540, 101550, 101520, 
    101490, 101480, 101430, 101360, 101310, 101260, 101220, 101180, 101120, 
    101050, 100960, 100910, 100840, 100770, 100680, 100630, 100570, 100510, 
    100460, 100430, 100410, 100390, 100370, 100360, 100370, 100390, 100410, 
    100410, 100400, 100400, 100390, 100380, 100380, 100400, 100400, 100440, 
    100470, 100490, 100480, 100480, 100470, 100460, 100460, 100470, 100450, 
    100480, 100480, 100490, 100530, 100590, 100610, 100640, 100690, 100710, 
    100740, 100770, 100790, 100800, 100800, 100850, 100860, 100860, 100820, 
    100770, 100740, 100700, 100710, 100690, 100670, 100640, 100620, 100600, 
    100570, 100540, 100460, 100370, 100330, 100280, 100250, 100270, 100230, 
    100210, 100210, 100200, 100170, 100160, 100130, 100160, 100150, 100130, 
    100140, 100180, 100220, 100260, 100310, 100360, 100400, 100400, 100390, 
    100390, 100420, 100400, 100390, 100360, 100370, 100380, 100400, 100450, 
    100490, 100540, 100570, 100590, 100600, 100630, 100650, 100680, 100720, 
    100740, 100740, 100760, 100770, 100790, 100810, 100840, 100860, 100910, 
    100940, 100990, 101060, 101130, 101170, 101220, 101280, 101320, 101360, 
    101360, 101400, 101420, 101470, 101500, 101540, 101570, 101580, 101600, 
    101620, 101630, 101620, 101620, 101620, 101620, 101610, 101610, 101630, 
    101620, 101600, 101540, 101510, 101480, 101470, 101440, 101410, 101360, 
    101340, 101320, 101300, 101310, 101320, 101290, 101250, 101210, 101200, 
    101200, 101160, 101160, 101150, 101140, 101140, 101190, 101240, 101250, 
    101220, 101200, 101220, 101240, 101250, 101260, 101290, 101320, 101340, 
    101350, 101360, 101360, 101340, 101360, 101380, 101400, 101390, 101400, 
    101440, 101480, 101500, 101510, 101560, 101610, 101610, 101650, 101650, 
    101670, 101710, 101740, 101750, 101790, 101820, 101820, 101830, 101850, 
    101870, 101890, 101910, 101920, 101930, 101950, 101960, 101980, 102000, 
    102020, 102040, 102050, 102040, 102040, 102040, 102050, 102070, 102070, 
    102090, 102100, 102110, 102110, 102120, 102120, 102140, 102150, 102170, 
    102170, 102170, 102210, 102210, 102220, 102230, 102240, 102260, 102270, 
    102230, 102240, 102230, 102220, 102230, 102250, 102230, 102270, 102270, 
    102280, 102300, 102320, 102340, 102350, 102360, 102360, 102380, 102400, 
    102470, 102490, 102530, 102550, 102530, 102540, 102550, 102550, 102550, 
    102540, 102530, 102570, 102580, 102600, 102600, 102620, 102630, 102640, 
    102670, 102720, 102730, 102750, 102760, 102770, 102800, 102830, 102890, 
    102930, 102960, 102990, 103040, 103070, 103100, 103140, 103170, 103180, 
    103210, 103250, 103290, 103330, 103370, 103400, 103410, 103440, 103450, 
    103460, 103480, 103470, 103460, 103480, 103500, 103500, 103510, 103520, 
    103520, 103520, 103520, 103510, 103510, 103500, 103490, 103490, 103490, 
    103490, 103500, 103490, 103480, 103450, 103420, 103420, 103400, 103390, 
    103380, 103350, 103330, 103320, 103320, 103310, 103320, 103300, 103300, 
    103280, 103270, 103270, 103270, 103270, 103260, 103260, 103270, 103270, 
    103250, 103240, 103230, 103220, 103210, 103190, 103190, 103190, 103200, 
    103170, 103160, 103150, 103140, 103130, 103120, 103130, 103120, 103100, 
    103100, 103100, 103100, 103110, 103110, 103120, 103120, 103120, 103110, 
    103100, 103090, 103100, 103120, 103120, 103110, 103120, 103130, 103120, 
    103100, 103080, 103100, 103090, 103070, 103030, 103000, 103000, 102990, 
    103010, 103040, 103040, 103060, 103080, 103070, 103060, 103030, 103030, 
    103010, 103000, 103000, 102990, 102970, 102960, 102980, 102960, 102940, 
    102920, 102900, 102880, 102860, 102860, 102850, 102850, 102860, 102850, 
    102890, 102860, 102830, 102820, 102790, 102750, 102720, 102730, 102710, 
    102690, 102680, 102660, 102650, 102620, 102580, 102560, 102530, 102500, 
    102480, 102520, 102510, 102490, 102470, 102470, 102420, 102410, 102400, 
    102420, 102390, 102360, 102360, 102360, 102360, 102340, 102350, 102350, 
    102340, 102330, 102310, 102260, 102240, 102200, 102170, 102130, 102080, 
    102030, 101990, 101950, 101890, 101830, 101740, 101620, 101480, 101380, 
    101260, 101110, 101000, 100880, 100760, 100670, 100570, 100440, 100320, 
    100210, 100130, 100050, 100010, 99930, 99870, 99810, 99710, 99630, 99570, 
    99500, 99520, 99540, 99540, 99520, 99520, 99550, 99610, 99660, 99720, 
    99760, 99810, 99830, 99850, 99830, 99780, 99730, 99660, 99630, 99600, 
    99550, 99490, 99410, 99310, 99200, 99090, 99030, 99020, 99040, 99040, 
    99060, 99130, 99200, 99260, 99320, 99350, 99410, 99490, 99550, 99620, 
    99680, 99740, 99810, 99900, 99950, 100000, 100050, 100100, 100160, 
    100180, 100210, 100210, 100260, 100270, 100270, 100320, 100350, 100380, 
    100440, 100470, 100510, 100540, 100560, 100560, 100620, 100630, 100640, 
    100660, 100690, 100720, 100760, 100770, 100810, 100810, 100820, 100830, 
    100830, 100840, 100840, 100860, 100900, 100890, 100910, 100910, 100910, 
    100890, 100920, 100960, 100950, 100990, 101030, 101090, 101080, 101100, 
    101110, 101130, 101130, 101170, 101160, 101160, 101150, 101170, 101150, 
    101160, 101180, 101140, 101130, 101130, 101100, 101090, 101070, 101070, 
    101040, 101040, 101040, 101030, 101050, 101080, 101100, 101120, 101160, 
    101180, 101210, 101190, 101230, 101210, 101260, 101260, 101260, 101290, 
    101340, 101350, 101380, 101370, 101420, 101430, 101460, 101490, 101520, 
    101550, 101570, 101610, 101640, 101640, 101660, 101650, 101650, 101650, 
    101650, 101650, 101650, 101660, 101650, 101640, 101640, 101620, 101620, 
    101600, 101570, 101540, 101530, 101540, 101540, 101550, 101540, 101550, 
    101540, 101540, 101520, 101490, 101450, 101430, 101400, 101360, 101330, 
    101300, 101260, 101220, 101190, 101150, 101130, 101080, 101020, 100970, 
    100940, 100900, 100860, 100820, 100810, 100790, 100760, 100730, 100680, 
    100630, 100580, 100540, 100520, 100500, 100450, 100430, 100400, 100340, 
    100300, 100250, 100210, 100150, 100100, 100050, 99990, 99930, 99870, 
    99810, 99760, 99710, 99620, 99550, 99520, 99490, 99460, 99430, 99420, 
    99430, 99440, 99460, 99460, 99490, 99510, 99520, 99580, 99610, 99620, 
    99680, 99740, 99820, 99910, 100020, 100110, 100250, 100360, 100490, 
    100610, 100700, 100790, 100880, 100970, 101030, 101110, 101150, 101200, 
    101250, 101290, 101320, 101270, 101310, 101280, 101240, 101230, 101210, 
    101210, 101170, 101150, 101150, 101180, 101200, 101190, 101210, 101260, 
    101330, 101400, 101520, 101640, 101740, 101910, 102040, 102150, 102210, 
    102310, 102380, 102430, 102430, 102470, 102470, 102440, 102400, 102400, 
    102410, 102360, 102320, 102250, 102180, 102120, 102060, 101990, 101930, 
    101890, 101850, 101830, 101780, 101730, 101670, 101610, 101560, 101500, 
    101430, 101380, 101330, 101250, 101210, 101160, 101110, 101110, 101110, 
    101110, 101090, 101090, 101080, 101090, 101140, 101210, 101270, 101380, 
    101490, 101530, 101580, 101630, 101680, 101730, 101770, 101830, 101840, 
    101880, 101940, 101990, 102040, 102070, 102090, 102090, 102110, 102110, 
    102130, 102120, 102110, 102090, 102100, 102100, 102090, 102040, 102010, 
    101980, 101960, 101930, 101890, 101850, 101800, 101780, 101730, 101720, 
    101680, 101620, 101560, 101490, 101450, 101370, 101310, 101250, 101180, 
    101140, 101100, 101060, 101030, 101000, 100950, 100920, 100890, 100860, 
    100800, 100790, 100760, 100770, 100760, 100760, 100770, 100800, 100790, 
    100780, 100770, 100780, 100810, 100850, 100860, 100870, 100900, 100950, 
    100960, 100980, 101030, 101050, 101060, 101090, 101120, 101160, 101180, 
    101210, 101260, 101270, 101310, 101360, 101410, 101430, 101480, 101520, 
    101550, 101580, 101580, 101620, 101650, 101680, 101720, 101730, 101740, 
    101750, 101760, 101770, 101790, 101800, 101810, 101810, 101810, 101840, 
    101850, 101870, 101890, 101890, 101890, 101880, 101900, 101910, 101930, 
    101930, 101960, 101980, 101990, 101980, 101980, 101960, 101960, 101950, 
    101930, 101900, 101880, 101850, 101830, 101810, 101800, 101770, 101740, 
    101710, 101660, 101620, 101580, 101560, 101510, 101460, 101420, 101380, 
    101330, 101280, 101240, 101200, 101160, 101120, 101090, 101060, 101040, 
    101020, 101020, 101020, 101000, 100940, 100920, 100900, 100890, 100850, 
    100790, 100750, 100700, 100690, 100670, 100670, 100650, 100630, 100640, 
    100610, 100580, 100570, 100570, 100560, 100540, 100530, 100530, 100530, 
    100530, 100540, 100520, 100480, 100460, 100440, 100390, 100380, 100370, 
    100340, 100340, 100310, 100290, 100280, 100270, 100240, 100240, 100240, 
    100230, 100210, 100210, 100220, 100240, 100270, 100290, 100300, 100300, 
    100310, 100310, 100330, 100350, 100360, 100360, 100370, 100380, 100380, 
    100400, 100410, 100400, 100400, 100400, 100390, 100380, 100370, 100370, 
    100380, 100400, 100420, 100460, 100470, 100460, 100480, 100480, 100460, 
    100460, 100430, 100430, 100430, 100420, 100410, 100400, 100380, 100310, 
    100270, 100250, 100200, 100150, 100140, 100140, 100140, 100150, 100150, 
    100160, 100170, 100180, 100190, 100200, 100220, 100320, 100280, 100300, 
    100310, 100330, 100320, 100340, 100360, 100370, 100370, 100380, 100370, 
    100370, 100360, 100360, 100350, 100350, 100360, 100370, 100380, 100360, 
    100360, 100340, 100330, 100330, 100330, 100330, 100320, 100310, 100310, 
    100290, 100290, 100290, 100260, 100250, 100220, 100210, 100190, 100180, 
    100170, 100170, 100170, 100180, 100180, 100180, 100180, 100180, 100180, 
    100170, 100140, 100150, 100160, 100150, 100140, 100130, 100130, 100110, 
    100110, 100090, 100090, 100080, 100060, 100050, 100050, 100080, 100090, 
    100110, 100110, 100110, 100140, 100150, 100140, 100150, 100160, 100170, 
    100190, 100210, 100230, 100250, 100250, 100270, 100280, 100300, 100310, 
    100330, 100360, 100370, 100400, 100440, 100450, 100480, 100500, 100510, 
    100560, 100560, 100550, 100540, 100570, 100560, 100590, 100590, 100580, 
    100580, 100590, 100590, 100550, 100520, 100510, 100470, 100440, 100420, 
    100420, 100430, 100410, 100430, 100420, 100420, 100420, 100410, 100430, 
    100460, 100480, 100530, 100580, 100620, 100650, 100690, 100740, 100790, 
    100810, 100840, 100870, 100860, 100860, 100880, 100900, 100930, 100950, 
    100960, 101000, 101030, 101030, 101020, 101010, 101000, 101000, 100990, 
    100970, 100980, 100990, 100980, 100970, 100980, 100980, 100980, 100960, 
    100930, 100900, 100880, 100880, 100870, 100880, 100900, 100900, 100900, 
    100890, 100850, 100830, 100830, 100790, 100770, 100750, 100730, 100720, 
    100730, 100710, 100710, 100690, 100650, 100610, 100550, 100490, 100440, 
    100390, 100350, 100320, 100290, 100250, 100230, 100200, 100160, 100110, 
    100020, 99930, 99900, 99860, 99790, 99740, 99700, 99660, 99600, 99550, 
    99510, 99470, 99450, 99430, 99390, 99340, 99300, 99270, 99240, 99230, 
    99190, 99170, 99170, 99180, 99160, 99170, 99200, 99230, 99270, 99300, 
    99330, 99370, 99400, 99400, 99410, 99460, 99480, 99500, 99530, 99550, 
    99570, 99600, 99590, 99570, 99560, 99550, 99510, 99460, 99420, 99360, 
    99280, 99160, 99090, 98990, 98880, 98850, 98730, 98550, 98410, 98280, 
    98200, 98130, 98060, 97990, 97920, 97890, 97900, 97890, 97890, 97870, 
    97840, 97820, 97790, 97770, 97710, 97700, 97680, 97710, 97730, 97770, 
    97800, 97780, 97810, 97800, 97790, 97800, 97840, 97860, 97910, 98000, 
    98080, 98170, 98210, 98250, 98280, 98310, 98340, 98370, 98380, 98380, 
    98380, 98360, 98350, 98330, 98350, 98310, 98300, 98290, 98280, 98260, 
    98240, 98230, 98200, 98200, 98210, 98190, 98170, 98160, 98140, 98100, 
    98120, 98160, 98150, 98130, 98130, 98170, 98270, 98370, 98500, 98620, 
    98710, 98800, 98870, 98940, 99040, 99090, 99180, 99260, 99340, 99410, 
    99480, 99550, 99630, 99700, 99760, 99810, 99870, 99920, 99970, 100010, 
    100050, 100090, 100120, 100140, 100150, 100170, 100110, 100100, 100090, 
    100080, 100060, 100060, 100050, 100010, 99990, 99970, 99990, 99960, 
    99870, 99830, 99780, 99720, 99650, 99600, 99540, 99540, 99510, 99480, 
    99440, 99430, 99400, 99370, 99330, 99320, 99300, 99280, 99260, 99260, 
    99230, 99220, 99190, 99160, 99130, 99070, 99030, 98970, 98910, 98890, 
    98860, 98840, 98810, 98780, 98780, 98810, 98840, 98860, 98880, 98930, 
    98970, 98990, 99060, 99110, 99170, 99220, 99270, 99280, 99290, 99320, 
    99350, 99400, 99460, 99490, 99530, 99550, 99580, 99620, 99620, 99630, 
    99600, 99590, 99590, 99570, 99560, 99540, 99540, 99540, 99520, 99480, 
    99440, 99420, 99410, 99390, 99340, 99330, 99330, 99360, 99360, 99380, 
    99400, 99420, 99410, 99410, 99440, 99460, 99500, 99560, 99630, 99710, 
    99790, 99900, 99950, 100000, 100020, 100100, 100140, 100170, 100230, 
    100270, 100290, 100350, 100390, 100450, 100480, 100520, 100570, 100600, 
    100630, 100640, 100660, 100690, 100690, 100740, 100780, 100750, 100760, 
    100720, 100700, 100600, 100530, 100440, 100330, 100260, 100150, 100060, 
    99980, 99840, 99690, 99530, 99370, 98990, 98910, 98580, 98160, 97810, 
    97390, 97050, 96820, 96600, 96440, 96320, 96210, 96150, 96070, 95990, 
    95970, 95980, 95990, 96070, 96140, 96240, 96310, 96380, 96480, 96550, 
    96610, 96690, 96790, 96910, 96960, 97060, 97150, 97210, 97260, 97320, 
    97370, 97400, 97400, 97390, 97400, 97420, 97410, 97450, 97430, 97450, 
    97450, 97450, 97490, 97490, 97530, 97580, 97620, 97710, 97730, 97760, 
    97830, 97860, 97930, 97980, 98040, 98110, 98170, 98210, 98280, 98350, 
    98430, 98500, 98550, 98610, 98640, 98660, 98680, 98710, 98750, 98790, 
    98830, 98850, 98860, 98910, 98950, 98990, 98980, 99030, 99050, 99060, 
    99080, 99090, 99110, 99110, 99120, 99130, 99130, 99100, 99070, 99050, 
    99030, 99000, 98980, 98970, 98960, 98950, 98970, 98990, 99010, 99030, 
    99020, 99050, 99100, 99130, 99150, 99180, 99210, 99230, 99270, 99290, 
    99320, 99360, 99360, 99390, 99430, 99470, 99530, 99540, 99570, 99610, 
    99620, 99670, 99710, 99710, 99730, 99720, 99760, 99800, 99820, 99840, 
    99860, 99890, 99940, 99950, 99990, 100020, 100060, 100070, 100070, 
    100090, 100080, 100070, 100050, 100070, 100070, 100090, 100120, 100140, 
    100140, 100110, 100080, 100050, 100020, 100010, 99940, 99890, 99800, 
    99770, 99730, 99670, 99610, 99510, 99450, 99380, 99330, 99240, 99180, 
    99130, 99020, 98970, 98850, 98770, 98650, 98490, 98390, 98270, 98230, 
    98160, 98160, 98180, 98230, 98180, 98160, 98170, 98170, 98170, 98110, 
    98160, 98180, 98170, 98140, 98060, 98000, 97870, 97910, 97820, 97890, 
    97970, 98100, 98280, 98450, 98610, 98730, 98780, 98840, 98910, 98960, 
    98980, 98990, 98980, 98980, 99010, 99060, 99110, 99190, 99260, 99340, 
    99470, 99560, 99660, 99720, 99800, 99840, 99960, 100050, 100130, 100210, 
    100280, 100340, 100420, 100460, 100520, 100530, 100560, 100540, 100560, 
    100590, 100630, 100630, 100650, 100660, 100690, 100690, 100740, 100770, 
    100780, 100780, 100790, 100820, 100860, 100870, 100880, 100880, 100890, 
    100920, 100910, 100900, 100900, 100870, 100820, 100790, 100740, 100680, 
    100670, 100650, 100600, 100560, 100570, 100530, 100500, 100480, 100460, 
    100430, 100420, 100400, 100410, 100430, 100410, 100420, 100400, 100350, 
    100290, 100230, 100200, 100160, 100100, 100050, 100030, 100010, 100000, 
    99990, 99950, 99930, 99920, 99940, 99970, 99990, 100010, 100060, 100100, 
    100140, 100180, 100220, 100260, 100290, 100340, 100390, 100430, 100450, 
    100490, 100490, 100530, 100570, 100600, 100610, 100600, 100590, 100590, 
    100590, 100580, 100550, 100510, 100480, 100450, 100410, 100400, 100360, 
    100320, 100260, 100210, 100180, 100150, 100090, 100040, 99980, 99930, 
    99940, 99870, 99840, 99790, 99750, 99680, 99640, 99580, 99540, 99500, 
    99460, 99410, 99360, 99310, 99240, 99200, 99190, 99160, 99140, 99100, 
    99050, 98990, 98980, 98980, 98980, 98990, 98960, 98940, 98930, 98920, 
    98950, 98980, 98960, 98980, 99020, 99000, 99020, 99080, 99110, 99100, 
    99170, 99210, 99270, 99310, 99360, 99410, 99460, 99500, 99540, 99600, 
    99650, 99710, 99760, 99780, 99790, 99790, 99810, 99820, 99870, 99910, 
    99950, 99980, 100010, 100070, 100070, 100080, 100100, 100050, 100060, 
    100100, 100090, 100070, 100040, 100010, 99970, 99960, 99920, 99900, 
    99860, 99800, 99720, 99650, 99560, 99490, 99440, 99410, 99360, 99300, 
    99260, 99200, 99150, 99130, 99090, 99060, 99030, 99000, 98980, 98970, 
    98980, 98990, 98980, 98980, 98990, 99010, 99030, 99030, 99030, 99040, 
    99060, 99090, 99130, 99160, 99180, 99170, 99210, 99210, 99240, 99260, 
    99250, 99270, 99310, 99350, 99390, 99400, 99420, 99450, 99450, 99460, 
    99470, 99490, 99480, 99470, 99500, 99530, 99560, 99620, 99660, 99660, 
    99690, 99690, 99740, 99760, 99760, 99780, 99860, 99940, 100020, 100070, 
    100150, 100210, 100240, 100290, 100320, 100350, 100400, 100400, 100440, 
    100460, 100530, 100580, 100600, 100600, 100640, 100670, 100670, 100650, 
    100650, 100650, 100650, 100680, 100680, 100700, 100690, 100680, 100680, 
    100710, 100720, 100720, 100730, 100740, 100760, 100810, 100830, 100820, 
    100840, 100850, 100870, 100870, 100900, 100880, 100880, 100880, 100880, 
    100900, 100910, 100930, 100930, 100910, 100900, 100890, 100870, 100860, 
    100840, 100840, 100850, 100850, 100870, 100880, 100930, 100930, 100940, 
    100980, 101000, 100980, 100950, 100990, 101010, 101040, 101020, 101040, 
    101050, 101050, 101070, 101080, 101100, 101100, 101070, 101070, 101090, 
    101110, 101110, 101100, 101060, 101040, 101050, 101040, 101030, 101030, 
    101050, 101080, 101090, 101100, 101150, 101150, 101170, 101210, 101220, 
    101240, 101240, 101240, 101220, 101230, 101230, 101240, 101220, 101210, 
    101220, 101230, 101210, 101220, 101190, 101160, 101130, 101110, 101090, 
    101080, 101080, 101080, 101030, 101010, 101010, 101020, 100980, 100960, 
    100930, 100870, 100850, 100810, 100760, 100710, 100660, 100570, 100500, 
    100430, 100330, 100210, 100100, 100010, 99930, 99860, 99810, 99730, 
    99650, 99560, 99500, 99480, 99440, 99450, 99490, 99490, 99520, 99510, 
    99500, 99520, 99530, 99530, 99560, 99550, 99520, 99500, 99540, 99580, 
    99600, 99610, 99610, 99620, 99620, 99650, 99650, 99680, 99710, 99740, 
    99810, 99910, 99990, 100090, 100160, 100260, 100350, 100420, 100500, 
    100560, 100620, 100680, 100720, 100780, 100800, 100830, 100870, 100900, 
    100930, 100950, 101000, 101030, 101000, 101010, 100990, 100990, 100980, 
    100910, 100850, 100810, 100750, 100720, 100700, 100680, 100640, 100550, 
    100440, 100340, 100290, 100290, 100310, 100330, 100350, 100380, 100370, 
    100320, 100270, 100340, 100340, 100340, 100350, 100250, 100270, 100280, 
    100250, 100220, 100170, 100100, 100050, 99980, 99940, 99860, 99810, 
    99800, 99750, 99670, 99590, 99530, 99450, 99370, 99280, 99210, 99120, 
    99030, 99000, 98910, 98810, 98730, 98650, 98550, 98520, 98460, 98360, 
    98330, 98380, 98450, 98450, 98480, 98450, 98440, 98390, 98340, 98300, 
    98260, 98170, 98100, 97960, 97850, 97780, 97730, 97730, 97660, 97530, 
    97480, 97490, 97450, 97480, 97490, 97530, 97540, 97580, 97550, 97520, 
    97490, 97480, 97530, 97590, 97710, 97810, 97970, 98090, 98170, 98250, 
    98380, 98470, 98540, 98670, 98810, 98950, 99060, 99160, 99250, 99330, 
    99440, 99560, 99640, 99740, 99840, 99930, 100000, 100060, 100110, 100120, 
    100130, 100120, 100110, 100140, 100160, 100190, 100220, 100260, 100250, 
    100250, 100280, 100270, 100270, 100260, 100250, 100250, 100250, 100250, 
    100270, 100230, 100190, 100170, 100150, 100150, 100140, 100160, 100190, 
    100200, 100220, 100220, 100270, 100280, 100300, 100270, 100280, 100270, 
    100260, 100240, 100220, 100220, 100190, 100180, 100160, 100160, 100160, 
    100160, 100150, 100160, 100160, 100150, 100160, 100200, 100210, 100230, 
    100230, 100220, 100240, 100230, 100250, 100250, 100240, 100220, 100240, 
    100260, 100280, 100290, 100310, 100330, 100360, 100350, 100360, 100390, 
    100370, 100390, 100390, 100400, 100420, 100460, 100460, 100500, 100510, 
    100580, 100600, 100610, 100620, 100620, 100630, 100640, 100670, 100690, 
    100730, 100730, 100740, 100730, 100770, 100830, 100850, 100860, 100860, 
    100880, 100910, 100890, 100850, 100850, 100890, 100870, 100840, 100880, 
    100850, 100860, 100840, 100840, 100880, 100910, 100890, 100890, 100900, 
    100930, 100950, 100970, 100970, 100970, 100980, 101020, 101030, 101070, 
    101100, 101160, 101180, 101200, 101240, 101270, 101270, 101280, 101330, 
    101320, 101360, 101370, 101440, 101460, 101500, 101490, 101470, 101460, 
    101450, 101470, 101460, 101450, 101480, 101470, 101490, 101490, 101450, 
    101420, 101430, 101380, 101330, 101360, 101340, 101320, 101300, 101290, 
    101270, 101240, 101190, 101150, 101100, 101060, 101020, 100990, 100980, 
    100970, 100940, 100930, 100930, 100880, 100860, 100830, 100790, 100760, 
    100740, 100720, 100670, 100690, 100670, 100670, 100670, 100640, 100590, 
    100570, 100550, 100550, 100530, 100510, 100500, 100470, 100490, 100500, 
    100520, 100510, 100500, 100480, 100510, 100500, 100560, 100560, 100590, 
    100610, 100610, 100630, 100660, 100660, 100660, 100690, 100670, 100690, 
    100670, 100670, 100670, 100670, 100680, 100670, 100670, 100650, 100600, 
    100580, 100570, 100530, 100510, 100490, 100490, 100470, 100460, 100480, 
    100490, 100500, 100450, 100410, 100410, 100430, 100450, 100470, 100480, 
    100490, 100520, 100560, 100600, 100630, 100660, 100700, 100730, 100760, 
    100800, 100820, 100830, 100880, 100930, 100970, 101000, 101030, 101060, 
    101080, 101090, 101130, 101150, 101160, 101200, 101220, 101240, 101270, 
    101300, 101350, 101370, 101390, 101430, 101460, 101470, 101490, 101540, 
    101570, 101620, 101670, 101710, 101740, 101760, 101770, 101790, 101790, 
    101800, 101830, 101880, 101900, 101930, 101960, 101970, 102000, 102040, 
    102030, 102040, 102040, 102070, 102070, 102090, 102120, 102160, 102210, 
    102240, 102260, 102290, 102280, 102300, 102300, 102300, 102310, 102310, 
    102310, 102320, 102320, 102290, 102240, 102200, 102160, 102110, 102050, 
    101990, 101930, 101870, 101800, 101770, 101770, 101750, 101720, 101700, 
    101670, 101650, 101640, 101640, 101650, 101670, 101680, 101720, 101740, 
    101770, 101810, 101830, 101830, 101830, 101840, 101860, 101870, 101870, 
    101860, 101910, 101950, 101950, 101950, 101920, 101900, 101870, 101860, 
    101850, 101830, 101810, 101850, 101860, 101870, 101890, 101890, 101860, 
    101840, 101790, 101760, 101750, 101740, 101730, 101710, 101720, 101750, 
    101740, 101740, 101730, 101710, 101700, 101670, 101640, 101600, 101600, 
    101600, 101580, 101550, 101530, 101510, 101500, 101490, 101470, 101450, 
    101430, 101450, 101420, 101420, 101440, 101470, 101490, 101500, 101510, 
    101530, 101560, 101560, 101570, 101590, 101610, 101630, 101650, 101660, 
    101680, 101670, 101700, 101710, 101720, 101750, 101740, 101750, 101760, 
    101760, 101800, 101810, 101820, 101830, 101850, 101890, 101920, 101920, 
    101950, 101950, 101960, 101980, 102000, 102020, 102050, 102060, 102050, 
    102060, 102090, 102090, 102080, 102090, 102110, 102140, 102160, 102180, 
    102200, 102220, 102230, 102240, 102240, 102230, 102220, 102230, 102230, 
    102230, 102240, 102260, 102280, 102300, 102290, 102300, 102310, 102300, 
    102290, 102270, 102270, 102280, 102280, 102300, 102310, 102340, 102360, 
    102360, 102370, 102370, 102380, 102390, 102420, 102440, 102470, 102500, 
    102520, 102540, 102520, 102540, 102530, 102530, 102520, 102520, 102520, 
    102510, 102520, 102530, 102520, 102530, 102510, 102510, 102500, 102450, 
    102410, 102410, 102400, 102420, 102380, 102370, 102340, 102330, 102330, 
    102310, 102230, 102200, 102130, 102130, 102120, 102090, 102060, 102030, 
    102000, 101970, 101900, 101800, 101740, 101660, 101580, 101510, 101450, 
    101350, 101220, 101140, 101110, 101060, 101000, 100920, 100830, 100770, 
    100670, 100630, 100600, 100600, 100600, 100590, 100600, 100590, 100610, 
    100590, 100610, 100620, 100640, 100660, 100650, 100680, 100730, 100740, 
    100750, 100770, 100790, 100800, 100800, 100800, 100810, 100800, 100810, 
    100830, 100870, 100900, 100910, 100910, 100910, 100910, 100920, 100930, 
    100950, 100970, 101000, 101040, 101100, 101150, 101200, 101240, 101270, 
    101330, 101350, 101380, 101390, 101390, 101410, 101450, 101490, 101540, 
    101590, 101640, 101680, 101700, 101710, 101730, 101750, 101790, 101830, 
    101840, 101890, 101940, 101960, 101970, 101980, 102000, 102030, 102050, 
    102060, 102060, 102050, 102040, 102040, 102040, 102010, 101990, 101950, 
    101950, 101940, 101930, 101940, 101950, 101970, 102010, 102070, 102110, 
    102200, 102290, 102360, 102400, 102430, 102460, 102470, 102450, 102440, 
    102460, 102500, 102540, 102550, 102570, 102570, 102560, 102550, 102570, 
    102570, 102560, 102500, 102460, 102450, 102410, 102370, 102340, 102310, 
    102280, 102230, 102180, 102140, 102100, 102070, 102060, 102040, 102030, 
    102050, 102030, 101980, 101960, 101950, 101930, 101920, 101910, 101880, 
    101850, 101860, 101870, 101860, 101840, 101800, 101770, 101750, 101740, 
    101740, 101700, 101660, 101650, 101650, 101680, 101670, 101640, 101580, 
    101520, 101450, 101420, 101390, 101380, 101340, 101320, 101280, 101280, 
    101290, 101250, 101220, 101230, 101210, 101210, 101220, 101260, 101290, 
    101280, 101280, 101300, 101310, 101300, 101280, 101260, 101250, 101240, 
    101240, 101230, 101230, 101200, 101160, 101160, 101150, 101100, 101080, 
    101080, 101030, 101000, 101020, 100970, 100960, 100940, 100930, 100910, 
    100940, 101010, 101080, 101180, 101200, 101300, 101410, 101530, 101580, 
    101670, 101740, 101820, 101870, 101910, 101940, 102000, 102040, 102060, 
    102090, 102140, 102160, 102180, 102220, 102260, 102300, 102330, 102350, 
    102360, 102340, 102340, 102340, 102320, 102280, 102320, 102360, 102360, 
    102280, 102240, 102230, 102190, 102170, 102110, 102070, 102030, 102000, 
    101960, 101920, 101890, 101860, 101820, 101730, 101640, 101590, 101520, 
    101450, 101420, 101410, 101450, 101510, 101540, 101540, 101540, 101540, 
    101520, 101480, 101490, 101520, 101540, 101550, 101560, 101610, 101640, 
    101700, 101730, 101750, 101770, 101780, 101790, 101830, 101840, 101850, 
    101850, 101840, 101850, 101840, 101810, 101780, 101750, 101670, 101610, 
    101550, 101510, 101460, 101400, 101340, 101290, 101210, 101150, 101080, 
    101030, 100980, 100940, 100910, 100880, 100840, 100810, 100790, 100770, 
    100750, 100730, 100730, 100760, 100790, 100810, 100800, 100820, 100830, 
    100860, 100880, 100930, 101000, 101040, 101060, 101100, 101150, 101180, 
    101220, 101250, 101300, 101360, 101400, 101430, 101460, 101490, 101530, 
    101540, 101570, 101610, 101610, 101620, 101640, 101670, 101680, 101700, 
    101710, 101710, 101700, 101700, 101710, 101700, 101710, 101700, 101670, 
    101670, 101690, 101670, 101680, 101670, 101630, 101640, 101630, 101620, 
    101630, 101610, 101620, 101650, 101680, 101730, 101780, 101800, 101830, 
    101840, 101860, 101900, 101950, 101990, 102020, 102070, 102160, 102190, 
    102220, 102270, 102360, 102390, 102380, 102450, 102480, 102550, 102550, 
    102650, 102730, 102800, 102810, 102900, 102960, 102970, 103000, 103040, 
    103090, 103150, 103190, 103220, 103260, 103320, 103370, 103400, 103410, 
    103420, 103450, 103460, 103460, 103470, 103460, 103480, 103490, 103480, 
    103440, 103440, 103400, 103370, 103350, 103320, 103290, 103260, 103220, 
    103180, 103170, 103140, 103080, 103040, 103000, 102940, 102870, 102830, 
    102780, 102730, 102690, 102660, 102620, 102600, 102580, 102540, 102500, 
    102450, 102390, 102330, 102270, 102220, 102170, 102120, 102070, 102010, 
    101980, 101920, 101850, 101810, 101750, 101710, 101650, 101580, 101530, 
    101510, 101460, 101440, 101430, 101390, 101350, 101320, 101290, 101260, 
    101230, 101220, 101210, 101200, 101200, 101220, 101210, 101230, 101250, 
    101210, 101180, 101190, 101190, 101190, 101210, 101220, 101290, 101330, 
    101400, 101410, 101430, 101490, 101540, 101590, 101640, 101650, 101680, 
    101740, 101750, 101790, 101830, 101870, 101860, 101850, 101870, 101900, 
    101890, 101880, 101910, 101920, 101920, 101950, 101990, 101980, 101980, 
    102020, 102060, 102080, 102090, 102110, 102140, 102130, 102150, 102160, 
    102170, 102160, 102170, 102150, 102140, 102110, 102100, 102090, 102080, 
    102070, 102080, 102120, 102150, 102160, 102170, 102170, 102160, 102130, 
    102110, 102090, 102070, 102050, 102030, 102030, 102020, 102020, 101970, 
    101940, 101910, 101870, 101830, 101790, 101760, 101730, 101720, 101730, 
    101680, 101620, 101580, 101560, 101520, 101430, 101370, 101320, 101280, 
    101250, 101200, 101160, 101070, 100990, 100870, 100740, 100620, 100530, 
    100420, 100340, 100270, 100220, 100180, 100180, 100160, 100150, 100150, 
    100130, 100120, 100110, 100090, 100080, 100060, 100090, 100110, 100130, 
    100140, 100150, 100130, 100150, 100160, 100160, 100150, 100160, 100190, 
    100210, 100250, 100290, 100330, 100360, 100370, 100360, 100380, 100370, 
    100370, 100370, 100390, 100420, 100420, 100400, 100400, 100410, 100410, 
    100410, 100420, 100450, 100460, 100500, 100500, 100530, 100580, 100600, 
    100630, 100650, 100670, 100700, 100720, 100720, 100750, 100780, 100800, 
    100820, 100850, 100880, 100890, 100910, 100920, 100930, 100940, 100950, 
    100940, 100940, 100940, 100930, 100930, 100930, 100940, 100910, 100880, 
    100850, 100840, 100810, 100780, 100750, 100760, 100730, 100710, 100720, 
    100710, 100690, 100660, 100670, 100660, 100630, 100620, 100610, 100580, 
    100580, 100570, 100570, 100570, 100560, 100550, 100540, 100570, 100580, 
    100540, 100530, 100460, 100420, 100400, 100360, 100350, 100310, 100290, 
    100270, 100250, 100220, 100190, 100170, 100140, 100120, 100100, 100090, 
    100090, 100060, 100060, 100040, 100010, 99980, 99940, 99920, 99890, 
    99890, 99910, 99930, 99910, 99880, 99840, 99810, 99820, 99790, 99760, 
    99730, 99700, 99680, 99670, 99660, 99660, 99650, 99640, 99610, 99600, 
    99580, 99510, 99470, 99440, 99400, 99360, 99320, 99290, 99210, 99150, 
    99130, 99100, 99080, 99030, 99000, 99010, 98960, 98940, 98910, 98890, 
    98850, 98770, 98740, 98660, 98590, 98580, 98550, 98480, 98440, 98420, 
    98390, 98360, 98360, 98370, 98410, 98470, 98540, 98620, 98730, 98810, 
    98900, 98970, 99010, 99060, 99070, 99080, 99120, 99160, 99220, 99260, 
    99320, 99390, 99470, 99530, 99570, 99610, 99650, 99680, 99670, 99720, 
    99760, 99800, 99830, 99910, 99980, 100030, 100130, 100200, 100280, 
    100360, 100420, 100420, 100440, 100470, 100570, 100580, 100600, 100640, 
    100650, 100680, 100730, 100760, 100770, 100770, 100770, 100760, 100780, 
    100780, 100770, 100740, 100740, 100770, 100750, 100690, 100690, 100660, 
    100590, 100510, 100470, 100420, 100350, 100330, 100270, 100260, 100330, 
    100330, 100270, 100280, 100300, 100370, 100430, 100470, 100480, 100570, 
    100610, 100630, 100640, 100630, 100610, 100600, 100570, 100540, 100500, 
    100490, 100440, 100430, 100430, 100410, 100380, 100350, 100330, 100320, 
    100310, 100270, 100260, 100240, 100260, 100260, 100270, 100270, 100260, 
    100250, 100240, 100220, 100200, 100200, 100190, 100170, 100170, 100170, 
    100170, 100160, 100140, 100110, 100080, 100050, 100030, 100010, 100000, 
    99980, 99950, 99950, 99940, 99960, 99970, 99970, 99970, 99950, 99960, 
    99930, 99950, 99950, 99940, 99960, 100000, 99990, 100000, 100010, 100030, 
    100040, 100070, 100090, 100130, 100170, 100220, 100270, 100340, 100400, 
    100460, 100530, 100590, 100640, 100710, 100740, 100770, 100840, 100910, 
    100960, 101000, 101060, 101120, 101170, 101220, 101270, 101320, 101320, 
    101330, 101330, 101380, 101410, 101440, 101530, 101590, 101630, 101680, 
    101720, 101750, 101770, 101800, 101840, 101870, 101890, 101900, 101930, 
    101930, 101940, 101930, 101930, 101940, 101930, 101900, 101910, 101930, 
    101920, 101940, 101950, 101960, 101950, 101930, 101940, 101920, 101890, 
    101860, 101830, 101820, 101800, 101780, 101760, 101730, 101720, 101680, 
    101640, 101610, 101540, 101500, 101470, 101440, 101400, 101380, 101340, 
    101330, 101290, 101230, 101170, 101140, 101090, 101080, 101070, 101040, 
    101030, 101020, 101010, 100990, 100950, 100920, 100880, 100850, 100780, 
    100730, 100720, 100690, 100710, 100680, 100640, 100660, 100630, 100610, 
    100580, 100570, 100560, 100510, 100480, 100480, 100460, 100460, 100470, 
    100450, 100430, 100410, 100380, 100340, 100300, 100270, 100260, 100230, 
    100220, 100210, 100200, 100170, 100130, 100110, 100070, 100030, 100010, 
    99980, 99930, 99890, 99860, 99830, 99800, 99740, 99710, 99670, 99630, 
    99580, 99550, 99520, 99480, 99450, 99440, 99420, 99420, 99400, 99410, 
    99410, 99400, 99370, 99340, 99320, 99320, 99300, 99300, 99280, 99290, 
    99290, 99270, 99270, 99240, 99200, 99170, 99160, 99130, 99070, 99120, 
    99100, 99100, 99100, 99090, 99080, 99040, 99080, 99120, 99140, 99150, 
    99180, 99190, 99200, 99270, 99330, 99330, 99310, 99290, 99260, 99270, 
    99280, 99310, 99350, 99410, 99480, 99550, 99630, 99710, 99780, 99850, 
    99920, 100000, 100070, 100150, 100240, 100340, 100450, 100550, 100640, 
    100740, 100830, 100910, 100990, 101060, 101110, 101180, 101220, 101290, 
    101370, 101430, 101530, 101590, 101650, 101700, 101730, 101760, 101780, 
    101810, 101800, 101750, 101720, 101700, 101640, 101590, 101560, 101510, 
    101460, 101410, 101390, 101360, 101360, 101370, 101370, 101350, 101370, 
    101360, 101370, 101340, 101330, 101330, 101310, 101310, 101310, 101300, 
    101290, 101270, 101250, 101230, 101250, 101250, 101270, 101330, 101350, 
    101350, 101400, 101440, 101470, 101470, 101520, 101560, 101580, 101600, 
    101650, 101690, 101750, 101790, 101820, 101880, 101910, 101940, 101990, 
    102000, 102010, 102040, 102040, 102050, 102080, 102090, 102110, 102140, 
    102170, 102220, 102240, 102240, 102220, 102220, 102220, 102210, 102190, 
    102180, 102110, 102040, 102010, 101990, 101960, 101900, 101830, 101760, 
    101700, 101620, 101540, 101480, 101420, 101360, 101330, 101280, 101240, 
    101190, 101120, 101060, 101000, 100950, 100870, 100770, 100680, 100590, 
    100440, 100320, 100190, 100090, 99970, 99850, 99710, 99520, 99380, 99260, 
    99220, 99220, 99310, 99330, 99310, 99310, 99310, 99310, 99430, 99440, 
    99480, 99530, 99370, 99390, 99440, 99470, 99510, 99510, 99550, 99600, 
    99640, 99680, 99740, 99810, 99900, 99990, 100080, 100170, 100250, 100330, 
    100430, 100460, 100520, 100580, 100630, 100680, 100720, 100750, 100780, 
    100790, 100750, 100690, 100660, 100630, 100640, 100660, 100710, 100740, 
    100780, 100820, 100870, 100920, 100940, 100940, 100970, 100970, 100960, 
    100940, 100890, 100820, 100780, 100740, 100690, 100670, 100610, 100550, 
    100500, 100430, 100340, 100210, 100090, 99970, 99870, 99760, 99670, 
    99530, 99420, 99270, 99100, 98990, 98900, 98780, 98650, 98500, 98350, 
    98250, 98170, 98080, 98040, 98040, 98020, 97980, 97940, 97960, 97910, 
    97860, 97840, 97810, 97820, 97770, 97820, 97820, 97770, 97730, 97700, 
    97720, 97720, 97720, 97710, 97750, 97780, 97790, 97780, 97780, 97830, 
    97790, 97810, 97800, 97830, 97880, 97940, 97980, 98050, 98120, 98170, 
    98200, 98260, 98270, 98360, 98370, 98390, 98400, 98450, 98490, 98520, 
    98560, 98580, 98620, 98620, 98630, 98630, 98620, 98600, 98590, 98590, 
    98600, 98620, 98630, 98610, 98620, 98610, 98620, 98630, 98640, 98630, 
    98620, 98620, 98630, 98650, 98650, 98670, 98690, 98690, 98730, 98730, 
    98750, 98760, 98800, 98860, 98910, 98990, 99030, 99080, 99130, 99190, 
    99250, 99300, 99380, 99430, 99480, 99530, 99580, 99630, 99690, 99720, 
    99740, 99780, 99810, 99830, 99850, 99860, 99840, 99830, 99810, 99810, 
    99830, 99820, 99810, 99800, 99790, 99750, 99700, 99640, 99610, 99590, 
    99600, 99600, 99630, 99630, 99660, 99690, 99710, 99780, 99840, 99910, 
    99980, 100050, 100140, 100240, 100300, 100390, 100460, 100520, 100580, 
    100640, 100680, 100690, 100720, 100750, 100770, 100800, 100840, 100910, 
    100920, 100930, 100940, 100940, 100910, 100840, 100810, 100800, 100790, 
    100780, 100720, 100680, 100630, 100580, 100510, 100450, 100410, 100410, 
    100390, 100380, 100380, 100380, 100380, 100370, 100380, 100380, 100390, 
    100390, 100400, 100410, 100410, 100420, 100450, 100490, 100540, 100590, 
    100600, 100570, 100560, 100570, 100600, 100590, 100570, 100560, 100570, 
    100580, 100580, 100600, 100610, 100610, 100620, 100620, 100630, 100620, 
    100620, 100620, 100660, 100680, 100700, 100690, 100690, 100730, 100720, 
    100730, 100730, 100720, 100720, 100730, 100730, 100750, 100770, 100780, 
    100780, 100770, 100770, 100760, 100770, 100760, 100790, 100800, 100820, 
    100830, 100850, 100840, 100860, 100870, 100880, 100890, 100900, 100880, 
    100870, 100860, 100870, 100860, 100900, 100900, 100860, 100820, 100820, 
    100760, 100750, 100710, 100660, 100650, 100600, 100560, 100530, 100520, 
    100520, 100500, 100500, 100450, 100470, 100440, 100440, 100400, 100410, 
    100380, 100370, 100370, 100360, 100310, 100270, 100260, 100230, 100200, 
    100150, 100150, 100170, 100190, 100230, 100280, 100330, 100350, 100350, 
    100350, 100320, 100320, 100310, 100310, 100300, 100320, 100330, 100330, 
    100320, 100300, 100290, 100310, 100300, 100310, 100330, 100330, 100340, 
    100360, 100390, 100410, 100430, 100440, 100450, 100470, 100510, 100500, 
    100510, 100540, 100550, 100580, 100600, 100590, 100590, 100580, 100570, 
    100580, 100560, 100530, 100510, 100480, 100470, 100450, 100410, 100350, 
    100300, 100250, 100200, 100140, 100090, 100000, 99950, 99860, 99780, 
    99700, 99650, 99590, 99520, 99430, 99360, 99260, 99170, 99080, 99020, 
    98960, 98920, 98890, 98870, 98860, 98850, 98830, 98810, 98820, 98820, 
    98830, 98840, 98860, 98880, 98900, 98910, 98910, 98940, 98940, 98940, 
    98950, 98950, 98970, 98980, 99020, 99050, 99090, 99120, 99140, 99180, 
    99220, 99250, 99280, 99300, 99350, 99380, 99420, 99450, 99480, 99530, 
    99540, 99580, 99600, 99640, 99680, 99710, 99750, 99770, 99800, 99830, 
    99860, 99880, 99890, 99880, 99880, 99850, 99810, 99790, 99770, 99780, 
    99770, 99760, 99770, 99770, 99760, 99770, 99760, 99760, 99780, 99800, 
    99810, 99820, 99840, 99860, 99880, 99910, 99920, 99950, 99960, 99980, 
    100020, 100070, 100120, 100190, 100280, 100370, 100450, 100520, 100600, 
    100680, 100740, 100810, 100880, 100930, 100990, 101020, 101050, 101030, 
    101010, 100980, 100970, 100960, 100970, 101030, 101120, 101220, 101330, 
    101430, 101530, 101660, 101750, 101790, 101830, 101870, 101880, 101890, 
    101830, 101820, 101710, 101650, 101610, 101530, 101480, 101410, 101360, 
    101340, 101350, 101360, 101390, 101430, 101490, 101580, 101660, 101750, 
    101850, 101960, 102010, 102030, 102160, 102200, 102220, 102240, 102230, 
    102230, 102240, 102230, 102230, 102140, 102090, 102020, 101920, 101860, 
    101730, 101600, 101480, 101350, 101190, 100990, 100850, 100800, 100750, 
    100770, 100790, 100780, 100750, 100730, 100730, 100730, 100700, 100660, 
    100640, 100670, 100660, 100660, 100670, 100590, 100530, 100500, 100450, 
    100460, 100480, 100550, 100580, 100660, 100690, 100730, 100790, 100830, 
    100880, 100950, 101000, 101080, 101120, 101220, 101260, 101330, 101360, 
    101380, 101410, 101460, 101460, 101500, 101480, 101490, 101550, 101560, 
    101610, 101610, 101590, 101630, 101620, 101650, 101670, 101680, 101660, 
    101650, 101680, 101700, 101720, 101720, 101720, 101730, 101700, 101690, 
    101670, 101670, 101660, 101650, 101670, 101700, 101710, 101710, 101670, 
    101660, 101670, 101680, 101670, 101650, 101620, 101600, 101580, 101580, 
    101590, 101590, 101570, 101550, 101540, 101520, 101500, 101510, 101510, 
    101460, 101470, 101490, 101540, 101540, 101510, 101450, 101430, 101410, 
    101380, 101340, 101270, 101180, 101100, 101040, 100980, 100930, 100880, 
    100790, 100750, 100700, 100630, 100590, 100530, 100490, 100480, 100470, 
    100430, 100390, 100410, 100410, 100420, 100420, 100450, 100480, 100470, 
    100440, 100430, 100470, 100500, 100540, 100550, 100550, 100570, 100590, 
    100610, 100620, 100640, 100640, 100640, 100650, 100680, 100720, 100740, 
    100740, 100710, 100710, 100720, 100730, 100720, 100720, 100720, 100720, 
    100740, 100740, 100720, 100720, 100710, 100700, 100700, 100680, 100650, 
    100590, 100570, 100540, 100510, 100490, 100470, 100430, 100370, 100340, 
    100290, 100210, 100160, 100090, 100020, 99950, 99890, 99810, 99720, 
    99650, 99580, 99530, 99520, 99500, 99500, 99500, 99540, 99550, 99580, 
    99640, 99650, 99680, 99730, 99770, 99810, 99840, 99840, 99860, 99880, 
    99940, 99970, 100000, 100050, 100090, 100130, 100160, 100200, 100240, 
    100260, 100300, 100340, 100380, 100410, 100460, 100500, 100560, 100590, 
    100620, 100660, 100720, 100750, 100790, 100810, 100880, 100920, 101000, 
    101060, 101130, 101170, 101210, 101250, 101290, 101320, 101360, 101390, 
    101430, 101490, 101530, 101610, 101660, 101720, 101750, 101780, 101800, 
    101830, 101860, 101890, 101940, 101990, 102020, 102030, 102060, 102100, 
    102120, 102130, 102130, 102150, 102150, 102160, 102150, 102180, 102190, 
    102200, 102220, 102170, 102140, 102130, 102130, 102100, 102080, 102070, 
    102090, 102090, 102070, 102080, 102080, 102060, 102050, 102020, 101970, 
    101910, 101880, 101800, 101760, 101710, 101660, 101610, 101590, 101560, 
    101530, 101490, 101450, 101410, 101370, 101320, 101280, 101250, 101220, 
    101170, 101100, 101030, 100960, 100880, 100800, 100720, 100630, 100560, 
    100510, 100440, 100360, 100260, 100160, 100070, 99970, 99900, 99820, 
    99730, 99650, 99580, 99520, 99460, 99420, 99380, 99310, 99290, 99270, 
    99260, 99270, 99260, 99270, 99310, 99340, 99360, 99380, 99390, 99410, 
    99410, 99400, 99380, 99330, 99270, 99250, 99240, 99250, 99230, 99240, 
    99240, 99260, 99300, 99320, 99370, 99410, 99450, 99500, 99520, 99560, 
    99600, 99620, 99640, 99650, 99660, 99680, 99700, 99710, 99730, 99740, 
    99770, 99780, 99830, 99870, 99900, 99950, 99970, 100010, 100000, 100030, 
    100090, 100110, 100140, 100170, 100220, 100250, 100270, 100250, 100220, 
    100210, 100240, 100230, 100240, 100220, 100210, 100210, 100210, 100210, 
    100200, 100210, 100210, 100190, 100190, 100180, 100180, 100170, 100180, 
    100200, 100220, 100230, 100230, 100220, 100260, 100270, 100290, 100320, 
    100360, 100380, 100380, 100410, 100440, 100440, 100440, 100470, 100480, 
    100490, 100500, 100520, 100530, 100540, 100580, 100610, 100630, 100620, 
    100640, 100680, 100710, 100740, 100770, 100790, 100820, 100840, 100830, 
    100820, 100830, 100850, 100880, 100860, 100810, 100820, 100800, 100810, 
    100800, 100800, 100790, 100770, 100740, 100720, 100690, 100620, 100580, 
    100490, 100420, 100320, 100210, 100100, 99960, 99850, 99730, 99590, 
    99420, 99300, 99110, 98960, 98800, 98710, 98590, 98470, 98340, 98220, 
    98130, 98000, 97880, 97790, 97670, 97510, 97450, 97400, 97420, 97440, 
    97490, 97530, 97580, 97650, 97690, 97750, 97750, 97900, 97970, 98040, 
    98120, 98210, 98320, 98410, 98510, 98580, 98650, 98760, 98840, 98920, 
    98980, 99050, 99110, 99160, 99220, 99260, 99330, 99380, 99400, 99410, 
    99420, 99440, 99440, 99440, 99410, 99370, 99320, 99280, 99240, 99230, 
    99200, 99160, 99120, 99090, 99060, 99010, 99000, 99010, 99040, 99050, 
    99070, 99110, 99170, 99240, 99320, 99400, 99490, 99580, 99660, 99780, 
    99890, 100000, 100110, 100200, 100320, 100440, 100540, 100630, 100740, 
    100810, 100840, 100840, 100860, 100860, 100860, 100870, 100840, 100790, 
    100780, 100750, 100680, 100610, 100550, 100500, 100480, 100480, 100490, 
    100470, 100500, 100520, 100550, 100550, 100500, 100490, 100460, 100420, 
    100380, 100330, 100290, 100250, 100200, 100140, 100070, 100010, 99960, 
    99900, 99890, 99910, 99940, 100010, 100080, 100190, 100290, 100390, 
    100450, 100570, 100670, 100770, 100900, 101030, 101100, 101250, 101350, 
    101450, 101540, 101630, 101700, 101770, 101810, 101830, 101880, 101890, 
    101910, 101950, 101970, 101970, 101980, 101980, 101980, 102000, 101980, 
    101990, 101970, 101920, 101930, 101930, 101920, 101890, 101840, 101830, 
    101790, 101770, 101720, 101650, 101660, 101660, 101660, 101680, 101700, 
    101710, 101730, 101770, 101820, 101830, 101880, 101950, 102000, 102040, 
    102090, 102170, 102220, 102250, 102290, 102370, 102420, 102460, 102480, 
    102490, 102520, 102530, 102540, 102580, 102610, 102600, 102590, 102580, 
    102570, 102560, 102520, 102500, 102460, 102450, 102450, 102420, 102400, 
    102390, 102390, 102370, 102340, 102310, 102300, 102280, 102260, 102250, 
    102260, 102270, 102290, 102290, 102290, 102310, 102300, 102300, 102290, 
    102290, 102290, 102290, 102300, 102300, 102290, 102270, 102270, 102250, 
    102260, 102240, 102160, 102120, 102160, 102140, 102130, 102110, 102090, 
    102070, 102020, 101980, 101940, 101900, 101870, 101830, 101750, 101740, 
    101710, 101680, 101660, 101660, 101640, 101650, 101650, 101640, 101630, 
    101630, 101630, 101640, 101670, 101700, 101750, 101800, 101830, 101880, 
    101910, 101920, 101940, 101980, 102000, 102040, 102100, 102160, 102190, 
    102240, 102270, 102320, 102390, 102410, 102450, 102460, 102470, 102490, 
    102520, 102540, 102540, 102540, 102540, 102530, 102500, 102470, 102420, 
    102360, 102320, 102250, 102200, 102170, 102140, 102130, 102140, 102150, 
    102140, 102120, 102140, 102130, 102100, 102110, 102110, 102140, 102160, 
    102130, 102100, 102080, 102070, 102060, 102050, 102030, 102020, 102020, 
    102020, 102020, 102010, 102010, 102000, 102000, 102000, 101980, 101960, 
    101950, 101920, 101900, 101900, 101880, 101870, 101890, 101840, 101830, 
    101820, 101810, 101790, 101810, 101810, 101800, 101820, 101820, 101830, 
    101820, 101860, 101840, 101850, 101870, 101890, 101920, 101930, 101950, 
    101970, 102020, 102040, 102070, 102090, 102110, 102140, 102160, 102180, 
    102220, 102240, 102270, 102280, 102320, 102350, 102360, 102400, 102420, 
    102440, 102450, 102450, 102470, 102490, 102500, 102500, 102520, 102530, 
    102540, 102560, 102560, 102550, 102540, 102550, 102520, 102520, 102500, 
    102490, 102500, 102490, 102480, 102470, 102450, 102430, 102420, 102400, 
    102360, 102360, 102350, 102340, 102330, 102320, 102300, 102290, 102270, 
    102260, 102250, 102220, 102210, 102200, 102200, 102200, 102200, 102200, 
    102210, 102220, 102230, 102230, 102250, 102260, 102270, 102270, 102280, 
    102280, 102280, 102310, 102330, 102330, 102330, 102310, 102300, 102320, 
    102310, 102300, 102310, 102310, 102320, 102330, 102320, 102330, 102330, 
    102330, 102330, 102370, 102380, 102360, 102350, 102360, 102360, 102360, 
    102370, 102400, 102430, 102470, 102480, 102510, 102530, 102560, 102580, 
    102610, 102630, 102630, 102650, 102680, 102690, 102670, 102640, 102660, 
    102670, 102690, 102690, 102690, 102690, 102680, 102660, 102620, 102590, 
    102550, 102540, 102490, 102440, 102410, 102380, 102330, 102300, 102270, 
    102240, 102210, 102160, 102130, 102090, 102030, 101990, 101950, 101880, 
    101820, 101750, 101680, 101620, 101540, 101470, 101420, 101370, 101350, 
    101310, 101280, 101290, 101360, 101390, 101420, 101450, 101470, 101490, 
    101480, 101460, 101440, 101430, 101410, 101380, 101350, 101310, 101260, 
    101220, 101190, 101130, 101090, 101020, 100970, 100920, 100900, 100880, 
    100860, 100840, 100830, 100820, 100820, 100800, 100790, 100760, 100740, 
    100730, 100730, 100730, 100740, 100750, 100750, 100770, 100750, 100770, 
    100760, 100770, 100760, 100740, 100750, 100750, 100770, 100780, 100780, 
    100750, 100740, 100740, 100700, 100700, 100710, 100710, 100710, 100720, 
    100740, 100740, 100750, 100740, 100750, 100750, 100760, 100740, 100720, 
    100700, 100700, 100690, 100700, 100700, 100690, 100670, 100670, 100660, 
    100670, 100660, 100650, 100640, 100630, 100640, 100640, 100680, 100680, 
    100700, 100700, 100720, 100720, 100720, 100710, 100720, 100730, 100730, 
    100760, 100780, 100790, 100830, 100850, 100870, 100890, 100900, 100910, 
    100930, 100920, 100940, 100960, 100990, 101020, 101030, 101030, 101040, 
    101030, 101020, 101020, 100990, 101000, 101000, 101000, 101000, 101010, 
    101020, 101040, 101030, 101040, 101030, 101040, 101050, 101080, 101100, 
    101130, 101140, 101170, 101180, 101200, 101210, 101220, 101240, 101250, 
    101250, 101270, 101280, 101300, 101320, 101350, 101380, 101410, 101410, 
    101420, 101420, 101430, 101440, 101460, 101470, 101470, 101500, 101500, 
    101520, 101530, 101520, 101520, 101490, 101490, 101500, 101480, 101470, 
    101470, 101470, 101450, 101430, 101430, 101440, 101440, 101420, 101360, 
    101320, 101270, 101240, 101160, 101120, 101080, 101020, 100970, 100960, 
    100940, 100920, 100900, 100870, 100840, 100810, 100770, 100730, 100680, 
    100630, 100580, 100530, 100450, 100340, 100240, 100120, 100010, 99930, 
    99820, 99720, 99640, 99570, 99530, 99490, 99470, 99440, 99400, 99330, 
    99380, 99410, 99520, 99660, 99710, 99710, 99740, 99810, 99820, 99800, 
    99840, 99850, 99900, 99900, 99920, 99950, 100000, 100060, 100100, 100180, 
    100230, 100310, 100390, 100460, 100520, 100600, 100700, 100780, 100860, 
    100940, 101010, 101090, 101150, 101190, 101230, 101280, 101320, 101350, 
    101420, 101480, 101530, 101550, 101580, 101590, 101600, 101610, 101590, 
    101570, 101550, 101540, 101530, 101500, 101500, 101480, 101440, 101420, 
    101400, 101360, 101330, 101300, 101280, 101270, 101260, 101250, 101250, 
    101240, 101260, 101240, 101250, 101230, 101190, 101170, 101160, 101160, 
    101170, 101180, 101160, 101150, 101150, 101140, 101120, 101100, 101110, 
    101140, 101120, 101100, 101110, 101120, 101080, 101040, 100990, 100960, 
    100920, 100910, 100870, 100810, 100750, 100710, 100720, 100700, 100700, 
    100760, 100780, 100840, 100890, 100960, 101000, 101040, 101100, 101160, 
    101240, 101300, 101370, 101440, 101500, 101560, 101590, 101640, 101650, 
    101710, 101730, 101770, 101790, 101860, 101900, 101950, 102000, 102040, 
    102080, 102110, 102130, 102150, 102180, 102200, 102250, 102300, 102350, 
    102400, 102410, 102440, 102470, 102480, 102500, 102480, 102500, 102520, 
    102530, 102540, 102560, 102600, 102620, 102630, 102620, 102630, 102620, 
    102600, 102580, 102570, 102560, 102570, 102580, 102560, 102560, 102560, 
    102550, 102540, 102540, 102530, 102550, 102550, 102580, 102590, 102620, 
    102630, 102650, 102660, 102690, 102730, 102760, 102770, 102790, 102810, 
    102840, 102880, 102920, 102970, 103000, 103040, 103080, 103110, 103120, 
    103140, 103170, 103190, 103210, 103240, 103270, 103290, 103310, 103340, 
    103360, 103370, 103370, 103390, 103390, 103390, 103390, 103420, 103430, 
    103460, 103480, 103480, 103470, 103500, 103490, 103470, 103480, 103480, 
    103490, 103480, 103490, 103500, 103490, 103480, 103470, 103470, 103440, 
    103400, 103370, 103350, 103320, 103290, 103270, 103250, 103220, 103200, 
    103200, 103170, 103150, 103150, 103110, 103090, 103080, 103080, 103070, 
    103040, 103070, 103030, 103000, 102960, 102890, 102840, 102790, 102750, 
    102690, 102700, 102730, 102730, 102730, 102730, 102720, 102710, 102720, 
    102690, 102680, 102670, 102660, 102610, 102580, 102550, 102530, 102500, 
    102490, 102440, 102390, 102340, 102330, 102300, 102290, 102290, 102270, 
    102240, 102260, 102260, 102230, 102220, 102210, 102200, 102220, 102220, 
    102240, 102280, 102310, 102310, 102320, 102320, 102310, 102260, 102250, 
    102240, 102210, 102190, 102180, 102150, 102140, 102100, 102090, 102050, 
    102010, 102010, 101980, 101950, 101920, 101910, 101910, 101890, 101870, 
    101850, 101840, 101780, 101760, 101710, 101680, 101640, 101580, 101560, 
    101530, 101510, 101490, 101460, 101440, 101440, 101430, 101410, 101380, 
    101380, 101400, 101410, 101410, 101420, 101430, 101420, 101430, 101420, 
    101430, 101440, 101450, 101460, 101460, 101440, 101450, 101480, 101490, 
    101500, 101510, 101530, 101520, 101540, 101540, 101550, 101560, 101580, 
    101610, 101640, 101680, 101700, 101720, 101740, 101760, 101780, 101780, 
    101780, 101780, 101810, 101820, 101830, 101830, 101840, 101840, 101840, 
    101840, 101850, 101830, 101830, 101800, 101780, 101770, 101770, 101790, 
    101750, 101720, 101680, 101660, 101630, 101600, 101580, 101560, 101540, 
    101510, 101490, 101480, 101460, 101420, 101390, 101380, 101380, 101370, 
    101360, 101370, 101410, 101450, 101520, 101550, 101600, 101640, 101700, 
    101750, 101800, 101840, 101890, 101940, 101990, 102020, 102070, 102110, 
    102180, 102210, 102250, 102290, 102310, 102330, 102340, 102380, 102420, 
    102460, 102490, 102520, 102530, 102560, 102570, 102570, 102580, 102570, 
    102550, 102530, 102500, 102500, 102490, 102480, 102460, 102460, 102430, 
    102400, 102400, 102360, 102320, 102300, 102270, 102240, 102210, 102170, 
    102170, 102140, 102120, 102100, 102080, 102050, 102040, 102010, 101990, 
    101950, 101960, 101940, 101940, 101920, 101920, 101890, 101870, 101870, 
    101850, 101830, 101830, 101810, 101810, 101820, 101800, 101780, 101790, 
    101810, 101810, 101800, 101770, 101770, 101760, 101770, 101790, 101810, 
    101820, 101820, 101840, 101850, 101860, 101860, 101860, 101870, 101850, 
    101870, 101860, 101870, 101840, 101840, 101820, 101800, 101760, 101750, 
    101740, 101690, 101670, 101660, 101650, 101630, 101600, 101590, 101590, 
    101590, 101580, 101560, 101570, 101540, 101550, 101540, 101530, 101560, 
    101570, 101580, 101600, 101630, 101640, 101670, 101680, 101680, 101710, 
    101740, 101760, 101820, 101880, 101900, 101920, 101930, 101960, 102000, 
    102010, 102040, 102060, 102090, 102120, 102150, 102170, 102180, 102200, 
    102210, 102210, 102220, 102210, 102200, 102190, 102180, 102190, 102200, 
    102160, 102130, 102110, 102070, 102060, 102030, 101970, 101940, 101890, 
    101860, 101830, 101780, 101760, 101730, 101690, 101670, 101650, 101650, 
    101600, 101560, 101550, 101550, 101570, 101590, 101590, 101590, 101580, 
    101590, 101600, 101580, 101580, 101560, 101570, 101570, 101580, 101590, 
    101590, 101560, 101550, 101540, 101530, 101510, 101480, 101460, 101420, 
    101410, 101420, 101400, 101400, 101390, 101380, 101350, 101350, 101350, 
    101360, 101360, 101370, 101390, 101410, 101440, 101450, 101470, 101490, 
    101500, 101520, 101520, 101530, 101550, 101570, 101600, 101610, 101650, 
    101630, 101640, 101630, 101640, 101630, 101630, 101620, 101590, 101570, 
    101530, 101500, 101480, 101410, 101370, 101340, 101280, 101220, 101150, 
    101140, 101080, 101010, 100970, 100920, 100900, 100840, 100780, 100740, 
    100720, 100660, 100640, 100620, 100610, 100590, 100570, 100550, 100490, 
    100410, 100370, 100320, 100350, 100430, 100450, 100500, 100480, 100450, 
    100420, 100430, 100420, 100490, 100540, 100570, 100590, 100620, 100650, 
    100710, 100750, 100760, 100860, 100910, 100960, 101020, 101070, 101140, 
    101140, 101220, 101270, 101310, 101340, 101370, 101420, 101490, 101510, 
    101600, 101560, 101580, 101600, 101630, 101610, 101600, 101590, 101580, 
    101550, 101520, 101490, 101450, 101410, 101360, 101310, 101260, 101190, 
    101140, 101100, 101060, 100980, 100910, 100870, 100810, 100770, 100720, 
    100690, 100680, 100670, 100640, 100640, 100650, 100650, 100680, 100690, 
    100740, 100760, 100790, 100830, 100870, 100910, 100910, 100930, 100940, 
    100930, 100930, 100960, 100980, 101010, 101020, 101060, 101080, 101090, 
    101090, 101120, 101130, 101160, 101160, 101170, 101190, 101230, 101280, 
    101310, 101360, 101370, 101400, 101380, 101400, 101390, 101390, 101380, 
    101380, 101410, 101380, 101360, 101370, 101400, 101380, 101370, 101360, 
    101360, 101360, 101360, 101400, 101410, 101430, 101460, 101490, 101510, 
    101530, 101590, 101590, 101640, 101680, 101700, 101720, 101740, 101790, 
    101820, 101820, 101820, 101850, 101880, 101880, 101890, 101910, 101940, 
    101930, 101950, 101950, 101960, 101940, 101940, 101920, 101910, 101900, 
    101900, 101900, 101890, 101870, 101870, 101860, 101840, 101820, 101810, 
    101780, 101780, 101780, 101780, 101780, 101760, 101750, 101770, 101770, 
    101780, 101790, 101790, 101790, 101820, 101830, 101840, 101860, 101880, 
    101900, 101920, 101940, 101980, 102000, 102040, 102060, 102080, 102110, 
    102150, 102170, 102210, 102230, 102240, 102270, 102270, 102280, 102280, 
    102290, 102290, 102310, 102340, 102360, 102350, 102360, 102380, 102380, 
    102390, 102390, 102390, 102400, 102410, 102420, 102440, 102450, 102460, 
    102460, 102480, 102480, 102490, 102470, 102470, 102470, 102460, 102480, 
    102470, 102470, 102470, 102470, 102470, 102470, 102470, 102470, 102470, 
    102460, 102460, 102460, 102480, 102500, 102500, 102500, 102500, 102490, 
    102490, 102470, 102450, 102460, 102460, 102450, 102430, 102410, 102400, 
    102390, 102360, 102360, 102320, 102320, 102300, 102270, 102240, 102220, 
    102220, 102190, 102180, 102150, 102130, 102120, 102100, 102100, 102070, 
    102050, 102030, 102030, 101980, 101950, 101940, 101910, 101890, 101870, 
    101850, 101830, 101830, 101800, 101780, 101750, 101740, 101730, 101700, 
    101680, 101670, 101680, 101680, 101680, 101680, 101680, 101680, 101670, 
    101670, 101670, 101660, 101660, 101660, 101650, 101660, 101680, 101660, 
    101680, 101670, 101690, 101690, 101690, 101700, 101720, 101720, 101720, 
    101710, 101700, 101710, 101700, 101690, 101690, 101710, 101710, 101710, 
    101720, 101710, 101710, 101710, 101700, 101710, 101710, 101710, 101700, 
    101700, 101700, 101700, 101690, 101690, 101670, 101660, 101630, 101610, 
    101560, 101530, 101500, 101480, 101450, 101430, 101400, 101360, 101320, 
    101300, 101280, 101250, 101220, 101180, 101140, 101130, 101110, 101070, 
    101050, 101050, 101030, 101020, 100990, 100960, 100940, 100930, 100910, 
    100900, 100880, 100860, 100850, 100840, 100810, 100780, 100770, 100780, 
    100740, 100730, 100740, 100740, 100740, 100740, 100740, 100740, 100750, 
    100760, 100780, 100780, 100770, 100750, 100760, 100770, 100780, 100790, 
    100800, 100800, 100820, 100840, 100840, 100870, 100890, 100910, 100930, 
    100950, 100980, 101000, 101010, 101050, 101080, 101100, 101120, 101160, 
    101200, 101230, 101260, 101320, 101370, 101400, 101440, 101470, 101470, 
    101490, 101550, 101590, 101610, 101600, 101630, 101630, 101670, 101670, 
    101690, 101720, 101730, 101740, 101740, 101730, 101730, 101730, 101710, 
    101710, 101710, 101700, 101700, 101690, 101680, 101650, 101640, 101620, 
    101620, 101600, 101590, 101610, 101640, 101640, 101660, 101660, 101670, 
    101670, 101670, 101680, 101660, 101670, 101660, 101640, 101640, 101660, 
    101650, 101630, 101620, 101610, 101620, 101590, 101580, 101580, 101580, 
    101590, 101580, 101610, 101630, 101650, 101650, 101660, 101670, 101670, 
    101690, 101690, 101680, 101700, 101730, 101750, 101760, 101790, 101800, 
    101820, 101840, 101830, 101830, 101830, 101830, 101860, 101870, 101890, 
    101910, 101930, 101910, 101920, 101920, 101920, 101910, 101910, 101910, 
    101910, 101940, 101940, 101940, 101940, 101930, 101910, 101930, 101940, 
    101900, 101910, 101900, 101890, 101880, 101900, 101900, 101920, 101930, 
    101930, 101940, 101950, 101960, 101970, 101990, 102010, 102030, 102050, 
    102110, 102140, 102170, 102180, 102210, 102240, 102270, 102290, 102340, 
    102380, 102420, 102470, 102500, 102510, 102540, 102540, 102540, 102560, 
    102560, 102570, 102580, 102590, 102600, 102620, 102640, 102660, 102680, 
    102710, 102730, 102730, 102730, 102720, 102730, 102760, 102780, 102810, 
    102840, 102820, 102830, 102830, 102830, 102840, 102820, 102820, 102810, 
    102810, 102800, 102840, 102830, 102820, 102820, 102790, 102760, 102710, 
    102690, 102640, 102610, 102550, 102520, 102490, 102470, 102430, 102400, 
    102370, 102310, 102270, 102250, 102200, 102190, 102140, 102110, 102130, 
    102060, 102000, 101970, 101910, 101830, 101760, 101680, 101620, 101550, 
    101480, 101430, 101340, 101260, 101190, 101150, 101110, 101080, 101040, 
    100990, 100950, 100930, 100940, 100930, 100960, 100970, 100980, 101030, 
    101050, 101050, 101070, 101070, 101070, 101080, 101060, 101060, 101060, 
    101010, 100980, 100930, 100890, 100830, 100780, 100740, 100700, 100670, 
    100640, 100620, 100600, 100630, 100630, 100660, 100710, 100730, 100780, 
    100820, 100820, 100880, 100930, 100980, 101050, 101090, 101160, 101170, 
    101210, 101250, 101290, 101310, 101350, 101360, 101400, 101430, 101480, 
    101510, 101560, 101590, 101620, 101650, 101670, 101670, 101670, 101680, 
    101700, 101720, 101750, 101790, 101800, 101800, 101820, 101830, 101830, 
    101850, 101840, 101850, 101880, 101890, 101910, 101920, 101960, 101980, 
    101980, 101990, 101990, 101980, 101990, 101980, 101970, 101970, 101990, 
    102020, 102040, 102050, 102060, 102050, 102030, 102040, 102030, 102040, 
    102050, 102060, 102070, 102100, 102110, 102130, 102130, 102160, 102170, 
    102170, 102170, 102170, 102160, 102180, 102200, 102220, 102240, 102230, 
    102230, 102230, 102220, 102200, 102190, 102180, 102190, 102180, 102170, 
    102170, 102170, 102180, 102160, 102110, 102080, 102010, 101940, 101900, 
    101860, 101850, 101830, 101790, 101730, 101700, 101690, 101670, 101610, 
    101560, 101510, 101500, 101470, 101430, 101410, 101380, 101360, 101360, 
    101380, 101370, 101340, 101340, 101310, 101320, 101320, 101310, 101330, 
    101320, 101350, 101340, 101360, 101360, 101350, 101350, 101360, 101360, 
    101370, 101400, 101430, 101450, 101470, 101500, 101510, 101530, 101560, 
    101590, 101590, 101610, 101640, 101670, 101710, 101730, 101760, 101750, 
    101750, 101750, 101750, 101760, 101770, 101780, 101790, 101830, 101880, 
    101890, 101900, 101930, 101960, 101980, 101980, 101980, 101980, 102000, 
    101980, 101970, 101980, 101930, 101910, 101870, 101850, 101770, 101690, 
    101620, 101600, 101590, 101600, 101620, 101640, 101630, 101600, 101600, 
    101590, 101560, 101540, 101510, 101490, 101450, 101430, 101440, 101450, 
    101440, 101450, 101460, 101480, 101490, 101490, 101500, 101530, 101540, 
    101560, 101590, 101610, 101630, 101630, 101600, 101580, 101580, 101580, 
    101550, 101510, 101510, 101490, 101480, 101480, 101480, 101500, 101500, 
    101520, 101510, 101540, 101580, 101590, 101620, 101650, 101690, 101740, 
    101780, 101800, 101820, 101850, 101890, 101920, 101940, 101950, 101980, 
    102000, 102020, 102040, 102060, 102070, 102060, 102040, 102000, 101960, 
    101910, 101870, 101820, 101790, 101750, 101700, 101650, 101590, 101540, 
    101480, 101430, 101370, 101300, 101240, 101220, 101180, 101150, 101100, 
    101050, 101020, 100970, 100940, 100910, 100880, 100870, 100860, 100850, 
    100810, 100820, 100810, 100790, 100770, 100770, 100730, 100690, 100640, 
    100590, 100530, 100490, 100490, 100480, 100470, 100440, 100420, 100430, 
    100430, 100430, 100430, 100470, 100470, 100510, 100520, 100590, 100650, 
    100700, 100740, 100810, 100890, 100960, 101010, 101070, 101110, 101130, 
    101180, 101200, 101210, 101200, 101230, 101220, 101190, 101170, 101130, 
    101130, 101100, 101070, 101060, 101040, 101010, 100990, 100970, 100960, 
    100950, 100920, 100910, 100900, 100890, 100870, 100860, 100860, 100870, 
    100880, 100880, 100890, 100910, 100920, 100940, 100940, 100930, 100920, 
    100940, 100980, 101000, 101020, 101040, 101050, 101060, 101040, 101060, 
    101060, 101050, 101060, 101070, 101080, 101090, 101110, 101140, 101170, 
    101180, 101160, 101140, 101140, 101150, 101150, 101150, 101170, 101160, 
    101170, 101160, 101150, 101150, 101140, 101140, 101140, 101140, 101150, 
    101170, 101190, 101210, 101240, 101270, 101270, 101300, 101300, 101300, 
    101320, 101340, 101350, 101360, 101380, 101400, 101430, 101440, 101450, 
    101470, 101460, 101460, 101460, 101450, 101450, 101470, 101480, 101490, 
    101480, 101510, 101490, 101480, 101480, 101460, 101460, 101430, 101420, 
    101410, 101410, 101420, 101420, 101420, 101430, 101400, 101400, 101390, 
    101380, 101370, 101360, 101340, 101350, 101330, 101320, 101300, 101270, 
    101230, 101190, 101150, 101120, 101090, 101010, 100940, 100900, 100880, 
    100850, 100820, 100800, 100760, 100720, 100690, 100630, 100580, 100530, 
    100490, 100440, 100400, 100370, 100320, 100280, 100250, 100210, 100160, 
    100130, 100100, 100060, 100040, 100020, 100000, 99980, 99990, 99990, 
    100010, 99980, 99970, 99960, 99960, 99980, 99980, 99990, 100000, 100010, 
    100020, 100050, 100060, 100070, 100080, 100100, 100110, 100130, 100150, 
    100180, 100190, 100210, 100250, 100270, 100290, 100310, 100350, 100360, 
    100400, 100430, 100440, 100510, 100560, 100610, 100630, 100690, 100780, 
    100830, 100880, 100920, 100970, 101000, 101050, 101090, 101130, 101180, 
    101230, 101260, 101270, 101270, 101280, 101270, 101270, 101270, 101260, 
    101270, 101310, 101340, 101350, 101360, 101370, 101390, 101400, 101410, 
    101410, 101360, 101380, 101400, 101430, 101460, 101480, 101500, 101510, 
    101530, 101530, 101530, 101530, 101620, 101630, 101590, 101590, 101640, 
    101590, 101580, 101650, 101670, 101660, 101660, 101660, 101680, 101700, 
    101720, 101740, 101770, 101810, 101830, 101840, 101850, 101860, 101880, 
    101890, 101930, 101950, 101850, 101870, 101880, 101920, 101930, 101940, 
    101940, 101920, 101910, 101920, 101920, 101900, 101900, 101910, 101920, 
    101920, 101890, 101890, 101890, 101890, 101870, 101860, 101850, 101840, 
    101840, 101860, 101870, 101890, 101880, 101850, 101840, 101800, 101770, 
    101740, 101730, 101760, 101770, 101800, 101820, 101830, 101850, 101860, 
    101870, 101870, 101880, 101910, 101950, 101980, 102020, 102050, 102070, 
    102100, 102100, 102100, 102100, 102100, 102090, 102070, 102050, 102040, 
    102060, 102050, 102040, 102030, 102100, 102090, 101960, 101930, 101900, 
    101870, 101850, 101840, 101840, 101830, 101810, 101780, 101760, 101740, 
    101730, 101710, 101690, 101670, 101670, 101670, 101680, 101670, 101660, 
    101670, 101670, 101690, 101700, 101720, 101770, 101760, 101780, 101810, 
    101830, 101910, 101940, 101970, 101990, 102030, 102070, 102100, 102130, 
    102150, 102140, 102150, 102090, 102110, 102130, 102150, 102130, 102100, 
    102090, 102080, 102070, 102060, 102040, 102030, 102000, 102000, 101980, 
    101950, 101940, 101920, 101900, 101860, 101810, 101780, 101750, 101730, 
    101720, 101720, 101720, 101720, 101720, 101660, 101650, 101630, 101610, 
    101590, 101590, 101580, 101560, 101540, 101500, 101480, 101470, 101480, 
    101450, 101420, 101390, 101360, 101350, 101350, 101330, 101320, 101310, 
    101310, 101290, 101250, 101220, 101210, 101200, 101170, 101170, 101160, 
    101150, 101140, 101150, 101130, 101100, 101100, 101090, 101070, 101050, 
    101030, 101020, 101010, 101020, 101010, 101000, 100960, 100930, 101090, 
    101080, 101060, 101020, 100990, 100970, 100810, 100800, 100810, 100770, 
    100770, 100750, 100730, 100710, 100700, 100690, 100680, 100670, 100670, 
    100670, 100650, 100670, 100680, 100680, 100680, 100690, 100700, 100700, 
    100690, 100690, 100690, 100710, 100710, 100710, 100710, 100710, 100700, 
    100700, 100720, 100730, 100740, 100750, 100760, 100770, 100780, 100780, 
    100780, 100760, 100760, 100760, 100770, 100770, 100780, 100790, 100800, 
    100800, 100820, 100850, 100850, 100860, 100870, 100880, 100900, 100920, 
    100940, 100970, 100990, 101010, 101020, 101010, 101030, 101060, 101050, 
    101090, 101120, 101150, 101170, 101180, 101180, 101160, 101150, 101160, 
    101190, 101190, 101170, 101150, 101150, 101140, 101120, 101130, 101130, 
    101130, 101160, 101160, 101140, 101180, 101150, 101130, 101130, 101090, 
    101060, 101040, 101050, 101040, 101010, 101000, 100970, 100960, 100960, 
    100960, 100960, 100950, 100940, 100940, 100930, 100930, 100920, 100920, 
    100910, 100880, 100860, 100860, 100850, 100830, 100830, 100790, 100780, 
    100780, 100770, 100800, 100800, 100790, 100770, 100760, 100730, 100740, 
    100830, 100810, 100820, 100830, 100850, 100880, 100920, 100960, 100860, 
    100870, 100880, 100900, 100930, 100960, 100990, 101020, 101040, 101060, 
    101090, 101130, 101150, 101190, 101190, 101190, 101240, 101300, 101330, 
    101480, 101500, 101530, 101560, 101560, 101470, 101470, 101460, 101460, 
    101450, 101450, 101450, 101440, 101440, 101420, 101400, 101380, 101360, 
    101370, 101350, 101320, 101290, 101290, 101300, 101300, 101290, 101290, 
    101290, 101300, 101280, 101240, 101200, 101300, 101250, 101210, 101110, 
    101100, 101160, 101070, 101060, 101040, 101000, 100970, 100950, 101000, 
    100990, 100880, 100880, 100890, 100880, 100880, 100890, 100890, 100870, 
    100850, 100800, 100780, 100720, 100700, 100690, 100690, 100700, 100700, 
    100670, 100650, 100650, 100650, 100720, 100710, 100700, 100670, 100690, 
    100710, 100690, 100680, 100670, 100660, 100670, 100690, 100680, 100700, 
    100720, 100750, 100790, 100810, 100830, 100840, 100850, 100860, 100860, 
    100870, 100890, 101070, 101090, 101030, 101060, 101100, 101030, 101060, 
    101090, 101120, 101140, 101160, 101180, 101200, 101200, 101220, 101240, 
    101260, 101270, 101290, 101310, 101330, 101340, 101360, 101400, 101420, 
    101440, 101490, 101520, 101560, 101590, 101620, 101650, 101680, 101710, 
    101720, 101720, 101720, 101750, 101770, 101790, 101800, 101820, 101840, 
    101850, 101860, 101860, 101840, 101840, 101840, 101840, 101850, 101860, 
    101880, 101910, 101890, 101890, 101910, 101900, 101890, 101880, 101870, 
    101860, 101850, 101860, 101870, 101870, 101860, 101860, 101850, 101840, 
    101810, 101780, 101750, 101740, 101730, 101740, 101740, 101740, 101740, 
    101830, 101800, 101720, 101700, 101680, 101660, 101640, 101620, 101600, 
    101590, 101570, 101550, 101520, 101490, 101470, 101430, 101390, 101340, 
    101310, 101280, 101230, 101180, 101130, 101090, 101050, 101020, 101000, 
    100920, 100890, 100880, 100810, 100790, 100770, 100740, 100690, 100680, 
    100670, 100630, 100610, 100590, 100560, 100530, 100560, 100560, 100550, 
    100530, 100510, 100480, 100490, 100470, 100480, 100490, 100490, 100510, 
    100560, 100630, 100670, 100690, 100710, 100730, 100750, 100780, 100780, 
    100800, 100820, 100860, 100900, 100940, 100990, 101060, 101140, 101180, 
    101240, 101320, 101360, 101390, 101430, 101460, 101460, 101450, 101450, 
    101450, 101440, 101410, 101390, 101310, 101240, 101180, 101090, 101000, 
    100920, 100820, 100760, 100750, 100640, 100690, 100730, 100780, 100810, 
    100850, 100860, 100900, 100900, 100940, 100970, 101030, 101050, 101060, 
    101060, 101080, 101080, 101080, 101070, 101080, 101060, 101040, 101010, 
    101000, 101010, 101020, 101020, 101010, 101030, 101020, 101020, 101050, 
    101040, 101050, 101090, 101110, 101120, 101140, 101170, 101190, 101200, 
    101220, 101220, 101230, 101220, 101240, 101250, 101260, 101270, 101300, 
    101300, 101320, 101310, 101290, 101270, 101260, 101250, 101240, 101230, 
    101220, 101220, 101240, 101230, 101220, 101200, 101150, 101110, 101100, 
    101110, 101070, 101060, 101050, 101040, 101020, 101000, 100990, 100990, 
    100980, 100980, 100950, 100950, 100940, 100920, 100910, 100900, 100900, 
    100910, 100910, 100900, 100890, 100880, 100870, 100860, 100910, 100900, 
    100890, 100870, 100870, 100880, 100870, 100850, 100760, 100750, 100750, 
    100740, 100740, 100750, 100770, 100790, 100830, 100850, 100940, 100960, 
    100980, 100990, 101000, 101020, 101030, 100930, 100950, 100990, 101010, 
    101030, 101050, 101070, 101080, 101090, 101110, 101120, 101120, 101140, 
    101150, 101180, 101200, 101200, 101200, 101180, 101160, 101190, 101160, 
    101130, 101130, 101080, 101050, 101020, 100990, 100980, 100950, 100890, 
    100830, 100760, 100700, 100650, 100580, 100560, 100520, 100480, 100450, 
    100380, 100310, 100240, 100170, 100110, 100030, 99970, 99940, 99950, 
    99900, 99890, 99890, 99920, 99930, 99950, 99980, 100060, 100120, 100200, 
    100340, 100430, 100540, 100650, 100700, 100780, 100830, 100930, 101000, 
    101050, 101100, 101140, 101200, 101260, 101310, 101320, 101380, 101400, 
    101420, 101430, 101400, 101410, 101410, 101390, 101400, 101390, 101360, 
    101340, 101330, 101300, 101260, 101210, 101150, 101100, 101060, 101000, 
    100930, 100860, 100790, 100700, 100610, 100520, 100400, 100290, 100160, 
    100050, 99970, 99920, 99880, 99850, 99830, 99810, 99800, 99790, 99780, 
    99780, 99780, 99770, 99790, 99820, 99840, 99860, 99880, 99940, 99960, 
    99960, 99960, 99970, 99980, 100000, 100020, 100030, 100030, 100010, 
    100020, 100030, 100030, 100020, 100010, 100000, 99990, 99970, 99970, 
    99970, 99970, 99970, 99970, 100040, 100050, 100050, 100040, 100030, 
    100000, 99860, 99830, 99800, 99770, 99740, 99730, 99680, 99680, 99680, 
    99690, 99710, 99740, 99780, 99840, 99880, 99920, 99960, 100020, 100080, 
    100150, 100370, 100350, 100440, 100520, 100610, 100680, 100720, 100790, 
    100820, 100870, 100900, 100940, 100970, 101000, 101010, 101020, 101020, 
    100960, 100870, 100820, 100710, 100740, 100680, 100600, 100520, 100410, 
    100270, 100160, 100060, 99920, 99790, 99750, 99530, 99390, 99210, 99040, 
    98840, 98660, 98450, 98300, 98250, 98250, 98240, 98230, 98220, 98230, 
    98260, 98340, 98400, 98470, 98550, 98680, 98800, 98950, 99100, 99190, 
    99370, 99600, 99780, 99960, 100090, 100210, 100310, 100380, 100450, 
    100510, 100590, 100680, 100730, 100820, 100890, 100950, 101020, 101120, 
    101200, 101190, 101270, 101320, 101360, 101470, 101510, 101630, 101650, 
    101670, 101730, 101750, 101770, 101770, 101790, 101760, 101760, 101740, 
    101720, 101700, 101660, 101630, 101600, 101530, 101440, 101360, 101310, 
    101230, 101170, 101130, 101090, 101040, 100990, 100930, 100860, 100790, 
    100690, 100640, 100570, 100520, 100500, 100490, 100470, 100450, 100380, 
    100300, 100220, 100140, 100070, 99980, 99980, 99930, 99910, 99900, 99900, 
    99900, 99850, 99890, 99950, 99900, 99870, 99880, 99920, 99960, 100000, 
    100040, 100080, 100050, 100130, 100190, 100170, 100150, 100140, 100130, 
    100120, 100110, 100110, 100130, 100170, 100200, 100230, 100240, 100210, 
    100210, 100150, 100130, 100520, 100520, 100520, 100520, 100500, 100460, 
    100070, 100040, 100010, 99980, 99950, 99930, 99910, 99890, 99860, 99850, 
    99880, 99910, 99930, 99970, 99980, 99990, 100010, 100020, 100060, 100070, 
    100100, 100160, 100180, 100190, 100210, 100240, 100260, 100290, 100320, 
    100350, 100380, 100430, 100450, 100480, 100500, 100520, 100570, 100590, 
    100620, 100700, 100760, 100800, 100830, 100850, 100860, 100860, 100870, 
    100900, 100930, 100960, 101000, 101060, 101080, 101100, 101180, 101180, 
    101200, 101240, 101280, 101320, 101300, 101370, 101410, 101450, 101510, 
    101560, 101600, 101650, 101690, 101730, 101770, 101820, 101880, 101940, 
    101990, 102160, 102180, 102180, 102150, 102180, 102190, 102170, 102210, 
    102240, 102240, 102250, 102240, 102250, 102250, 102220, 102210, 102200, 
    102190, 102140, 102120, 102100, 102090, 102080, 102060, 102020, 101990, 
    101980, 101940, 101930, 101940, 101950, 101970, 101980, 102000, 102010, 
    102030, 102040, 102010, 102000, 101990, 101980, 101960, 101940, 101950, 
    101940, 101930, 101910, 101890, 101860, 101830, 101800, 101780, 101750, 
    101720, 101700, 101690, 101680, 101680, 101670, 101640, 101600, 101520, 
    101470, 101390, 101370, 101350, 101280, 101250, 101210, 101190, 101160, 
    101140, 101050, 101000, 100940, 100910, 100880, 100830, 100780, 100740, 
    100720, 100710, 100670, 100620, 100550, 100520, 100470, 100400, 100320, 
    100240, 100170, 100080, 100010, 99920, 99840, 99750, 99650, 99650, 99440, 
    99340, 99270, 99170, 99070, 99010, 98920, 98850, 98830, 98800, 98760, 
    98720, 98710, 98650, 98610, 98590, 98570, 98550, 98540, 98520, 98510, 
    98490, 98480, 98480, 98510, 98550, 98590, 98630, 98650, 98700, 98710, 
    98720, 98790, 98870, 98930, 98960, 99000, 99130, 99080, 99130, 99180, 
    99230, 99270, 99310, 99340, 99380, 99410, 99450, 99460, 99490, 99510, 
    99520, 99550, 99560, 99580, 99610, 99690, 99680, 99710, 99700, 99720, 
    99730, 99770, 99780, 99800, 99790, 99820, 99910, 99880, 99910, 99930, 
    99930, 99950, 99970, 99990, 100020, 100060, 100110, 100160, 100200, 
    100240, 100300, 100340, 100400, 100460, 100510, 100550, 100590, 100640, 
    100700, 100750, 100810, 100870, 100950, 100990, 101050, 101120, 101180, 
    101270, 101300, 101340, 101350, 101330, 101350, 101330, 101300, 101280, 
    101270, 101300, 101480, 101410, 101460, 101490, 101520, 101540, 101580, 
    101610, 101620, 101630, 101640, 101770, 101770, 101750, 101760, 101710, 
    101640, 101630, 101580, 101550, 101510, 101460, 101410, 101320, 101260, 
    101190, 101100, 101020, 100930, 100850, 100770, 100670, 100570, 100470, 
    100360, 100250, 100150, 100090, 100050, 100040, 100070, 100100, 100090, 
    100130, 100180, 100230, 100260, 100290, 100320, 100460, 100390, 100430, 
    100480, 100620, 100620, 100700, 100790, 100870, 100950, 101100, 101100, 
    101180, 101260, 101350, 101410, 101470, 101580, 101630, 101680, 101720, 
    101770, 101790, 101760, 101740, 101750, 101740, 101730, 101740, 101750, 
    101750, 101690, 101620, 101590, 101550, 101480, 101400, 101350, 101270, 
    101290, 101330, 101290, 101300, 101290, 101270, 101280, 101250, 101300, 
    101270, 101280, 101290, 101310, 101330, 101360, 101380, 101390, 101460, 
    101540, 101600, 101650, 101750, 101760, 101770, 101810, 101830, 101840, 
    101830, 101800, 101690, 101640, 101520, 101340, 101250, 101190, 101170, 
    101240, 101360, 101450, 101570, 101690, 101810, 101910, 101990, 102090, 
    102180, 102270, 102320, 102410, 102480, 102580, 102660, 102730, 102790, 
    102820, 102850, 102890, 102950, 103020, 103070, 103120, 103190, 103250, 
    103280, 103310, 103340, 103380, 103400, 103380, 103370, 103420, 103460, 
    103490, 103520, 103540, 103550, 103590, 103630, 103660, 103670, 103660, 
    103700, 103710, 103690, 103760, 103750, 103680, 103700, 103710, 103710, 
    103700, 103690, 103680, 103670, 103650, 103650, 103650, 103640, 103650, 
    103630, 103600, 103590, 103570, 103550, 103530, 103510, 103490, 103460, 
    103420, 103400, 103380, 103340, 103310, 103280, 103230, 103170, 103120, 
    103080, 103120, 103000, 102970, 102940, 102890, 102860, 102820, 102770, 
    102720, 102670, 102610, 102550, 102520, 102490, 102490, 102460, 102380, 
    102340, 102290, 102250, 102200, 102140, 102080, 102040, 102010, 102010, 
    101990, 101970, 101960, 101970, 101970, 101950, 101920, 101920, 101920, 
    101910, 101930, 101950, 101970, 101980, 102020, 102040, 102040, 102030, 
    102020, 102020, 102000, 101990, 101990, 101990, 101980, 101970, 101970, 
    101980, 101960, 101960, 101940, 101920, 101910, 101910, 101900, 101890, 
    101880, 101860, 101850, 101810, 101770, 101740, 101730, 101680, 101640, 
    101600, 101570, 101540, 101500, 101460, 101430, 101420, 101420, 101410, 
    101410, 101400, 101440, 101450, 101470, 101500, 101540, 101570, 101580, 
    101590, 101610, 101630, 101640, 101640, 101630, 101630, 101620, 101610, 
    101620, 101640, 101650, 101680, 101700, 101730, 101740, 101760, 101780, 
    101810, 101830, 101860, 101880, 101900, 101920, 101930, 101940, 101940, 
    101930, 101930, 101950, 101930, 101930, 101930, 101930, 101950, 101970, 
    101980, 101980, 101990, 101990, 101990, 101990, 102000, 102020, 102040, 
    102060, 102070, 102150, 102190, 102270, 102310, 102340, 102360, 102390, 
    102410, 102410, 102410, 102420, 102440, 102430, 102440, 102440, 102420, 
    102390, 102370, 102340, 102300, 102260, 102250, 102240, 102200, 102160, 
    102230, 102200, 102060, 102020, 101980, 101960, 101910, 101880, 101850, 
    101830, 101810, 101800, 101770, 101740, 101720, 101690, 101630, 101620, 
    101590, 101560, 101540, 101510, 101570, 101440, 101400, 101360, 101300, 
    101280, 101230, 101210, 101190, 101170, 101170, 101180, 101200, 101240, 
    101260, 101290, 101330, 101380, 101390, 101420, 101440, 101410, 101490, 
    101520, 101550, 101580, 101600, 101610, 101630, 101650, 101680, 101690, 
    101710, 101870, 101760, 101780, 101800, 101830, 101860, 101890, 101910, 
    101930, 101940, 101940, 102070, 102070, 102120, 102100, 102050, 102010, 
    101990, 101830, 101810, 101790, 101770, 101720, 101660, 101640, 101610, 
    101590, 101600, 101580, 101580, 101570, 101560, 101540, 101530, 101540, 
    101540, 101760, 101700, 101710, 101700, 101530, 101530, 101530, 101520, 
    101520, 101490, 101470, 101450, 101450, 101450, 101440, 101440, 101480, 
    101500, 101520, 101530, 101530, 101530, 101550, 101550, 101570, 101580, 
    101590, 101610, 101620, 101640, 101650, 101660, 101640, 101620, 101640, 
    101650, 101640, 101620, 101640, 101670, 101700, 101730, 101740, 101780, 
    101790, 101770, 101910, 101730, 101700, 101670, 101850, 101820, 101590, 
    101560, 101560, 101530, 101500, 101450, 101390, 101370, 101330, 101290, 
    101260, 101310, 101290, 101200, 101180, 101150, 101110, 101050, 101010, 
    100970, 100930, 100890, 100850, 100940, 100910, 100880, 100870, 100830, 
    100800, 100760, 100640, 100620, 100600, 100570, 100520, 100580, 100590, 
    100620, 100670, 100710, 100710, 100700, 100700, 100700, 100700, 100720, 
    100710, 100690, 100660, 100660, 100610, 100690, 100660, 100470, 100420, 
    100370, 100350, 100320, 100300, 100310, 100350, 100350, 100340, 100320, 
    100300, 100300, 100410, 100310, 100320, 100340, 100340, 100350, 100370, 
    100360, 100330, 100310, 100300, 100230, 100240, 100170, 100140, 100190, 
    100200, 100200, 100210, 100220, 100230, 100270, 100280, 100320, 100360, 
    100400, 100410, 100480, 100500, 100520, 100530, 100540, 100540, 100540, 
    100480, 100420, 100360, 100310, 100230, 100160, 100110, 100060, 100010, 
    100000, 99940, 99910, 99880, 99840, 99820, 99780, 99750, 99840, 99700, 
    99660, 99620, 99580, 99530, 99500, 99480, 99460, 99420, 99400, 99530, 
    99380, 99370, 99350, 99350, 99350, 99350, 99380, 99410, 99410, 99430, 
    99620, 99660, 99660, 99540, 99580, 99640, 99680, 99730, 99780, 99830, 
    99900, 99950, 99990, 100020, 100090, 100170, 100250, 100320, 100370, 
    100430, 100460, 100510, 100540, 100550, 100600, 100620, 100670, 100720, 
    100760, 100810, 100830, 100920, 100930, 100950, 100860, 100860, 100860, 
    100850, 100830, 100860, 100890, 100900, 100930, 100940, 100960, 100970, 
    100980, 101010, 101010, 101010, 101030, 101050, 101060, 101080, 101090, 
    101130, 101160, 101180, 101210, 101210, 101240, 101280, 101320, 101370, 
    101420, 101480, 101540, 101550, 101590, 101610, 101640, 101660, 101680, 
    101680, 101710, 101730, 101750, 101780, 101790, 101800, 101800, 101820, 
    101820, 101810, 101810, 101820, 101840, 101840, 101860, 101870, 101870, 
    101850, 101860, 101830, 101790, 101750, 101730, 101690, 101680, 101640, 
    101630, 101620, 101570, 101530, 101500, 101460, 101430, 101400, 101360, 
    101340, 101330, 101330, 101310, 101280, 101250, 101250, 101220, 101190, 
    101170, 101120, 101070, 101030, 101000, 100970, 100950, 100910, 100880, 
    100840, 100790, 100750, 100700, 100670, 100620, 100600, 100570, 100520, 
    100510, 100490, 100480, 100460, 100430, 100380, 100360, 100360, 100370, 
    100350, 100340, 100340, 100340, 100320, 100300, 100290, 100280, 100260, 
    100260, 100250, 100240, 100230, 100260, 100270, 100280, 100280, 100300, 
    100290, 100310, 100330, 100340, 100350, 100370, 100390, 100450, 100500, 
    100540, 100570, 100600, 100620, 100620, 100620, 100640, 100660, 100690, 
    100690, 100660, 100680, 100670, 100670, 100650, 100630, 100610, 100600, 
    100570, 100540, 100530, 100510, 100470, 100420, 100390, 100340, 100280, 
    100250, 100190, 100140, 100100, 100040, 100010, 100000, 99970, 99980, 
    99990, 100010, 100010, 100000, 100020, 100040, 100050, 100110, 100180, 
    100220, 100290, 100360, 100420, 100470, 100540, 100630, 100660, 100710, 
    100750, 100760, 100810, 100830, 100870, 100900, 100920, 100970, 100970, 
    101010, 101000, 101000, 101020, 101020, 101000, 100990, 100980, 100950, 
    100910, 100860, 100770, 100690, 100660, 100630, 100570, 100490, 100460, 
    100430, 100350, 100290, 100240, 100190, 100130, 100070, 100000, 99900, 
    99770, 99650, 99550, 99460, 99350, 99290, 99200, 99090, 98980, 98860, 
    98770, 98700, 98610, 98550, 98460, 98400, 98420, 98430, 98420, 98540, 
    98630, 98700, 98740, 98820, 98890, 98950, 99010, 99020, 99050, 99150, 
    99220, 99300, 99390, 99460, 99520, 99590, 99700, 99780, 99850, 99920, 
    100040, 100100, 100130, 100200, 100250, 100300, 100300, 100300, 100330, 
    100350, 100370, 100390, 100370, 100380, 100420, 100440, 100460, 100490, 
    100500, 100510, 100530, 100550, 100560, 100600, 100630, 100670, 100720, 
    100770, 100830, 100900, 100940, 101000, 101050, 101090, 101130, 101160, 
    101180, 101160, 101160, 101180, 101190, 101210, 101200, 101210, 101210, 
    101230, 101260, 101300, 101340, 101370, 101440, 101500, 101550, 101610, 
    101630, 101660, 101670, 101710, 101750, 101770, 101810, 101850, 101880, 
    101900, 101950, 102010, 102040, 102050, 102080, 102120, 102160, 102210, 
    102260, 102320, 102380, 102440, 102490, 102520, 102550, 102570, 102610, 
    102640, 102670, 102700, 102690, 102710, 102710, 102750, 102770, 102780, 
    102790, 102750, 102790, 102770, 102800, 102830, 102840, 102860, 102900, 
    102940, 102990, 103020, 103030, 103030, 103050, 103070, 103070, 103080, 
    103120, 103150, 103180, 103200, 103240, 103260, 103270, 103280, 103280, 
    103270, 103280, 103270, 103280, 103280, 103250, 103210, 103200, 103190, 
    103130, 103070, 103020, 102980, 102900, 102840, 102760, 102660, 102550, 
    102450, 102340, 102190, 102060, 101900, 101710, 101530, 101340, 101180, 
    101100, 100950, 100770, 100700, 100580, 100580, 100560, 100570, 100540, 
    100530, 100590, 100710, 100760, 100800, 100890, 100940, 100980, 101040, 
    101140, 101190, 101220, 101270, 101350, 101390, 101430, 101510, 101550, 
    101550, 101540, 101550, 101560, 101540, 101480, 101480, 101470, 101460, 
    101420, 101400, 101370, 101320, 101260, 101140, 101020, 100960, 100860, 
    100750, 100620, 100490, 100350, 100240, 100130, 100060, 100020, 99960, 
    99960, 99970, 99980, 99980, 99990, 100010, 100030, 100080, 100080, 
    100110, 100110, 100110, 100110, 100120, 100110, 100110, 100110, 100150, 
    100190, 100170, 100210, 100250, 100280, 100300, 100340, 100330, 100390, 
    100420, 100450, 100510, 100540, 100580, 100630, 100620, 100650, 100660, 
    100640, 100670, 100640, 100620, 100620, 100650, 100680, 100700, 100740, 
    100840, 100910, 101020, 101130, 101240, 101340, 101480, 101580, 101680, 
    101770, 101870, 101910, 102000, 102050, 102120, 102110, 102140, 102160, 
    102120, 102140, 102090, 102070, 102000, 102020, 101990, 101900, 101850, 
    101790, 101700, 101610, 101570, 101560, 101540, 101500, 101440, 101430, 
    101370, 101340, 101260, 101180, 101120, 101050, 100990, 100910, 100880, 
    100800, 100780, 100820, 100800, 100900, 100960, 100970, 101000, 101050, 
    101070, 101120, 101140, 101170, 101200, 101260, 101280, 101300, 101310, 
    101320, 101280, 101280, 101260, 101230, 101170, 101140, 101130, 101110, 
    101140, 101090, 101060, 101040, 101120, 101090, 101110, 101140, 101170, 
    101200, 101180, 101170, 101160, 101130, 101120, 101080, 101030, 101040, 
    101050, 101010, 100990, 100990, 100980, 100930, 100920, 100850, 100840, 
    100740, 100620, 100520, 100420, 100330, 100210, 100080, 99960, 99850, 
    99810, 99910, 100030, 100110, 100220, 100330, 100500, 100640, 100610, 
    100680, 100760, 100860, 100880, 100900, 100920, 100940, 100950, 100920, 
    100880, 100860, 100810, 100800, 100820, 100810, 100790, 100790, 100750, 
    100760, 100750, 100760, 100770, 100780, 100780, 100790, 100820, 100880, 
    100900, 100890, 100870, 100910, 100910, 100920, 100920, 100900, 100920, 
    100930, 100920, 100910, 100920, 100930, 100930, 100920, 100880, 100850, 
    100780, 100750, 100740, 100750, 100680, 100660, 100610, 100540, 100530, 
    100470, 100390, 100290, 100220, 100200, 100170, 100130, 100110, 100070, 
    100080, 100060, 100010, 99920, 99840, 99770, 99690, 99630, 99580, 99560, 
    99550, 99480, 99380, 99320, 99280, 99220, 99180, 99180, 99230, 99280, 
    99310, 99390, 99480, 99550, 99640, 99710, 99750, 99770, 99790, 99800, 
    99800, 99770, 99740, 99690, 99670, 99630, 99590, 99600, 99700, 99810, 
    99940, 100110, 100240, 100420, 100610, 100820, 101070, 101310, 101520, 
    101700, 101860, 102010, 102110, 102230, 102320, 102400, 102460, 102540, 
    102610, 102700, 102730, 102810, 102820, 102870, 102880, 102880, 102900, 
    102940, 102980, 103010, 103030, 103030, 103050, 103080, 103080, 103110, 
    103100, 103090, 103100, 103100, 103120, 103120, 103140, 103140, 103130, 
    103120, 103110, 103110, 103090, 103070, 103060, 103000, 102970, 102910, 
    102870, 102820, 102780, 102740, 102710, 102680, 102650, 102600, 102540, 
    102510, 102480, 102470, 102460, 102440, 102420, 102410, 102370, 102340, 
    102300, 102230, 102210, 102200, 102150, 102160, 102220, 102190, 102120, 
    102120, 102090, 102030, 102000, 101960, 101890, 101830, 101800, 101810, 
    101810, 101770, 101770, 101730, 101670, 101600, 101560, 101530, 101480, 
    101420, 101370, 101350, 101330, 101310, 101280, 101310, 101230, 101150, 
    101150, 101120, 101060, 101070, 101050, 101030, 100990, 101000, 101050, 
    101040, 101020, 101050, 101060, 101090, 101100, 101150, 101090, 101110, 
    101170, 101240, 101310, 101360, 101400, 101440, 101550, 101610, 101650, 
    101720, 101720, 101720, 101770, 101780, 101780, 101780, 101780, 101780, 
    101770, 101770, 101730, 101700, 101660, 101630, 101600, 101560, 101540, 
    101510, 101460, 101410, 101330, 101270, 101170, 101080, 101000, 100930, 
    100790, 100710, 100650, 100530, 100380, 100260, 100140, 100030, 99890, 
    99800, 99650, 99530, 99420, 99320, 99240, 99130, 99060, 98970, 98900, 
    98770, 98670, 98580, 98490, 98470, 98350, 98250, 98220, 98170, 98110, 
    98020, 97970, 97890, 97840, 97790, 97730, 97630, 97580, 97540, 97470, 
    97420, 97390, 97340, 97310, 97250, 97170, 97160, 97160, 97130, 97200, 
    97220, 97230, 97260, 97330, 97370, 97430, 97520, 97530, 97640, 97680, 
    97790, 97880, 97980, 98050, 98150, 98220, 98300, 98330, 98330, 98370, 
    98430, 98520, 98520, 98550, 98580, 98630, 98690, 98740, 98750, 98730, 
    98790, 98790, 98810, 98820, 98800, 98830, 98870, 98890, 98900, 98910, 
    98900, 98890, 98900, 98880, 98880, 98850, 98850, 98850, 98850, 98870, 
    98880, 98890, 98890, 98890, 98890, 98900, 98930, 98930, 98940, 98980, 
    99020, 99020, 99030, 99050, 99060, 99050, 99050, 99030, 99030, 99040, 
    99050, 99070, 99130, 99170, 99230, 99270, 99270, 99290, 99290, 99290, 
    99310, 99340, 99340, 99350, 99380, 99380, 99350, 99330, 99320, 99290, 
    99210, 99170, 99120, 99080, 99010, 98990, 98930, 98850, 98770, 98650, 
    98580, 98480, 98410, 98280, 98140, 98000, 97870, 97850, 97810, 97790, 
    97690, 97650, 97600, 97530, 97530, 97500, 97490, 97480, 97480, 97480, 
    97490, 97500, 97520, 97520, 97510, 97500, 97530, 97530, 97510, 97520, 
    97520, 97530, 97510, 97500, 97510, 97490, 97460, 97450, 97460, 97480, 
    97480, 97470, 97460, 97500, 97550, 97580, 97650, 97710, 97800, 97870, 
    97940, 98000, 98050, 98100, 98170, 98230, 98290, 98340, 98360, 98370, 
    98400, 98420, 98420, 98440, 98480, 98520, 98540, 98580, 98660, 98710, 
    98750, 98760, 98790, 98820, 98830, 98820, 98840, 98820, 98810, 98810, 
    98820, 98820, 98790, 98780, 98770, 98770, 98730, 98710, 98700, 98690, 
    98700, 98670, 98660, 98650, 98630, 98610, 98590, 98590, 98560, 98520, 
    98500, 98460, 98440, 98400, 98390, 98350, 98340, 98340, 98340, 98320, 
    98340, 98320, 98320, 98310, 98310, 98320, 98320, 98300, 98290, 98280, 
    98280, 98290, 98310, 98300, 98340, 98360, 98400, 98440, 98480, 98520, 
    98580, 98650, 98700, 98730, 98750, 98780, 98810, 98850, 98870, 98930, 
    99030, 99120, 99180, 99230, 99270, 99330, 99350, 99390, 99440, 99520, 
    99540, 99590, 99650, 99670, 99720, 99750, 99750, 99800, 99810, 99820, 
    99850, 99870, 99870, 99900, 99900, 99920, 99890, 99880, 99870, 99820, 
    99800, 99790, 99730, 99690, 99660, 99640, 99580, 99570, 99530, 99470, 
    99390, 99360, 99300, 99260, 99210, 99180, 99160, 99180, 99230, 99320, 
    99370, 99410, 99420, 99420, 99440, 99460, 99490, 99500, 99470, 99450, 
    99470, 99470, 99480, 99510, 99550, 99560, 99590, 99610, 99630, 99650, 
    99690, 99730, 99810, 99860, 99940, 99950, 99980, 100010, 100070, 100100, 
    100140, 100180, 100220, 100230, 100290, 100330, 100350, 100400, 100430, 
    100470, 100490, 100500, 100530, 100520, 100540, 100570, 100600, 100600, 
    100640, 100620, 100630, 100630, 100630, 100660, 100660, 100670, 100650, 
    100630, 100630, 100640, 100630, 100620, 100620, 100630, 100600, 100600, 
    100580, 100560, 100550, 100570, 100600, 100610, 100590, 100560, 100550, 
    100530, 100540, 100540, 100560, 100560, 100550, 100560, 100580, 100550, 
    100540, 100530, 100570, 100550, 100580, 100580, 100570, 100590, 100590, 
    100590, 100630, 100650, 100670, 100640, 100640, 100650, 100660, 100650, 
    100670, 100660, 100680, 100700, 100710, 100720, 100740, 100730, 100750, 
    100750, 100750, 100750, 100740, 100730, 100730, 100770, 100780, 100820, 
    100830, 100850, 100870, 100880, 100890, 100910, 100920, 100930, 100940, 
    100950, 100950, 101010, 101050, 101060, 101100, 101130, 101160, 101190, 
    101200, 101210, 101210, 101270, 101300, 101360, 101400, 101420, 101480, 
    101510, 101540, 101590, 101600, 101630, 101640, 101660, 101670, 101710, 
    101750, 101750, 101740, 101770, 101800, 101790, 101820, 101870, 101860, 
    101860, 101900, 101940, 101940, 101980, 102010, 102030, 102050, 102080, 
    102090, 102100, 102120, 102140, 102170, 102200, 102220, 102230, 102250, 
    102280, 102270, 102290, 102300, 102300, 102280, 102280, 102290, 102290, 
    102290, 102270, 102230, 102190, 102170, 102140, 102140, 102110, 102070, 
    102030, 102010, 102000, 101960, 101910, 101860, 101810, 101780, 101720, 
    101630, 101540, 101490, 101410, 101330, 101280, 101240, 101200, 101150, 
    101070, 101020, 100960, 100910, 100830, 100780, 100700, 100630, 100580, 
    100500, 100400, 100310, 100250, 100170, 100090, 100010, 100000, 99910, 
    99890, 99940, 99980, 100020, 100050, 100070, 100050, 100040, 100080, 
    100120, 100080, 100070, 100050, 100040, 100050, 100050, 100020, 99970, 
    99930, 99810, 99720, 99600, 99520, 99310, 99160, 99000, 98900, 98800, 
    98710, 98530, 98410, 98220, 98110, 97960, 97880, 97780, 97750, 97680, 
    97640, 97620, 97620, 97670, 97730, 97780, 97850, 97870, 97880, 97910, 
    97970, 98090, 98170, 98250, 98290, 98360, 98380, 98440, 98490, 98530, 
    98560, 98580, 98600, 98640, 98650, 98660, 98670, 98670, 98660, 98660, 
    98650, 98620, 98580, 98580, 98580, 98580, 98580, 98560, 98520, 98490, 
    98450, 98430, 98390, 98360, 98310, 98280, 98260, 98220, 98190, 98160, 
    98130, 98090, 98080, 98070, 98030, 98010, 97960, 97940, 97930, 97940, 
    97940, 97930, 97920, 97910, 97890, 97890, 97910, 97930, 97920, 97950, 
    97980, 98020, 98100, 98180, 98240, 98310, 98380, 98460, 98530, 98640, 
    98750, 98850, 99000, 99120, 99250, 99340, 99430, 99540, 99640, 99760, 
    99850, 99930, 100020, 100070, 100140, 100240, 100330, 100410, 100480, 
    100550, 100620, 100700, 100780, 100840, 100910, 100970, 101040, 101120, 
    101190, 101240, 101290, 101340, 101400, 101440, 101480, 101520, 101560, 
    101610, 101660, 101700, 101740, 101790, 101840, 101860, 101880, 101930, 
    101930, 101950, 101950, 101970, 102010, 102040, 102020, 102040, 102030, 
    102050, 102040, 102040, 102020, 102040, 102000, 101950, 101960, 101920, 
    101870, 101840, 101820, 101740, 101680, 101610, 101500, 101420, 101290, 
    101170, 101100, 101020, 100920, 100820, 100740, 100650, 100530, 100420, 
    100310, 100250, 100160, 100080, 100050, 100000, 99930, 99870, 99820, 
    99760, 99720, 99670, 99640, 99580, 99540, 99510, 99490, 99440, 99440, 
    99430, 99370, 99340, 99270, 99180, 99100, 99080, 99050, 99050, 99070, 
    99110, 99160, 99250, 99330, 99360, 99410, 99430, 99490, 99530, 99560, 
    99610, 99620, 99600, 99630, 99660, 99650, 99640, 99670, 99690, 99670, 
    99680, 99690, 99680, 99670, 99610, 99540, 99540, 99540, 99510, 99470, 
    99450, 99450, 99410, 99520, 99590, 99640, 99680, 99760, 99790, 99820, 
    99910, 99970, 99990, 100010, 100050, 100100, 100180, 100210, 100290, 
    100340, 100390, 100450, 100470, 100510, 100550, 100570, 100590, 100620, 
    100640, 100640, 100650, 100620, 100630, 100610, 100590, 100580, 100550, 
    100540, 100540, 100540, 100520, 100530, 100540, 100550, 100580, 100560, 
    100560, 100590, 100600, 100600, 100610, 100620, 100680, 100710, 100730, 
    100760, 100780, 100820, 100840, 100860, 100880, 100900, 100920, 100960, 
    100970, 100990, 100990, 101000, 101030, 101050, 101060, 101080, 101080, 
    101060, 101030, 101030, 101020, 101030, 101030, 101040, 101030, 101000, 
    100970, 100930, 100900, 100870, 100860, 100820, 100800, 100780, 100730, 
    100700, 100650, 100590, 100540, 100500, 100430, 100370, 100340, 100300, 
    100260, 100260, 100290, 100330, 100350, 100390, 100470, 100490, 100540, 
    100530, 100530, 100500, 100500, 100490, 100500, 100510, 100530, 100550, 
    100530, 100530, 100520, 100510, 100500, 100460, 100440, 100470, 100530, 
    100510, 100520, 100540, 100550, 100560, 100590, 100590, 100590, 100580, 
    100580, 100580, 100600, 100600, 100610, 100610, 100620, 100630, 100620, 
    100620, 100600, 100580, 100590, 100570, 100580, 100570, 100550, 100550, 
    100550, 100540, 100550, 100570, 100580, 100600, 100660, 100710, 100750, 
    100800, 100850, 100880, 100930, 100940, 100960, 100970, 100980, 100980, 
    101000, 101040, 101060, 101090, 101110, 101120, 101110, 101090, 101110, 
    101110, 101090, 101100, 101130, 101090, 101110, 101130, 101150, 101170, 
    101190, 101200, 101230, 101250, 101240, 101260, 101290, 101330, 101370, 
    101410, 101440, 101470, 101500, 101520, 101530, 101560, 101580, 101610, 
    101620, 101650, 101700, 101750, 101790, 101800, 101810, 101810, 101820, 
    101820, 101790, 101780, 101770, 101730, 101670, 101620, 101520, 101460, 
    101340, 101220, 101150, 101100, 101050, 101040, 101050, 101110, 101190, 
    101320, 101330, 101440, 101470, 101490, 101440, 101400, 101330, 101230, 
    101100, 100990, 100870, 100730, 100600, 100470, 100350, 100240, 100140, 
    100050, 100050, 100000, 100000, 100020, 100080, 100100, 100150, 100190, 
    100180, 100190, 100220, 100250, 100280, 100230, 100370, 100470, 100540, 
    100630, 100730, 100820, 100910, 100980, 101040, 101160, 101240, 101310, 
    101390, 101470, 101540, 101600, 101670, 101740, 101790, 101830, 101850, 
    101920, 101950, 101990, 102040, 102080, 102090, 102090, 102090, 102080, 
    102020, 101960, 101860, 101750, 101620, 101530, 101390, 101220, 101040, 
    100860, 100760, 100700, 100610, 100570, 100510, 100410, 100350, 100260, 
    100200, 100240, 100250, 100300, 100300, 100310, 100270, 100240, 100210, 
    100230, 100210, 100240, 100240, 100180, 100180, 100200, 100170, 100170, 
    100170, 100160, 100200, 100190, 100200, 100240, 100260, 100270, 100280, 
    100300, 100340, 100380, 100260, 100250, 100260, 100290, 100300, 100290, 
    100270, 100260, 100260, 100220, 100220, 100210, 100170, 100130, 100110, 
    100090, 100090, 100100, 100100, 100110, 100120, 100140, 100190, 100220, 
    100230, 100220, 100260, 100290, 100330, 100340, 100390, 100430, 100450, 
    100490, 100520, 100550, 100580, 100600, 100620, 100630, 100670, 100690, 
    100730, 100770, 100820, 100850, 100870, 100910, 100910, 100940, 100940, 
    100940, 100900, 100920, 100910, 100910, 100890, 100870, 100880, 100820, 
    100820, 100800, 100760, 100740, 100750, 100710, 100690, 100710, 100670, 
    100700, 100700, 100710, 100680, 100710, 100720, 100760, 100810, 100840, 
    100830, 100860, 100890, 100890, 100920, 100970, 100950, 101000, 100990, 
    100980, 101010, 101030, 101060, 101080, 101110, 101170, 101220, 101210, 
    101220, 101250, 101260, 101330, 101330, 101340, 101330, 101310, 101310, 
    101370, 101390, 101390, 101380, 101380, 101410, 101430, 101460, 101460, 
    101470, 101530, 101560, 101590, 101620, 101630, 101630, 101640, 101640, 
    101660, 101630, 101570, 101530, 101520, 101510, 101460, 101470, 101470, 
    101430, 101390, 101360, 101320, 101320, 101310, 101290, 101290, 101320, 
    101350, 101380, 101370, 101390, 101410, 101410, 101420, 101450, 101450, 
    101470, 101470, 101490, 101530, 101550, 101560, 101570, 101620, 101620, 
    101630, 101660, 101670, 101680, 101730, 101780, 101790, 101780, 101830, 
    101800, 101790, 101800, 101820, 101820, 101810, 101800, 101790, 101800, 
    101820, 101840, 101850, 101830, 101840, 101840, 101840, 101840, 101850, 
    101850, 101870, 101900, 101930, 101950, 101970, 101990, 102010, 102020, 
    102030, 102060, 102060, 102090, 102090, 102130, 102150, 102190, 102180, 
    102170, 102170, 102160, 102150, 102150, 102130, 102150, 102180, 102180, 
    102220, 102230, 102260, 102270, 102270, 102290, 102280, 102310, 102360, 
    102350, 102380, 102380, 102380, 102410, 102440, 102430, 102430, 102440, 
    102440, 102450, 102480, 102510, 102560, 102590, 102630, 102650, 102640, 
    102630, 102650, 102670, 102700, 102700, 102690, 102680, 102620, 102630, 
    102610, 102570, 102530, 102490, 102470, 102410, 102390, 102250, 102220, 
    102160, 102100, 102040, 101990, 101930, 101860, 101780, 101700, 101620, 
    101580, 101520, 101480, 101390, 101300, 101260, 101220, 101160, 101100, 
    101000, 100930, 100860, 100820, 100730, 100690, 100630, 100570, 100510, 
    100440, 100360, 100240, 100130, 100000, 99870, 99710, 99550, 99400, 
    99200, 99010, 98870, 98710, 98520, 98370, 98180, 97970, 97740, 97510, 
    97290, 97100, 96920, 96750, 96640, 96590, 96570, 96620, 96680, 96730, 
    96750, 96780, 96870, 96970, 97100, 97260, 97500, 97670, 97860, 98070, 
    98230, 98380, 98500, 98600, 98690, 98750, 98770, 98820, 98870, 98900, 
    98930, 99120, 99140, 99000, 99020, 99010, 99010, 99010, 98970, 98990, 
    98980, 98960, 98930, 98920, 98810, 98760, 98750, 98720, 98690, 98660, 
    98640, 98640, 98640, 98640, 98630, 98610, 98620, 98630, 98650, 98700, 
    98750, 98730, 98760, 98810, 98870, 98920, 99000, 99050, 99100, 99120, 
    99100, 99100, 99120, 99140, 99180, 99220, 99220, 99250, 99250, 99250, 
    99260, 99270, 99310, 99310, 99300, 99280, 99300, 99310, 99330, 99350, 
    99390, 99400, 99370, 99310, 99290, 99250, 99210, 99280, 99140, 99100, 
    99000, 98940, 98890, 98810, 98740, 98650, 98560, 98460, 98410, 98400, 
    98360, 98300, 98240, 98230, 98260, 98280, 98290, 98290, 98310, 98340, 
    98360, 98370, 98400, 98440, 98500, 98580, 98650, 98680, 98730, 98740, 
    98740, 98780, 98810, 98830, 98810, 98830, 98830, 98850, 98880, 98880, 
    98870, 98850, 98840, 98820, 98790, 98810, 98810, 98790, 98750, 98720, 
    98720, 98700, 98670, 98660, 98630, 98600, 98580, 98550, 98580, 98570, 
    98580, 98590, 98600, 98590, 98580, 98600, 98620, 98630, 98650, 98670, 
    98660, 98680, 98740, 98770, 98820, 98850, 98850, 98890, 98930, 98980, 
    99020, 99060, 99080, 99120, 99160, 99190, 99220, 99260, 99280, 99310, 
    99340, 99380, 99390, 99430, 99470, 99510, 99590, 99660, 99730, 99780, 
    99860, 99930, 100010, 100080, 100160, 100210, 100270, 100360, 100470, 
    100560, 100630, 100710, 100740, 100790, 100820, 100870, 100890, 100900, 
    100930, 100940, 101010, 101030, 101040, 101090, 101140, 101180, 101210, 
    101280, 101360, 101390, 101470, 101520, 101600, 101640, 101700, 101720, 
    101750, 101790, 101780, 101740, 101740, 101650, 101530, 101400, 101270, 
    101070, 100860, 100690, 100440, 100210, 99960, 99680, 99420, 99170, 
    98890, 98690, 98530, 98450, 98390, 98370, 98370, 98340, 98310, 98280, 
    98280, 98250, 98230, 98190, 98150, 98140, 98130, 98110, 98140, 98160, 
    98170, 98150, 98070, 98040, 97990, 98070, 98090, 98170, 98320, 98380, 
    98450, 98450, 98470, 98470, 98430, 98420, 98380, 98360, 98390, 98340, 
    98330, 98290, 98240, 98160, 98110, 98020, 98040, 98020, 98040, 98080, 
    98130, 98210, 98240, 98250, 98270, 98300, 98320, 98350, 98400, 98420, 
    98490, 98510, 98550, 98620, 98660, 98700, 98780, 98820, 98870, 98900, 
    98930, 98940, 98940, 98960, 98990, 99030, 99060, 99080, 99110, 99110, 
    99100, 99110, 99120, 99130, 99150, 99180, 99170, 99200, 99240, 99300, 
    99330, 99290, 99300, 99330, 99320, 99320, 99300, 99320, 99340, 99360, 
    99340, 99340, 99350, 99350, 99340, 99340, 99380, 99380, 99400, 99390, 
    99430, 99460, 99480, 99480, 99470, 99460, 99450, 99420, 99370, 99340, 
    99320, 99310, 99300, 99280, 99260, 99250, 99230, 99200, 99170, 99150, 
    99130, 99130, 99130, 99110, 99090, 99110, 99120, 99090, 99080, 99070, 
    99050, 99050, 99040, 99030, 99010, 98990, 99000, 99000, 98980, 98940, 
    98910, 98880, 98870, 98840, 98810, 98810, 98800, 98780, 98790, 98790, 
    98780, 98810, 98840, 98840, 98820, 98840, 98880, 98900, 98950, 98990, 
    99020, 99070, 99120, 99130, 99190, 99240, 99270, 99300, 99380, 99450, 
    99480, 99550, 99600, 99660, 99730, 99770, 99820, 99840, 99870, 99900, 
    99920, 99970, 100010, 100050, 100100, 100160, 100190, 100230, 100240, 
    100260, 100290, 100320, 100330, 100340, 100360, 100400, 100430, 100440, 
    100480, 100450, 100450, 100440, 100380, 100410, 100380, 100370, 100380, 
    100320, 100290, 100280, 100260, 100220, 100110, 100010, 99870, 99830, 
    99770, 99700, 99680, 99690, 99660, 99640, 99640, 99590, 99540, 99510, 
    99510, 99500, 99490, 99470, 99510, 99560, 99590, 99620, 99660, 99750, 
    99800, 99870, 99930, 100000, 100050, 100110, 100160, 100250, 100320, 
    100410, 100520, 100610, 100690, 100760, 100830, 100900, 100970, 101020, 
    101110, 101140, 101190, 101270, 101320, 101370, 101380, 101410, 101420, 
    101390, 101380, 101370, 101380, 101380, 101360, 101370, 101410, 101340, 
    101220, 101200, 101240, 101190, 101110, 101100, 101020, 100980, 100920, 
    100850, 100820, 100760, 100700, 100690, 100640, 100550, 100510, 100470, 
    100410, 100380, 100380, 100360, 100370, 100320, 100300, 100290, 100250, 
    100210, 100190, 100170, 100130, 100070, 100080, 100020, 100010, 99970, 
    99890, 99870, 99880, 99840, 99790, 99720, 99680, 99670, 99670, 99670, 
    99640, 99630, 99590, 99610, 99580, 99570, 99550, 99570, 99510, 99480, 
    99500, 99540, 99580, 99590, 99590, 99620, 99610, 99610, 99610, 99600, 
    99600, 99590, 99630, 99650, 99690, 99690, 99660, 99670, 99640, 99600, 
    99600, 99550, 99520, 99480, 99400, 99430, 99340, 99300, 99250, 99200, 
    99150, 99110, 99090, 99100, 99100, 99130, 99170, 99220, 99240, 99310, 
    99340, 99380, 99420, 99440, 99500, 99570, 99640, 99710, 99790, 99840, 
    99880, 99930, 99980, 100120, 100170, 100210, 100240, 100270, 100340, 
    100380, 100390, 100400, 100410, 100410, 100390, 100390, 100400, 100390, 
    100350, 100310, 100350, 100310, 100270, 100230, 100200, 100170, 100080, 
    100040, 99990, 99930, 99900, 99870, 99880, 99860, 99840, 99820, 99830, 
    99880, 99880, 99870, 99910, 99920, 99920, 99940, 99920, 99900, 99900, 
    99880, 99830, 99760, 99660, 99580, 99540, 99460, 99360, 99290, 99180, 
    99130, 99060, 98970, 98930, 98870, 98760, 98700, 98640, 98580, 98530, 
    98500, 98510, 98450, 98410, 98360, 98320, 98290, 98250, 98210, 98170, 
    98110, 98060, 97980, 97950, 97910, 97890, 97840, 97780, 97690, 97520, 
    97380, 97250, 97110, 96900, 96700, 96970, 96780, 96660, 96520, 96350, 
    96200, 96080, 95960, 95840, 95710, 95600, 95500, 95380, 95280, 95220, 
    95200, 95180, 95180, 95210, 95260, 95310, 95310, 95300, 95290, 95530, 
    95520, 95520, 95510, 95530, 95540, 95560, 95590, 95630, 95650, 95690, 
    95720, 95910, 95960, 96020, 96080, 96170, 96230, 96300, 96390, 96480, 
    96560, 96650, 96750, 96880, 96950, 97030, 97130, 97200, 97290, 97380, 
    97450, 97530, 97590, 97640, 97710, 97770, 97850, 97910, 98090, 98180, 
    98240, 98340, 98450, 98550, 98630, 98700, 98650, 98720, 98820, 98920, 
    99030, 99110, 99170, 99260, 99350, 99430, 99490, 99570, 99530, 99610, 
    99680, 99780, 99880, 99970, 100040, 100110, 100180, 100220, 100260, 
    100250, 100290, 100310, 100360, 100390, 100360, 100370, 100350, 100320, 
    100310, 100260, 100220, 100160, 100200, 100090, 100030, 99960, 99840, 
    99640, 99450, 99300, 99120, 98910, 98740, 98620, 98630, 98600, 98650, 
    98770, 98930, 99090, 99270, 99450, 99640, 99870, 99940, 100180, 100240, 
    100330, 100470, 100530, 100530, 100510, 100470, 100370, 100280, 100200, 
    100150, 100080, 100060, 100040, 100010, 100010, 100060, 100130, 100240, 
    100380, 100590, 100810, 100960, 101140, 101460, 101580, 101670, 101840, 
    101910, 101930, 101950, 102010, 101990, 101980, 101870, 101810, 101690, 
    101530, 101360, 101200, 101000, 100820, 100630, 100440, 100210, 100050, 
    99860, 99760, 99680, 99610, 99580, 99540, 99490, 99420, 99330, 99120, 
    98840, 98570, 98200, 97950, 97780, 98080, 98170, 98150, 98190, 98280, 
    98470, 98680, 98930, 99240, 99690, 100010, 100230, 100500, 100720, 
    100950, 101150, 101290, 101470, 101520, 101560, 101650, 101620, 101590, 
    101450, 101510, 101510, 101470, 101460, 101440, 101420, 101410, 101370, 
    101370, 101390, 101400, 101360, 101430, 101490, 101530, 101590, 101660, 
    101680, 101710, 101690, 101690, 101700, 101700, 101730, 101770, 101800, 
    101830, 101850, 101900, 102010, 101910, 101910, 101920, 101910, 101930, 
    101930, 101930, 101930, 101960, 101950, 101930, 101890, 101880, 101870, 
    101840, 101810, 101790, 101800, 101830, 101860, 101880, 101920, 101940, 
    101950, 101970, 101970, 101990, 102180, 102190, 102050, 102090, 102120, 
    102170, 102220, 102250, 102250, 102270, 102290, 102290, 102310, 102360, 
    102360, 102330, 102350, 102370, 102390, 102380, 102390, 102520, 102420, 
    102440, 102390, 102430, 102450, 102470, 102490, 102570, 102590, 102570, 
    102550, 102540, 102550, 102500, 102490, 102470, 102480, 102450, 102430, 
    102420, 102390, 102430, 102410, 102300, 102280, 102250, 102200, 102170, 
    102160, 102130, 102120, 102080, 102070, 102010, 101960, 101890, 101810, 
    101780, 101700, 101640, 101550, 101490, 101450, 101550, 101280, 101460, 
    101140, 101110, 101060, 100990, 101220, 101180, 100880, 100870, 101130, 
    101110, 101100, 100870, 100880, 100890, 100920, 100930, 100940, 100940, 
    101180, 101000, 101020, 101220, 101090, 101130, 101170, 101350, 101220, 
    101220, 101410, 101290, 101330, 101540, 101400, 101590, 101480, 101510, 
    101530, 101550, 101580, 101630, 101650, 101660, 101630, 101760, 101680, 
    101720, 101730, 101810, 101720, 101730, 101730, 101730, 101730, 101740, 
    101710, 101690, 101690, 101690, 101670, 101670, 101670, 101680, 101650, 
    101640, 101630, 101600, 101590, 101580, 101570, 101570, 101550, 101520, 
    101450, 101460, 101440, 101430, 101430, 101460, 101400, 101360, 101300, 
    101250, 101210, 101180, 101120, 101010, 100930, 100830, 100790, 100720, 
    100650, 100590, 100530, 100650, 100490, 100440, 100340, 100250, 100170, 
    100100, 100090, 100090, 100050, 100020, 99960, 99920, 99940, 99960, 
    99990, 100010, 100020, 100080, 100110, 100140, 100140, 100190, 100150, 
    100180, 100120, 100040, 100010, 99950, 99900, 99830, 99790, 99750, 99710, 
    99660, 99620, 99450, 99410, 99330, 99230, 99160, 99100, 99080, 99050, 
    99000, 98960, 98940, 98930, 98920, 98910, 98900, 98900, 99000, 98890, 
    98910, 98930, 98940, 98970, 98990, 99010, 99030, 99060, 99080, 99150, 
    99210, 99260, 99320, 99370, 99430, 99490, 99540, 99580, 99610, 99620, 
    99660, 99660, 99650, 99680, 99720, 99740, 99850, 99900, 99920, 99910, 
    99900, 99900, 99890, 99850, 99830, 100050, 100020, 100070, 100100, 
    100090, 100090, 100050, 100010, 99980, 99910, 99820, 99820, 99910, 99840, 
    99800, 99750, 99700, 99680, 99630, 99590, 99490, 99470, 99430, 99420, 
    99370, 99320, 99220, 99210, 99250, 99180, 99200, 99260, 99160, 99140, 
    99380, 99390, 99340, 99300, 99440, 99430, 99530, 99500, 99560, 99580, 
    99700, 99750, 99760, 99840, 99890, 99910, 99950, 100000, 100050, 100080, 
    100140, 100240, 100180, 100200, 100200, 100230, 100260, 100290, 100300, 
    100280, 100290, 100280, 100260, 100230, 100210, 100240, 100230, 100180, 
    100140, 100140, 100150, 100200, 100180, 100100, 100140, 100160, 100180, 
    100220, 100230, 100230, 100290, 100280, 100360, 100420, 100500, 100530, 
    100600, 100670, 100700, 100790, 100870, 100940, 101040, 101100, 101190, 
    101260, 101330, 101360, 101480, 101530, 101590, 101630, 101710, 101710, 
    101770, 101860, 101880, 101940, 101970, 102000, 102000, 102010, 102030, 
    102070, 102110, 102140, 102170, 102170, 102200, 102240, 102270, 102310, 
    102340, 102380, 102420, 102440, 102440, 102440, 102460, 102460, 102480, 
    102500, 102540, 102600, 102620, 102630, 102640, 102630, 102650, 102650, 
    102690, 102700, 102720, 102700, 102770, 102680, 102660, 102760, 102590, 
    102560, 102580, 102590, 102600, 102540, 102510, 102470, 102460, 102400, 
    102340, 102320, 102260, 102240, 102190, 102100, 102080, 102060, 101970, 
    101910, 101780, 101820, 101600, 101510, 101410, 101320, 101230, 101160, 
    101250, 100990, 100940, 100860, 100770, 100680, 100610, 100540, 100420, 
    100350, 100260, 100200, 100170, 100110, 100040, 99970, 99900, 99840, 
    99790, 99890, 99680, 99640, 99710, 99570, 99530, 99480, 99440, 99360, 
    99260, 99200, 99110, 99050, 98970, 98940, 98900, 98870, 98830, 98810, 
    98790, 98760, 98820, 98800, 98810, 98870, 98840, 98850, 98900, 98960, 
    99020, 99060, 99120, 99180, 99230, 99290, 99340, 99380, 99430, 99480, 
    99540, 99570, 99600, 99620, 99630, 99660, 99650, 99740, 99770, 99680, 
    99710, 99710, 99700, 99700, 99810, 99690, 99690, 99680, 99690, 99700, 
    99720, 99730, 99730, 99710, 99690, 99680, 99660, 99660, 99650, 99640, 
    99590, 99540, 99500, 99460, 99410, 99360, 99350, 99290, 99220, 99210, 
    99180, 99170, 99170, 99180, 99170, 99190, 99210, 99220, 99250, 99280, 
    99310, 99350, 99410, 99460, 99500, 99540, 99690, 99730, 99770, 99780, 
    99830, 99870, 99910, 99950, 100000, 100020, 100090, 100110, 100140, 
    100140, 100140, 100170, 100170, 100220, 100240, 100230, 100250, 100260, 
    100250, 100260, 100250, 100250, 100250, 100240, 100260, 100250, 100260, 
    100270, 100240, 100250, 100250, 100220, 100210, 100190, 100170, 100170, 
    100170, 100140, 100110, 100070, 100060, 100030, 100010, 99960, 99940, 
    99920, 99900, 99890, 99830, 99820, 99780, 99730, 99720, 99630, 99580, 
    99520, 99490, 99480, 99470, 99480, 99490, 99670, 99710, 99780, 99850, 
    99930, 99990, 100030, 100080, 100120, 100160, 100190, 100230, 100250, 
    100270, 100310, 100320, 100340, 100360, 100360, 100370, 100370, 100360, 
    100380, 100380, 100360, 100340, 100350, 100340, 100300, 100280, 100270, 
    99990, 99950, 99910, 99870, 99800, 99740, 99650, 99570, 99460, 99370, 
    99400, 99380, 99420, 99470, 99560, 99630, 99720, 99860, 100010, 100130, 
    100270, 100420, 100540, 100650, 100770, 100840, 100860, 100910, 100960, 
    101020, 101070, 101070, 101040, 100940, 100820, 100770, 100660, 100530, 
    100370, 100250, 100150, 100080, 100010, 99900, 99810, 99710, 99610, 
    99540, 99470, 99410, 99360, 99320, 99330, 99320, 99360, 99400, 99430, 
    99500, 99590, 99680, 99760, 99840, 99920, 99970, 100050, 100130, 100200, 
    100280, 100350, 100400, 100480, 100570, 100620, 100700, 100730, 100770, 
    100790, 100810, 100820, 100830, 100830, 100800, 100760, 100750, 100730, 
    100720, 100680, 100650, 100670, 100690, 100720, 100750, 100770, 100830, 
    100870, 100900, 100950, 101000, 101080, 101120, 101150, 101200, 101250, 
    101260, 101320, 101310, 101290, 101320, 101320, 101330, 101300, 101320, 
    101310, 101280, 101250, 101200, 101140, 101010, 100850, 100780, 100680, 
    100610, 100550, 100500, 100450, 100400, 100340, 100330, 100360, 100340, 
    100320, 100340, 100340, 100320, 100310, 100320, 100330, 100340, 100390, 
    100380, 100380, 100340, 100320, 100310, 100270, 100280, 100240, 100240, 
    100260, 100200, 100200, 100220, 100330, 100380, 100440, 100460, 100490, 
    100720, 100830, 100900, 100990, 101030, 101110, 101200, 101300, 101390, 
    101520, 101830, 101940, 102050, 102110, 102210, 102430, 102500, 102600, 
    102630, 102690, 102740, 102750, 102730, 102690, 102660, 102610, 102570, 
    102520, 102490, 102460, 102420, 102440, 102390, 102420, 102380, 102340, 
    102260, 102200, 102020, 101980, 101920, 101890, 101820, 101860, 101870, 
    101910, 101950, 102010, 102020, 102000, 101980, 101920, 101970, 101970, 
    101970, 101970, 101990, 101960, 101960, 101960, 101930, 101870, 101840, 
    101840, 101790, 101810, 101780, 101740, 101670, 101700, 101700, 101680, 
    101710, 101720, 101700, 101680, 101650, 101670, 101670, 101710, 101700, 
    101710, 101720, 101720, 101730, 101740, 101740, 101740, 101750, 101770, 
    101790, 101820, 101830, 101800, 101830, 101850, 101880, 101890, 101900, 
    101910, 101880, 101870, 101870, 101880, 101870, 101840, 101830, 101820, 
    101810, 101820, 101810, 101820, 101820, 101820, 101810, 101820, 101820, 
    101840, 101860, 101890, 101900, 101910, 101900, 101900, 101900, 101890, 
    101900, 101930, 101940, 101950, 101890, 101910, 101910, 101910, 101900, 
    101890, 101890, 101890, 101870, 101870, 101850, 101860, 101850, 101860, 
    101850, 101860, 101860, 101840, 101830, 101810, 101810, 101810, 101800, 
    101790, 101770, 101750, 101740, 101720, 101710, 101680, 101650, 101630, 
    101610, 101540, 101230, 101260, 101260, 101250, 101260, 101280, 101300, 
    101310, 101330, 101330, 101340, 101360, 101370, 101400, 101410, 101440, 
    101450, 101460, 101490, 101510, 101530, 101570, 101610, 101630, 101670, 
    101700, 101710, 101720, 101730, 101710, 101700, 101700, 101690, 101680, 
    101650, 101630, 101620, 101650, 101650, 101650, 101640, 101660, 101660, 
    101660, 101670, 101630, 101630, 101640, 101660, 101620, 101620, 101620, 
    101620, 101620, 101620, 101610, 101610, 101610, 101560, 101540, 101540, 
    101540, 101530, 101520, 101490, 101470, 101460, 101460, 101450, 101440, 
    101440, 101440, 101430, 101420, 101440, 101470, 101470, 101480, 101480, 
    101510, 101520, 101540, 101560, 101600, 101600, 101610, 101640, 101660, 
    101660, 101690, 101730, 101750, 101740, 101760, 101790, 101820, 101860, 
    101890, 101910, 101900, 101910, 101920, 101940, 101970, 101970, 101980, 
    101970, 101950, 101950, 101930, 101920, 101910, 101920, 101900, 101900, 
    101880, 101850, 101830, 101820, 101800, 101790, 101710, 101670, 101640, 
    101620, 101610, 101590, 101560, 101530, 101510, 101470, 101440, 101420, 
    101390, 101370, 101340, 101330, 101310, 101280, 101270, 101250, 101210, 
    101150, 101120, 101070, 101030, 101000, 100970, 100940, 100910, 100880, 
    100850, 100740, 100710, 100690, 100680, 100660, 100660, 100650, 100650, 
    100640, 100630, 100620, 100620, 100610, 100570, 100560, 100550, 100580, 
    100590, 100600, 100600, 100610, 100600, 100610, 100610, 100630, 100650, 
    100670, 100710, 100740, 100760, 100790, 100800, 100810, 100830, 100820, 
    100830, 100850, 100860, 100890, 100910, 100920, 100930, 100930, 100960, 
    100980, 100980, 100990, 101000, 101010, 101030, 101070, 101100, 101110, 
    101120, 101140, 101160, 101190, 101210, 101220, 101250, 101280, 101410, 
    101420, 101450, 101490, 101530, 101540, 101560, 101570, 101610, 101650, 
    101660, 101710, 101750, 101760, 101790, 101800, 101810, 101820, 101820, 
    101830, 101830, 101830, 101850, 101840, 101840, 101830, 101770, 101740, 
    101730, 101710, 101720, 101720, 101720, 101730, 101700, 101690, 101680, 
    101660, 101640, 101620, 101610, 101580, 101550, 101540, 101530, 101490, 
    101460, 101440, 101440, 101430, 101410, 101380, 101350, 101320, 101280, 
    101230, 101220, 101190, 101150, 101140, 101110, 101080, 101070, 101080, 
    101070, 101070, 101020, 101010, 101030, 101050, 101080, 101110, 101120, 
    101150, 101180, 101220, 101250, 101290, 101320, 101350, 101380, 101410, 
    101450, 101470, 101480, 101480, 101500, 101510, 101530, 101560, 101580, 
    101600, 101630, 101640, 101630, 101620, 101610, 101630, 101630, 101630, 
    101650, 101650, 101650, 101640, 101620, 101590, 101570, 101560, 101550, 
    101540, 101520, 101520, 101500, 101480, 101470, 101430, 101410, 101410, 
    101380, 101380, 101360, 101340, 101340, 101330, 101350, 101360, 101350, 
    101340, 101340, 101330, 101330, 101320, 101360, 101360, 101360, 101360, 
    101310, 101310, 101270, 101210, 101180, 101180, 101170, 101130, 101090, 
    101060, 101030, 100980, 100920, 100920, 100900, 100890, 100860, 100850, 
    100830, 100790, 100730, 100710, 100640, 100610, 100570, 100530, 100500, 
    100470, 100440, 100420, 100380, 100350, 100310, 100270, 100220, 100170, 
    100100, 100060, 100000, 99950, 99920, 99810, 99750, 99730, 99710, 99700, 
    99660, 99630, 99630, 99630, 99650, 99650, 99680, 99700, 99710, 99720, 
    99730, 99720, 99740, 99750, 99770, 99800, 99860, 99870, 99910, 99940, 
    99920, 99950, 99960, 99980, 99990, 100030, 100070, 100090, 100120, 
    100160, 100190, 100220, 100250, 100280, 100310, 100480, 100520, 100550, 
    100610, 100700, 100730, 100930, 100940, 100950, 100970, 101000, 101020, 
    101030, 101040, 101100, 101110, 101130, 101140, 101150, 101180, 101220, 
    101240, 101270, 101290, 101300, 101360, 101370, 101390, 101410, 101430, 
    101430, 101470, 101530, 101570, 101580, 101600, 101630, 101650, 101670, 
    101730, 101750, 101830, 101860, 101900, 101920, 101940, 101980, 102000, 
    102000, 102020, 102030, 102060, 102100, 102130, 102150, 102150, 102190, 
    102190, 102180, 102190, 102200, 102190, 102200, 102190, 102180, 102190, 
    102190, 102160, 102150, 102130, 102090, 102070, 102060, 102040, 102000, 
    101980, 101980, 101990, 101940, 101920, 101890, 101850, 101820, 101810, 
    101780, 101770, 101750, 101730, 101700, 101680, 101660, 101650, 101620, 
    101590, 101580, 101560, 101530, 101530, 101510, 101480, 101460, 101450, 
    101420, 101410, 101380, 101340, 101310, 101310, 101340, 101350, 101360, 
    101370, 101360, 101340, 101330, 101310, 101300, 101300, 101280, 101280, 
    101260, 101250, 101260, 101260, 101250, 101210, 101190, 101180, 101160, 
    101130, 101130, 101130, 101130, 101130, 101140, 101150, 101150, 101140, 
    101140, 101160, 101150, 101130, 101140, 101140, 101160, 101150, 101220, 
    101240, 101240, 101270, 101300, 101290, 101330, 101330, 101370, 101370, 
    101400, 101430, 101460, 101490, 101510, 101550, 101590, 101620, 101660, 
    101690, 101660, 101720, 101740, 101770, 101760, 101790, 101850, 101870, 
    101880, 101880, 101880, 101870, 101870, 101860, 101870, 101860, 101840, 
    101820, 101800, 101770, 101810, 101770, 101740, 101710, 101680, 101650, 
    101610, 101550, 101530, 101510, 101510, 101450, 101410, 101380, 101360, 
    101360, 101310, 101260, 101240, 101220, 101170, 101130, 101110, 101080, 
    101080, 101030, 100980, 100960, 100890, 100840, 100810, 100790, 100720, 
    100640, 100600, 100530, 100460, 100380, 100330, 100230, 100190, 100130, 
    100090, 100020, 99980, 99940, 99910, 99860, 99850, 99780, 99800, 99800, 
    99770, 99760, 99760, 99740, 99730, 99740, 99710, 99690, 99670, 99640, 
    99630, 99580, 99590, 99610, 99580, 99540, 99560, 99540, 99570, 99600, 
    99610, 99620, 99570, 99640, 99630, 99610, 99590, 99510, 99500, 99580, 
    99600, 99630, 99600, 99640, 99630, 99620, 99590, 99610, 99640, 99660, 
    99690, 99740, 99760, 99790, 99820, 99860, 99880, 99920, 99940, 99990, 
    100020, 100090, 100120, 100150, 100200, 100230, 100270, 100300, 100340, 
    100360, 100390, 100390, 100450, 100480, 100520, 100530, 100570, 100580, 
    100610, 100640, 100660, 100650, 100660, 100660, 100680, 100690, 100690, 
    100690, 100690, 100710, 100720, 100700, 100700, 100690, 100690, 100690, 
    100710, 100740, 100760, 100780, 100790, 100800, 100810, 100800, 100790, 
    100790, 100770, 100750, 100740, 100740, 100740, 100720, 100700, 100690, 
    100660, 100640, 100620, 100590, 100540, 100510, 100500, 100480, 100470, 
    100450, 100410, 100410, 100380, 100330, 100310, 100290, 100270, 100270, 
    100250, 100230, 100210, 100220, 100210, 100190, 100170, 100150, 100140, 
    100130, 100110, 100100, 100090, 100090, 100110, 100110, 100090, 100080, 
    100070, 100040, 100040, 100010, 100000, 99980, 99950, 99910, 99890, 
    99880, 99880, 99870, 99850, 99850, 99870, 99890, 99910, 99910, 99920, 
    99950, 99970, 100010, 100020, 100040, 100080, 100120, 100150, 100180, 
    100200, 100210, 100230, 100250, 100280, 100290, 100310, 100300, 100340, 
    100320, 100300, 100290, 100300, 100300, 100270, 100220, 100250, 100240, 
    100250, 100230, 100200, 100120, 100030, 99950, 99870, 99720, 99630, 
    99620, 99550, 99590, 99600, 99560, 99540, 99560, 99490, 99450, 99450, 
    99510, 99420, 99410, 99450, 99500, 99470, 99530, 99530, 99450, 99400, 
    99370, 99410, 99370, 99400, 99430, 99450, 99480, 99530, 99540, 99580, 
    99560, 99580, 99570, 99570, 99610, 99640, 99600, 99610, 99580, 99610, 
    99650, 99690, 99700, 99730, 99740, 99760, 99800, 99800, 99830, 99870, 
    99870, 99910, 99950, 99930, 99950, 99960, 99960, 100000, 100020, 100040, 
    100020, 100030, 100040, 100120, 100170, 100220, 100290, 100340, 100380, 
    100420, 100480, 100530, 100560, 100620, 100640, 100660, 100680, 100700, 
    100720, 100780, 100830, 100850, 100910, 100960, 100980, 101020, 101070, 
    101110, 101130, 101150, 101160, 101160, 101160, 101150, 101140, 101110, 
    101090, 101080, 101060, 101040, 101030, 101030, 101010, 100990, 100990, 
    100970, 100960, 100940, 100930, 100930, 100940, 100920, 100910, 100900, 
    100900, 100890, 100880, 100850, 100830, 100820, 100810, 100800, 100800, 
    100790, 100770, 100760, 100750, 100730, 100730, 100720, 100700, 100680, 
    100660, 100650, 100630, 100640, 100640, 100640, 100620, 100600, 100590, 
    100560, 100530, 100510, 100500, 100500, 100490, 100490, 100490, 100480, 
    100490, 100490, 100480, 100480, 100500, 100510, 100530, 100560, 100580, 
    100610, 100630, 100660, 100690, 100690, 100710, 100730, 100750, 100760, 
    100770, 100810, 100830, 100850, 100880, 100890, 100920, 100930, 100950, 
    100970, 100990, 101010, 101030, 101060, 101080, 101100, 101120, 101130, 
    101130, 101130, 101150, 101160, 101150, 101160, 101170, 101190, 101200, 
    101200, 101210, 101230, 101250, 101260, 101260, 101250, 101240, 101240, 
    101250, 101250, 101250, 101260, 101270, 101260, 101260, 101260, 101250, 
    101260, 101260, 101280, 101300, 101320, 101340, 101360, 101380, 101400, 
    101420, 101430, 101470, 101460, 101510, 101520, 101550, 101590, 101630, 
    101650, 101680, 101730, 101760, 101770, 101810, 101820, 101840, 101870, 
    101920, 101950, 102000, 102020, 102050, 102060, 102090, 102090, 102100, 
    102110, 102110, 102130, 102150, 102140, 102140, 102140, 102150, 102150, 
    102170, 102180, 102160, 102140, 102140, 102130, 102140, 102170, 102190, 
    102190, 102200, 102220, 102200, 102220, 102210, 102200, 102190, 102190, 
    102190, 102190, 102180, 102190, 102170, 102160, 102140, 102110, 102070, 
    102050, 102060, 102050, 102050, 102050, 102040, 102040, 102040, 102060, 
    102040, 102010, 102000, 101980, 101950, 101950, 101940, 101920, 101920, 
    101910, 101900, 101870, 101850, 101840, 101840, 101820, 101810, 101800, 
    101790, 101790, 101790, 101780, 101750, 101730, 101710, 101720, 101690, 
    101660, 101630, 101630, 101620, 101600, 101590, 101580, 101560, 101550, 
    101540, 101510, 101500, 101480, 101440, 101420, 101440, 101420, 101420, 
    101430, 101430, 101420, 101420, 101400, 101410, 101390, 101400, 101410, 
    101420, 101400, 101420, 101400, 101360, 101370, 101380, 101360, 101360, 
    101350, 101330, 101320, 101310, 101270, 101260, 101250, 101240, 101210, 
    101200, 101200, 101180, 101150, 101140, 101110, 101120, 101110, 101110, 
    101110, 101110, 101100, 101090, 101090, 101090, 101100, 101110, 101130, 
    101160, 101180, 101200, 101220, 101250, 101290, 101320, 101350, 101360, 
    101390, 101410, 101440, 101470, 101490, 101540, 101570, 101600, 101630, 
    101650, 101670, 101700, 101710, 101720, 101720, 101730, 101760, 101770, 
    101790, 101780, 101780, 101770, 101760, 101760, 101760, 101750, 101750, 
    101770, 101760, 101780, 101780, 101790, 101800, 101800, 101790, 101780, 
    101760, 101750, 101730, 101720, 101710, 101720, 101740, 101740, 101710, 
    101680, 101670, 101680, 101670, 101690, 101690, 101700, 101740, 101780, 
    101800, 101810, 101820, 101850, 101850, 101880, 101880, 101890, 101890, 
    101890, 101890, 101910, 101940, 101940, 101950, 101970, 101980, 101980, 
    101980, 101990, 102000, 102030, 102020, 102030, 102040, 102050, 102030, 
    102000, 101980, 101950, 101900, 101860, 101850, 101850, 101820, 101800, 
    101780, 101760, 101730, 101720, 101680, 101650, 101620, 101590, 101560, 
    101540, 101540, 101520, 101500, 101500, 101460, 101430, 101430, 101410, 
    101420, 101410, 101420, 101440, 101470, 101470, 101500, 101520, 101520, 
    101530, 101530, 101560, 101580, 101610, 101610, 101660, 101680, 101720, 
    101750, 101780, 101800, 101820, 101870, 101900, 101900, 101910, 101940, 
    101970, 102010, 102030, 102060, 102060, 102080, 102070, 102080, 102070, 
    102070, 102070, 102070, 102090, 102110, 102150, 102150, 102170, 102190, 
    102190, 102210, 102230, 102250, 102260, 102280, 102280, 102290, 102300, 
    102300, 102310, 102330, 102360, 102370, 102370, 102390, 102390, 102430, 
    102450, 102480, 102510, 102530, 102540, 102560, 102580, 102580, 102610, 
    102630, 102630, 102650, 102640, 102650, 102660, 102660, 102660, 102670, 
    102680, 102700, 102690, 102660, 102660, 102650, 102630, 102610, 102600, 
    102580, 102600, 102590, 102560, 102510, 102510, 102490, 102490, 102430, 
    102420, 102410, 102410, 102400, 102390, 102350, 102340, 102330, 102270, 
    102240, 102200, 102130, 102080, 102030, 102000, 101970, 101950, 101940, 
    101930, 101890, 101900, 101880, 101870, 101880, 101850, 101890, 101890, 
    101900, 101930, 101940, 101950, 101970, 102000, 102010, 102020, 102070, 
    102080, 102080, 102140, 102180, 102180, 102220, 102250, 102260, 102250, 
    102260, 102240, 102250, 102260, 102260, 102270, 102260, 102270, 102270, 
    102270, 102290, 102280, 102270, 102290, 102300, 102310, 102300, 102300, 
    102280, 102280, 102270, 102260, 102260, 102250, 102260, 102240, 102240, 
    102210, 102230, 102210, 102210, 102230, 102210, 102200, 102210, 102200, 
    102180, 102170, 102140, 102150, 102160, 102180, 102170, 102140, 102130, 
    102120, 102110, 102090, 102080, 102080, 102080, 102090, 102110, 102100, 
    102120, 102130, 102130, 102110, 102090, 102100, 102130, 102170, 102180, 
    102190, 102200, 102210, 102220, 102220, 102240, 102250, 102250, 102240, 
    102260, 102280, 102300, 102320, 102340, 102350, 102360, 102360, 102370, 
    102370, 102360, 102360, 102370, 102360, 102360, 102360, 102380, 102380, 
    102360, 102350, 102340, 102330, 102330, 102330, 102320, 102320, 102320, 
    102300, 102280, 102260, 102250, 102240, 102230, 102220, 102190, 102160, 
    102130, 102110, 102080, 102060, 102050, 102030, 102000, 101980, 101960, 
    101930, 101890, 101870, 101850, 101810, 101780, 101750, 101740, 101720, 
    101690, 101660, 101630, 101600, 101590, 101560, 101530, 101520, 101490, 
    101470, 101440, 101430, 101420, 101420, 101410, 101410, 101400, 101380, 
    101380, 101350, 101340, 101330, 101330, 101340, 101340, 101330, 101320, 
    101310, 101290, 101250, 101210, 101190, 101140, 101160, 101160, 101150, 
    101120, 101090, 101060, 101040, 101000, 100910, 100830, 100760, 100730, 
    100720, 100710, 100750, 100720, 100820, 100840, 100890, 100900, 100930, 
    100910, 100950, 100940, 100980, 100950, 100950, 100920, 100960, 101040, 
    101050, 101090, 101070, 101100, 101110, 101140, 101200, 101210, 101250, 
    101250, 101270, 101280, 101260, 101280, 101300, 101310, 101340, 101360, 
    101380, 101390, 101400, 101390, 101400, 101390, 101390, 101390, 101390, 
    101390, 101400, 101420, 101440, 101450, 101460, 101480, 101480, 101500, 
    101520, 101530, 101510, 101480, 101480, 101440, 101420, 101390, 101380, 
    101370, 101370, 101380, 101370, 101400, 101390, 101380, 101360, 101390, 
    101400, 101400, 101400, 101430, 101440, 101460, 101480, 101490, 101490, 
    101490, 101480, 101480, 101500, 101540, 101550, 101560, 101580, 101600, 
    101600, 101630, 101610, 101610, 101620, 101630, 101640, 101630, 101640, 
    101670, 101680, 101680, 101660, 101660, 101670, 101650, 101640, 101640, 
    101640, 101670, 101680, 101690, 101700, 101690, 101690, 101690, 101680, 
    101660, 101660, 101660, 101630, 101620, 101620, 101620, 101620, 101620, 
    101620, 101610, 101610, 101590, 101570, 101540, 101530, 101510, 101490, 
    101480, 101470, 101470, 101470, 101480, 101490, 101470, 101470, 101460, 
    101460, 101460, 101470, 101470, 101460, 101460, 101480, 101470, 101470, 
    101440, 101420, 101400, 101390, 101400, 101360, 101360, 101330, 101320, 
    101250, 101240, 101210, 101170, 101110, 101100, 101050, 101050, 101010, 
    100960, 100910, 100880, 100860, 100830, 100770, 100700, 100660, 100600, 
    100640, 100580, 100560, 100530, 100510, 100520, 100490, 100450, 100440, 
    100410, 100390, 100370, 100350, 100400, 100400, 100380, 100370, 100360, 
    100350, 100340, 100340, 100310, 100310, 100310, 100300, 100270, 100260, 
    100270, 100270, 100270, 100270, 100260, 100270, 100270, 100280, 100290, 
    100300, 100330, 100350, 100360, 100380, 100400, 100420, 100440, 100480, 
    100520, 100530, 100570, 100600, 100620, 100660, 100700, 100730, 100770, 
    100810, 100840, 100890, 100940, 100970, 101010, 101070, 101130, 101180, 
    101230, 101280, 101350, 101400, 101440, 101480, 101530, 101580, 101610, 
    101640, 101680, 101730, 101760, 101790, 101820, 101850, 101890, 101920, 
    101940, 101970, 101990, 102010, 102030, 102060, 102100, 102120, 102120, 
    102130, 102130, 102120, 102140, 102150, 102140, 102160, 102170, 102180, 
    102180, 102180, 102180, 102160, 102160, 102130, 102100, 102090, 102080, 
    102070, 102040, 102040, 101990, 101950, 101980, 101950, 101930, 101940, 
    101880, 101850, 101830, 101800, 101770, 101710, 101690, 101610, 101520, 
    101500, 101530, 101530, 101450, 101380, 101340, 101310, 101300, 101260, 
    101260, 101270, 101230, 101280, 101280, 101290, 101310, 101330, 101360, 
    101350, 101370, 101380, 101400, 101420, 101440, 101450, 101460, 101480, 
    101490, 101530, 101570, 101600, 101640, 101660, 101690, 101710, 101750, 
    101780, 101810, 101830, 101870, 101900, 101920, 101940, 101970, 102000, 
    102020, 102030, 102020, 102030, 102040, 102050, 102050, 102040, 102050, 
    102070, 102090, 102090, 102110, 102120, 102110, 102100, 102100, 102110, 
    102090, 102080, 102060, 102020, 102020, 102040, 102030, 102010, 101970, 
    101990, 101960, 101950, 101950, 101940, 101900, 101910, 101970, 101980, 
    101990, 102010, 102040, 102040, 102060, 102040, 102030, 102040, 102070, 
    102100, 102100, 102120, 102120, 102130, 102140, 102150, 102150, 102150, 
    102140, 102120, 102120, 102130, 102160, 102180, 102200, 102200, 102180, 
    102170, 102150, 102150, 102120, 102120, 102090, 102080, 102080, 102090, 
    102080, 102080, 102080, 102070, 102060, 102010, 101970, 101950, 101940, 
    101950, 101970, 101970, 101970, 101950, 101930, 101910, 101890, 101880, 
    101900, 101880, 101870, 101880, 101880, 101890, 101900, 101900, 101900, 
    101910, 101930, 101940, 101950, 101970, 102020, 102050, 102070, 102100, 
    102120, 102130, 102150, 102170, 102180, 102200, 102210, 102230, 102240, 
    102250, 102280, 102290, 102290, 102300, 102290, 102290, 102290, 102290, 
    102280, 102260, 102230, 102210, 102200, 102180, 102130, 102130, 102100, 
    102070, 102030, 101990, 101980, 101920, 101870, 101810, 101790, 101780, 
    101740, 101700, 101670, 101560, 101540, 101470, 101420, 101380, 101350, 
    101330, 101320, 101310, 101290, 101270, 101250, 101240, 101230, 101220, 
    101190, 101170, 101150, 101140, 101110, 101080, 101090, 101070, 101050, 
    101050, 101020, 101020, 101010, 101010, 101000, 101000, 101000, 101010, 
    101030, 101010, 101010, 101020, 101020, 101020, 101020, 101010, 101020, 
    101030, 101030, 101060, 101080, 101100, 101110, 101130, 101140, 101120, 
    101140, 101150, 101150, 101150, 101170, 101180, 101190, 101180, 101190, 
    101200, 101210, 101190, 101170, 101150, 101170, 101180, 101170, 101170, 
    101170, 101180, 101170, 101150, 101130, 101110, 101120, 101110, 101080, 
    101090, 101100, 101090, 101090, 101110, 101110, 101110, 101110, 101110, 
    101110, 101110, 101120, 101130, 101130, 101130, 101160, 101170, 101180, 
    101190, 101180, 101180, 101180, 101180, 101180, 101200, 101220, 101240, 
    101260, 101290, 101300, 101310, 101340, 101350, 101370, 101380, 101390, 
    101410, 101420, 101440, 101470, 101480, 101490, 101510, 101510, 101510, 
    101510, 101510, 101500, 101510, 101510, 101510, 101520, 101520, 101520, 
    101500, 101520, 101520, 101500, 101480, 101480, 101510, 101500, 101500, 
    101480, 101470, 101470, 101460, 101430, 101410, 101420, 101420, 101440, 
    101450, 101460, 101460, 101460, 101460, 101450, 101430, 101410, 101400, 
    101380, 101360, 101340, 101320, 101300, 101290, 101290, 101260, 101250, 
    101220, 101190, 101160, 101120, 101090, 101080, 101060, 101060, 101060, 
    101040, 101020, 101010, 101010, 101000, 101020, 101020, 101010, 101020, 
    101030, 101040, 101030, 101040, 101060, 101080, 101100, 101130, 101160, 
    101190, 101210, 101250, 101290, 101340, 101400, 101470, 101530, 101580, 
    101650, 101700, 101750, 101790, 101820, 101850, 101930, 101970, 102040, 
    102120, 102180, 102210, 102260, 102310, 102350, 102380, 102400, 102430, 
    102450, 102500, 102530, 102550, 102590, 102620, 102620, 102600, 102610, 
    102630, 102640, 102670, 102680, 102710, 102730, 102760, 102780, 102790, 
    102790, 102800, 102800, 102800, 102790, 102780, 102750, 102730, 102720, 
    102700, 102710, 102680, 102650, 102590, 102560, 102560, 102540, 102500, 
    102490, 102490, 102500, 102480, 102450, 102450, 102410, 102370, 102330, 
    102280, 102240, 102180, 102150, 102100, 102050, 102020, 102010, 101970, 
    101960, 101910, 101880, 101840, 101770, 101690, 101610, 101570, 101530, 
    101520, 101490, 101480, 101430, 101410, 101330, 101330, 101330, 101310, 
    101280, 101280, 101300, 101280, 101270, 101310, 101320, 101300, 101320, 
    101310, 101280, 101260, 101240, 101240, 101230, 101240, 101230, 101230, 
    101260, 101260, 101250, 101240, 101240, 101260, 101280, 101290, 101310, 
    101310, 101300, 101300, 101320, 101230, 101150, 101070, 101020, 101050, 
    101040, 101070, 101050, 101060, 101110, 101110, 101130, 101160, 101180, 
    101180, 101200, 101190, 101200, 101230, 101260, 101270, 101270, 101250, 
    101240, 101230, 101260, 101240, 101250, 101260, 101260, 101280, 101320, 
    101340, 101360, 101380, 101420, 101470, 101540, 101570, 101620, 101680, 
    101730, 101800, 101820, 101870, 101910, 101940, 101980, 102040, 102050, 
    102080, 102120, 102150, 102190, 102250, 102280, 102300, 102340, 102350, 
    102390, 102410, 102420, 102440, 102450, 102470, 102510, 102550, 102560, 
    102600, 102620, 102620, 102650, 102670, 102680, 102680, 102680, 102690, 
    102680, 102710, 102710, 102710, 102710, 102700, 102670, 102630, 102590, 
    102570, 102500, 102470, 102370, 102340, 102310, 102190, 102110, 102030, 
    101940, 101850, 101780, 101680, 101590, 101520, 101500, 101480, 101480, 
    101460, 101430, 101420, 101410, 101410, 101390, 101410, 101420, 101410, 
    101420, 101430, 101450, 101450, 101480, 101480, 101480, 101490, 101510, 
    101500, 101500, 101520, 101530, 101560, 101590, 101610, 101630, 101660, 
    101670, 101680, 101690, 101730, 101730, 101750, 101760, 101780, 101790, 
    101830, 101820, 101820, 101810, 101820, 101840, 101840, 101850, 101830, 
    101850, 101880, 101880, 101890, 101910, 101920, 101910, 101910, 101920, 
    101920, 101910, 101910, 101900, 101900, 101900, 101890, 101900, 101890, 
    101890, 101870, 101850, 101840, 101820, 101790, 101770, 101750, 101740, 
    101730, 101710, 101690, 101670, 101670, 101670, 101670, 101650, 101640, 
    101640, 101650, 101650, 101680, 101690, 101690, 101720, 101730, 101720, 
    101720, 101730, 101740, 101750, 101750, 101770, 101790, 101800, 101810, 
    101820, 101830, 101810, 101800, 101790, 101780, 101790, 101820, 101820, 
    101830, 101850, 101870, 101850, 101830, 101820, 101800, 101800, 101800, 
    101780, 101790, 101790, 101760, 101720, 101740, 101720, 101670, 101620, 
    101570, 101500, 101450, 101420, 101420, 101360, 101320, 101250, 101210, 
    101200, 101180, 101120, 101050, 101050, 101040, 101000, 100990, 100960, 
    100940, 100900, 100900, 100880, 100880, 100880, 100920, 100910, 100910, 
    100930, 100940, 100980, 100990, 101000, 101030, 101020, 101040, 101030, 
    101020, 101010, 100990, 100980, 100970, 100980, 100950, 100930, 100920, 
    100900, 100880, 100870, 100840, 100800, 100810, 100810, 100810, 100800, 
    100780, 100760, 100730, 100730, 100720, 100740, 100750, 100730, 100720, 
    100770, 100780, 100780, 100820, 100840, 100880, 100910, 100910, 100960, 
    100980, 101020, 101080, 101100, 101190, 101200, 101240, 101330, 101370, 
    101430, 101490, 101530, 101560, 101630, 101650, 101670, 101710, 101760, 
    101790, 101830, 101840, 101880, 101900, 101930, 101970, 101990, 102020, 
    102050, 102070, 102060, 102060, 102070, 102080, 102070, 102070, 102050, 
    102030, 102010, 101990, 101960, 101940, 101950, 101930, 101910, 101880, 
    101860, 101830, 101800, 101760, 101700, 101670, 101640, 101590, 101540, 
    101490, 101460, 101420, 101380, 101340, 101320, 101280, 101230, 101180, 
    101150, 101130, 101110, 101090, 101080, 101060, 101050, 101050, 101050, 
    101040, 101010, 101000, 100970, 100980, 100990, 101000, 100960, 100960, 
    100960, 100930, 100890, 100840, 100800, 100760, 100730, 100720, 100690, 
    100660, 100640, 100620, 100610, 100610, 100600, 100580, 100570, 100560, 
    100570, 100580, 100580, 100600, 100620, 100630, 100640, 100660, 100680, 
    100700, 100710, 100740, 100780, 100820, 100860, 100900, 100920, 100950, 
    100980, 101000, 101030, 101040, 101060, 101070, 101090, 101110, 101130, 
    101130, 101140, 101140, 101130, 101120, 101130, 101120, 101100, 101110, 
    101090, 101090, 101090, 101080, 101080, 101060, 101050, 101020, 101000, 
    101000, 100990, 100960, 100940, 100910, 100900, 100850, 100800, 100750, 
    100710, 100680, 100640, 100570, 100540, 100470, 100390, 100310, 100240, 
    100160, 100080, 99980, 99860, 99770, 99710, 99720, 99730, 99770, 99820, 
    99890, 99920, 99970, 100010, 100030, 100060, 100100, 100120, 100110, 
    100150, 100200, 100240, 100240, 100260, 100300, 100340, 100350, 100350, 
    100340, 100380, 100390, 100400, 100420, 100450, 100480, 100520, 100530, 
    100550, 100570, 100580, 100610, 100610, 100590, 100630, 100660, 100690, 
    100750, 100820, 100870, 100930, 100990, 101070, 101120, 101180, 101210, 
    101240, 101260, 101300, 101330, 101330, 101300, 101280, 101280, 101230, 
    101160, 101080, 101040, 100970, 100910, 100890, 100870, 100870, 100860, 
    100860, 100870, 100890, 100910, 100920, 100890, 100890, 100910, 100940, 
    100950, 100980, 101010, 101010, 101010, 101000, 100990, 100950, 100900, 
    100850, 100820, 100740, 100720, 100680, 100620, 100520, 100460, 100430, 
    100410, 100420, 100450, 100450, 100520, 100550, 100670, 100710, 100780, 
    100830, 100870, 100920, 100980, 101050, 101130, 101240, 101290, 101360, 
    101400, 101420, 101430, 101450, 101490, 101480, 101460, 101440, 101420, 
    101400, 101380, 101370, 101330, 101310, 101310, 101290, 101270, 101250, 
    101270, 101340, 101360, 101380, 101400, 101470, 101510, 101550, 101540, 
    101600, 101620, 101640, 101680, 101690, 101690, 101710, 101720, 101730, 
    101720, 101740, 101730, 101710, 101690, 101670, 101640, 101590, 101550, 
    101490, 101450, 101400, 101360, 101350, 101310, 101270, 101210, 101160, 
    101130, 101110, 101090, 101070, 101070, 101050, 101060, 101090, 101100, 
    101110, 101130, 101140, 101190, 101220, 101270, 101360, 101400, 101460, 
    101520, 101570, 101630, 101670, 101730, 101760, 101780, 101800, 101820, 
    101840, 101870, 101890, 101910, 101910, 101920, 101930, 101910, 101910, 
    101890, 101860, 101840, 101850, 101860, 101830, 101820, 101790, 101780, 
    101760, 101740, 101710, 101670, 101660, 101640, 101590, 101530, 101490, 
    101470, 101440, 101390, 101350, 101330, 101300, 101290, 101260, 101270, 
    101250, 101250, 101260, 101280, 101300, 101300, 101300, 101330, 101350, 
    101350, 101360, 101390, 101390, 101400, 101400, 101420, 101430, 101440, 
    101460, 101470, 101500, 101510, 101490, 101510, 101520, 101500, 101490, 
    101490, 101500, 101520, 101520, 101540, 101550, 101530, 101510, 101490, 
    101460, 101420, 101440, 101440, 101440, 101440, 101430, 101400, 101370, 
    101350, 101340, 101350, 101350, 101360, 101380, 101420, 101430, 101430, 
    101410, 101420, 101420, 101410, 101410, 101400, 101360, 101330, 101330, 
    101350, 101350, 101320, 101340, 101340, 101350, 101340, 101320, 101300, 
    101300, 101290, 101280, 101290, 101280, 101300, 101300, 101300, 101310, 
    101310, 101320, 101330, 101320, 101340, 101390, 101430, 101470, 101490, 
    101540, 101590, 101620, 101660, 101660, 101670, 101680, 101680, 101730, 
    101790, 101850, 101860, 101900, 101910, 101900, 101880, 101880, 101870, 
    101850, 101830, 101810, 101780, 101760, 101720, 101680, 101630, 101600, 
    101540, 101470, 101440, 101390, 101350, 101300, 101270, 101270, 101210, 
    101190, 101160, 101120, 101070, 101030, 101020, 100990, 100970, 101000, 
    101020, 101000, 101000, 100970, 100970, 100970, 100980, 100980, 100980, 
    101010, 101050, 101060, 101050, 101060, 101070, 101110, 101140, 101150, 
    101160, 101160, 101180, 101180, 101220, 101230, 101250, 101260, 101260, 
    101250, 101250, 101250, 101240, 101240, 101250, 101270, 101280, 101270, 
    101280, 101290, 101290, 101290, 101290, 101290, 101280, 101270, 101280, 
    101270, 101270, 101270, 101270, 101280, 101290, 101270, 101280, 101270, 
    101260, 101260, 101270, 101280, 101300, 101300, 101330, 101360, 101380, 
    101390, 101390, 101410, 101430, 101450, 101460, 101490, 101530, 101530, 
    101560, 101590, 101610, 101650, 101660, 101680, 101710, 101740, 101760, 
    101790, 101820, 101870, 101920, 101950, 101990, 102030, 102060, 102080, 
    102110, 102140, 102180, 102230, 102280, 102300, 102330, 102350, 102380, 
    102400, 102430, 102460, 102490, 102520, 102560, 102590, 102610, 102640, 
    102680, 102710, 102740, 102770, 102780, 102800, 102810, 102840, 102840, 
    102840, 102830, 102790, 102780, 102770, 102760, 102720, 102660, 102600, 
    102530, 102460, 102380, 102300, 102210, 102120, 102050, 101950, 101850, 
    101740, 101650, 101530, 101430, 101310, 101200, 101110, 101060, 101000, 
    100950, 100930, 100880, 100810, 100730, 100640, 100540, 100440, 100310, 
    100240, 100110, 99980, 99810, 99630, 99420, 99180, 98880, 98540, 98190, 
    97890, 97540, 97240, 97020, 96800, 96660, 96620, 96610, 96590, 96600, 
    96620, 96640, 96700, 96780, 96880, 97010, 97150, 97320, 97500, 97670, 
    97820, 97950, 98100, 98250, 98350, 98460, 98570, 98680, 98790, 98860, 
    98950, 99030, 99090, 99140, 99190, 99210, 99270, 99320, 99360, 99400, 
    99420, 99460, 99500, 99540, 99560, 99570, 99600, 99620, 99630, 99660, 
    99670, 99670, 99660, 99680, 99700, 99700, 99700, 99730, 99700, 99720, 
    99720, 99740, 99720, 99730, 99730, 99770, 99790, 99800, 99820, 99850, 
    99870, 99880, 99900, 99920, 99950, 99950, 99970, 99980, 100010, 100030, 
    100030, 100060, 100100, 100120, 100140, 100170, 100200, 100240, 100270, 
    100310, 100350, 100400, 100450, 100480, 100510, 100540, 100560, 100590, 
    100610, 100630, 100640, 100660, 100690, 100730, 100750, 100770, 100800, 
    100840, 100870, 100870, 100900, 100940, 100960, 101010, 101070, 101110, 
    101150, 101190, 101240, 101290, 101330, 101380, 101420, 101460, 101500, 
    101560, 101610, 101660, 101710, 101750, 101820, 101880, 101930, 102000, 
    102050, 102100, 102160, 102220, 102270, 102320, 102370, 102440, 102520, 
    102540, 102550, 102570, 102630, 102620, 102670, 102690, 102730, 102740, 
    102760, 102770, 102790, 102800, 102740, 102750, 102730, 102710, 102700, 
    102710, 102730, 102740, 102750, 102750, 102760, 102780, 102810, 102790, 
    102800, 102830, 102850, 102870, 102890, 102900, 102900, 102900, 102920, 
    102950, 102950, 102950, 102980, 103010, 103050, 103070, 103120, 103170, 
    103150, 103160, 103170, 103190, 103210, 103210, 103190, 103180, 103170, 
    103180, 103210, 103190, 103170, 103130, 103110, 103100, 103100, 103080, 
    103070, 103050, 103040, 103040, 103050, 103040, 103030, 103010, 102980, 
    102940, 102940, 102900, 102870, 102860, 102860, 102820, 102820, 102800, 
    102790, 102760, 102730, 102710, 102660, 102630, 102560, 102540, 102540, 
    102540, 102540, 102540, 102520, 102500, 102510, 102520, 102510, 102470, 
    102460, 102420, 102380, 102350, 102320, 102270, 102250, 102220, 102170, 
    102140, 102090, 102050, 102020, 101990, 101960, 101930, 101880, 101850, 
    101800, 101740, 101680, 101620, 101560, 101500, 101400, 101320, 101240, 
    101160, 101080, 101050, 100990, 100940, 100940, 100910, 100880, 100840, 
    100810, 100770, 100730, 100700, 100680, 100630, 100570, 100530, 100500, 
    100450, 100430, 100410, 100370, 100360, 100350, 100340, 100340, 100350, 
    100340, 100360, 100390, 100420, 100460, 100490, 100530, 100560, 100600, 
    100640, 100680, 100720, 100740, 100760, 100780, 100780, 100820, 100820, 
    100840, 100860, 100880, 100870, 100880, 100880, 100890, 100900, 100890, 
    100910, 100910, 100910, 100920, 100930, 100930, 100950, 100970, 101000, 
    101020, 101050, 101060, 101100, 101110, 101120, 101130, 101170, 101180, 
    101200, 101230, 101270, 101270, 101260, 101270, 101240, 101190, 101160, 
    101120, 101070, 101000, 100970, 100900, 100850, 100790, 100720, 100640, 
    100570, 100530, 100510, 100460, 100460, 100450, 100420, 100400, 100360, 
    100330, 100310, 100270, 100180, 100090, 100060, 99990, 99860, 99730, 
    99590, 99510, 99410, 99300, 99180, 99070, 98970, 98880, 98770, 98660, 
    98540, 98460, 98380, 98310, 98250, 98180, 98120, 98120, 98150, 98140, 
    98190, 98250, 98310, 98380, 98460, 98550, 98630, 98710, 98780, 98830, 
    98910, 98980, 99030, 99110, 99170, 99230, 99300, 99370, 99440, 99500, 
    99560, 99610, 99690, 99750, 99810, 99870, 99930, 100000, 100070, 100150, 
    100220, 100290, 100340, 100380, 100440, 100500, 100530, 100510, 100570, 
    100570, 100600, 100640, 100630, 100660, 100660, 100670, 100660, 100660, 
    100690, 100660, 100640, 100640, 100620, 100600, 100560, 100510, 100460, 
    100380, 100310, 100210, 100140, 100050, 99990, 99910, 99850, 99800, 
    99730, 99640, 99550, 99540, 99500, 99460, 99410, 99380, 99320, 99300, 
    99260, 99230, 99230, 99230, 99200, 99200, 99260, 99270, 99300, 99320, 
    99340, 99390, 99490, 99580, 99610, 99710, 99760, 99870, 99960, 100060, 
    100150, 100240, 100340, 100430, 100510, 100590, 100660, 100710, 100740, 
    100780, 100790, 100830, 100850, 100860, 100850, 100830, 100800, 100770, 
    100740, 100720, 100710, 100680, 100640, 100580, 100520, 100490, 100470, 
    100430, 100390, 100350, 100310, 100260, 100190, 100140, 100100, 100070, 
    100040, 100000, 99970, 99930, 99880, 99850, 99830, 99800, 99740, 99690, 
    99640, 99630, 99630, 99610, 99560, 99530, 99540, 99550, 99560, 99580, 
    99550, 99530, 99530, 99530, 99530, 99510, 99510, 99500, 99480, 99490, 
    99480, 99480, 99480, 99490, 99500, 99500, 99510, 99510, 99510, 99510, 
    99540, 99530, 99540, 99530, 99510, 99510, 99470, 99460, 99410, 99390, 
    99390, 99370, 99340, 99340, 99260, 99220, 99210, 99180, 99110, 99080, 
    99080, 99040, 99020, 99050, 99050, 99020, 98980, 98920, 98850, 98760, 
    98660, 98530, 98440, 98350, 98260, 98160, 98070, 98020, 98010, 97920, 
    97840, 97780, 97750, 97710, 97650, 97630, 97630, 97640, 97690, 97710, 
    97780, 97840, 97890, 97990, 98050, 98130, 98220, 98320, 98400, 98500, 
    98570, 98670, 98780, 98860, 98950, 99040, 99120, 99180, 99250, 99310, 
    99370, 99460, 99540, 99650, 99740, 99820, 99860, 99940, 100010, 100110, 
    100190, 100250, 100310, 100380, 100450, 100510, 100580, 100630, 100680, 
    100710, 100750, 100780, 100780, 100800, 100810, 100840, 100870, 100900, 
    100920, 100940, 100950, 100950, 100940, 100930, 100940, 100950, 100960, 
    100980, 100990, 101040, 101060, 101090, 101140, 101200, 101250, 101290, 
    101330, 101370, 101450, 101530, 101580, 101610, 101660, 101720, 101800, 
    101850, 101900, 101940, 101990, 102030, 102050, 102050, 102100, 102110, 
    102150, 102160, 102150, 102130, 102080, 102030, 101990, 101970, 101940, 
    101940, 101930, 101920, 101900, 101910, 101890, 101880, 101850, 101840, 
    101830, 101820, 101780, 101750, 101700, 101620, 101570, 101480, 101410, 
    101330, 101260, 101220, 101140, 101050, 100950, 100880, 100830, 100830, 
    100830, 100830, 100830, 100820, 100830, 100890, 100920, 100940, 100920, 
    100900, 100920, 100850, 100840, 100840, 100840, 100810, 100780, 100740, 
    100700, 100670, 100670, 100690, 100710, 100720, 100740, 100700, 100680, 
    100640, 100590, 100510, 100440, 100310, 100240, 100100, 100040, 99910, 
    99720, 99570, 99480, 99350, 99200, 99090, 98980, 98860, 98730, 98670, 
    98590, 98530, 98480, 98450, 98410, 98400, 98400, 98400, 98390, 98400, 
    98400, 98400, 98420, 98450, 98460, 98470, 98470, 98490, 98530, 98580, 
    98570, 98570, 98570, 98610, 98650, 98700, 98700, 98730, 98780, 98840, 
    98860, 98890, 98940, 99010, 99050, 99130, 99200, 99260, 99320, 99390, 
    99440, 99490, 99530, 99580, 99590, 99620, 99650, 99670, 99710, 99740, 
    99770, 99760, 99740, 99740, 99730, 99740, 99740, 99720, 99690, 99680, 
    99660, 99650, 99630, 99630, 99630, 99660, 99660, 99650, 99680, 99690, 
    99710, 99750, 99800, 99850, 99880, 99930, 99990, 100070, 100120, 100180, 
    100210, 100260, 100310, 100380, 100430, 100490, 100550, 100610, 100690, 
    100740, 100810, 100850, 100890, 100950, 101010, 101070, 101130, 101190, 
    101250, 101300, 101370, 101380, 101460, 101520, 101560, 101590, 101620, 
    101640, 101690, 101720, 101730, 101780, 101820, 101830, 101820, 101840, 
    101860, 101860, 101850, 101850, 101850, 101860, 101820, 101800, 101790, 
    101790, 101720, 101710, 101660, 101620, 101580, 101560, 101540, 101520, 
    101480, 101470, 101440, 101390, 101340, 101270, 101220, 101170, 101120, 
    101100, 101100, 101080, 101040, 100970, 100930, 100930, 100870, 100830, 
    100760, 100700, 100650, 100610, 100570, 100500, 100510, 100480, 100380, 
    100280, 100160, 100080, 100010, 99920, 99860, 99780, 99700, 99620, 99530, 
    99440, 99370, 99320, 99250, 99200, 99170, 99120, 99090, 99100, 99090, 
    99100, 99090, 99060, 99050, 99050, 99090, 99080, 99050, 99040, 99030, 
    99060, 99100, 99120, 99180, 99230, 99260, 99260, 99280, 99300, 99320, 
    99360, 99350, 99360, 99390, 99410, 99440, 99420, 99390, 99370, 99360, 
    99340, 99310, 99310, 99300, 99280, 99290, 99300, 99320, 99280, 99330, 
    99300, 99240, 99290, 99270, 99200, 99180, 99160, 99220, 99270, 99290, 
    99320, 99370, 99460, 99480, 99520, 99570, 99610, 99720, 99800, 99870, 
    99940, 100040, 100100, 100120, 100210, 100260, 100320, 100380, 100460, 
    100510, 100560, 100620, 100690, 100770, 100810, 100850, 100890, 100920, 
    100990, 101040, 101080, 101140, 101180, 101260, 101350, 101400, 101480, 
    101550, 101600, 101640, 101700, 101750, 101780, 101850, 101900, 101960, 
    102010, 102050, 102080, 102100, 102130, 102180, 102200, 102210, 102210, 
    102230, 102210, 102220, 102240, 102220, 102250, 102230, 102190, 102150, 
    102120, 102080, 102060, 102030, 102010, 101980, 101970, 101920, 101890, 
    101860, 101820, 101710, 101610, 101550, 101520, 101390, 101380, 101320, 
    101280, 101230, 101170, 101140, 101080, 101040, 100980, 100920, 100850, 
    100740, 100650, 100600, 100530, 100420, 100370, 100270, 100150, 100070, 
    99920, 99790, 99630, 99500, 99420, 99340, 99250, 99190, 99140, 99090, 
    99040, 99010, 99010, 99040, 99040, 99030, 99030, 99020, 99020, 99030, 
    99060, 99030, 99030, 99020, 99030, 99010, 99020, 99020, 99060, 99080, 
    99080, 99060, 99080, 99080, 99050, 99030, 99010, 99000, 99000, 99010, 
    99000, 99020, 99040, 99060, 99090, 99110, 99120, 99140, 99150, 99150, 
    99160, 99170, 99200, 99220, 99240, 99250, 99250, 99250, 99240, 99250, 
    99270, 99290, 99320, 99340, 99390, 99430, 99490, 99540, 99600, 99630, 
    99650, 99690, 99740, 99750, 99780, 99850, 99880, 99920, 99970, 100030, 
    100050, 100070, 100110, 100130, 100160, 100180, 100180, 100190, 100200, 
    100200, 100230, 100220, 100180, 100190, 100170, 100160, 100150, 100130, 
    100110, 100100, 100100, 100090, 100080, 100080, 100030, 99990, 99940, 
    99910, 99860, 99810, 99750, 99720, 99680, 99650, 99620, 99620, 99580, 
    99550, 99530, 99530, 99530, 99520, 99480, 99460, 99480, 99450, 99470, 
    99470, 99460, 99470, 99480, 99470, 99500, 99490, 99520, 99510, 99550, 
    99560, 99610, 99640, 99650, 99670, 99680, 99700, 99710, 99730, 99760, 
    99810, 99860, 99900, 99940, 99970, 99980, 99970, 100000, 100010, 100030, 
    100070, 100030, 100060, 100010, 99990, 100000, 99970, 99920, 99860, 
    99770, 99700, 99580, 99410, 99300, 99200, 99100, 99010, 98880, 98790, 
    98790, 98780, 98800, 98880, 98960, 99050, 99110, 99170, 99220, 99240, 
    99240, 99220, 99210, 99210, 99220, 99200, 99220, 99250, 99280, 99280, 
    99350, 99390, 99430, 99480, 99480, 99510, 99520, 99540, 99560, 99580, 
    99650, 99660, 99670, 99660, 99720, 99740, 99790, 99800, 99800, 99820, 
    99820, 99860, 99860, 99870, 99930, 99910, 99900, 99930, 99930, 99930, 
    99910, 99950, 99960, 99930, 99880, 99860, 99850, 99870, 99890, 99900, 
    99910, 99910, 99900, 99850, 99870, 99850, 99820, 99820, 99820, 99800, 
    99800, 99820, 99800, 99780, 99730, 99740, 99720, 99690, 99660, 99630, 
    99610, 99580, 99560, 99530, 99480, 99430, 99400, 99360, 99320, 99280, 
    99230, 99180, 99130, 99100, 99020, 98990, 98950, 98900, 98860, 98820, 
    98780, 98740, 98660, 98590, 98560, 98540, 98510, 98540, 98490, 98470, 
    98440, 98410, 98390, 98410, 98400, 98400, 98470, 98470, 98490, 98510, 
    98520, 98570, 98600, 98650, 98690, 98750, 98800, 98850, 98870, 98910, 
    98950, 98940, 98970, 98970, 99010, 99020, 99080, 99070, 99080, 99090, 
    99100, 99160, 99210, 99230, 99260, 99260, 99260, 99240, 99250, 99250, 
    99250, 99220, 99200, 99200, 99190, 99200, 99170, 99130, 99100, 99060, 
    99020, 98970, 98940, 98900, 98910, 98990, 98910, 99000, 98990, 99010, 
    99020, 98990, 99020, 99030, 99050, 99070, 99050, 99050, 99080, 99110, 
    99150, 99180, 99190, 99200, 99210, 99210, 99210, 99250, 99270, 99300, 
    99310, 99310, 99310, 99290, 99280, 99300, 99340, 99380, 99430, 99480, 
    99550, 99570, 99610, 99630, 99620, 99620, 99610, 99600, 99580, 99610, 
    99630, 99650, 99690, 99750, 99790, 99830, 99890, 99900, 99920, 99960, 
    99990, 100020, 100030, 100060, 100090, 100140, 100150, 100180, 100210, 
    100230, 100250, 100250, 100260, 100260, 100270, 100260, 100280, 100280, 
    100280, 100260, 100240, 100210, 100160, 100100, 100060, 100020, 99980, 
    99920, 99850, 99780, 99710, 99640, 99570, 99510, 99460, 99410, 99330, 
    99250, 99180, 99110, 99020, 98980, 98920, 98850, 98780, 98740, 98690, 
    98630, 98610, 98550, 98520, 98480, 98450, 98450, 98430, 98380, 98350, 
    98310, 98300, 98260, 98260, 98240, 98190, 98190, 98160, 98130, 98110, 
    98120, 98120, 98150, 98130, 98130, 98120, 98080, 98110, 98090, 98070, 
    98080, 98070, 98060, 98040, 98020, 97990, 97970, 97930, 97890, 97850, 
    97830, 97780, 97680, 97590, 97540, 97520, 97530, 97600, 97650, 97670, 
    97670, 97730, 97830, 97920, 97910, 97990, 98000, 98040, 98070, 98100, 
    98130, 98180, 98210, 98220, 98290, 98340, 98360, 98390, 98420, 98400, 
    98410, 98430, 98420, 98480, 98510, 98560, 98620, 98690, 98760, 98790, 
    98840, 98900, 98950, 99000, 99070, 99110, 99180, 99210, 99280, 99360, 
    99440, 99510, 99560, 99640, 99700, 99770, 99850, 99920, 99960, 100060, 
    100120, 100190, 100250, 100340, 100430, 100510, 100560, 100650, 100700, 
    100750, 100800, 100850, 100900, 100930, 101000, 101050, 101080, 101120, 
    101130, 101140, 101130, 101110, 101100, 101080, 101060, 101040, 101030, 
    101010, 100960, 100930, 100890, 100830, 100800, 100790, 100750, 100700, 
    100690, 100690, 100670, 100690, 100690, 100680, 100690, 100660, 100650, 
    100630, 100620, 100590, 100550, 100540, 100540, 100530, 100490, 100470, 
    100440, 100420, 100360, 100280, 100190, 100100, 100010, 99920, 99830, 
    99740, 99620, 99490, 99430, 99330, 99230, 99210, 99190, 99200, 99220, 
    99190, 99200, 99210, 99290, 99320, 99360, 99370, 99390, 99400, 99400, 
    99410, 99420, 99470, 99480, 99520, 99560, 99590, 99550, 99610, 99620, 
    99650, 99680, 99660, 99670, 99710, 99750, 99770, 99810, 99830, 99820, 
    99850, 99890, 99890, 99890, 99900, 99930, 99930, 99970, 100020, 100050, 
    100080, 100080, 100100, 100120, 100130, 100110, 100080, 100110, 100130, 
    100130, 100130, 100130, 100130, 100130, 100110, 100090, 100090, 100060, 
    100050, 100030, 100040, 100070, 100080, 100080, 100080, 100080, 100060, 
    100080, 100080, 100070, 100050, 100040, 100030, 100040, 100040, 100030, 
    100000, 99980, 99970, 99980, 99970, 99960, 99950, 99940, 99930, 99920, 
    99920, 99880, 99880, 99880, 99840, 99850, 99860, 99850, 99870, 99900, 
    99910, 99960, 100020, 100060, 100090, 100100, 100150, 100200, 100270, 
    100320, 100380, 100410, 100450, 100510, 100540, 100540, 100560, 100550, 
    100600, 100640, 100680, 100740, 100790, 100850, 100920, 100980, 101050, 
    101130, 101210, 101290, 101360, 101400, 101500, 101560, 101600, 101670, 
    101720, 101770, 101840, 101880, 101910, 101940, 101970, 102030, 102030, 
    102050, 102060, 102060, 102080, 102090, 102120, 102130, 102130, 102120, 
    102110, 102100, 102060, 102050, 102030, 101990, 101960, 101970, 101950, 
    101910, 101850, 101770, 101740, 101660, 101600, 101550, 101420, 101350, 
    101230, 101160, 101100, 101020, 100930, 100800, 100700, 100580, 100420, 
    100290, 100160, 100060, 99930, 99840, 99710, 99640, 99510, 99330, 99180, 
    99030, 98880, 98730, 98570, 98440, 98320, 98250, 98160, 98010, 97900, 
    97790, 97740, 97630, 97510, 97490, 97460, 97380, 97330, 97190, 97070, 
    97260, 97290, 97370, 97430, 97420, 97380, 97340, 97280, 97330, 97290, 
    97220, 97230, 97190, 97180, 97190, 97250, 97220, 97160, 97140, 97120, 
    97050, 97040, 97080, 97090, 97090, 97070, 97070, 97080, 97070, 97040, 
    97030, 97020, 96970, 96990, 96990, 96950, 96930, 96890, 96890, 96890, 
    96880, 96860, 96840, 96830, 96830, 96850, 96860, 96890, 96900, 96920, 
    96930, 96940, 96970, 97000, 97030, 97060, 97100, 97160, 97220, 97300, 
    97360, 97410, 97480, 97550, 97630, 97700, 97790, 97890, 98010, 98130, 
    98260, 98360, 98470, 98540, 98650, 98730, 98780, 98850, 98850, 98920, 
    98980, 99030, 99080, 99110, 99130, 99130, 99170, 99230, 99210, 99210, 
    99160, 99120, 99110, 99100, 99040, 99020, 98980, 98920, 98870, 98820, 
    98740, 98630, 98550, 98480, 98390, 98370, 98380, 98380, 98350, 98330, 
    98310, 98290, 98240, 98210, 98170, 98110, 98060, 98030, 98020, 97990, 
    97960, 97920, 97890, 97870, 97860, 97810, 97770, 97740, 97710, 97670, 
    97650, 97620, 97580, 97540, 97570, 97570, 97570, 97570, 97590, 97570, 
    97580, 97620, 97660, 97700, 97740, 97740, 97710, 97710, 97730, 97780, 
    97830, 97860, 97870, 97930, 97960, 98030, 98080, 98130, 98190, 98260, 
    98330, 98390, 98430, 98460, 98530, 98580, 98610, 98700, 98740, 98820, 
    98890, 98910, 98940, 98980, 99000, 99060, 99130, 99180, 99250, 99320, 
    99390, 99470, 99540, 99610, 99690, 99770, 99860, 99930, 100000, 100050, 
    100140, 100210, 100290, 100390, 100470, 100560, 100650, 100670, 100730, 
    100780, 100790, 100830, 100820, 100680, 100530, 100490, 100450, 100420, 
    100410, 100440, 100450, 100490, 100530, 100620, 100740, 100870, 100980, 
    101040, 101190, 101280, 101380, 101460, 101480, 101480, 101510, 101530, 
    101550, 101630, 101630, 101620, 101640, 101650, 101600, 101550, 101490, 
    101430, 101370, 101360, 101360, 101280, 101230, 101190, 101140, 101070, 
    100980, 100840, 100750, 100720, 100620, 100540, 100480, 100410, 100370, 
    100340, 100250, 100140, 100030, 99940, 99830, 99710, 99680, 99690, 99710, 
    99740, 99770, 99890, 99990, 100090, 100150, 100230, 100240, 100280, 
    100280, 100240, 100280, 100260, 100270, 100260, 100250, 100140, 100050, 
    99940, 99820, 99660, 99620, 99460, 99480, 99490, 99570, 99590, 99640, 
    99670, 99690, 99700, 99790, 99890, 100010, 100120, 100230, 100350, 
    100470, 100580, 100680, 100760, 100810, 100890, 100840, 100840, 100840, 
    100840, 100830, 100810, 100730, 100680, 100620, 100510, 100390, 100320, 
    100280, 100330, 100310, 100340, 100430, 100460, 100570, 100670, 100700, 
    100730, 100760, 100720, 100670, 100610, 100620, 100530, 100390, 100350, 
    100330, 100330, 100360, 100510, 100680, 100850, 101040, 101200, 101390, 
    101560, 101710, 101890, 102060, 102140, 102130, 102090, 102020, 102020, 
    101890, 101810, 101740, 101690, 101580, 101530, 101460, 101400, 101320, 
    101250, 101230, 101160, 101200, 101300, 101300, 101340, 101350, 101370, 
    101410, 101440, 101420, 101450, 101430, 101420, 101410, 101420, 101450, 
    101480, 101500, 101530, 101530, 101530, 101560, 101610, 101610, 101630, 
    101680, 101710, 101730, 101780, 101830, 101890, 101920, 101960, 102010, 
    102060, 102090, 102120, 102150, 102170, 102210, 102220, 102250, 102270, 
    102270, 102260, 102240, 102240, 102250, 102240, 102220, 102210, 102190, 
    102190, 102170, 102150, 102140, 102120, 102090, 102060, 102040, 102030, 
    101990, 101950, 101940, 101940, 101960, 101950, 101940, 101930, 101910, 
    101910, 101900, 101930, 101950, 101960, 101990, 102010, 102040, 102060, 
    102080, 102090, 102100, 102120, 102140, 102150, 102150, 102180, 102210, 
    102230, 102260, 102300, 102310, 102330, 102310, 102340, 102340, 102330, 
    102340, 102320, 102330, 102340, 102340, 102290, 102260, 102240, 102200, 
    102190, 102150, 102110, 102070, 102010, 101980, 101950, 101960, 101960, 
    101950, 101940, 101930, 101940, 101940, 101950, 101960, 101960, 101980, 
    102000, 102030, 102050, 102050, 102070, 102080, 102100, 102110, 102130, 
    102140, 102150, 102160, 102160, 102190, 102190, 102180, 102180, 102190, 
    102180, 102170, 102170, 102170, 102170, 102160, 102170, 102180, 102200, 
    102200, 102190, 102190, 102210, 102200, 102200, 102180, 102170, 102190, 
    102220, 102250, 102280, 102270, 102270, 102290, 102280, 102270, 102260, 
    102290, 102300, 102320, 102340, 102390, 102430, 102450, 102480, 102480, 
    102490, 102520, 102540, 102560, 102590, 102630, 102690, 102750, 102790, 
    102830, 102870, 102920, 102960, 102980, 103020, 103050, 103080, 103130, 
    103170, 103230, 103250, 103270, 103300, 103300, 103330, 103350, 103380, 
    103380, 103370, 103380, 103400, 103420, 103410, 103420, 103410, 103380, 
    103370, 103340, 103300, 103260, 103240, 103170, 103130, 103090, 103030, 
    102980, 102910, 102840, 102760, 102690, 102610, 102550, 102470, 102410, 
    102370, 102340, 102330, 102290, 102250, 102200, 102160, 102100, 102060, 
    102030, 101990, 101930, 101870, 101820, 101760, 101690, 101600, 101540, 
    101460, 101380, 101290, 101170, 101060, 100980, 100940, 100910, 100940, 
    100940, 100900, 100860, 100860, 100880, 100890, 100910, 100950, 100960, 
    101000, 101040, 101080, 101150, 101170, 101190, 101210, 101260, 101300, 
    101310, 101330, 101350, 101370, 101410, 101450, 101480, 101480, 101470, 
    101470, 101500, 101520, 101510, 101510, 101520, 101510, 101530, 101530, 
    101530, 101550, 101530, 101540, 101520, 101530, 101520, 101510, 101520, 
    101530, 101590, 101660, 101670, 101660, 101700, 101730, 101720, 101740, 
    101720, 101730, 101740, 101740, 101770, 101810, 101860, 101900, 101920, 
    101910, 101910, 101920, 101930, 101920, 101930, 101870, 101870, 101880, 
    101860, 101880, 101830, 101800, 101770, 101720, 101690, 101670, 101610, 
    101600, 101570, 101530, 101470, 101430, 101360, 101320, 101260, 101220, 
    101180, 101170, 101170, 101140, 101120, 101120, 101130, 101110, 101160, 
    101170, 101180, 101190, 101180, 101200, 101190, 101170, 101180, 101190, 
    101190, 101180, 101170, 101150, 101140, 101140, 101120, 101090, 101100, 
    101090, 101080, 101080, 101060, 101050, 101030, 101020, 100990, 100970, 
    100960, 100930, 100910, 100890, 100870, 100850, 100800, 100790, 100760, 
    100740, 100710, 100680, 100650, 100650, 100640, 100630, 100630, 100660, 
    100650, 100640, 100610, 100590, 100600, 100630, 100660, 100650, 100650, 
    100700, 100720, 100720, 100750, 100760, 100770, 100770, 100780, 100770, 
    100740, 100710, 100700, 100700, 100680, 100680, 100620, 100550, 100460, 
    100440, 100420, 100390, 100310, 100280, 100240, 100200, 100170, 100140, 
    100090, 100030, 100020, 99970, 99980, 99960, 99950, 99930, 99940, 99950, 
    100010, 100040, 100050, 100070, 100080, 100100, 100120, 100120, 100100, 
    100090, 100080, 100100, 100110, 100090, 100110, 100120, 100130, 100160, 
    100190, 100250, 100280, 100310, 100370, 100400, 100480, 100560, 100600, 
    100650, 100680, 100700, 100750, 100770, 100820, 100850, 100850, 100900, 
    100880, 100940, 100950, 100940, 100950, 100970, 100960, 100970, 100920, 
    100890, 100870, 100860, 100860, 100860, 100860, 100860, 100880, 100860, 
    100850, 100860, 100870, 100860, 100850, 100870, 100910, 100910, 100920, 
    100940, 100960, 100990, 101000, 100990, 100990, 100980, 100990, 100990, 
    101040, 101090, 101150, 101150, 101170, 101190, 101230, 101260, 101270, 
    101300, 101270, 101270, 101280, 101280, 101240, 101190, 101120, 101070, 
    101000, 100920, 100860, 100790, 100700, 100630, 100610, 100540, 100480, 
    100440, 100420, 100350, 100290, 100210, 100130, 100060, 99980, 99950, 
    99880, 99830, 99760, 99700, 99630, 99550, 99500, 99440, 99370, 99320, 
    99260, 99200, 99170, 99160, 99120, 99080, 99070, 99030, 98960, 98930, 
    98900, 98870, 98820, 98790, 98790, 98760, 98740, 98720, 98700, 98690, 
    98650, 98620, 98590, 98540, 98510, 98480, 98530, 98490, 98440, 98390, 
    98350, 98330, 98320, 98330, 98290, 98300, 98280, 98250, 98220, 98190, 
    98140, 98110, 98060, 98010, 97970, 97930, 97920, 97910, 97900, 97920, 
    97940, 97960, 97970, 97960, 97980, 97950, 97930, 97930, 97950, 97940, 
    97950, 97970, 97990, 97980, 97970, 97990, 97970, 97970, 97960, 98000, 
    98040, 98100, 98100, 98130, 98220, 98290, 98390, 98430, 98480, 98530, 
    98540, 98600, 98660, 98750, 98760, 98800, 98840, 98870, 98880, 98920, 
    98970, 98960, 98970, 99010, 98990, 98970, 98970, 98980, 99030, 99060, 
    99040, 99050, 99020, 98980, 98960, 98980, 99000, 99010, 99000, 99030, 
    99030, 99050, 99040, 99100, 99020, 99100, 99130, 99130, 99140, 99190, 
    99200, 99230, 99250, 99290, 99260, 99320, 99310, 99310, 99310, 99300, 
    99270, 99300, 99320, 99320, 99370, 99420, 99400, 99450, 99490, 99460, 
    99450, 99470, 99550, 99520, 99530, 99550, 99480, 99510, 99560, 99650, 
    99680, 99730, 99750, 99830, 99890, 99860, 99890, 99910, 99980, 100010, 
    100020, 100040, 100080, 100110, 100110, 100140, 100210, 100220, 100230, 
    100270, 100320, 100350, 100380, 100380, 100450, 100510, 100540, 100540, 
    100540, 100550, 100560, 100600, 100700, 100690, 100720, 100810, 100910, 
    100960, 100970, 101030, 101090, 101150, 101170, 101170, 101230, 101220, 
    101260, 101280, 101320, 101360, 101380, 101400, 101440, 101420, 101390, 
    101370, 101350, 101370, 101360, 101310, 101280, 101260, 101230, 101190, 
    101140, 101080, 101030, 101000, 100990, 100980, 100950, 100900, 100870, 
    100830, 100790, 100770, 100740, 100680, 100640, 100640, 100620, 100610, 
    100590, 100590, 100560, 100540, 100530, 100530, 100530, 100510, 100500, 
    100490, 100520, 100520, 100540, 100550, 100540, 100510, 100530, 100510, 
    100500, 100490, 100500, 100500, 100530, 100520, 100500, 100500, 100480, 
    100460, 100460, 100460, 100450, 100440, 100440, 100460, 100460, 100450, 
    100430, 100420, 100400, 100390, 100360, 100330, 100310, 100300, 100310, 
    100280, 100290, 100260, 100230, 100200, 100160, 100130, 100100, 100070, 
    100040, 100010, 99980, 99960, 99960, 99940, 99920, 99870, 99820, 99770, 
    99750, 99740, 99710, 99660, 99630, 99590, 99560, 99530, 99430, 99330, 
    99260, 99190, 99110, 99040, 98960, 98880, 98900, 98770, 98790, 98780, 
    98780, 98710, 98690, 98630, 98600, 98560, 98530, 98530, 98500, 98510, 
    98520, 98530, 98530, 98580, 98600, 98600, 98630, 98670, 98670, 98710, 
    98710, 98720, 98750, 98770, 98830, 98850, 98850, 98860, 98890, 98900, 
    98930, 98920, 98940, 98960, 98980, 99000, 99020, 99030, 99040, 99080, 
    99100, 99120, 99140, 99140, 99150, 99180, 99240, 99260, 99280, 99300, 
    99330, 99340, 99360, 99380, 99400, 99410, 99430, 99460, 99490, 99500, 
    99540, 99560, 99620, 99670, 99720, 99760, 99800, 99840, 99900, 99990, 
    100050, 100140, 100200, 100250, 100310, 100350, 100390, 100430, 100450, 
    100470, 100480, 100490, 100500, 100540, 100550, 100560, 100560, 100560, 
    100570, 100590, 100590, 100590, 100600, 100590, 100650, 100660, 100680, 
    100690, 100700, 100700, 100700, 100690, 100640, 100600, 100550, 100510, 
    100470, 100430, 100440, 100450, 100470, 100480, 100490, 100540, 100560, 
    100580, 100620, 100670, 100740, 100780, 100830, 100850, 100850, 100870, 
    100900, 100900, 100910, 100900, 100910, 100920, 100930, 100980, 100900, 
    100910, 100850, 100780, 100700, 100700, 100680, 100630, 100600, 100580, 
    100560, 100560, 100580, 100620, 100640, 100660, 100690, 100720, 100740, 
    100740, 100740, 100760, 100790, 100780, 100750, 100730, 100710, 100690, 
    100680, 100670, 100650, 100620, 100610, 100610, 100620, 100630, 100640, 
    100650, 100670, 100680, 100670, 100680, 100700, 100700, 100700, 100730, 
    100760, 100750, 100780, 100800, 100790, 100790, 100770, 100730, 100670, 
    100640, 100600, 100570, 100540, 100480, 100450, 100440, 100370, 100290, 
    100250, 100230, 100180, 100120, 100080, 100060, 100050, 100060, 100080, 
    100090, 100080, 100090, 100140, 100150, 100180, 100190, 100220, 100270, 
    100320, 100350, 100380, 100420, 100420, 100400, 100360, 100310, 100290, 
    100230, 100170, 100170, 100170, 100160, 100100, 100040, 99960, 99880, 
    99820, 99750, 99660, 99580, 99560, 99530, 99520, 99490, 99440, 99400, 
    99360, 99280, 99240, 99190, 99190, 99150, 99110, 99070, 99070, 99060, 
    99030, 99000, 99000, 98980, 98960, 98940, 98930, 98890, 98920, 98970, 
    98990, 99040, 99090, 99150, 99160, 99190, 99220, 99270, 99320, 99370, 
    99420, 99480, 99540, 99630, 99690, 99740, 99790, 99840, 99890, 99940, 
    99980, 100020, 100040, 100050, 100100, 100120, 100120, 100150, 100160, 
    100140, 100130, 100110, 100090, 100040, 100000, 99990, 99930, 99890, 
    99890, 99840, 99830, 99780, 99720, 99670, 99680, 99690, 99710, 99710, 
    99690, 99730, 99750, 99800, 99820, 99830, 99850, 99930, 99970, 100020, 
    100090, 100150, 100190, 100240, 100300, 100350, 100380, 100430, 100480, 
    100520, 100560, 100590, 100610, 100630, 100670, 100720, 100710, 100710, 
    100710, 100650, 100650, 100670, 100730, 100740, 100780, 100820, 100850, 
    100890, 100940, 101000, 101060, 101120, 101200, 101250, 101300, 101330, 
    101360, 101390, 101450, 101490, 101530, 101540, 101530, 101550, 101580, 
    101600, 101600, 101580, 101580, 101580, 101580, 101600, 101600, 101590, 
    101580, 101560, 101540, 101550, 101530, 101490, 101480, 101500, 101500, 
    101480, 101490, 101470, 101430, 101410, 101410, 101390, 101400, 101410, 
    101410, 101400, 101430, 101440, 101420, 101410, 101410, 101390, 101400, 
    101410, 101400, 101410, 101420, 101460, 101440, 101450, 101480, 101510, 
    101510, 101500, 101470, 101480, 101490, 101480, 101490, 101510, 101500, 
    101490, 101460, 101440, 101400, 101360, 101320, 101300, 101290, 101250, 
    101220, 101190, 101190, 101170, 101140, 101100, 101070, 101050, 101030, 
    101010, 100970, 100910, 100890, 100890, 100850, 100830, 100810, 100780, 
    100760, 100750, 100740, 100730, 100720, 100700, 100710, 100700, 100700, 
    100720, 100720, 100710, 100700, 100690, 100670, 100670, 100660, 100650, 
    100640, 100630, 100630, 100630, 100630, 100600, 100580, 100560, 100540, 
    100530, 100500, 100480, 100470, 100450, 100460, 100450, 100460, 100450, 
    100460, 100460, 100450, 100440, 100440, 100420, 100400, 100380, 100330, 
    100290, 100280, 100240, 100220, 100190, 100160, 100150, 100120, 100120, 
    100090, 100080, 100080, 100090, 100130, 100130, 100150, 100160, 100160, 
    100160, 100170, 100180, 100150, 100130, 100090, 100050, 99990, 99940, 
    99880, 99790, 99690, 99580, 99500, 99470, 99390, 99370, 99350, 99370, 
    99430, 99480, 99520, 99510, 99490, 99530, 99520, 99550, 99570, 99600, 
    99640, 99660, 99720, 99780, 99820, 99850, 99860, 99860, 99860, 99860, 
    99870, 99860, 99890, 99920, 99950, 99970, 100000, 99990, 99990, 99990, 
    100000, 100000, 100010, 100040, 100070, 100080, 100100, 100130, 100120, 
    100120, 100170, 100170, 100180, 100200, 100230, 100240, 100230, 100270, 
    100290, 100290, 100310, 100290, 100270, 100270, 100270, 100270, 100240, 
    100210, 100210, 100210, 100220, 100230, 100210, 100200, 100170, 100160, 
    100140, 100140, 100120, 100130, 100080, 100090, 100080, 100080, 100080, 
    100120, 100170, 100220, 100230, 100280, 100340, 100380, 100420, 100460, 
    100490, 100490, 100490, 100510, 100510, 100520, 100530, 100540, 100560, 
    100570, 100600, 100610, 100660, 100660, 100680, 100710, 100730, 100750, 
    100780, 100810, 100830, 100870, 100910, 100940, 100980, 101010, 101040, 
    101040, 101050, 101060, 101050, 101070, 101080, 101080, 101100, 101100, 
    101140, 101130, 101110, 101100, 101100, 101080, 101080, 101080, 101080, 
    101090, 101080, 101090, 101100, 101100, 101100, 101100, 101120, 101140, 
    101170, 101180, 101210, 101230, 101250, 101290, 101320, 101340, 101350, 
    101360, 101370, 101400, 101410, 101440, 101460, 101490, 101510, 101530, 
    101550, 101580, 101590, 101580, 101580, 101580, 101580, 101560, 101570, 
    101550, 101570, 101590, 101570, 101580, 101560, 101530, 101520, 101500, 
    101510, 101520, 101510, 101480, 101460, 101440, 101420, 101410, 101410, 
    101400, 101410, 101410, 101410, 101390, 101410, 101390, 101410, 101410, 
    101430, 101460, 101470, 101470, 101460, 101480, 101460, 101430, 101440, 
    101440, 101400, 101380, 101350, 101310, 101300, 101310, 101300, 101260, 
    101240, 101190, 101160, 101140, 101110, 101080, 101050, 101060, 101000, 
    100950, 100860, 100750, 100700, 100610, 100500, 100410, 100370, 100320, 
    100300, 100280, 100350, 100380, 100410, 100440, 100480, 100510, 100540, 
    100510, 100500, 100520, 100520, 100520, 100530, 100500, 100530, 100500, 
    100500, 100460, 100470, 100470, 100440, 100380, 100360, 100310, 100260, 
    100210, 100150, 100040, 99900, 99720, 99540, 99390, 99240, 99160, 99220, 
    99230, 99240, 99250, 99200, 99180, 99180, 99170, 99100, 99070, 99110, 
    99150, 99340, 99550, 99730, 99950, 100120, 100310, 100440, 100580, 
    100680, 100720, 100740, 100740, 100700, 100660, 100500, 100350, 100190, 
    99930, 99660, 99380, 99050, 98750, 98510, 98270, 98110, 97980, 97900, 
    97880, 97910, 97970, 98060, 98180, 98300, 98460, 98650, 98850, 99070, 
    99260, 99460, 99600, 99720, 99850, 99950, 100070, 100200, 100280, 100400, 
    100480, 100550, 100580, 100630, 100620, 100650, 100650, 100680, 100730, 
    100750, 100790, 100800, 100850, 100890, 100890, 100880, 100900, 100890, 
    100930, 100970, 101000, 101030, 101060, 101160, 101230, 101280, 101330, 
    101370, 101430, 101490, 101510, 101530, 101560, 101590, 101620, 101640, 
    101680, 101740, 101770, 101790, 101790, 101820, 101820, 101810, 101830, 
    101800, 101820, 101840, 101840, 101870, 101880, 101870, 101860, 101830, 
    101820, 101790, 101790, 101750, 101720, 101700, 101710, 101670, 101740, 
    101700, 101690, 101660, 101630, 101600, 101520, 101530, 101520, 101520, 
    101500, 101490, 101490, 101460, 101420, 101400, 101370, 101340, 101300, 
    101280, 101260, 101240, 101220, 101220, 101210, 101190, 101160, 101160, 
    101190, 101170, 101170, 101140, 101120, 101130, 101140, 101150, 101150, 
    101150, 101140, 101130, 101140, 101170, 101130, 101130, 101150, 101190, 
    101210, 101230, 101240, 101240, 101230, 101240, 101220, 101230, 101220, 
    101210, 101190, 101190, 101160, 101160, 101160, 101140, 101090, 101050, 
    101040, 101020, 100990, 100980, 100950, 100930, 100940, 100920, 100910, 
    100890, 100860, 100830, 100810, 100810, 100780, 100770, 100760, 100740, 
    100730, 100730, 100710, 100700, 100690, 100670, 100670, 100650, 100640, 
    100640, 100640, 100650, 100650, 100660, 100690, 100690, 100710, 100740, 
    100740, 100780, 100770, 100810, 100830, 100840, 100870, 100900, 100910, 
    100930, 100950, 100950, 100950, 100970, 100970, 100980, 100970, 101010, 
    101020, 101050, 101050, 101070, 101100, 101110, 101130, 101110, 101100, 
    101100, 101070, 101050, 101030, 101010, 101020, 101000, 100980, 100940, 
    100930, 100910, 100890, 100870, 100860, 100860, 100860, 100860, 100850, 
    100850, 100820, 100810, 100810, 100810, 100800, 100790, 100790, 100790, 
    100790, 100770, 100750, 100740, 100720, 100730, 100710, 100690, 100670, 
    100670, 100640, 100610, 100590, 100590, 100570, 100550, 100550, 100550, 
    100530, 100530, 100530, 100520, 100530, 100550, 100570, 100570, 100560, 
    100560, 100560, 100560, 100550, 100540, 100520, 100510, 100490, 100470, 
    100460, 100440, 100420, 100390, 100350, 100320, 100280, 100230, 100190, 
    100170, 100150, 100080, 100040, 99980, 99950, 99870, 99800, 99760, 99710, 
    99640, 99580, 99500, 99450, 99380, 99340, 99270, 99220, 99100, 98990, 
    98920, 98750, 98630, 98510, 98420, 98340, 98270, 98170, 98130, 98070, 
    97990, 97930, 97830, 97760, 97680, 97660, 97600, 97540, 97490, 97440, 
    97390, 97330, 97310, 97310, 97320, 97300, 97350, 97380, 97420, 97490, 
    97580, 97680, 97790, 97900, 98020, 98130, 98240, 98320, 98380, 98420, 
    98500, 98560, 98650, 98740, 98790, 98840, 98880, 98920, 98960, 98980, 
    99000, 99020, 99040, 99050, 99090, 99090, 99110, 99100, 99110, 99120, 
    99140, 99160, 99160, 99180, 99200, 99250, 99250, 99290, 99310, 99310, 
    99330, 99340, 99340, 99350, 99350, 99340, 99340, 99350, 99350, 99340, 
    99370, 99400, 99410, 99430, 99450, 99470, 99510, 99530, 99580, 99630, 
    99660, 99710, 99750, 99810, 99870, 99910, 99970, 100010, 100090, 100120, 
    100160, 100210, 100250, 100310, 100380, 100440, 100510, 100580, 100630, 
    100650, 100690, 100740, 100780, 100830, 100880, 100940, 100990, 101020, 
    101070, 101090, 101150, 101170, 101190, 101250, 101290, 101330, 101350, 
    101390, 101430, 101430, 101450, 101480, 101490, 101510, 101530, 101530, 
    101540, 101560, 101580, 101590, 101610, 101630, 101640, 101660, 101640, 
    101660, 101670, 101670, 101680, 101690, 101700, 101710, 101720, 101730, 
    101710, 101700, 101690, 101700, 101700, 101710, 101720, 101740, 101750, 
    101750, 101780, 101780, 101770, 101750, 101740, 101710, 101700, 101720, 
    101720, 101750, 101740, 101760, 101770, 101790, 101780, 101770, 101770, 
    101750, 101730, 101740, 101740, 101740, 101770, 101800, 101830, 101830, 
    101850, 101860, 101850, 101860, 101860, 101870, 101870, 101890, 101920, 
    101930, 101920, 101900, 101870, 101850, 101850, 101830, 101820, 101820, 
    101810, 101820, 101810, 101800, 101800, 101790, 101780, 101760, 101740, 
    101710, 101680, 101670, 101660, 101640, 101640, 101650, 101650, 101620, 
    101590, 101570, 101530, 101530, 101520, 101520, 101510, 101510, 101520, 
    101520, 101530, 101520, 101500, 101480, 101490, 101480, 101480, 101480, 
    101470, 101460, 101460, 101470, 101480, 101490, 101520, 101540, 101550, 
    101560, 101590, 101620, 101640, 101670, 101690, 101700, 101710, 101720, 
    101730, 101730, 101720, 101720, 101720, 101740, 101740, 101740, 101750, 
    101740, 101760, 101760, 101730, 101710, 101720, 101710, 101710, 101700, 
    101710, 101710, 101700, 101710, 101700, 101660, 101660, 101630, 101610, 
    101610, 101620, 101600, 101580, 101580, 101560, 101560, 101550, 101540, 
    101490, 101450, 101420, 101390, 101370, 101340, 101330, 101290, 101260, 
    101230, 101220, 101220, 101190, 101200, 101200, 101220, 101240, 101270, 
    101300, 101350, 101390, 101420, 101400, 101420, 101490, 101490, 101520, 
    101550, 101580, 101600, 101640, 101650, 101670, 101710, 101720, 101700, 
    101730, 101760, 101760, 101810, 101790, 101810, 101810, 101840, 101870, 
    101880, 101880, 101890, 101920, 101930, 101950, 101970, 101980, 101930, 
    101950, 101970, 102010, 102030, 101990, 102020, 102020, 102030, 102020, 
    102000, 101990, 102000, 102010, 102040, 102070, 102060, 102120, 102110, 
    102140, 102180, 102200, 102210, 102210, 102190, 102200, 102180, 102190, 
    102210, 102220, 102210, 102200, 102220, 102190, 102170, 102150, 102130, 
    102110, 102090, 102100, 102080, 102040, 102010, 101970, 101930, 101870, 
    101860, 101770, 101730, 101680, 101610, 101560, 101510, 101430, 101400, 
    101370, 101310, 101260, 101230, 101220, 101190, 101180, 101160, 101150, 
    101150, 101140, 101130, 101130, 101120, 101130, 101120, 101100, 101090, 
    101070, 101040, 101120, 101120, 101140, 101140, 101190, 101190, 101180, 
    101220, 101220, 101250, 101240, 101240, 101280, 101270, 101290, 101330, 
    101320, 101330, 101350, 101320, 101340, 101340, 101360, 101340, 101370, 
    101380, 101400, 101400, 101430, 101440, 101430, 101440, 101430, 101420, 
    101430, 101440, 101460, 101470, 101460, 101470, 101470, 101470, 101480, 
    101500, 101480, 101480, 101480, 101510, 101520, 101530, 101540, 101550, 
    101550, 101540, 101550, 101540, 101550, 101560, 101580, 101590, 101610, 
    101610, 101600, 101570, 101570, 101570, 101560, 101530, 101510, 101490, 
    101470, 101460, 101460, 101410, 101420, 101380, 101360, 101350, 101310, 
    101300, 101280, 101250, 101220, 101200, 101180, 101160, 101170, 101160, 
    101140, 101110, 101080, 101060, 101060, 101020, 101010, 101000, 100980, 
    100940, 100920, 100900, 100880, 100850, 100830, 100810, 100780, 100770, 
    100790, 100760, 100770, 100780, 100800, 100810, 100820, 100840, 100860, 
    100870, 100880, 100900, 100910, 100910, 100940, 100950, 100970, 101010, 
    101030, 101040, 101060, 101070, 101070, 101090, 101100, 101110, 101110, 
    101120, 101120, 101140, 101140, 101140, 101150, 101130, 101130, 101130, 
    101140, 101140, 101150, 101160, 101170, 101190, 101220, 101220, 101230, 
    101240, 101250, 101250, 101260, 101260, 101280, 101300, 101330, 101350, 
    101360, 101380, 101400, 101410, 101420, 101450, 101470, 101500, 101530, 
    101550, 101570, 101590, 101600, 101630, 101630, 101640, 101640, 101620, 
    101630, 101610, 101600, 101600, 101580, 101550, 101520, 101490, 101480, 
    101450, 101440, 101430, 101420, 101410, 101420, 101420, 101410, 101410, 
    101380, 101390, 101370, 101360, 101340, 101320, 101320, 101330, 101340, 
    101330, 101320, 101340, 101320, 101330, 101310, 101290, 101270, 101260, 
    101250, 101250, 101250, 101240, 101230, 101200, 101190, 101170, 101160, 
    101160, 101160, 101170, 101170, 101190, 101220, 101260, 101280, 101300, 
    101320, 101340, 101360, 101400, 101450, 101470, 101510, 101580, 101640, 
    101670, 101720, 101780, 101830, 101860, 101910, 101950, 101980, 102020, 
    102040, 102100, 102150, 102180, 102220, 102260, 102290, 102310, 102320, 
    102350, 102360, 102390, 102430, 102460, 102490, 102540, 102590, 102640, 
    102690, 102730, 102750, 102770, 102830, 102860, 102900, 102960, 103020, 
    103060, 103110, 103160, 103200, 103230, 103270, 103310, 103350, 103390, 
    103440, 103490, 103530, 103570, 103590, 103610, 103600, 103620, 103580, 
    103580, 103620, 103610, 103610, 103590, 103590, 103580, 103590, 103550, 
    103560, 103580, 103530, 103490, 103460, 103470, 103470, 103500, 103510, 
    103500, 103500, 103480, 103490, 103480, 103450, 103430, 103410, 103410, 
    103380, 103370, 103360, 103370, 103360, 103310, 103290, 103260, 103210, 
    103160, 103120, 103090, 103080, 103070, 103060, 103030, 103000, 103010, 
    103030, 103020, 103010, 103020, 103030, 103070, 103120, 103170, 103200, 
    103240, 103310, 103350, 103370, 103400, 103430, 103460, 103480, 103520, 
    103550, 103570, 103590, 103610, 103620, 103640, 103670, 103680, 103660, 
    103630, 103620, 103590, 103570, 103540, 103550, 103520, 103510, 103490, 
    103470, 103450, 103430, 103410, 103380, 103360, 103330, 103300, 103290, 
    103260, 103220, 103170, 103120, 103100, 103050, 103000, 102930, 102850, 
    102810, 102770, 102730, 102680, 102630, 102590, 102530, 102490, 102450, 
    102400, 102350, 102270, 102220, 102180, 102140, 102130, 102130, 102110, 
    102100, 102070, 102040, 102030, 102010, 101990, 101980, 101960, 101960, 
    101950, 101940, 101950, 101970, 101980, 101980, 101960, 101940, 101910, 
    101920, 101930, 101930, 101960, 101980, 101980, 101990, 101980, 101980, 
    101980, 101970, 101960, 101950, 101950, 101960, 101980, 102010, 102020, 
    102030, 102040, 102040, 102030, 102040, 102060, 102090, 102120, 102160, 
    102210, 102230, 102260, 102280, 102310, 102340, 102340, 102340, 102360, 
    102380, 102400, 102430, 102460, 102470, 102490, 102480, 102480, 102470, 
    102490, 102480, 102450, 102450, 102460, 102470, 102470, 102450, 102430, 
    102420, 102410, 102380, 102340, 102300, 102290, 102260, 102230, 102210, 
    102200, 102180, 102160, 102130, 102120, 102100, 102080, 102070, 102050, 
    102080, 102110, 102140, 102160, 102190, 102190, 102210, 102220, 102240, 
    102240, 102270, 102280, 102280, 102290, 102290, 102300, 102300, 102280, 
    102270, 102250, 102220, 102180, 102160, 102140, 102130, 102120, 102130, 
    102140, 102110, 102110, 102100, 102090, 102080, 102050, 102030, 101990, 
    101970, 101950, 101910, 101920, 101920, 101900, 101880, 101850, 101830, 
    101810, 101810, 101800, 101780, 101790, 101780, 101770, 101760, 101760, 
    101770, 101750, 101720, 101680, 101660, 101620, 101620, 101600, 101570, 
    101560, 101540, 101500, 101470, 101450, 101440, 101440, 101410, 101410, 
    101410, 101410, 101430, 101440, 101470, 101480, 101500, 101530, 101540, 
    101550, 101550, 101580, 101620, 101620, 101660, 101690, 101730, 101750, 
    101790, 101810, 101840, 101840, 101860, 101880, 101900, 101920, 101940, 
    101960, 101980, 101980, 101990, 101990, 101990, 101990, 101980, 101960, 
    101950, 101930, 101930, 101930, 101930, 101920, 101910, 101900, 101900, 
    101890, 101860, 101880, 101890, 101890, 101890, 101910, 101910, 101900, 
    101900, 101900, 101890, 101870, 101850, 101810, 101820, 101820, 101810, 
    101740, 101720, 101730, 101710, 101710, 101700, 101660, 101620, 101570, 
    101530, 101510, 101470, 101450, 101420, 101360, 101270, 101230, 101170, 
    101130, 101130, 101100, 101080, 101070, 101050, 101050, 101020, 100930, 
    100850, 100820, 100730, 100680, 100660, 100590, 100600, 100590, 100610, 
    100630, 100670, 100710, 100760, 100830, 100900, 100940, 100990, 101050, 
    101100, 101130, 101170, 101210, 101240, 101280, 101340, 101360, 101390, 
    101420, 101410, 101420, 101450, 101470, 101480, 101490, 101520, 101540, 
    101530, 101540, 101550, 101530, 101530, 101530, 101500, 101480, 101450, 
    101450, 101420, 101420, 101400, 101380, 101340, 101310, 101240, 101210, 
    101140, 101090, 101030, 101010, 100990, 100940, 100880, 100830, 100770, 
    100720, 100660, 100570, 100530, 100470, 100390, 100320, 100250, 100200, 
    100150, 100110, 100060, 100020, 99990, 99990, 99970, 99950, 99930, 99910, 
    99910, 99910, 99920, 99910, 99900, 99890, 99890, 99880, 99890, 99900, 
    99910, 99910, 99920, 99930, 99930, 99940, 99930, 99920, 99920, 99930, 
    99930, 99950, 99980, 99990, 100020, 100040, 100050, 100040, 100050, 
    100040, 100040, 100040, 100030, 100040, 100040, 100050, 100050, 100040, 
    100030, 100020, 100000, 99970, 99940, 99930, 99950, 99960, 99970, 99990, 
    100010, 100010, 99990, 99970, 99930, 99930, 99880, 99870, 99860, 99840, 
    99830, 99820, 99770, 99750, 99740, 99730, 99700, 99650, 99620, 99530, 
    99550, 99600, 99610, 99630, 99680, 99680, 99710, 99730, 99710, 99700, 
    99700, 99700, 99700, 99690, 99690, 99710, 99710, 99680, 99700, 99710, 
    99690, 99700, 99730, 99780, 99830, 99840, 99870, 99920, 99970, 99990, 
    100030, 100070, 100110, 100140, 100170, 100190, 100230, 100270, 100300, 
    100330, 100380, 100410, 100440, 100450, 100480, 100500, 100520, 100550, 
    100580, 100610, 100640, 100670, 100710, 100740, 100780, 100810, 100850, 
    100890, 100930, 100970, 101020, 101060, 101090, 101170, 101220, 101280, 
    101320, 101360, 101400, 101420, 101440, 101480, 101470, 101490, 101520, 
    101530, 101530, 101550, 101590, 101630, 101660, 101670, 101710, 101720, 
    101740, 101780, 101800, 101830, 101870, 101890, 101910, 101940, 101950, 
    101960, 101970, 101980, 102000, 102020, 102030, 102040, 102050, 102050, 
    102010, 101990, 101950, 101920, 101890, 101870, 101860, 101820, 101810, 
    101780, 101760, 101750, 101690, 101650, 101630, 101580, 101570, 101580, 
    101580, 101590, 101600, 101620, 101620, 101630, 101620, 101610, 101590, 
    101580, 101560, 101550, 101570, 101580, 101590, 101590, 101560, 101570, 
    101570, 101560, 101550, 101550, 101540, 101550, 101560, 101550, 101540, 
    101530, 101530, 101530, 101530, 101520, 101510, 101500, 101520, 101510, 
    101530, 101540, 101550, 101550, 101550, 101570, 101580, 101610, 101620, 
    101610, 101620, 101640, 101650, 101670, 101690, 101690, 101690, 101700, 
    101720, 101730, 101720, 101730, 101720, 101720, 101720, 101710, 101690, 
    101700, 101710, 101700, 101690, 101680, 101670, 101620, 101580, 101540, 
    101510, 101490, 101470, 101430, 101390, 101360, 101330, 101290, 101260, 
    101250, 101210, 101170, 101140, 101120, 101110, 101110, 101110, 101060, 
    101040, 101000, 100980, 100930, 100860, 100770, 100720, 100610, 100530, 
    100480, 100430, 100430, 100490, 100520, 100520, 100520, 100520, 100560, 
    100570, 100590, 100600, 100620, 100640, 100640, 100640, 100630, 100650, 
    100620, 100600, 100610, 100620, 100690, 100750, 100840, 100950, 101040, 
    101160, 101260, 101390, 101450, 101560, 101620, 101750, 101850, 101960, 
    102070, 102160, 102250, 102370, 102480, 102500, 102570, 102670, 102710, 
    102770, 102830, 102890, 102940, 103010, 103050, 103080, 103120, 103160, 
    103190, 103210, 103220, 103230, 103250, 103270, 103270, 103280, 103290, 
    103280, 103270, 103250, 103220, 103210, 103180, 103140, 103130, 103110, 
    103080, 103060, 103030, 102990, 102950, 102920, 102860, 102810, 102770, 
    102720, 102670, 102620, 102570, 102510, 102460, 102400, 102330, 102280, 
    102220, 102160, 102110, 102040, 101990, 101940, 101890, 101840, 101810, 
    101770, 101750, 101720, 101690, 101640, 101620, 101590, 101580, 101570, 
    101560, 101550, 101550, 101540, 101540, 101540, 101560, 101590, 101620, 
    101660, 101720, 101790, 101870, 101920, 101960, 102020, 102070, 102100, 
    102140, 102130, 102140, 102130, 102150, 102130, 102130, 102130, 102080, 
    102040, 102010, 101960, 101890, 101830, 101770, 101720, 101650, 101620, 
    101580, 101500, 101440, 101370, 101320, 101270, 101230, 101210, 101170, 
    101200, 101180, 101220, 101220, 101250, 101270, 101250, 101280, 101320, 
    101340, 101330, 101350, 101390, 101410, 101440, 101460, 101490, 101510, 
    101530, 101540, 101540, 101570, 101550, 101540, 101570, 101560, 101530, 
    101560, 101570, 101530, 101550, 101570, 101560, 101580, 101560, 101550, 
    101580, 101580, 101580, 101590, 101660, 101700, 101740, 101750, 101770, 
    101800, 101820, 101860, 101890, 101930, 101990, 102030, 102070, 102090, 
    102110, 102140, 102150, 102160, 102170, 102170, 102190, 102210, 102250, 
    102260, 102260, 102280, 102290, 102310, 102310, 102280, 102270, 102240, 
    102230, 102210, 102200, 102190, 102150, 102130, 102110, 102080, 102060, 
    102020, 101990, 101960, 101930, 101920, 101910, 101890, 101870, 101850, 
    101820, 101770, 101770, 101750, 101720, 101680, 101650, 101630, 101620, 
    101580, 101570, 101550, 101540, 101520, 101500, 101470, 101440, 101420, 
    101410, 101410, 101390, 101380, 101360, 101360, 101340, 101340, 101320, 
    101310, 101300, 101300, 101310, 101320, 101320, 101340, 101350, 101390, 
    101400, 101420, 101410, 101420, 101420, 101410, 101430, 101450, 101490, 
    101530, 101550, 101560, 101570, 101570, 101550, 101560, 101560, 101560, 
    101570, 101580, 101580, 101570, 101550, 101540, 101510, 101500, 101490, 
    101470, 101460, 101450, 101450, 101460, 101440, 101430, 101420, 101450, 
    101450, 101400, 101400, 101400, 101400, 101390, 101370, 101390, 101410, 
    101410, 101410, 101400, 101390, 101370, 101340, 101320, 101290, 101260, 
    101230, 101190, 101160, 101120, 101080, 101040, 100980, 100940, 100910, 
    100870, 100820, 100790, 100760, 100700, 100670, 100630, 100620, 100620, 
    100620, 100630, 100650, 100650, 100640, 100650, 100680, 100710, 100730, 
    100760, 100790, 100830, 100840, 100860, 100850, 100860, 100880, 100890, 
    100910, 100930, 100950, 100970, 101010, 101020, 101030, 101040, 101040, 
    101050, 101040, 101040, 101040, 101060, 101070, 101070, 101070, 101070, 
    101080, 101070, 101070, 101090, 101080, 101080, 101100, 101130, 101140, 
    101160, 101170, 101180, 101220, 101240, 101240, 101250, 101250, 101270, 
    101300, 101340, 101360, 101380, 101400, 101440, 101450, 101460, 101470, 
    101500, 101530, 101550, 101570, 101610, 101640, 101660, 101690, 101710, 
    101730, 101750, 101760, 101780, 101810, 101810, 101830, 101850, 101880, 
    101870, 101870, 101870, 101890, 101890, 101890, 101890, 101900, 101870, 
    101830, 101830, 101800, 101790, 101770, 101750, 101710, 101670, 101580, 
    101520, 101510, 101480, 101400, 101320, 101210, 101180, 101130, 101030, 
    100950, 100870, 100790, 100730, 100650, 100640, 100610, 100590, 100580, 
    100560, 100590, 100560, 100530, 100520, 100470, 100450, 100440, 100430, 
    100410, 100410, 100410, 100430, 100450, 100490, 100490, 100510, 100520, 
    100520, 100530, 100550, 100570, 100610, 100640, 100660, 100680, 100670, 
    100680, 100690, 100710, 100740, 100760, 100760, 100770, 100800, 100800, 
    100820, 100840, 100860, 100870, 100890, 100900, 100930, 100940, 100970, 
    100960, 100970, 101030, 101080, 101070, 101060, 101040, 101030, 100980, 
    100950, 100920, 100900, 100880, 100870, 100860, 100860, 100850, 100830, 
    100820, 100800, 100780, 100760, 100750, 100740, 100720, 100730, 100720, 
    100740, 100730, 100730, 100720, 100700, 100680, 100650, 100620, 100610, 
    100590, 100590, 100580, 100570, 100570, 100550, 100550, 100540, 100530, 
    100550, 100520, 100520, 100510, 100500, 100500, 100500, 100490, 100460, 
    100470, 100430, 100430, 100430, 100420, 100400, 100400, 100420, 100420, 
    100440, 100460, 100490, 100530, 100570, 100600, 100600, 100620, 100600, 
    100640, 100660, 100670, 100700, 100710, 100710, 100720, 100750, 100750, 
    100750, 100770, 100790, 100800, 100820, 100850, 100860, 100880, 100870, 
    100890, 100890, 100910, 100910, 100900, 100860, 100830, 100840, 100840, 
    100840, 100820, 100810, 100830, 100810, 100790, 100790, 100770, 100750, 
    100760, 100760, 100760, 100730, 100740, 100730, 100750, 100740, 100730, 
    100730, 100710, 100700, 100680, 100650, 100650, 100630, 100620, 100590, 
    100560, 100540, 100520, 100500, 100490, 100500, 100470, 100480, 100490, 
    100530, 100580, 100590, 100630, 100650, 100640, 100680, 100690, 100710, 
    100730, 100750, 100770, 100800, 100780, 100790, 100780, 100780, 100770, 
    100780, 100770, 100760, 100760, 100760, 100790, 100810, 100840, 100850, 
    100890, 100890, 100920, 100950, 100960, 100970, 101000, 101030, 101070, 
    101120, 101140, 101180, 101200, 101230, 101260, 101280, 101290, 101310, 
    101350, 101390, 101420, 101460, 101480, 101510, 101540, 101560, 101570, 
    101580, 101580, 101600, 101610, 101620, 101620, 101630, 101650, 101640, 
    101650, 101640, 101620, 101610, 101620, 101590, 101570, 101550, 101550, 
    101560, 101530, 101520, 101510, 101490, 101420, 101390, 101370, 101330, 
    101290, 101270, 101250, 101220, 101170, 101140, 101130, 101090, 101060, 
    101010, 100970, 100940, 100920, 100920, 100930, 100970, 100990, 101010, 
    101010, 101000, 101020, 101020, 101040, 101050, 101070, 101090, 101110, 
    101140, 101150, 101160, 101150, 101160, 101140, 101150, 101130, 101140, 
    101150, 101140, 101150, 101150, 101150, 101150, 101150, 101170, 101160, 
    101160, 101160, 101170, 101180, 101180, 101200, 101240, 101260, 101280, 
    101290, 101310, 101310, 101350, 101380, 101380, 101400, 101420, 101450, 
    101460, 101480, 101510, 101510, 101520, 101520, 101540, 101550, 101560, 
    101590, 101580, 101600, 101610, 101620, 101640, 101640, 101650, 101660, 
    101660, 101640, 101630, 101630, 101640, 101650, 101630, 101640, 101640, 
    101610, 101610, 101580, 101560, 101540, 101500, 101480, 101480, 101460, 
    101470, 101470, 101440, 101420, 101400, 101370, 101370, 101370, 101370, 
    101370, 101360, 101360, 101370, 101380, 101370, 101380, 101370, 101360, 
    101350, 101350, 101330, 101330, 101340, 101340, 101340, 101320, 101310, 
    101310, 101300, 101280, 101250, 101220, 101200, 101170, 101140, 101090, 
    101080, 101050, 101030, 101000, 100970, 100950, 100920, 100890, 100870, 
    100850, 100840, 100830, 100840, 100850, 100840, 100820, 100790, 100760, 
    100700, 100650, 100640, 100600, 100550, 100510, 100460, 100400, 100340, 
    100300, 100250, 100200, 100150, 100010, 99960, 99900, 99790, 99650, 
    99500, 99320, 99180, 99210, 99020, 99080, 99120, 99110, 99050, 99040, 
    99100, 99160, 99230, 99330, 99450, 99550, 99650, 99720, 99820, 99930, 
    99990, 100080, 100160, 100240, 100310, 100410, 100490, 100540, 100600, 
    100670, 100700, 100750, 100810, 100860, 100930, 101000, 101080, 101150, 
    101210, 101280, 101350, 101380, 101430, 101470, 101500, 101550, 101590, 
    101630, 101700, 101740, 101770, 101790, 101810, 101850, 101870, 101850, 
    101850, 101870, 101890, 101910, 101930, 101930, 101940, 101940, 101930, 
    101910, 101930, 101920, 101920, 101900, 101920, 101940, 101940, 101930, 
    101900, 101890, 101900, 101890, 101870, 101840, 101820, 101820, 101840, 
    101820, 101810, 101830, 101850, 101840, 101850, 101840, 101800, 101790, 
    101800, 101820, 101830, 101850, 101850, 101870, 101880, 101880, 101910, 
    101890, 101900, 101920, 101940, 101970, 102000, 102020, 102060, 102090, 
    102110, 102140, 102170, 102160, 102160, 102170, 102180, 102200, 102230, 
    102240, 102240, 102240, 102240, 102230, 102250, 102240, 102230, 102220, 
    102190, 102190, 102190, 102190, 102170, 102160, 102170, 102160, 102140, 
    102130, 102100, 102040, 102010, 102000, 101980, 101960, 101940, 101930, 
    101910, 101890, 101870, 101840, 101830, 101780, 101750, 101740, 101740, 
    101760, 101730, 101740, 101720, 101690, 101680, 101660, 101620, 101610, 
    101600, 101570, 101570, 101520, 101510, 101560, 101560, 101560, 101550, 
    101500, 101480, 101440, 101390, 101380, 101410, 101370, 101380, 101340, 
    101320, 101280, 101230, 101180, 101120, 101120, 101110, 101090, 101090, 
    101110, 101130, 101080, 101070, 101060, 101060, 101050, 101020, 101000, 
    101020, 101030, 101050, 101110, 101130, 101170, 101170, 101170, 101180, 
    101150, 101140, 101120, 101100, 101080, 101080, 101070, 101060, 101000, 
    100970, 100990, 100910, 100900, 100910, 100910, 100910, 100930, 100950, 
    100950, 100970, 101010, 101000, 101030, 101060, 101080, 101060, 101020, 
    101010, 101020, 101050, 101030, 101010, 101010, 101000, 100970, 100940, 
    100900, 100880, 100880, 100890, 100880, 100830, 100800, 100780, 100780, 
    100760, 100750, 100740, 100720, 100720, 100700, 100700, 100720, 100730, 
    100730, 100740, 100750, 100740, 100730, 100740, 100740, 100730, 100720, 
    100710, 100710, 100700, 100720, 100720, 100730, 100740, 100750, 100730, 
    100730, 100760, 100760, 100750, 100740, 100750, 100760, 100760, 100760, 
    100750, 100750, 100760, 100760, 100750, 100730, 100720, 100740, 100720, 
    100730, 100740, 100760, 100780, 100780, 100780, 100790, 100800, 100810, 
    100830, 100840, 100850, 100860, 100900, 100900, 100930, 100950, 100950, 
    100950, 100960, 100950, 100950, 100950, 100960, 100960, 100970, 100970, 
    100980, 100970, 100960, 100960, 100940, 100910, 100920, 100910, 100900, 
    100910, 100900, 100910, 100890, 100870, 100850, 100800, 100760, 100750, 
    100740, 100710, 100720, 100700, 100700, 100700, 100690, 100660, 100610, 
    100570, 100560, 100520, 100480, 100430, 100410, 100410, 100370, 100380, 
    100380, 100360, 100270, 100200, 100100, 100030, 99990, 99950, 99920, 
    99880, 99890, 99900, 99940, 99930, 99950, 99950, 99940, 99950, 99930, 
    99940, 99950, 99940, 99910, 99880, 99890, 99880, 99880, 99850, 99840, 
    99820, 99830, 99830, 99820, 99820, 99820, 99840, 99870, 99890, 99910, 
    99920, 99930, 99940, 99990, 100040, 100090, 100130, 100180, 100230, 
    100280, 100340, 100410, 100440, 100510, 100540, 100590, 100640, 100690, 
    100750, 100810, 100860, 100920, 100980, 101030, 101070, 101090, 101120, 
    101170, 101240, 101290, 101330, 101380, 101420, 101480, 101540, 101580, 
    101600, 101620, 101640, 101650, 101660, 101700, 101700, 101710, 101720, 
    101740, 101750, 101770, 101770, 101750, 101760, 101770, 101780, 101790, 
    101790, 101800, 101840, 101850, 101850, 101830, 101840, 101820, 101790, 
    101790, 101800, 101810, 101810, 101820, 101820, 101800, 101800, 101810, 
    101800, 101780, 101780, 101770, 101760, 101750, 101770, 101760, 101770, 
    101750, 101740, 101750, 101740, 101710, 101690, 101650, 101650, 101620, 
    101600, 101580, 101560, 101550, 101520, 101480, 101430, 101390, 101350, 
    101330, 101320, 101330, 101350, 101400, 101420, 101430, 101430, 101470, 
    101510, 101550, 101580, 101610, 101640, 101670, 101710, 101730, 101740, 
    101780, 101800, 101830, 101850, 101860, 101870, 101890, 101920, 101930, 
    101980, 102010, 102030, 102040, 102070, 102070, 102080, 102090, 102090, 
    102120, 102130, 102160, 102180, 102210, 102220, 102230, 102250, 102260, 
    102260, 102270, 102260, 102260, 102260, 102280, 102310, 102330, 102350, 
    102340, 102350, 102350, 102350, 102350, 102340, 102330, 102340, 102330, 
    102310, 102310, 102280, 102260, 102260, 102240, 102230, 102210, 102190, 
    102180, 102160, 102150, 102140, 102170, 102180, 102150, 102140, 102130, 
    102140, 102130, 102120, 102090, 102070, 102070, 102080, 102090, 102080, 
    102070, 102060, 102030, 101990, 101970, 101960, 101920, 101890, 101870, 
    101860, 101840, 101810, 101760, 101740, 101690, 101670, 101640, 101590, 
    101560, 101530, 101500, 101490, 101480, 101460, 101450, 101440, 101420, 
    101400, 101420, 101420, 101430, 101420, 101420, 101420, 101430, 101430, 
    101430, 101450, 101440, 101450, 101450, 101470, 101470, 101470, 101480, 
    101500, 101520, 101500, 101460, 101410, 101380, 101340, 101300, 101260, 
    101230, 101170, 101080, 101010, 101020, 101020, 101030, 101050, 101050, 
    101050, 101060, 101060, 101060, 101050, 101040, 101050, 101080, 101100, 
    101110, 101090, 101080, 101060, 101060, 101050, 101070, 101060, 101060, 
    101070, 101090, 101090, 101110, 101150, 101150, 101160, 101160, 101170, 
    101160, 101180, 101190, 101200, 101220, 101240, 101260, 101280, 101290, 
    101300, 101290, 101300, 101310, 101330, 101360, 101370, 101420, 101450, 
    101460, 101470, 101510, 101490, 101490, 101510, 101500, 101480, 101480, 
    101490, 101490, 101490, 101480, 101470, 101470, 101440, 101410, 101380, 
    101370, 101350, 101360, 101370, 101410, 101420, 101400, 101390, 101380, 
    101370, 101350, 101320, 101300, 101280, 101250, 101240, 101230, 101220, 
    101190, 101170, 101140, 101120, 101090, 101060, 101040, 101020, 101010, 
    101030, 101040, 101040, 101010, 100980, 100970, 100950, 100930, 100900, 
    100880, 100860, 100830, 100840, 100820, 100810, 100810, 100800, 100790, 
    100790, 100770, 100740, 100720, 100710, 100700, 100710, 100700, 100710, 
    100710, 100710, 100700, 100680, 100660, 100640, 100620, 100600, 100590, 
    100590, 100570, 100570, 100580, 100570, 100570, 100550, 100520, 100510, 
    100460, 100440, 100440, 100420, 100420, 100420, 100420, 100400, 100380, 
    100360, 100360, 100360, 100350, 100360, 100350, 100360, 100370, 100370, 
    100380, 100380, 100370, 100360, 100360, 100340, 100330, 100320, 100300, 
    100290, 100270, 100250, 100240, 100210, 100180, 100150, 100130, 100100, 
    100070, 100050, 100050, 100040, 100030, 100020, 100010, 100000, 99970, 
    99960, 99950, 99940, 99930, 99920, 99910, 99910, 99920, 99940, 99930, 
    99930, 99920, 99920, 99900, 99900, 99890, 99890, 99910, 99930, 99960, 
    99990, 100020, 100050, 100080, 100080, 100100, 100120, 100190, 100200, 
    100230, 100270, 100290, 100300, 100320, 100320, 100330, 100340, 100320, 
    100350, 100350, 100340, 100340, 100340, 100380, 100370, 100360, 100320, 
    100310, 100290, 100310, 100300, 100300, 100300, 100290, 100290, 100270, 
    100250, 100250, 100250, 100230, 100210, 100190, 100160, 100130, 100120, 
    100130, 100120, 100080, 100090, 100080, 100060, 100050, 100080, 100050, 
    100080, 100080, 100120, 100140, 100190, 100200, 100250, 100270, 100300, 
    100330, 100360, 100390, 100420, 100440, 100470, 100490, 100510, 100530, 
    100550, 100550, 100560, 100560, 100560, 100570, 100610, 100610, 100630, 
    100650, 100670, 100710, 100710, 100730, 100740, 100710, 100720, 100720, 
    100710, 100710, 100700, 100680, 100680, 100660, 100670, 100670, 100640, 
    100620, 100610, 100590, 100560, 100540, 100540, 100520, 100510, 100500, 
    100490, 100490, 100490, 100500, 100500, 100490, 100500, 100520, 100560, 
    100590, 100590, 100620, 100640, 100660, 100680, 100690, 100690, 100710, 
    100700, 100710, 100730, 100740, 100730, 100720, 100720, 100710, 100680, 
    100640, 100610, 100550, 100520, 100480, 100440, 100440, 100400, 100380, 
    100380, 100390, 100430, 100490, 100500, 100580, 100630, 100670, 100710, 
    100760, 100790, 100850, 100910, 100970, 101030, 101090, 101140, 101180, 
    101240, 101280, 101300, 101350, 101390, 101440, 101450, 101460, 101460, 
    101450, 101430, 101430, 101430, 101430, 101430, 101430, 101420, 101420, 
    101420, 101430, 101440, 101440, 101440, 101460, 101490, 101530, 101550, 
    101590, 101590, 101600, 101650, 101670, 101670, 101650, 101650, 101640, 
    101610, 101600, 101620, 101600, 101560, 101510, 101500, 101450, 101380, 
    101290, 101230, 101130, 101000, 100910, 100810, 100740, 100680, 100640, 
    100590, 100550, 100530, 100500, 100480, 100500, 100500, 100520, 100560, 
    100600, 100650, 100720, 100790, 100900, 100970, 101010, 101110, 101180, 
    101220, 101270, 101330, 101360, 101360, 101380, 101340, 101330, 101280, 
    101210, 101110, 101150, 101130, 101110, 101090, 101070, 101070, 101080, 
    101070, 101040, 101040, 101040, 101060, 101100, 101130, 101180, 101250, 
    101290, 101340, 101370, 101390, 101390, 101370, 101340, 101310, 101290, 
    101280, 101280, 101260, 101270, 101250, 101240, 101220, 101190, 101150, 
    101140, 101110, 101070, 101030, 101000, 100960, 100920, 100890, 100840, 
    100790, 100740, 100690, 100600, 100510, 100450, 100380, 100340, 100300, 
    100220, 100180, 100160, 100090, 100070, 100090, 100110, 100100, 100090, 
    100120, 100150, 100170, 100200, 100200, 100180, 100230, 100230, 100240, 
    100280, 100310, 100360, 100380, 100410, 100460, 100530, 100550, 100570, 
    100590, 100630, 100680, 100740, 100740, 100730, 100710, 100730, 100720, 
    100760, 100720, 100700, 100680, 100640, 100590, 100580, 100610, 100620, 
    100640, 100680, 100690, 100750, 100790, 100870, 100960, 101040, 101120, 
    101230, 101330, 101430, 101520, 101600, 101680, 101730, 101790, 101860, 
    101920, 101950, 101980, 101990, 102010, 102030, 102050, 102070, 102080, 
    102060, 102080, 102110, 102100, 102060, 102040, 102020, 102000, 101960, 
    101900, 101800, 101750, 101680, 101630, 101570, 101490, 101420, 101370, 
    101290, 101180, 101080, 101020, 100960, 100870, 100790, 100750, 100670, 
    100590, 100510, 100410, 100310, 100220, 100160, 100110, 100090, 100090, 
    100120, 100190, 100250, 100280, 100330, 100330, 100380, 100420, 100460, 
    100530, 100590, 100640, 100680, 100760, 100830, 100860, 100910, 100950, 
    100980, 100990, 100980, 100970, 100970, 100950, 100970, 100970, 101040, 
    101070, 101080, 101100, 101120, 101090, 101110, 101110, 101100, 101080, 
    101080, 101070, 101050, 101030, 100990, 100930, 100900, 100830, 100780, 
    100730, 100700, 100670, 100620, 100590, 100570, 100530, 100510, 100480, 
    100450, 100410, 100350, 100290, 100210, 100150, 100090, 99990, 99890, 
    99790, 99730, 99670, 99670, 99640, 99610, 99580, 99530, 99450, 99330, 
    99230, 99130, 99060, 99010, 98950, 98890, 98850, 98760, 98680, 98620, 
    98500, 98430, 98330, 98310, 98260, 98170, 98140, 98050, 97970, 97940, 
    97920, 97900, 97900, 97940, 97990, 98060, 98110, 98180, 98230, 98290, 
    98350, 98440, 98510, 98580, 98660, 98750, 98850, 98960, 99050, 99110, 
    99170, 99250, 99310, 99340, 99400, 99440, 99460, 99480, 99520, 99550, 
    99570, 99570, 99550, 99550, 99490, 99460, 99410, 99410, 99370, 99360, 
    99330, 99300, 99270, 99230, 99200, 99150, 99110, 99080, 99050, 99060, 
    99060, 99090, 99090, 99110, 99120, 99120, 99130, 99130, 99130, 99130, 
    99170, 99170, 99190, 99200, 99220, 99250, 99260, 99260, 99240, 99240, 
    99210, 99190, 99170, 99180, 99150, 99140, 99120, 99110, 99110, 99090, 
    99080, 99060, 99080, 99090, 99080, 99080, 99100, 99110, 99100, 99110, 
    99110, 99100, 99120, 99140, 99140, 99160, 99190, 99230, 99270, 99330, 
    99400, 99460, 99520, 99570, 99630, 99690, 99780, 99860, 99930, 99990, 
    100040, 100110, 100180, 100240, 100280, 100350, 100420, 100470, 100500, 
    100540, 100580, 100620, 100650, 100690, 100720, 100750, 100760, 100780, 
    100810, 100830, 100830, 100840, 100840, 100850, 100870, 100860, 100850, 
    100860, 100860, 100870, 100880, 100870, 100860, 100870, 100890, 100900, 
    100900, 100900, 100900, 100910, 100930, 100950, 100970, 100980, 100980, 
    101020, 101030, 101050, 101070, 101100, 101120, 101130, 101160, 101200, 
    101220, 101250, 101270, 101280, 101310, 101340, 101370, 101360, 101360, 
    101360, 101370, 101380, 101410, 101380, 101370, 101370, 101360, 101350, 
    101340, 101320, 101290, 101260, 101230, 101230, 101230, 101200, 101160, 
    101130, 101110, 101070, 101040, 101010, 100990, 100970, 100950, 100930, 
    100900, 100880, 100820, 100780, 100750, 100730, 100690, 100670, 100650, 
    100620, 100600, 100560, 100570, 100560, 100570, 100540, 100550, 100540, 
    100570, 100590, 100620, 100660, 100710, 100760, 100790, 100840, 100890, 
    100920, 100960, 101010, 101040, 101070, 101120, 101170, 101210, 101240, 
    101280, 101320, 101340, 101340, 101390, 101420, 101440, 101480, 101530, 
    101570, 101610, 101630, 101650, 101670, 101660, 101690, 101700, 101700, 
    101720, 101750, 101770, 101790, 101820, 101840, 101850, 101860, 101860, 
    101880, 101900, 101890, 101880, 101920, 101950, 101960, 102000, 102000, 
    101980, 101990, 101990, 101980, 101980, 102030, 102040, 102070, 102080, 
    102080, 102070, 102070, 102070, 102070, 102060, 102050, 102020, 102000, 
    101970, 101970, 101970, 101940, 101900, 101880, 101860, 101840, 101790, 
    101760, 101740, 101720, 101700, 101700, 101690, 101680, 101650, 101640, 
    101620, 101560, 101520, 101510, 101500, 101490, 101500, 101500, 101460, 
    101500, 101460, 101440, 101460, 101480, 101480, 101470, 101470, 101460, 
    101470, 101510, 101530, 101490, 101520, 101540, 101540, 101540, 101550, 
    101540, 101560, 101580, 101620, 101630, 101660, 101670, 101670, 101670, 
    101670, 101680, 101700, 101680, 101690, 101690, 101700, 101720, 101730, 
    101710, 101680, 101660, 101680, 101660, 101620, 101590, 101550, 101510, 
    101480, 101470, 101440, 101400, 101370, 101250, 101170, 101110, 100990, 
    100870, 100750, 100610, 100480, 100400, 100320, 100220, 100110, 99990, 
    99870, 99800, 99720, 99630, 99520, 99420, 99300, 99220, 99160, 99110, 
    99080, 99090, 99100, 99110, 99130, 99160, 99190, 99260, 99270, 99340, 
    99430, 99550, 99620, 99710, 99830, 99940, 100080, 100210, 100290, 100380, 
    100460, 100580, 100690, 100800, 100880, 100950, 100990, 101070, 101140, 
    101230, 101280, 101330, 101400, 101480, 101530, 101580, 101630, 101670, 
    101690, 101720, 101750, 101770, 101790, 101830, 101830, 101860, 101860, 
    101860, 101850, 101840, 101810, 101820, 101820, 101820, 101800, 101770, 
    101740, 101710, 101690, 101640, 101600, 101530, 101410, 101390, 101370, 
    101320, 101230, 101130, 101050, 100980, 100890, 100810, 100770, 100720, 
    100640, 100600, 100500, 100500, 100460, 100430, 100420, 100410, 100410, 
    100430, 100460, 100480, 100480, 100480, 100480, 100470, 100450, 100400, 
    100310, 100210, 100120, 100020, 99880, 99710, 99540, 99390, 99190, 99070, 
    99000, 98890, 98820, 98870, 98970, 99030, 99120, 99310, 99410, 99570, 
    99760, 100020, 100160, 100250, 100270, 100390, 100450, 100510, 100570, 
    100600, 100610, 100620, 100630, 100660, 100680, 100710, 100760, 100830, 
    100890, 100970, 101040, 101080, 101110, 101150, 101160, 101200, 101220, 
    101220, 101230, 101240, 101280, 101320, 101310, 101320, 101310, 101330, 
    101350, 101390, 101420, 101470, 101530, 101570, 101560, 101560, 101510, 
    101470, 101380, 101300, 101140, 100970, 100770, 100670, 100640, 100710, 
    100790, 100830, 100860, 100840, 100880, 100910, 100930, 100960, 101010, 
    101110, 101170, 101180, 101210, 101240, 101260, 101250, 101200, 101150, 
    101090, 101050, 101060, 101060, 101090, 101140, 101180, 101210, 101270, 
    101330, 101420, 101500, 101560, 101620, 101680, 101740, 101770, 101840, 
    101880, 101910, 101940, 101910, 101910, 101900, 101860, 101860, 101800, 
    101760, 101750, 101710, 101680, 101660, 101660, 101640, 101640, 101650, 
    101650, 101640, 101650, 101670, 101700, 101700, 101690, 101680, 101670, 
    101670, 101640, 101630, 101640, 101650, 101650, 101670, 101680, 101700, 
    101710, 101710, 101720, 101720, 101700, 101670, 101650, 101630, 101620, 
    101620, 101620, 101620, 101640, 101650, 101650, 101650, 101630, 101640, 
    101640, 101640, 101650, 101650, 101680, 101700, 101710, 101710, 101740, 
    101740, 101740, 101760, 101790, 101820, 101840, 101850, 101850, 101880, 
    101900, 101920, 101930, 101930, 101920, 101950, 101940, 101930, 101920, 
    101920, 101940, 101940, 101940, 101920, 101880, 101830, 101770, 101720, 
    101690, 101640, 101580, 101520, 101440, 101370, 101300, 101220, 101110, 
    101040, 100970, 100860, 100790, 100760, 100720, 100700, 100690, 100710, 
    100720, 100740, 100720, 100710, 100710, 100680, 100660, 100620, 100600, 
    100550, 100560, 100560, 100540, 100510, 100470, 100440, 100410, 100390, 
    100380, 100360, 100330, 100330, 100340, 100350, 100370, 100360, 100360, 
    100350, 100350, 100350, 100350, 100360, 100330, 100310, 100340, 100360, 
    100340, 100310, 100320, 100320, 100290, 100260, 100240, 100230, 100210, 
    100170, 100150, 100130, 100090, 100040, 100010, 99970, 99910, 99830, 
    99770, 99740, 99660, 99600, 99520, 99430, 99390, 99310, 99210, 99150, 
    99100, 99060, 99010, 98930, 98900, 98840, 98840, 98820, 98840, 98840, 
    98870, 98860, 98900, 98890, 98900, 98920, 98930, 98930, 98970, 98980, 
    98980, 99020, 99040, 98990, 98990, 99010, 99000, 98980, 98950, 98960, 
    98980, 98960, 98970, 98950, 98950, 98910, 98940, 98930, 98960, 99000, 
    99050, 99100, 99110, 99130, 99120, 99160, 99180, 99190, 99190, 99220, 
    99230, 99260, 99290, 99340, 99420, 99480, 99530, 99580, 99640, 99690, 
    99750, 99810, 99880, 99940, 100000, 100060, 100140, 100240, 100330, 
    100420, 100510, 100610, 100700, 100800, 100910, 101020, 101120, 101200, 
    101290, 101370, 101420, 101430, 101430, 101400, 101390, 101450, 101460, 
    101510, 101580, 101660, 101710, 101860, 102000, 102130, 102250, 102360, 
    102410, 102410, 102440, 102450, 102410, 102370, 102350, 102320, 102270, 
    102210, 102120, 102010, 101950, 101890, 101860, 101820, 101820, 101760, 
    101690, 101600, 101510, 101460, 101390, 101290, 101180, 101050, 100900, 
    100730, 100630, 100570, 100510, 100490, 100510, 100530, 100580, 100620, 
    100620, 100630, 100690, 100790, 100870, 100990, 101110, 101230, 101360, 
    101500, 101620, 101750, 101890, 102050, 102210, 102280, 102350, 102470, 
    102550, 102590, 102680, 102740, 102740, 102740, 102770, 102750, 102750, 
    102710, 102690, 102630, 102520, 102430, 102310, 102210, 102080, 101950, 
    101830, 101690, 101560, 101480, 101340, 101200, 101130, 101070, 101010, 
    100980, 101010, 101180, 101220, 101260, 101290, 101240, 101230, 101230, 
    101390, 101450, 101630, 101740, 101870, 101960, 102080, 102160, 102250, 
    102330, 102390, 102440, 102470, 102500, 102540, 102590, 102650, 102660, 
    102680, 102710, 102740, 102760, 102790, 102830, 102860, 102880, 102900, 
    102920, 102940, 102960, 102950, 102970, 102950, 102930, 102890, 102890, 
    102870, 102860, 102820, 102780, 102730, 102680, 102620, 102580, 102540, 
    102480, 102460, 102420, 102380, 102320, 102300, 102210, 102170, 102130, 
    102090, 102010, 101950, 101930, 101860, 101850, 101820, 101830, 101830, 
    101820, 101790, 101790, 101800, 101770, 101770, 101780, 101780, 101770, 
    101760, 101750, 101740, 101710, 101670, 101620, 101560, 101500, 101420, 
    101330, 101240, 101200, 101130, 101080, 100980, 100890, 100800, 100750, 
    100720, 100730, 100740, 100760, 100800, 100870, 100930, 100980, 101040, 
    101100, 101150, 101200, 101260, 101280, 101310, 101340, 101380, 101420, 
    101480, 101530, 101570, 101600, 101630, 101650, 101660, 101680, 101680, 
    101710, 101730, 101760, 101790, 101810, 101830, 101840, 101870, 101900, 
    101920, 101950, 101980, 101970, 102000, 102040, 102070, 102090, 102110, 
    102150, 102150, 102180, 102220, 102220, 102220, 102220, 102250, 102240, 
    102240, 102240, 102230, 102250, 102230, 102190, 102120, 102070, 101970, 
    101890, 101810, 101720, 101620, 101510, 101430, 101350, 101290, 101200, 
    101120, 101080, 101010, 100920, 100870, 100830, 100760, 100680, 100660, 
    100600, 100540, 100500, 100430, 100360, 100270, 100170, 100090, 100050, 
    100030, 100110, 100140, 100200, 100180, 100170, 100300, 100430, 100510, 
    100500, 100550, 100620, 100650, 100740, 100840, 100880, 100950, 100960, 
    101100, 101200, 101280, 101360, 101430, 101470, 101500, 101560, 101600, 
    101640, 101650, 101660, 101640, 101660, 101630, 101610, 101590, 101550, 
    101550, 101530, 101530, 101540, 101570, 101580, 101580, 101560, 101570, 
    101600, 101600, 101610, 101610, 101630, 101620, 101630, 101640, 101640, 
    101640, 101630, 101620, 101610, 101600, 101580, 101580, 101600, 101620, 
    101630, 101620, 101600, 101600, 101600, 101600, 101630, 101630, 101630, 
    101660, 101680, 101690, 101690, 101680, 101650, 101660, 101660, 101640, 
    101640, 101660, 101640, 101620, 101620, 101630, 101630, 101630, 101630, 
    101610, 101590, 101580, 101570, 101550, 101540, 101530, 101540, 101540, 
    101540, 101530, 101500, 101490, 101470, 101470, 101460, 101450, 101440, 
    101460, 101450, 101450, 101420, 101440, 101460, 101410, 101400, 101410, 
    101410, 101390, 101390, 101410, 101440, 101480, 101510, 101520, 101490, 
    101450, 101420, 101390, 101370, 101360, 101320, 101280, 101240, 101140, 
    101130, 100990, 100960, 100930, 100880, 100830, 100820, 100790, 100810, 
    100820, 100920, 100950, 101020, 101050, 101090, 101170, 101220, 101340, 
    101420, 101500, 101550, 101650, 101730, 101790, 101830, 101830, 101820, 
    101860, 101860, 101840, 101850, 101850, 101910, 101950, 102040, 102120, 
    102220, 102300, 102380, 102450, 102530, 102610, 102660, 102700, 102710, 
    102760, 102790, 102800, 102800, 102790, 102790, 102790, 102800, 102780, 
    102800, 102810, 102850, 102850, 102860, 102840, 102890, 102910, 102890, 
    102880, 102900, 102900, 102900, 102890, 102920, 102960, 102940, 102970, 
    102970, 102940, 102930, 102890, 102860, 102830, 102800, 102760, 102730, 
    102720, 102710, 102690, 102680, 102620, 102570, 102540, 102480, 102420, 
    102350, 102290, 102230, 102150, 102070, 102010, 101950, 101880, 101820, 
    101750, 101680, 101600, 101530, 101470, 101410, 101360, 101320, 101280, 
    101240, 101210, 101170, 101130, 101090, 101070, 101040, 101030, 101040, 
    101030, 101040, 101030, 101010, 100980, 100960, 100920, 100910, 100900, 
    100900, 100880, 100890, 100890, 100870, 100860, 100840, 100840, 100830, 
    100800, 100770, 100740, 100700, 100660, 100660, 100670, 100690, 100710, 
    100720, 100740, 100740, 100730, 100750, 100760, 100780, 100800, 100820, 
    100870, 100910, 100930, 100940, 100970, 100990, 100970, 100960, 100970, 
    100950, 100920, 100910, 100910, 100930, 100950, 100950, 100950, 100970, 
    101000, 101020, 101030, 101060, 101080, 101110, 101150, 101210, 101260, 
    101250, 101310, 101330, 101340, 101400, 101460, 101540, 101570, 101690, 
    101730, 101760, 101800, 101840, 101870, 101890, 101950, 101990, 102100, 
    102140, 102200, 102260, 102330, 102400, 102450, 102540, 102620, 102670, 
    102710, 102760, 102780, 102810, 102820, 102860, 102900, 102930, 102960, 
    102990, 103040, 103080, 103110, 103130, 103150, 103170, 103200, 103220, 
    103230, 103270, 103280, 103300, 103310, 103320, 103340, 103340, 103340, 
    103330, 103310, 103320, 103340, 103350, 103360, 103340, 103330, 103320, 
    103300, 103280, 103250, 103220, 103210, 103200, 103210, 103210, 103210, 
    103210, 103200, 103200, 103210, 103190, 103180, 103190, 103190, 103220, 
    103220, 103230, 103230, 103240, 103230, 103220, 103200, 103190, 103180, 
    103190, 103180, 103150, 103160, 103160, 103150, 103140, 103110, 103090, 
    103050, 103020, 102990, 102960, 102920, 102890, 102860, 102830, 102810, 
    102790, 102760, 102720, 102700, 102680, 102670, 102640, 102610, 102610, 
    102610, 102590, 102620, 102630, 102630, 102630, 102640, 102660, 102680, 
    102690, 102680, 102690, 102730, 102740, 102750, 102760, 102780, 102800, 
    102810, 102820, 102830, 102840, 102840, 102860, 102870, 102900, 102920, 
    102940, 102940, 102940, 102940, 102940, 102960, 102960, 102970, 102970, 
    102980, 102960, 102960, 102960, 102940, 102910, 102890, 102870, 102830, 
    102820, 102770, 102720, 102690, 102640, 102620, 102580, 102530, 102490, 
    102440, 102390, 102340, 102300, 102260, 102220, 102200, 102190, 102170, 
    102160, 102160, 102150, 102160, 102170, 102180, 102210, 102240, 102260, 
    102280, 102320, 102330, 102330, 102340, 102350, 102340, 102340, 102330, 
    102330, 102310, 102260, 102230, 102200, 102140, 102080, 102000, 101910, 
    101850, 101790, 101720, 101650, 101560, 101510, 101470, 101420, 101360, 
    101300, 101230, 101170, 101080, 101020, 100930, 100880, 100800, 100730, 
    100660, 100590, 100500, 100430, 100350, 100280, 100180, 100120, 100050, 
    99960, 99870, 99790, 99700, 99650, 99580, 99530, 99460, 99390, 99310, 
    99200, 99130, 99040, 98990, 98910, 98880, 98750, 98670, 98610, 98510, 
    98440, 98390, 98380, 98380, 98450, 98590, 98730, 98940, 99120, 99230, 
    99380, 99580, 99730, 99800, 99920, 100050, 100100, 100180, 100240, 
    100280, 100340, 100340, 100370, 100400, 100430, 100460, 100510, 100580, 
    100620, 100660, 100720, 100780, 100880, 100970, 101070, 101180, 101240, 
    101250, 101350, 101420, 101470, 101520, 101560, 101600, 101660, 101710, 
    101770, 101770, 101810, 101830, 101840, 101870, 101900, 101920, 101970, 
    102020, 102050, 102110, 102130, 102150, 102170, 102200, 102210, 102210, 
    102210, 102200, 102180, 102160, 102140, 102130, 102130, 102100, 102060, 
    101990, 101970, 101920, 101890, 101840, 101790, 101800, 101790, 101770, 
    101740, 101720, 101670, 101610, 101620, 101580, 101560, 101500, 101470, 
    101450, 101410, 101390, 101370, 101340, 101260, 101210, 101170, 101120, 
    101090, 101020, 100960, 100950, 100930, 100900, 100870, 100830, 100780, 
    100760, 100740, 100740, 100710, 100700, 100690, 100690, 100640, 100610, 
    100600, 100570, 100550, 100520, 100500, 100460, 100420, 100380, 100360, 
    100330, 100320, 100290, 100260, 100260, 100230, 100180, 100180, 100160, 
    100120, 100080, 100030, 99970, 99910, 99850, 99760, 99640, 99560, 99460, 
    99400, 99250, 99190, 99100, 98980, 98840, 98640, 98370, 98170, 97950, 
    97740, 97570, 97390, 97260, 97200, 97150, 97100, 96950, 96910, 96890, 
    96920, 96980, 97100, 97200, 97300, 97390, 97480, 97480, 97550, 97600, 
    97660, 97720, 97830, 97920, 98010, 98120, 98210, 98280, 98370, 98390, 
    98440, 98500, 98510, 98540, 98520, 98510, 98470, 98430, 98340, 98220, 
    98070, 97990, 97910, 97840, 97800, 97760, 97690, 97630, 97560, 97540, 
    97450, 97390, 97380, 97400, 97430, 97510, 97870, 97870, 98130, 98380, 
    98640, 98880, 99080, 99260, 99380, 99540, 99690, 99760, 99880, 100000, 
    100100, 100160, 100250, 100360, 100470, 100580, 100650, 100740, 100820, 
    100910, 101000, 101100, 101170, 101230, 101290, 101340, 101370, 101400, 
    101420, 101460, 101480, 101500, 101500, 101520, 101530, 101530, 101520, 
    101500, 101490, 101480, 101470, 101470, 101460, 101430, 101380, 101360, 
    101340, 101340, 101330, 101330, 101260, 101210, 101170, 101120, 101080, 
    101030, 100980, 100910, 100900, 100880, 100840, 100820, 100800, 100760, 
    100710, 100650, 100610, 100580, 100530, 100490, 100440, 100410, 100370, 
    100350, 100330, 100330, 100300, 100300, 100300, 100320, 100330, 100350, 
    100340, 100330, 100350, 100330, 100340, 100360, 100380, 100450, 100480, 
    100520, 100550, 100610, 100650, 100670, 100690, 100700, 100740, 100740, 
    100810, 100840, 100870, 100910, 100960, 101010, 101070, 101100, 101150, 
    101170, 101200, 101230, 101290, 101310, 101340, 101380, 101400, 101430, 
    101430, 101430, 101440, 101450, 101460, 101470, 101480, 101500, 101500, 
    101540, 101580, 101590, 101600, 101630, 101650, 101640, 101640, 101640, 
    101640, 101650, 101670, 101700, 101700, 101700, 101660, 101660, 101670, 
    101660, 101660, 101660, 101670, 101670, 101670, 101660, 101680, 101710, 
    101710, 101720, 101720, 101700, 101720, 101710, 101700, 101710, 101720, 
    101740, 101740, 101740, 101740, 101770, 101780, 101770, 101760, 101750, 
    101750, 101770, 101760, 101780, 101810, 101840, 101880, 101900, 101890, 
    101890, 101900, 101900, 101890, 101880, 101880, 101890, 101890, 101900, 
    101890, 101890, 101860, 101820, 101800, 101780, 101740, 101710, 101690, 
    101660, 101630, 101630, 101610, 101590, 101540, 101510, 101470, 101460, 
    101450, 101430, 101450, 101470, 101520, 101550, 101530, 101500, 101480, 
    101510, 101510, 101510, 101540, 101540, 101550, 101550, 101560, 101580, 
    101600, 101580, 101570, 101600, 101590, 101600, 101620, 101620, 101640, 
    101680, 101690, 101690, 101710, 101750, 101760, 101780, 101770, 101850, 
    101890, 101900, 101940, 101960, 101980, 101990, 102020, 102040, 102050, 
    102030, 102020, 102000, 101990, 101980, 101960, 101940, 101930, 101900, 
    101860, 101800, 101730, 101680, 101620, 101570, 101520, 101450, 101380, 
    101330, 101270, 101230, 101170, 101110, 101060, 100980, 100930, 100870, 
    100790, 100740, 100710, 100690, 100670, 100660, 100640, 100610, 100580, 
    100530, 100500, 100460, 100450, 100410, 100390, 100360, 100330, 100360, 
    100420, 100460, 100460, 100490, 100510, 100490, 100540, 100560, 100590, 
    100610, 100640, 100640, 100650, 100670, 100640, 100670, 100730, 100780, 
    100850, 100860, 100880, 100890, 100930, 100990, 101010, 101040, 101100, 
    101110, 101130, 101170, 101200, 101230, 101230, 101260, 101290, 101330, 
    101380, 101420, 101420, 101440, 101480, 101500, 101540, 101560, 101570, 
    101610, 101650, 101680, 101710, 101760, 101800, 101820, 101840, 101850, 
    101880, 101900, 101930, 101970, 101980, 102000, 102000, 101990, 101990, 
    101990, 101980, 101980, 101960, 101920, 101910, 101890, 101870, 101850, 
    101820, 101800, 101760, 101720, 101670, 101630, 101600, 101550, 101510, 
    101450, 101410, 101370, 101320, 101260, 101200, 101140, 101100, 101060, 
    101030, 100990, 100960, 100970, 100960, 100980, 100960, 100930, 100920, 
    100890, 100860, 100830, 100810, 100760, 100710, 100720, 100680, 100630, 
    100590, 100550, 100490, 100420, 100380, 100330, 100300, 100280, 100250, 
    100210, 100160, 100130, 100090, 100040, 99980, 99910, 99850, 99870, 
    99850, 99890, 99920, 99940, 99990, 100070, 100140, 100160, 100220, 
    100280, 100340, 100370, 100420, 100440, 100460, 100480, 100510, 100580, 
    100620, 100700, 100770, 100900, 101010, 101090, 101150, 101220, 101320, 
    101350, 101370, 101370, 101410, 101430, 101440, 101410, 101400, 101370, 
    101340, 101310, 101290, 101270, 101240, 101200, 101180, 101140, 101090, 
    101050, 101020, 100990, 100960, 100940, 100910, 100900, 100890, 100910, 
    100930, 100920, 100920, 100910, 100890, 100890, 100890, 100890, 100880, 
    100890, 100860, 100880, 100870, 100850, 100830, 100780, 100760, 100740, 
    100690, 100660, 100610, 100550, 100510, 100480, 100450, 100390, 100340, 
    100310, 100260, 100180, 100110, 100040, 99990, 99960, 99950, 99920, 
    99970, 100010, 100040, 100070, 100100, 100140, 100210, 100260, 100280, 
    100330, 100390, 100470, 100510, 100540, 100630, 100710, 100740, 100810, 
    100850, 100860, 100910, 101000, 101060, 101120, 101200, 101290, 101350, 
    101410, 101470, 101520, 101530, 101570, 101580, 101620, 101650, 101670, 
    101720, 101740, 101740, 101780, 101780, 101780, 101760, 101770, 101780, 
    101780, 101790, 101820, 101810, 101780, 101780, 101740, 101700, 101670, 
    101630, 101590, 101550, 101530, 101480, 101450, 101400, 101350, 101300, 
    101250, 101210, 101160, 101100, 101040, 101000, 100980, 100950, 100930, 
    100930, 100900, 100890, 100880, 100880, 100850, 100820, 100780, 100780, 
    100760, 100730, 100720, 100730, 100710, 100710, 100730, 100700, 100700, 
    100680, 100640, 100620, 100650, 100660, 100670, 100650, 100680, 100680, 
    100680, 100650, 100640, 100640, 100650, 100670, 100690, 100720, 100740, 
    100770, 100790, 100800, 100790, 100810, 100800, 100800, 100790, 100800, 
    100830, 100820, 100820, 100820, 100830, 100820, 100850, 100860, 100860, 
    100850, 100850, 100860, 100890, 100890, 100880, 100870, 100810, 100780, 
    100750, 100720, 100700, 100680, 100660, 100630, 100620, 100620, 100610, 
    100580, 100570, 100550, 100520, 100510, 100480, 100450, 100410, 100370, 
    100360, 100330, 100270, 100240, 100220, 100180, 100160, 100130, 100130, 
    100080, 100080, 100070, 100080, 100110, 100150, 100150, 100130, 100100, 
    100080, 100060, 100030, 99960, 99860, 99820, 99780, 99750, 99700, 99640, 
    99590, 99530, 99500, 99480, 99450, 99420, 99420, 99440, 99490, 99540, 
    99620, 99700, 99750, 99840, 99940, 100000, 100040, 100070, 100090, 
    100140, 100200, 100240, 100220, 100170, 100200, 100130, 100070, 100040, 
    100000, 99960, 99900, 99840, 99800, 99750, 99710, 99670, 99630, 99610, 
    99580, 99540, 99500, 99470, 99440, 99410, 99380, 99360, 99330, 99300, 
    99290, 99290, 99290, 99290, 99290, 99280, 99290, 99290, 99310, 99310, 
    99330, 99340, 99350, 99390, 99420, 99440, 99450, 99470, 99490, 99540, 
    99620, 99680, 99760, 99800, 99820, 99850, 99900, 99810, 99780, 99710, 
    99670, 99590, 99460, 99310, 99170, 98900, 98690, 98450, 98110, 97870, 
    97600, 97320, 97060, 96830, 96620, 96530, 96630, 96640, 96700, 96750, 
    96800, 96860, 96910, 96980, 97010, 97100, 97260, 97430, 97530, 97610, 
    97740, 97880, 97990, 98100, 98150, 98140, 98150, 98150, 98140, 98130, 
    98110, 98080, 98060, 97990, 97850, 97660, 97460, 97160, 96880, 96640, 
    96500, 96480, 96510, 96440, 96420, 96450, 96500, 96490, 96500, 96490, 
    96370, 96330, 96320, 96370, 96430, 96460, 96540, 96560, 96600, 96650, 
    96660, 96700, 96670, 96660, 96680, 96700, 96670, 96760, 96800, 96830, 
    96850, 96850, 96840, 96840, 96810, 96780, 96830, 96820, 96820, 96850, 
    96870, 96850, 96840, 96870, 96900, 96920, 96940, 96980, 97010, 97080, 
    97130, 97160, 97230, 97260, 97290, 97320, 97380, 97410, 97450, 97470, 
    97510, 97530, 97550, 97570, 97590, 97580, 97580, 97580, 97590, 97600, 
    97610, 97620, 97630, 97700, 97740, 97760, 97780, 97790, 97840, 97890, 
    97920, 97930, 97950, 97980, 98000, 98030, 98070, 98100, 98140, 98150, 
    98180, 98190, 98210, 98210, 98230, 98250, 98250, 98270, 98280, 98320, 
    98340, 98320, 98310, 98300, 98300, 98280, 98230, 98200, 98150, 98140, 
    98150, 98110, 98070, 98050, 98030, 97990, 97950, 97920, 97900, 97890, 
    97900, 97890, 97920, 97990, 98010, 98010, 97990, 97990, 98030, 98040, 
    98150, 98270, 98390, 98530, 98690, 98850, 98970, 99090, 99230, 99370, 
    99460, 99600, 99740, 99880, 99950, 100080, 100250, 100350, 100470, 
    100550, 100630, 100750, 100830, 100880, 100910, 100940, 101000, 101070, 
    101120, 101190, 101240, 101250, 101260, 101290, 101280, 101270, 101260, 
    101190, 101100, 100970, 100810, 100640, 100450, 100290, 100070, 99780, 
    99570, 99350, 99150, 98910, 98710, 98540, 98390, 98320, 98240, 98240, 
    98150, 98220, 98200, 98310, 98380, 98490, 98600, 98730, 98850, 98950, 
    99020, 99110, 99190, 99220, 99290, 99420, 99460, 99590, 99700, 99780, 
    99890, 99960, 100040, 100080, 100110, 100130, 100170, 100180, 100130, 
    100100, 100130, 100140, 100200, 100260, 100250, 100260, 100250, 100280, 
    100230, 100270, 100330, 100380, 100440, 100520, 100550, 100590, 100640, 
    100650, 100680, 100730, 100790, 100830, 100860, 100920, 101000, 101070, 
    101140, 101240, 101310, 101400, 101490, 101600, 101660, 101710, 101770, 
    101800, 101910, 101970, 102050, 102130, 102140, 102170, 102190, 102210, 
    102220, 102250, 102260, 102260, 102240, 102260, 102300, 102300, 102300, 
    102280, 102250, 102240, 102250, 102250, 102260, 102240, 102260, 102250, 
    102250, 102220, 102190, 102150, 102130, 102100, 102060, 102010, 101950, 
    101930, 101910, 101890, 101890, 101850, 101820, 101770, 101730, 101710, 
    101660, 101640, 101610, 101570, 101570, 101530, 101540, 101540, 101530, 
    101520, 101560, 101570, 101570, 101570, 101590, 101610, 101650, 101700, 
    101720, 101730, 101770, 101800, 101820, 101830, 101800, 101840, 101830, 
    101810, 101820, 101860, 101870, 101860, 101870, 101850, 101800, 101760, 
    101740, 101700, 101660, 101610, 101590, 101510, 101420, 101380, 101290, 
    101210, 101120, 101080, 101040, 100970, 100940, 100910, 100890, 100870, 
    100900, 100860, 100800, 100720, 100630, 100510, 100360, 100170, 99960, 
    99790, 99700, 99570, 99420, 99250, 99110, 99000, 98860, 98790, 98740, 
    98810, 98880, 98850, 98840, 98920, 98980, 98990, 99030, 99070, 99080, 
    99100, 99150, 99160, 99140, 99130, 99130, 99100, 99050, 99000, 98890, 
    98800, 98690, 98610, 98580, 98460, 98480, 98500, 98510, 98490, 98580, 
    98620, 98660, 98700, 98720, 98760, 98790, 98780, 98870, 98910, 98950, 
    99000, 99020, 99060, 99080, 99100, 99110, 99170, 99200, 99210, 99240, 
    99290, 99380, 99400, 99430, 99430, 99430, 99430, 99440, 99440, 99420, 
    99390, 99350, 99350, 99350, 99350, 99350, 99350, 99330, 99310, 99310, 
    99300, 99280, 99290, 99320, 99330, 99330, 99380, 99400, 99410, 99440, 
    99480, 99500, 99460, 99500, 99530, 99560, 99570, 99580, 99610, 99640, 
    99660, 99650, 99690, 99700, 99720, 99700, 99710, 99700, 99700, 99690, 
    99720, 99710, 99690, 99700, 99680, 99690, 99690, 99680, 99660, 99620, 
    99620, 99580, 99580, 99600, 99590, 99550, 99500, 99480, 99430, 99380, 
    99330, 99320, 99260, 99250, 99210, 99170, 99130, 99100, 99040, 98990, 
    98950, 98880, 98830, 98770, 98720, 98660, 98650, 98610, 98580, 98540, 
    98520, 98520, 98540, 98550, 98540, 98560, 98600, 98620, 98660, 98720, 
    98760, 98800, 98870, 98890, 98940, 98980, 99020, 99060, 99070, 99110, 
    99160, 99210, 99270, 99300, 99310, 99330, 99350, 99330, 99320, 99350, 
    99370, 99410, 99440, 99480, 99490, 99530, 99540, 99540, 99550, 99550, 
    99540, 99540, 99530, 99540, 99570, 99590, 99610, 99600, 99610, 99620, 
    99600, 99620, 99620, 99620, 99620, 99620, 99620, 99620, 99620, 99630, 
    99630, 99650, 99600, 99590, 99570, 99540, 99540, 99560, 99590, 99620, 
    99640, 99640, 99640, 99660, 99680, 99710, 99730, 99740, 99760, 99790, 
    99830, 99890, 99900, 99930, 99950, 99990, 100050, 100080, 100100, 100130, 
    100180, 100230, 100260, 100300, 100340, 100380, 100430, 100480, 100540, 
    100550, 100540, 100560, 100570, 100590, 100560, 100610, 100630, 100610, 
    100570, 100490, 100410, 100330, 100230, 100070, 99900, 99730, 99530, 
    99310, 99070, 98810, 98580, 98350, 98140, 97970, 97800, 97780, 97760, 
    97690, 97740, 97700, 97670, 97610, 97540, 97430, 97340, 97270, 97160, 
    97120, 96910, 96890, 96980, 96990, 96980, 96910, 96930, 96880, 97010, 
    97030, 97060, 97150, 97270, 97450, 97630, 97860, 98090, 98300, 98440, 
    98550, 98570, 98610, 98640, 98630, 98590, 98520, 98460, 98400, 98380, 
    98370, 98350, 98350, 98330, 98340, 98370, 98420, 98410, 98370, 98400, 
    98360, 98310, 98270, 98220, 98150, 98060, 98010, 97950, 97890, 97840, 
    97820, 97830, 97860, 97890, 97930, 97970, 98000, 98060, 98150, 98160, 
    98180, 98220, 98260, 98320, 98360, 98440, 98450, 98470, 98500, 98530, 
    98530, 98510, 98500, 98560, 98580, 98670, 98770, 98860, 98940, 98980, 
    99050, 99120, 99150, 99210, 99280, 99360, 99410, 99530, 99670, 99800, 
    99870, 99930, 99960, 99970, 99990, 99930, 100020, 100130, 100200, 100280, 
    100400, 100420, 100490, 100580, 100680, 100780, 100900, 100950, 101080, 
    101140, 101200, 101210, 101270, 101330, 101370, 101400, 101410, 101420, 
    101440, 101440, 101420, 101400, 101420, 101440, 101450, 101410, 101410, 
    101390, 101370, 101350, 101320, 101320, 101290, 101260, 101250, 101250, 
    101230, 101200, 101170, 101150, 101110, 101080, 101070, 101030, 101000, 
    100970, 100950, 100940, 100930, 100890, 100850, 100830, 100790, 100730, 
    100680, 100650, 100580, 100510, 100430, 100390, 100330, 100310, 100260, 
    100190, 100070, 99990, 99900, 99810, 99710, 99600, 99480, 99390, 99270, 
    99120, 99000, 98910, 98750, 98620, 98490, 98390, 98330, 98330, 98360, 
    98390, 98410, 98430, 98430, 98430, 98410, 98380, 98380, 98370, 98330, 
    98310, 98270, 98290, 98350, 98370, 98360, 98380, 98430, 98480, 98510, 
    98560, 98660, 98730, 98850, 98960, 99090, 99270, 99410, 99570, 99730, 
    99860, 100030, 100160, 100340, 100490, 100610, 100760, 100880, 100960, 
    101080, 101160, 101210, 101260, 101270, 101280, 101290, 101300, 101320, 
    101320, 101330, 101340, 101310, 101270, 101260, 101180, 101160, 101090, 
    101050, 100980, 100960, 100920, 100860, 100790, 100680, 100600, 100490, 
    100410, 100370, 100310, 100250, 100240, 100250, 100340, 100420, 100470, 
    100540, 100620, 100690, 100750, 100810, 100820, 100850, 100880, 100900, 
    100920, 100930, 100920, 100900, 100910, 100930, 100920, 100930, 100900, 
    100890, 100880, 100910, 100930, 100950, 100940, 100920, 100860, 100830, 
    100760, 100660, 100650, 100580, 100490, 100440, 100420, 100370, 100330, 
    100290, 100240, 100190, 100100, 100060, 100070, 100090, 100080, 100070, 
    100090, 100120, 100110, 100110, 100110, 100120, 100140, 100160, 100180, 
    100220, 100290, 100330, 100370, 100440, 100460, 100500, 100540, 100580, 
    100620, 100700, 100760, 100790, 100900, 100950, 100930, 101010, 101060, 
    101100, 101100, 101130, 101170, 101230, 101340, 101400, 101420, 101470, 
    101560, 101660, 101740, 101790, 101860, 101910, 102010, 102050, 102080, 
    102100, 102150, 102180, 102230, 102270, 102300, 102300, 102280, 102290, 
    102290, 102300, 102270, 102250, 102210, 102210, 102200, 102170, 102130, 
    102080, 102030, 101970, 101900, 101820, 101740, 101680, 101610, 101530, 
    101450, 101380, 101300, 101240, 101190, 101110, 101080, 101030, 100970, 
    100920, 100850, 100830, 100800, 100820, 100810, 100780, 100740, 100730, 
    100720, 100690, 100640, 100620, 100610, 100580, 100570, 100560, 100530, 
    100500, 100470, 100450, 100440, 100420, 100390, 100340, 100310, 100280, 
    100270, 100240, 100210, 100180, 100170, 100150, 100100, 100080, 100030, 
    100000, 99980, 99980, 99990, 100000, 100020, 100050, 100090, 100140, 
    100190, 100240, 100300, 100340, 100450, 100520, 100610, 100700, 100730, 
    100760, 100770, 100810, 100820, 100780, 100780, 100740, 100680, 100650, 
    100650, 100610, 100620, 100620, 100650, 100650, 100630, 100600, 100580, 
    100590, 100570, 100560, 100590, 100640, 100670, 100680, 100640, 100620, 
    100630, 100660, 100680, 100690, 100730, 100730, 100770, 100780, 100830, 
    100860, 100870, 100920, 100930, 101020, 101080, 101120, 101150, 101200, 
    101260, 101330, 101410, 101430, 101480, 101530, 101590, 101600, 101640, 
    101650, 101660, 101630, 101620, 101600, 101580, 101540, 101480, 101440, 
    101430, 101430, 101420, 101400, 101390, 101450, 101540, 101610, 101660, 
    101730, 101780, 101770, 101830, 101860, 101900, 101970, 102050, 102140, 
    102190, 102210, 102280, 102430, 102500, 102540, 102540, 102600, 102600, 
    102680, 102700, 102810, 102870, 102930, 102960, 102990, 103030, 103000, 
    102950, 102940, 102970, 103000, 103020, 103020, 103060, 103080, 103120, 
    103150, 103150, 103180, 103230, 103230, 103200, 103200, 103190, 103230, 
    103210, 103220, 103190, 103240, 103290, 103280, 103290, 103280, 103320, 
    103310, 103330, 103350, 103330, 103310, 103280, 103230, 103220, 103190, 
    103140, 103080, 103050, 102990, 102910, 102850, 102820, 102750, 102680, 
    102600, 102470, 102350, 102220, 102100, 101990, 101860, 101700, 101580, 
    101460, 101410, 101370, 101310, 101310, 101350, 101360, 101410, 101430, 
    101430, 101440, 101400, 101390, 101370, 101320, 101230, 101150, 101010, 
    100870, 100690, 100560, 100410, 100250, 100210, 100050, 99920, 99760, 
    99570, 99470, 99260, 99010, 98790, 98570, 98290, 98070, 97910, 97850, 
    97830, 97840, 97890, 97990, 98120, 98340, 98590, 98810, 98970, 99120, 
    99300, 99420, 99470, 99480, 99580, 99610, 99700, 99690, 99640, 99620, 
    99630, 99630, 99640, 99700, 99800, 99930, 100050, 100190, 100330, 100510, 
    100660, 100820, 100930, 101100, 101300, 101440, 101610, 101750, 101880, 
    102020, 102150, 102260, 102360, 102450, 102510, 102540, 102610, 102700, 
    102720, 102690, 102690, 102760, 102680, 102580, 102500, 102400, 102300, 
    102230, 102120, 101980, 101890, 101760, 101670, 101560, 101470, 101390, 
    101260, 101150, 101040, 100940, 100870, 100800, 100730, 100690, 100640, 
    100620, 100630, 100680, 100730, 100760, 100820, 100890, 100920, 100940, 
    101040, 101080, 101190, 101240, 101250, 101240, 101270, 101320, 101330, 
    101310, 101300, 101300, 101340, 101330, 101320, 101320, 101300, 101270, 
    101260, 101220, 101210, 101210, 101200, 101220, 101210, 101180, 101170, 
    101150, 101120, 101100, 101080, 101050, 101030, 101020, 101000, 101000, 
    101010, 101020, 101010, 101000, 101010, 100990, 100970, 100960, 100950, 
    100950, 100960, 100950, 100960, 100960, 100950, 100900, 100880, 100850, 
    100830, 100820, 100760, 100720, 100730, 100720, 100720, 100690, 100670, 
    100620, 100560, 100530, 100470, 100410, 100370, 100310, 100240, 100190, 
    100130, 100040, 99970, 99900, 99820, 99730, 99580, 99470, 99360, 99220, 
    99090, 99000, 98910, 98760, 98600, 98420, 98280, 98240, 98230, 98270, 
    98270, 98270, 98280, 98270, 98290, 98330, 98330, 98310, 98310, 98290, 
    98320, 98260, 98220, 98210, 98160, 98110, 98040, 97940, 97850, 97850, 
    97830, 97840, 97870, 97900, 97930, 97990, 98000, 97990, 97980, 98000, 
    98020, 98100, 98120, 98190, 98300, 98410, 98520, 98700, 98820, 99000, 
    99170, 99310, 99510, 99550, 99620, 99750, 99830, 99960, 99940, 99980, 
    99990, 100090, 100150, 100140, 100120, 100070, 100080, 100060, 100000, 
    99990, 99960, 99960, 99960, 99950, 99910, 99900, 99960, 99960, 99910, 
    99920, 99940, 99920, 99860, 99880, 99860, 99860, 99850, 99870, 99860, 
    99830, 99850, 99870, 99840, 99860, 99840, 99840, 99830, 99830, 99810, 
    99840, 99800, 99790, 99740, 99720, 99700, 99670, 99630, 99640, 99610, 
    99650, 99690, 99710, 99740, 99790, 99820, 99890, 99920, 99970, 99990, 
    100060, 100050, 100120, 100170, 100250, 100270, 100300, 100320, 100340, 
    100400, 100410, 100450, 100470, 100510, 100520, 100570, 100600, 100630, 
    100670, 100720, 100750, 100760, 100780, 100830, 100860, 100890, 100960, 
    101010, 101070, 101100, 101130, 101170, 101210, 101220, 101270, 101320, 
    101360, 101400, 101430, 101470, 101510, 101560, 101600, 101620, 101650, 
    101650, 101700, 101720, 101760, 101790, 101840, 101890, 101920, 101930, 
    101950, 101970, 102010, 102040, 102060, 102100, 102150, 102200, 102220, 
    102240, 102250, 102250, 102220, 102180, 102190, 102200, 102200, 102170, 
    102130, 102110, 102100, 102070, 101990, 101960, 101920, 101880, 101810, 
    101760, 101720, 101670, 101650, 101600, 101520, 101460, 101400, 101350, 
    101270, 101240, 101200, 101190, 101150, 101100, 101050, 101050, 101050, 
    101040, 101020, 100980, 100960, 100920, 100890, 100910, 100910, 100900, 
    100880, 100860, 100890, 100880, 100890, 100880, 100860, 100840, 100820, 
    100800, 100810, 100840, 100780, 100760, 100750, 100750, 100760, 100770, 
    100780, 100780, 100760, 100740, 100730, 100720, 100730, 100720, 100710, 
    100730, 100740, 100740, 100710, 100710, 100700, 100690, 100700, 100710, 
    100720, 100710, 100730, 100750, 100780, 100810, 100830, 100830, 100880, 
    100930, 100980, 101020, 101060, 101120, 101180, 101220, 101270, 101300, 
    101330, 101380, 101400, 101420, 101450, 101460, 101470, 101500, 101530, 
    101550, 101590, 101620, 101600, 101610, 101630, 101630, 101630, 101630, 
    101620, 101600, 101560, 101530, 101510, 101500, 101440, 101370, 101290, 
    101250, 101220, 101160, 101130, 101070, 101070, 101050, 101020, 101000, 
    100990, 100970, 100940, 100930, 100890, 100880, 100860, 100810, 100780, 
    100750, 100730, 100660, 100620, 100600, 100550, 100540, 100540, 100550, 
    100560, 100570, 100600, 100630, 100700, 100760, 100830, 100890, 100980, 
    101100, 101180, 101260, 101370, 101430, 101470, 101510, 101560, 101600, 
    101630, 101650, 101670, 101630, 101650, 101600, 101530, 101500, 101500, 
    101490, 101470, 101480, 101460, 101430, 101370, 101400, 101350, 101310, 
    101270, 101250, 101250, 101220, 101240, 101260, 101260, 101250, 101240, 
    101240, 101190, 101160, 101130, 101080, 101030, 101000, 100970, 100960, 
    100900, 100860, 100800, 100760, 100740, 100710, 100700, 100710, 100730, 
    100730, 100710, 100700, 100690, 100690, 100680, 100660, 100650, 100640, 
    100660, 100680, 100690, 100760, 100820, 100870, 100930, 100980, 101010, 
    101030, 101060, 101050, 101090, 101110, 101140, 101180, 101190, 101200, 
    101230, 101230, 101210, 101210, 101220, 101230, 101240, 101260, 101270, 
    101270, 101250, 101250, 101240, 101240, 101220, 101190, 101150, 101090, 
    101030, 101000, 100930, 100850, 100770, 100650, 100540, 100360, 100180, 
    99980, 99750, 99690, 99590, 99570, 99540, 99520, 99500, 99490, 99620, 
    99750, 99830, 99920, 99970, 100030, 100110, 100150, 100200, 100220, 
    100290, 100310, 100330, 100350, 100320, 100280, 100230, 100180, 100110, 
    100050, 100010, 99980, 99950, 99930, 99860, 99880, 99840, 99840, 99820, 
    99780, 99800, 99830, 99860, 99910, 99940, 100000, 100050, 100200, 100220, 
    100290, 100410, 100550, 100600, 100680, 100730, 100830, 100900, 100930, 
    100960, 100970, 100970, 101020, 101040, 101040, 101010, 100990, 100940, 
    100890, 100790, 100700, 100600, 100510, 100400, 100270, 100140, 100030, 
    99920, 99850, 99810, 99780, 99750, 99720, 99660, 99610, 99550, 99510, 
    99500, 99470, 99460, 99430, 99410, 99380, 99330, 99270, 99190, 99100, 
    98970, 98840, 98710, 98610, 98510, 98440, 98340, 98230, 98180, 98080, 
    98020, 97930, 97860, 97800, 97710, 97630, 97560, 97510, 97490, 97460, 
    97450, 97470, 97450, 97450, 97480, 97510, 97560, 97600, 97620, 97650, 
    97710, 97810, 97810, 97830, 97870, 97910, 97950, 98000, 98050, 98100, 
    98140, 98170, 98190, 98240, 98280, 98320, 98330, 98360, 98390, 98430, 
    98470, 98480, 98470, 98510, 98520, 98540, 98470, 98520, 98530, 98490, 
    98490, 98480, 98500, 98510, 98450, 98460, 98450, 98470, 98490, 98450, 
    98410, 98380, 98390, 98380, 98350, 98320, 98300, 98300, 98300, 98350, 
    98350, 98380, 98380, 98360, 98390, 98360, 98370, 98370, 98400, 98410, 
    98420, 98410, 98420, 98430, 98430, 98420, 98410, 98420, 98420, 98400, 
    98380, 98390, 98400, 98380, 98370, 98380, 98360, 98350, 98360, 98340, 
    98340, 98340, 98330, 98360, 98360, 98380, 98360, 98370, 98370, 98380, 
    98410, 98420, 98430, 98460, 98500, 98510, 98530, 98540, 98550, 98560, 
    98570, 98580, 98560, 98540, 98530, 98530, 98540, 98530, 98550, 98570, 
    98610, 98630, 98670, 98720, 98750, 98760, 98800, 98850, 98900, 98950, 
    99000, 99050, 99110, 99160, 99230, 99270, 99300, 99360, 99380, 99450, 
    99530, 99560, 99590, 99660, 99700, 99760, 99800, 99850, 99880, 99920, 
    99950, 99960, 99970, 100000, 100010, 100050, 100080, 100100, 100110, 
    100110, 100110, 100110, 100140, 100160, 100150, 100150, 100140, 100140, 
    100140, 100130, 100120, 100120, 100090, 100050, 100010, 100010, 99990, 
    99960, 99920, 99910, 99890, 99880, 99860, 99830, 99790, 99750, 99690, 
    99650, 99590, 99550, 99490, 99470, 99400, 99340, 99320, 99270, 99200, 
    99150, 99130, 99130, 99140, 99130, 99160, 99190, 99220, 99260, 99280, 
    99310, 99320, 99390, 99450, 99530, 99610, 99720, 99750, 99840, 99900, 
    99970, 99970, 100000, 100020, 100030, 99990, 100020, 100010, 100010, 
    100000, 99990, 100010, 100010, 100000, 99990, 99950, 99940, 99940, 99980, 
    100000, 100030, 100040, 100070, 100090, 100140, 100170, 100180, 100190, 
    100160, 100150, 100110, 100070, 100000, 99930, 99940, 99830, 99740, 
    99630, 99550, 99390, 99230, 99080, 98940, 98780, 98650, 98560, 98470, 
    98400, 98340, 98320, 98320, 98350, 98400, 98450, 98500, 98570, 98650, 
    98760, 98900, 99090, 99270, 99360, 99580, 99720, 99820, 99890, 99970, 
    100010, 100090, 100140, 100160, 100230, 100250, 100200, 100230, 100240, 
    100250, 100260, 100240, 100250, 100280, 100320, 100380, 100470, 100470, 
    100560, 100630, 100630, 100730, 100820, 100860, 100870, 100920, 100980, 
    101000, 101050, 101120, 101200, 101170, 101220, 101220, 101290, 101290, 
    101370, 101420, 101420, 101430, 101500, 101500, 101500, 101520, 101510, 
    101500, 101450, 101430, 101490, 101490, 101520, 101550, 101550, 101540, 
    101530, 101500, 101490, 101460, 101440, 101380, 101360, 101320, 101280, 
    101260, 101250, 101230, 101200, 101160, 101120, 101080, 101060, 101040, 
    101050, 101080, 101080, 101080, 101080, 101060, 101060, 101020, 101000, 
    100960, 100950, 100940, 100930, 100950, 100950, 100940, 100940, 100930, 
    100970, 101000, 101020, 101030, 101030, 101020, 101010, 101000, 101000, 
    100960, 100960, 100960, 100960, 100970, 100950, 100930, 100910, 100910, 
    100920, 100920, 100920, 100900, 100920, 100910, 100890, 100880, 100850, 
    100840, 100850, 100840, 100820, 100850, 100840, 100850, 100860, 100860, 
    100870, 100920, 100930, 100950, 100980, 100990, 101020, 101030, 101050, 
    101090, 101120, 101140, 101180, 101170, 101210, 101230, 101260, 101280, 
    101300, 101320, 101330, 101370, 101400, 101440, 101470, 101500, 101530, 
    101540, 101530, 101540, 101540, 101530, 101530, 101510, 101510, 101480, 
    101460, 101450, 101430, 101340, 101240, 101210, 101170, 101130, 101070, 
    100980, 100910, 100860, 100810, 100770, 100700, 100630, 100540, 100460, 
    100410, 100360, 100330, 100300, 100260, 100220, 100210, 100170, 100130, 
    100180, 100160, 100150, 100150, 100220, 100250, 100340, 100430, 100470, 
    100530, 100560, 100600, 100640, 100660, 100660, 100680, 100710, 100710, 
    100700, 100730, 100750, 100730, 100720, 100730, 100720, 100730, 100740, 
    100770, 100790, 100790, 100810, 100830, 100810, 100800, 100790, 100790, 
    100770, 100800, 100800, 100790, 100780, 100790, 100810, 100880, 100930, 
    100950, 100970, 101020, 101040, 101060, 101040, 101030, 101010, 101020, 
    101030, 101030, 101030, 101030, 101020, 101020, 101020, 101010, 101020, 
    101030, 101060, 101060, 101120, 101130, 101140, 101150, 101180, 101200, 
    101220, 101260, 101280, 101310, 101360, 101330, 101340, 101350, 101350, 
    101380, 101400, 101410, 101430, 101450, 101480, 101510, 101530, 101550, 
    101560, 101580, 101570, 101580, 101590, 101580, 101600, 101620, 101630, 
    101640, 101640, 101660, 101670, 101660, 101650, 101650, 101610, 101580, 
    101570, 101550, 101530, 101520, 101520, 101520, 101510, 101520, 101520, 
    101500, 101480, 101440, 101410, 101390, 101340, 101340, 101300, 101280, 
    101290, 101270, 101240, 101180, 101140, 101110, 101100, 101100, 101110, 
    101100, 101110, 101130, 101120, 101100, 101090, 101060, 101040, 101020, 
    100980, 100950, 100940, 100900, 100880, 100880, 100840, 100830, 100810, 
    100790, 100810, 100790, 100810, 100830, 100860, 100900, 100910, 100940, 
    100930, 100940, 101000, 101010, 101040, 101060, 101090, 101110, 101150, 
    101170, 101190, 101220, 101270, 101300, 101320, 101340, 101390, 101420, 
    101450, 101460, 101510, 101540, 101580, 101610, 101650, 101680, 101720, 
    101740, 101770, 101800, 101820, 101820, 101840, 101870, 101900, 101950, 
    101980, 101980, 102000, 102030, 102050, 102080, 102080, 102090, 102110, 
    102150, 102200, 102220, 102240, 102260, 102280, 102290, 102290, 102310, 
    102310, 102310, 102320, 102310, 102320, 102350, 102360, 102360, 102360, 
    102360, 102370, 102350, 102330, 102310, 102300, 102310, 102300, 102300, 
    102300, 102300, 102290, 102270, 102250, 102250, 102210, 102190, 102160, 
    102130, 102130, 102110, 102070, 102030, 101980, 101940, 101880, 101850, 
    101820, 101830, 101890, 101970, 102050, 102090, 102140, 102170, 102200, 
    102240, 102320, 102330, 102370, 102370, 102380, 102390, 102400, 102420, 
    102420, 102440, 102450, 102450, 102460, 102480, 102500, 102520, 102510, 
    102500, 102480, 102490, 102480, 102490, 102510, 102480, 102450, 102460, 
    102430, 102420, 102400, 102420, 102430, 102430, 102440, 102460, 102440, 
    102410, 102420, 102410, 102390, 102400, 102380, 102360, 102360, 102350, 
    102320, 102310, 102290, 102300, 102300, 102280, 102290, 102270, 102280, 
    102270, 102260, 102260, 102260, 102260, 102230, 102220, 102220, 102210, 
    102200, 102190, 102160, 102130, 102120, 102100, 102090, 102070, 102030, 
    102020, 102000, 101970, 101970, 101950, 101920, 101920, 101910, 101920, 
    101920, 101910, 101890, 101890, 101900, 101930, 101930, 101900, 101900, 
    101920, 101930, 101930, 101940, 101950, 101980, 101970, 101950, 101950, 
    101950, 101930, 101930, 101920, 101930, 101920, 101900, 101920, 101910, 
    101910, 101900, 101880, 101850, 101810, 101780, 101770, 101760, 101760, 
    101750, 101730, 101720, 101720, 101690, 101680, 101650, 101620, 101600, 
    101580, 101570, 101550, 101530, 101510, 101510, 101490, 101450, 101420, 
    101400, 101360, 101350, 101340, 101330, 101350, 101360, 101370, 101360, 
    101320, 101320, 101290, 101250, 101240, 101250, 101260, 101300, 101340, 
    101380, 101370, 101370, 101370, 101340, 101340, 101320, 101270, 101260, 
    101260, 101220, 101270, 101260, 101250, 101240, 101230, 101240, 101250, 
    101240, 101280, 101350, 101400, 101450, 101420, 101510, 101540, 101550, 
    101590, 101600, 101600, 101650, 101670, 101690, 101690, 101720, 101750, 
    101790, 101790, 101780, 101800, 101810, 101800, 101780, 101780, 101790, 
    101800, 101810, 101830, 101840, 101840, 101830, 101820, 101800, 101810, 
    101780, 101770, 101730, 101740, 101770, 101790, 101810, 101790, 101790, 
    101780, 101760, 101740, 101740, 101780, 101780, 101800, 101810, 101840, 
    101860, 101860, 101870, 101840, 101850, 101830, 101810, 101800, 101810, 
    101800, 101800, 101800, 101800, 101820, 101790, 101780, 101770, 101750, 
    101740, 101740, 101730, 101730, 101740, 101750, 101730, 101720, 101700, 
    101670, 101640, 101630, 101610, 101580, 101570, 101560, 101540, 101540, 
    101530, 101520, 101520, 101500, 101500, 101510, 101500, 101490, 101470, 
    101480, 101500, 101510, 101520, 101520, 101540, 101550, 101570, 101570, 
    101590, 101580, 101580, 101600, 101610, 101630, 101630, 101650, 101650, 
    101640, 101630, 101610, 101600, 101580, 101560, 101530, 101510, 101450, 
    101380, 101300, 101240, 101180, 101140, 101110, 101050, 101030, 101010, 
    100980, 100990, 101010, 101020, 101010, 101020, 101040, 101040, 101040, 
    101040, 101020, 101000, 100980, 100980, 100960, 100940, 100910, 100860, 
    100820, 100770, 100700, 100660, 100590, 100550, 100520, 100500, 100480, 
    100520, 100580, 100680, 100770, 100870, 100920, 100990, 100990, 101030, 
    101050, 101060, 101080, 101080, 101070, 101070, 101100, 101100, 101200, 
    101210, 101250, 101300, 101340, 101370, 101410, 101460, 101490, 101580, 
    101640, 101720, 101820, 101930, 102060, 102180, 102290, 102380, 102500, 
    102600, 102670, 102710, 102770, 102840, 102850, 102870, 102880, 102890, 
    102910, 102930, 102960, 103000, 103010, 103030, 103040, 103030, 103000, 
    102960, 102920, 102900, 102900, 102880, 102840, 102820, 102810, 102760, 
    102700, 102670, 102640, 102620, 102540, 102470, 102410, 102370, 102320, 
    102320, 102260, 102230, 102190, 102170, 102130, 102090, 102070, 102040, 
    102020, 102010, 102000, 102020, 102030, 102030, 102020, 102030, 102020, 
    102050, 102070, 102110, 102160, 102220, 102250, 102310, 102360, 102420, 
    102470, 102530, 102580, 102590, 102610, 102650, 102670, 102690, 102700, 
    102710, 102710, 102690, 102710, 102720, 102720, 102690, 102650, 102610, 
    102550, 102530, 102440, 102380, 102280, 102170, 102030, 101910, 101790, 
    101700, 101590, 101520, 101460, 101370, 101330, 101250, 101230, 101170, 
    101130, 101120, 101090, 101060, 101000, 101030, 101010, 101020, 100990, 
    101000, 101010, 100950, 100990, 101050, 101100, 101130, 101170, 101240, 
    101330, 101350, 101450, 101560, 101610, 101680, 101770, 101820, 101900, 
    101990, 102050, 102110, 102160, 102260, 102340, 102440, 102510, 102560, 
    102620, 102690, 102730, 102770, 102770, 102800, 102800, 102820, 102850, 
    102850, 102870, 102880, 102880, 102870, 102860, 102840, 102800, 102780, 
    102770, 102760, 102760, 102770, 102820, 102770, 102860, 102890, 102920, 
    102910, 102920, 102970, 102970, 102970, 102990, 103030, 103020, 103000, 
    103040, 103020, 103020, 103040, 103050, 103060, 103040, 103050, 103070, 
    103090, 103110, 103120, 103110, 103110, 103120, 103100, 103100, 103130, 
    103140, 103190, 103180, 103200, 103200, 103220, 103230, 103210, 103220, 
    103230, 103240, 103250, 103250, 103230, 103270, 103270, 103280, 103280, 
    103310, 103290, 103270, 103270, 103250, 103220, 103210, 103200, 103200, 
    103190, 103160, 103160, 103130, 103110, 103090, 103080, 103060, 103030, 
    103040, 103060, 103070, 103080, 103100, 103120, 103160, 103180, 103210, 
    103230, 103260, 103300, 103330, 103380, 103400, 103430, 103440, 103460, 
    103460, 103450, 103440, 103420, 103390, 103460, 103340, 103330, 103310, 
    103310, 103290, 103260, 103230, 103210, 103190, 103160, 103130, 103100, 
    103070, 103060, 103070, 103060, 103030, 103000, 102990, 102960, 102940, 
    102920, 102890, 102850, 102850, 102850, 102860, 102870, 102860, 102850, 
    102840, 102840, 102840, 102830, 102820, 102840, 102840, 102850, 102860, 
    102860, 102880, 102890, 102890, 102890, 102910, 102900, 102890, 102880, 
    102900, 102890, 102900, 102920, 102930, 102940, 102930, 102930, 102930, 
    102920, 102900, 102900, 102900, 102910, 102920, 102940, 102940, 102940, 
    102940, 102940, 102960, 102940, 102930, 102930, 102940, 102960, 102980, 
    102980, 102990, 103010, 103030, 103040, 103030, 103050, 103060, 103050, 
    103060, 103060, 103070, 103090, 103100, 103080, 103060, 103070, 103070, 
    103070, 103080, 103070, 103060, 103040, 103030, 103010, 102980, 102960, 
    102910, 102860, 102810, 102740, 102670, 102570, 102440, 102360, 102270, 
    102190, 102120, 102050, 101920, 101810, 101690, 101670, 101650, 101640, 
    101610, 101590, 101590, 101580, 101620, 101620, 101660, 101670, 101700, 
    101740, 101770, 101790, 101830, 101850, 101880, 101890, 101920, 101940, 
    101950, 101960, 101980, 101980, 101960, 101940, 101960, 101970, 101980, 
    102020, 102020, 102020, 102020, 102020, 102010, 102020, 102030, 102020, 
    102030, 102030, 102050, 102080, 102080, 102100, 102110, 102120, 102100, 
    102120, 102110, 102120, 102120, 102130, 102120, 102150, 102160, 102170, 
    102180, 102180, 102170, 102150, 102140, 102140, 102140, 102110, 102110, 
    102110, 102100, 102090, 102070, 102060, 102040, 102020, 102000, 101990, 
    101980, 101980, 101980, 101980, 101990, 102000, 102000, 102000, 102000, 
    101990, 101970, 101960, 101940, 101940, 101950, 101950, 101960, 101940, 
    101930, 101930, 101930, 101940, 101930, 101920, 101930, 101950, 101960, 
    101990, 101990, 101990, 101980, 101990, 102000, 101980, 101960, 101950, 
    101950, 101940, 101950, 101950, 101950, 101930, 101910, 101900, 101860, 
    101850, 101810, 101780, 101760, 101760, 101750, 101770, 101770, 101760, 
    101730, 101710, 101670, 101630, 101620, 101610, 101570, 101550, 101530, 
    101510, 101510, 101490, 101480, 101450, 101440, 101400, 101370, 101330, 
    101290, 101280, 101240, 101210, 101180, 101150, 101090, 101050, 100980, 
    100930, 100890, 100840, 100790, 100770, 100770, 100770, 100790, 100810, 
    100790, 100770, 100790, 100790, 100800, 100830, 100820, 100820, 100840, 
    100880, 100880, 100880, 100900, 100910, 100920, 100930, 100930, 100950, 
    100960, 101010, 101010, 101030, 101040, 101050, 101060, 101070, 101070, 
    101060, 101060, 101060, 101040, 101050, 101090, 101100, 101090, 101110, 
    101100, 101090, 101090, 101090, 101090, 101120, 101110, 101110, 101100, 
    101100, 101130, 101130, 101150, 101150, 101150, 101150, 101170, 101170, 
    101160, 101190, 101200, 101210, 101220, 101230, 101250, 101260, 101280, 
    101300, 101320, 101330, 101350, 101350, 101350, 101370, 101380, 101380, 
    101390, 101410, 101430, 101440, 101440, 101460, 101480, 101520, 101540, 
    101570, 101590, 101610, 101630, 101650, 101660, 101660, 101680, 101670, 
    101690, 101690, 101700, 101710, 101720, 101730, 101730, 101740, 101720, 
    101720, 101710, 101710, 101690, 101680, 101670, 101680, 101680, 101660, 
    101640, 101640, 101660, 101660, 101650, 101640, 101640, 101660, 101700, 
    101710, 101750, 101790, 101820, 101850, 101890, 101910, 101920, 101940, 
    101960, 102010, 102030, 102060, 102070, 102110, 102130, 102140, 102150, 
    102160, 102150, 102140, 102150, 102140, 102150, 102150, 102160, 102160, 
    102160, 102150, 102150, 102140, 102110, 102090, 102080, 102080, 102090, 
    102110, 102110, 102130, 102140, 102140, 102130, 102130, 102130, 102120, 
    102110, 102130, 102150, 102140, 102110, 102080, 102020, 101960, 101920, 
    101900, 101830, 101780, 101730, 101650, 101620, 101570, 101500, 101460, 
    101410, 101320, 101220, 101260, 101180, 101130, 101080, 101110, 101110, 
    101110, 101110, 101120, 101140, 101150, 101220, 101230, 101260, 101290, 
    101340, 101370, 101400, 101430, 101390, 101370, 101390, 101380, 101380, 
    101490, 101510, 101520, 101490, 101600, 101660, 101680, 101750, 101760, 
    101790, 101820, 101880, 101900, 101890, 101910, 101940, 101920, 101930, 
    101920, 101920, 101920, 101910, 101910, 101920, 101940, 101950, 102010, 
    102040, 102040, 102090, 102120, 102150, 102250, 102320, 102370, 102390, 
    102430, 102470, 102500, 102570, 102610, 102640, 102680, 102720, 102750, 
    102780, 102820, 102820, 102870, 102900, 102930, 102960, 102990, 103010, 
    103020, 103030, 103020, 103010, 103020, 103030, 103030, 103020, 103020, 
    103000, 103010, 103010, 102990, 102970, 102970, 102960, 102940, 102940, 
    102910, 102880, 102840, 102800, 102770, 102740, 102710, 102690, 102660, 
    102610, 102580, 102550, 102510, 102480, 102440, 102420, 102420, 102410, 
    102390, 102360, 102350, 102340, 102350, 102340, 102340, 102340, 102330, 
    102320, 102310, 102310, 102320, 102330, 102320, 102340, 102350, 102360, 
    102390, 102380, 102380, 102400, 102390, 102400, 102430, 102460, 102450, 
    102420, 102420, 102440, 102440, 102450, 102440, 102410, 102410, 102380, 
    102390, 102360, 102330, 102320, 102310, 102290, 102270, 102260, 102220, 
    102190, 102160, 102160, 102140, 102100, 102050, 102030, 102000, 101980, 
    101960, 101930, 101910, 101900, 101890, 101820, 101810, 101780, 101760, 
    101750, 101720, 101680, 101680, 101660, 101640, 101660, 101630, 101650, 
    101650, 101630, 101680, 101710, 101710, 101730, 101760, 101790, 101800, 
    101820, 101850, 101890, 101930, 101940, 101980, 102010, 102030, 102050, 
    102070, 102070, 102060, 102060, 102070, 102080, 102080, 102050, 102040, 
    102060, 102090, 102100, 102110, 102120, 102170, 102180, 102210, 102240, 
    102270, 102280, 102310, 102330, 102380, 102420, 102430, 102430, 102460, 
    102500, 102520, 102560, 102590, 102620, 102630, 102650, 102690, 102710, 
    102730, 102740, 102740, 102740, 102740, 102770, 102800, 102820, 102840, 
    102860, 102870, 102880, 102900, 102910, 102900, 102920, 102920, 102930, 
    102950, 102920, 102910, 102920, 102910, 102910, 102910, 102890, 102870, 
    102830, 102820, 102820, 102790, 102770, 102730, 102730, 102730, 102720, 
    102700, 102700, 102680, 102690, 102680, 102680, 102680, 102660, 102650, 
    102660, 102650, 102640, 102630, 102600, 102550, 102500, 102470, 102450, 
    102410, 102380, 102340, 102290, 102240, 102220, 102180, 102130, 102080, 
    102020, 101980, 101940, 101910, 101890, 101870, 101830, 101800, 101760, 
    101730, 101690, 101650, 101620, 101580, 101550, 101520, 101500, 101470, 
    101450, 101430, 101400, 101340, 101300, 101260, 101220, 101190, 101170, 
    101150, 101140, 101120, 101100, 101100, 101080, 101060, 101050, 101020, 
    101000, 100990, 100970, 100950, 100940, 100930, 100920, 100880, 100870, 
    100860, 100860, 100830, 100800, 100780, 100790, 100790, 100780, 100750, 
    100740, 100740, 100720, 100700, 100670, 100620, 100600, 100570, 100550, 
    100530, 100500, 100450, 100430, 100400, 100380, 100350, 100310, 100270, 
    100240, 100220, 100220, 100190, 100180, 100190, 100180, 100150, 100150, 
    100150, 100160, 100160, 100170, 100180, 100170, 100180, 100170, 100190, 
    100180, 100180, 100180, 100180, 100160, 100140, 100130, 100130, 100120, 
    100140, 100150, 100160, 100160, 100140, 100130, 100130, 100110, 100100, 
    100080, 100090, 100090, 100090, 100100, 100110, 100130, 100150, 100180, 
    100210, 100220, 100250, 100270, 100320, 100370, 100400, 100440, 100480, 
    100530, 100560, 100570, 100600, 100630, 100660, 100690, 100720, 100750, 
    100790, 100810, 100830, 100860, 100870, 100890, 100900, 100890, 100900, 
    100910, 100910, 100900, 100900, 100920, 100920, 100920, 100920, 100910, 
    100880, 100860, 100840, 100830, 100810, 100790, 100800, 100780, 100790, 
    100790, 100790, 100760, 100730, 100710, 100690, 100690, 100710, 100720, 
    100730, 100730, 100750, 100740, 100750, 100750, 100760, 100740, 100730, 
    100730, 100730, 100740, 100740, 100750, 100750, 100760, 100750, 100740, 
    100720, 100710, 100690, 100680, 100700, 100690, 100690, 100720, 100710, 
    100700, 100690, 100690, 100670, 100670, 100670, 100660, 100650, 100630, 
    100640, 100630, 100630, 100620, 100650, 100660, 100670, 100680, 100680, 
    100700, 100730, 100790, 100820, 100840, 100840, 100860, 100860, 100880, 
    100900, 100940, 100940, 100960, 100980, 100990, 101000, 101020, 101040, 
    101030, 101050, 101050, 101070, 101070, 101080, 101100, 101110, 101130, 
    101150, 101130, 101130, 101160, 101180, 101160, 101170, 101160, 101170, 
    101180, 101180, 101180, 101180, 101170, 101200, 101200, 101200, 101200, 
    101190, 101190, 101200, 101210, 101220, 101200, 101190, 101180, 101180, 
    101190, 101180, 101160, 101150, 101140, 101120, 101110, 101110, 101110, 
    101110, 101110, 101100, 101110, 101130, 101130, 101130, 101120, 101130, 
    101130, 101120, 101140, 101150, 101160, 101150, 101150, 101130, 101140, 
    101140, 101110, 101100, 101090, 101060, 101030, 101020, 101030, 101040, 
    101030, 101030, 101030, 101000, 100990, 100980, 100990, 100990, 100980, 
    101000, 101000, 100990, 100990, 100990, 100990, 100980, 100990, 100970, 
    100950, 100960, 100970, 100980, 100970, 100990, 100990, 100990, 100990, 
    100950, 100950, 100940, 100940, 100930, 100910, 100930, 100930, 100930, 
    100910, 100900, 100860, 100860, 100860, 100850, 100830, 100810, 100810, 
    100780, 100760, 100750, 100720, 100700, 100670, 100640, 100610, 100570, 
    100540, 100520, 100500, 100490, 100470, 100450, 100430, 100390, 100360, 
    100360, 100330, 100320, 100300, 100300, 100300, 100280, 100270, 100270, 
    100260, 100240, 100240, 100240, 100230, 100230, 100230, 100230, 100230, 
    100240, 100250, 100240, 100250, 100250, 100240, 100240, 100260, 100260, 
    100230, 100220, 100210, 100220, 100200, 100180, 100170, 100140, 100110, 
    100070, 100050, 100030, 99990, 99990, 99990, 99970, 99940, 99910, 99900, 
    99890, 99860, 99830, 99840, 99830, 99850, 99860, 99880, 99890, 99950, 
    99960, 99980, 100020, 100050, 100090, 100120, 100160, 100210, 100260, 
    100290, 100350, 100390, 100420, 100480, 100530, 100600, 100660, 100720, 
    100780, 100850, 100900, 100990, 101060, 101120, 101190, 101240, 101300, 
    101340, 101370, 101390, 101430, 101470, 101480, 101530, 101560, 101590, 
    101610, 101630, 101640, 101660, 101690, 101710, 101700, 101720, 101750, 
    101780, 101810, 101820, 101820, 101840, 101820, 101810, 101800, 101770, 
    101760, 101750, 101720, 101710, 101720, 101690, 101680, 101660, 101630, 
    101610, 101580, 101540, 101510, 101490, 101490, 101470, 101480, 101490, 
    101470, 101460, 101430, 101420, 101400, 101390, 101370, 101360, 101370, 
    101370, 101380, 101350, 101350, 101350, 101350, 101350, 101340, 101340, 
    101320, 101320, 101330, 101310, 101330, 101340, 101340, 101340, 101340, 
    101330, 101300, 101270, 101230, 101200, 101190, 101170, 101160, 101180, 
    101170, 101170, 101120, 101070, 101050, 100980, 100970, 100930, 100880, 
    100850, 100830, 100760, 100700, 100680, 100640, 100610, 100580, 100540, 
    100500, 100460, 100450, 100420, 100390, 100380, 100340, 100320, 100290, 
    100270, 100230, 100190, 100170, 100150, 100140, 100150, 100150, 100140, 
    100150, 100140, 100140, 100120, 100140, 100150, 100150, 100160, 100170, 
    100200, 100240, 100270, 100300, 100320, 100350, 100380, 100420, 100430, 
    100450, 100480, 100500, 100540, 100570, 100630, 100700, 100720, 100730, 
    100760, 100780, 100790, 100780, 100810, 100820, 100860, 100900, 100940, 
    100970, 100980, 100980, 100990, 100990, 100980, 100990, 100980, 100970, 
    100980, 101000, 101010, 101010, 101010, 100990, 100960, 100940, 100930, 
    100910, 100900, 100890, 100860, 100840, 100820, 100800, 100760, 100710, 
    100690, 100660, 100610, 100570, 100540, 100500, 100460, 100420, 100410, 
    100380, 100340, 100300, 100260, 100240, 100210, 100180, 100160, 100130, 
    100110, 100130, 100130, 100150, 100160, 100130, 100130, 100120, 100130, 
    100140, 100150, 100170, 100190, 100220, 100260, 100290, 100340, 100360, 
    100390, 100410, 100430, 100450, 100470, 100480, 100510, 100520, 100530, 
    100540, 100550, 100540, 100540, 100540, 100540, 100570, 100580, 100620, 
    100650, 100670, 100710, 100760, 100760, 100780, 100790, 100790, 100810, 
    100840, 100860, 100880, 100910, 100920, 100920, 100930, 100930, 100930, 
    100940, 100940, 100950, 100940, 100940, 100940, 100930, 100940, 100950, 
    100950, 100940, 100930, 100910, 100890, 100900, 100880, 100860, 100850, 
    100830, 100810, 100800, 100800, 100810, 100800, 100770, 100760, 100750, 
    100740, 100740, 100730, 100740, 100740, 100750, 100740, 100730, 100720, 
    100720, 100700, 100700, 100680, 100690, 100690, 100700, 100700, 100700, 
    100690, 100680, 100700, 100700, 100700, 100710, 100730, 100740, 100740, 
    100760, 100740, 100750, 100720, 100720, 100720, 100690, 100660, 100640, 
    100610, 100600, 100570, 100520, 100510, 100450, 100410, 100390, 100360, 
    100310, 100270, 100250, 100210, 100170, 100160, 100130, 100100, 100090, 
    100090, 100090, 100100, 100090, 100090, 100070, 100040, 100030, 100110, 
    100170, 100250, 100320, 100380, 100410, 100500, 100570, 100620, 100720, 
    100790, 100890, 100990, 101050, 101130, 101190, 101200, 101210, 101260, 
    101270, 101310, 101340, 101370, 101390, 101400, 101410, 101440, 101450, 
    101450, 101430, 101410, 101380, 101390, 101380, 101340, 101300, 101270, 
    101230, 101250, 101190, 101160, 101070, 101010, 100950, 100870, 100810, 
    100750, 100620, 100520, 100450, 100390, 100330, 100280, 100220, 100130, 
    100060, 100040, 100010, 100010, 100030, 100030, 100020, 100060, 100090, 
    100110, 100110, 100120, 100110, 100090, 100050, 100020, 100050, 100030, 
    100070, 100090, 100140, 100160, 100200, 100280, 100290, 100310, 100360, 
    100440, 100510, 100570, 100590, 100640, 100720, 100780, 100810, 100840, 
    100880, 100880, 100930, 100990, 100980, 101010, 101040, 101060, 101080, 
    101090, 101090, 101070, 101090, 101060, 101010, 100990, 100970, 100950, 
    100940, 100940, 100930, 100900, 100850, 100850, 100820, 100790, 100800, 
    100780, 100790, 100780, 100780, 100770, 100780, 100800, 100820, 100840, 
    100850, 100870, 100890, 100930, 100970, 101000, 101040, 101060, 101100, 
    101120, 101130, 101120, 101140, 101160, 101130, 101120, 101080, 101040, 
    100980, 100920, 100860, 100790, 100730, 100680, 100620, 100610, 100630, 
    100650, 100660, 100670, 100680, 100710, 100750, 100770, 100820, 100860, 
    100910, 100920, 100940, 100970, 101010, 101060, 101130, 101180, 101240, 
    101300, 101380, 101450, 101490, 101530, 101550, 101580, 101620, 101670, 
    101720, 101780, 101830, 101850, 101880, 101910, 101930, 101950, 101980, 
    101990, 101990, 101970, 101960, 101980, 101980, 101990, 102010, 101980, 
    101940, 101880, 101830, 101790, 101740, 101700, 101670, 101590, 101570, 
    101540, 101520, 101540, 101590, 101630, 101660, 101690, 101750, 101790, 
    101810, 101840, 101850, 101910, 101980, 101990, 101980, 101950, 101960, 
    101970, 101980, 101980, 101970, 101970, 101960, 101960, 101960, 101960, 
    101930, 101930, 101920, 101890, 101880, 101870, 101850, 101840, 101810, 
    101780, 101760, 101720, 101670, 101600, 101570, 101550, 101490, 101470, 
    101470, 101450, 101420, 101370, 101350, 101340, 101340, 101330, 101310, 
    101300, 101290, 101300, 101330, 101350, 101370, 101390, 101410, 101400, 
    101400, 101400, 101410, 101430, 101440, 101460, 101480, 101490, 101510, 
    101540, 101550, 101550, 101550, 101540, 101530, 101520, 101510, 101490, 
    101460, 101430, 101410, 101410, 101370, 101330, 101310, 101270, 101240, 
    101190, 101160, 101140, 101110, 101100, 101060, 101020, 100990, 100970, 
    100920, 100880, 100870, 100850, 100840, 100800, 100770, 100740, 100720, 
    100710, 100690, 100680, 100680, 100650, 100620, 100610, 100610, 100580, 
    100580, 100570, 100570, 100550, 100540, 100530, 100520, 100500, 100500, 
    100530, 100550, 100570, 100610, 100640, 100680, 100720, 100760, 100810, 
    100840, 100880, 100910, 100930, 101020, 101040, 101060, 101090, 101150, 
    101180, 101190, 101210, 101220, 101250, 101250, 101270, 101290, 101290, 
    101310, 101340, 101350, 101370, 101370, 101390, 101400, 101380, 101400, 
    101410, 101400, 101420, 101440, 101460, 101480, 101480, 101500, 101480, 
    101460, 101440, 101450, 101430, 101430, 101430, 101430, 101470, 101470, 
    101460, 101460, 101440, 101450, 101440, 101420, 101420, 101440, 101450, 
    101440, 101450, 101460, 101430, 101420, 101390, 101350, 101330, 101310, 
    101280, 101260, 101270, 101240, 101230, 101190, 101180, 101160, 101130, 
    101110, 101080, 101060, 101070, 101060, 101080, 101090, 101100, 101100, 
    101090, 101060, 101030, 101010, 101010, 100990, 100960, 100930, 100970, 
    100970, 100940, 100920, 100910, 100910, 100910, 100880, 100850, 100840, 
    100830, 100840, 100830, 100860, 100860, 100880, 100890, 100890, 100900, 
    100900, 100910, 100920, 100920, 100930, 100940, 100970, 100980, 101010, 
    101010, 101000, 101000, 100990, 100990, 100990, 101010, 101020, 101040, 
    101040, 101040, 101080, 101130, 101110, 101090, 101090, 101100, 101100, 
    101080, 101080, 101090, 101090, 101090, 101090, 101110, 101100, 101090, 
    101070, 101050, 101020, 101020, 101030, 101030, 101050, 101060, 101070, 
    101070, 101080, 101090, 101090, 101090, 101100, 101100, 101110, 101110, 
    101100, 101110, 101130, 101140, 101140, 101140, 101130, 101130, 101110, 
    101110, 101110, 101130, 101150, 101150, 101180, 101190, 101190, 101200, 
    101220, 101220, 101220, 101230, 101240, 101250, 101270, 101280, 101320, 
    101350, 101370, 101390, 101410, 101420, 101410, 101400, 101410, 101440, 
    101440, 101450, 101460, 101470, 101480, 101490, 101470, 101480, 101470, 
    101470, 101480, 101510, 101530, 101540, 101560, 101570, 101580, 101590, 
    101580, 101560, 101570, 101560, 101550, 101550, 101560, 101570, 101580, 
    101580, 101580, 101580, 101580, 101580, 101560, 101550, 101550, 101540, 
    101550, 101550, 101560, 101560, 101560, 101560, 101550, 101550, 101540, 
    101540, 101530, 101560, 101560, 101580, 101590, 101610, 101640, 101650, 
    101660, 101660, 101660, 101660, 101680, 101700, 101720, 101730, 101770, 
    101800, 101820, 101840, 101870, 101880, 101890, 101890, 101890, 101910, 
    101940, 101980, 102000, 102030, 102050, 102070, 102070, 102080, 102080, 
    102070, 102080, 102100, 102100, 102100, 102110, 102110, 102110, 102100, 
    102080, 102050, 102030, 101990, 101970, 101950, 101960, 101930, 101910, 
    101880, 101830, 101810, 101780, 101730, 101700, 101670, 101660, 101660, 
    101650, 101650, 101650, 101630, 101640, 101630, 101610, 101600, 101580, 
    101570, 101560, 101530, 101530, 101510, 101500, 101500, 101480, 101470, 
    101440, 101420, 101400, 101370, 101350, 101330, 101330, 101330, 101310, 
    101300, 101270, 101220, 101190, 101170, 101140, 101130, 101130, 101130, 
    101100, 101090, 101060, 101030, 100990, 100930, 100890, 100840, 100780, 
    100750, 100690, 100660, 100620, 100620, 100580, 100560, 100520, 100480, 
    100490, 100490, 100450, 100420, 100390, 100360, 100310, 100310, 100290, 
    100270, 100250, 100230, 100210, 100200, 100190, 100180, 100160, 100160, 
    100140, 100100, 100090, 100070, 100040, 100000, 99970, 99940, 99940, 
    99910, 99900, 99870, 99850, 99830, 99810, 99780, 99760, 99740, 99690, 
    99650, 99620, 99550, 99530, 99500, 99490, 99460, 99440, 99420, 99390, 
    99380, 99370, 99350, 99350, 99330, 99310, 99310, 99310, 99300, 99330, 
    99330, 99340, 99360, 99360, 99370, 99400, 99430, 99450, 99470, 99490, 
    99510, 99540, 99580, 99610, 99620, 99620, 99590, 99590, 99610, 99600, 
    99600, 99590, 99580, 99580, 99570, 99550, 99520, 99510, 99510, 99490, 
    99470, 99480, 99510, 99500, 99510, 99510, 99550, 99620, 99730, 99860, 
    99970, 100140, 100260, 100350, 100470, 100570, 100670, 100780, 100870, 
    100910, 100950, 100950, 100990, 101000, 101010, 101020, 101030, 101030, 
    101060, 101070, 101090, 101100, 101140, 101170, 101190, 101220, 101240, 
    101260, 101290, 101300, 101340, 101360, 101360, 101380, 101400, 101410, 
    101430, 101430, 101420, 101450, 101480, 101490, 101520, 101540, 101540, 
    101540, 101510, 101500, 101500, 101500, 101490, 101500, 101500, 101510, 
    101520, 101510, 101500, 101520, 101500, 101500, 101490, 101480, 101460, 
    101460, 101460, 101460, 101440, 101430, 101410, 101390, 101350, 101330, 
    101280, 101260, 101230, 101230, 101230, 101210, 101210, 101190, 101190, 
    101180, 101170, 101130, 101090, 101060, 101050, 101030, 101030, 101030, 
    101030, 101000, 101000, 100980, 100980, 100940, 100920, 100920, 100890, 
    100880, 100860, 100880, 100880, 100870, 100870, 100870, 100870, 100860, 
    100840, 100830, 100830, 100830, 100830, 100840, 100850, 100870, 100870, 
    100870, 100880, 100860, 100840, 100820, 100810, 100800, 100830, 100850, 
    100880, 100900, 100920, 100950, 100980, 101000, 101040, 101040, 101080, 
    101110, 101130, 101180, 101220, 101270, 101320, 101350, 101370, 101390, 
    101400, 101420, 101440, 101460, 101490, 101520, 101560, 101600, 101610, 
    101650, 101680, 101670, 101660, 101680, 101710, 101720, 101720, 101720, 
    101750, 101770, 101780, 101800, 101810, 101800, 101810, 101810, 101800, 
    101810, 101800, 101820, 101840, 101830, 101840, 101860, 101860, 101850, 
    101840, 101840, 101850, 101850, 101840, 101840, 101830, 101810, 101760, 
    101740, 101690, 101650, 101600, 101580, 101560, 101550, 101500, 101460, 
    101410, 101380, 101350, 101340, 101310, 101270, 101250, 101170, 101140, 
    101100, 101080, 101070, 101070, 101030, 100960, 100970, 100950, 100940, 
    100890, 100870, 100830, 100820, 100820, 100800, 100780, 100760, 100740, 
    100720, 100660, 100620, 100600, 100570, 100550, 100530, 100520, 100510, 
    100470, 100460, 100450, 100460, 100480, 100470, 100490, 100510, 100540, 
    100580, 100610, 100640, 100660, 100700, 100700, 100700, 100680, 100690, 
    100690, 100680, 100650, 100630, 100640, 100650, 100670, 100660, 100640, 
    100630, 100610, 100600, 100560, 100520, 100480, 100450, 100410, 100350, 
    100290, 100250, 100190, 100130, 100080, 100020, 99990, 99940, 99920, 
    99910, 99870, 99870, 99860, 99840, 99810, 99780, 99750, 99750, 99720, 
    99710, 99680, 99640, 99620, 99590, 99580, 99550, 99540, 99530, 99520, 
    99500, 99480, 99460, 99450, 99450, 99440, 99440, 99430, 99410, 99420, 
    99390, 99350, 99310, 99250, 99220, 99190, 99140, 99130, 99100, 99050, 
    99010, 98960, 98930, 98900, 98870, 98850, 98840, 98830, 98850, 98850, 
    98900, 98930, 98980, 99010, 99050, 99090, 99130, 99170, 99150, 99210, 
    99240, 99270, 99300, 99330, 99360, 99410, 99460, 99500, 99520, 99570, 
    99620, 99680, 99730, 99790, 99860, 99930, 99980, 100060, 100140, 100190, 
    100240, 100290, 100340, 100390, 100410, 100460, 100500, 100560, 100590, 
    100600, 100630, 100680, 100690, 100710, 100720, 100720, 100730, 100750, 
    100780, 100770, 100770, 100770, 100750, 100760, 100760, 100750, 100750, 
    100740, 100750, 100750, 100770, 100780, 100780, 100770, 100790, 100780, 
    100780, 100780, 100780, 100790, 100780, 100780, 100770, 100780, 100780, 
    100780, 100790, 100790, 100760, 100730, 100720, 100700, 100680, 100650, 
    100610, 100560, 100540, 100530, 100480, 100390, 100290, 100190, 100120, 
    100060, 100020, 99970, 99940, 99940, 99900, 99840, 99800, 99750, 99710, 
    99660, 99670, 99670, 99730, 99840, 100010, 100100, 100190, 100300, 
    100390, 100460, 100550, 100630, 100710, 100800, 100890, 100970, 101070, 
    101170, 101270, 101350, 101410, 101480, 101530, 101570, 101630, 101680, 
    101760, 101840, 101900, 101970, 102030, 102060, 102090, 102080, 102080, 
    102110, 102140, 102130, 102170, 102180, 102210, 102260, 102270, 102280, 
    102280, 102280, 102250, 102250, 102250, 102230, 102230, 102260, 102250, 
    102260, 102270, 102270, 102260, 102260, 102250, 102230, 102220, 102230, 
    102200, 102190, 102200, 102220, 102220, 102200, 102160, 102140, 102120, 
    102090, 102030, 101990, 101960, 101940, 101910, 101900, 101880, 101850, 
    101800, 101790, 101760, 101720, 101680, 101660, 101660, 101670, 101650, 
    101650, 101610, 101570, 101540, 101520, 101510, 101500, 101500, 101480, 
    101480, 101490, 101510, 101530, 101550, 101540, 101590, 101610, 101630, 
    101630, 101650, 101700, 101740, 101760, 101800, 101820, 101840, 101870, 
    101890, 101910, 101950, 101950, 101940, 101930, 101890, 101890, 101900, 
    101910, 101910, 101910, 101900, 101930, 101950, 101990, 102000, 102010, 
    102040, 102060, 102070, 102040, 102010, 102010, 102030, 102030, 102020, 
    102000, 101980, 101960, 101930, 101920, 101890, 101860, 101830, 101840, 
    101830, 101800, 101800, 101780, 101750, 101720, 101710, 101700, 101700, 
    101690, 101680, 101640, 101630, 101600, 101590, 101590, 101590, 101580, 
    101570, 101510, 101490, 101480, 101490, 101470, 101450, 101400, 101380, 
    101350, 101320, 101320, 101320, 101320, 101290, 101300, 101270, 101260, 
    101260, 101260, 101240, 101230, 101250, 101230, 101230, 101200, 101230, 
    101200, 101240, 101240, 101180, 101190, 101160, 101130, 101140, 101130, 
    101130, 101150, 101170, 101210, 101230, 101260, 101280, 101310, 101310, 
    101340, 101360, 101380, 101400, 101400, 101440, 101480, 101500, 101560, 
    101560, 101560, 101580, 101590, 101630, 101680, 101700, 101690, 101730, 
    101770, 101820, 101840, 101860, 101880, 101910, 101930, 101970, 102030, 
    102020, 102070, 102100, 102110, 102140, 102170, 102200, 102200, 102230, 
    102240, 102250, 102280, 102280, 102300, 102300, 102300, 102290, 102280, 
    102250, 102260, 102240, 102220, 102190, 102200, 102160, 102140, 102110, 
    102080, 102060, 102030, 102000, 101990, 101960, 101960, 101940, 101930, 
    101910, 101890, 101870, 101860, 101870, 101880, 101860, 101840, 101800, 
    101790, 101790, 101780, 101760, 101740, 101730, 101720, 101680, 101660, 
    101630, 101600, 101540, 101510, 101450, 101440, 101400, 101370, 101320, 
    101300, 101280, 101250, 101180, 101120, 101040, 100980, 100940, 100880, 
    100820, 100780, 100750, 100710, 100690, 100670, 100660, 100670, 100670, 
    100700, 100720, 100790, 100820, 100870, 100940, 100960, 101020, 101060, 
    101110, 101170, 101200, 101270, 101300, 101330, 101370, 101390, 101400, 
    101430, 101460, 101480, 101520, 101510, 101480, 101450, 101410, 101380, 
    101390, 101390, 101370, 101330, 101290, 101230, 101210, 101180, 101150, 
    101150, 101130, 101100, 101120, 101140, 101170, 101190, 101200, 101180, 
    101190, 101160, 101170, 101160, 101140, 101160, 101200, 101230, 101300, 
    101430, 101550, 101680, 101810, 101950, 102050, 102180, 102300, 102380, 
    102470, 102560, 102630, 102700, 102770, 102850, 102900, 102950, 103000, 
    103010, 103020, 103050, 103030, 103070, 103090, 103100, 103130, 103120, 
    103110, 103090, 103080, 103040, 103030, 103010, 103000, 102990, 102980, 
    102980, 102990, 102970, 102970, 102950, 102940, 102910, 102930, 102910, 
    102890, 102890, 102870, 102880, 102870, 102870, 102860, 102840, 102810, 
    102760, 102730, 102670, 102630, 102600, 102560, 102510, 102460, 102420, 
    102360, 102280, 102230, 102170, 102120, 102070, 102000, 101950, 101890, 
    101870, 101850, 101830, 101820, 101790, 101780, 101760, 101750, 101720, 
    101710, 101720, 101710, 101700, 101670, 101650, 101620, 101550, 101450, 
    101350, 101170, 101070, 100990, 101010, 101010, 101040, 101060, 101040, 
    101040, 100970, 100910, 100910, 100880, 100880, 100990, 101010, 101100, 
    101180, 101310, 101400, 101470, 101580, 101660, 101740, 101800, 101870, 
    101940, 102050, 102140, 102230, 102340, 102440, 102490, 102570, 102670, 
    102710, 102730, 102790, 102850, 102880, 102890, 102870, 102870, 102830, 
    102800, 102730, 102640, 102580, 102550, 102540, 102520, 102490, 102500, 
    102480, 102500, 102480, 102440, 102360, 102320, 102220, 102100, 102000, 
    101980, 101900, 101850, 101890, 101840, 101860, 101850, 101840, 101890, 
    101940, 101970, 101990, 102030, 102070, 102080, 102120, 102180, 102240, 
    102270, 102290, 102300, 102300, 102310, 102340, 102370, 102370, 102390, 
    102410, 102390, 102400, 102370, 102340, 102310, 102340, 102370, 102410, 
    102420, 102480, 102520, 102550, 102580, 102570, 102560, 102550, 102580, 
    102580, 102590, 102610, 102620, 102650, 102680, 102690, 102710, 102730, 
    102750, 102760, 102770, 102760, 102730, 102760, 102800, 102820, 102890, 
    102960, 102970, 102920, 102900, 102900, 102890, 102890, 102890, 102900, 
    102920, 102910, 102900, 102910, 102920, 102940, 102940, 102950, 102960, 
    102930, 102950, 102880, 102890, 102880, 102860, 102820, 102780, 102730, 
    102690, 102650, 102620, 102590, 102590, 102610, 102610, 102610, 102580, 
    102560, 102540, 102530, 102520, 102510, 102500, 102530, 102540, 102560, 
    102580, 102630, 102660, 102660, 102640, 102660, 102670, 102680, 102670, 
    102680, 102690, 102690, 102680, 102660, 102610, 102600, 102540, 102520, 
    102500, 102500, 102440, 102430, 102400, 102340, 102370, 102370, 102350, 
    102300, 102260, 102210, 102190, 102150, 102110, 102090, 102080, 102110, 
    102080, 102030, 102030, 102010, 101970, 101930, 101890, 101860, 101820, 
    101790, 101710, 101650, 101570, 101540, 101490, 101450, 101400, 101350, 
    101290, 101210, 101130, 101070, 101010, 100960, 100920, 100880, 100810, 
    100790, 100780, 100730, 100640, 100540, 100490, 100490, 100510, 100480, 
    100430, 100340, 100350, 100360, 100310, 100280, 100250, 100230, 100210, 
    100190, 100180, 100150, 100140, 100130, 100110, 100110, 100100, 100100, 
    100080, 100060, 100020, 100000, 100000, 99990, 99990, 100010, 99990, 
    99990, 99980, 99990, 100000, 100000, 100010, 100040, 100070, 100090, 
    100100, 100110, 100150, 100170, 100190, 100200, 100220, 100200, 100210, 
    100210, 100210, 100220, 100250, 100280, 100310, 100330, 100360, 100360, 
    100360, 100380, 100400, 100420, 100440, 100480, 100500, 100530, 100570, 
    100600, 100640, 100680, 100710, 100750, 100780, 100820, 100840, 100860, 
    100910, 100960, 101010, 101060, 101080, 101120, 101160, 101190, 101240, 
    101280, 101290, 101320, 101350, 101370, 101400, 101410, 101410, 101410, 
    101430, 101440, 101430, 101450, 101460, 101460, 101470, 101490, 101510, 
    101530, 101530, 101540, 101540, 101560, 101580, 101590, 101580, 101570, 
    101590, 101580, 101590, 101600, 101620, 101610, 101600, 101590, 101600, 
    101600, 101600, 101580, 101580, 101590, 101610, 101620, 101610, 101620, 
    101630, 101620, 101600, 101570, 101580, 101570, 101570, 101560, 101570, 
    101580, 101560, 101530, 101530, 101520, 101510, 101510, 101510, 101480, 
    101470, 101470, 101480, 101530, 101580, 101600, 101640, 101650, 101680, 
    101710, 101730, 101730, 101750, 101770, 101780, 101780, 101780, 101780, 
    101780, 101760, 101740, 101740, 101740, 101740, 101740, 101730, 101750, 
    101780, 101810, 101820, 101810, 101810, 101810, 101820, 101820, 101820, 
    101820, 101830, 101840, 101850, 101850, 101840, 101830, 101800, 101790, 
    101790, 101780, 101800, 101800, 101790, 101800, 101810, 101790, 101780, 
    101770, 101770, 101750, 101730, 101730, 101730, 101730, 101730, 101720, 
    101700, 101700, 101700, 101670, 101630, 101600, 101580, 101560, 101560, 
    101560, 101540, 101550, 101590, 101610, 101600, 101570, 101560, 101550, 
    101540, 101530, 101510, 101500, 101490, 101470, 101450, 101440, 101430, 
    101430, 101440, 101440, 101430, 101430, 101440, 101450, 101480, 101500, 
    101530, 101530, 101530, 101470, 101460, 101440, 101400, 101380, 101380, 
    101340, 101340, 101350, 101340, 101330, 101300, 101280, 101240, 101230, 
    101200, 101160, 101200, 101170, 101190, 101170, 101150, 101170, 101170, 
    101160, 101170, 101140, 101090, 101070, 101090, 101050, 101050, 101070, 
    101080, 101100, 101120, 101130, 101160, 101170, 101180, 101150, 101180, 
    101200, 101210, 101240, 101240, 101260, 101250, 101230, 101230, 101200, 
    101180, 101160, 101130, 101100, 101060, 101050, 101030, 101010, 100970, 
    100960, 100920, 100880, 100810, 100810, 100790, 100770, 100760, 100750, 
    100760, 100750, 100750, 100720, 100720, 100720, 100730, 100750, 100760, 
    100790, 100820, 100840, 100860, 100860, 100860, 100890, 100890, 100920, 
    100940, 100980, 101020, 101070, 101110, 101160, 101200, 101220, 101240, 
    101270, 101310, 101330, 101350, 101380, 101400, 101450, 101490, 101510, 
    101530, 101550, 101590, 101610, 101630, 101660, 101680, 101720, 101750, 
    101790, 101820, 101850, 101890, 101910, 101940, 101970, 101980, 102000, 
    102000, 102000, 102020, 102020, 102030, 102020, 102050, 102050, 102020, 
    102020, 102020, 102030, 102020, 102010, 102000, 101990, 101990, 101990, 
    101980, 102000, 101970, 101960, 101940, 101910, 101860, 101810, 101760, 
    101710, 101670, 101630, 101590, 101530, 101480, 101440, 101400, 101390, 
    101350, 101350, 101340, 101340, 101350, 101370, 101400, 101420, 101450, 
    101470, 101500, 101520, 101540, 101570, 101600, 101590, 101630, 101640, 
    101660, 101680, 101690, 101700, 101690, 101720, 101720, 101730, 101740, 
    101740, 101760, 101780, 101790, 101780, 101790, 101810, 101810, 101810, 
    101840, 101850, 101850, 101870, 101900, 101910, 101940, 101950, 101970, 
    101950, 101960, 101970, 101970, 101970, 101930, 101900, 101870, 101840, 
    101830, 101770, 101740, 101700, 101610, 101560, 101530, 101460, 101400, 
    101340, 101300, 101240, 101180, 101180, 101140, 101070, 100990, 100990, 
    100960, 100930, 100930, 100900, 100840, 100800, 100770, 100740, 100740, 
    100690, 100670, 100690, 100720, 100740, 100790, 100840, 100870, 100920, 
    100980, 101030, 101060, 101100, 101150, 101180, 101170, 101180, 101160, 
    101150, 101160, 101150, 101120, 101100, 101050, 100990, 100980, 100910, 
    100860, 100790, 100760, 100720, 100710, 100700, 100690, 100650, 100660, 
    100640, 100650, 100640, 100640, 100600, 100620, 100620, 100630, 100620, 
    100640, 100650, 100670, 100670, 100620, 100590, 100600, 100570, 100540, 
    100520, 100560, 100560, 100540, 100540, 100490, 100440, 100420, 100400, 
    100390, 100310, 100240, 100150, 100130, 100070, 100020, 99910, 99800, 
    99700, 99620, 99540, 99450, 99390, 99300, 99210, 99110, 99010, 98900, 
    98840, 98780, 98720, 98640, 98570, 98500, 98490, 98480, 98500, 98500, 
    98500, 98510, 98530, 98550, 98540, 98550, 98550, 98590, 98610, 98640, 
    98640, 98660, 98680, 98740, 98750, 98750, 98740, 98760, 98820, 98860, 
    98850, 98890, 98930, 98950, 99000, 99030, 99080, 99130, 99180, 99190, 
    99160, 99180, 99170, 99140, 99190, 99210, 99290, 99330, 99360, 99370, 
    99320, 99360, 99520, 99400, 99530, 99530, 99630, 99630, 99630, 99650, 
    99690, 99690, 99590, 99510, 99590, 99530, 99530, 99590, 99540, 99600, 
    99630, 99700, 99670, 99680, 99630, 99620, 99600, 99600, 99580, 99550, 
    99560, 99570, 99580, 99580, 99670, 99680, 99700, 99690, 99690, 99690, 
    99690, 99710, 99700, 99700, 99710, 99690, 99650, 99650, 99630, 99620, 
    99640, 99630, 99630, 99630, 99630, 99660, 99670, 99690, 99730, 99750, 
    99770, 99750, 99750, 99740, 99750, 99780, 99780, 99750, 99750, 99740, 
    99760, 99780, 99760, 99730, 99730, 99710, 99700, 99700, 99680, 99680, 
    99680, 99700, 99680, 99650, 99640, 99590, 99550, 99490, 99470, 99420, 
    99390, 99360, 99320, 99260, 99200, 99170, 99140, 99080, 99000, 98970, 
    98940, 98890, 98860, 98830, 98790, 98760, 98730, 98670, 98630, 98600, 
    98570, 98530, 98490, 98470, 98440, 98420, 98390, 98380, 98360, 98360, 
    98330, 98290, 98280, 98280, 98260, 98260, 98270, 98280, 98300, 98320, 
    98320, 98330, 98340, 98310, 98320, 98320, 98270, 98270, 98230, 98260, 
    98260, 98260, 98260, 98260, 98290, 98290, 98330, 98370, 98420, 98490, 
    98590, 98720, 98900, 99020, 99120, 99180, 99290, 99390, 99450, 99510, 
    99550, 99650, 99700, 99750, 99790, 99870, 99920, 99980, 99970, 100050, 
    100040, 100070, 100100, 100150, 100190, 100240, 100310, 100390, 100460, 
    100490, 100550, 100580, 100640, 100700, 100750, 100760, 100810, 100860, 
    100910, 100950, 100990, 101020, 101040, 101080, 101130, 101160, 101180, 
    101200, 101240, 101280, 101320, 101360, 101390, 101440, 101450, 101470, 
    101500, 101540, 101580, 101600, 101640, 101680, 101710, 101750, 101800, 
    101800, 101820, 101850, 101890, 101930, 101970, 101990, 102010, 102040, 
    102080, 102130, 102180, 102220, 102220, 102260, 102270, 102280, 102280, 
    102270, 102270, 102270, 102240, 102210, 102210, 102170, 102180, 102120, 
    102080, 102040, 101990, 101950, 101900, 101830, 101840, 101800, 101720, 
    101690, 101660, 101620, 101580, 101510, 101410, 101360, 101270, 101200, 
    101180, 101170, 101100, 101030, 101020, 100920, 100870, 100810, 100750, 
    100670, 100600, 100620, 100610, 100560, 100540, 100520, 100500, 100450, 
    100460, 100470, 100490, 100480, 100450, 100430, 100420, 100440, 100400, 
    100410, 100390, 100370, 100430, 100490, 100540, 100600, 100610, 100580, 
    100550, 100530, 100500, 100500, 100540, 100550, 100480, 100450, 100460, 
    100430, 100430, 100400, 100380, 100340, 100300, 100300, 100290, 100290, 
    100240, 100170, 100140, 100120, 100050, 100050, 99980, 100000, 100020, 
    100010, 100020, 100020, 100020, 100010, 99970, 99940, 99960, 99970, 
    99990, 100000, 99990, 100010, 100020, 100020, 100000, 100000, 99990, 
    99980, 99970, 99990, 100030, 100060, 100080, 100110, 100080, 100090, 
    100120, 100130, 100130, 100150, 100160, 100160, 100170, 100170, 100190, 
    100230, 100230, 100250, 100260, 100280, 100280, 100290, 100300, 100310, 
    100330, 100340, 100330, 100330, 100360, 100370, 100380, 100370, 100380, 
    100390, 100410, 100420, 100440, 100460, 100460, 100480, 100500, 100530, 
    100530, 100550, 100570, 100590, 100610, 100620, 100640, 100660, 100690, 
    100690, 100690, 100730, 100740, 100750, 100750, 100740, 100740, 100750, 
    100740, 100740, 100760, 100780, 100820, 100850, 100860, 100880, 100880, 
    100880, 100940, 100970, 101000, 101030, 101070, 101110, 101150, 101180, 
    101200, 101210, 101210, 101200, 101240, 101280, 101320, 101330, 101360, 
    101370, 101400, 101410, 101430, 101430, 101440, 101440, 101450, 101510, 
    101530, 101550, 101550, 101540, 101530, 101540, 101540, 101540, 101560, 
    101540, 101570, 101570, 101590, 101600, 101590, 101590, 101580, 101580, 
    101580, 101590, 101570, 101550, 101540, 101520, 101520, 101520, 101490, 
    101480, 101480, 101460, 101440, 101450, 101470, 101480, 101490, 101500, 
    101510, 101530, 101540, 101540, 101540, 101570, 101550, 101580, 101590, 
    101620, 101650, 101760, 101750, 101830, 101870, 101910, 101980, 102000, 
    102030, 102070, 102080, 102100, 102110, 102150, 102190, 102240, 102250, 
    102280, 102300, 102330, 102310, 102330, 102330, 102370, 102380, 102410, 
    102460, 102490, 102530, 102560, 102590, 102600, 102620, 102610, 102610, 
    102600, 102620, 102630, 102680, 102710, 102740, 102750, 102760, 102780, 
    102820, 102830, 102840, 102840, 102880, 102950, 103000, 103030, 103050, 
    103070, 103110, 103150, 103200, 103250, 103280, 103330, 103360, 103380, 
    103450, 103500, 103530, 103540, 103530, 103550, 103570, 103570, 103620, 
    103640, 103670, 103740, 103770, 103800, 103850, 103830, 103820, 103800, 
    103810, 103750, 103740, 103710, 103710, 103730, 103750, 103760, 103770, 
    103760, 103730, 103720, 103700, 103690, 103690, 103670, 103670, 103680, 
    103710, 103740, 103770, 103770, 103790, 103820, 103810, 103810, 103820, 
    103840, 103860, 103870, 103850, 103860, 103840, 103820, 103810, 103780, 
    103810, 103780, 103730, 103710, 103700, 103720, 103730, 103720, 103690, 
    103640, 103610, 103610, 103620, 103570, 103540, 103520, 103500, 103470, 
    103460, 103410, 103380, 103350, 103310, 103290, 103270, 103250, 103180, 
    103170, 103150, 103140, 103130, 103120, 103070, 103040, 103010, 102980, 
    102950, 102920, 102900, 102880, 102850, 102830, 102780, 102750, 102720, 
    102680, 102640, 102610, 102540, 102500, 102460, 102400, 102350, 102290, 
    102270, 102260, 102230, 102160, 102110, 102020, 101970, 101910, 101870, 
    101830, 101790, 101740, 101700, 101650, 101610, 101580, 101520, 101470, 
    101410, 101350, 101290, 101230, 101190, 101160, 101120, 101090, 101050, 
    101000, 100940, 100880, 100820, 100780, 100730, 100690, 100650, 100610, 
    100600, 100570, 100520, 100490, 100420, 100380, 100350, 100320, 100290, 
    100300, 100320, 100320, 100360, 100410, 100450, 100470, 100500, 100520, 
    100560, 100590, 100610, 100650, 100690, 100730, 100760, 100810, 100830, 
    100840, 100870, 100910, 100960, 100980, 100980, 101000, 101010, 101030, 
    101040, 101070, 101060, 101060, 101070, 101130, 101140, 101120, 101140, 
    101180, 101250, 101300, 101300, 101330, 101340, 101360, 101360, 101350, 
    101340, 101340, 101330, 101320, 101300, 101280, 101280, 101310, 101300, 
    101300, 101290, 101280, 101280, 101290, 101300, 101300, 101300, 101300, 
    101260, 101250, 101250, 101230, 101190, 101150, 101110, 101060, 101030, 
    101000, 100970, 100930, 100880, 100860, 100850, 100790, 100670, 100580, 
    100490, 100390, 100360, 100320, 100220, 100120, 100020, 99900, 99800, 
    99720, 99590, 99460, 99380, 99340, 99280, 99300, 99280, 99280, 99300, 
    99310, 99270, 99250, 99230, 99200, 99160, 99130, 99090, 99070, 99050, 
    99070, 99050, 99050, 99050, 99050, 99030, 99020, 99010, 99010, 99020, 
    99010, 98980, 98970, 98950, 98940, 98940, 98900, 98840, 98850, 98800, 
    98760, 98760, 98710, 98680, 98670, 98650, 98660, 98680, 98670, 98650, 
    98630, 98600, 98590, 98560, 98560, 98560, 98560, 98570, 98590, 98580, 
    98560, 98580, 98570, 98630, 98660, 98710, 98830, 98900, 99000, 99060, 
    99140, 99240, 99310, 99430, 99510, 99570, 99620, 99670, 99740, 99770, 
    99820, 99870, 99910, 99950, 100000, 100030, 100100, 100120, 100200, 
    100230, 100270, 100300, 100350, 100360, 100390, 100420, 100430, 100440, 
    100430, 100460, 100470, 100470, 100480, 100520, 100540, 100550, 100560, 
    100570, 100590, 100580, 100600, 100600, 100590, 100610, 100620, 100650, 
    100660, 100670, 100660, 100670, 100660, 100640, 100630, 100620, 100620, 
    100610, 100620, 100640, 100640, 100670, 100680, 100710, 100740, 100750, 
    100780, 100810, 100840, 100860, 100870, 100880, 100890, 100920, 100950, 
    100930, 100950, 100970, 100980, 101010, 101000, 101010, 101050, 101040, 
    101070, 101090, 101110, 101110, 101120, 101100, 101100, 101090, 101080, 
    101070, 101080, 101080, 101080, 101130, 101190, 101200, 101200, 101250, 
    101290, 101300, 101300, 101350, 101370, 101380, 101420, 101480, 101530, 
    101530, 101560, 101570, 101610, 101620, 101660, 101690, 101760, 101810, 
    101850, 101900, 101930, 101950, 101900, 101900, 101910, 101890, 101890, 
    101920, 101940, 101930, 101950, 101980, 102020, 102040, 102020, 101990, 
    101950, 101890, 101860, 101830, 101820, 101790, 101770, 101770, 101750, 
    101710, 101660, 101630, 101600, 101550, 101510, 101480, 101460, 101440, 
    101410, 101410, 101390, 101380, 101350, 101330, 101290, 101280, 101220, 
    101210, 101200, 101200, 101180, 101180, 101190, 101220, 101220, 101260, 
    101250, 101250, 101250, 101240, 101230, 101200, 101170, 101160, 101200, 
    101140, 101060, 100990, 100940, 100910, 100870, 100850, 100840, 100810, 
    100790, 100740, 100690, 100640, 100620, 100610, 100560, 100550, 100490, 
    100450, 100430, 100350, 100290, 100240, 100190, 100130, 100070, 100020, 
    99990, 99910, 99890, 99830, 99800, 99750, 99710, 99650, 99640, 99620, 
    99560, 99530, 99470, 99430, 99420, 99380, 99360, 99330, 99320, 99300, 
    99270, 99250, 99260, 99240, 99240, 99250, 99280, 99320, 99340, 99350, 
    99360, 99370, 99400, 99380, 99400, 99380, 99410, 99410, 99460, 99460, 
    99520, 99550, 99580, 99590, 99630, 99620, 99700, 99760, 99810, 99820, 
    99900, 99930, 99930, 100060, 100060, 100110, 100130, 100140, 100170, 
    100160, 100170, 100180, 100190, 100170, 100170, 100200, 100210, 100240, 
    100270, 100260, 100260, 100260, 100250, 100250, 100250, 100250, 100240, 
    100240, 100240, 100240, 100250, 100240, 100240, 100230, 100220, 100210, 
    100200, 100180, 100160, 100160, 100150, 100150, 100150, 100120, 100110, 
    100080, 100080, 100070, 100040, 100040, 100020, 100020, 99990, 99960, 
    99940, 99910, 99890, 99880, 99840, 99830, 99810, 99830, 99740, 99700, 
    99700, 99740, 99740, 99740, 99750, 99760, 99760, 99760, 99790, 99830, 
    99890, 99930, 99970, 99990, 100030, 100060, 100080, 100120, 100170, 
    100220, 100240, 100260, 100280, 100310, 100350, 100380, 100410, 100460, 
    100490, 100540, 100560, 100560, 100570, 100600, 100600, 100570, 100540, 
    100530, 100520, 100530, 100540, 100530, 100490, 100430, 100350, 100270, 
    100150, 100030, 99910, 99850, 99680, 99570, 99410, 99140, 98890, 98600, 
    98250, 97960, 97580, 97220, 96930, 96710, 96510, 96290, 96120, 95920, 
    95800, 95720, 95660, 95590, 95550, 95490, 95460, 95480, 95530, 95580, 
    95640, 95730, 95800, 95850, 95860, 95830, 95830, 95920, 96020, 96100, 
    96170, 96230, 96310, 96380, 96390, 96560, 96620, 96680, 96700, 96740, 
    96800, 96850, 96910, 96980, 97050, 97120, 97200, 97290, 97360, 97450, 
    97540, 97600, 97680, 97760, 97830, 97900, 97950, 98010, 98100, 98160, 
    98250, 98340, 98370, 98430, 98510, 98620, 98690, 98760, 98810, 98890, 
    98930, 98960, 98970, 99020, 99010, 99010, 98990, 98980, 98970, 98950, 
    98930, 98900, 98890, 98910, 98930, 98960, 98990, 99030, 99090, 99140, 
    99180, 99230, 99220, 99230, 99280, 99360, 99420, 99490, 99570, 99620, 
    99660, 99750, 99820, 99850, 99890, 99950, 100020, 100050, 100110, 100150, 
    100180, 100220, 100230, 100260, 100310, 100310, 100330, 100350, 100360, 
    100400, 100400, 100430, 100420, 100430, 100430, 100470, 100500, 100520, 
    100570, 100590, 100650, 100690, 100720, 100760, 100810, 100860, 100920, 
    100990, 101080, 101120, 101190, 101240, 101330, 101370, 101390, 101440, 
    101470, 101490, 101480, 101510, 101560, 101600, 101650, 101670, 101690, 
    101690, 101660, 101700, 101690, 101680, 101700, 101700, 101690, 101660, 
    101610, 101470, 101370, 101250, 101150, 100980, 100860, 100750, 100650, 
    100630, 100600, 100570, 100510, 100510, 100480, 100520, 100530, 100510, 
    100490, 100560, 100620, 100620, 100620, 100620, 100600, 100530, 100510, 
    100510, 100440, 100380, 100280, 100130, 99940, 99780, 99580, 99350, 
    99110, 98850, 98540, 98290, 98390, 98590, 98690, 98650, 98680, 98760, 
    98790, 98780, 98830, 98900, 98910, 98950, 99000, 98990, 99050, 99110, 
    99170, 99250, 99330, 99420, 99530, 99610, 99670, 99730, 99800, 99840, 
    99910, 99970, 100010, 100080, 100170, 100240, 100310, 100380, 100420, 
    100490, 100530, 100570, 100650, 100700, 100720, 100760, 100830, 100870, 
    100910, 100960, 100970, 100960, 100970, 101000, 101000, 100990, 101010, 
    101060, 101070, 101070, 101080, 101080, 101060, 101040, 101040, 101020, 
    101030, 101010, 100990, 100960, 100950, 100960, 100940, 100920, 100900, 
    100860, 100860, 100850, 100850, 100870, 100870, 100890, 100900, 100920, 
    100930, 100920, 100910, 100910, 100910, 100910, 100900, 100890, 100890, 
    100870, 100850, 100860, 100840, 100800, 100780, 100780, 100760, 100720, 
    100700, 100680, 100660, 100680, 100670, 100650, 100610, 100580, 100550, 
    100520, 100490, 100510, 100480, 100480, 100490, 100500, 100510, 100520, 
    100520, 100530, 100500, 100510, 100510, 100490, 100470, 100480, 100500, 
    100510, 100550, 100580, 100580, 100600, 100600, 100620, 100620, 100630, 
    100640, 100650, 100660, 100670, 100670, 100680, 100690, 100680, 100660, 
    100650, 100650, 100650, 100650, 100670, 100670, 100710, 100730, 100740, 
    100750, 100780, 100800, 100790, 100810, 100810, 100810, 100820, 100830, 
    100830, 100840, 100830, 100840, 100840, 100830, 100830, 100820, 100800, 
    100790, 100790, 100780, 100800, 100830, 100850, 100820, 100830, 100830, 
    100780, 100810, 100800, 100800, 100820, 100830, 100840, 100840, 100850, 
    100890, 100900, 100890, 100880, 100860, 100850, 100860, 100870, 100900, 
    100920, 100930, 100890, 100890, 100840, 100810, 100750, 100700, 100630, 
    100590, 100560, 100530, 100500, 100470, 100440, 100370, 100330, 100240, 
    100220, 100180, 100150, 100130, 100130, 100150, 100180, 100280, 100280, 
    100340, 100320, 100320, 100300, 100370, 100400, 100450, 100460, 100460, 
    100460, 100480, 100410, 100360, 100350, 100310, 100250, 100190, 100140, 
    100090, 100070, 99990, 100000, 99990, 99950, 99890, 99840, 99820, 99830, 
    99810, 99810, 99830, 99810, 99830, 99850, 99900, 99870, 99870, 99890, 
    99950, 99990, 100050, 100070, 100110, 100190, 100290, 100380, 100500, 
    100550, 100620, 100710, 100770, 100810, 100840, 100890, 100950, 101000, 
    101040, 101060, 101060, 101080, 101090, 101150, 101140, 101150, 101160, 
    101170, 101200, 101200, 101210, 101220, 101240, 101230, 101220, 101240, 
    101260, 101290, 101260, 101300, 101320, 101360, 101370, 101380, 101370, 
    101400, 101400, 101380, 101410, 101430, 101440, 101430, 101410, 101420, 
    101430, 101430, 101450, 101470, 101490, 101460, 101460, 101460, 101460, 
    101480, 101480, 101500, 101520, 101540, 101560, 101540, 101550, 101560, 
    101540, 101540, 101530, 101520, 101540, 101530, 101550, 101600, 101630, 
    101630, 101640, 101660, 101640, 101590, 101580, 101520, 101490, 101440, 
    101380, 101340, 101310, 101260, 101200, 101150, 101080, 101030, 100940, 
    100900, 100850, 100790, 100730, 100700, 100710, 100720, 100730, 100770, 
    100830, 100870, 100920, 100950, 100990, 101020, 100970, 100940, 100890, 
    100800, 100720, 100600, 100480, 100380, 100300, 100200, 100090, 100010, 
    99920, 99780, 99690, 99540, 99510, 99450, 99320, 99230, 99190, 99100, 
    99010, 98930, 98830, 98750, 98710, 98700, 98770, 98860, 98920, 98980, 
    99140, 99170, 99250, 99320, 99370, 99440, 99450, 99490, 99530, 99560, 
    99550, 99530, 99460, 99430, 99400, 99380, 99360, 99370, 99350, 99330, 
    99270, 99230, 99190, 99180, 99190, 99200, 99190, 99200, 99240, 99280, 
    99320, 99360, 99390, 99390, 99380, 99480, 99490, 99510, 99540, 99580, 
    99610, 99650, 99700, 99740, 99750, 99750, 99750, 99720, 99720, 99710, 
    99740, 99620, 99690, 99710, 99730, 99720, 99730, 99740, 99770, 99780, 
    99810, 99830, 99850, 99780, 99840, 99890, 99930, 99950, 100010, 100060, 
    100100, 100160, 100210, 100260, 100290, 100380, 100450, 100530, 100620, 
    100720, 100780, 100830, 100870, 100940, 101010, 101030, 101060, 101090, 
    101110, 101120, 101170, 101230, 101270, 101280, 101310, 101340, 101300, 
    101270, 101250, 101250, 101260, 101270, 101270, 101270, 101220, 101140, 
    101110, 101090, 100990, 100970, 100990, 101030, 101120, 101190, 101310, 
    101410, 101480, 101530, 101570, 101610, 101620, 101630, 101650, 101740, 
    101760, 101770, 101780, 101800, 101820, 101810, 101800, 101790, 101800, 
    101790, 101780, 101790, 101770, 101740, 101740, 101750, 101700, 101660, 
    101630, 101600, 101540, 101490, 101460, 101370, 101300, 101260, 101220, 
    101190, 101180, 101120, 101080, 101060, 101060, 101060, 101080, 101070, 
    101100, 101150, 101210, 101260, 101290, 101320, 101360, 101390, 101420, 
    101450, 101460, 101520, 101560, 101590, 101630, 101650, 101650, 101640, 
    101640, 101640, 101640, 101640, 101640, 101750, 101750, 101740, 101720, 
    101730, 101730, 101700, 101660, 101640, 101600, 101570, 101560, 101610, 
    101610, 101610, 101640, 101670, 101680, 101680, 101690, 101700, 101670, 
    101650, 101670, 101730, 101730, 101730, 101730, 101740, 101740, 101740, 
    101760, 101760, 101770, 101760, 101760, 101780, 101810, 101840, 101860, 
    101860, 101880, 101870, 101840, 101800, 101770, 101760, 101750, 101740, 
    101740, 101730, 101710, 101700, 101640, 101620, 101600, 101580, 101550, 
    101510, 101500, 101450, 101440, 101420, 101400, 101390, 101380, 101370, 
    101330, 101320, 101300, 101260, 101250, 101170, 101170, 101190, 101180, 
    101160, 101160, 101140, 101130, 101130, 101110, 101080, 101060, 101070, 
    101060, 101110, 101140, 101120, 101120, 101100, 101100, 101080, 101100, 
    101110, 101090, 101080, 101080, 101080, 101100, 101100, 101090, 101090, 
    101090, 101070, 101040, 101010, 101020, 100910, 100930, 100920, 100930, 
    100910, 100900, 100930, 100980, 100990, 101010, 101050, 101100, 101070, 
    101070, 101060, 101060, 101110, 101150, 101190, 101210, 101210, 101210, 
    101210, 101190, 101260, 101260, 101280, 101280, 101300, 101280, 101280, 
    101230, 101170, 101130, 101070, 101040, 100970, 100920, 100870, 100830, 
    100800, 100780, 100750, 100700, 100660, 100630, 100600, 100580, 100630, 
    100640, 100640, 100670, 100700, 100720, 100760, 100780, 100780, 100790, 
    100810, 100870, 100960, 101020, 101030, 101080, 101130, 101180, 101230, 
    101250, 101270, 101290, 101310, 101350, 101220, 101270, 101320, 101360, 
    101380, 101400, 101430, 101470, 101470, 101470, 101480, 101520, 101540, 
    101590, 101620, 101630, 101650, 101670, 101700, 101720, 101740, 101760, 
    101770, 101750, 101670, 101690, 101710, 101740, 101770, 101810, 101820, 
    101820, 101780, 101750, 101770, 101820, 101770, 101770, 101760, 101780, 
    101790, 101810, 101810, 101830, 101860, 101860, 101840, 101830, 101790, 
    101840, 101890, 101950, 101990, 101980, 101990, 102050, 102110, 102130, 
    102110, 102100, 102170, 102220, 102270, 102340, 102390, 102420, 102420, 
    102450, 102510, 102550, 102560, 102570, 102590, 102610, 102650, 102680, 
    102730, 102730, 102710, 102690, 102680, 102660, 102650, 102630, 102580, 
    102560, 102550, 102550, 102510, 102480, 102440, 102390, 102320, 102280, 
    102260, 102210, 102120, 102110, 102080, 102040, 102010, 101970, 101930, 
    101900, 101860, 101770, 101720, 101660, 101650, 101630, 101600, 101580, 
    101570, 101550, 101530, 101500, 101440, 101420, 101420, 101420, 101340, 
    101360, 101370, 101390, 101390, 101380, 101360, 101330, 101290, 101280, 
    101230, 101180, 101100, 101050, 101020, 100940, 100850, 100820, 100750, 
    100680, 100610, 100540, 100440, 100350, 100180, 100040, 99930, 99900, 
    99870, 99830, 99780, 99720, 99670, 99660, 99650, 99610, 99440, 99260, 
    99110, 98940, 98740, 98370, 97970, 97650, 97360, 97260, 97330, 97350, 
    97310, 97360, 97450, 97540, 97660, 97820, 97990, 98120, 98240, 98360, 
    98430, 98510, 98600, 98690, 98760, 98810, 98870, 98950, 99030, 99140, 
    99300, 99460, 99640, 99790, 100040, 100230, 100420, 100570, 100650, 
    100690, 100700, 100710, 100700, 100680, 100770, 100900, 101090, 101150, 
    101170, 101190, 101220, 101200, 101160, 101070, 100930, 100770, 100620, 
    100510, 100250, 100110, 99930, 99730, 99510, 99340, 99220, 99100, 99010, 
    98920, 98860, 98790, 98830, 98780, 98740, 98700, 98670, 98640, 98620, 
    98560, 98520, 98490, 98500, 98510, 98580, 98590, 98630, 98680, 98720, 
    98790, 98840, 98890, 98960, 99010, 99030, 99060, 99160, 99200, 99230, 
    99260, 99270, 99260, 99270, 99270, 99250, 99200, 99160, 99130, 99300, 
    99330, 99390, 99430, 99480, 99540, 99610, 99670, 99710, 99710, 99710, 
    99760, 99780, 99770, 99750, 99700, 99630, 99530, 99540, 99520, 99530, 
    99520, 99480, 99460, 99460, 99470, 99420, 99360, 99310, 99220, 99080, 
    98890, 98750, 98650, 98540, 98480, 98450, 98510, 98640, 98790, 98910, 
    99060, 99200, 99260, 99260, 99270, 99260, 99310, 99160, 99040, 99180, 
    99440, 99680, 99800, 99930, 100020, 100130, 100240, 100360, 100450, 
    100500, 100560, 100620, 100670, 100700, 100730, 100770, 100800, 100830, 
    100880, 100920, 100950, 100930, 100960, 101000, 101060, 101100, 101120, 
    101130, 101140, 101160, 101180, 101190, 101210, 101290, 101310, 101350, 
    101370, 101380, 101400, 101430, 101440, 101450, 101430, 101420, 101420, 
    101400, 101400, 101430, 101450, 101460, 101470, 101450, 101420, 101380, 
    101350, 101350, 101360, 101350, 101360, 101360, 101350, 101340, 101340, 
    101340, 101350, 101370, 101370, 101360, 101330, 101350, 101370, 101410, 
    101440, 101470, 101490, 101500, 101510, 101510, 101510, 101510, 101530, 
    101580, 101580, 101570, 101550, 101560, 101590, 101600, 101610, 101620, 
    101610, 101600, 101610, 101700, 101720, 101760, 101760, 101780, 101800, 
    101810, 101830, 101840, 101880, 101880, 101890, 101890, 101930, 101960, 
    101980, 102000, 102020, 102050, 102090, 102090, 102070, 102060, 102070, 
    102170, 102200, 102220, 102260, 102300, 102340, 102380, 102390, 102380, 
    102390, 102390, 102430, 102480, 102500, 102520, 102560, 102570, 102580, 
    102600, 102630, 102650, 102660, 102660, 102680, 102650, 102670, 102700, 
    102740, 102780, 102820, 102840, 102880, 102930, 102970, 103020, 103040, 
    103020, 103060, 103100, 103120, 103150, 103170, 103170, 103190, 103220, 
    103220, 103220, 103210, 103180, 103200, 103210, 103240, 103260, 103270, 
    103280, 103290, 103290, 103290, 103280, 103270, 103230, 103220, 103210, 
    103220, 103220, 103210, 103200, 103200, 103210, 103200, 103180, 103150, 
    103210, 103210, 103220, 103240, 103270, 103260, 103250, 103250, 103240, 
    103220, 103190, 103160, 103150, 103110, 103080, 103060, 103040, 103010, 
    103010, 103010, 103010, 102990, 102960, 102940, 103000, 102990, 102990, 
    102990, 103000, 103020, 103030, 103030, 103050, 103060, 103070, 103090, 
    103170, 103220, 103230, 103210, 103200, 103220, 103260, 103290, 103260, 
    103230, 103220, 103230, 103220, 103210, 103210, 103260, 103290, 103310, 
    103310, 103320, 103310, 103310, 103310, 103330, 103300, 103340, 103370, 
    103400, 103420, 103430, 103470, 103480, 103480, 103470, 103460, 103440, 
    103460, 103480, 103510, 103510, 103520, 103520, 103520, 103540, 103540, 
    103550, 103540, 103570, 103670, 103690, 103720, 103720, 103690, 103700, 
    103690, 103660, 103650, 103610, 103560, 103510, 103430, 103400, 103380, 
    103400, 103380, 103370, 103360, 103350, 103320, 103290, 103270, 103250, 
    103270, 103250, 103240, 103260, 103280, 103340, 103400, 103470, 103550, 
    103610, 103710, 103800, 103860, 103960, 104050, 104120, 104200, 104150, 
    104230, 104290, 104300, 104310, 104310, 104350, 104360, 104400, 104450, 
    104470, 104490, 104490, 104470, 104390, 104380, 104350, 104300, 104240, 
    104220, 104190, 104140, 104080, 104000, 103930, 103900, 103870, 103780, 
    103730, 103720, 103720, 103770, 103670, 103610, 103590, 103590, 103580, 
    103590, 103640, 103690, 103720, 103710, 103700, 103840, 103880, 103860, 
    103870, 103860, 103770, 103660, 103570, 103430, 103360, 103260, 103220, 
    103190, 103210, 103150, 103060, 102990, 102960, 102880, 102760, 102650, 
    102550, 102440, 102360, 102220, 102120, 102040, 101960, 101840, 101690, 
    101550, 101390, 101280, 101220, 101160, 101130, 101450, 101510, 101600, 
    101690, 101770, 101930, 102110, 102260, 102400, 102500, 102600, 102750, 
    102750, 102850, 102960, 103060, 103040, 103130, 103210, 103260, 103350, 
    103380, 103420, 103470, 103520, 103560, 103580, 103610, 103650, 103680, 
    103660, 103640, 103630, 103610, 103620, 103610, 103610, 103620, 103620, 
    103620, 103630, 103640, 103620, 103610, 103590, 103580, 103610, 103590, 
    103580, 103520, 103540, 103530, 103510, 103510, 103480, 103460, 103450, 
    103410, 103350, 103290, 103250, 103230, 103200, 103180, 103180, 103170, 
    103160, 103130, 103090, 103060, 103020, 103020, 102970, 102940, 102920, 
    102900, 102900, 102900, 102880, 102890, 102900, 102890, 102880, 102880, 
    102910, 102880, 102910, 102940, 102960, 102960, 102990, 102990, 103010, 
    103030, 103030, 103020, 103030, 103010, 103040, 103060, 103090, 103110, 
    103110, 103120, 103140, 103140, 103150, 103170, 103170, 103200, 103220, 
    103250, 103280, 103310, 103300, 103300, 103290, 103300, 103300, 103300, 
    103290, 103280, 103290, 103300, 103310, 103290, 103270, 103240, 103230, 
    103220, 103200, 103190, 103180, 103190, 103190, 103200, 103190, 103180, 
    103160, 103160, 103150, 103140, 103150, 103140, 103150, 103120, 103100, 
    103090, 103080, 103060, 103040, 103030, 103020, 103010, 103000, 102980, 
    102960, 102940, 102940, 102960, 102950, 102960, 102950, 102930, 102920, 
    102910, 102900, 102890, 102870, 102870, 102850, 102860, 102840, 102830, 
    102830, 102810, 102800, 102800, 102780, 102780, 102780, 102790, 102810, 
    102830, 102840, 102840, 102830, 102840, 102840, 102840, 102840, 102820, 
    102820, 102840, 102850, 102860, 102870, 102860, 102850, 102840, 102840, 
    102850, 102840, 102850, 102870, 102870, 102890, 102930, 102930, 102930, 
    102940, 102950, 102950, 102970, 102970, 102970, 102960, 102970, 102990, 
    103020, 103040, 103040, 103040, 103050, 103050, 103060, 103060, 103050, 
    103060, 103080, 103110, 103130, 103130, 103130, 103150, 103160, 103150, 
    103150, 103140, 103150, 103170, 103200, 103200, 103200, 103200, 103200, 
    103180, 103170, 103150, 103150, 103150, 103160, 103160, 103160, 103160, 
    103180, 103180, 103180, 103160, 103160, 103140, 103130, 103130, 103110, 
    103100, 103100, 103100, 103100, 103080, 103050, 103020, 102980, 102960, 
    102940, 102910, 102880, 102840, 102820, 102810, 102810, 102770, 102740, 
    102710, 102670, 102650, 102630, 102610, 102580, 102590, 102600, 102600, 
    102610, 102590, 102550, 102530, 102500, 102470, 102450, 102450, 102440, 
    102440, 102440, 102450, 102470, 102460, 102450, 102460, 102460, 102460, 
    102460, 102460, 102460, 102470, 102470, 102480, 102510, 102530, 102520, 
    102520, 102510, 102510, 102510, 102520, 102510, 102520, 102540, 102560, 
    102570, 102580, 102570, 102570, 102580, 102570, 102580, 102590, 102580, 
    102590, 102590, 102580, 102580, 102600, 102580, 102580, 102580, 102590, 
    102560, 102550, 102570, 102570, 102580, 102610, 102650, 102640, 102680, 
    102670, 102680, 102710, 102710, 102720, 102720, 102740, 102730, 102740, 
    102750, 102750, 102740, 102760, 102740, 102730, 102720, 102710, 102700, 
    102720, 102710, 102710, 102670, 102670, 102660, 102620, 102650, 102600, 
    102570, 102520, 102480, 102400, 102370, 102360, 102320, 102290, 102250, 
    102200, 102140, 102080, 102050, 101990, 101950, 101910, 101870, 101830, 
    101800, 101800, 101770, 101680, 101630, 101590, 101520, 101430, 101310, 
    101230, 101140, 101040, 100930, 100800, 100660, 100490, 100300, 100130, 
    99930, 99720, 99530, 99340, 99160, 98990, 98830, 98680, 98500, 98400, 
    98270, 98200, 98160, 98130, 98120, 98080, 98150, 98240, 98330, 98460, 
    98610, 98730, 98870, 99080, 99360, 99570, 99690, 99940, 100180, 100310, 
    100510, 100670, 100820, 100950, 101080, 101220, 101370, 101500, 101610, 
    101670, 101700, 101790, 101870, 101910, 101930, 101980, 102000, 102030, 
    102050, 102080, 102120, 102130, 102190, 102200, 102220, 102240, 102230, 
    102240, 102230, 102230, 102200, 102190, 102140, 102110, 102070, 102060, 
    102030, 101980, 101930, 101880, 101790, 101730, 101700, 101670, 101610, 
    101590, 101550, 101510, 101450, 101420, 101360, 101310, 101300, 101260, 
    101240, 101180, 101130, 101120, 101080, 101070, 101040, 100990, 100930, 
    100910, 100880, 100850, 100820, 100780, 100780, 100770, 100730, 100740, 
    100750, 100770, 100770, 100770, 100800, 100850, 100880, 100920, 100920, 
    100950, 100960, 101000, 101030, 101060, 101060, 101060, 101060, 101050, 
    101020, 101010, 100990, 100970, 100930, 100890, 100840, 100810, 100770, 
    100740, 100730, 100710, 100710, 100660, 100660, 100640, 100660, 100650, 
    100670, 100680, 100700, 100700, 100700, 100720, 100730, 100740, 100770, 
    100750, 100730, 100720, 100740, 100740, 100740, 100750, 100780, 100810, 
    100830, 100900, 100960, 101040, 101090, 101110, 101160, 101190, 101210, 
    101240, 101230, 101260, 101250, 101300, 101400, 101440, 101460, 101500, 
    101550, 101580, 101590, 101610, 101620, 101600, 101630, 101670, 101690, 
    101750, 101800, 101850, 101880, 101890, 101890, 101910, 101910, 101910, 
    101920, 101920, 101910, 101910, 101910, 101930, 101970, 101990, 102010, 
    102020, 102050, 102050, 102030, 102020, 101990, 101980, 101920, 101880, 
    101840, 101780, 101720, 101690, 101580, 101550, 101550, 101520, 101490, 
    101460, 101440, 101430, 101430, 101460, 101440, 101430, 101400, 101400, 
    101380, 101360, 101350, 101360, 101320, 101310, 101330, 101330, 101330, 
    101310, 101290, 101270, 101250, 101250, 101230, 101200, 101210, 101200, 
    101190, 101180, 101210, 101180, 101210, 101190, 101150, 101100, 101040, 
    101000, 100980, 100940, 100870, 100810, 100760, 100690, 100620, 100570, 
    100530, 100510, 100490, 100490, 100480, 100490, 100540, 100580, 100610, 
    100650, 100700, 100740, 100770, 100810, 100840, 100870, 100920, 100960, 
    101000, 101020, 101050, 101080, 101110, 101120, 101140, 101160, 101190, 
    101190, 101220, 101240, 101270, 101300, 101330, 101340, 101330, 101320, 
    101310, 101330, 101300, 101310, 101300, 101310, 101310, 101320, 101310, 
    101310, 101290, 101280, 101250, 101240, 101230, 101210, 101210, 101190, 
    101190, 101190, 101190, 101180, 101170, 101130, 101120, 101110, 101100, 
    101100, 101100, 101120, 101130, 101140, 101150, 101150, 101160, 101160, 
    101160, 101170, 101180, 101190, 101210, 101240, 101260, 101290, 101310, 
    101330, 101360, 101370, 101380, 101370, 101400, 101430, 101460, 101490, 
    101530, 101580, 101610, 101650, 101670, 101690, 101730, 101760, 101790, 
    101850, 101930, 102020, 102070, 102130, 102190, 102220, 102270, 102320, 
    102350, 102380, 102420, 102460, 102490, 102520, 102550, 102600, 102650, 
    102650, 102670, 102690, 102710, 102740, 102750, 102790, 102850, 102870, 
    102860, 102900, 102920, 102930, 102940, 102920, 102930, 102920, 102930, 
    102950, 102980, 102990, 103000, 102990, 103020, 103000, 102980, 102950, 
    102940, 102950, 102920, 102930, 102920, 102900, 102890, 102890, 102870, 
    102840, 102830, 102810, 102780, 102790, 102750, 102720, 102710, 102710, 
    102710, 102690, 102690, 102680, 102680, 102650, 102640, 102610, 102610, 
    102590, 102570, 102570, 102540, 102520, 102520, 102490, 102460, 102430, 
    102410, 102390, 102370, 102340, 102330, 102330, 102320, 102290, 102260, 
    102250, 102210, 102180, 102140, 102100, 102090, 102070, 102040, 102010, 
    101990, 101980, 101950, 101930, 101890, 101860, 101830, 101810, 101800, 
    101800, 101800, 101780, 101780, 101760, 101750, 101760, 101770, 101750, 
    101760, 101750, 101770, 101770, 101760, 101790, 101820, 101820, 101840, 
    101840, 101830, 101820, 101830, 101830, 101840, 101860, 101880, 101890, 
    101900, 101900, 101920, 101920, 101930, 101950, 101940, 101940, 101930, 
    101960, 101950, 101930, 101940, 101930, 101940, 101950, 101950, 101940, 
    101930, 101930, 101910, 101900, 101890, 101900, 101880, 101880, 101860, 
    101850, 101860, 101840, 101830, 101820, 101810, 101810, 101800, 101800, 
    101760, 101750, 101720, 101720, 101700, 101700, 101680, 101660, 101620, 
    101600, 101580, 101530, 101510, 101480, 101450, 101400, 101360, 101300, 
    101230, 101160, 101080, 101010, 100940, 100870, 100740, 100620, 100510, 
    100400, 100300, 100220, 100160, 100030, 100110, 100120, 100190, 100180, 
    100240, 100280, 100320, 100370, 100440, 100500, 100590, 100650, 100710, 
    100780, 100870, 100950, 100980, 101030, 101090, 101130, 101170, 101200, 
    101200, 101210, 101200, 101180, 101170, 101170, 101180, 101120, 101070, 
    101090, 101050, 101020, 100940, 100910, 100890, 100840, 100830, 100780, 
    100730, 100650, 100590, 100480, 100440, 100440, 100430, 100430, 100460, 
    100500, 100550, 100670, 100730, 100810, 100830, 100890, 100910, 100930, 
    100990, 101020, 100970, 101010, 100990, 100940, 100960, 100910, 100850, 
    100740, 100600, 100500, 100410, 100350, 100290, 100230, 100200, 100190, 
    100210, 100220, 100260, 100300, 100340, 100380, 100420, 100440, 100470, 
    100530, 100590, 100660, 100740, 100820, 100880, 100960, 101030, 101120, 
    101200, 101280, 101330, 101360, 101410, 101470, 101510, 101550, 101620, 
    101670, 101680, 101720, 101740, 101760, 101780, 101810, 101810, 101820, 
    101850, 101870, 101870, 101850, 101830, 101800, 101760, 101690, 101630, 
    101580, 101560, 101580, 101640, 101690, 101720, 101780, 101820, 101860, 
    101870, 101900, 101900, 101890, 101900, 101910, 101920, 101930, 101900, 
    101870, 101860, 101840, 101780, 101730, 101680, 101620, 101570, 101560, 
    101530, 101480, 101430, 101370, 101340, 101310, 101280, 101250, 101250, 
    101220, 101220, 101230, 101250, 101260, 101250, 101250, 101230, 101220, 
    101220, 101190, 101160, 101120, 101110, 101090, 101090, 101070, 101060, 
    101040, 101020, 101030, 101050, 101070, 101080, 101140, 101230, 101310, 
    101370, 101440, 101500, 101560, 101610, 101680, 101740, 101780, 101840, 
    101870, 101940, 102010, 102070, 102130, 102160, 102160, 102160, 102220, 
    102260, 102290, 102310, 102300, 102290, 102340, 102370, 102430, 102440, 
    102490, 102520, 102540, 102530, 102560, 102590, 102600, 102640, 102650, 
    102690, 102750, 102780, 102810, 102820, 102830, 102840, 102860, 102880, 
    102900, 102880, 102890, 102890, 102890, 102890, 102880, 102860, 102840, 
    102820, 102780, 102720, 102660, 102610, 102570, 102510, 102480, 102430, 
    102380, 102320, 102270, 102200, 102150, 102080, 102040, 101980, 101920, 
    101860, 101820, 101790, 101750, 101690, 101640, 101570, 101490, 101430, 
    101380, 101320, 101280, 101240, 101200, 101170, 101140, 101090, 101050, 
    101010, 100960, 100900, 100840, 100790, 100750, 100720, 100680, 100650, 
    100610, 100520, 100510, 100510, 100530, 100550, 100580, 100600, 100600, 
    100610, 100630, 100660, 100680, 100730, 100760, 100780, 100830, 100870, 
    100900, 100920, 100950, 100970, 101000, 101010, 101030, 101030, 101050, 
    101040, 101060, 101060, 101090, 101100, 101120, 101120, 101130, 101130, 
    101130, 101130, 101080, 101060, 101020, 100990, 100960, 100910, 100870, 
    100830, 100800, 100770, 100750, 100730, 100700, 100650, 100630, 100640, 
    100660, 100680, 100710, 100700, 100710, 100730, 100750, 100770, 100760, 
    100770, 100760, 100760, 100760, 100750, 100770, 100770, 100780, 100780, 
    100770, 100750, 100720, 100700, 100690, 100680, 100700, 100690, 100690, 
    100690, 100690, 100690, 100690, 100690, 100680, 100660, 100650, 100640, 
    100630, 100650, 100660, 100670, 100670, 100690, 100700, 100710, 100710, 
    100720, 100720, 100740, 100750, 100770, 100790, 100800, 100830, 100850, 
    100860, 100890, 100900, 100910, 100930, 100940, 100970, 100990, 101020, 
    101050, 101070, 101090, 101120, 101150, 101160, 101180, 101200, 101220, 
    101240, 101270, 101310, 101340, 101360, 101370, 101380, 101410, 101420, 
    101430, 101430, 101450, 101460, 101480, 101500, 101520, 101550, 101560, 
    101580, 101580, 101590, 101590, 101610, 101620, 101630, 101660, 101660, 
    101650, 101640, 101630, 101620, 101600, 101590, 101580, 101560, 101540, 
    101510, 101500, 101490, 101480, 101440, 101380, 101340, 101310, 101290, 
    101250, 101230, 101210, 101180, 101170, 101170, 101150, 101120, 101090, 
    101070, 101060, 101050, 101050, 101020, 101020, 101040, 101060, 101070, 
    101090, 101100, 101100, 101120, 101150, 101170, 101180, 101170, 101200, 
    101200, 101200, 101210, 101250, 101260, 101270, 101280, 101300, 101300, 
    101290, 101300, 101320, 101330, 101350, 101380, 101390, 101400, 101420, 
    101450, 101470, 101480, 101460, 101490, 101500, 101510, 101520, 101550, 
    101570, 101590, 101600, 101610, 101630, 101650, 101680, 101700, 101690, 
    101720, 101750, 101760, 101780, 101800, 101810, 101860, 101870, 101900, 
    101920, 101900, 101900, 101900, 101940, 101940, 101960, 101980, 102000, 
    102000, 102020, 102030, 102020, 102030, 102030, 102040, 102050, 102070, 
    102100, 102140, 102150, 102140, 102150, 102150, 102100, 102070, 102030, 
    102000, 102000, 102000, 101990, 101970, 102010, 102000, 102000, 101990, 
    101970, 101960, 101920, 101900, 101890, 101880, 101840, 101810, 101770, 
    101770, 101740, 101700, 101660, 101640, 101610, 101590, 101570, 101490, 
    101430, 101380, 101360, 101330, 101290, 101260, 101200, 101120, 101100, 
    101040, 101010, 100980, 100980, 100930, 100910, 100930, 100930, 100970, 
    100970, 100980, 100980, 100990, 101010, 101010, 101010, 100980, 100940, 
    100920, 100890, 100860, 100780, 100720, 100660, 100610, 100510, 100440, 
    100420, 100340, 100250, 100200, 100110, 100000, 99880, 99800, 99720, 
    99710, 99840, 99910, 99950, 99980, 100010, 100030, 100050, 100060, 
    100040, 100030, 99990, 99950, 99860, 99800, 99730, 99670, 99600, 99430, 
    99280, 99170, 99130, 99110, 98110, 99140, 99230, 99310, 99380, 99460, 
    99540, 99600, 99670, 99740, 99800, 99880, 99950, 100010, 100080, 100130, 
    100220, 100270, 100320, 100350, 100410, 100410, 100420, 100430, 100430, 
    100400, 100380, 100360, 100370, 100390, 100420, 100420, 100400, 100420, 
    100390, 100340, 100290, 100260, 100240, 100230, 100220, 100240, 100240, 
    100250, 100260, 100310, 100320, 100380, 100460, 100520, 100590, 100640, 
    100690, 100750, 100810, 100860, 100900, 100910, 100930, 100900, 100890, 
    100910, 100850, 100780, 100690, 100600, 100510, 100420, 100300, 100180, 
    100030, 99870, 99690, 99540, 99430, 99330, 99290, 99290, 99280, 99320, 
    99400, 99490, 99630, 99740, 99870, 99980, 100110, 100230, 100340, 100450, 
    100550, 100660, 100750, 100850, 100920, 100990, 101080, 101160, 101200, 
    101260, 101300, 101370, 101400, 101420, 101420, 101410, 101400, 101420, 
    101420, 101410, 101390, 101400, 101390, 101350, 101330, 101300, 101250, 
    101170, 101060, 100970, 100820, 100720, 100660, 100600, 100550, 100520, 
    100500, 100520, 100540, 100570, 100600, 100620, 100660, 100720, 100780, 
    100860, 100940, 101030, 101100, 101190, 101250, 101320, 101390, 101440, 
    101520, 101580, 101650, 101710, 101780, 101830, 101870, 101900, 101950, 
    101940, 101910, 101890, 101840, 101790, 101720, 101640, 101600, 101540, 
    101500, 101450, 101420, 101430, 101420, 101380, 101490, 101560, 101680, 
    101790, 101890, 102000, 102030, 102160, 102250, 102340, 102420, 102460, 
    102490, 102520, 102570, 102610, 102670, 102670, 102670, 102680, 102720, 
    102730, 102710, 102670, 102610, 102570, 102520, 102480, 102430, 102390, 
    102330, 102280, 102230, 102170, 102120, 102040, 101950, 101920, 101880, 
    101840, 101800, 101770, 101740, 101700, 101650, 101630, 101580, 101520, 
    101490, 101450, 101430, 101430, 101380, 101400, 101380, 101350, 101290, 
    101260, 101250, 101190, 101120, 101090, 101110, 101120, 101120, 101120, 
    101120, 101100, 101110, 101090, 101070, 101070, 101030, 101000, 100980, 
    100950, 100890, 100840, 100760, 100670, 100580, 100530, 100440, 100370, 
    100280, 100140, 100080, 100040, 100050, 100080, 100100, 100050, 100040, 
    100020, 100030, 100080, 100070, 100070, 100080, 100090, 100100, 100090, 
    100090, 100080, 100100, 100090, 100090, 100090, 100110, 100110, 100130, 
    100150, 100160, 100150, 100160, 100140, 100140, 100140, 100120, 100080, 
    100060, 100040, 100030, 100010, 100010, 99980, 99950, 99930, 99900, 
    99870, 99850, 99810, 99800, 99800, 99810, 99810, 99800, 99800, 99790, 
    99780, 99810, 99810, 99830, 99830, 99860, 99850, 99870, 99890, 99910, 
    99950, 99980, 100000, 100050, 100090, 100120, 100130, 100150, 100160, 
    100200, 100210, 100230, 100210, 100220, 100200, 100180, 100170, 100120, 
    100070, 100010, 99920, 99900, 99880, 99840, 99800, 99790, 99790, 99800, 
    99800, 99840, 99850, 99890, 99910, 99970, 100030, 100080, 100130, 100190, 
    100250, 100290, 100340, 100380, 100430, 100460, 100490, 100540, 100580, 
    100610, 100640, 100670, 100690, 100710, 100710, 100710, 100730, 100730, 
    100730, 100730, 100760, 100760, 100760, 100780, 100800, 100810, 100830, 
    100840, 100860, 100880, 100910, 100940, 100980, 101030, 101060, 101110, 
    101160, 101200, 101240, 101270, 101310, 101310, 101320, 101360, 101380, 
    101410, 101490, 101530, 101550, 101580, 101580, 101570, 101530, 101500, 
    101450, 101400, 101370, 101330, 101280, 101200, 101120, 101040, 100970, 
    100890, 100820, 100770, 100720, 100680, 100630, 100590, 100560, 100530, 
    100510, 100510, 100510, 100510, 100530, 100560, 100580, 100610, 100670, 
    100690, 100710, 100770, 100810, 100880, 100930, 101000, 101020, 101050, 
    101070, 101110, 101100, 101140, 101130, 101110, 101060, 101020, 100950, 
    100870, 100780, 100700, 100630, 100520, 100430, 100390, 100380, 100360, 
    100350, 100360, 100360, 100400, 100440, 100490, 100540, 100620, 100690, 
    100790, 100850, 100920, 100970, 101030, 101090, 101150, 101220, 101280, 
    101340, 101400, 101440, 101440, 101470, 101500, 101540, 101560, 101540, 
    101500, 101460, 101420, 101420, 101440, 101400, 101380, 101400, 101410, 
    101380, 101350, 101280, 101210, 101150, 101070, 100990, 100940, 100870, 
    100820, 100780, 100740, 100720, 100720, 100760, 100770, 100810, 100850, 
    100900, 100930, 100990, 101040, 101100, 101170, 101220, 101240, 101270, 
    101320, 101340, 101360, 101380, 101400, 101400, 101440, 101440, 101440, 
    101440, 101450, 101440, 101450, 101520, 101590, 101620, 101660, 101690, 
    101740, 101780, 101810, 101850, 101880, 101860, 101850, 101850, 101860, 
    101860, 101870, 101890, 101900, 101940, 101960, 102000, 102040, 102060, 
    102090, 102150, 102210, 102250, 102290, 102350, 102390, 102400, 102420, 
    102430, 102430, 102430, 102400, 102370, 102350, 102310, 102270, 102230, 
    102180, 102140, 102090, 102030, 101940, 101870, 101780, 101690, 101570, 
    101480, 101360, 101260, 101180, 101080, 100970, 100870, 100790, 100660, 
    100570, 100500, 100420, 100380, 100350, 100320, 100300, 100300, 100280, 
    100270, 100290, 100310, 100310, 100330, 100350, 100360, 100370, 100390, 
    100410, 100420, 100440, 100470, 100410, 100410, 100390, 100390, 100380, 
    100350, 100350, 100330, 100280, 100260, 100230, 100190, 100170, 100150, 
    100110, 100080, 100070, 100050, 100040, 100030, 100020, 100010, 100020, 
    100010, 100000, 99980, 99980, 99980, 99980, 99980, 99980, 99980, 99950, 
    99930, 99910, 99900, 99890, 99880, 99850, 99840, 99830, 99810, 99840, 
    99840, 99840, 99830, 99840, 99860, 99880, 99910, 99920, 99950, 99980, 
    100010, 100060, 100100, 100140, 100180, 100220, 100290, 100340, 100400, 
    100470, 100550, 100610, 100680, 100750, 100840, 100910, 100980, 101040, 
    101110, 101180, 101210, 101250, 101270, 101290, 101340, 101360, 101370, 
    101420, 101450, 101450, 101450, 101480, 101480, 101480, 101490, 101500, 
    101500, 101500, 101490, 101480, 101480, 101480, 101490, 101500, 101470, 
    101470, 101450, 101430, 101380, 101360, 101360, 101320, 101310, 101270, 
    101250, 101250, 101210, 101160, 101140, 101080, 101050, 101060, 101030, 
    101010, 100980, 100950, 100960, 100920, 100890, 100860, 100830, 100800, 
    100780, 100730, 100710, 100670, 100660, 100620, 100600, 100610, 100580, 
    100520, 100470, 100450, 100400, 100340, 100300, 100230, 100200, 100150, 
    100100, 100020, 99950, 99890, 99850, 99830, 99770, 99760, 99760, 99730, 
    99700, 99700, 99690, 99730, 99760, 99800, 99830, 99860, 99920, 99990, 
    100060, 100120, 100190, 100270, 100330, 100400, 100460, 100490, 100540, 
    100610, 100660, 100710, 100770, 100840, 100890, 100940, 101000, 101040, 
    101080, 101110, 101170, 101180, 101230, 101260, 101300, 101330, 101350, 
    101360, 101370, 101390, 101400, 101400, 101400, 101380, 101390, 101390, 
    101410, 101410, 101410, 101430, 101420, 101420, 101420, 101410, 101420, 
    101420, 101430, 101430, 101430, 101440, 101440, 101440, 101430, 101460, 
    101470, 101490, 101500, 101510, 101520, 101520, 101520, 101520, 101530, 
    101540, 101540, 101540, 101550, 101540, 101520, 101510, 101500, 101500, 
    101480, 101480, 101470, 101450, 101420, 101400, 101370, 101320, 101300, 
    101260, 101240, 101220, 101220, 101170, 101130, 101080, 101020, 101010, 
    100990, 100920, 100850, 100790, 100760, 100730, 100710, 100670, 100610, 
    100600, 100570, 100540, 100480, 100460, 100420, 100370, 100320, 100270, 
    100210, 100160, 100090, 100050, 100020, 99970, 99920, 99870, 99830, 
    99790, 99760, 99730, 99720, 99710, 99720, 99710, 99700, 99710, 99720, 
    99730, 99730, 99750, 99760, 99760, 99770, 99810, 99840, 99860, 99890, 
    99910, 99960, 99980, 100010, 100030, 100050, 100070, 100120, 100160, 
    100200, 100240, 100270, 100320, 100350, 100380, 100420, 100440, 100480, 
    100520, 100560, 100610, 100650, 100700, 100720, 100760, 100790, 100820, 
    100850, 100870, 100870, 100850, 100890, 100900, 100900, 100890, 100840, 
    100770, 100730, 100690, 100560, 100470, 100350, 100300, 100290, 100170, 
    100110, 100020, 99990, 100000, 99990, 100020, 99970, 99930, 99940, 99940, 
    99930, 99920, 99880, 99870, 99860, 99850, 99840, 99810, 99730, 99730, 
    99720, 99710, 99690, 99620, 99570, 99520, 99490, 99460, 99430, 99420, 
    99410, 99390, 99410, 99450, 99530, 99610, 99680, 99770, 99860, 99930, 
    100020, 100090, 100140, 100220, 100240, 100270, 100330, 100380, 100440, 
    100500, 100560, 100640, 100690, 100740, 100810, 100860, 100920, 100950, 
    100990, 101050, 101100, 101120, 101130, 101140, 101150, 101140, 101130, 
    101080, 101090, 101060, 101030, 101000, 100970, 100930, 100870, 100820, 
    100760, 100690, 100590, 100530, 100480, 100440, 100380, 100400, 100320, 
    100230, 100130, 100020, 99940, 99870, 99830, 99730, 99680, 99660, 99620, 
    99590, 99560, 99540, 99520, 99500, 99500, 99510, 99530, 99550, 99590, 
    99640, 99690, 99770, 99830, 99900, 99970, 100050, 100130, 100200, 100250, 
    100300, 100350, 100410, 100440, 100480, 100530, 100570, 100600, 100620, 
    100660, 100690, 100730, 100730, 100740, 100770, 100830, 100850, 100890, 
    100920, 100940, 100970, 101000, 101030, 101040, 101070, 101060, 101080, 
    101090, 101110, 101120, 101120, 101140, 101150, 101150, 101160, 101140, 
    101170, 101170, 101190, 101180, 101180, 101200, 101220, 101230, 101220, 
    101200, 101200, 101200, 101190, 101170, 101160, 101160, 101170, 101170, 
    101160, 101160, 101140, 101140, 101130, 101110, 101100, 101090, 101080, 
    101070, 101110, 101120, 101080, 101070, 101050, 101030, 101000, 100970, 
    100930, 100850, 100820, 100770, 100750, 100700, 100670, 100610, 100570, 
    100540, 100500, 100480, 100410, 100330, 100300, 100250, 100200, 100150, 
    100120, 100090, 100030, 99980, 99920, 99920, 99900, 99850, 99820, 99810, 
    99820, 99830, 99830, 99820, 99820, 99820, 99820, 99830, 99830, 99840, 
    99850, 99860, 99890, 99900, 99900, 99920, 99920, 99890, 99860, 99830, 
    99800, 99770, 99760, 99730, 99700, 99670, 99630, 99580, 99550, 99520, 
    99480, 99440, 99380, 99330, 99300, 99270, 99230, 99190, 99180, 99110, 
    99080, 99080, 99070, 99040, 99020, 99030, 99040, 99050, 99080, 99110, 
    99130, 99140, 99170, 99200, 99210, 99230, 99270, 99300, 99360, 99450, 
    99500, 99570, 99620, 99640, 99680, 99730, 99760, 99790, 99830, 99870, 
    99900, 99950, 100000, 100040, 100070, 100110, 100140, 100160, 100190, 
    100220, 100240, 100250, 100290, 100310, 100350, 100370, 100390, 100390, 
    100410, 100420, 100420, 100420, 100430, 100450, 100450, 100470, 100500, 
    100500, 100500, 100550, 100530, 100520, 100530, 100540, 100540, 100550, 
    100580, 100590, 100630, 100630, 100660, 100690, 100690, 100710, 100720, 
    100720, 100730, 100750, 100760, 100810, 100820, 100860, 100860, 100910, 
    100910, 100970, 101000, 101030, 101060, 101060, 101070, 101080, 101100, 
    101090, 101080, 101080, 101110, 101120, 101100, 101110, 101100, 101120, 
    101150, 101180, 101170, 101190, 101180, 101180, 101170, 101140, 101110, 
    101090, 101050, 101020, 100990, 100960, 100920, 100880, 100810, 100750, 
    100690, 100620, 100560, 100480, 100430, 100390, 100410, 100430, 100480, 
    100580, 100650, 100740, 100800, 100860, 100910, 100960, 101010, 101080, 
    101130, 101190, 101270, 101310, 101370, 101410, 101450, 101480, 101490, 
    101510, 101510, 101530, 101540, 101540, 101570, 101550, 101540, 101540, 
    101560, 101540, 101540, 101520, 101520, 101540, 101540, 101560, 101540, 
    101530, 101570, 101560, 101550, 101540, 101530, 101530, 101540, 101530, 
    101520, 101490, 101500, 101510, 101510, 101510, 101490, 101480, 101490, 
    101460, 101440, 101430, 101430, 101440, 101420, 101430, 101420, 101410, 
    101380, 101390, 101390, 101390, 101380, 101380, 101380, 101380, 101370, 
    101380, 101380, 101370, 101350, 101340, 101330, 101310, 101290, 101310, 
    101320, 101320, 101320, 101330, 101330, 101330, 101340, 101300, 101270, 
    101260, 101260, 101260, 101280, 101290, 101310, 101300, 101310, 101330, 
    101310, 101310, 101330, 101330, 101350, 101350, 101380, 101390, 101390, 
    101400, 101410, 101430, 101430, 101410, 101400, 101370, 101370, 101360, 
    101340, 101340, 101350, 101320, 101310, 101310, 101290, 101260, 101200, 
    101160, 101150, 101140, 101120, 101100, 101090, 101080, 101080, 101100, 
    101110, 101110, 101080, 101050, 101030, 101000, 100960, 100910, 100880, 
    100840, 100790, 100730, 100670, 100640, 100600, 100540, 100470, 100440, 
    100410, 100390, 100360, 100330, 100370, 100390, 100380, 100400, 100390, 
    100400, 100400, 100430, 100490, 100470, 100440, 100430, 100460, 100490, 
    100500, 100530, 100550, 100590, 100620, 100660, 100700, 100740, 100750, 
    100780, 100790, 100790, 100800, 100770, 100770, 100750, 100720, 100670, 
    100650, 100630, 100610, 100560, 100520, 100460, 100410, 100340, 100300, 
    100250, 100200, 100210, 100220, 100260, 100280, 100220, 100180, 100150, 
    100100, 100040, 99990, 99940, 99940, 99910, 99910, 99960, 99940, 100000, 
    100030, 100120, 100160, 100250, 100320, 100390, 100440, 100500, 100560, 
    100630, 100690, 100690, 100700, 100680, 100690, 100700, 100710, 100730, 
    100760, 100790, 100820, 100860, 100890, 100920, 100950, 100940, 100970, 
    100950, 100950, 100920, 100860, 100810, 100750, 100660, 100550, 100490, 
    100410, 100340, 100290, 100240, 100250, 100230, 100240, 100260, 100290, 
    100300, 100340, 100380, 100410, 100430, 100460, 100470, 100500, 100500, 
    100540, 100580, 100640, 100680, 100750, 100800, 100840, 100890, 100920, 
    100940, 100950, 100960, 100950, 100940, 100940, 100940, 100910, 100870, 
    100850, 100810, 100750, 100690, 100590, 100530, 100460, 100390, 100370, 
    100330, 100280, 100260, 100240, 100220, 100220, 100240, 100260, 100300, 
    100330, 100380, 100430, 100490, 100510, 100590, 100620, 100660, 100700, 
    100730, 100740, 100760, 100760, 100780, 100780, 100780, 100780, 100760, 
    100770, 100760, 100740, 100720, 100690, 100650, 100630, 100610, 100580, 
    100590, 100590, 100600, 100550, 100520, 100530, 100490, 100460, 100410, 
    100370, 100370, 100400, 100420, 100460, 100490, 100540, 100600, 100650, 
    100670, 100700, 100770, 100840, 100880, 100920, 100950, 101010, 101030, 
    101070, 101140, 101170, 101190, 101190, 101210, 101230, 101260, 101280, 
    101310, 101310, 101340, 101350, 101350, 101370, 101390, 101420, 101440, 
    101460, 101490, 101530, 101580, 101620, 101670, 101710, 101750, 101790, 
    101810, 101830, 101860, 101840, 101850, 101840, 101840, 101840, 101810, 
    101810, 101800, 101770, 101740, 101720, 101690, 101680, 101680, 101690, 
    101730, 101740, 101730, 101740, 101760, 101780, 101740, 101740, 101720, 
    101690, 101680, 101620, 101580, 101510, 101420, 101350, 101310, 101230, 
    101130, 101050, 100980, 100850, 100780, 100700, 100620, 100570, 100500, 
    100490, 100510, 100500, 100490, 100450, 100390, 100370, 100310, 100280, 
    100250, 100190, 100170, 100160, 100170, 100180, 100200, 100200, 100200, 
    100190, 100180, 100200, 100220, 100250, 100290, 100320, 100360, 100400, 
    100440, 100480, 100510, 100540, 100570, 100620, 100640, 100690, 100740, 
    100790, 100860, 100920, 100960, 100990, 101000, 101050, 101080, 101110, 
    101130, 101150, 101160, 101170, 101150, 101140, 101090, 101070, 101030, 
    101000, 100990, 100950, 100910, 100880, 100860, 100840, 100800, 100740, 
    100690, 100630, 100600, 100570, 100540, 100530, 100530, 100510, 100480, 
    100490, 100470, 100460, 100420, 100410, 100370, 100350, 100340, 100320, 
    100290, 100290, 100310, 100290, 100280, 100250, 100230, 100190, 100180, 
    100160, 100110, 100130, 100090, 100090, 100070, 100030, 100010, 99980, 
    99950, 99920, 99940, 99950, 99960, 99980, 100000, 100030, 100080, 100140, 
    100230, 100280, 100310, 100350, 100380, 100420, 100510, 100560, 100590, 
    100640, 100680, 100740, 100780, 100800, 100810, 100820, 100850, 100850, 
    100850, 100840, 100820, 100790, 100780, 100760, 100710, 100680, 100640, 
    100590, 100570, 100550, 100530, 100500, 100500, 100520, 100550, 100550, 
    100570, 100550, 100540, 100520, 100520, 100560, 100610, 100660, 100750, 
    100870, 100930, 100990, 100990, 101040, 101070, 101090, 101080, 101110, 
    101110, 101150, 101160, 101190, 101210, 101240, 101270, 101270, 101280, 
    101280, 101310, 101290, 101340, 101420, 101490, 101600, 101660, 101680, 
    101740, 101760, 101750, 101790, 101780, 101770, 101730, 101680, 101610, 
    101540, 101480, 101420, 101370, 101350, 101360, 101340, 101340, 101370, 
    101390, 101400, 101450, 101450, 101480, 101530, 101550, 101580, 101590, 
    101630, 101630, 101660, 101660, 101660, 101680, 101690, 101670, 101650, 
    101650, 101640, 101650, 101650, 101660, 101640, 101650, 101680, 101740, 
    101780, 101790, 101820, 101850, 101870, 101860, 101870, 101910, 101910, 
    101970, 102020, 102060, 102070, 102110, 102140, 102170, 102190, 102200, 
    102200, 102220, 102210, 102200, 102200, 102210, 102220, 102220, 102220, 
    102240, 102230, 102230, 102220, 102180, 102160, 102160, 102160, 102160, 
    102160, 102140, 102130, 102110, 102110, 102100, 102070, 102030, 102000, 
    101980, 101980, 101990, 101990, 101960, 101950, 101920, 101880, 101880, 
    101840, 101780, 101800, 101810, 101860, 101870, 101870, 101880, 101860, 
    101860, 101860, 101860, 101860, 101870, 101870, 101830, 101820, 101830, 
    101860, 101870, 101850, 101840, 101850, 101830, 101790, 101740, 101760, 
    101760, 101760, 101770, 101750, 101720, 101710, 101720, 101710, 101700, 
    101720, 101720, 101730, 101750, 101740, 101760, 101760, 101760, 101780, 
    101830, 101850, 101890, 101930, 101950, 101960, 101990, 101990, 102000, 
    101990, 102000, 102000, 101990, 101990, 102000, 101980, 101970, 101950, 
    101920, 101930, 101920, 101920, 101920, 101890, 101880, 101850, 101830, 
    101810, 101780, 101760, 101720, 101690, 101670, 101640, 101640, 101610, 
    101590, 101560, 101540, 101510, 101480, 101450, 101410, 101390, 101390, 
    101380, 101360, 101340, 101330, 101300, 101270, 101260, 101230, 101210, 
    101200, 101200, 101200, 101190, 101200, 101170, 101200, 101190, 101200, 
    101210, 101200, 101210, 101230, 101260, 101280, 101320, 101340, 101350, 
    101350, 101370, 101370, 101380, 101350, 101310, 101340, 101320, 101320, 
    101320, 101320, 101290, 101270, 101250, 101210, 101180, 101110, 101040, 
    101010, 100980, 100970, 100940, 100910, 100880, 100850, 100820, 100800, 
    100750, 100720, 100690, 100630, 100610, 100560, 100510, 100490, 100410, 
    100360, 100320, 100210, 100240, 100210, 100170, 100150, 100100, 100040, 
    99990, 99940, 99910, 99860, 99860, 99840, 99800, 99760, 99740, 99730, 
    99760, 99720, 99790, 99840, 99800, 99840, 99900, 99900, 99910, 99950, 
    99940, 99950, 99970, 100010, 100040, 100060, 100100, 100110, 100130, 
    100150, 100160, 100170, 100200, 100230, 100260, 100270, 100300, 100330, 
    100340, 100340, 100350, 100370, 100360, 100360, 100370, 100380, 100410, 
    100420, 100430, 100430, 100440, 100470, 100480, 100490, 100490, 100510, 
    100520, 100530, 100570, 100590, 100640, 100670, 100690, 100700, 100730, 
    100770, 100770, 100780, 100800, 100830, 100860, 100890, 100920, 100950, 
    100980, 100990, 101010, 101020, 101040, 101060, 101070, 101070, 101090, 
    101120, 101150, 101160, 101180, 101180, 101190, 101200, 101190, 101190, 
    101160, 101170, 101180, 101170, 101190, 101170, 101160, 101150, 101140, 
    101120, 101090, 101080, 101060, 101060, 101050, 101040, 101040, 101030, 
    101000, 101010, 101010, 100990, 100960, 100950, 100940, 100930, 100920, 
    100910, 100930, 100930, 100930, 100930, 100930, 100910, 100900, 100880, 
    100890, 100910, 100910, 100920, 100930, 100910, 100910, 100910, 100910, 
    100900, 100910, 100900, 100880, 100870, 100850, 100860, 100850, 100850, 
    100840, 100840, 100840, 100830, 100830, 100820, 100810, 100800, 100790, 
    100770, 100770, 100760, 100790, 100780, 100800, 100800, 100800, 100790, 
    100780, 100770, 100760, 100760, 100780, 100790, 100810, 100810, 100820, 
    100810, 100810, 100800, 100800, 100790, 100780, 100780, 100790, 100810, 
    100820, 100840, 100830, 100850, 100850, 100850, 100850, 100850, 100860, 
    100870, 100880, 100890, 100910, 100910, 100920, 100930, 100930, 100940, 
    100950, 100970, 100980, 100980, 101000, 101030, 101040, 101060, 101080, 
    101110, 101100, 101110, 101120, 101140, 101150, 101160, 101170, 101180, 
    101190, 101170, 101160, 101150, 101140, 101150, 101110, 101090, 101070, 
    101090, 101070, 101050, 101030, 101020, 100990, 100960, 100920, 100870, 
    100820, 100770, 100720, 100680, 100640, 100620, 100530, 100470, 100430, 
    100380, 100300, 100260, 100180, 100090, 100000, 99920, 99840, 99710, 
    99590, 99540, 99420, 99270, 99150, 98990, 98820, 98680, 98600, 98580, 
    98520, 98500, 98470, 98480, 98470, 98460, 98460, 98430, 98440, 98430, 
    98430, 98460, 98470, 98460, 98480, 98490, 98490, 98480, 98490, 98490, 
    98480, 98490, 98500, 98500, 98510, 98520, 98520, 98550, 98560, 98570, 
    98590, 98590, 98590, 98590, 98610, 98610, 98620, 98630, 98660, 98660, 
    98660, 98670, 98680, 98680, 98670, 98670, 98680, 98710, 98730, 98740, 
    98760, 98770, 98770, 98810, 98840, 98870, 98920, 98950, 98980, 99040, 
    99100, 99150, 99170, 99200, 99260, 99270, 99290, 99300, 99320, 99390, 
    99430, 99480, 99500, 99560, 99600, 99640, 99680, 99700, 99750, 99800, 
    99820, 99850, 99880, 99940, 99970, 99990, 100030, 100050, 100060, 100050, 
    100090, 100120, 100140, 100140, 100150, 100170, 100190, 100220, 100250, 
    100280, 100310, 100320, 100350, 100400, 100470, 100490, 100510, 100550, 
    100580, 100610, 100640, 100680, 100690, 100710, 100730, 100740, 100780, 
    100800, 100830, 100850, 100890, 100920, 100950, 100960, 101000, 101020, 
    101000, 101010, 101040, 101050, 101050, 101050, 101060, 101070, 101090, 
    101100, 101090, 101090, 101090, 101090, 101090, 101100, 101110, 101110, 
    101130, 101130, 101130, 101150, 101150, 101160, 101150, 101160, 101170, 
    101160, 101170, 101180, 101190, 101200, 101200, 101190, 101190, 101160, 
    101120, 101090, 101090, 101070, 101040, 100990, 100940, 100870, 100850, 
    100810, 100760, 100760, 100660, 100630, 100550, 100480, 100430, 100360, 
    100310, 100270, 100220, 100170, 100120, 100060, 100040, 100010, 99980, 
    99960, 99950, 99940, 99950, 99960, 99970, 100000, 100030, 100050, 100090, 
    100140, 100180, 100220, 100260, 100310, 100370, 100400, 100460, 100490, 
    100520, 100530, 100560, 100560, 100580, 100610, 100630, 100640, 100640, 
    100650, 100660, 100670, 100680, 100690, 100700, 100700, 100710, 100730, 
    100730, 100730, 100740, 100750, 100770, 100790, 100820, 100830, 100860, 
    100880, 100910, 100950, 100990, 101030, 101060, 101120, 101160, 101190, 
    101220, 101250, 101280, 101310, 101350, 101380, 101400, 101410, 101410, 
    101410, 101420, 101390, 101370, 101330, 101300, 101260, 101240, 101200, 
    101180, 101170, 101220, 101220, 101220, 101230, 101200, 101180, 101160, 
    101130, 101060, 101000, 100940, 100840, 100810, 100770, 100720, 100650, 
    100570, 100490, 100390, 100280, 100190, 100080, 99980, 99860, 99720, 
    99610, 99440, 99240, 99070, 98920, 98750, 98720, 98920, 99070, 99100, 
    99180, 99150, 99100, 99090, 99090, 99180, 99180, 99150, 99190, 99230, 
    99290, 99400, 99530, 99630, 99750, 99830, 99900, 100050, 100200, 100330, 
    100450, 100520, 100550, 100670, 100720, 100830, 100900, 100980, 101010, 
    101010, 101020, 101030, 101020, 100990, 100990, 100970, 100950, 100950, 
    100970, 101000, 101020, 101010, 100990, 100960, 100950, 100940, 100900, 
    100890, 100850, 100840, 100810, 100770, 100680, 100630, 100550, 100510, 
    100460, 100410, 100380, 100370, 100390, 100390, 100390, 100380, 100360, 
    100350, 100320, 100280, 100260, 100220, 100200, 100180, 100150, 100140, 
    100140, 100140, 100130, 100100, 100030, 99980, 99950, 99920, 99830, 
    99790, 99660, 99540, 99420, 99300, 99200, 99130, 99080, 99080, 99110, 
    99170, 99240, 99320, 99400, 99490, 99600, 99690, 99780, 99890, 99980, 
    100080, 100190, 100300, 100400, 100500, 100610, 100700, 100800, 100900, 
    101000, 101080, 101130, 101210, 101260, 101340, 101420, 101500, 101580, 
    101650, 101700, 101740, 101770, 101820, 101840, 101850, 101880, 101900, 
    101920, 101910, 101900, 101870, 101830, 101770, 101710, 101640, 101560, 
    101480, 101420, 101370, 101320, 101250, 101190, 101110, 101070, 101050, 
    100980, 100990, 101050, 101080, 101130, 101150, 101180, 101200, 101260, 
    101310, 101360, 101410, 101450, 101500, 101540, 101600, 101650, 101710, 
    101770, 101820, 101870, 101910, 101940, 101980, 102010, 102030, 102030, 
    102040, 102040, 101990, 101990, 101970, 101940, 101900, 101840, 101780, 
    101760, 101710, 101680, 101620, 101580, 101570, 101560, 101570, 101560, 
    101570, 101600, 101590, 101600, 101580, 101590, 101570, 101580, 101600, 
    101580, 101570, 101550, 101520, 101510, 101490, 101460, 101440, 101400, 
    101390, 101350, 101330, 101330, 101320, 101310, 101310, 101330, 101330, 
    101320, 101340, 101350, 101340, 101370, 101380, 101410, 101440, 101470, 
    101510, 101550, 101580, 101610, 101630, 101660, 101670, 101680, 101680, 
    101690, 101700, 101690, 101690, 101680, 101700, 101730, 101740, 101710, 
    101690, 101660, 101670, 101660, 101670, 101670, 101650, 101630, 101610, 
    101610, 101620, 101610, 101580, 101560, 101570, 101590, 101590, 101610, 
    101610, 101600, 101570, 101580, 101560, 101550, 101550, 101510, 101480, 
    101480, 101460, 101420, 101420, 101380, 101360, 101320, 101300, 101280, 
    101250, 101210, 101170, 101140, 101100, 101090, 101050, 101010, 100990, 
    100980, 100950, 100920, 100890, 100880, 100850, 100810, 100800, 100800, 
    100840, 100830, 100780, 100780, 100810, 100800, 100820, 100810, 100840, 
    100850, 100840, 100850, 100860, 100860, 100850, 100850, 100830, 100800, 
    100770, 100730, 100710, 100700, 100700, 100680, 100670, 100660, 100650, 
    100640, 100620, 100600, 100560, 100540, 100500, 100470, 100450, 100440, 
    100430, 100410, 100410, 100390, 100370, 100370, 100380, 100360, 100380, 
    100430, 100460, 100490, 100530, 100540, 100570, 100600, 100610, 100620, 
    100620, 100630, 100630, 100650, 100680, 100700, 100700, 100720, 100710, 
    100690, 100690, 100710, 100720, 100730, 100720, 100740, 100780, 100830, 
    100880, 100920, 100930, 100940, 100980, 101000, 101020, 101060, 101090, 
    101130, 101170, 101200, 101240, 101270, 101290, 101310, 101330, 101340, 
    101370, 101410, 101420, 101440, 101460, 101490, 101500, 101520, 101540, 
    101550, 101560, 101560, 101560, 101590, 101600, 101620, 101620, 101630, 
    101640, 101630, 101610, 101600, 101600, 101590, 101580, 101580, 101590, 
    101550, 101540, 101530, 101500, 101470, 101430, 101370, 101370, 101340, 
    101310, 101310, 101290, 101290, 101290, 101270, 101260, 101230, 101220, 
    101220, 101220, 101220, 101220, 101220, 101240, 101240, 101240, 101250, 
    101270, 101260, 101270, 101280, 101280, 101300, 101310, 101340, 101360, 
    101390, 101400, 101420, 101430, 101430, 101430, 101460, 101470, 101480, 
    101510, 101510, 101500, 101500, 101490, 101480, 101490, 101480, 101470, 
    101450, 101460, 101460, 101460, 101460, 101440, 101420, 101410, 101360, 
    101320, 101310, 101280, 101280, 101230, 101210, 101190, 101170, 101120, 
    101100, 101100, 101060, 101040, 101040, 101010, 100990, 100960, 100940, 
    100940, 100920, 100890, 100830, 100810, 100830, 100810, 100780, 100770, 
    100730, 100690, 100660, 100630, 100620, 100650, 100640, 100630, 100640, 
    100640, 100590, 100560, 100560, 100560, 100570, 100560, 100550, 100530, 
    100530, 100520, 100520, 100530, 100550, 100570, 100580, 100570, 100580, 
    100560, 100520, 100510, 100480, 100450, 100470, 100490, 100470, 100430, 
    100410, 100400, 100400, 100390, 100410, 100350, 100340, 100280, 100280, 
    100230, 100170, 100100, 100050, 99980, 99880, 99820, 99750, 99630, 99500, 
    99360, 99260, 99130, 99100, 99030, 98900, 98790, 98750, 98650, 98560, 
    98400, 98260, 98130, 98090, 98020, 97920, 97890, 97900, 97870, 97830, 
    97830, 97790, 97760, 97720, 97730, 97730, 97750, 97740, 97720, 97720, 
    97720, 97710, 97690, 97680, 97670, 97680, 97690, 97710, 97730, 97730, 
    97750, 97770, 97790, 97790, 97810, 97830, 97870, 97890, 97920, 97950, 
    97990, 98040, 98090, 98120, 98170, 98200, 98240, 98260, 98270, 98280, 
    98300, 98330, 98370, 98400, 98410, 98400, 98420, 98420, 98430, 98430, 
    98430, 98460, 98480, 98510, 98540, 98590, 98640, 98670, 98690, 98720, 
    98760, 98800, 98820, 98860, 98880, 98930, 98960, 98970, 99000, 99020, 
    99030, 99040, 99050, 99050, 99060, 99080, 99100, 99130, 99160, 99200, 
    99230, 99240, 99260, 99270, 99290, 99330, 99350, 99380, 99400, 99440, 
    99450, 99450, 99460, 99470, 99480, 99490, 99510, 99490, 99520, 99510, 
    99510, 99520, 99520, 99530, 99530, 99550, 99550, 99550, 99550, 99550, 
    99550, 99550, 99540, 99550, 99570, 99570, 99580, 99580, 99580, 99610, 
    99640, 99690, 99730, 99760, 99790, 99830, 99860, 99910, 99940, 99960, 
    99970, 100010, 100020, 100050, 100050, 100090, 100120, 100160, 100190, 
    100240, 100250, 100260, 100270, 100310, 100330, 100330, 100370, 100420, 
    100450, 100480, 100520, 100570, 100630, 100670, 100720, 100760, 100810, 
    100840, 100880, 100920, 100950, 100980, 100980, 101010, 101030, 101020, 
    101010, 100980, 100970, 100950, 100910, 100880, 100870, 100850, 100830, 
    100810, 100790, 100760, 100740, 100690, 100640, 100590, 100550, 100530, 
    100510, 100490, 100480, 100460, 100460, 100440, 100430, 100420, 100420, 
    100420, 100420, 100420, 100430, 100430, 100420, 100410, 100410, 100420, 
    100420, 100430, 100440, 100450, 100460, 100480, 100480, 100480, 100540, 
    100570, 100600, 100580, 100600, 100650, 100660, 100650, 100650, 100680, 
    100680, 100680, 100700, 100730, 100760, 100760, 100760, 100760, 100750, 
    100750, 100740, 100730, 100700, 100700, 100670, 100660, 100610, 100590, 
    100570, 100530, 100510, 100490, 100460, 100430, 100410, 100410, 100420, 
    100420, 100410, 100410, 100400, 100400, 100380, 100360, 100330, 100290, 
    100270, 100230, 100170, 100140, 100090, 100030, 100000, 99920, 99830, 
    99720, 99640, 99570, 99510, 99460, 99400, 99320, 99260, 99170, 99100, 
    99020, 98950, 98880, 98800, 98740, 98690, 98630, 98580, 98550, 98500, 
    98500, 98500, 98480, 98480, 98480, 98470, 98490, 98540, 98590, 98650, 
    98690, 98760, 98810, 98850, 98890, 98900, 98920, 98950, 98960, 99000, 
    99030, 99070, 99100, 99100, 99120, 99140, 99160, 99190, 99220, 99230, 
    99240, 99250, 99320, 99360, 99380, 99400, 99430, 99460, 99440, 99410, 
    99410, 99410, 99400, 99390, 99370, 99350, 99350, 99310, 99270, 99230, 
    99190, 99140, 99100, 99080, 99050, 99020, 99010, 98990, 99000, 98980, 
    98970, 98950, 98930, 98900, 98900, 98890, 98880, 98890, 98880, 98880, 
    98870, 98870, 98860, 98850, 98830, 98820, 98800, 98780, 98770, 98780, 
    98790, 98820, 98830, 98840, 98840, 98850, 98870, 98880, 98900, 98920, 
    98950, 98980, 99020, 99060, 99100, 99150, 99180, 99230, 99280, 99330, 
    99380, 99440, 99510, 99550, 99650, 99730, 99790, 99870, 99950, 100010, 
    100090, 100150, 100190, 100270, 100350, 100420, 100500, 100570, 100630, 
    100690, 100700, 100750, 100790, 100800, 100820, 100870, 100910, 100980, 
    101050, 101130, 101200, 101240, 101290, 101340, 101410, 101460, 101500, 
    101530, 101570, 101610, 101640, 101660, 101700, 101710, 101700, 101670, 
    101630, 101630, 101630, 101650, 101650, 101670, 101700, 101720, 101750, 
    101760, 101780, 101770, 101770, 101770, 101770, 101760, 101740, 101700, 
    101670, 101630, 101570, 101530, 101480, 101420, 101420, 101350, 101310, 
    101230, 101160, 101120, 101060, 100960, 100850, 100790, 100730, 100620, 
    100510, 100400, 100270, 100120, 100030, 99900, 99800, 99700, 99490, 
    99390, 99210, 99150, 99080, 99050, 98970, 98910, 98820, 98770, 98690, 
    98640, 98560, 98530, 98550, 98610, 98660, 98730, 98880, 98940, 98990, 
    99010, 99050, 99110, 99100, 99110, 99090, 99100, 99090, 99060, 99020, 
    99010, 99010, 99020, 99020, 99020, 99050, 99060, 99090, 99110, 99110, 
    99110, 99130, 99140, 99140, 99150, 99160, 99160, 99160, 99160, 99150, 
    99160, 99150, 99180, 99200, 99210, 99230, 99270, 99320, 99400, 99450, 
    99510, 99550, 99580, 99660, 99720, 99780, 99850, 99900, 99960, 100020, 
    100060, 100110, 100160, 100190, 100220, 100250, 100270, 100280, 100300, 
    100300, 100320, 100330, 100350, 100350, 100350, 100330, 100330, 100300, 
    100260, 100250, 100210, 100170, 100140, 100110, 100080, 100050, 100030, 
    100000, 99970, 99920, 99890, 99860, 99820, 99800, 99800, 99820, 99830, 
    99820, 99830, 99840, 99840, 99860, 99880, 99900, 99940, 99970, 99990, 
    100020, 100060, 100130, 100190, 100230, 100280, 100330, 100400, 100450, 
    100490, 100550, 100610, 100680, 100750, 100820, 100880, 100940, 101020, 
    101040, 101080, 101080, 101120, 101150, 101150, 101160, 101190, 101190, 
    101160, 101140, 101120, 101090, 101050, 101000, 100950, 100930, 100910, 
    100830, 100810, 100770, 100730, 100650, 100560, 100450, 100350, 100250, 
    100170, 100060, 99970, 99850, 99750, 99670, 99590, 99480, 99410, 99310, 
    99180, 99080, 99080, 99000, 98940, 98880, 98840, 98780, 98720, 98660, 
    98650, 98600, 98520, 98480, 98400, 98340, 98300, 98260, 98200, 98160, 
    98130, 98130, 98080, 98080, 98070, 98060, 98050, 98050, 98110, 98120, 
    98150, 98180, 98240, 98290, 98300, 98320, 98350, 98400, 98430, 98480, 
    98520, 98570, 98670, 98710, 98760, 98850, 98950, 99050, 99110, 99230, 
    99340, 99430, 99530, 99640, 99800, 99930, 100070, 100120, 100200, 100260, 
    100380, 100430, 100510, 100550, 100640, 100670, 100760, 100800, 100870, 
    100870, 100940, 100980, 101020, 101070, 101090, 101130, 101200, 101220, 
    101240, 101270, 101300, 101330, 101370, 101390, 101420, 101450, 101440, 
    101460, 101530, 101530, 101580, 101590, 101610, 101630, 101640, 101680, 
    101700, 101710, 101770, 101790, 101850, 101840, 101890, 101950, 102000, 
    102050, 102090, 102120, 102140, 102170, 102190, 102230, 102260, 102280, 
    102320, 102360, 102400, 102420, 102450, 102500, 102540, 102580, 102630, 
    102690, 102760, 102820, 102880, 102910, 102950, 102980, 103000, 103060, 
    103100, 103090, 103130, 103150, 103170, 103160, 103140, 103130, 103110, 
    103080, 103040, 103030, 103000, 102950, 102920, 102830, 102850, 102830, 
    102810, 102750, 102690, 102670, 102610, 102580, 102550, 102500, 102440, 
    102370, 102330, 102280, 102210, 102170, 102110, 102050, 101970, 101900, 
    101850, 101790, 101710, 101650, 101610, 101550, 101490, 101430, 101310, 
    101240, 101160, 101070, 101000, 100910, 100790, 100700, 100630, 100560, 
    100500, 100420, 100310, 100220, 100140, 100070, 100020, 99990, 99950, 
    99950, 99980, 100050, 100140, 100210, 100260, 100320, 100360, 100390, 
    100370, 100370, 100400, 100510, 100610, 100740, 100870, 100970, 101030, 
    101170, 101300, 101350, 101470, 101570, 101700, 101840, 101930, 102030, 
    102120, 102110, 102110, 102150, 102140, 102080, 102050, 102000, 101960, 
    101910, 101880, 101830, 101790, 101780, 101750, 101680, 101640, 101580, 
    101500, 101430, 101370, 101310, 101280, 101240, 101230, 101200, 101150, 
    101120, 101110, 101080, 101060, 101060, 101070, 101080, 101070, 101070, 
    101070, 101070, 101100, 101090, 101090, 101120, 101110, 101130, 101140, 
    101150, 101200, 101270, 101290, 101350, 101390, 101430, 101460, 101510, 
    101540, 101560, 101580, 101610, 101640, 101660, 101680, 101720, 101770, 
    101760, 101780, 101810, 101830, 101870, 101900, 101920, 101950, 102000, 
    102050, 102060, 102080, 102100, 102110, 102120, 102120, 102110, 102120, 
    102150, 102130, 102110, 102090, 102070, 102050, 101980, 101940, 101910, 
    101830, 101790, 101760, 101720, 101680, 101650, 101640, 101620, 101600, 
    101600, 101550, 101520, 101450, 101420, 101420, 101420, 101390, 101380, 
    101350, 101310, 101270, 101220, 101140, 101080, 101000, 100930, 100830, 
    100730, 100680, 100670, 100640, 100570, 100570, 100540, 100510, 100440, 
    100370, 100340, 100280, 100200, 100140, 100110, 100080, 100020, 100000, 
    99940, 99900, 99850, 99820, 99820, 99820, 99870, 99910, 99950, 99960, 
    100020, 100050, 100090, 100140, 100230, 100230, 100260, 100340, 100390, 
    100470, 100490, 100550, 100610, 100660, 100660, 100680, 100730, 100750, 
    100770, 100810, 100820, 100860, 100960, 101020, 101080, 101120, 101160, 
    101220, 101250, 101320, 101390, 101450, 101550, 101610, 101680, 101740, 
    101820, 101860, 101950, 101990, 102040, 102070, 102070, 102080, 102100, 
    102130, 102150, 102200, 102290, 102360, 102420, 102470, 102500, 102530, 
    102540, 102560, 102590, 102640, 102650, 102670, 102680, 102710, 102720, 
    102740, 102750, 102770, 102800, 102800, 102810, 102850, 102890, 102910, 
    102920, 102950, 102960, 102950, 102960, 102980, 102920, 102890, 102890, 
    102870, 102850, 102850, 102850, 102800, 102810, 102780, 102750, 102730, 
    102690, 102620, 102570, 102540, 102530, 102490, 102440, 102400, 102360, 
    102320, 102250, 102190, 102160, 102080, 102040, 101970, 101930, 101880, 
    101810, 101720, 101650, 101580, 101510, 101400, 101320, 101280, 101230, 
    101180, 101120, 101090, 101020, 100970, 100900, 100830, 100780, 100750, 
    100670, 100590, 100520, 100500, 100500, 100490, 100450, 100430, 100460, 
    100450, 100450, 100490, 100520, 100530, 100510, 100560, 100530, 100540, 
    100540, 100580, 100600, 100620, 100620, 100630, 100640, 100680, 100700, 
    100700, 100710, 100740, 100740, 100730, 100760, 100760, 100770, 100780, 
    100760, 100740, 100740, 100750, 100720, 100710, 100700, 100710, 100700, 
    100720, 100710, 100760, 100780, 100790, 100820, 100860, 100890, 100910, 
    100990, 101010, 101030, 101040, 101060, 101070, 101100, 101130, 101140, 
    101170, 101200, 101230, 101260, 101260, 101270, 101310, 101320, 101350, 
    101350, 101370, 101380, 101380, 101380, 101400, 101420, 101420, 101420, 
    101430, 101430, 101420, 101400, 101370, 101340, 101320, 101300, 101250, 
    101230, 101170, 101140, 101100, 101050, 101010, 100960, 100930, 100870, 
    100840, 100800, 100750, 100690, 100620, 100560, 100520, 100470, 100420, 
    100410, 100400, 100390, 100430, 100420, 100470, 100510, 100540, 100560, 
    100620, 100660, 100690, 100730, 100760, 100800, 100870, 100920, 100990, 
    101030, 101120, 101210, 101230, 101290, 101330, 101390, 101440, 101500, 
    101520, 101530, 101570, 101550, 101560, 101560, 101570, 101570, 101560, 
    101550, 101580, 101610, 101660, 101720, 101780, 101870, 101950, 102050, 
    102180, 102260, 102350, 102460, 102490, 102540, 102610, 102720, 102810, 
    102910, 102940, 103020, 103160, 103130, 103170, 103130, 103090, 102990, 
    102910, 102800, 102620, 102480, 102340, 102210, 102090, 101970, 101810, 
    101650, 101500, 101310, 101220, 101170, 101150, 101170, 101150, 101100, 
    101100, 101060, 100980, 100900, 100840, 100720, 100620, 100450, 100300, 
    100120, 99950, 99900, 99790, 99700, 99580, 99500, 99510, 99490, 99630, 
    99700, 99780, 99790, 99810, 99830, 99870, 99900, 100040, 100210, 100390, 
    100570, 100800, 101110, 101390, 101690, 101790, 102070, 102200, 102340, 
    102410, 102530, 102580, 102690, 102740, 102800, 102880, 102950, 102970, 
    102990, 102970, 102920, 102850, 102740, 102710, 102610, 102500, 102390, 
    102240, 102120, 101990, 101830, 101810, 101780, 101760, 101760, 101740, 
    101740, 101820, 101860, 101920, 101980, 102020, 102050, 102090, 102110, 
    102120, 102160, 102190, 102190, 102180, 102210, 102200, 102160, 102120, 
    102090, 102020, 101980, 101940, 101880, 101770, 101660, 101570, 101460, 
    101340, 101270, 101140, 101010, 100890, 100780, 100620, 100460, 100330, 
    100190, 100090, 99980, 99850, 99730, 99630, 99530, 99460, 99420, 99390, 
    99420, 99460, 99550, 99660, 99770, 99860, 99990, 100070, 100160, 100230, 
    100330, 100450, 100530, 100600, 100630, 100710, 100780, 100850, 100910, 
    100930, 100990, 101030, 101060, 101070, 101110, 101080, 101100, 101120, 
    101120, 101160, 101190, 101240, 101260, 101300, 101310, 101310, 101300, 
    101330, 101360, 101410, 101420, 101460, 101460, 101470, 101480, 101490, 
    101510, 101520, 101530, 101540, 101560, 101580, 101630, 101640, 101670, 
    101680, 101680, 101690, 101700, 101700, 101710, 101690, 101710, 101720, 
    101740, 101750, 101770, 101750, 101760, 101770, 101790, 101800, 101760, 
    101770, 101780, 101770, 101800, 101810, 101810, 101810, 101800, 101780, 
    101750, 101710, 101660, 101620, 101570, 101530, 101470, 101420, 101340, 
    101250, 101140, 101050, 100980, 100880, 100750, 100620, 100490, 100400, 
    100260, 100190, 100060, 100000, 100030, 100000, 99970, 99980, 99930, 
    99840, 99830, 99810, 99790, 99750, 99710, 99690, 99650, 99620, 99590, 
    99570, 99590, 99620, 99660, 99660, 99700, 99710, 99740, 99750, 99700, 
    99650, 99610, 99450, 99260, 99400, 99650, 99750, 99740, 99810, 99950, 
    99990, 99980, 99930, 99910, 99890, 99970, 99980, 100020, 100090, 100190, 
    100250, 100260, 100240, 100200, 100270, 100210, 100220, 100270, 100250, 
    100290, 100220, 100240, 100240, 100250, 100250, 100240, 100250, 100240, 
    100260, 100290, 100300, 100340, 100340, 100350, 100390, 100360, 100390, 
    100390, 100370, 100330, 100340, 100360, 100420, 100410, 100410, 100440, 
    100440, 100430, 100450, 100460, 100450, 100480, 100470, 100460, 100400, 
    100410, 100400, 100410, 100390, 100390, 100380, 100350, 100320, 100310, 
    100280, 100290, 100250, 100220, 100200, 100200, 100140, 100130, 100080, 
    100010, 99970, 99910, 99860, 99790, 99750, 99700, 99670, 99660, 99690, 
    99690, 99700, 99690, 99670, 99670, 99670, 99660, 99620, 99610, 99620, 
    99640, 99630, 99620, 99650, 99630, 99610, 99550, 99550, 99550, 99510, 
    99490, 99460, 99470, 99470, 99480, 99440, 99410, 99390, 99350, 99330, 
    99290, 99270, 99270, 99290, 99250, 99230, 99240, 99220, 99220, 99190, 
    99190, 99180, 99150, 99170, 99170, 99180, 99190, 99200, 99210, 99220, 
    99210, 99250, 99270, 99290, 99290, 99290, 99260, 99310, 99310, 99300, 
    99280, 99260, 99230, 99210, 99210, 99200, 99170, 99140, 99130, 99110, 
    99110, 99120, 99120, 99110, 99070, 99060, 99070, 99060, 99090, 99100, 
    99100, 99100, 99130, 99170, 99210, 99230, 99250, 99270, 99300, 99330, 
    99340, 99360, 99380, 99410, 99420, 99470, 99490, 99510, 99510, 99520, 
    99530, 99530, 99540, 99520, 99490, 99470, 99490, 99490, 99440, 99370, 
    99340, 99300, 99280, 99290, 99230, 99210, 99180, 99170, 99150, 99140, 
    99120, 99080, 99090, 99100, 99100, 99090, 99080, 99100, 99100, 99110, 
    99110, 99140, 99160, 99150, 99160, 99190, 99190, 99220, 99230, 99250, 
    99270, 99300, 99340, 99350, 99380, 99400, 99410, 99400, 99410, 99420, 
    99440, 99450, 99450, 99460, 99500, 99570, 99570, 99610, 99640, 99660, 
    99700, 99730, 99780, 99820, 99880, 99930, 100000, 100070, 100130, 100170, 
    100190, 100210, 100280, 100340, 100380, 100400, 100420, 100430, 100480, 
    100520, 100570, 100590, 100630, 100680, 100720, 100750, 100810, 100830, 
    100870, 100900, 100960, 101000, 100990, 100950, 100910, 100850, 100830, 
    100810, 100840, 100890, 100890, 100890, 100910, 100920, 100930, 100930, 
    100870, 100790, 100720, 100630, 100560, 100480, 100420, 100310, 100230, 
    100120, 100020, 99910, 99900, 99900, 99940, 100050, 100170, 100260, 
    100310, 100360, 100450, 100540, 100600, 100620, 100680, 100720, 100700, 
    100740, 100700, 100690, 100680, 100680, 100670, 100640, 100610, 100550, 
    100510, 100470, 100390, 100320, 100230, 100170, 100040, 99960, 99820, 
    99650, 99440, 99160, 98920, 98760, 98680, 98680, 98660, 98650, 98690, 
    98780, 98890, 98960, 99040, 99080, 99080, 99100, 99090, 99050, 99000, 
    98950, 99000, 99070, 99140, 99250, 99310, 99380, 99480, 99600, 99740, 
    99910, 100010, 100080, 100170, 100260, 100310, 100380, 100400, 100440, 
    100430, 100410, 100400, 100350, 100310, 100220, 100150, 100070, 99950, 
    99840, 99740, 99640, 99580, 99490, 99440, 99400, 99380, 99370, 99380, 
    99420, 99400, 99420, 99440, 99430, 99450, 99440, 99440, 99440, 99430, 
    99420, 99380, 99340, 99360, 99440, 99550, 99710, 99890, 99940, 100020, 
    100150, 100230, 100350, 100420, 100540, 100630, 100690, 100770, 100800, 
    100850, 100860, 100870, 100880, 100880, 100870, 100880, 100920, 101000, 
    101030, 101040, 101090, 101150, 101190, 101210, 101270, 101340, 101430, 
    101480, 101570, 101630, 101730, 101810, 101900, 101960, 102040, 102090, 
    102110, 102160, 102280, 102340, 102390, 102440, 102470, 102510, 102550, 
    102560, 102580, 102580, 102580, 102560, 102540, 102530, 102500, 102460, 
    102450, 102410, 102330, 102220, 102090, 102020, 102000, 101940, 101880, 
    101840, 101820, 101830, 101780, 101710, 101660, 101610, 101510, 101460, 
    101430, 101420, 101390, 101410, 101400, 101380, 101370, 101360, 101330, 
    101330, 101310, 101340, 101390, 101420, 101450, 101460, 101450, 101500, 
    101520, 101550, 101560, 101580, 101580, 101560, 101540, 101510, 101490, 
    101490, 101500, 101480, 101450, 101410, 101370, 101360, 101310, 101290, 
    101250, 101250, 101240, 101210, 101210, 101190, 101170, 101150, 101110, 
    101060, 101020, 101010, 100990, 100950, 100900, 100880, 100840, 100820, 
    100790, 100780, 100730, 100710, 100670, 100620, 100580, 100510, 100450, 
    100370, 100310, 100250, 100180, 100100, 100020, 99940, 99850, 99750, 
    99620, 99430, 99280, 99150, 99010, 98900, 98830, 98710, 98600, 98520, 
    98470, 98390, 98340, 98350, 98310, 98360, 98450, 98550, 98700, 98810, 
    98920, 99020, 99150, 99250, 99340, 99410, 99500, 99600, 99670, 99750, 
    99870, 99930, 100000, 100020, 100040, 100080, 100150, 100200, 100270, 
    100340, 100360, 100420, 100440, 100500, 100520, 100550, 100550, 100520, 
    100520, 100490, 100410, 100330, 100290, 100260, 100210, 100130, 100040, 
    100000, 99940, 99880, 99850, 99820, 99790, 99770, 99770, 99750, 99750, 
    99750, 99750, 99770, 99790, 99800, 99830, 99870, 99890, 99890, 99940, 
    99970, 100000, 100040, 100050, 100060, 100100, 100070, 100060, 100040, 
    100070, 100050, 100040, 100030, 100020, 100020, 100010, 100000, 100000, 
    100020, 100020, 100020, 100030, 100050, 100090, 100130, 100140, 100150, 
    100140, 100200, 100220, 100240, 100240, 100250, 100260, 100260, 100270, 
    100310, 100360, 100380, 100380, 100410, 100410, 100460, 100460, 100480, 
    100490, 100500, 100530, 100540, 100580, 100590, 100610, 100620, 100640, 
    100630, 100660, 100660, 100670, 100670, 100670, 100640, 100590, 100540, 
    100530, 100430, 100410, 100360, 100340, 100320, 100310, 100310, 100330, 
    100340, 100410, 100430, 100430, 100400, 100340, 100260, 100180, 100110, 
    100000, 99900, 99820, 99780, 99690, 99600, 99500, 99420, 99350, 99340, 
    99350, 99350, 99390, 99440, 99520, 99600, 99660, 99740, 99800, 99840, 
    99870, 99920, 99960, 99990, 99990, 99990, 100040, 100120, 100190, 100260, 
    100330, 100400, 100470, 100550, 100600, 100660, 100660, 100680, 100690, 
    100710, 100730, 100740, 100750, 100740, 100730, 100720, 100710, 100710, 
    100700, 100690, 100690, 100730, 100760, 100790, 100810, 100840, 100860, 
    100870, 100870, 100840, 100820, 100820, 100830, 100840, 100820, 100810, 
    100770, 100760, 100730, 100700, 100650, 100560, 100510, 100450, 100420, 
    100370, 100360, 100380, 100400, 100440, 100470, 100520, 100550, 100590, 
    100630, 100690, 100740, 100810, 100880, 100940, 100990, 101030, 101080, 
    101110, 101170, 101210, 101270, 101310, 101350, 101390, 101450, 101520, 
    101570, 101600, 101660, 101710, 101730, 101720, 101780, 101770, 101790, 
    101830, 101830, 101830, 101820, 101790, 101770, 101760, 101700, 101630, 
    101580, 101510, 101410, 101280, 101160, 101030, 100920, 100830, 100740, 
    100660, 100580, 100520, 100470, 100420, 100360, 100370, 100350, 100370, 
    100390, 100400, 100420, 100490, 100530, 100560, 100630, 100670, 100700, 
    100740, 100750, 100760, 100800, 100850, 100860, 100880, 100900, 100880, 
    100890, 100910, 100920, 100970, 101000, 100980, 100990, 100970, 100970, 
    100960, 100930, 100880, 100830, 100800, 100780, 100750, 100720, 100700, 
    100690, 100710, 100700, 100690, 100670, 100680, 100700, 100650, 100610, 
    100590, 100530, 100520, 100520, 100480, 100380, 100280, 100290, 100260, 
    100180, 100100, 100040, 100010, 99980, 100000, 99940, 99920, 99870, 
    99860, 99870, 99850, 99840, 99800, 99790, 99760, 99760, 99760, 99710, 
    99680, 99700, 99760, 99710, 99720, 99730, 99750, 99740, 99730, 99730, 
    99750, 99800, 99830, 99850, 99840, 99820, 99850, 99890, 99970, 100050, 
    100080, 100090, 100100, 100090, 100080, 100110, 100170, 100150, 100150, 
    100240, 100320, 100400, 100510, 100590, 100660, 100760, 100840, 100920, 
    100970, 101040, 101050, 101080, 101110, 101170, 101240, 101280, 101290, 
    101300, 101320, 101320, 101320, 101310, 101270, 101250, 101210, 101130, 
    101090, 101030, 100950, 100880, 100810, 100760, 100670, 100580, 100500, 
    100410, 100310, 100230, 100200, 100170, 100180, 100140, 100100, 100100, 
    100100, 100080, 100050, 99960, 99900, 99860, 99780, 99750, 99620, 99480, 
    99350, 99240, 99060, 98880, 98720, 98530, 98490, 98380, 98310, 98230, 
    98210, 98160, 98070, 98070, 98140, 98280, 98380, 98500, 98640, 98750, 
    98900, 99020, 99060, 99270, 99340, 99530, 99680, 99810, 99770, 99890, 
    99980, 100030, 100060, 100050, 100120, 100120, 100130, 100140, 100160, 
    100210, 100220, 100200, 100220, 100250, 100260, 100300, 100300, 100290, 
    100280, 100280, 100270, 100220, 100180, 100170, 100180, 100180, 100140, 
    100120, 100100, 100070, 100040, 100020, 100000, 99960, 99930, 99880, 
    99840, 99800, 99760, 99720, 99690, 99650, 99600, 99570, 99550, 99500, 
    99490, 99460, 99420, 99370, 99330, 99300, 99290, 99280, 99270, 99300, 
    99320, 99370, 99390, 99420, 99410, 99420, 99470, 99520, 99570, 99600, 
    99610, 99650, 99690, 99730, 99750, 99770, 99790, 99820, 99890, 99920, 
    99960, 99990, 100010, 100050, 100090, 100110, 100130, 100160, 100170, 
    100190, 100220, 100250, 100290, 100280, 100280, 100260, 100250, 100250, 
    100280, 100270, 100260, 100270, 100280, 100280, 100290, 100300, 100300, 
    100300, 100300, 100320, 100320, 100310, 100310, 100290, 100290, 100290, 
    100300, 100300, 100300, 100290, 100270, 100280, 100290, 100260, 100260, 
    100270, 100260, 100260, 100280, 100270, 100240, 100240, 100220, 100200, 
    100190, 100190, 100180, 100190, 100190, 100190, 100200, 100200, 100180, 
    100170, 100170, 100180, 100180, 100190, 100200, 100190, 100210, 100230, 
    100240, 100230, 100200, 100190, 100180, 100180, 100180, 100210, 100200, 
    100180, 100170, 100170, 100170, 100150, 100130, 100090, 100070, 100060, 
    100040, 100020, 100000, 99970, 99980, 99990, 100000, 100000, 100000, 
    99990, 99990, 99970, 99970, 99960, 99960, 99960, 99960, 99960, 99990, 
    100030, 100040, 100060, 100040, 100050, 100050, 100080, 100120, 100160, 
    100190, 100240, 100250, 100270, 100330, 100360, 100400, 100440, 100470, 
    100520, 100550, 100590, 100640, 100690, 100730, 100790, 100830, 100870, 
    100900, 100950, 100980, 101020, 101060, 101090, 101150, 101200, 101260, 
    101290, 101310, 101330, 101360, 101390, 101420, 101440, 101470, 101490, 
    101500, 101540, 101580, 101600, 101630, 101650, 101660, 101690, 101700, 
    101700, 101720, 101750, 101780, 101830, 101860, 101880, 101910, 101910, 
    101920, 101930, 101960, 101970, 102000, 102010, 102000, 102010, 102050, 
    102070, 102070, 102080, 102100, 102120, 102130, 102140, 102160, 102200, 
    102250, 102270, 102310, 102330, 102350, 102370, 102400, 102410, 102440, 
    102450, 102480, 102520, 102540, 102570, 102620, 102640, 102650, 102650, 
    102690, 102710, 102720, 102720, 102740, 102780, 102800, 102820, 102820, 
    102850, 102860, 102850, 102860, 102890, 102890, 102890, 102900, 102910, 
    102930, 102930, 102950, 102950, 102940, 102940, 102930, 102910, 102910, 
    102890, 102870, 102880, 102880, 102860, 102820, 102810, 102780, 102760, 
    102760, 102720, 102740, 102720, 102710, 102670, 102650, 102640, 102620, 
    102590, 102550, 102540, 102530, 102520, 102490, 102460, 102440, 102460, 
    102460, 102460, 102460, 102450, 102440, 102410, 102430, 102430, 102420, 
    102410, 102410, 102400, 102400, 102390, 102380, 102370, 102330, 102300, 
    102290, 102250, 102200, 102180, 102150, 102130, 102090, 102050, 101990, 
    101960, 101900, 101850, 101820, 101770, 101750, 101680, 101650, 101590, 
    101550, 101520, 101500, 101460, 101420, 101370, 101330, 101290, 101250, 
    101200, 101170, 101140, 101130, 101140, 101160, 101150, 101160, 101190, 
    101190, 101210, 101210, 101200, 101190, 101190, 101200, 101240, 101240, 
    101260, 101280, 101300, 101350, 101360, 101380, 101420, 101430, 101430, 
    101460, 101480, 101500, 101510, 101470, 101500, 101510, 101510, 101500, 
    101500, 101520, 101520, 101530, 101540, 101540, 101530, 101520, 101510, 
    101510, 101500, 101480, 101510, 101440, 101450, 101430, 101430, 101420, 
    101410, 101400, 101360, 101310, 101330, 101300, 101290, 101280, 101250, 
    101240, 101240, 101240, 101240, 101230, 101210, 101190, 101150, 101120, 
    101090, 101080, 101050, 101020, 101010, 100990, 100950, 100910, 100880, 
    100830, 100800, 100770, 100700, 100660, 100650, 100670, 100720, 100790, 
    100860, 100900, 100950, 100990, 101050, 101100, 101160, 101210, 101270, 
    101320, 101390, 101460, 101550, 101610, 101660, 101730, 101780, 101820, 
    101900, 101960, 102030, 102100, 102180, 102240, 102310, 102340, 102370, 
    102400, 102430, 102460, 102510, 102550, 102600, 102630, 102680, 102720, 
    102760, 102790, 102780, 102800, 102810, 102840, 102850, 102870, 102900, 
    102910, 102940, 102970, 102960, 102960, 102960, 102940, 102930, 102930, 
    102910, 102890, 102890, 102890, 102880, 102860, 102860, 102830, 102780, 
    102720, 102680, 102660, 102620, 102580, 102540, 102500, 102460, 102440, 
    102420, 102400, 102400, 102380, 102360, 102330, 102320, 102310, 102330, 
    102350, 102370, 102390, 102400, 102410, 102390, 102360, 102340, 102330, 
    102330, 102340, 102330, 102330, 102340, 102320, 102320, 102300, 102280, 
    102270, 102240, 102220, 102220, 102200, 102200, 102210, 102210, 102200, 
    102210, 102200, 102170, 102150, 102120, 102110, 102100, 102090, 102110, 
    102120, 102130, 102130, 102130, 102130, 102130, 102140, 102140, 102130, 
    102140, 102130, 102150, 102150, 102170, 102180, 102190, 102210, 102210, 
    102180, 102190, 102180, 102190, 102190, 102200, 102220, 102210, 102210, 
    102230, 102210, 102190, 102160, 102140, 102080, 102050, 102020, 102000, 
    102020, 101990, 101970, 101920, 101900, 101840, 101790, 101730, 101660, 
    101620, 101560, 101500, 101470, 101410, 101370, 101310, 101260, 101190, 
    101170, 101130, 101100, 101050, 101020, 101020, 101000, 100990, 100970, 
    100960, 100960, 100960, 100930, 100880, 100860, 100850, 100810, 100800, 
    100800, 100810, 100810, 100810, 100830, 100830, 100850, 100820, 100810, 
    100830, 100830, 100860, 100870, 100870, 100870, 100860, 100850, 100840, 
    100840, 100850, 100830, 100810, 100780, 100800, 100780, 100770, 100750, 
    100720, 100690, 100640, 100620, 100610, 100570, 100570, 100570, 100550, 
    100540, 100550, 100550, 100530, 100510, 100500, 100480, 100450, 100440, 
    100420, 100420, 100400, 100380, 100360, 100340, 100320, 100300, 100280, 
    100250, 100220, 100190, 100190, 100190, 100200, 100210, 100210, 100200, 
    100200, 100220, 100200, 100190, 100170, 100160, 100150, 100150, 100140, 
    100140, 100140, 100160, 100150, 100140, 100170, 100180, 100170, 100190, 
    100210, 100220, 100250, 100280, 100320, 100330, 100340, 100370, 100420, 
    100450, 100460, 100470, 100490, 100510, 100510, 100550, 100560, 100600, 
    100620, 100600, 100620, 100640, 100650, 100670, 100680, 100700, 100700, 
    100740, 100740, 100770, 100780, 100790, 100800, 100780, 100770, 100740, 
    100720, 100700, 100690, 100670, 100630, 100610, 100580, 100560, 100530, 
    100510, 100490, 100460, 100450, 100450, 100440, 100470, 100480, 100490, 
    100500, 100500, 100500, 100470, 100490, 100490, 100460, 100430, 100420, 
    100400, 100380, 100360, 100320, 100280, 100240, 100210, 100160, 100080, 
    100000, 99920, 99850, 99810, 99750, 99710, 99640, 99570, 99530, 99490, 
    99460, 99440, 99440, 99420, 99420, 99430, 99470, 99510, 99560, 99610, 
    99650, 99680, 99770, 99820, 99880, 99920, 99970, 100050, 100100, 100140, 
    100200, 100240, 100270, 100310, 100350, 100350, 100380, 100410, 100420, 
    100430, 100460, 100500, 100510, 100490, 100450, 100440, 100410, 100400, 
    100400, 100390, 100400, 100410, 100440, 100470, 100490, 100520, 100540, 
    100580, 100630, 100710, 100780, 100840, 100920, 100980, 101050, 101090, 
    101140, 101180, 101220, 101270, 101340, 101390, 101420, 101470, 101500, 
    101580, 101630, 101690, 101720, 101780, 101810, 101830, 101830, 101850, 
    101860, 101840, 101830, 101820, 101820, 101840, 101840, 101790, 101780, 
    101750, 101700, 101680, 101650, 101650, 101620, 101590, 101580, 101550, 
    101520, 101490, 101430, 101400, 101350, 101300, 101270, 101250, 101230, 
    101220, 101180, 101140, 101110, 101080, 101060, 101000, 100960, 100890, 
    100850, 100810, 100760, 100740, 100730, 100730, 100690, 100670, 100650, 
    100640, 100630, 100610, 100600, 100620, 100640, 100640, 100660, 100680, 
    100690, 100670, 100670, 100670, 100680, 100690, 100700, 100710, 100730, 
    100740, 100770, 100790, 100760, 100750, 100730, 100650, 100610, 100540, 
    100480, 100430, 100390, 100340, 100340, 100340, 100370, 100380, 100400, 
    100440, 100490, 100520, 100570, 100630, 100650, 100680, 100710, 100690, 
    100680, 100730, 100710, 100650, 100570, 100470, 100360, 100180, 100020, 
    99920, 99840, 99770, 99740, 99650, 99600, 99570, 99500, 99460, 99340, 
    99210, 99090, 98940, 98770, 98610, 98460, 98310, 98220, 98140, 98100, 
    98100, 98080, 98080, 98080, 98110, 98130, 98170, 98230, 98280, 98340, 
    98410, 98510, 98600, 98670, 98800, 98920, 99010, 99120, 99230, 99320, 
    99400, 99480, 99530, 99600, 99660, 99660, 99720, 99720, 99720, 99740, 
    99730, 99710, 99640, 99570, 99520, 99470, 99390, 99300, 99300, 99260, 
    99260, 99270, 99310, 99390, 99460, 99560, 99650, 99750, 99930, 100050, 
    100160, 100330, 100530, 100710, 100820, 100930, 101050, 101150, 101250, 
    101320, 101410, 101430, 101460, 101510, 101560, 101590, 101630, 101620, 
    101640, 101630, 101630, 101580, 101560, 101530, 101520, 101530, 101530, 
    101570, 101560, 101550, 101560, 101560, 101530, 101500, 101430, 101380, 
    101370, 101360, 101370, 101380, 101360, 101320, 101180, 101120, 101060, 
    100990, 100910, 100790, 100680, 100630, 100630, 100620, 100610, 100580, 
    100570, 100580, 100590, 100590, 100620, 100650, 100660, 100750, 100800, 
    100830, 100890, 100940, 100970, 101000, 101040, 101060, 101060, 101020, 
    101000, 101000, 100990, 100960, 100970, 100940, 100940, 100920, 100910, 
    100910, 100850, 100830, 100870, 100860, 100880, 100900, 100950, 100950, 
    101020, 101070, 101070, 101120, 101100, 101110, 101150, 101170, 101150, 
    101190, 101150, 101200, 101240, 101230, 101260, 101260, 101260, 101240, 
    101270, 101270, 101240, 101220, 101260, 101240, 101200, 101180, 101120, 
    101070, 101010, 100990, 100920, 100870, 100780, 100720, 100660, 100580, 
    100470, 100350, 100250, 100200, 100190, 100170, 100120, 100100, 100100, 
    100080, 100110, 100090, 100110, 100120, 100050, 100040, 100030, 100040, 
    99990, 99960, 99940, 99920, 99900, 99900, 99880, 99880, 99880, 99870, 
    99870, 99860, 99940, 99960, 99990, 100060, 100040, 100100, 100100, 
    100100, 100050, 100120, 100120, 100130, 100170, 100180, 100180, 100210, 
    100240, 100250, 100240, 100160, 100170, 100110, 100100, 100040, 99930, 
    99900, 99850, 99780, 99770, 99700, 99710, 99660, 99630, 99620, 99590, 
    99560, 99540, 99500, 99480, 99430, 99400, 99350, 99320, 99290, 99240, 
    99200, 99210, 99200, 99220, 99240, 99260, 99260, 99300, 99350, 99370, 
    99360, 99320, 99370, 99340, 99350, 99340, 99320, 99350, 99390, 99460, 
    99510, 99520, 99530, 99560, 99560, 99570, 99570, 99620, 99630, 99700, 
    99820, 99880, 100010, 100130, 100190, 100240, 100320, 100430, 100470, 
    100470, 100520, 100560, 100580, 100570, 100580, 100620, 100670, 100640, 
    100710, 100740, 100740, 100700, 100750, 100760, 100780, 100790, 100790, 
    100810, 100810, 100830, 100850, 100860, 100880, 100880, 100870, 100880, 
    100870, 100880, 100890, 100880, 100910, 100890, 100880, 100860, 100860, 
    100860, 100880, 100880, 100920, 100930, 100940, 100940, 100950, 100940, 
    100900, 100890, 100870, 100850, 100810, 100800, 100780, 100740, 100710, 
    100690, 100650, 100630, 100600, 100540, 100490, 100480, 100450, 100410, 
    100410, 100350, 100350, 100300, 100270, 100210, 100150, 100120, 100070, 
    100030, 100030, 100030, 100000, 99990, 99990, 99970, 99960, 99970, 99950, 
    99940, 99950, 99970, 99970, 99990, 100000, 100020, 100030, 100040, 
    100060, 100080, 100080, 100100, 100110, 100120, 100150, 100190, 100230, 
    100260, 100280, 100300, 100330, 100360, 100400, 100420, 100450, 100450, 
    100500, 100530, 100550, 100570, 100600, 100600, 100600, 100600, 100600, 
    100600, 100610, 100600, 100590, 100590, 100580, 100580, 100580, 100570, 
    100560, 100520, 100510, 100480, 100470, 100470, 100450, 100430, 100410, 
    100430, 100400, 100360, 100370, 100360, 100330, 100320, 100330, 100330, 
    100330, 100370, 100360, 100360, 100340, 100350, 100330, 100320, 100340, 
    100320, 100310, 100300, 100310, 100320, 100350, 100370, 100350, 100320, 
    100310, 100300, 100280, 100240, 100220, 100190, 100190, 100150, 100140, 
    100140, 100130, 100090, 100060, 100060, 100040, 100020, 100010, 99990, 
    99990, 100000, 100010, 100010, 99990, 99980, 99950, 99930, 99910, 99920, 
    99910, 99880, 99900, 99870, 99890, 99910, 99910, 99900, 99910, 99930, 
    99920, 99880, 99900, 99940, 99960, 99990, 100000, 100030, 100050, 100050, 
    100070, 100090, 100120, 100140, 100170, 100200, 100230, 100280, 100300, 
    100330, 100350, 100370, 100390, 100440, 100440, 100450, 100440, 100460, 
    100480, 100500, 100510, 100510, 100530, 100540, 100540, 100550, 100560, 
    100580, 100580, 100590, 100610, 100640, 100600, 100580, 100590, 100590, 
    100600, 100560, 100570, 100540, 100520, 100490, 100500, 100510, 100480, 
    100500, 100500, 100430, 100460, 100480, 100490, 100480, 100470, 100440, 
    100430, 100440, 100460, 100450, 100450, 100460, 100430, 100370, 100330, 
    100270, 100200, 100030, 99910, 99790, 99670, 99580, 99410, 99230, 99150, 
    98980, 99030, 99130, 99220, 99270, 99470, 99680, 99860, 100010, 100070, 
    100120, 100250, 100310, 100370, 100390, 100430, 100490, 100580, 100630, 
    100660, 100730, 100730, 100710, 100650, 100610, 100550, 100450, 100370, 
    100300, 100280, 100140, 100060, 99890, 99690, 99560, 99440, 99310, 99170, 
    99020, 98900, 98760, 98680, 98590, 98580, 98550, 98570, 98590, 98630, 
    98710, 98790, 98870, 98950, 99000, 99050, 99090, 99160, 99210, 99230, 
    99210, 99220, 99190, 99170, 99170, 99110, 99070, 99040, 99030, 99010, 
    98970, 98940, 98880, 98850, 98840, 98810, 98760, 98710, 98670, 98640, 
    98590, 98540, 98460, 98400, 98370, 98290, 98210, 98100, 97990, 97970, 
    97920, 97900, 97880, 97870, 97880, 97900, 97900, 97930, 97980, 98030, 
    98110, 98160, 98170, 98210, 98230, 98270, 98260, 98240, 98220, 98170, 
    98100, 98090, 98050, 98020, 97990, 97930, 97920, 97940, 97930, 97910, 
    97900, 97910, 97930, 97980, 98010, 98080, 98100, 98130, 98180, 98240, 
    98300, 98360, 98440, 98500, 98560, 98650, 98700, 98760, 98830, 98900, 
    99000, 99030, 99120, 99170, 99200, 99230, 99250, 99280, 99330, 99360, 
    99390, 99360, 99340, 99380, 99400, 99390, 99350, 99310, 99290, 99280, 
    99320, 99460, 99520, 99590, 99630, 99790, 99860, 99920, 100030, 100110, 
    100150, 100200, 100280, 100350, 100410, 100480, 100600, 100630, 100700, 
    100730, 100770, 100760, 100810, 100840, 100810, 100800, 100790, 100790, 
    100790, 100790, 100790, 100760, 100730, 100650, 100580, 100530, 100460, 
    100390, 100340, 100280, 100210, 100180, 100130, 100090, 100030, 99950, 
    99910, 99860, 99820, 99770, 99720, 99680, 99650, 99620, 99590, 99560, 
    99480, 99440, 99450, 99420, 99390, 99310, 99280, 99220, 99200, 99160, 
    99090, 99020, 98980, 98890, 98820, 98750, 98670, 98640, 98590, 98520, 
    98470, 98470, 98450, 98390, 98340, 98290, 98220, 98170, 98110, 98050, 
    97960, 97890, 97810, 97730, 97680, 97590, 97560, 97630, 97650, 97630, 
    97610, 97630, 97640, 97700, 97780, 97860, 97880, 97870, 97930, 97950, 
    97900, 98040, 98090, 98170, 98230, 98340, 98410, 98470, 98560, 98670, 
    98740, 98790, 98870, 98910, 99000, 99070, 99110, 99140, 99180, 99210, 
    99240, 99240, 99250, 99250, 99270, 99270, 99340, 99370, 99410, 99430, 
    99460, 99460, 99460, 99470, 99450, 99440, 99440, 99410, 99450, 99490, 
    99460, 99440, 99430, 99450, 99490, 99480, 99470, 99500, 99530, 99520, 
    99530, 99510, 99530, 99570, 99560, 99570, 99610, 99610, 99620, 99620, 
    99640, 99630, 99660, 99660, 99670, 99690, 99700, 99750, 99760, 99780, 
    99810, 99820, 99830, 99810, 99790, 99790, 99820, 99800, 99840, 99870, 
    99900, 99910, 99950, 99950, 99950, 99990, 100000, 99980, 100010, 100040, 
    100100, 100140, 100160, 100170, 100210, 100240, 100270, 100310, 100330, 
    100360, 100400, 100430, 100470, 100510, 100550, 100570, 100590, 100600, 
    100640, 100640, 100650, 100660, 100690, 100730, 100790, 100800, 100830, 
    100870, 100890, 100920, 100940, 100950, 101000, 101020, 101050, 101090, 
    101120, 101200, 101230, 101240, 101250, 101310, 101340, 101330, 101370, 
    101380, 101410, 101440, 101460, 101520, 101510, 101520, 101510, 101490, 
    101420, 101360, 101230, 101090, 100980, 100840, 100650, 100520, 100360, 
    100190, 100030, 99990, 99910, 99930, 99970, 100040, 100060, 100090, 
    100140, 100200, 100270, 100370, 100460, 100590, 100640, 100730, 100770, 
    100790, 100800, 100810, 100820, 100820, 100810, 100680, 100650, 100610, 
    100580, 100550, 100540, 100540, 100560, 100610, 100650, 100730, 100800, 
    100880, 100940, 101040, 101210, 101310, 101440, 101580, 101700, 101830, 
    101940, 102010, 102110, 102180, 102240, 102290, 102370, 102440, 102530, 
    102570, 102630, 102690, 102720, 102760, 102780, 102790, 102800, 102810, 
    102790, 102800, 102800, 102820, 102840, 102870, 102940, 102990, 103000, 
    103020, 103040, 103080, 103120, 103190, 103230, 103240, 103270, 103290, 
    103300, 103330, 103360, 103390, 103400, 103420, 103410, 103420, 103400, 
    103400, 103390, 103390, 103390, 103310, 103240, 103200, 103160, 103130, 
    103030, 102960, 102910, 102810, 102710, 102600, 102520, 102450, 102420, 
    102390, 102340, 102310, 102290, 102240, 102210, 102170, 102140, 102100, 
    102060, 102030, 101980, 101910, 101860, 101810, 101770, 101740, 101690, 
    101620, 101580, 101520, 101490, 101460, 101430, 101420, 101400, 101400, 
    101400, 101390, 101390, 101410, 101430, 101450, 101450, 101480, 101510, 
    101550, 101580, 101600, 101610, 101630, 101660, 101680, 101710, 101780, 
    101830, 101890, 101960, 102010, 102050, 102100, 102130, 102160, 102180, 
    102200, 102210, 102240, 102250, 102280, 102270, 102260, 102270, 102270, 
    102250, 102230, 102190, 102170, 102150, 102120, 102090, 102040, 102020, 
    101970, 101960, 101920, 101850, 101810, 101760, 101730, 101680, 101650, 
    101640, 101610, 101550, 101560, 101520, 101500, 101450, 101420, 101390, 
    101390, 101360, 101360, 101390, 101410, 101390, 101400, 101410, 101380, 
    101380, 101320, 101320, 101250, 101240, 101270, 101290, 101290, 101270, 
    101270, 101300, 101320, 101240, 101150, 101090, 101000, 100950, 100870, 
    100770, 100770, 100730, 100740, 100770, 100830, 100840, 100840, 100880, 
    100910, 100940, 100980, 101040, 101090, 101150, 101200, 101280, 101400, 
    101500, 101600, 101700, 101790, 101890, 101950, 102040, 102130, 102160, 
    102170, 102180, 102160, 102120, 102060, 102000, 101970, 101940, 101880, 
    101820, 101770, 101700, 101630, 101630, 101590, 101540, 101550, 101520, 
    101490, 101520, 101540, 101590, 101610, 101620, 101630, 101620, 101560, 
    101500, 101470, 101450, 101400, 101320, 101270, 101250, 101240, 101250, 
    101240, 101300, 101340, 101410, 101450, 101510, 101560, 101640, 101720, 
    101780, 101850, 101890, 101920, 101940, 101920, 101940, 101910, 101870, 
    101830, 101810, 101750, 101680, 101660, 101640, 101640, 101570, 101540, 
    101530, 101520, 101480, 101440, 101440, 101450, 101450, 101450, 101450, 
    101450, 101450, 101430, 101440, 101430, 101400, 101350, 101290, 101260, 
    101230, 101230, 101260, 101230, 101180, 101160, 101180, 101170, 101130, 
    101110, 101110, 101120, 101110, 101080, 101050, 101020, 100930, 100830, 
    100730, 100620, 100530, 100450, 100330, 100210, 100170, 100150, 100150, 
    100140, 100170, 100300, 100450, 100570, 100670, 100740, 100800, 100840, 
    100800, 100830, 100860, 100830, 100810, 100750, 100660, 100570, 100520, 
    100410, 100290, 100220, 100190, 100140, 100110, 100070, 100000, 99960, 
    99940, 99930, 99940, 99930, 99930, 99950, 99980, 100040, 100080, 100100, 
    100140, 100170, 100240, 100370, 100450, 100530, 100620, 100690, 100770, 
    100860, 100940, 101010, 101090, 101160, 101190, 101230, 101270, 101310, 
    101350, 101400, 101430, 101450, 101440, 101450, 101440, 101430, 101390, 
    101340, 101330, 101300, 101260, 101200, 101180, 101170, 101140, 101130, 
    101080, 101050, 101040, 101020, 101020, 101040, 101050, 101070, 101100, 
    101120, 101150, 101170, 101210, 101250, 101290, 101330, 101360, 101400, 
    101450, 101480, 101530, 101580, 101640, 101690, 101740, 101830, 101900, 
    101960, 102040, 102100, 102160, 102210, 102250, 102330, 102390, 102400, 
    102430, 102460, 102440, 102450, 102420, 102420, 102390, 102400, 102440, 
    102450, 102460, 102460, 102470, 102480, 102490, 102500, 102490, 102470, 
    102470, 102480, 102490, 102490, 102490, 102490, 102460, 102460, 102430, 
    102400, 102350, 102300, 102290, 102250, 102240, 102230, 102250, 102240, 
    102240, 102240, 102250, 102260, 102270, 102290, 102310, 102330, 102360, 
    102390, 102450, 102490, 102520, 102560, 102610, 102640, 102670, 102680, 
    102710, 102720, 102750, 102770, 102800, 102800, 102810, 102810, 102780, 
    102770, 102750, 102730, 102710, 102700, 102700, 102700, 102700, 102690, 
    102660, 102630, 102620, 102600, 102560, 102530, 102510, 102470, 102460, 
    102440, 102410, 102380, 102360, 102350, 102350, 102360, 102360, 102370, 
    102380, 102410, 102430, 102450, 102490, 102510, 102530, 102550, 102580, 
    102610, 102600, 102600, 102620, 102640, 102680, 102690, 102700, 102700, 
    102700, 102690, 102680, 102630, 102590, 102540, 102500, 102440, 102400, 
    102350, 102280, 102220, 102110, 102010, 101910, 101830, 101730, 101680, 
    101700, 101730, 101830, 101910, 101920, 101930, 102010, 102050, 102100, 
    102120, 102110, 102100, 102090, 102130, 102120, 102140, 102100, 102080, 
    102050, 102050, 101980, 102010, 101970, 101950, 101920, 101850, 101850, 
    101840, 101850, 101850, 101800, 101770, 101730, 101690, 101660, 101630, 
    101620, 101620, 101660, 101700, 101740, 101760, 101800, 101860, 101800, 
    101860, 101940, 102020, 102110, 102130, 102280, 102360, 102490, 102530, 
    102590, 102560, 102560, 102610, 102650, 102730, 102710, 102730, 102750, 
    102730, 102710, 102720, 102690, 102580, 102440, 102390, 102280, 102130, 
    101970, 101810, 101740, 101600, 101450, 101350, 101290, 101220, 101160, 
    101080, 101130, 101070, 101030, 101010, 101000, 100990, 101010, 101050, 
    101090, 101140, 101130, 101140, 101200, 101180, 101250, 101280, 101280, 
    101320, 101350, 101380, 101380, 101450, 101480, 101530, 101550, 101640, 
    101700, 101770, 101820, 101910, 101940, 101990, 102050, 102070, 102130, 
    102130, 102170, 102170, 102200, 102240, 102280, 102250, 102290, 102320, 
    102350, 102340, 102340, 102330, 102340, 102330, 102340, 102300, 102310, 
    102300, 102290, 102290, 102290, 102300, 102280, 102260, 102240, 102220, 
    102210, 102170, 102160, 102130, 102080, 102070, 102060, 102040, 102010, 
    102040, 102070, 102080, 102070, 102070, 102100, 102110, 102130, 102130, 
    102140, 102160, 102180, 102160, 102140, 102150, 102190, 102240, 102280, 
    102290, 102320, 102370, 102380, 102390, 102440, 102460, 102460, 102470, 
    102520, 102520, 102520, 102530, 102540, 102540, 102550, 102520, 102520, 
    102520, 102540, 102530, 102560, 102590, 102610, 102640, 102680, 102660, 
    102710, 102730, 102730, 102730, 102740, 102770, 102790, 102810, 102830, 
    102810, 102800, 102790, 102770, 102750, 102730, 102700, 102680, 102620, 
    102600, 102570, 102500, 102470, 102440, 102400, 102360, 102310, 102250, 
    102170, 102080, 102040, 102020, 101970, 101990, 101980, 101980, 101940, 
    101950, 101950, 101960, 101970, 101990, 102000, 102020, 102040, 102090, 
    102120, 102200, 102270, 102340, 102390, 102440, 102480, 102520, 102550, 
    102580, 102610, 102660, 102720, 102750, 102780, 102810, 102820, 102840, 
    102870, 102890, 102920, 102950, 102990, 103030, 103060, 103090, 103100, 
    103110, 103120, 103110, 103110, 103110, 103100, 103100, 103120, 103120, 
    103120, 103120, 103100, 103090, 103090, 103070, 103060, 103050, 103060, 
    103070, 103070, 103090, 103090, 103090, 103110, 103130, 103130, 103090, 
    103080, 103090, 103110, 103090, 103110, 103150, 103160, 103140, 103170, 
    103160, 103090, 103060, 103050, 103020, 103000, 102990, 102970, 102970, 
    102940, 102930, 102850, 102800, 102770, 102740, 102650, 102600, 102550, 
    102500, 102460, 102450, 102420, 102360, 102310, 102200, 102060, 102000, 
    101970, 101890, 101800, 101770, 101720, 101700, 101660, 101610, 101550, 
    101490, 101440, 101400, 101350, 101310, 101260, 101230, 101200, 101180, 
    101150, 101100, 101080, 101000, 100960, 100930, 100890, 100830, 100780, 
    100750, 100740, 100730, 100730, 100700, 100710, 100710, 100710, 100730, 
    100740, 100740, 100750, 100770, 100800, 100820, 100860, 100870, 100890, 
    100920, 100970, 101020, 101060, 101070, 101090, 101110, 101130, 101180, 
    101200, 101230, 101250, 101270, 101330, 101340, 101370, 101410, 101390, 
    101410, 101480, 101550, 101600, 101640, 101690, 101760, 101830, 101880, 
    101930, 101970, 101990, 102040, 102080, 102130, 102170, 102200, 102220, 
    102230, 102270, 102280, 102300, 102310, 102340, 102350, 102380, 102390, 
    102410, 102420, 102440, 102460, 102470, 102500, 102520, 102510, 102510, 
    102560, 102560, 102570, 102580, 102610, 102620, 102640, 102670, 102690, 
    102720, 102720, 102730, 102740, 102770, 102790, 102820, 102860, 102870, 
    102880, 102900, 102910, 102930, 102890, 102920, 102910, 102910, 102930, 
    102950, 102970, 102980, 102960, 102940, 102940, 102940, 102940, 102960, 
    102960, 102960, 102970, 102980, 103020, 103030, 103040, 103040, 103070, 
    103080, 103070, 103050, 103040, 103030, 103030, 103040, 103020, 103030, 
    103020, 103010, 102980, 102970, 102970, 102960, 102970, 102980, 102990, 
    103000, 103010, 103030, 103020, 103030, 103030, 103040, 103040, 103040, 
    103030, 103020, 103030, 103030, 103010, 103000, 103020, 103020, 103010, 
    102990, 102980, 102970, 102960, 102960, 102960, 102960, 102960, 102960, 
    102970, 102950, 102950, 102950, 102940, 102960, 102980, 103000, 103020, 
    103060, 103090, 103100, 103150, 103150, 103160, 103140, 103150, 103150, 
    103130, 103130, 103110, 103090, 103070, 103040, 103030, 102990, 102980, 
    102930, 102890, 102860, 102810, 102790, 102760, 102720, 102750, 102720, 
    102690, 102680, 102630, 102590, 102550, 102530, 102490, 102440, 102430, 
    102380, 102360, 102340, 102290, 102230, 102170, 102110, 102060, 102010, 
    101970, 101950, 101910, 101860, 101820, 101790, 101710, 101740, 101720, 
    101710, 101700, 101680, 101670, 101640, 101620, 101640, 101650, 101640, 
    101640, 101640, 101650, 101650, 101610, 101630, 101620, 101640, 101670, 
    101700, 101710, 101740, 101760, 101790, 101770, 101750, 101760, 101730, 
    101700, 101680, 101660, 101620, 101590, 101560, 101530, 101510, 101480, 
    101460, 101440, 101410, 101380, 101340, 101330, 101310, 101300, 101330, 
    101360, 101350, 101350, 101350, 101390, 101380, 101410, 101450, 101490, 
    101550, 101550, 101630, 101690, 101700, 101710, 101710, 101710, 101710, 
    101730, 101770, 101780, 101790, 101800, 101820, 101840, 101860, 101870, 
    101870, 101890, 101900, 101900, 101910, 101920, 101930, 101910, 101910, 
    101900, 101890, 101860, 101840, 101810, 101780, 101780, 101770, 101760, 
    101760, 101740, 101710, 101660, 101640, 101610, 101560, 101500, 101500, 
    101460, 101420, 101400, 101390, 101380, 101380, 101380, 101390, 101400, 
    101400, 101410, 101410, 101400, 101410, 101420, 101440, 101460, 101470, 
    101500, 101510, 101540, 101570, 101610, 101640, 101700, 101770, 101820, 
    101880, 101920, 101960, 102010, 102040, 102070, 102100, 102140, 102170, 
    102210, 102240, 102270, 102260, 102260, 102290, 102310, 102330, 102350, 
    102350, 102290, 102280, 102260, 102240, 102300, 102250, 102200, 102150, 
    102120, 102110, 102100, 102080, 102040, 102010, 101950, 101920, 101870, 
    101840, 101800, 101820, 101750, 101650, 101620, 101630, 101710, 101920, 
    101680, 101670, 101610, 101690, 101660, 101640, 101660, 101730, 101750, 
    101760, 101760, 101740, 101760, 101790, 101790, 101790, 101770, 101760, 
    101760, 101800, 101800, 101810, 101810, 101780, 101780, 101780, 101750, 
    101770, 101820, 101830, 101850, 101850, 101780, 101780, 101740, 101700, 
    101680, 101650, 101650, 101630, 101600, 101570, 101530, 101520, 101490, 
    101440, 101400, 101350, 101300, 101280, 101250, 101270, 101250, 101240, 
    101250, 101230, 101190, 101160, 101140, 101140, 101130, 101130, 101140, 
    101130, 101110, 101110, 101100, 101090, 101100, 101080, 101060, 101060, 
    101030, 101040, 101030, 101040, 101050, 101040, 101040, 101030, 101040, 
    101010, 100990, 100960, 100920, 100900, 100870, 100870, 100850, 100850, 
    100830, 100830, 100840, 100820, 100830, 100840, 100830, 100850, 100850, 
    100870, 100880, 100880, 100900, 100920, 100920, 100920, 100930, 100930, 
    100930, 100930, 100940, 100940, 100970, 100980, 100990, 101000, 100990, 
    100990, 100980, 100990, 100990, 101000, 101030, 101030, 101050, 101070, 
    101060, 101080, 101060, 101040, 101040, 101040, 101060, 101070, 101080, 
    101090, 101100, 101110, 101100, 101080, 101110, 101120, 101110, 101110, 
    101120, 101130, 101150, 101160, 101180, 101170, 101190, 101200, 101230, 
    101240, 101250, 101280, 101300, 101310, 101330, 101360, 101380, 101410, 
    101440, 101460, 101490, 101480, 101490, 101500, 101520, 101560, 101560, 
    101610, 101610, 101630, 101670, 101680, 101680, 101680, 101660, 101650, 
    101650, 101660, 101690, 101720, 101750, 101760, 101760, 101760, 101780, 
    101770, 101810, 101830, 101840, 101840, 101880, 101910, 101920, 101960, 
    101980, 101990, 102010, 102030, 102050, 102070, 102090, 102130, 102180, 
    102210, 102230, 102240, 102270, 102270, 102290, 102300, 102310, 102310, 
    102330, 102350, 102350, 102350, 102380, 102370, 102370, 102380, 102360, 
    102360, 102360, 102340, 102350, 102340, 102360, 102360, 102370, 102360, 
    102350, 102340, 102330, 102290, 102260, 102250, 102230, 102250, 102260, 
    102270, 102310, 102290, 102280, 102300, 102320, 102340, 102350, 102370, 
    102390, 102390, 102420, 102460, 102480, 102490, 102500, 102500, 102500, 
    102500, 102480, 102480, 102480, 102490, 102500, 102520, 102520, 102520, 
    102530, 102520, 102530, 102540, 102530, 102520, 102520, 102520, 102530, 
    102540, 102550, 102570, 102560, 102580, 102610, 102600, 102600, 102620, 
    102630, 102680, 102690, 102750, 102770, 102780, 102800, 102800, 102810, 
    102800, 102770, 102800, 102760, 102780, 102760, 102750, 102770, 102730, 
    102710, 102690, 102630, 102590, 102560, 102510, 102470, 102390, 102350, 
    102310, 102250, 102220, 102170, 102100, 102090, 102070, 102070, 102050, 
    102020, 102020, 101980, 101990, 101970, 101930, 101900, 101900, 101850, 
    101810, 101840, 101830, 101850, 101880, 101910, 101940, 101960, 101930, 
    101910, 101860, 101810, 101800, 101750, 101720, 101640, 101560, 101520, 
    101450, 101410, 101340, 101290, 101230, 101160, 101120, 101100, 101080, 
    101040, 101020, 101020, 101020, 101040, 101060, 101080, 101080, 101060, 
    101080, 101080, 101100, 101120, 101140, 101140, 101130, 101160, 101150, 
    101130, 101060, 101020, 101000, 101000, 100990, 101060, 100990, 100990, 
    101010, 100980, 100950, 100930, 100910, 100900, 100910, 100920, 100930, 
    100900, 100900, 100870, 100870, 100900, 100880, 100890, 100900, 100890, 
    100870, 100880, 100880, 100880, 100890, 100890, 100910, 100940, 100970, 
    100980, 100990, 100980, 100970, 100980, 100970, 100970, 100950, 100950, 
    100940, 100930, 100910, 100890, 100880, 100870, 100850, 100840, 100830, 
    100810, 100780, 100810, 100810, 100810, 100800, 100830, 100850, 100880, 
    100890, 100880, 100890, 100920, 100910, 100910, 100900, 100880, 100870, 
    100870, 100860, 100840, 100830, 100810, 100780, 100760, 100770, 100780, 
    100820, 100840, 100870, 100890, 100900, 100900, 100910, 100910, 100910, 
    100920, 100930, 100960, 101000, 101020, 101030, 101080, 101100, 101130, 
    101140, 101150, 101170, 101190, 101220, 101260, 101290, 101330, 101360, 
    101390, 101410, 101430, 101450, 101470, 101470, 101470, 101490, 101520, 
    101530, 101560, 101570, 101570, 101570, 101570, 101560, 101550, 101530, 
    101510, 101490, 101480, 101480, 101490, 101460, 101440, 101440, 101420, 
    101420, 101400, 101380, 101380, 101370, 101370, 101370, 101380, 101390, 
    101370, 101390, 101400, 101380, 101370, 101340, 101330, 101330, 101350, 
    101360, 101360, 101350, 101370, 101380, 101390, 101400, 101400, 101400, 
    101400, 101400, 101410, 101400, 101440, 101460, 101470, 101480, 101500, 
    101510, 101510, 101530, 101520, 101540, 101570, 101590, 101610, 101640, 
    101660, 101680, 101680, 101700, 101710, 101690, 101700, 101700, 101710, 
    101700, 101730, 101720, 101710, 101710, 101690, 101680, 101650, 101620, 
    101590, 101560, 101520, 101510, 101480, 101450, 101430, 101380, 101360, 
    101340, 101290, 101250, 101210, 101190, 101160, 101140, 101110, 101080, 
    101070, 101020, 101000, 100960, 100930, 100890, 100850, 100820, 100810, 
    100810, 100770, 100760, 100760, 100740, 100720, 100690, 100680, 100640, 
    100630, 100630, 100620, 100610, 100650, 100610, 100600, 100610, 100570, 
    100560, 100520, 100490, 100470, 100470, 100440, 100400, 100370, 100350, 
    100300, 100270, 100210, 100150, 100100, 100020, 99960, 99890, 99830, 
    99780, 99720, 99650, 99600, 99560, 99500, 99470, 99420, 99400, 99390, 
    99420, 99450, 99470, 99520, 99560, 99570, 99590, 99640, 99660, 99670, 
    99690, 99680, 99680, 99700, 99710, 99720, 99790, 99820, 99860, 99880, 
    99940, 100000, 100070, 100100, 100160, 100190, 100240, 100290, 100310, 
    100340, 100370, 100390, 100380, 100420, 100440, 100440, 100430, 100450, 
    100430, 100430, 100430, 100370, 100360, 100380, 100350, 100330, 100380, 
    100440, 100420, 100420, 100450, 100470, 100500, 100520, 100550, 100560, 
    100600, 100640, 100650, 100650, 100710, 100800, 100860, 100930, 100980, 
    101000, 101070, 101090, 101090, 101160, 101180, 101250, 101270, 101290, 
    101310, 101290, 101270, 101240, 101200, 101210, 101200, 101130, 101020, 
    100970, 100900, 100870, 100820, 100710, 100690, 100640, 100580, 100560, 
    100570, 100510, 100490, 100440, 100410, 100450, 100420, 100400, 100420, 
    100470, 100480, 100510, 100570, 100590, 100600, 100580, 100570, 100580, 
    100550, 100540, 100490, 100410, 100460, 100500, 100500, 100470, 100490, 
    100470, 100500, 100520, 100510, 100490, 100510, 100530, 100580, 100670, 
    100730, 100740, 100770, 100790, 100810, 100830, 100880, 100910, 100940, 
    100950, 100970, 101030, 101080, 101120, 101190, 101230, 101290, 101340, 
    101370, 101410, 101450, 101470, 101510, 101560, 101600, 101620, 101660, 
    101680, 101710, 101740, 101750, 101780, 101800, 101840, 101850, 101860, 
    101890, 101890, 101920, 101920, 101940, 101960, 101990, 101990, 101980, 
    102020, 102000, 101990, 101990, 101990, 101990, 101950, 102000, 102000, 
    101980, 101950, 101890, 101840, 101800, 101800, 101800, 101760, 101720, 
    101670, 101650, 101630, 101610, 101660, 101640, 101640, 101590, 101580, 
    101630, 101570, 101630, 101650, 101680, 101720, 101770, 101800, 101830, 
    101830, 101810, 101820, 101850, 101870, 101870, 101890, 101920, 101950, 
    101980, 101990, 102010, 102050, 102070, 102060, 102080, 102120, 102150, 
    102130, 102110, 102150, 102180, 102220, 102260, 102290, 102310, 102330, 
    102340, 102370, 102370, 102370, 102370, 102360, 102370, 102390, 102410, 
    102420, 102430, 102450, 102450, 102450, 102440, 102430, 102440, 102450, 
    102440, 102450, 102440, 102420, 102410, 102370, 102360, 102340, 102320, 
    102310, 102300, 102300, 102310, 102290, 102290, 102280, 102270, 102240, 
    102230, 102240, 102240, 102240, 102240, 102220, 102230, 102240, 102240, 
    102230, 102210, 102190, 102170, 102170, 102140, 102400, 102140, 102150, 
    102120, 102100, 102060, 102030, 102010, 101980, 101950, 101930, 101870, 
    101840, 101810, 101790, 101760, 101720, 101700, 101650, 101600, 101580, 
    101530, 101510, 101480, 101450, 101460, 101460, 101450, 101430, 101420, 
    101400, 101380, 101360, 101360, 101350, 101350, 101350, 101340, 101350, 
    101340, 101320, 101320, 101310, 101310, 101310, 101300, 101300, 101290, 
    101310, 101330, 101330, 101340, 101330, 101350, 101350, 101350, 101330, 
    101340, 101320, 101310, 101310, 101310, 101320, 101330, 101320, 101330, 
    101330, 101330, 101340, 101320, 101320, 101300, 101310, 101280, 101290, 
    101330, 101330, 101340, 101360, 101370, 101380, 101390, 101410, 101410, 
    101420, 101440, 101450, 101470, 101480, 101470, 101450, 101460, 101450, 
    101470, 101460, 101450, 101470, 101500, 101550, 101550, 101550, 101550, 
    101560, 101530, 101510, 101510, 101520, 101510, 101490, 101500, 101490, 
    101500, 101510, 101510, 101510, 101530, 101520, 101530, 101530, 101530, 
    101520, 101530, 101570, 101580, 101580, 101560, 101550, 101550, 101570, 
    101580, 101580, 101600, 101600, 101620, 101640, 101650, 101650, 101650, 
    101660, 101660, 101660, 101660, 101670, 101670, 101670, 101690, 101700, 
    101710, 101710, 101710, 101710, 101730, 101720, 101710, 101730, 101730, 
    101720, 101750, 101760, 101780, 101810, 101820, 101820, 101840, 101850, 
    101860, 101870, 101890, 101890, 101910, 101950, 101990, 102000, 101440, 
    101990, 102010, 102030, 102050, 102080, 102120, 102130, 102150, 102170, 
    102210, 102250, 102240, 102250, 102250, 102250, 102240, 102220, 102210, 
    102190, 102170, 102140, 102120, 102120, 102060, 102030, 101990, 101950, 
    101870, 101820, 101750, 101660, 101580, 101510, 101410, 101350, 101300, 
    101210, 101120, 101010, 100940, 100830, 100750, 100700, 100640, 100600, 
    100570, 100590, 100580, 100580, 100580, 100600, 100640, 100720, 100800, 
    100850, 100900, 100960, 101020, 101130, 101190, 101240, 101290, 101340, 
    101360, 101370, 101390, 101420, 101450, 101460, 101480, 101480, 101510, 
    101510, 101490, 101480, 101470, 101470, 101470, 101450, 101450, 101450, 
    101410, 101410, 101400, 101400, 101360, 101320, 101290, 101280, 101270, 
    101260, 101270, 101260, 101250, 101250, 101260, 101250, 101230, 101210, 
    101210, 101200, 101160, 101150, 101140, 101140, 101160, 101180, 101200, 
    101210, 101230, 101220, 101250, 101260, 101240, 101230, 101240, 101250, 
    101250, 101250, 101260, 101250, 101250, 101220, 101200, 101200, 101170, 
    101170, 101160, 101170, 101170, 101160, 101190, 101160, 101140, 101140, 
    101140, 101110, 101090, 101090, 101090, 101100, 101090, 101110, 101130, 
    101100, 101090, 101070, 101030, 101020, 101030, 101040, 101040, 101040, 
    101070, 101110, 101130, 101130, 101160, 101180, 101180, 101200, 101240, 
    101260, 101290, 101340, 101400, 101420, 101450, 101460, 101500, 101520, 
    101520, 101540, 101560, 101560, 101600, 101630, 101660, 101660, 101670, 
    101680, 101660, 101660, 101670, 101660, 101650, 101660, 101630, 101650, 
    101670, 101680, 101670, 101630, 101600, 101600, 101620, 101640, 101660, 
    101690, 101720, 101740, 101770, 101790, 101840, 101910, 101980, 102000, 
    102000, 102000, 102020, 102030, 102060, 102080, 102110, 102130, 102150, 
    102160, 102160, 102150, 102160, 102180, 102210, 102220, 102240, 102280, 
    102270, 102290, 102300, 102310, 102310, 102310, 102300, 102300, 102310, 
    102330, 102340, 102360, 102380, 102390, 102400, 102400, 102390, 102410, 
    102410, 102420, 102430, 102460, 102500, 102550, 102590, 102650, 102690, 
    102720, 102760, 102800, 102830, 102840, 102890, 102940, 102960, 103010, 
    103070, 103100, 103110, 103130, 103180, 103180, 103210, 103220, 103230, 
    103270, 103280, 103310, 103330, 103350, 103370, 103380, 103370, 103380, 
    103370, 103350, 103340, 103330, 103310, 103320, 103340, 103330, 103320, 
    103320, 103320, 103300, 103280, 103300, 103300, 103300, 103290, 103310, 
    103330, 103350, 103360, 103400, 103410, 103410, 103400, 103400, 103400, 
    103420, 103410, 103400, 103400, 103400, 103380, 103370, 103360, 103350, 
    103310, 103320, 103310, 103270, 103250, 103230, 103220, 103200, 103180, 
    103140, 103080, 103030, 103000, 102940, 102900, 102870, 102840, 102810, 
    102760, 102750, 102720, 102680, 102640, 102610, 102600, 102560, 102560, 
    102540, 102520, 102500, 102450, 102440, 102410, 102390, 102350, 102320, 
    102280, 102250, 102210, 102190, 102190, 102170, 102150, 102150, 102140, 
    102130, 102100, 102080, 102080, 102070, 102120, 102150, 102170, 102210, 
    102260, 102300, 102320, 102340, 102370, 102380, 102400, 102400, 102410, 
    102440, 102440, 102440, 102450, 102460, 102440, 102460, 102450, 102440, 
    102420, 102390, 102370, 102360, 102310, 102300, 102310, 102310, 102290, 
    102280, 102280, 102260, 102240, 102230, 102220, 102200, 102210, 102210, 
    102190, 102180, 102180, 102170, 102160, 102150, 102130, 102140, 102130, 
    102110, 102120, 102120, 102140, 102140, 102150, 102160, 102150, 102140, 
    102140, 102140, 102130, 102130, 102130, 102120, 102110, 102110, 102090, 
    102080, 102080, 102060, 102070, 102040, 102070, 102060, 102070, 102070, 
    102090, 102090, 102070, 102080, 102070, 102050, 102030, 102020, 102020, 
    102020, 102000, 101980, 101980, 101980, 101960, 101940, 101910, 101890, 
    101880, 101850, 101840, 101830, 101830, 101830, 101840, 101860, 101870, 
    101880, 101890, 101900, 101920, 101920, 101920, 101920, 101930, 101920, 
    101930, 101940, 101940, 101920, 101940, 101930, 101940, 101920, 101920, 
    101930, 101930, 101920, 101930, 101940, 101940, 101930, 101910, 101900, 
    101880, 101850, 101830, 101810, 101790, 101770, 101750, 101740, 101720, 
    101700, 101680, 101660, 101640, 101660, 101660, 101660, 101670, 101710, 
    101740, 101740, 101760, 101770, 101780, 101770, 101780, 101760, 101770, 
    101780, 101790, 101800, 101820, 101830, 101840, 101830, 101810, 101790, 
    101790, 101780, 101760, 101740, 101740, 101740, 101740, 101740, 101730, 
    101740, 101740, 101720, 101720, 101720, 101730, 101720, 101730, 101730, 
    101730, 101750, 101750, 101750, 101760, 101750, 101750, 101750, 101760, 
    101760, 101760, 101770, 101770, 101790, 101800, 101810, 101820, 101820, 
    101810, 101800, 101790, 101780, 101780, 101790, 101790, 101810, 101830, 
    101830, 101840, 101850, 101870, 101870, 101860, 101840, 101840, 101860, 
    101870, 101900, 101900, 101900, 101900, 101900, 101910, 101880, 101870, 
    101870, 101880, 101880, 101880, 101860, 101880, 101870, 101880, 101870, 
    101850, 101840, 101820, 101850, 101850, 101890, 101880, 101900, 101860, 
    101870, 101870, 101870, 101860, 101850, 101840, 101810, 101780, 101770, 
    101760, 101770, 101740, 101710, 101680, 101650, 101630, 101620, 101620, 
    101610, 101600, 101610, 101620, 101600, 101610, 101620, 101620, 101610, 
    101590, 101560, 101550, 101540, 101520, 101500, 101500, 101500, 101480, 
    101470, 101460, 101420, 101410, 101400, 101380, 101380, 101360, 101340, 
    101370, 101310, 101320, 101320, 101300, 101250, 101240, 101190, 101170, 
    101140, 101110, 101080, 101060, 101030, 101010, 100980, 100930, 100890, 
    100850, 100790, 100740, 100680, 100610, 100590, 100600, 100520, 100500, 
    100410, 100320, 100290, 100250, 100210, 100210, 100200, 100200, 100180, 
    100160, 100160, 100140, 100110, 100080, 100050, 100040, 100020, 99970, 
    99940, 99920, 99890, 99870, 99870, 99850, 99830, 99830, 99820, 99810, 
    99790, 99780, 99780, 99760, 99750, 99760, 99740, 99710, 99700, 99690, 
    99700, 99690, 99700, 99710, 99720, 99730, 99760, 99790, 99810, 99850, 
    99860, 99880, 99880, 99890, 99890, 99880, 99900, 99910, 99920, 99930, 
    99940, 99940, 99940, 99920, 99880, 99850, 99820, 99810, 99800, 99810, 
    99820, 99830, 99870, 99880, 99890, 99910, 99930, 99950, 100000, 100020, 
    100060, 100060, 100100, 100130, 100170, 100200, 100230, 100260, 100280, 
    100280, 100310, 100340, 100380, 100400, 100410, 100440, 100480, 100520, 
    100550, 100570, 100590, 100600, 100620, 100640, 100660, 100690, 100700, 
    100720, 100730, 100760, 100770, 100790, 100800, 100810, 100850, 100850, 
    100860, 100880, 100900, 100910, 100930, 100940, 100950, 100950, 100950, 
    100970, 100970, 100960, 100980, 101000, 101000, 100980, 100980, 100980, 
    100960, 100980, 100980, 100970, 100960, 100960, 100940, 100910, 100910, 
    100890, 100880, 100850, 100820, 100790, 100750, 100730, 100690, 100650, 
    100610, 100540, 100490, 100420, 100360, 100320, 100270, 100220, 100190, 
    100180, 100140, 100130, 100140, 100120, 100120, 100160, 100150, 100170, 
    100230, 100260, 100290, 100340, 100410, 100480, 100520, 100580, 100640, 
    100700, 100770, 100840, 100880, 100970, 101010, 101040, 101110, 101160, 
    101190, 101240, 101290, 101340, 101380, 101430, 101470, 101500, 101520, 
    101530, 101540, 101550, 101570, 101580, 101590, 101620, 101620, 101620, 
    101630, 101630, 101640, 101630, 101620, 101630, 101630, 101650, 101650, 
    101670, 101680, 101700, 101710, 101700, 101700, 101720, 101650, 101710, 
    101750, 101770, 101780, 101800, 101850, 101850, 101850, 101850, 101850, 
    101860, 101880, 101900, 101920, 101930, 101950, 101940, 101950, 101960, 
    101960, 101970, 101730, 101830, 101860, 101920, 101930, 101990, 102000, 
    102000, 102000, 101990, 101980, 101980, 101960, 101930, 101900, 101860, 
    101840, 101830, 101830, 101810, 101800, 101790, 101790, 101760, 101740, 
    101730, 101720, 101710, 101870, 101700, 101700, 101690, 101690, 101680, 
    101680, 101680, 101670, 101660, 101660, 101680, 101690, 101710, 101770, 
    101800, 101820, 101840, 101860, 101880, 101910, 101920, 101960, 101690, 
    101740, 101990, 102030, 102080, 102110, 102150, 102170, 102170, 102180, 
    102160, 102160, 102170, 102190, 102190, 102180, 102160, 102170, 102050, 
    102010, 102060, 102120, 102160, 102190, 102180, 101930, 101850, 101840, 
    101770, 101750, 101670, 101570, 101530, 101480, 101430, 101320, 101260, 
    101190, 101110, 101100, 101060, 101000, 100960, 100930, 100880, 100850, 
    100820, 100810, 101870, 101370, 100770, 100760, 100750, 100760, 100800, 
    100840, 100860, 100870, 100860, 100840, 100810, 100790, 100800, 100830, 
    100870, 100890, 100920, 100960, 100990, 100990, 101000, 101010, 101050, 
    101060, 101060, 101070, 101080, 101060, 101050, 101050, 101000, 101000, 
    100960, 100890, 100870, 100820, 100750, 100720, 100660, 100640, 100590, 
    100570, 100540, 100520, 100500, 100460, 100450, 100440, 100410, 100460, 
    100450, 100420, 100440, 100440, 100400, 100360, 100360, 100350, 100330, 
    100330, 100340, 100330, 100320, 100290, 100280, 100350, 100360, 100360, 
    100380, 100390, 100350, 100420, 100430, 100480, 100510, 100540, 100580, 
    100620, 100620, 100660, 100680, 100690, 100700, 100710, 100760, 100790, 
    100790, 100800, 100810, 100800, 100790, 100790, 100800, 100790, 100760, 
    100720, 100740, 100780, 100760, 100750, 100740, 100740, 100730, 100720, 
    100710, 100700, 100710, 100710, 100730, 100720, 100730, 100770, 100790, 
    100780, 100740, 100740, 100740, 100730, 100710, 100720, 100700, 100740, 
    100730, 100730, 100660, 100670, 100640, 100640, 100630, 100660, 100620, 
    100610, 100610, 100640, 100710, 100640, 100670, 100620, 100630, 100600, 
    100570, 100540, 100500, 100490, 100470, 100450, 100440, 100350 ;

 air_pressure_at_sea_level_qnh = 1007, 1007.1, 1006.7, 1006.7, 1006.8, 
    1006.8, 1006.7, 1006.6, 1007.2, 1007.1, 1007.3, 1007.5, 1007.5, 1007.5, 
    1007.5, 1007.5, 1007.5, 1007.6, 1007.8, 1007.9, 1006.9, 1007, 1006.8, 
    1006.8, 1006.6, 1006.6, 1006.5, 1006.4, 1006.4, 1006.3, 1006.3, 1006.2, 
    1006.6, 1006.6, 1006.5, 1006.5, 1006.5, 1006.4, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 1003, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 1007.6, 1007.6, 1008, 1008, 1008.3, 1008.7, 1009.1, 
    1009.4, 1009.6, 1009.8, 1009.9, 1010.1, 1010.2, 1010.3, 1010.4, 1010.2, 
    1010.2, 1010.3, 1010.6, 1010.5, 1010.6, 1010.7, 1010.7, 1010.5, 1010.4, 
    1010.2, 1010.1, 1009.9, 1010, 1010, 1010, 1010.2, 1010.1, 1010, 1010.2, 
    1010.1, 1010.3, 1010.6, 1010.9, 1011.2, 1011.7, 1012.3, 1012.9, 1013.5, 
    1014.1, 1014.7, 1015.2, 1015.8, 1016.4, 1017, 1017.4, 1017.8, 1018.4, 
    1018.8, 1018.9, 1019.5, 1019.7, 1020, 1020.3, 1020.6, 1020.7, 1020.5, 
    1020.7, 1020.8, _, 1022.3, 1022.6, 1023.1, 1023.4, 1023.7, 1024.1, 
    1024.4, 1024.5, 1024.5, 1024.6, 1025, 1025.2, 1025.5, 1025.9, 1026.3, 
    1026.2, 1026.2, 1026.3, 1026.6, 1026.5, 1026.1, 1025.9, 1025.8, 1025.4, 
    1025.9, 1025.8, 1025.5, 1026.1, 1026, 1025.8, 1025.6, 1025.6, 1025.6, 
    1024.7, 1024.5, 1024.3, 1024.1, 1024.1, 1024.1, 1024.2, 1024.3, 1024.4, 
    1024.1, 1024.2, 1023.8, 1023.7, 1023.7, 1024, 1024.4, 1024.7, 1025.1, 
    1025.3, 1025.5, 1025.7, 1025.9, 1025.7, 1025.9, 1026.1, 1026.5, 1026.6, 
    1027, 1027.3, 1027.8, 1028.3, 1028.6, 1028.8, 1029, 1029.3, 1029.7, 
    1029.5, 1030, 1030.3, 1030.5, 1030.9, 1031.6, 1031.8, 1032.3, 1032.5, 
    1032.7, 1014.8, 1033.1, 1033.6, 1033.6, 1033.9, 1034.1, 1034.5, 1034.7, 
    1034.8, 1035.1, 1034.9, 1035, 1035.1, 1035.2, 1035.1, 1035.1, 1034.9, 
    1035, 1034.9, 1034.7, 1034.6, 1034.3, 1034.1, 1034.3, 1034.4, 1034.1, 
    1034, 1033.9, 1034, 1034.2, 1034.1, 1034, 1034.2, 1034.2, 1034, 1034, 
    1033.9, 1033.6, 1033.6, 1033.7, 1033.6, 1033.7, 1033.8, 1034.1, 1034.4, 
    1034.4, 1034.4, 1034.4, 1034.5, 1034.5, 1034.6, 1034.4, 1034.5, 1034.6, 
    1035, 1035.1, 1035.2, 1034.9, 1035.1, 1035.3, 1035.3, 1035.4, 1035.1, 
    1035.1, 1035, 1034.8, 1035, 1035, 1035, 1034.9, 1034.9, 1034.8, 1034.8, 
    1034.8, 1034.8, 1035, 1035.2, 1035.2, 1035.4, 1035.5, 1035.9, 1035.8, 
    1035.8, 1036.1, 1036.1, 1036.3, 1036.4, 1036.5, 1036.5, 1036.4, 1036.9, 
    1037.2, 1037.3, 1037.4, 1037.5, 1037.4, 1037, 1036.9, 1036.4, 1036, 
    1035.9, 1035.7, 1035.5, 1035.1, 1034.8, 1034.4, 1033.8, 1033.4, 1033.1, 
    1032.7, 1032.3, 1031.9, 1031.2, 1030.8, 1030.5, 1030.3, 1029.9, 1029.7, 
    1029.2, 1028.7, 1028.1, 1027.7, 1027.2, 1026.7, 1026.2, 1025.8, 1025.3, 
    1025.1, 1024.5, 1024.3, 1023.8, 1023.7, 1023.6, 1023.5, 1023.2, 1023.2, 
    1023.5, 1023.7, 1023.9, 1024.1, 1024.6, 1024.7, 1024.7, 1024.8, 1024.9, 
    1024.9, 1024.7, 1024.6, 1024.6, 1024.7, 1024.6, 1024.8, 1024.9, 1024.8, 
    1024.8, 1024.7, 1024.5, 1024.6, 1024.6, 1024.3, 1024.3, 1024, 1024.1, 
    1024, 1024.1, 1024, 1023.9, 1023.7, 1023.4, 1023.4, 1023.4, 1023.2, 
    1023.2, 1023.2, 1023.3, 1023.3, 1023.2, 1023, 1022.9, 1022.7, 1022.5, 
    1022.2, 1022, 1021.4, 1021.3, 1021, 1021.1, 1021.2, 1021.2, 1020.8, 
    1020.5, 1020.3, 1020.1, 1019.8, 1019.5, 1019.4, 1019.2, 1019, 1018.8, 
    1018.5, 1018.4, 1018.2, 1017.8, 1017.4, 1017, 1016.9, 1016.8, 1016.4, 
    1016.1, 1016.1, 1016.1, 1016, 1015.8, 1015.6, 1015.6, 1015.2, 1015, 
    1014.9, 1014.5, 1014.4, 1014.4, 1014, 1013.7, 1013.3, 1013.1, 1012.6, 
    1012, 1011.5, 1011.3, 1011, 1010.7, 1010.4, 1010.2, 1010.1, 1009.9, 
    1010.1, 1010, 1009.8, 1009.7, 1009.6, 1009.5, 1009.4, 1009.4, 1009.2, 
    1008.9, 1009.2, 1009.7, 1009.5, 1010.1, 1010.3, 1010.7, 1011.2, 1011.8, 
    1012.3, 1012.9, 1013.4, 1013.7, 1014.5, 1015.4, 1016.1, 1016.6, 1017.1, 
    1017.4, 1017.7, 1018.2, 1018.9, 1019.6, 1020.2, 1020.7, 1021.4, 1022.3, 
    1023, 1023.5, 1024.1, 1024.7, 1025.2, 1025.8, 1026.5, 1027.1, 1027.7, 
    1028.3, 1029, 1029.7, 1030.4, 1030.9, 1031.3, 1031.6, 1031.8, 1032.1, 
    1032.1, 1031.6, 1031.5, 1031.3, 1030.7, 1030.5, 1030.2, 1029.6, 1029, 
    1027.9, 1026.7, 1025.9, 1025, 1023.4, 1022.2, 1021.2, 1020.2, 1019.7, 
    1019.4, 1019.3, 1019.2, 1019.2, 1018.9, 1019.1, 1019.1, 1019.2, 1019.2, 
    1019, 1019.2, 1019.2, 1019.5, 1019.8, 1020.2, 1020.5, 1020.9, 1021.2, 
    1021.7, 1021.8, 1021.9, 1022.1, 1022.5, 1022.4, 1022.4, 1022.6, 1022.8, 
    1022.7, 1022.8, 1022.8, 1023.1, 1023.4, 1023.7, 1023.5, 1023.9, 1024.2, 
    1024.8, 1025.3, 1025.7, 1025.9, 1026, 1026.3, 1026.6, 1026.8, 1027.2, 
    1027.4, 1027.7, 1028.2, 1028.9, 1029.4, 1029.6, 1029.9, 1030.3, 1030.7, 
    1030.8, 1031, 1031.4, 1031.7, 1031.9, 1032, 1032.3, 1032.2, 1032, 1031.8, 
    1031.3, 1030.9, 1030.5, 1030.1, 1029.5, 1029.1, 1028.8, 1028.3, 1027.9, 
    1027.5, 1027.3, 1026.7, 1026.2, 1025.8, 1025.2, 1024.7, 1024.3, 1023.9, 
    1023.4, 1023.1, 1023.1, 1022.7, 1022.5, 1022.1, 1021.8, 1021.4, 1021.2, 
    1021.1, 1020.7, 1020.5, 1020.4, 1020.6, 1020.6, 1020.3, 1020.2, 1020.1, 
    1020, 1020, 1019.9, 1019.6, 1019.6, 1019.4, 1019.8, 1020.2, 1020.3, 
    1020.2, 1020.4, 1020.4, 1020.8, 1020.9, 1021, 1021.2, 1021.4, 1021.5, 
    1021.8, 1022.1, 1022.2, 1022.2, 1021.9, 1021.1, 1020.7, 1020.1, 1019.3, 
    1018, 1016.8, 1015.6, 1014.4, 1013.1, 1012.3, 1011.4, 1010.5, 1009.7, 
    1009, 1008.5, 1007.7, 1006.5, 1005.7, 1005.1, 1005, 1005.2, 1005.3, 
    1005.5, 1005.5, 1005.7, 1005.7, 1005.9, 1005.9, 1006, 1006, 1006.1, 
    1005.9, 1005.8, 1005.5, 1005.3, 1005, 1004.8, 1004.6, 1004.7, 1004.5, 
    1004.3, 1004.7, 1005.2, 1006, 1007.1, 1008, 1008.9, 1010, 1011.1, 1012.4, 
    1013.6, 1014.6, 1015.5, 1016.5, 1017.1, 1018.2, 1019, 1019.7, 1020.5, 
    1020.7, 1021.5, 1022.2, 1022.7, 1023.1, 1023.6, 1024.2, 1024.7, 1025.3, 
    1026.1, 1026.8, 1027.4, 1028, 1028.5, 1029, 1029.5, 1030.1, 1030.5, 
    1030.9, 1031.2, 1031.5, 1032, 1032, 1032.1, 1032.2, 1031.9, 1031.7, 
    1031.5, 1031, 1030.2, 1029.5, 1028.5, 1027.4, 1026, 1024.6, 1023.5, 
    1022.5, 1021, 1019.4, 1018.3, 1017.5, 1016.6, 1016.5, 1017.1, 1018.1, 
    1019.3, 1019.7, 1020.5, 1021.5, 1021.8, 1023, 1023.5, 1024.3, 1025.1, 
    1025.2, 1025.8, 1026.5, 1027.2, 1028, 1028.5, 1028.7, 1029, 1029.2, 
    1029.4, 1029.9, 1030, 1030.2, 1030.4, 1030.4, 1030.3, 1030.4, 1030.4, 
    1030.3, 1030, 1029.8, 1029.6, 1029.2, 1028.9, 1028.6, 1028.3, 1028, 
    1027.7, 1027.4, 1027, 1026.1, 1025, 1023.8, 1022.9, 1021.5, 1020.3, 
    1018.5, 1017.3, 1016, 1014.9, 1014.1, 1012.8, 1011.9, 1010.9, 1010, 
    1009.8, 1009.4, 1009, 1008.3, 1007.9, 1007.3, 1007.3, 1007.3, 1006.7, 
    1006.6, 1006.1, 1005, 1004.1, 1003.9, 1003.8, 1003.9, 1004.5, 1004.6, 
    1005.2, 1006, 1006, 1005.9, 1006.9, 1008.7, 1009.7, 1010.8, 1012, 1013.1, 
    1014.3, 1015.4, 1016.4, 1017.8, 1019.2, 1020.2, 1021.1, 1022, 1022.7, 
    1023.3, 1023.8, 1024.3, 1024.2, 1024.6, 1025, 1024.8, 1024.8, 1024.5, 
    1024.1, 1023.4, 1022.7, 1022.1, 1021.3, 1020.5, 1019.7, 1019, 1018.4, 
    1017.8, 1017, 1016.5, 1015.5, 1014.8, 1014.1, 1013.2, 1012.6, 1011.9, 
    1010.8, 1010.1, 1009.5, 1008.8, 1007.8, 1007.2, 1006.5, 1006.2, 1005.7, 
    1005.3, 1004.8, 1004.4, 1003.7, 1003.3, 1002.8, 1002.3, 1001.5, 1000.9, 
    1000.1, 999.4, 998.8, 998.6, 998.4, 998.3, 998.3, 998.4, 998.6, 998.9, 
    998.8, 998.9, 998.9, 998.8, 998.9, 998.8, 998.8, 998.5, 998.4, 998.6, 
    998.6, 998.5, 998.3, 998, 997.5, 996.9, 996.4, 995.4, 995, 995, 994.6, 
    993.8, 992.9, 992.7, 992.5, 992.2, 991.7, 991, 990.6, 990.3, 990, 989.6, 
    989.1, 988.6, 988.3, 988.2, 987.9, 987.6, 987, 986.6, 986.4, 986.5, 
    986.5, 986.6, 986.7, 986.9, 987.2, 987.7, 988.2, 988.4, 988.6, 988.8, 
    989.3, 989.8, 990.4, 991, 991.3, 991.7, 992.4, 993.3, 993.9, 994.5, 995, 
    995.7, 996.6, 997.4, 998.3, 999, 999.9, 1000.4, 1001, 1001.6, 1002.2, 
    1002.8, 1003.3, 1003.5, 1004.1, 1004.4, 1004.5, 1004.6, 1004.8, 1005.1, 
    1005.1, 1005.3, 1005.2, 1005.1, 1005, 1004.4, 1004, 1003.1, 1001.9, 
    1000.9, 1000.3, 999.9, 999.6, 999.4, 999.1, 998.9, 998.8, 999.2, 999.7, 
    1000.2, 1000.4, 1000.4, 1000.6, 1001.4, 1001.9, 1002.8, 1003.6, 1004.2, 
    1004.5, 1004.8, 1005.3, 1005.2, 1005.6, 1005.9, 1006.1, 1006.4, 1006.5, 
    1006.9, 1007.2, 1007.1, 1007, 1006.8, 1006.1, 1005.1, 1004.3, 1003.8, 
    1003.5, 1003.1, 1003, 1003.2, 1003.1, 1003.1, 1003, 1002.3, 1001.8, 
    1001.2, 1001.1, 1001.1, 1001.1, 1000.9, 1000.8, 1000.6, 1000.7, 1000.5, 
    1000.2, 999.6, 999.5, 998.6, 998.1, 997.8, 997.4, 997.1, 996.7, 996.3, 
    996.2, 995.6, 995.3, 995.5, 995.1, 994.9, 995, 994.9, 994.6, 994.3, 
    993.5, 994.5, 994, 994, 994.4, 994.6, 994.7, 994.6, 994.9, 995.3, 995.3, 
    995.7, 995.9, 996.2, 996, 995.7, 995.5, 995.7, 995.6, 995.6, 995.2, 
    995.4, 995.3, 995.3, 995.2, 995.5, 995.5, 995.4, 995.3, 995, 994.9, 
    994.7, 994.2, 994.4, 994.6, 994.8, 995, 994.9, 995.2, 995, 994.9, 994.8, 
    994.4, 993.9, 993.5, 993, 992.5, 992.4, 992.1, 992, 991.6, 991.3, 990.9, 
    990.6, 990.4, 990.4, 990.2, 990, 990.2, 990.5, 990.6, 991.1, 991.8, 
    992.2, 992.5, 993, 993.5, 994.1, 994.6, 995.2, 995.5, 996.1, 996.6, 
    997.1, 997.7, 998.6, 999.2, 999.9, 1000.5, 1001.2, 1001.7, 1002.5, 
    1003.1, 1003.7, 1004.5, 1005.3, 1005.9, 1006.6, 1007.1, 1007.6, 1008.1, 
    1008.6, 1009.2, 1009.8, 1010.1, 1010.7, 1011.4, 1012, 1012.5, 1012.9, 
    1013.3, 1013.8, 1014.2, 1014.7, 1014.9, 1015.2, 1015.3, 1015.6, 1015.8, 
    1015.8, 1016, 1016.2, 1016.2, 1016, 1015.8, 1015.3, 1014.9, 1014.3, 
    1013.6, 1012.9, 1012, 1010.7, 1009.5, 1008.3, 1007.2, 1005.9, 1004.3, 
    1002.1, 1000.3, 998.2, 997.2, 996.6, 996.1, 995.7, 995.3, 995, 994.8, 
    994.8, 994.2, 993.6, 993.1, 992.6, 992, 991.7, 991.3, 991.1, 990.8, 991, 
    991.2, 991.7, 992, 992.5, 992.7, 992.8, 993.2, 993.4, 993.5, 993.8, 
    993.8, 993.5, 993.3, 993.2, 993.9, 994.4, 995.5, 996.3, 996.7, 997, 
    997.9, 998.3, 999, 999.1, 999.3, 999.3, 999.6, 999.9, 1000.1, 1000.4, 
    1000.7, 1001.3, 1001.7, 1002.1, 1002.8, 1003.3, 1003.8, 1004.5, 1005.1, 
    1005.8, 1006.8, 1007.5, 1008, 1008.8, 1009.7, 1010.1, 1010.7, 1011.7, 
    1012, 1012.5, 1012.9, 1013.2, 1013.2, 1013.9, 1014.3, 1014.7, 1015, 
    1015.3, 1015.4, 1015.3, 1015.3, 1015.2, 1014.6, 1014.3, 1013.9, 1013.5, 
    1012.7, 1012.6, 1012.1, 1011.9, 1012.2, 1012, 1011.8, 1011.3, 1011.8, 
    1011.9, 1011.8, 1011.7, 1011.7, 1011.2, 1010.6, 1010, 1009.1, 1008.1, 
    1007.1, 1005.9, 1004.9, 1004.3, 1003.1, 1002.5, 1002.1, 1000.9, 999.9, 
    998.7, 997.5, 995.9, 994.1, 993.2, 993, 993, 993.1, 992.9, 992.9, 993.5, 
    994, 994.9, 995.7, 996.4, 997.2, 997.4, 998.1, 998.5, 998.7, 999.4, 
    1000.2, 1000.7, 1001.5, 1002.8, 1003.8, 1004.9, 1005.6, 1006.8, 1007.6, 
    1008.8, 1009.8, 1010.5, 1011.3, 1012.1, 1012.9, 1013.7, 1014.3, 1014.8, 
    1015.2, 1015.7, 1015.9, 1016.2, 1016.4, 1016.7, 1016.8, 1017.1, 1017.3, 
    1017.6, 1017.8, 1018, 1018.1, 1018.2, 1018.4, 1018.5, 1018.9, 1019, 1019, 
    1019.1, 1019.3, 1019.5, 1019.8, 1020.2, 1020.3, 1020.7, 1020.7, 1021, 
    1021.2, 1021.1, 1020.9, 1021.1, 1021.3, 1021.4, 1021.5, 1022, 1022.1, 
    1022.3, 1022.1, 1022.2, 1022.2, 1022.2, 1022.5, 1022.4, 1022.8, 1023.3, 
    1023.5, 1023.7, 1023.8, 1024.1, 1024.2, 1024.3, 1024.2, 1024.3, 1024.3, 
    1024, 1023.8, 1023.7, 1023.5, 1023.4, 1023.2, 1023.1, 1022.8, 1022.5, 
    1022, 1021.7, 1021.1, 1020.7, 1020.5, 1020.3, 1020, 1019.6, 1019.2, 
    1018.7, 1018.2, 1017.3, 1016.7, 1016.2, 1015.5, 1014.5, 1013.6, 1012.8, 
    1011.8, 1010.8, 1009.4, 1008.7, 1007.7, 1006.9, 1005.8, 1004.9, 1004.2, 
    1003.7, 1003.1, 1002.8, 1002.8, 1003, 1003.1, 1003.1, 1003.1, 1003.1, 
    1003.1, 1003, 1003.1, 1003.3, 1003.4, 1003.6, 1003.5, 1003.6, 1003.6, 
    1003.4, 1003.1, 1002.9, 1002.6, 1002.2, 1002.2, 1002.2, 1002.1, 1002.2, 
    1002.1, 1002.2, 1002.1, 1001.8, 1001.4, 1001, 1001.2, 1001, 1001.1, 
    1000.9, 1000.6, 1000.5, 999.9, 999.8, 1000.2, 1000.4, 1001.3, 1002, 
    1002.9, 1003.6, 1004.1, 1004.6, 1005.1, 1005.7, 1006.2, 1006.7, 1007.4, 
    1007.7, 1008.2, 1009, 1009.5, 1010.1, 1010.7, 1011.2, 1011.9, 1012.6, 
    1013.4, 1014.1, 1014.4, 1014.5, 1014.9, 1015, 1015.3, 1015.5, 1015.7, 
    1015.7, 1016, 1016.3, 1016.3, 1016.3, 1016.3, 1016, 1015.9, 1015.7, 
    1015.6, 1015.1, 1014.5, 1014, 1013.5, 1013.2, 1012.5, 1011.7, 1011, 
    1010.3, 1009.4, 1008.3, 1007.5, 1006.6, 1005.6, 1004.5, 1003.3, 1002.5, 
    1001.3, 999.8, 999.2, 998.2, 996.9, 996.1, 995.6, 995.2, 994.9, 994.7, 
    995, 995.3, 995.8, 996.1, 996.7, 997.3, 997.9, 998.6, 999.4, 1000.6, 
    1001.9, 1002.8, 1003.6, 1004.9, 1006, 1007, 1007.9, 1008.9, 1010.4, 
    1011.3, 1011.6, 1012.2, 1012.9, 1013.5, 1014, 1014.7, 1015.1, 1015, 
    1015.1, 1015.3, 1015.4, 1015.6, 1015.2, 1015.2, 1015, 1014.9, 1014.9, 
    1014.8, 1014.8, 1014.7, 1014.4, 1014.3, 1014.1, 1014.1, 1013.9, 1014, 
    1014.6, 1014.9, 1015.3, 1015.6, 1015.8, 1016, 1016.3, 1016.9, 1017.2, 
    1017.6, 1017.3, 1017.4, 1017.6, 1017.8, 1018.4, 1019, 1019.8, 1020.3, 
    1020.9, 1021.2, 1021.2, 1021.4, 1021.4, 1021.5, 1021.8, 1022.1, 1022.1, 
    1022.2, 1022.3, 1022.4, 1022.4, 1022.1, 1021.8, 1021.7, 1021.8, 1021.5, 
    1021, 1020.8, 1020.5, 1019.9, 1019.4, 1019.2, 1018.7, 1017.9, 1017.7, 
    1017, 1016.2, 1015.7, 1015.2, 1014.5, 1014, 1013.7, 1013.4, 1013.1, 
    1012.9, 1012.6, 1012.3, 1012, 1011.9, 1011.9, 1011.9, 1011.8, 1011.8, 
    1011.6, 1011.4, 1011.1, 1011, 1010.8, 1010.4, 1010.3, 1010.2, 1010.1, 
    1010, 1009.8, 1009.7, 1009.4, 1009, 1009, 1009, 1008.8, 1008.8, 1009.1, 
    1009.2, 1009.1, 1008.9, 1008.8, 1008.8, 1008.8, 1008.7, 1008.7, 1008.6, 
    1008.5, 1008.6, 1008.8, 1008.6, 1008.4, 1008.2, 1008.1, 1008, 1007.9, 
    1007.9, 1007.7, 1007.6, 1007.5, 1007.6, 1007.3, 1007.1, 1006.9, 1006.8, 
    1006.9, 1007, 1006.9, 1007, 1007.1, 1007.1, 1007.1, 1006.8, 1006.6, 
    1006.5, 1006.4, 1006.3, 1006.2, 1006.3, 1006.3, 1006.3, 1006.3, 1006.1, 
    1006, 1006.1, 1006.1, 1006, 1005.9, 1006, 1006, 1006, 1006, 1006.2, 
    1006.2, 1006.3, 1006.2, 1006.2, 1006.2, 1006.2, 1006.1, 1005.9, 1005.8, 
    1005.8, 1005.8, 1005.9, 1005.8, 1005.8, 1005.8, 1005.7, 1005.7, 1005.7, 
    1005.7, 1005.7, 1005.7, 1006, 1006.3, 1006.4, 1006.5, 1006.4, 1006.2, 
    1006.4, 1006.3, 1006, 1006.1, 1006.1, 1006, 1005.9, 1005.7, 1005.4, 
    1005.3, 1005.2, 1005, 1004.8, 1004.5, 1004.1, 1003.7, 1003.4, 1003.3, 
    1003.2, 1003.1, 1003, 1002.8, 1002.4, 1002.2, 1002.1, 1001.9, 1001.8, 
    1001.6, 1001.6, 1001.6, 1001.7, 1001.8, 1001.8, 1001.7, 1001.7, 1001.7, 
    1001.7, 1002, 1001.9, 1001.5, 1000.9, 1000.7, 1000.8, 1000.9, 1001, 1001, 
    1001.1, 1001.1, 1001.3, 1001.7, 1001.7, 1001.7, 1001.8, 1002.1, 1002.3, 
    1002.8, 1003.1, 1003.3, 1003.4, 1003.2, 1003.3, 1003.5, 1003.5, 1003.2, 
    1003.1, 1003.4, 1003.5, 1003.8, 1004.1, 1004.4, 1004.8, 1004.7, 1005, 
    1004.9, 1004.7, 1004.8, 1004.6, 1004.5, 1004.5, 1004.5, 1004.5, 1004.5, 
    1004.5, 1004.7, 1004.7, 1004.6, 1004.4, 1004.5, 1004.4, 1004.4, 1004.1, 
    1004.1, 1003.6, 1003.4, 1003.3, 1003.1, 1002.8, 1002.7, 1002.6, 1002.5, 
    1002.5, 1002.1, 1002.2, 1002.2, 1002.2, 1002, 1001.8, 1001.9, 1002.1, 
    1002.1, 1001.7, 1001.8, 1001.8, 1001.9, 1002.2, 1002.4, 1002.5, 1002.6, 
    1002.8, 1002.7, 1002.9, 1003, 1003, 1002.8, 1003, 1002.9, 1003, 1003.2, 
    1003.4, 1003.3, 1003.2, 1003.2, 1003.1, 1003, 1002.8, 1002.7, 1002.8, 
    1002.7, 1002.7, 1002.5, 1002.4, 1002.4, 1002.2, 1002.1, 1002.2, 1002.2, 
    1002.2, 1002.1, 1002.2, 1002.3, 1002.3, 1002.6, 1003.1, 1003.5, 1003.9, 
    1004.1, 1004.5, 1005, 1005.5, 1005.8, 1006.2, 1006.7, 1007.2, 1007.8, 
    1008.2, 1008.5, 1008.9, 1009.2, 1009.5, 1009.9, 1010.6, 1011.1, 1011.6, 
    1012, 1012.5, 1013, 1013.5, 1013.6, 1014, 1014.3, 1014.6, 1015, 1015.4, 
    1015.6, 1015.8, 1015.8, 1016.2, 1016.2, 1016.4, 1016.2, 1016.2, 1015.9, 
    1015.8, 1015.9, 1015.8, 1015.9, 1015.8, 1015.6, 1015.5, 1015.5, 1015.3, 
    1015.2, 1015, 1014.9, 1014.7, 1014.4, 1014.2, 1014, 1013.8, 1013.9, 
    1013.9, 1013.9, 1013.9, 1014, 1014, 1014.1, 1014.1, 1014.2, 1014.1, 
    1013.9, 1013.8, 1013.5, 1013.4, 1013.4, 1013.4, 1013.6, 1013.7, 1013.7, 
    1013.5, 1013.3, 1012.9, 1012.9, 1013, 1012.4, 1012.5, 1012.6, 1012.3, 
    1012.6, 1012.5, 1012.4, 1012.3, 1012.2, 1012, 1012, 1011.9, 1011.8, 
    1011.8, 1011.8, 1011.6, 1011.5, 1011.5, 1011.3, 1011.1, 1010.8, 1010.4, 
    1010.1, 1009.9, 1010, 1010, 1009.9, 1009.7, 1009.3, 1009.2, 1009.2, 
    1009.4, 1009.8, 1010.3, 1010.8, 1011, 1011.5, 1011.9, 1012.5, 1012.9, 
    1013.4, 1013.8, 1014.6, 1015.3, 1015.8, 1016.2, 1016.4, 1016.3, 1016.5, 
    1016.5, 1016.3, 1016.6, 1015.9, 1015.3, 1014.4, 1013.4, 1012.1, 1011.2, 
    1010.9, 1011.3, 1011.6, 1011.7, 1012.6, 1013.5, 1014.3, 1015, 1016, 
    1016.8, 1017.4, 1018.1, 1018.7, 1019.1, 1019.5, 1019.9, 1020.2, 1020.5, 
    1020.5, 1020.7, 1020.6, 1020.5, 1020.6, 1020.6, 1020.6, 1020.4, 1020.6, 
    1020.7, 1021.1, 1021.4, 1021.5, 1021.8, 1022.2, 1023, 1023.4, 1023.6, 
    1023.6, 1023.8, 1024.3, 1024.7, 1025.4, 1025.8, 1026, 1026.4, 1026.4, 
    1026.5, 1026.4, 1026.5, 1026.4, 1026.4, 1026.4, 1026.1, 1026.1, 1025.8, 
    1025.2, 1024.7, 1024.1, 1023.4, 1023.2, 1022.9, 1022.6, 1022.6, 1022.4, 
    1022.1, 1022.4, 1022.5, 1022.4, 1022.4, 1022, 1021.7, 1021.4, 1021, 
    1020.5, 1020.1, 1019.6, 1018.9, 1018.4, 1017.9, 1017.5, 1016.5, 1015.7, 
    1015, 1014.1, 1013.4, 1012.7, 1012, 1011.6, 1011.2, 1010.9, 1010.4, 
    1009.9, 1009.4, 1009, 1008.7, 1008.4, 1008, 1007.9, 1007.9, 1007.8, 
    1008.1, 1008.4, 1008.9, 1009.2, 1009.4, 1009.3, 1009.4, 1009.4, 1009.5, 
    1009.5, 1010.1, 1010.6, 1011.4, 1012.5, 1013.5, 1014.9, 1015.6, 1016.4, 
    1017, 1017.7, 1018.3, 1018.5, 1019, 1019.4, 1020.2, 1020.7, 1021, 1021.2, 
    1021.1, 1021.1, 1021.4, 1021.8, 1022, 1022.1, 1022.1, 1021.9, 1022.1, 
    1022.3, 1022.6, 1022.7, 1022.5, 1022.1, 1021.5, 1020.5, 1019.9, 1019.7, 
    1019.8, 1019.8, 1019.6, 1019.3, 1019.1, 1018.7, 1018.1, 1017.7, 1017.5, 
    1017.4, 1017.1, 1016.8, 1016.7, 1016.6, 1016.6, 1016.5, 1016.5, 1016.2, 
    1016, 1016, 1015.8, 1015.8, 1016.1, 1016.3, 1016.4, 1016.8, 1017.4, 
    1017.7, 1018.3, 1018.8, 1019.2, 1019.6, 1019.8, 1019.8, 1020.2, 1020.6, 
    1021.1, 1021.7, 1022.3, 1022.8, 1023.3, 1023.7, 1023.8, 1024, 1024.3, 
    1024.3, 1024.4, 1024.3, 1024.1, 1024, 1023.8, 1023.5, 1023.3, 1023.1, 
    1022.5, 1022.6, 1022.4, 1022.2, 1022.4, 1022.4, 1022.6, 1022.8, 1023, 
    1023.3, 1023.4, 1023.3, 1023.3, 1023.3, 1023.3, 1022.8, 1022.6, 1022.1, 
    1022, 1021.9, 1021.5, 1021.2, 1020.7, 1020.4, 1019.7, 1018.9, 1018.6, 
    1018.1, 1017.4, 1016.6, 1015.7, 1014.9, 1014.5, 1013.8, 1013.2, 1012.5, 
    1012, 1011.8, 1011.8, 1012.2, 1012.7, 1013.5, 1014.3, 1015.1, 1015.9, 
    1016.9, 1017.6, 1018.4, 1019.2, 1019.6, 1021.1, 1020.7, 1021.1, 1021.5, 
    1022.3, 1022.9, 1023.6, 1024, 1024.5, 1025, 1025.3, 1025.7, 1026.1, 
    1026.5, 1026.7, 1026.7, 1027, 1027.2, 1027.2, 1027, 1027, 1026.4, 1025.6, 
    1024.8, 1024.5, 1024.4, 1023.8, 1022.9, 1021.9, 1020.9, 1020, 1019.2, 
    1018.8, 1018.4, 1018.2, 1018.4, 1018.1, 1018, 1018.2, 1018.3, 1018.6, 
    1018.8, 1019, 1019.2, 1019.7, 1019.9, 1020, 1020.5, 1020.9, 1021, 1021.2, 
    1021.3, 1021.5, 1021.5, 1021.5, 1021.5, 1021.7, 1021.8, 1021.7, 1021.3, 
    1020.9, 1020.8, 1020.5, 1020.1, 1019.4, 1019.1, 1019, 1019, 1018.5, 
    1018.3, 1018, 1018, 1018, 1017.8, 1017.9, 1018, 1018.1, 1018.4, 1018.8, 
    1019.4, 1019.7, 1020.1, 1020.4, 1020.6, 1020.7, 1020.7, 1020.7, 1020.5, 
    1020.3, 1020.2, 1019.9, 1019.4, 1019.1, 1018.5, 1018, 1017.2, 1016.3, 
    1015.4, 1014.4, 1013.2, 1012.2, 1011.1, 1009.9, 1009.2, 1009, 1008.2, 
    1007.4, 1006.7, 1006.5, 1006.3, 1006.4, 1006.5, 1006.3, 1006.3, 1006.6, 
    1007, 1007.9, 1008.6, 1009.2, 1009.7, 1010, 1010.7, 1011.5, 1012.5, 
    1013.4, 1014.2, 1015.3, 1016.2, 1017.1, 1018, 1018.8, 1019.5, 1020.4, 
    1020.9, 1021.4, 1022.1, 1022.2, 1022.5, 1022.7, 1022.8, 1022.8, 1022.6, 
    1022.5, 1022.1, 1021.3, 1020.6, 1020, 1019.2, 1019, 1018.6, 1018.2, 
    1018.2, 1018.5, 1018.3, 1018.3, 1018.2, 1018, 1018.2, 1018.2, 1018.5, 
    1018.7, 1019.1, 1019.6, 1019.9, 1020.2, 1020.2, 1020.4, 1020.2, 1020.2, 
    1020.2, 1020.4, 1020.3, 1020.2, 1020.3, 1020.5, 1020.8, 1021.2, 1021.1, 
    1021.2, 1021.2, 1021.3, 1021.5, 1021.4, 1021.1, 1020.8, 1020.6, 1020.7, 
    1020.7, 1020.3, 1020.1, 1020.1, 1019.9, 1019.6, 1019.4, 1019.1, 1018.9, 
    1018.7, 1018.7, 1018.4, 1018.4, 1018.2, 1018, 1017.7, 1018, 1017.7, 
    1017.5, 1017.5, 1017.2, 1016.7, 1016.3, 1015.9, 1015.9, 1015.8, 1015.6, 
    1015.4, 1015.1, 1015, 1014.9, 1014.8, 1014.8, 1014.8, 1014.7, 1014.8, 
    1015.2, 1015.4, 1015.5, 1015.8, 1015.8, 1015.7, 1015.8, 1015.9, 1016, 
    1016.1, 1016.2, 1016.4, 1016.6, 1016.7, 1017, 1017.1, 1017, 1017, 1017.2, 
    1017.2, 1017, 1016.8, 1016.7, 1016.8, 1017, 1017.3, 1017.4, 1017.7, 
    1017.9, 1018.4, 1018.5, 1018.8, 1018.9, 1019.2, 1019.4, 1019.4, 1019.7, 
    1019.7, 1019.6, 1019.6, 1019.3, 1019.1, 1018.9, 1018.8, 1018.6, 1018.7, 
    1018.7, 1019.1, 1019.3, 1019.6, 1019.6, 1019.6, 1019.6, 1019.6, 1019.7, 
    1019.7, 1019.7, 1019.5, 1019.3, 1019.1, 1018.6, 1018.3, 1018.1, 1018.1, 
    1018.3, 1017.8, 1018.6, 1019, 1020.4, 1021.4, 1021.2, 1021.9, 1022.4, 
    1023.3, 1023.3, 1023.5, 1024.2, 1025.1, 1025.8, 1026.2, 1026.6, 1027.4, 
    1028.1, 1028.3, 1028.7, 1029.3, 1029.2, 1029.5, 1029.2, 1029.6, 1029.6, 
    1029.1, 1028.8, 1028.5, 1028.5, 1028.7, 1029, 1029.1, 1028.9, 1028.6, 
    1028.3, 1028, 1027.8, 1027.5, 1027.4, 1027.2, 1027, 1026.7, 1026.7, 
    1026.5, 1026.2, 1025.7, 1025.4, 1025, 1024.7, 1024.6, 1024.4, 1024.2, 
    1024.4, 1024.6, 1024.7, 1024.7, 1025, 1025.4, 1025.5, 1025.8, 1025.9, 
    1026.4, 1026.6, 1027, 1027.4, 1027.9, 1028.2, 1028.5, 1029.1, 1029.5, 
    1029.5, 1029.9, 1030.1, 1030.3, 1030.4, 1030.5, 1030.8, 1030.8, 1031, 
    1031.2, 1031.1, 1030.9, 1030.6, 1030.2, 1029.6, 1029.3, 1028.6, 1028, 
    1027.6, 1027.2, 1026.9, 1026.4, 1026.2, 1026.2, 1025.9, 1025.8, 1025.5, 
    1025.2, 1024.8, 1024.7, 1024.1, 1023.9, 1024, 1023.7, 1023.3, 1023.6, 
    1023.3, 1023.2, 1022.7, 1022.5, 1022.5, 1023, 1023, 1023.1, 1022.9, 
    1022.6, 1022.3, 1022.2, 1022.1, 1021.9, 1021.5, 1021, 1020.9, 1020.6, 
    1020.8, 1021, 1021, 1020.9, 1021.2, 1021.9, 1022.5, 1023, 1023.5, 1023.8, 
    1024, 1024, 1024.2, 1024.5, 1024.9, 1025, 1025.1, 1025.2, 1025.4, 1025.5, 
    1025.6, 1025.7, 1025.7, 1025.8, 1027.4, 1027.4, 1027.4, 1026, 1026.2, 
    1026.2, 1026, 1025.8, 1025.5, 1025.2, 1025.2, 1024.9, 1024.2, 1024.1, 
    1023.6, 1023.6, 1023.2, 1022.5, 1022.4, 1022.6, 1022.9, 1022.5, 1022.4, 
    1022.2, 1022.2, 1022.3, 1022.3, 1022.7, 1022.7, 1022.8, 1022.5, 1022.3, 
    1022.3, 1022.3, 1021.9, 1021.9, 1021.4, 1021, 1020.9, 1020.7, 1020.3, 
    1019.8, 1019.4, 1019, 1018.5, 1018, 1017.3, 1016.7, 1016.2, 1015.8, 
    1015.3, 1014.8, 1014.5, 1014, 1013.4, 1012.9, 1012.5, 1012.2, 1011.6, 
    1011.3, 1010.7, 1010.5, 1010.3, 1010, 1009.6, 1009.2, 1008.8, 1008.5, 
    1008.1, 1007.6, 1007.1, 1006.7, 1006.2, 1006, 1005.7, 1005.2, 1004.7, 
    1004.4, 1004, 1003.7, 1003.4, 1003.3, 1003.4, 1003.5, 1003.8, 1003.9, 
    1003.8, 1003.7, 1004.1, 1004.9, 1005.3, 1005.5, 1005.6, 1005.9, 1005.9, 
    1006.2, 1006.8, 1007.5, 1008.1, 1008.6, 1009, 1009.3, 1009.4, 1009.5, 
    1009.6, 1009.6, 1009.8, 1010, 1010.3, 1010.7, 1011, 1011.2, 1011.2, 
    1011.1, 1011.1, 1011.1, 1011.4, 1012, 1012.4, 1012.7, 1013.2, 1013.5, 
    1014.1, 1014.6, 1015.2, 1015.9, 1016.5, 1017.3, 1017.8, 1018.5, 1019, 
    1019.8, 1021, 1022.2, 1023.2, 1024.3, 1024.8, 1025.5, 1026.2, 1026.8, 
    1027.2, 1027.7, 1028.3, 1028.9, 1029.5, 1030.2, 1030.7, 1031, 1031.2, 
    1031.6, 1032, 1032.3, 1032.7, 1032.8, 1033.1, 1033.4, 1033.9, 1034.5, 
    1035.4, 1035.9, 1036.6, 1037.2, 1037.7, 1038.2, 1039, 1039.5, 1040.4, 
    1041.2, 1042, 1042.7, 1043.3, 1044.2, 1044.4, 1045, 1045.9, 1046.3, 
    1046.4, 1046.8, 1047.1, 1047.4, 1047.5, 1047.7, 1048.2, 1048.9, 1049.3, 
    1049.9, 1051.1, 1051.3, 1051.6, 1052, 1052.4, 1052.7, 1052.9, 1053.1, 
    1053.1, 1053, 1052.9, 1052.8, 1052.9, 1053, 1053.3, 1053.2, 1053.2, 
    1053.3, 1053.8, 1054.3, 1054.6, 1054.9, 1055.1, 1055.2, 1055.2, 1055.7, 
    1055.8, 1056, 1055.9, 1056, 1056.1, 1056.4, 1056.9, 1057.2, 1057.3, 
    1057.4, 1057.4, 1057.4, 1057.4, 1057.1, 1057, 1057, 1057, 1056.9, 1056.7, 
    1056.7, 1056.5, 1056.2, 1057.8, 1055.7, 1055.4, 1055.2, 1054.6, 1054.6, 
    1054.4, 1054.1, 1053.8, 1053.4, 1053.1, 1052.7, 1052.3, 1051.7, 1051.1, 
    1050.7, 1050.2, 1049.5, 1048.9, 1048.7, 1048.2, 1048, 1047.5, 1046.8, 
    1047.5, 1047, 1044.6, 1043.8, 1043.3, 1042.6, 1042, 1041.5, 1040.9, 
    1040.3, 1039.7, 1038.9, 1038.3, 1037.8, 1037.6, 1037, 1037, 1036.3, 1036, 
    1036, 1035.8, 1035.4, 1035, 1034.6, 1034.5, 1034.3, 1033.8, 1033.9, 
    1033.5, 1033, 1033.2, 1033.5, 1033.8, 1033.8, 1034, 1033.8, 1033.5, 
    1033.3, 1033, 1033, 1032.8, 1032.5, 1032.1, 1031.2, 1031, 1030.8, 1030.3, 
    1029.9, 1029.4, 1028.9, 1028.8, 1028.6, 1028.5, 1028.7, 1028.8, 1029, 
    1029.3, 1029.5, 1029.7, 1029.7, 1029.6, 1029.7, 1030, 1030.2, 1030.3, 
    1030.2, 1030.4, 1030.7, 1030.9, 1030.9, 1030.6, 1030.5, 1031.9, 1030.2, 
    1030.2, 1030.1, 1029.9, 1029.6, 1029.5, 1029.5, 1029.3, 1029.3, 1028.9, 
    1028.7, 1028.4, 1028, 1027.8, 1027.4, 1027, 1026.6, 1026.3, 1026.3, 
    1026.2, 1026, 1025.7, 1025.2, 1024.9, 1024.8, 1024.4, 1024.3, 1024, 
    1023.6, 1023.3, 1023.1, 1022.6, 1022.4, 1022, 1021.5, 1021, 1020.5, 
    1019.9, 1019.4, 1018.9, 1018.6, 1018, 1017.4, 1017, 1016.2, 1015.5, 
    1014.6, 1013.8, 1013, 1012, 1011.8, 1011.1, 1011.1, 1011.4, 1011.9, 
    1011.4, 1011.9, 1012.3, 1012.7, 1012.8, 1012.9, 1012.3, 1013.2, 1013.5, 
    1013.2, 1013, 1013.1, 1012.6, 1012, 1012, 1011.7, 1012, 1012.1, 1012.5, 
    1012.9, 1013.5, 1013.8, 1014.4, 1015, 1015.5, 1016.1, 1016.5, 1016.8, 
    1017.3, 1017.5, 1017.7, 1017.9, 1018.1, 1018.2, 1018.3, 1018.5, 1018.4, 
    1018.4, 1018.2, 1018, 1017.9, 1017.8, 1017.4, 1017.4, 1017.4, 1017.2, 
    1016.9, 1016.8, 1016.7, 1016.6, 1016.4, 1016.1, 1015.8, 1015.4, 1015.3, 
    1015, 1014.6, 1014.4, 1014.3, 1013.9, 1013.7, 1013.5, 1013.4, 1013.4, 
    1013, 1012.6, 1012.2, 1011.9, 1011.5, 1011.2, 1010.8, 1010.6, 1010.3, 
    1009.9, 1009.9, 1009.6, 1009.1, 1008.8, 1008.5, 1008.2, 1007.8, 1007.4, 
    1006.8, 1006.4, 1006, 1005.8, 1005.5, 1005.1, 1004.7, 1004.3, 1003.8, 
    1003.5, 1003.3, 1002.7, 1002.4, 1002.4, 1002.3, 1002.2, 1001.9, 1001.9, 
    1001.7, 1001.7, 1001.7, 1001.9, 1001.9, 1001.7, 1001.7, 1001.7, 1001.7, 
    1001.8, 1001.9, 1002, 1002, 1002.1, 1002.1, 1002, 1002.2, 1002.3, 1002.5, 
    1002.9, 1003.1, 1003.4, 1003.7, 1004.2, 1004.4, 1004.5, 1004.8, 1005, 
    1005.3, 1005.8, 1006.3, 1006.7, 1007.2, 1007.7, 1008.1, 1008.5, 1010.8, 
    1009.1, 1009.4, 1010, 1010.2, 1010.6, 1011.1, 1011.5, 1012.1, 1012.5, 
    1012.7, 1013, 1013.5, 1013.6, 1013.7, 1013.9, 1014.1, 1014.1, 1014.3, 
    1014.6, 1014.9, 1014.8, 1014.9, 1015.7, 1015.3, 1015.4, 1015.3, 1015.4, 
    1015.4, 1015.4, 1015.7, 1015.8, 1016, 1016.4, 1016.6, 1016.7, 1016.8, 
    1016.9, 1017, 1017.2, 1017.6, 1017.8, 1018.1, 1018.4, 1019, 1019.4, 
    1019.5, 1019.8, 1019.9, 1020.1, 1020.3, 1020.6, 1021, 1021.3, 1021.4, 
    1021.7, 1022, 1022, 1022.1, 1022.7, 1022.8, 1022.9, 1022.8, 1022.7, 
    1022.2, 1022.9, 1023.5, 1023.4, 1023.9, 1024.3, 1024.5, 1024.4, 1024.8, 
    1025.2, 1025.4, 1025.3, 1025.4, 1025.4, 1025.4, 1025.2, 1025.7, 1025.6, 
    1025.5, 1025.2, 1024.8, 1024.6, 1024.5, 1024.6, 1025.9, 1026.8, 1027.5, 
    1027.9, 1028.1, 1028.2, 1028.2, 1028, 1027.8, 1027.6, 1027.2, 1026.4, 
    1026.1, 1025.7, 1025.5, 1024.9, 1024.4, 1023.8, 1023.2, 1022.3, 1021.4, 
    1020.7, 1019.8, 1018.9, 1018.2, 1017.8, 1017.3, 1017, 1017.2, 1017, 
    1016.9, 1016.9, 1017, 1017.1, 1017, 1017, 1017.2, 1017.6, 1018.2, 1018.5, 
    1018.7, 1018.7, 1018.8, 1018.7, 1018.3, 1018.2, 1017.8, 1017.6, 1017.1, 
    1016.7, 1016.6, 1016.5, 1016.2, 1015.7, 1015.5, 1015.1, 1015, 1014.8, 
    1014.4, 1013.8, 1013.3, 1012.8, 1012.5, 1012.3, 1011.9, 1011.6, 1011.3, 
    1011, 1010.7, 1010.6, 1010.4, 1010.2, 1010.2, 1009.8, 1009.9, 1010, 
    1010.1, 1010.4, 1010.5, 1010.5, 1010.6, 1010.6, 1010.5, 1010.7, 1010.7, 
    1010.8, 1010.8, 1011, 1011.1, 1011.1, 1011, 1011, 1011, 1011, 1010.8, 
    1010.7, 1010.6, 1010.7, 1010.8, 1010.9, 1011, 1010.8, 1010.8, 1010.7, 
    1010.4, 1010.4, 1010.3, 1010.4, 1010.4, 1010.3, 1010.3, 1010.4, 1010.5, 
    1010.4, 1010.4, 1010.4, 1010.5, 1010.6, 1010.4, 1010.2, 1010.3, 1010.5, 
    1010.9, 1011.2, 1011.5, 1011.4, 1011.3, 1011.6, 1011.6, 1011.8, 1011.5, 
    1011.9, 1012.2, 1012.4, 1012.7, 1012.9, 1013.3, 1013.8, 1014.1, 1014.2, 
    1014.4, 1014.8, 1015.1, 1015.1, 1015.2, 1015.7, 1016, 1016.4, 1016.5, 
    1016.5, 1016.4, 1016.4, 1016.4, 1016.6, 1016.7, 1016.5, 1016.2, 1016, 
    1016.1, 1016, 1015.9, 1015.7, 1015.4, 1015.2, 1015, 1015, 1014.9, 1014.5, 
    1014.4, 1014.3, 1014.3, 1014.3, 1014.4, 1014.4, 1014.4, 1014.3, 1014.2, 
    1014.2, 1014, 1014, 1013.8, 1013.8, 1014, 1014.2, 1014.2, 1014.1, 1014, 
    1013.7, 1013.5, 1013.5, 1013.3, 1013.2, 1013.1, 1012.9, 1012.6, 1012.6, 
    1012.5, 1012.3, 1012.1, 1012, 1011.8, 1011.7, 1011.5, 1011.4, 1011.2, 
    1011, 1010.9, 1010.9, 1010.7, 1010.7, 1010.7, 1010.5, 1010.4, 1010.3, 
    1010.3, 1010, 1010, 1009.8, 1009.9, 1009.8, 1009.8, 1009.7, 1009.5, 
    1009.5, 1009.4, 1009.3, 1009.5, 1009.4, 1009.3, 1009.3, 1009.3, 1009.3, 
    1009.4, 1009.5, 1009.6, 1009.6, 1009.7, 1010, 1010.2, 1010.3, 1010.6, 
    1010.7, 1010.8, 1011, 1011.1, 1011.3, 1011.6, 1011.8, 1011.7, 1011.7, 
    1011.9, 1011.7, 1011.6, 1011.8, 1011.8, 1011.9, 1011.6, 1011.6, 1011.3, 
    1011.1, 1011, 1010.6, 1010.1, 1009.7, 1009.2, 1008.8, 1008.4, 1007.9, 
    1007.6, 1007.1, 1006.7, 1006.2, 1005.8, 1005.4, 1004.8, 1004.4, 1004.1, 
    1003.7, 1003.6, 1003.4, 1003.2, 1003.2, 1003, 1003, 1003, 1003, 1003, 
    1003.3, 1003.1, 1003.4, 1003.5, 1003.8, 1003.8, 1004.1, 1004.3, 1004.6, 
    1004.8, 1004.9, 1004.9, 1004.7, 1004.5, 1004.7, 1004.8, 1004.8, 1004.7, 
    1004.7, 1004.7, 1005, 1004.8, 1004.8, 1004.6, 1004.6, 1004.5, 1004.6, 
    1004.6, 1004.7, 1004.6, 1004.4, 1004.3, 1004.3, 1004.3, 1004, 1003.8, 
    1003.7, 1003.8, 1003.9, 1004.1, 1004.5, 1004.7, 1004.7, 1005.1, 1005.2, 
    1005.5, 1005.7, 1006.3, 1006.7, 1006.9, 1007.3, 1008.8, 1008.3, 1008.7, 
    1009, 1009.3, 1009.8, 1010.3, 1010.7, 1011, 1011.5, 1012.1, 1012.4, 
    1012.8, 1013.4, 1013.9, 1014.3, 1014.7, 1015.1, 1015.3, 1015.8, 1015.8, 
    1016, 1016.4, 1016.6, 1016.7, 1016.9, 1017.3, 1017.5, 1017.4, 1017.5, 
    1017.5, 1017.4, 1017.4, 1017.3, 1017.1, 1017, 1016.9, 1016.7, 1016.2, 
    1015.8, 1015.4, 1015.1, 1014.7, 1014.3, 1013.5, 1012.4, 1011.6, 1010.8, 
    1009.6, 1008.1, 1006.7, 1004.6, 1003, 1001.5, 1000, 998.2, 997.2, 996.4, 
    996, 995.9, 995.8, 995.9, 996.1, 996.5, 996.6, 996.5, 996.2, 996, 995.6, 
    995.2, 994.9, 994.5, 994, 993.4, 992.9, 992.6, 992.2, 991.7, 991.5, 
    991.3, 991.2, 991.1, 991.1, 991.1, 991.8, 991.3, 991.5, 991.9, 992.1, 
    992.3, 992.5, 992.8, 992.6, 992.7, 992.8, 992.9, 993.2, 993.2, 993.1, 
    993.1, 993, 992.6, 992.4, 991.9, 992, 991.6, 991.3, 991.1, 990.6, 990.5, 
    990.2, 990, 990, 990.1, 990.1, 990.3, 990.5, 990.6, 990.9, 991.3, 991.6, 
    991.9, 992.3, 992.7, 993, 993.3, 993.5, 994, 994.3, 994.6, 995.1, 995.4, 
    995.7, 995.9, 996.1, 996.3, 996.6, 996.9, 997.2, 997.3, 997.6, 997.9, 
    998.4, 998.7, 999.1, 999.5, 999.7, 1000, 1000.2, 1000.5, 1000.7, 1000.7, 
    1000.8, 1001, 1001.1, 1001.4, 1001.5, 1001.4, 1001.4, 1001.3, 1001.1, 
    1000.9, 1000.9, 1000.9, 1000.9, 1000.9, 1001.1, 1001.4, 1001.6, 1001.9, 
    1002.1, 1002.6, 1002.8, 1003.1, 1003.5, 1003.6, 1003.9, 1004.2, 1004.6, 
    1004.9, 1005.5, 1005.8, 1006.2, 1006.7, 1007.4, 1007.9, 1008.3, 1008.7, 
    1009.1, 1009.5, 1009.7, 1010.1, 1010.5, 1010.9, 1011.2, 1011.3, 1011.6, 
    1011.9, 1011.9, 1011.9, 1011.8, 1011.6, 1011.4, 1011.3, 1011.1, 1011.2, 
    1011.1, 1010.8, 1010.7, 1010.5, 1010.6, 1010.2, 1009.8, 1009.5, 1009.1, 
    1008.7, 1008.1, 1007.6, 1007.4, 1007.1, 1006.5, 1006.4, 1006.1, 1005.8, 
    1005.7, 1005.6, 1005.3, 1005.4, 1005.5, 1005.6, 1005.6, 1005.9, 1006.2, 
    1006.4, 1006.8, 1006.9, 1007.2, 1007.1, 1007.3, 1007.6, 1007.7, 1007.9, 
    1008.2, 1008.3, 1008.5, 1008.6, 1008.5, 1008.5, 1008.8, 1008.8, 1008.8, 
    1008.7, 1009, 1009.3, 1009.5, 1009.6, 1009.9, 1010.1, 1010.3, 1010.5, 
    1010.4, 1010.4, 1010.6, 1010.9, 1011.1, 1011.3, 1011.6, 1011.9, 1011.9, 
    1011.9, 1011.9, 1012, 1012.2, 1012.1, 1012.2, 1012.4, 1012.3, 1012.5, 
    1012.8, 1012.8, 1012.7, 1012.6, 1012.3, 1012.3, 1012, 1012, 1011.8, 
    1011.5, 1011.4, 1011.2, 1011.1, 1010.8, 1010.6, 1010.4, 1010.1, 1009.9, 
    1009.6, 1009.4, 1009.3, 1009.5, 1009.5, 1009.5, 1009.4, 1009.2, 1009, 
    1008.9, 1008.8, 1008.6, 1008.4, 1008, 1007.7, 1007.1, 1007.1, 1006.8, 
    1006.3, 1006.3, 1005.9, 1005.5, 1005.2, 1005, 1004.6, 1004.5, 1004.7, 
    1004.7, 1004.7, 1004.9, 1005.2, 1005.3, 1005.4, 1005.6, 1005.7, 1006, 
    1006.2, 1006.2, 1006.4, 1006.6, 1006.6, 1007.1, 1007.5, 1007.8, 1008.2, 
    1008.6, 1008.8, 1009.1, 1009.3, 1009.7, 1010, 1010.1, 1010.4, 1010.9, 
    1011.4, 1011.6, 1011.7, 1012, 1012.1, 1012.2, 1012.5, 1012.5, 1012.4, 
    1012.9, 1013.2, 1013.3, 1013.7, 1014, 1014.1, 1014.2, 1014.3, 1014.1, 
    1014.1, 1014.1, 1014.1, 1014.2, 1014.4, 1014.6, 1014.6, 1014.8, 1015.1, 
    1015.1, 1015.5, 1015.8, 1015.8, 1015.8, 1015.9, 1015.9, 1016.1, 1016.2, 
    1016.4, 1016.6, 1016.4, 1016.3, 1015.9, 1015.7, 1015.5, 1015.4, 1015.2, 
    1014.8, 1014.6, 1014.4, 1014.3, 1014.2, 1013.9, 1013.6, 1013.3, 1012.9, 
    1012.3, 1011.9, 1011.6, 1011.2, 1011, 1010.8, 1010.4, 1010, 1009.6, 
    1009.4, 1009.1, 1008.9, 1008.6, 1008.2, 1007.6, 1007.3, 1006.8, 1006.6, 
    1006.1, 1005.9, 1005.6, 1005.5, 1005.4, 1005.2, 1005.1, 1005.2, 1005.2, 
    1005.5, 1005.8, 1006.1, 1006.4, 1006.6, 1006.9, 1007.2, 1007.5, 1007.7, 
    1008, 1008.3, 1008.6, 1009.3, 1009.6, 1010.2, 1010.6, 1011, 1011.6, 
    1011.8, 1012.2, 1012.5, 1012.7, 1013, 1013.1, 1013.6, 1014, 1014.4, 
    1014.8, 1015.2, 1015.3, 1015.6, 1016, 1016, 1015.9, 1016.1, 1016.2, 
    1016.3, 1016.3, 1016.4, 1016.3, 1016.2, 1016.2, 1016, 1015.9, 1015.6, 
    1015.5, 1015.3, 1015, 1014.9, 1014.6, 1014.6, 1014.5, 1014.3, 1014, 
    1013.8, 1013.3, 1012.8, 1012.5, 1011.4, 1011.2, 1010.5, 1010.2, 1009.9, 
    1009.8, 1009.8, 1009.7, 1009.8, 1009.9, 1009.7, 1009.6, 1009.5, 1009.5, 
    1009.5, 1009.8, 1010, 1010.2, 1010.6, 1010.8, 1011.1, 1011.2, 1011.4, 
    1011.5, 1011.9, 1012.3, 1012.8, 1013, 1013.3, 1013.8, 1014.3, 1014.7, 
    1015, 1015.5, 1016, 1016.4, 1016.6, 1017, 1017.5, 1018, 1018.7, 1019, 
    1019.3, 1019.4, 1019.8, 1020.1, 1020.2, 1020.4, 1020.6, 1020.8, 1021.1, 
    1021.5, 1021.8, 1022, 1022.1, 1022.6, 1022.9, 1023.1, 1023.4, 1023.5, 
    1024, 1024.2, 1024.4, 1024.9, 1025.3, 1025.9, 1026.2, 1026.6, 1026.8, 
    1027.2, 1027.5, 1027.9, 1028.1, 1028.3, 1028.6, 1028.9, 1029.1, 1029.4, 
    1029.7, 1029.7, 1029.7, 1029.8, 1029.8, 1029.7, 1029.7, 1029.5, 1029.7, 
    1029.7, 1029.7, 1029.7, 1029.6, 1029.4, 1029.3, 1029, 1028.7, 1028.4, 
    1028.2, 1028.2, 1028, 1027.9, 1027.9, 1027.7, 1027.6, 1027.4, 1027.3, 
    1027.1, 1027, 1026.8, 1026.4, 1026.3, 1026.1, 1026, 1026, 1026, 1025.9, 
    1025.6, 1025.3, 1025.1, 1024.9, 1024.6, 1024.4, 1024.4, 1024.5, 1024.6, 
    1024.5, 1024.4, 1024.3, 1024.4, 1024.5, 1024.3, 1024.5, 1024.5, 1024.4, 
    1024.6, 1024.9, 1025.2, 1025.5, 1025.8, 1026, 1026.2, 1026.5, 1026.8, 
    1027.3, 1027.7, 1028, 1028.3, 1028.7, 1029.1, 1029.5, 1029.8, 1030.2, 
    1030.5, 1030.7, 1030.6, 1030.8, 1031, 1031.2, 1031.2, 1031.3, 1031.2, 
    1031.1, 1031.1, 1031.4, 1031.2, 1030.6, 1030.6, 1030.3, 1029.6, 1028.9, 
    1028.6, 1028.2, 1027.7, 1027.4, 1026.7, 1025.8, 1025.5, 1024.4, 1022.8, 
    1021.9, 1020.7, 1019.3, 1018.1, 1017.1, 1016, 1015.1, 1014.3, 1013.5, 
    1012.7, 1012, 1011.5, 1010.7, 1010.1, 1009.8, 1009.6, 1009.7, 1009.9, 
    1010, 1010.6, 1011.1, 1011.7, 1012, 1012.8, 1013.4, 1013.9, 1014.5, 
    1014.8, 1015.4, 1015.9, 1016.7, 1017.5, 1018.3, 1019.1, 1020, 1020.6, 
    1021.3, 1022, 1022.7, 1023.1, 1023.5, 1023.7, 1024.4, 1025, 1025.4, 
    1025.8, 1025.7, 1025.9, 1026.1, 1026, 1025.9, 1025.8, 1025.7, 1025.7, 
    1025.6, 1025.4, 1025.3, 1025.3, 1025, 1025, 1024.6, 1024.3, 1023.9, 
    1023.6, 1023.4, 1023.4, 1023.4, 1023.5, 1023.6, 1023.5, 1023.5, 1023.3, 
    1023.1, 1022.7, 1022.5, 1022.3, 1022, 1021.5, 1021.5, 1021.5, 1021.3, 
    1021, 1020.7, 1020.4, 1020, 1019.9, 1019.7, 1019.4, 1019.2, 1019.4, 
    1019.3, 1019.5, 1019.6, 1019.6, 1019.5, 1019.3, 1019.3, 1019.4, 1019.6, 
    1020, 1020.1, 1020.4, 1021, 1021.2, 1021.7, 1021.7, 1021.9, 1021.8, 
    1022.1, 1022.1, 1022.1, 1022.1, 1022.4, 1022.4, 1022.7, 1022.9, 1023.1, 
    1023.3, 1023.1, 1023.2, 1023.3, 1023.5, 1023.6, 1023.4, 1023.4, 1023.7, 
    1024, 1024, 1023.8, 1023.5, 1023.3, 1022.7, 1022.3, 1021.7, 1021.4, 
    1020.8, 1020.5, 1020.1, 1019.7, 1019.2, 1018.8, 1018.4, 1017.6, 1016.9, 
    1016, 1014.9, 1014, 1013.1, 1012.3, 1011.5, 1010.8, 1010.1, 1009.5, 
    1008.9, 1008, 1007.6, 1006.8, 1005.8, 1004.8, 1004.2, 1003.5, 1002.7, 
    1002.2, 1002, 1001.7, 1001.3, 1001, 1000.6, 1000.9, 1001, 1001.2, 1001.5, 
    1001.6, 1002.3, 1003, 1003.7, 1004.3, 1005.6, 1006.5, 1007.4, 1008.2, 
    1008.9, 1009.5, 1010.2, 1011.2, 1012.2, 1013.2, 1014.1, 1015, 1015.8, 
    1016.5, 1017.3, 1018, 1018.6, 1019.2, 1019.8, 1020.5, 1021, 1021.3, 
    1021.4, 1021.8, 1022.1, 1022.3, 1022.1, 1022.3, 1022.1, 1021.9, 1021.7, 
    1021.9, 1021.8, 1021.7, 1021.8, 1021.7, 1021.5, 1021.4, 1021.4, 1021.1, 
    1020.8, 1020.8, 1020.6, 1020.4, 1020.2, 1020, 1020, 1019.9, 1019.8, 
    1019.6, 1019.1, 1019, 1018.7, 1018.4, 1018.1, 1018, 1017.9, 1017.7, 
    1017.8, 1017.9, 1018, 1018, 1017.8, 1017.5, 1017.4, 1017.4, 1017.4, 
    1017.4, 1017.7, 1018.1, 1018.6, 1019.1, 1019.9, 1020.6, 1020.8, 1021.3, 
    1021.7, 1022, 1022.6, 1023.1, 1023.5, 1023.9, 1024.3, 1024.7, 1025.1, 
    1025.2, 1025.2, 1025.3, 1025.5, 1025.7, 1025.5, 1025.4, 1025.5, 1025.3, 
    1024.8, 1024.2, 1023.6, 1022.4, 1021.7, 1021.4, 1020.9, 1020.4, 1020.5, 
    1021, 1021.4, 1021.9, 1022.5, 1022.9, 1023.2, 1023.4, 1023.9, 1024.1, 
    1023.9, 1023.5, 1023.3, 1023.1, 1023.1, 1023.1, 1023, 1022.7, 1022.4, 
    1022, 1021.5, 1020.9, 1020.6, 1020.1, 1019.5, 1019, 1018.5, 1018.1, 
    1017.7, 1017.6, 1017.3, 1017.1, 1016.5, 1016.3, 1016, 1015.7, 1015.5, 
    1015.7, 1015.5, 1015.5, 1015.6, 1015.7, 1015.8, 1016.1, 1015.9, 1016.2, 
    1016.3, 1016.5, 1016.6, 1017, 1017.5, 1018, 1018.3, 1018.7, 1018.9, 
    1019.3, 1019.6, 1019.8, 1020.1, 1020.4, 1020.8, 1021, 1021.4, 1022, 
    1022.2, 1022.7, 1022.8, 1023.1, 1023.4, 1023.7, 1023.9, 1024.1, 1024.3, 
    1024.6, 1024.9, 1025.2, 1025.5, 1025.8, 1025.8, 1025.9, 1025.7, 1025.7, 
    1025.5, 1025.6, 1025.6, 1025.6, 1025.5, 1025.6, 1025.7, 1025.6, 1025.6, 
    1025.5, 1025.2, 1025.1, 1024.7, 1024.3, 1023.9, 1023.5, 1023.4, 1023.7, 
    1023.6, 1023, 1022.8, 1022.5, 1022, 1021.4, 1021.3, 1020.8, 1020.3, 
    1020.1, 1019.7, 1019.6, 1019.2, 1018.5, 1017.9, 1017.1, 1016.4, 1016.2, 
    1015.3, 1014.6, 1014.4, 1014, 1014.3, 1014.3, 1014.4, 1014.4, 1014.3, 
    1013.9, 1013.4, 1012.3, 1011.5, 1010.7, 1010.4, 1010.2, 1009.9, 1010.2, 
    1010.7, 1011.3, 1011.5, 1011.9, 1011.9, 1012.8, 1013, 1013.9, 1014.4, 
    1014.7, 1015.5, 1015.9, 1016.6, 1017, 1017.2, 1017.2, 1017.4, 1017.9, 
    1018.4, 1018.5, 1019.1, 1019.4, 1019.5, 1019.7, 1019.8, 1019.7, 1019.2, 
    1018.5, 1017.6, 1017, 1016.5, 1015.9, 1015.6, 1015.4, 1014.7, 1014.3, 
    1014.4, 1014.5, 1014.1, 1014, 1013.5, 1013.1, 1012.9, 1012.8, 1012.7, 
    1012.7, 1012.7, 1012.8, 1013.1, 1013, 1013, 1012.8, 1012.8, 1012.9, 
    1012.9, 1013.1, 1013.2, 1013.4, 1014, 1014.1, 1014.2, 1014.3, 1014.1, 
    1014.5, 1014.2, 1014.1, 1014.3, 1014, 1013.6, 1013.2, 1012.8, 1012.8, 
    1012.1, 1011.4, 1010.7, 1009.9, 1009.1, 1008.1, 1007.6, 1007.3, 1006.8, 
    1007.3, 1007.7, 1008.2, 1008.9, 1010.2, 1011.3, 1012.1, 1013, 1013.6, 
    1014.4, 1014.7, 1015, 1015.2, 1015.4, 1015.8, 1016.1, 1016.4, 1016.5, 
    1016.6, 1016.7, 1016.7, 1016.6, 1016.6, 1016.5, 1016.7, 1016.5, 1016.5, 
    1016.8, 1016.6, 1016.5, 1016.1, 1015.8, 1015.6, 1015.3, 1014.8, 1014.3, 
    1013.8, 1013.3, 1013, 1012.7, 1012, 1011.4, 1010.9, 1010.2, 1009.5, 
    1008.9, 1008.3, 1007.7, 1007.6, 1007.5, 1007.4, 1007.3, 1007.3, 1007.5, 
    1007.8, 1007.9, 1008, 1008.1, 1008.3, 1008.4, 1008.5, 1009.1, 1009.5, 
    1010, 1010.5, 1010.9, 1011, 1011, 1011.3, 1011.4, 1011.2, 1011.4, 1011.5, 
    1011.5, 1011.3, 1011.6, 1011.6, 1011.4, 1011.4, 1011.4, 1011.7, 1011.9, 
    1012.1, 1011.9, 1012.4, 1012.6, 1012.9, 1013.1, 1013.5, 1013.7, 1013.9, 
    1014.1, 1014.2, 1014.2, 1014.3, 1014.3, 1014.3, 1014.4, 1014.5, 1014.6, 
    1014.7, 1014.6, 1014.5, 1014.1, 1013.8, 1013.3, 1012.8, 1012.3, 1012, 
    1011.8, 1011.6, 1011.4, 1011, 1010.7, 1010.1, 1009.7, 1009.1, 1008.8, 
    1008.4, 1008, 1008, 1007.9, 1007.9, 1008, 1008, 1008, 1007.8, 1007.7, 
    1007.8, 1008.1, 1008.2, 1008.5, 1008.6, 1008.7, 1009.1, 1009.2, 1009.3, 
    1009.4, 1009.4, 1009.2, 1008.9, 1008.8, 1008.5, 1008.3, 1008.1, 1007.9, 
    1007.8, 1007.4, 1007.3, 1006.6, 1006.2, 1006, 1005.9, 1005.5, 1005.2, 
    1004.8, 1004.1, 1003.6, 1003.7, 1003.5, 1003.2, 1002.7, 1002.4, 1002.3, 
    1001.9, 1001.5, 1001, 1000.8, 1000.6, 1000.6, 1000.9, 1001, 1001.1, 
    1001.3, 1001.3, 1001.3, 1001.4, 1001.4, 1001.5, 1001.4, 1001.2, 1001.1, 
    1001.2, 1001.1, 1001.2, 1001.4, 1001.6, 1001.9, 1002, 1002.2, 1002.2, 
    1002.2, 1002.6, 1002.9, 1003.3, 1003.5, 1003.9, 1004.2, 1004.5, 1004.7, 
    1004.9, 1005, 1005.2, 1005.3, 1005.3, 1005.4, 1005.5, 1005.7, 1005.8, 
    1005.8, 1005.9, 1005.9, 1005.9, 1005.7, 1005.7, 1005.6, 1005.6, 1005.4, 
    1005.5, 1005.3, 1005.3, 1005.4, 1005.5, 1005.5, 1005.3, 1004.9, 1004.5, 
    1004.1, 1003.9, 1003.8, 1003.9, 1003.8, 1003.8, 1003.7, 1003.6, 1003.3, 
    1002.9, 1002.5, 1002.4, 1002.1, 1001.7, 1001.6, 1001.7, 1001.9, 1002.1, 
    1002.4, 1002.4, 1002.7, 1003, 1002.9, 1002.6, 1002.8, 1003, 1003.2, 
    1003.4, 1003.5, 1003.6, 1003.9, 1004.2, 1004.4, 1004.8, 1005, 1005, 
    1005.1, 1005.3, 1005.8, 1005.9, 1006.2, 1006.1, 1006.3, 1006.5, 1006.8, 
    1007.1, 1007, 1007.4, 1007.4, 1007.5, 1007.5, 1007.6, 1007.9, 1008.3, 
    1008.7, 1009.3, 1009.5, 1009.8, 1010, 1010.1, 1010.2, 1010.3, 1010.4, 
    1010.6, 1010.8, 1011.1, 1011, 1011.2, 1011.1, 1011, 1010.6, 1010.7, 
    1010.2, 1009.8, 1009.7, 1009.5, 1009.7, 1009.8, 1009.7, 1009.6, 1009.4, 
    1009.3, 1009.3, 1009.3, 1009.2, 1009.3, 1009.2, 1009.2, 1009.3, 1009.1, 
    1009, 1008.6, 1008.5, 1008.3, 1008.3, 1008, 1007.9, 1007.8, 1007.9, 
    1007.9, 1008, 1007.9, 1007.7, 1007.7, 1007.9, 1008, 1007.9, 1007.9, 
    1008.1, 1008.1, 1008, 1008.3, 1008.4, 1008.7, 1008.8, 1008.9, 1009, 1009, 
    1009.3, 1009.3, 1009.7, 1010, 1010.4, 1010.8, 1011.1, 1011.3, 1011.4, 
    1011.3, 1011.2, 1011, 1011, 1010.9, 1010.6, 1010.1, 1009.8, 1009.7, 
    1009.5, 1009.3, 1008.8, 1008.5, 1008.3, 1007.7, 1007.2, 1006.7, 1006, 
    1005.3, 1004.9, 1004.5, 1003.7, 1003.3, 1002.7, 1002.3, 1001.7, 1001.3, 
    1000.9, 1000.4, 1000.2, 1000.1, 999.8, 999.9, 999.8, 999.7, 999.6, 999.6, 
    999.6, 999.6, 999.6, 1000, 1000.2, 1000.3, 1000.8, 1001.2, 1001.8, 
    1002.5, 1002.7, 1002.9, 1003.7, 1004.2, 1004.8, 1005.2, 1005.5, 1006.1, 
    1007.2, 1008, 1008.9, 1009.7, 1010.5, 1011.1, 1011.9, 1012.5, 1012.9, 
    1013.5, 1014, 1013.3, 1013.8, 1014.2, 1015.4, 1015.6, 1015.7, 1015.9, 
    1015.8, 1015.9, 1015.9, 1015.9, 1016, 1015.9, 1015.8, 1015.7, 1015.5, 
    1015.5, 1015.5, 1015.4, 1015.3, 1015, 1014.9, 1014.6, 1014.2, 1013.8, 
    1013.7, 1013.6, 1013.5, 1013.4, 1013.2, 1013.1, 1013, 1012.9, 1012.8, 
    1012.5, 1012.3, 1012.3, 1012.3, 1012.6, 1012.8, 1012.6, 1012.4, 1012.2, 
    1012.1, 1011.6, 1011.3, 1011.1, 1011.3, 1011.5, 1011.7, 1012, 1012.3, 
    1012.6, 1012.8, 1012.9, 1013.2, 1013.4, 1013.2, 1013.2, 1013.4, 1013.4, 
    1013.5, 1013.8, 1014.1, 1014.4, 1014.7, 1014.9, 1015.2, 1015.3, 1015.2, 
    1015.1, 1014.9, 1015, 1014.9, 1014.8, 1014.6, 1014.3, 1013.9, 1014, 
    1013.9, 1013.8, 1013.4, 1013.1, 1013.2, 1013.1, 1013.3, 1013.8, 1014.4, 
    1015, 1015.6, 1015.9, 1016, 1016, 1015.8, 1015.6, 1015.4, 1015.1, 1015.1, 
    1014.7, 1014.3, 1014.2, 1013.8, 1013.3, 1012.8, 1012, 1011.3, 1010.6, 
    1010, 1009.6, 1009.1, 1008.6, 1008.2, 1007.9, 1007.6, 1007.7, 1007.6, 
    1007.6, 1007.5, 1007.8, 1008, 1008.3, 1009.1, 1009.5, 1010.1, 1010.3, 
    1010.5, 1010.9, 1010.6, 1010.4, 1010.1, 1010.1, 1009.5, 1009.1, 1008.4, 
    1007.8, 1007.8, 1007.3, 1006.4, 1006.2, 1005.7, 1005.6, 1005.3, 1005, 
    1004.9, 1004.8, 1005.7, 1006.3, 1007.1, 1007.2, 1007.4, 1007.6, 1007.3, 
    1007.3, 1007.3, 1007.3, 1007.1, 1007, 1007, 1007.2, 1007.3, 1007.3, 
    1007.2, 1007, 1007, 1007.2, 1007, 1006.6, 1006.1, 1005.9, 1005.9, 1006.2, 
    1006.9, 1007.4, 1007.8, 1008.3, 1008.6, 1008.7, 1009.1, 1009.3, 1009.8, 
    1010.1, 1010.1, 1010.4, 1010.6, 1010.8, 1010.8, 1010.8, 1010.8, 1010.8, 
    1010.7, 1010.8, 1011.1, 1011, 1011.4, 1011.9, 1012.2, 1012.2, 1011.9, 
    1011.9, 1011.9, 1011.7, 1011.5, 1011.5, 1011.3, 1011.2, 1011.1, 1011.1, 
    1011.1, 1010.7, 1010.2, 1010, 1009.5, 1009.4, 1009.1, 1008.7, 1008.3, 
    1007.9, 1007.5, 1007.3, 1007.4, 1007, 1006.8, 1006.5, 1005.9, 1005.6, 
    1005.4, 1005, 1004.7, 1004.2, 1003.9, 1004, 1003.7, 1003.4, 1003.5, 
    1003.3, 1003.3, 1003.4, 1003.3, 1003.2, 1003.2, 1003.2, 1003.2, 1003.2, 
    1003.4, 1003.4, 1003.4, 1003.3, 1003.4, 1003.5, 1003.7, 1003.8, 1003.8, 
    1004.1, 1004.6, 1004.9, 1005.3, 1005.6, 1006, 1006.4, 1006.5, 1006.6, 
    1006.7, 1006.8, 1007, 1007.2, 1007.1, 1006.9, 1006.7, 1006.6, 1006.5, 
    1006.2, 1005.8, 1005.7, 1005.5, 1005.3, 1005.1, 1005.2, 1005.6, 1006.1, 
    1006.3, 1006.7, 1006.9, 1006.8, 1006.5, 1006.2, 1005.9, 1005.8, 1005.9, 
    1005.8, 1005.8, 1006, 1006.2, 1006.2, 1006.1, 1006.2, 1005.9, 1005.6, 
    1005.2, 1004.6, 1004.2, 1003.9, 1003.4, 1003.2, 1002.9, 1002.6, 1002.4, 
    1002, 1001.8, 1001.3, 1000.6, 999.9, 999.9, 1000.1, 1000.6, 1001.3, 
    1001.7, 1001.9, 1002.2, 1002.3, 1002, 1001.7, 1001.4, 1001.3, 1001, 
    1000.8, 1000.8, 1000.5, 1000.4, 1000.5, 1000.3, 1000, 999.8, 999.6, 
    999.6, 999.4, 999.3, 999.2, 999.1, 999.1, 999.1, 999.2, 999.1, 999, 
    998.9, 999, 999, 998.9, 998.8, 998.8, 998.8, 999, 999.1, 999.1, 999, 
    998.8, 998.5, 998.3, 997.9, 997.8, 997.8, 997.6, 997.3, 997.2, 997.2, 
    997.2, 996.8, 996.6, 996.5, 996.4, 996.2, 996.1, 996.1, 996, 996, 996.2, 
    996.2, 996.4, 996.7, 996.8, 997, 997, 997.1, 997.4, 997.5, 997.8, 998.1, 
    998.5, 999.1, 999.2, 999.6, 999.9, 1000.4, 1000.7, 1001.1, 1001.4, 
    1001.8, 1002.2, 1002.6, 1003, 1003.3, 1003.8, 1004.2, 1004.7, 1005, 
    1005.4, 1005.8, 1006.1, 1006.2, 1006.7, 1007.1, 1007.7, 1008.2, 1008.8, 
    1009.3, 1009.9, 1010.3, 1010.7, 1011.2, 1011.5, 1011.9, 1012.3, 1012.8, 
    1013.2, 1013.8, 1014.2, 1014.7, 1015.1, 1015.3, 1015.5, 1015.7, 1015.9, 
    1016.1, 1016.1, 1016.1, 1016.3, 1016.3, 1016.3, 1016.2, 1016.2, 1016.2, 
    1016, 1015.9, 1015.7, 1015.5, 1015.4, 1015.2, 1014.7, 1014.4, 1014.1, 
    1014, 1013.6, 1013.3, 1012.9, 1012.5, 1012.1, 1011.7, 1011.6, 1011.3, 
    1011, 1011.1, 1010.8, 1010.4, 1010.2, 1009.7, 1009.6, 1009.3, 1008.9, 
    1008.4, 1008, 1007.6, 1007.3, 1007, 1006.8, 1006.5, 1006.2, 1006.1, 
    1005.3, 1005.1, 1004.8, 1004.6, 1004.2, 1004, 1003.4, 1003.1, 1002.6, 
    1002.4, 1002.7, 1002.1, 1001.7, 1001.4, 1001.1, 1000.9, 1000.2, 1000.1, 
    999.8, 999.5, 999.2, 999.2, 998.8, 998.5, 998, 997.8, 997.6, 997.3, 997, 
    997.1, 996.8, 997, 997.1, 997, 997.3, 997.7, 998, 998, 998.2, 998.4, 
    998.3, 998.3, 998.6, 998.9, 999.3, 999.7, 1000.1, 1000.4, 1000.8, 1001.1, 
    1001.5, 1001.7, 1002.3, 1002.9, 1003.4, 1003.7, 1004.3, 1004.6, 1005.1, 
    1005.5, 1005.7, 1006, 1006.3, 1006.5, 1006.9, 1007.2, 1007.8, 1008, 
    1008.5, 1008.9, 1009.3, 1009.7, 1010, 1010.2, 1010.4, 1010.7, 1010.8, 
    1011, 1011.1, 1011.5, 1011.7, 1011.9, 1012, 1012.1, 1012.2, 1012.2, 
    1012.2, 1012.5, 1012.8, 1013, 1013.2, 1013.3, 1013.5, 1013.8, 1013.9, 
    1014.1, 1014.2, 1014.3, 1014.5, 1014.8, 1015, 1015.4, 1015.7, 1016, 
    1016.3, 1016.7, 1017, 1017, 1017.3, 1017.4, 1017.2, 1017.3, 1017.5, 
    1017.7, 1018, 1017.8, 1018, 1017.9, 1017.9, 1017.9, 1017.9, 1017.8, 
    1017.7, 1017.4, 1016.8, 1016.4, 1016.1, 1015.5, 1015.2, 1014.4, 1013.7, 
    1013.1, 1012.5, 1011.5, 1010.5, 1009.5, 1009, 1007.8, 1007, 1006.5, 
    1006.1, 1005.2, 1004.7, 1004.3, 1003.2, 1002.4, 1001.7, 1001.2, 1000.5, 
    999.9, 999.6, 999.4, 999.3, 999.3, 999.4, 999.4, 999.6, 999.9, 1000, 
    1000.1, 1000.2, 1000.9, 1001.6, 1002.7, 1003.2, 1003.8, 1004.4, 1005.1, 
    1005.6, 1006.1, 1006.8, 1007.3, 1007.6, 1007.6, 1008, 1008.5, 1008.8, 
    1009, 1009.2, 1009.4, 1009.7, 1009.8, 1010.1, 1010.6, 1011, 1011.3, 
    1011.2, 1011.3, 1011.5, 1011.6, 1011.6, 1011.7, 1011.8, 1011.9, 1012.1, 
    1012.3, 1012.7, 1013.1, 1013.3, 1013.6, 1013.9, 1014.3, 1014.4, 1014.5, 
    1014.7, 1014.8, 1015, 1015.1, 1015, 1015.1, 1015.3, 1015.6, 1015.7, 
    1015.6, 1015.8, 1015.9, 1016, 1015.8, 1016.1, 1016.3, 1016.4, 1016.5, 
    1016.8, 1017, 1017.1, 1017.3, 1017.4, 1017.5, 1017.3, 1017.3, 1017.5, 
    1017.6, 1017.5, 1017.5, 1017.2, 1017.2, 1017.1, 1017.1, 1017.3, 1017.5, 
    1017.2, 1017, 1016.7, 1016.7, 1016.7, 1016.7, 1016.5, 1016.5, 1016.4, 
    1016.4, 1016.4, 1016.3, 1016.2, 1015.9, 1015.7, 1015.7, 1015.6, 1015.4, 
    1015.2, 1015.1, 1014.9, 1014.9, 1014.9, 1014.8, 1014.8, 1014.7, 1014.7, 
    1014.8, 1014.7, 1014.7, 1014.8, 1014.8, 1014.7, 1014.7, 1014.7, 1014.6, 
    1014.4, 1014.1, 1013.7, 1013.4, 1013.1, 1012.8, 1012.5, 1012.3, 1012.2, 
    1012.1, 1011.9, 1011.4, 1011, 1010.6, 1010.5, 1010.2, 1009.7, 1009.6, 
    1009.5, 1009.4, 1009.3, 1009, 1009, 1008.9, 1009, 1008.8, 1008.7, 1008.8, 
    1008.8, 1009, 1009.1, 1009.1, 1009.1, 1009.5, 1009.7, 1009.7, 1009.9, 
    1009.9, 1009.9, 1010, 1010.3, 1010.8, 1011.3, 1011.6, 1011.8, 1012.3, 
    1012.6, 1012.9, 1013.3, 1013.5, 1013.8, 1013.8, 1014, 1014.4, 1014.6, 
    1014.7, 1014.7, 1014.8, 1014.7, 1014.6, 1014.4, 1014.4, 1014.3, 1014.4, 
    1014.3, 1014.4, 1014.3, 1014.5, 1014.5, 1014.7, 1014.5, 1014.5, 1014.6, 
    1014.6, 1014.4, 1014.3, 1014.5, 1014.6, 1014.7, 1015, 1015.1, 1015.1, 
    1015, 1014.9, 1014.9, 1014.9, 1014.8, 1014.9, 1014.9, 1015.2, 1015.2, 
    1015.2, 1015.2, 1015.2, 1015.1, 1015, 1014.9, 1014.5, 1014.3, 1014.4, 
    1014.4, 1014.2, 1014.1, 1014.1, 1014, 1013.6, 1013.5, 1013.2, 1013.1, 
    1012.8, 1012.7, 1012.7, 1012.5, 1012.3, 1012.3, 1012.3, 1012.4, 1012.5, 
    1012.5, 1012.5, 1012.1, 1012, 1011.8, 1011.7, 1011.5, 1011.6, 1011.4, 
    1011.5, 1011.5, 1011.5, 1011.6, 1011.6, 1011.7, 1011.6, 1011.3, 1011.1, 
    1010.9, 1011, 1010.4, 1010.3, 1010.3, 1010.1, 1009.7, 1009.3, 1008.8, 
    1008.4, 1008, 1007.6, 1006.9, 1006.5, 1005.8, 1005.5, 1004.7, 1003.6, 
    1002.5, 1002, 1001.5, 1001.1, 1000.8, 1001, 1000.5, 1000.5, 1000.7, 
    1001.4, 1001.6, 1001.9, 1002.1, 1002.7, 1003.3, 1003.8, 1004.4, 1004.9, 
    1005.5, 1006.2, 1006.8, 1007.4, 1007.9, 1008.5, 1008.9, 1009.4, 1009.8, 
    1010.3, 1010.7, 1011.2, 1011.6, 1012, 1012.6, 1013, 1013.7, 1014.2, 
    1014.8, 1015, 1015.3, 1015.3, 1015.6, 1015.7, 1015.9, 1016, 1016.1, 
    1016.4, 1016.4, 1016.5, 1016.6, 1016.5, 1016.4, 1016.4, 1016.3, 1016.3, 
    1016.3, 1016.2, 1016.2, 1016.6, 1016.8, 1016.9, 1016.6, 1016.5, 1015.9, 
    1016, 1015.9, 1016, 1016.3, 1016.3, 1016.1, 1016.4, 1016.2, 1016.2, 
    1016.2, 1015.9, 1015.7, 1015.7, 1015.4, 1015.3, 1015.2, 1015.2, 1014.7, 
    1014.5, 1014.3, 1014.3, 1014.4, 1014.1, 1013.9, 1013.5, 1013.5, 1013.5, 
    1013.4, 1013.6, 1013.7, 1013.8, 1013.7, 1013.7, 1013.8, 1013.7, 1013.8, 
    1014.1, 1014.3, 1014.4, 1014.5, 1014.7, 1014.9, 1015, 1015.2, 1015.3, 
    1015.3, 1015.4, 1015.3, 1015.2, 1015.2, 1015, 1015.1, 1015.2, 1015, 1015, 
    1015.1, 1014.9, 1014.5, 1014.3, 1014, 1013.6, 1013.3, 1013.2, 1013, 
    1012.7, 1012.4, 1012.4, 1012.1, 1012.1, 1011.5, 1011, 1010.7, 1010.3, 
    1009.7, 1009.1, 1008.4, 1008.1, 1007.7, 1007.5, 1006.8, 1006.2, 1005.7, 
    1005.5, 1005.1, 1005, 1005, 1004.8, 1004.8, 1005, 1005.2, 1005.4, 1005.8, 
    1005.9, 1006.3, 1006.3, 1006.5, 1006.9, 1006.9, 1007.1, 1007.3, 1007.6, 
    1007.8, 1008, 1008.1, 1008, 1008.2, 1008, 1008, 1008, 1008, 1007.9, 
    1008.1, 1008, 1008, 1008, 1008, 1008, 1007.9, 1007.8, 1007.8, 1007.6, 
    1007.8, 1007.8, 1007.9, 1007.8, 1008, 1008.1, 1008.1, 1008.1, 1008, 1008, 
    1008, 1007.7, 1007.7, 1007.7, 1007.2, 1006.8, 1006.5, 1006.3, 1006, 
    1005.7, 1005.2, 1004.9, 1004.3, 1003.2, 1002.7, 1001.8, 1001.4, 1000.9, 
    1000.7, 1000.7, 1001, 1001.2, 1001.2, 1001.5, 1001.8, 1002.1, 1002.6, 
    1003.1, 1003.8, 1004.2, 1004.7, 1004.8, 1005.2, 1005.5, 1005.4, 1005.4, 
    1005.1, 1004.7, 1004.4, 1004, 1003.5, 1003.3, 1003, 1002.8, 1002.3, 
    1001.8, 1001.4, 1001.1, 1000.4, 999.7, 999.1, 998.6, 998.1, 997.7, 997.3, 
    997, 996.9, 996.5, 995.7, 995, 994.5, 994.2, 994.1, 993.9, 993.8, 993.9, 
    994, 994.1, 994.3, 994.4, 994.7, 994.9, 995.1, 995.1, 995.6, 995.8, 
    996.3, 996.6, 996.7, 996.8, 997, 997.1, 997.2, 997.1, 997, 996.8, 996.6, 
    996.2, 996.1, 996.2, 996.1, 996.2, 996.3, 996.4, 996.6, 997, 997.4, 
    997.7, 998.6, 999.3, 1000, 1000.6, 1001.4, 1001.9, 1002.5, 1002.9, 
    1003.6, 1004, 1004.4, 1004.7, 1005, 1005.2, 1005.4, 1005.3, 1005.4, 
    1005.2, 1004.4, 1003.7, 1002.7, 1001.7, 1000.6, 1000, 999.2, 998.5, 
    997.9, 997.7, 997.6, 997.7, 998, 998.5, 999.4, 999.9, 1000.4, 1001, 
    1001.5, 1001.6, 1001.9, 1002.2, 1002.7, 1003, 1003.2, 1003.4, 1003.4, 
    1003.3, 1003.4, 1003.5, 1003.4, 1003.3, 1003.2, 1003.1, 1003.1, 1002.9, 
    1003.1, 1003, 1003.2, 1003, 1002.8, 1002.7, 1002.5, 1002.6, 1002.9, 1003, 
    1003.2, 1003.3, 1003.5, 1003.6, 1003.8, 1004.1, 1004.4, 1004.5, 1004.8, 
    1005, 1005.2, 1005.4, 1005.6, 1005.9, 1006.1, 1006.2, 1006.5, 1006.5, 
    1006.4, 1006.1, 1006.1, 1006.2, 1006.5, 1006.4, 1006.8, 1006.7, 1006.4, 
    1006.2, 1005.8, 1005.8, 1005.6, 1005.4, 1005, 1005.2, 1005.1, 1005.5, 
    1005.7, 1005.4, 1005.8, 1006, 1006.3, 1005.9, 1005.7, 1005.8, 1005.6, 
    1005.2, 1005.2, 1005.4, 1005, 1004.9, 1004.7, 1004.3, 1004.1, 1004, 1004, 
    1004, 1004, 1004.1, 1003.8, 1004, 1004.2, 1004.1, 1004, 1003.8, 1003.9, 
    1004.1, 1004.5, 1004.5, 1004.1, 1003.8, 1004, 1004.2, 1004.2, 1004.1, 
    1003.8, 1003.3, 1003, 1002.5, 1002, 1002.1, 1002.1, 1001.9, 1001.7, 
    1001.9, 1002.1, 1002.2, 1001.8, 1001.6, 1001.5, 1001, 1000.6, 1000.2, 
    1000, 999.6, 999.4, 999.2, 998.9, 998.9, 998.8, 998.7, 998.7, 998.7, 
    998.6, 998.7, 998.7, 998.9, 998.7, 998.8, 999, 999.3, 999.4, 999.4, 
    999.8, 999.9, 999.9, 999.9, 1000.1, 1000, 1000.1, 1000.1, 1000.2, 1000.7, 
    1000.7, 1001.1, 1001.2, 1001.3, 1001.4, 1001.6, 1001.6, 1001.8, 1001.8, 
    1001.9, 1002.2, 1002.4, 1002.6, 1002.7, 1003, 1003.4, 1003.6, 1003.8, 
    1003.8, 1003.7, 1003.9, 1004.3, 1004.7, 1004.8, 1005.1, 1005.5, 1005.7, 
    1006, 1006.2, 1006.5, 1006.7, 1006.7, 1007, 1007.2, 1007.3, 1007.6, 
    1007.7, 1007.8, 1008, 1008, 1007.9, 1007.8, 1007.5, 1007.2, 1006.8, 
    1006.6, 1006.6, 1006.1, 1005.7, 1005.4, 1004.7, 1003.9, 1003.2, 1002.7, 
    1002.1, 1001.5, 1001.3, 1001.3, 1001.3, 1001.1, 1002.2, 1003.2, 1004.5, 
    1005.7, 1006.9, 1007.9, 1008.9, 1009.9, 1010.6, 1011.5, 1012.4, 1013.3, 
    1014, 1014.4, 1014.9, 1015.5, 1015.8, 1016.1, 1016.5, 1016.7, 1017.1, 
    1017.3, 1017.8, 1018, 1018.3, 1018.5, 1018.5, 1018.5, 1018.5, 1018.6, 
    1018.3, 1018.3, 1018.2, 1018.1, 1017.9, 1017.7, 1017.4, 1016.7, 1016.2, 
    1015.8, 1015.3, 1014.6, 1013.8, 1013.1, 1012.2, 1011.7, 1010.9, 1010, 
    1009.3, 1008.7, 1008.5, 1008.1, 1007.2, 1005.9, 1005, 1004.4, 1004, 
    1003.6, 1003.1, 1002.8, 1002.2, 1001.4, 1000.4, 999.4, 998, 996.8, 996.3, 
    995.7, 994.8, 994.1, 993.5, 993.2, 992.6, 992.5, 992.3, 992.2, 992.3, 
    992.5, 992.6, 992.8, 992.6, 993.2, 993.5, 993.8, 994.1, 994.3, 994.5, 
    994.8, 995, 995.1, 995.1, 995.2, 995.3, 995.3, 995.4, 995.3, 995.5, 
    995.5, 995.6, 995.6, 995.4, 995.4, 995.4, 995.5, 995.5, 995.3, 995.3, 
    995.3, 995.2, 994.8, 994.7, 994.5, 994.2, 994, 993.9, 993.5, 993.2, 993, 
    992.8, 992.5, 992.3, 991.8, 991.8, 991.6, 991.3, 991, 990.8, 991.1, 991, 
    990.8, 990.4, 990.4, 990.2, 990.2, 990.4, 990.6, 990.8, 991, 991.2, 
    991.9, 992.3, 992.7, 993.1, 993.3, 993.8, 994.7, 995, 995.9, 996.4, 
    997.2, 997.3, 998.2, 999.1, 999.7, 1000.5, 1001.1, 1001.6, 1002.4, 
    1002.9, 1003.7, 1004.1, 1004.6, 1005, 1005.7, 1006.3, 1006.8, 1007.3, 
    1007.9, 1008.4, 1009, 1009.4, 1009.6, 1010.1, 1010.5, 1010.7, 1011, 
    1011.2, 1011.5, 1011.6, 1012, 1012.5, 1012.8, 1013.1, 1013.4, 1013.5, 
    1013.9, 1013.9, 1014.1, 1014.4, 1014.6, 1014.8, 1015.1, 1015.3, 1015.5, 
    1015.5, 1015.6, 1015.7, 1015.6, 1015.9, 1015.6, 1015.9, 1015.8, 1016.1, 
    1016.1, 1016.2, 1016.2, 1016.2, 1016.1, 1016, 1015.8, 1015.8, 1015.7, 
    1015.7, 1015.6, 1015.6, 1015.6, 1015.7, 1015.6, 1015.4, 1015.3, 1015.2, 
    1015.2, 1015.1, 1015, 1014.9, 1015, 1015, 1015.2, 1015.1, 1015, 1015.1, 
    1015, 1015, 1015, 1015.1, 1014.9, 1014.7, 1014.6, 1014.8, 1014.9, 1014.9, 
    1015, 1014.9, 1014.5, 1014, 1013.8, 1013.6, 1013.5, 1013.2, 1013, 1012.9, 
    1013, 1013.2, 1013.2, 1013.1, 1012.6, 1012.2, 1011.8, 1011.2, 1010.9, 
    1010.3, 1009.8, 1009.8, 1009.5, 1009.3, 1008.7, 1008.3, 1008, 1007.8, 
    1007.7, 1007.6, 1007.5, 1007.5, 1007.3, 1007.3, 1007.4, 1007.3, 1007.2, 
    1007.1, 1006.5, 1006.1, 1005.6, 1005.3, 1005.1, 1005, 1005, 1005, 1004.6, 
    1004.7, 1004.6, 1004.1, 1003.6, 1003.2, 1002.6, 1002.3, 1002.6, 1002.8, 
    1002.9, 1002.9, 1002.7, 1002.6, 1002, 1001.9, 1001.4, 1001.3, 1001, 
    1000.9, 1000.7, 1000.7, 1000.5, 1000.2, 999.8, 1000, 1000, 1000.1, 
    1000.4, 1000.6, 1000.6, 1000.7, 1000.8, 1000.9, 1000.9, 1001.2, 1001.3, 
    1001.5, 1001.4, 1001.4, 1001.6, 1001.9, 1001.9, 1001.9, 1001.6, 1001.4, 
    1001.3, 1001.2, 1000.9, 1000.7, 1000.4, 1000, 999.4, 999, 998.6, 998.5, 
    998.6, 998.8, 999.4, 999.7, 1000.2, 1000.8, 1001.6, 1002.2, 1002.5, 
    1002.9, 1003.2, 1003.3, 1003.7, 1003.8, 1003.7, 1003.4, 1002.9, 1001.9, 
    1001, 1000.5, 1000.2, 999.3, 999.1, 998.9, 998.7, 999.2, 999.7, 1000.3, 
    1001, 1002, 1002.9, 1003.7, 1004.3, 1004.7, 1005.2, 1005.7, 1006.2, 
    1006.4, 1006.9, 1007, 1007.2, 1007.3, 1007, 1006.9, 1006.7, 1006.2, 
    1006.1, 1006.1, 1006, 1006.2, 1006.3, 1007, 1007.5, 1008.2, 1008.9, 
    1009.2, 1010, 1010.3, 1011.2, 1011.3, 1012.4, 1013.1, 1013.6, 1014, 
    1014.5, 1014.9, 1015.1, 1015.5, 1015.7, 1015.7, 1015.7, 1015.9, 1015.7, 
    1016.1, 1015.8, 1015.4, 1015.5, 1015, 1014.9, 1014.8, 1014.3, 1013.6, 
    1013.1, 1012.6, 1012.1, 1011.8, 1011.2, 1010.5, 1009.6, 1009, 1008.4, 
    1007.6, 1006.8, 1006.3, 1005.7, 1005.1, 1004.6, 1004.3, 1004.1, 1004.1, 
    1003.7, 1003.7, 1003.7, 1003.9, 1004.1, 1004.1, 1004, 1004, 1003.9, 
    1003.8, 1003.8, 1004, 1004, 1004.4, 1004.7, 1004.9, 1004.8, 1004.8, 
    1004.6, 1004.6, 1004.6, 1004.7, 1004.5, 1004.8, 1004.8, 1004.9, 1005.3, 
    1005.9, 1006.1, 1006.4, 1006.9, 1007.1, 1007.4, 1007.6, 1007.9, 1008, 
    1008, 1008.5, 1008.6, 1008.6, 1008.2, 1007.7, 1007.4, 1007, 1007.1, 
    1006.9, 1006.7, 1006.4, 1006.2, 1006, 1005.7, 1005.4, 1004.7, 1003.7, 
    1003.3, 1002.8, 1002.6, 1002.8, 1002.3, 1002.1, 1002.1, 1002, 1001.7, 
    1001.6, 1001.3, 1001.6, 1001.5, 1001.3, 1001.5, 1001.8, 1002.2, 1002.6, 
    1003.1, 1003.6, 1004.1, 1004, 1003.9, 1004, 1004.2, 1004, 1003.9, 1003.6, 
    1003.7, 1003.8, 1004.1, 1004.5, 1004.9, 1005.4, 1005.8, 1005.9, 1006, 
    1006.3, 1006.5, 1006.8, 1007.2, 1007.4, 1007.4, 1007.6, 1007.7, 1007.9, 
    1008.1, 1008.4, 1008.6, 1009.1, 1009.4, 1009.9, 1010.6, 1011.3, 1011.7, 
    1012.2, 1012.8, 1013.2, 1013.6, 1013.6, 1014, 1014.2, 1014.6, 1015, 
    1015.4, 1015.7, 1015.8, 1015.9, 1016.2, 1016.3, 1016.2, 1016.1, 1016.2, 
    1016.2, 1016.1, 1016.1, 1016.3, 1016.2, 1016, 1015.4, 1015.1, 1014.8, 
    1014.7, 1014.3, 1014.1, 1013.6, 1013.3, 1013.2, 1013, 1013.1, 1013.2, 
    1012.9, 1012.4, 1012.1, 1012, 1012, 1011.6, 1011.6, 1011.8, 1011.4, 
    1011.4, 1011.9, 1012.4, 1012.5, 1012.2, 1012, 1011.8, 1012.4, 1012.5, 
    1012.6, 1012.9, 1013.2, 1013.4, 1013.4, 1013.6, 1013.6, 1013.4, 1013.6, 
    1013.8, 1014, 1013.9, 1014, 1014.4, 1014.8, 1015, 1015.1, 1015.6, 1016.1, 
    1016.1, 1016.4, 1016.5, 1016.7, 1017.1, 1017.3, 1017.5, 1017.9, 1018.2, 
    1018.2, 1018.3, 1018.5, 1018.7, 1018.9, 1019.1, 1019.2, 1019.3, 1019.5, 
    1019.6, 1019.8, 1020, 1020.2, 1020.4, 1020.4, 1020.4, 1020.4, 1020.4, 
    1020.5, 1020.6, 1020.7, 1020.9, 1021, 1021.1, 1021.1, 1021.2, 1021.2, 
    1021.4, 1021.5, 1021.8, 1021.8, 1021.8, 1022.2, 1022.2, 1022.4, 1022.4, 
    1022.5, 1022.7, 1022.8, 1022.4, 1022.5, 1022.4, 1022.3, 1022.4, 1022.6, 
    1022.4, 1022.8, 1022.8, 1022.9, 1023.1, 1023.3, 1023.5, 1023.6, 1023.7, 
    1023.7, 1023.9, 1024.1, 1024.7, 1025, 1025.4, 1025.6, 1025.4, 1025.4, 
    1025.6, 1025.6, 1025.6, 1025.5, 1025.4, 1025.8, 1025.9, 1026.1, 1026.1, 
    1026.3, 1026.4, 1026.5, 1026.8, 1027.3, 1027.4, 1027.6, 1027.7, 1027.8, 
    1028.1, 1028.3, 1029, 1029.4, 1029.6, 1030, 1030.5, 1030.8, 1031.1, 
    1031.4, 1031.8, 1031.9, 1032.2, 1032.6, 1033, 1033.4, 1033.8, 1034, 
    1034.2, 1034.4, 1034.6, 1034.6, 1034.8, 1034.7, 1034.6, 1034.8, 1035, 
    1035, 1035.1, 1035.3, 1035.2, 1035.2, 1035.3, 1035.1, 1035.2, 1035, 
    1034.9, 1034.9, 1034.9, 1034.9, 1035, 1035, 1034.8, 1034.6, 1034.3, 
    1034.2, 1034.1, 1034, 1033.8, 1033.5, 1033.3, 1033.2, 1033.3, 1033.2, 
    1033.2, 1033, 1033, 1032.8, 1032.8, 1032.7, 1032.8, 1032.8, 1032.6, 
    1032.6, 1032.7, 1032.7, 1032.6, 1032.5, 1032.4, 1032.3, 1032.2, 1032, 
    1031.9, 1031.9, 1032, 1031.7, 1031.6, 1031.5, 1031.4, 1031.3, 1031.2, 
    1031.3, 1031.2, 1031, 1031, 1031.1, 1031, 1031.2, 1031.1, 1031.3, 1031.3, 
    1031.2, 1031.1, 1031, 1030.9, 1031.1, 1031.2, 1031.3, 1031.1, 1031.2, 
    1031.3, 1031.2, 1031.1, 1030.8, 1031, 1030.9, 1030.8, 1030.4, 1030.1, 
    1030.1, 1029.9, 1030.2, 1030.5, 1030.4, 1030.7, 1030.8, 1030.7, 1030.6, 
    1030.3, 1030.3, 1030.1, 1030.1, 1030.1, 1029.9, 1029.7, 1029.7, 1029.8, 
    1029.6, 1029.4, 1029.3, 1029.1, 1028.9, 1028.7, 1028.7, 1028.6, 1028.6, 
    1028.6, 1028.6, 1029, 1028.7, 1028.4, 1028.3, 1028, 1027.6, 1027.3, 
    1027.3, 1027.2, 1027, 1026.9, 1026.7, 1026.6, 1026.3, 1025.9, 1025.7, 
    1025.4, 1025.1, 1024.9, 1025.3, 1025.2, 1025, 1024.8, 1024.8, 1024.3, 
    1024.2, 1024.1, 1024.3, 1024, 1023.7, 1023.7, 1023.7, 1023.7, 1023.5, 
    1023.6, 1023.6, 1023.5, 1023.4, 1023.2, 1022.7, 1022.5, 1022.1, 1021.8, 
    1021.3, 1020.8, 1020.3, 1019.9, 1019.5, 1018.9, 1018.3, 1017.4, 1016.1, 
    1014.8, 1013.8, 1012.6, 1011.1, 1010, 1008.8, 1007.6, 1006.7, 1005.7, 
    1004.4, 1003.2, 1002.1, 1001.3, 1000.5, 1000.1, 999.3, 998.7, 998.1, 
    997.1, 996.3, 995.7, 995, 995.2, 995.4, 995.4, 995.2, 995.2, 995.5, 
    996.1, 996.6, 997.2, 997.6, 998.1, 998.3, 998.5, 998.3, 997.8, 997.3, 
    996.6, 996.3, 996, 995.5, 994.9, 994.1, 993, 992, 990.8, 990.2, 990.1, 
    990.3, 990.3, 990.5, 991.2, 991.9, 992.5, 993.1, 993.4, 994.1, 994.9, 
    995.5, 996.2, 996.7, 997.4, 998.1, 999, 999.5, 1000, 1000.5, 1000.9, 
    1001.6, 1001.8, 1002, 1002.1, 1002.6, 1002.7, 1002.7, 1003.2, 1003.5, 
    1003.8, 1004.4, 1004.7, 1005, 1005.3, 1005.6, 1005.6, 1006.1, 1006.3, 
    1006.3, 1006.6, 1006.9, 1007.2, 1007.5, 1007.7, 1008.1, 1008.1, 1008.1, 
    1008.3, 1008.3, 1008.3, 1008.4, 1008.5, 1008.9, 1008.9, 1009, 1009.1, 
    1009, 1008.9, 1009.1, 1009.6, 1009.5, 1009.9, 1010.2, 1010.8, 1010.8, 
    1011, 1011.1, 1011.2, 1011.3, 1011.7, 1011.5, 1011.6, 1011.5, 1011.7, 
    1011.5, 1011.5, 1011.8, 1011.4, 1011.3, 1011.3, 1011, 1010.9, 1010.7, 
    1010.7, 1010.4, 1010.3, 1010.4, 1010.3, 1010.5, 1010.8, 1011, 1011.2, 
    1011.5, 1011.8, 1012.1, 1011.9, 1012.2, 1012.1, 1012.6, 1012.6, 1012.6, 
    1012.9, 1013.3, 1013.5, 1013.8, 1013.7, 1014.2, 1014.3, 1014.6, 1014.8, 
    1015.2, 1015.5, 1015.7, 1016.1, 1016.3, 1016.3, 1016.5, 1016.5, 1016.5, 
    1016.5, 1016.4, 1016.5, 1016.5, 1016.5, 1016.4, 1016.4, 1016.3, 1016.1, 
    1016.1, 1016, 1015.7, 1015.4, 1015.3, 1015.3, 1015.4, 1015.4, 1015.4, 
    1015.5, 1015.4, 1015.3, 1015.2, 1014.9, 1014.4, 1014.3, 1014, 1013.6, 
    1013.3, 1013, 1012.5, 1012.2, 1011.9, 1011.5, 1011.3, 1010.7, 1010.1, 
    1009.7, 1009.4, 1009, 1008.6, 1008.2, 1008.1, 1007.9, 1007.6, 1007.3, 
    1006.8, 1006.3, 1005.7, 1005.4, 1005.2, 1004.9, 1004.5, 1004.3, 1004, 
    1003.4, 1003, 1002.5, 1002.1, 1001.5, 1001, 1000.5, 999.9, 999.3, 998.6, 
    998, 997.6, 997.1, 996.2, 995.5, 995.2, 994.9, 994.6, 994.3, 994.2, 
    994.3, 994.3, 994.6, 994.6, 994.9, 995, 995.2, 995.7, 996.1, 996.2, 
    996.8, 997.4, 998.2, 999.1, 1000.1, 1001.1, 1002.5, 1003.6, 1004.9, 
    1006.1, 1006.9, 1007.8, 1008.7, 1009.6, 1010.2, 1011.1, 1011.4, 1012, 
    1012.5, 1012.9, 1013.1, 1012.7, 1013, 1012.7, 1012.4, 1012.2, 1012, 
    1012.1, 1011.6, 1011.4, 1011.4, 1011.7, 1011.9, 1011.8, 1012.1, 1012.5, 
    1013.2, 1014, 1015.1, 1016.3, 1017.4, 1019, 1020.3, 1021.5, 1022.1, 
    1023.1, 1023.8, 1024.3, 1024.3, 1024.7, 1024.7, 1024.5, 1024.1, 1024, 
    1024.1, 1023.6, 1023.2, 1022.5, 1021.8, 1021.1, 1020.5, 1019.9, 1019.2, 
    1018.8, 1018.4, 1018.2, 1017.8, 1017.3, 1016.7, 1016.1, 1015.6, 1014.9, 
    1014.2, 1013.8, 1013.2, 1012.4, 1012, 1011.5, 1011.1, 1011.1, 1011.1, 
    1011.1, 1010.9, 1010.8, 1010.8, 1010.9, 1011.4, 1012, 1012.7, 1013.7, 
    1014.9, 1015.3, 1015.8, 1016.3, 1016.8, 1017.2, 1017.7, 1018.2, 1018.4, 
    1018.7, 1019.3, 1019.8, 1020.3, 1020.6, 1020.8, 1020.8, 1021, 1021, 
    1021.2, 1021.1, 1021, 1020.8, 1020.9, 1020.9, 1020.8, 1020.4, 1020, 
    1019.7, 1019.5, 1019.2, 1018.9, 1018.4, 1018, 1017.7, 1017.3, 1017.1, 
    1016.8, 1016.2, 1015.5, 1014.8, 1014.4, 1013.7, 1013, 1012.5, 1011.8, 
    1011.4, 1011, 1010.6, 1010.2, 1009.9, 1009.4, 1009.2, 1008.8, 1008.6, 
    1008, 1007.8, 1007.6, 1007.6, 1007.5, 1007.6, 1007.6, 1007.9, 1007.8, 
    1007.7, 1007.7, 1007.7, 1008, 1008.5, 1008.5, 1008.7, 1008.9, 1009.4, 
    1009.6, 1009.8, 1010.2, 1010.5, 1010.5, 1010.9, 1011.1, 1011.5, 1011.8, 
    1012, 1012.6, 1012.7, 1013.1, 1013.6, 1014, 1014.3, 1014.7, 1015.1, 
    1015.5, 1015.7, 1015.8, 1016.1, 1016.4, 1016.7, 1017.1, 1017.2, 1017.4, 
    1017.4, 1017.5, 1017.6, 1017.8, 1017.9, 1018.1, 1018.1, 1018, 1018.3, 
    1018.4, 1018.6, 1018.8, 1018.8, 1018.8, 1018.8, 1018.9, 1019, 1019.2, 
    1019.3, 1019.5, 1019.8, 1019.8, 1019.7, 1019.7, 1019.6, 1019.5, 1019.5, 
    1019.2, 1019, 1018.7, 1018.5, 1018.2, 1018.1, 1017.9, 1017.6, 1017.3, 
    1017, 1016.5, 1016.1, 1015.8, 1015.5, 1015, 1014.5, 1014.1, 1013.7, 
    1013.3, 1012.8, 1012.4, 1012, 1011.5, 1011.2, 1010.8, 1010.6, 1010.4, 
    1010.2, 1010.1, 1010.1, 1010, 1009.4, 1009.1, 1008.9, 1008.9, 1008.5, 
    1007.9, 1007.4, 1007, 1006.8, 1006.6, 1006.6, 1006.5, 1006.3, 1006.3, 
    1006, 1005.7, 1005.7, 1005.6, 1005.6, 1005.3, 1005.3, 1005.2, 1005.2, 
    1005.3, 1005.3, 1005.1, 1004.8, 1004.6, 1004.3, 1003.9, 1003.8, 1003.7, 
    1003.3, 1003.3, 1003, 1002.8, 1002.8, 1002.6, 1002.4, 1002.4, 1002.3, 
    1002.2, 1002.1, 1002.1, 1002.1, 1002.3, 1002.6, 1002.9, 1002.9, 1003, 
    1003.1, 1003.1, 1003.3, 1003.4, 1003.5, 1003.5, 1003.7, 1003.7, 1003.7, 
    1003.9, 1004, 1003.9, 1003.9, 1003.9, 1003.9, 1003.8, 1003.6, 1003.6, 
    1003.8, 1003.9, 1004.2, 1004.5, 1004.6, 1004.5, 1004.7, 1004.7, 1004.5, 
    1004.5, 1004.3, 1004.2, 1004.2, 1004.1, 1004, 1003.9, 1003.7, 1003, 
    1002.7, 1002.4, 1001.9, 1001.5, 1001.3, 1001.3, 1001.3, 1001.4, 1001.5, 
    1001.6, 1001.6, 1001.8, 1001.8, 1001.9, 1002.1, 1003.1, 1002.7, 1003, 
    1003, 1003.2, 1003.1, 1003.4, 1003.5, 1003.6, 1003.7, 1003.7, 1003.6, 
    1003.6, 1003.5, 1003.5, 1003.4, 1003.4, 1003.5, 1003.6, 1003.7, 1003.6, 
    1003.5, 1003.4, 1003.3, 1003.3, 1003.3, 1003.2, 1003.1, 1003, 1003, 
    1002.9, 1002.8, 1002.8, 1002.6, 1002.5, 1002.2, 1002.1, 1001.9, 1001.8, 
    1001.7, 1001.7, 1001.7, 1001.7, 1001.8, 1001.8, 1001.8, 1001.7, 1001.7, 
    1001.6, 1001.4, 1001.5, 1001.5, 1001.4, 1001.4, 1001.3, 1001.2, 1001.1, 
    1001, 1000.9, 1000.8, 1000.7, 1000.5, 1000.5, 1000.5, 1000.8, 1000.9, 
    1001.1, 1001, 1001.1, 1001.4, 1001.5, 1001.4, 1001.5, 1001.6, 1001.7, 
    1001.9, 1002.1, 1002.3, 1002.4, 1002.4, 1002.7, 1002.8, 1003, 1003, 
    1003.3, 1003.5, 1003.6, 1003.9, 1004.4, 1004.5, 1004.8, 1005, 1005, 
    1005.5, 1005.5, 1005.5, 1005.4, 1005.7, 1005.6, 1005.9, 1005.9, 1005.8, 
    1005.7, 1005.8, 1005.8, 1005.5, 1005.1, 1005, 1004.7, 1004.3, 1004.2, 
    1004.2, 1004.2, 1004.1, 1004.2, 1004.1, 1004.2, 1004.1, 1004, 1004.3, 
    1004.6, 1004.8, 1005.3, 1005.7, 1006.1, 1006.5, 1006.8, 1007.4, 1007.9, 
    1008, 1008.3, 1008.6, 1008.5, 1008.6, 1008.7, 1008.9, 1009.2, 1009.4, 
    1009.5, 1009.9, 1010.2, 1010.2, 1010.1, 1010.1, 1009.9, 1009.9, 1009.9, 
    1009.7, 1009.7, 1009.8, 1009.8, 1009.6, 1009.8, 1009.7, 1009.7, 1009.6, 
    1009.3, 1009, 1008.7, 1008.7, 1008.6, 1008.7, 1008.9, 1008.9, 1008.9, 
    1008.9, 1008.4, 1008.2, 1008.2, 1007.9, 1007.6, 1007.5, 1007.3, 1007.2, 
    1007.3, 1007.1, 1007, 1006.8, 1006.5, 1006.1, 1005.4, 1004.8, 1004.3, 
    1003.9, 1003.4, 1003.2, 1002.9, 1002.4, 1002.2, 1002, 1001.6, 1001, 
    1000.1, 999.3, 999, 998.6, 997.8, 997.4, 997, 996.5, 996, 995.4, 995, 
    994.7, 994.5, 994.2, 993.9, 993.2, 992.9, 992.6, 992.2, 992.1, 991.8, 
    991.5, 991.6, 991.7, 991.5, 991.6, 991.9, 992.2, 992.6, 992.8, 993.2, 
    993.6, 993.9, 994, 994.1, 994.6, 994.8, 995, 995.2, 995.4, 995.7, 995.9, 
    995.9, 995.7, 995.6, 995.5, 995, 994.6, 994.2, 993.5, 992.6, 991.5, 
    990.8, 989.8, 988.7, 988.4, 987.2, 985.5, 984, 982.7, 981.9, 981.2, 
    980.5, 979.8, 979.1, 978.8, 978.9, 978.9, 978.8, 978.6, 978.3, 978.1, 
    977.8, 977.6, 977, 976.9, 976.7, 977, 977.2, 977.6, 977.9, 977.7, 978, 
    977.9, 977.8, 977.9, 978.3, 978.4, 979, 979.9, 980.6, 981.5, 981.9, 
    982.4, 982.6, 983, 983.2, 983.5, 983.7, 983.7, 983.7, 983.5, 983.4, 
    983.2, 983.4, 983, 982.8, 982.7, 982.7, 982.5, 982.2, 982.1, 981.8, 
    981.9, 981.9, 981.8, 981.6, 981.5, 981.3, 980.9, 981, 981.5, 981.4, 
    981.2, 981.2, 981.6, 982.6, 983.6, 984.9, 986.1, 986.9, 987.8, 988.5, 
    989.3, 990.2, 990.7, 991.6, 992.4, 993.2, 994.1, 994.8, 995.4, 996.3, 
    996.9, 997.6, 998.1, 998.6, 999.1, 999.6, 1000.1, 1000.4, 1000.9, 1001.1, 
    1001.3, 1001.4, 1001.6, 1001, 1000.9, 1000.8, 1000.8, 1000.5, 1000.6, 
    1000.5, 1000, 999.9, 999.6, 999.8, 999.6, 998.6, 998.2, 997.8, 997.1, 
    996.4, 996, 995.4, 995.4, 995.1, 994.8, 994.4, 994.2, 994, 993.6, 993.2, 
    993.1, 992.9, 992.7, 992.5, 992.5, 992.2, 992, 991.8, 991.5, 991.1, 
    990.6, 990.2, 989.6, 989, 988.8, 988.5, 988.3, 988, 987.7, 987.7, 988, 
    988.4, 988.5, 988.7, 989.2, 989.5, 989.8, 990.5, 991, 991.6, 992.1, 
    992.6, 992.7, 992.8, 993.1, 993.4, 994, 994.5, 994.8, 995.2, 995.4, 
    995.8, 996.1, 996.1, 996.2, 996, 995.8, 995.8, 995.6, 995.5, 995.3, 
    995.4, 995.3, 995.1, 994.7, 994.4, 994.1, 994, 993.8, 993.3, 993.2, 
    993.1, 993.4, 993.5, 993.6, 993.9, 994.1, 994.1, 994, 994.4, 994.6, 
    994.9, 995.5, 996.3, 997.1, 997.8, 998.9, 999.5, 999.9, 1000.2, 1000.9, 
    1001.3, 1001.6, 1002.2, 1002.7, 1002.8, 1003.5, 1003.9, 1004.5, 1004.7, 
    1005.1, 1005.6, 1005.9, 1006.2, 1006.3, 1006.5, 1006.8, 1006.8, 1007.3, 
    1007.7, 1007.4, 1007.5, 1007.2, 1006.9, 1005.9, 1005.2, 1004.3, 1003.2, 
    1002.6, 1001.5, 1000.6, 999.7, 998.4, 996.8, 995.3, 993.5, 989.8, 988.7, 
    985.7, 981.5, 978, 973.8, 970.5, 968.1, 966, 964.3, 963, 962, 961.3, 
    960.5, 959.7, 959.6, 959.6, 959.8, 960.5, 961.3, 962.2, 962.9, 963.6, 
    964.6, 965.4, 966, 967, 967.9, 969.1, 969.5, 970.5, 971.4, 972, 972.5, 
    973.1, 973.6, 973.9, 973.8, 973.8, 973.9, 974.1, 974, 974.4, 974.2, 
    974.4, 974.2, 974.3, 974.8, 974.7, 975.1, 975.7, 976, 976.9, 977.1, 
    977.5, 978.1, 978.4, 979.1, 979.7, 980.3, 981, 981.6, 982, 982.7, 983.3, 
    984.1, 984.8, 985.4, 985.9, 986.3, 986.5, 986.6, 987, 987, 987.8, 988.2, 
    988.3, 988.4, 989, 989.4, 989.7, 989.7, 990.2, 990.3, 990.5, 990.6, 
    990.7, 990.9, 991, 991, 991.1, 991.1, 990.8, 990.5, 990.3, 990.1, 989.9, 
    989.7, 989.6, 989.5, 989.4, 989.5, 989.8, 989.9, 990.1, 990.1, 990.4, 
    990.9, 991.2, 991.4, 991.7, 992, 992.2, 992.6, 992.8, 993, 993.5, 993.5, 
    993.9, 994.2, 994.7, 995.3, 995.4, 995.7, 996.1, 996.1, 996.7, 997.1, 
    997.1, 997.2, 997.2, 997.5, 997.9, 998.1, 998.3, 998.5, 998.8, 999.3, 
    999.5, 999.8, 1000.1, 1000.5, 1000.6, 1000.6, 1000.9, 1000.8, 1000.6, 
    1000.5, 1000.6, 1000.7, 1000.9, 1001.1, 1001.4, 1001.4, 1001, 1000.8, 
    1000.4, 1000.2, 1000.1, 999.4, 998.8, 998, 997.6, 997.3, 996.6, 996, 995, 
    994.5, 993.8, 993.2, 992.3, 991.7, 991.2, 990.1, 989.6, 988.4, 987.6, 
    986.4, 984.8, 983.8, 982.6, 982.2, 981.5, 981.5, 981.7, 982.2, 981.7, 
    981.5, 981.6, 981.6, 981.6, 981.1, 981.5, 981.7, 981.6, 981.3, 980.5, 
    979.9, 978.7, 979, 978.1, 978.8, 979.6, 980.9, 982.7, 984.4, 986, 987.2, 
    987.7, 988.3, 989, 989.5, 989.7, 989.8, 989.7, 989.7, 990, 990.5, 991, 
    991.8, 992.5, 993.3, 994.7, 995.6, 996.6, 997.2, 998, 998.4, 999.6, 
    1000.4, 1001.3, 1002.1, 1002.7, 1003.4, 1004.1, 1004.5, 1005.2, 1005.3, 
    1005.6, 1005.3, 1005.5, 1005.9, 1006.2, 1006.2, 1006.4, 1006.6, 1006.9, 
    1006.8, 1007.3, 1007.6, 1007.7, 1007.7, 1007.9, 1008.1, 1008.5, 1008.6, 
    1008.7, 1008.7, 1008.8, 1009.1, 1009, 1008.9, 1008.9, 1008.6, 1008.1, 
    1007.8, 1007.3, 1006.7, 1006.6, 1006.4, 1005.9, 1005.5, 1005.6, 1005.2, 
    1004.9, 1004.7, 1004.5, 1004.2, 1004.1, 1003.9, 1004, 1004.2, 1004, 
    1004.1, 1003.9, 1003.4, 1002.8, 1002.2, 1001.9, 1001.5, 1000.9, 1000.4, 
    1000.2, 1000, 999.9, 999.8, 999.4, 999.2, 999.1, 999.3, 999.6, 999.8, 
    1000, 1000.5, 1000.9, 1001.3, 1001.7, 1002.1, 1002.5, 1002.8, 1003.3, 
    1003.8, 1004.2, 1004.4, 1004.8, 1004.8, 1005.2, 1005.6, 1005.9, 1006, 
    1005.9, 1005.8, 1005.8, 1005.8, 1005.7, 1005.4, 1004.9, 1004.7, 1004.4, 
    1004, 1003.8, 1003.5, 1003.1, 1002.5, 1002, 1001.7, 1001.4, 1000.8, 
    1000.3, 999.7, 999.2, 999.2, 998.6, 998.3, 997.8, 997.4, 996.7, 996.3, 
    995.7, 995.3, 994.9, 994.5, 994, 993.4, 992.9, 992.2, 991.8, 991.7, 
    991.4, 991.2, 990.8, 990.4, 989.7, 989.6, 989.6, 989.6, 989.7, 989.4, 
    989.3, 989.1, 989, 989.3, 989.6, 989.4, 989.7, 990, 989.8, 990, 990.6, 
    990.9, 990.8, 991.5, 991.9, 992.5, 993, 993.4, 994, 994.6, 994.9, 995.4, 
    995.9, 996.4, 997, 997.5, 997.7, 997.8, 997.8, 998, 998.1, 998.6, 999, 
    999.4, 999.7, 1000, 1000.6, 1000.6, 1000.7, 1000.9, 1000.4, 1000.5, 
    1000.9, 1000.8, 1000.7, 1000.3, 1000, 999.6, 999.5, 999.1, 998.9, 998.5, 
    997.9, 997.1, 996.4, 995.5, 994.8, 994.4, 994, 993.5, 992.8, 992.4, 
    991.8, 991.4, 991.2, 990.8, 990.4, 990.1, 989.8, 989.6, 989.5, 989.6, 
    989.7, 989.6, 989.6, 989.8, 989.9, 990.1, 990.1, 990.1, 990.2, 990.4, 
    990.7, 991.1, 991.4, 991.6, 991.5, 991.9, 992, 992.2, 992.4, 992.3, 
    992.5, 992.9, 993.3, 993.8, 993.9, 994.1, 994.4, 994.5, 994.5, 994.6, 
    994.8, 994.7, 994.6, 994.9, 995.2, 995.5, 996.1, 996.5, 996.5, 996.8, 
    996.8, 997.3, 997.5, 997.5, 997.7, 998.5, 999.3, 1000.1, 1000.6, 1001.4, 
    1002.1, 1002.3, 1002.8, 1003.2, 1003.5, 1004, 1004, 1004.3, 1004.6, 
    1005.2, 1005.7, 1005.9, 1006, 1006.4, 1006.6, 1006.6, 1006.5, 1006.5, 
    1006.4, 1006.4, 1006.7, 1006.7, 1006.9, 1006.8, 1006.7, 1006.7, 1007, 
    1007.1, 1007.1, 1007.2, 1007.3, 1007.5, 1007.9, 1008.2, 1008.1, 1008.3, 
    1008.4, 1008.6, 1008.6, 1008.8, 1008.7, 1008.7, 1008.7, 1008.7, 1008.9, 
    1009, 1009.2, 1009.2, 1009, 1008.9, 1008.8, 1008.6, 1008.5, 1008.4, 
    1008.3, 1008.4, 1008.4, 1008.6, 1008.7, 1009.2, 1009.2, 1009.3, 1009.7, 
    1009.9, 1009.7, 1009.4, 1009.8, 1010, 1010.3, 1010.1, 1010.3, 1010.4, 
    1010.4, 1010.6, 1010.7, 1010.9, 1010.9, 1010.6, 1010.6, 1010.8, 1011, 
    1011, 1010.9, 1010.5, 1010.3, 1010.4, 1010.3, 1010.2, 1010.2, 1010.4, 
    1010.7, 1010.8, 1010.9, 1011.4, 1011.5, 1011.6, 1012, 1012.1, 1012.3, 
    1012.3, 1012.3, 1012.1, 1012.2, 1012.2, 1012.3, 1012.1, 1012, 1012.1, 
    1012.3, 1012, 1012.1, 1011.8, 1011.5, 1011.3, 1011, 1010.8, 1010.7, 
    1010.7, 1010.7, 1010.3, 1010.1, 1010, 1010.1, 1009.8, 1009.6, 1009.2, 
    1008.7, 1008.4, 1008, 1007.6, 1007, 1006.5, 1005.7, 1005, 1004.2, 1003.2, 
    1002.1, 1001, 1000, 999.3, 998.6, 998, 997.2, 996.4, 995.6, 995, 994.7, 
    994.3, 994.4, 994.9, 994.9, 995.2, 995.1, 995, 995.2, 995.3, 995.3, 
    995.6, 995.5, 995.2, 995, 995.4, 995.7, 995.9, 996, 996, 996.2, 996.2, 
    996.5, 996.5, 996.7, 997.1, 997.3, 998.1, 999.1, 999.9, 1000.8, 1001.5, 
    1002.6, 1003.4, 1004.2, 1005, 1005.6, 1006.2, 1006.7, 1007.1, 1007.7, 
    1008, 1008.3, 1008.7, 1008.9, 1009.3, 1009.4, 1009.9, 1010.2, 1010, 1010, 
    1009.8, 1009.8, 1009.7, 1009, 1008.4, 1008, 1007.4, 1007.1, 1007, 1006.8, 
    1006.3, 1005.5, 1004.4, 1003.4, 1002.9, 1002.9, 1003.1, 1003.3, 1003.5, 
    1003.8, 1003.7, 1003.2, 1002.7, 1003.4, 1003.4, 1003.4, 1003.5, 1002.5, 
    1002.7, 1002.7, 1002.5, 1002.1, 1001.7, 1001, 1000.5, 999.8, 999.4, 
    998.6, 998.1, 997.9, 997.5, 996.7, 995.8, 995.3, 994.5, 993.6, 992.7, 
    992, 991.1, 990.1, 989.8, 989, 988, 987.3, 986.4, 985.4, 985.1, 984.5, 
    983.5, 983.2, 983.7, 984.4, 984.4, 984.7, 984.4, 984.3, 983.8, 983.3, 
    983, 982.6, 981.6, 980.9, 979.5, 978.4, 977.8, 977.3, 977.2, 976.5, 
    975.2, 974.8, 974.8, 974.5, 974.8, 974.9, 975.2, 975.3, 975.8, 975.5, 
    975.2, 974.9, 974.7, 975.2, 975.8, 977, 978, 979.6, 980.8, 981.6, 982.8, 
    984, 984.6, 985.3, 986.6, 988, 989.4, 990.5, 991.5, 992.4, 993.2, 994.4, 
    995.6, 996.4, 997.5, 998.4, 999.3, 1000, 1000.5, 1001.1, 1001.1, 1001.3, 
    1001.2, 1001.1, 1001.4, 1001.6, 1001.9, 1002.2, 1002.6, 1002.5, 1002.5, 
    1002.8, 1002.7, 1002.7, 1002.6, 1002.5, 1002.5, 1002.5, 1002.5, 1002.7, 
    1002.3, 1001.9, 1001.7, 1001.5, 1001.4, 1001.4, 1001.6, 1001.8, 1002, 
    1002.1, 1002.2, 1002.7, 1002.8, 1003, 1002.7, 1002.8, 1002.7, 1002.5, 
    1002.3, 1002.2, 1002.2, 1001.9, 1001.8, 1001.6, 1001.6, 1001.6, 1001.5, 
    1001.5, 1001.6, 1001.5, 1001.5, 1001.5, 1001.9, 1002, 1002.3, 1002.3, 
    1002.2, 1002.3, 1002.3, 1002.5, 1002.5, 1002.3, 1002.1, 1002.4, 1002.6, 
    1002.8, 1002.9, 1003.1, 1003.3, 1003.5, 1003.5, 1003.6, 1003.8, 1003.6, 
    1003.9, 1003.9, 1004, 1004.2, 1004.5, 1004.6, 1004.9, 1005, 1005.7, 1006, 
    1006.1, 1006.2, 1006.2, 1006.1, 1006.4, 1006.6, 1006.9, 1007.2, 1007.3, 
    1007.4, 1007.3, 1007.6, 1008.3, 1008.5, 1008.6, 1008.6, 1008.8, 1009, 
    1008.8, 1008.5, 1008.5, 1008.9, 1008.6, 1008.4, 1008.7, 1008.4, 1008.5, 
    1008.4, 1008.3, 1008.8, 1009, 1008.9, 1008.9, 1009, 1009.3, 1009.5, 
    1009.6, 1009.6, 1009.6, 1009.8, 1010.1, 1010.2, 1010.7, 1011, 1011.5, 
    1011.7, 1012, 1012.3, 1012.6, 1012.6, 1012.7, 1013.2, 1013.1, 1013.5, 
    1013.6, 1014.3, 1014.6, 1014.9, 1014.8, 1014.6, 1014.6, 1014.4, 1014.6, 
    1014.5, 1014.4, 1014.7, 1014.6, 1014.8, 1014.8, 1014.4, 1014.1, 1014.2, 
    1013.7, 1013.2, 1013.5, 1013.4, 1013.1, 1012.9, 1012.9, 1012.6, 1012.3, 
    1011.8, 1011.4, 1010.9, 1010.5, 1010.2, 1009.8, 1009.7, 1009.6, 1009.4, 
    1009.3, 1009.2, 1008.7, 1008.5, 1008.2, 1007.9, 1007.5, 1007.4, 1007.1, 
    1006.7, 1006.9, 1006.6, 1006.6, 1006.6, 1006.3, 1005.8, 1005.6, 1005.4, 
    1005.4, 1005.2, 1005.1, 1005, 1004.7, 1004.8, 1004.9, 1005.1, 1005.1, 
    1004.9, 1004.8, 1005.1, 1004.9, 1005.5, 1005.6, 1005.9, 1006.1, 1006, 
    1006.3, 1006.5, 1006.6, 1006.5, 1006.8, 1006.6, 1006.9, 1006.6, 1006.7, 
    1006.6, 1006.7, 1006.8, 1006.6, 1006.6, 1006.4, 1005.9, 1005.8, 1005.6, 
    1005.3, 1005, 1004.9, 1004.9, 1004.6, 1004.5, 1004.8, 1004.9, 1005, 
    1004.4, 1004.1, 1004.1, 1004.3, 1004.5, 1004.6, 1004.7, 1004.9, 1005.2, 
    1005.5, 1006, 1006.2, 1006.6, 1007, 1007.2, 1007.6, 1007.9, 1008.2, 
    1008.2, 1008.7, 1009.3, 1009.7, 1010, 1010.2, 1010.5, 1010.7, 1010.8, 
    1011.2, 1011.4, 1011.5, 1011.9, 1012.1, 1012.4, 1012.6, 1012.9, 1013.4, 
    1013.6, 1013.8, 1014.2, 1014.5, 1014.6, 1014.8, 1015.3, 1015.6, 1016.1, 
    1016.6, 1017, 1017.3, 1017.5, 1017.6, 1017.8, 1017.8, 1017.9, 1018.2, 
    1018.7, 1018.9, 1019.2, 1019.5, 1019.6, 1019.9, 1020.3, 1020.3, 1020.3, 
    1020.3, 1020.6, 1020.6, 1020.8, 1021.1, 1021.7, 1022.1, 1022.4, 1022.6, 
    1022.9, 1022.8, 1023, 1023, 1023, 1023.1, 1023.1, 1023.1, 1023.2, 1023.2, 
    1022.9, 1022.4, 1022, 1021.5, 1021, 1020.4, 1019.8, 1019.3, 1018.6, 1018, 
    1017.7, 1017.7, 1017.4, 1017.2, 1016.9, 1016.6, 1016.5, 1016.4, 1016.3, 
    1016.4, 1016.7, 1016.8, 1017.2, 1017.4, 1017.7, 1018, 1018.2, 1018.3, 
    1018.3, 1018.4, 1018.5, 1018.6, 1018.6, 1018.6, 1019, 1019.4, 1019.5, 
    1019.5, 1019.2, 1019, 1018.6, 1018.5, 1018.4, 1018.3, 1018.1, 1018.5, 
    1018.6, 1018.7, 1018.9, 1018.8, 1018.5, 1018.4, 1017.8, 1017.5, 1017.5, 
    1017.3, 1017.2, 1017.1, 1017.1, 1017.4, 1017.3, 1017.3, 1017.2, 1017.1, 
    1016.9, 1016.6, 1016.3, 1015.9, 1015.9, 1015.9, 1015.7, 1015.5, 1015.2, 
    1015, 1014.9, 1014.8, 1014.6, 1014.4, 1014.3, 1014.4, 1014.1, 1014.1, 
    1014.3, 1014.7, 1014.8, 1014.9, 1015, 1015.3, 1015.5, 1015.5, 1015.7, 
    1015.8, 1016, 1016.3, 1016.4, 1016.5, 1016.7, 1016.7, 1016.9, 1017, 
    1017.1, 1017.4, 1017.3, 1017.4, 1017.5, 1017.5, 1017.9, 1018, 1018.1, 
    1018.2, 1018.4, 1018.8, 1019.1, 1019.1, 1019.4, 1019.4, 1019.5, 1019.7, 
    1019.9, 1020.1, 1020.4, 1020.5, 1020.4, 1020.5, 1020.8, 1020.8, 1020.7, 
    1020.8, 1021, 1021.3, 1021.4, 1021.8, 1021.9, 1022.2, 1022.3, 1022.4, 
    1022.4, 1022.2, 1022.2, 1022.3, 1022.3, 1022.3, 1022.4, 1022.6, 1022.7, 
    1023, 1022.8, 1022.9, 1023, 1022.9, 1022.8, 1022.7, 1022.7, 1022.7, 
    1022.8, 1022.9, 1023.1, 1023.4, 1023.5, 1023.5, 1023.6, 1023.7, 1023.8, 
    1023.9, 1024.1, 1024.4, 1024.6, 1024.9, 1025.1, 1025.3, 1025.2, 1025.3, 
    1025.3, 1025.2, 1025.1, 1025.2, 1025.1, 1025, 1025.2, 1025.2, 1025.1, 
    1025.3, 1025.1, 1025.1, 1025, 1024.5, 1024.1, 1024.1, 1024, 1024.2, 
    1023.7, 1023.7, 1023.4, 1023.3, 1023.3, 1023, 1022.2, 1022, 1021.2, 
    1021.1, 1021.1, 1020.8, 1020.5, 1020.2, 1019.9, 1019.6, 1018.9, 1018, 
    1017.3, 1016.5, 1015.7, 1015, 1014.5, 1013.4, 1012.1, 1011.4, 1011.1, 
    1010.5, 1010, 1009.1, 1008.3, 1007.7, 1006.7, 1006.3, 1005.9, 1006, 1006, 
    1005.9, 1005.9, 1005.8, 1006.1, 1005.9, 1006.1, 1006.2, 1006.4, 1006.5, 
    1006.5, 1006.8, 1007.2, 1007.4, 1007.5, 1007.7, 1007.9, 1007.3, 1008, 
    1008, 1008, 1008, 1008.1, 1008.3, 1008.6, 1008.8, 1009.1, 1009.1, 1009.1, 
    1009.1, 1009.2, 1009.3, 1009.5, 1009.7, 1010, 1010.4, 1010.9, 1011.4, 
    1011.9, 1012.3, 1012.7, 1013.3, 1013.5, 1013.8, 1013.8, 1013.8, 1014, 
    1014.5, 1014.9, 1015.4, 1015.8, 1016.4, 1016.7, 1016.9, 1017, 1017.3, 
    1017.5, 1017.8, 1018.2, 1018.4, 1018.9, 1019.3, 1019.5, 1019.7, 1019.8, 
    1019.9, 1020.2, 1020.4, 1020.5, 1020.5, 1020.4, 1020.3, 1020.4, 1020.3, 
    1020, 1019.8, 1019.4, 1019.5, 1019.3, 1019.2, 1019.3, 1019.4, 1019.7, 
    1020.1, 1020.7, 1021, 1022, 1022.9, 1023.6, 1024.1, 1024.4, 1024.6, 
    1024.7, 1024.5, 1024.4, 1024.6, 1025, 1025.4, 1025.5, 1025.7, 1025.7, 
    1025.6, 1025.5, 1025.7, 1025.7, 1025.6, 1025, 1024.6, 1024.5, 1024.1, 
    1023.8, 1023.5, 1023.1, 1022.8, 1022.3, 1021.9, 1021.3, 1020.9, 1020.6, 
    1020.5, 1020.3, 1020.3, 1020.5, 1020.3, 1019.8, 1019.6, 1019.5, 1019.2, 
    1019.2, 1019.1, 1018.7, 1018.5, 1018.5, 1018.7, 1018.5, 1018.4, 1018, 
    1017.7, 1017.5, 1017.4, 1017.3, 1017, 1016.6, 1016.5, 1016.4, 1016.7, 
    1016.7, 1016.4, 1015.8, 1015.2, 1014.5, 1014.2, 1013.9, 1013.8, 1013.4, 
    1013.2, 1012.8, 1012.8, 1012.9, 1012.5, 1012.2, 1012.2, 1012.1, 1012, 
    1012.1, 1012.5, 1012.9, 1012.8, 1012.8, 1013, 1013.1, 1012.9, 1012.7, 
    1012.6, 1012.4, 1012.3, 1012.4, 1012.3, 1012.3, 1012, 1011.6, 1011.6, 
    1011.4, 1011, 1010.8, 1010.8, 1010.3, 1010, 1010.2, 1009.7, 1009.6, 
    1009.4, 1009.3, 1009.1, 1009.4, 1010, 1010.8, 1011.7, 1012, 1012.9, 
    1014.1, 1015.2, 1015.7, 1016.6, 1017.4, 1018.1, 1018.6, 1019, 1019.3, 
    1019.9, 1020.3, 1020.5, 1020.8, 1021.3, 1021.4, 1021.8, 1022.2, 1022.6, 
    1023, 1023.3, 1023.5, 1023.6, 1023.4, 1023.4, 1023.4, 1023.2, 1022.8, 
    1023.2, 1023.5, 1023.5, 1022.8, 1022.4, 1022.3, 1021.9, 1021.7, 1021, 
    1020.6, 1020.2, 1019.9, 1019.6, 1019.1, 1018.8, 1018.5, 1018.1, 1017.2, 
    1016.3, 1015.8, 1015.1, 1014.5, 1014.2, 1014.1, 1014.4, 1015, 1015.4, 
    1015.4, 1015.4, 1015.4, 1015.2, 1014.8, 1014.8, 1015.2, 1015.4, 1015.5, 
    1015.5, 1016, 1016.4, 1017, 1017.2, 1017.4, 1017.7, 1017.7, 1017.8, 
    1018.2, 1018.3, 1018.4, 1018.4, 1018.3, 1018.5, 1018.3, 1018, 1017.7, 
    1017.4, 1016.6, 1016, 1015.5, 1015.1, 1014.5, 1013.9, 1013.3, 1012.8, 
    1012, 1011.5, 1010.8, 1010.3, 1009.8, 1009.3, 1009.1, 1008.8, 1008.4, 
    1008, 1007.9, 1007.7, 1007.5, 1007.3, 1007.3, 1007.6, 1007.9, 1008.1, 
    1008, 1008.2, 1008.3, 1008.6, 1008.8, 1009.3, 1010, 1010.4, 1010.6, 1011, 
    1011.5, 1011.8, 1012.2, 1012.5, 1013, 1013.6, 1014, 1014.3, 1014.5, 
    1014.8, 1015.2, 1015.4, 1015.6, 1016, 1016.1, 1016.2, 1016.3, 1016.7, 
    1016.8, 1017, 1017.1, 1017.1, 1016.9, 1016.9, 1017.1, 1017, 1017, 1017, 
    1016.6, 1016.6, 1016.9, 1016.6, 1016.7, 1016.7, 1016.3, 1016.4, 1016.3, 
    1016.2, 1016.2, 1016.1, 1016.2, 1016.5, 1016.7, 1017.2, 1017.7, 1017.9, 
    1018.2, 1018.4, 1018.6, 1018.9, 1019.4, 1019.9, 1020.2, 1020.7, 1021.7, 
    1021.9, 1022.3, 1022.8, 1023.6, 1023.9, 1023.9, 1024.5, 1024.8, 1025.6, 
    1025.5, 1026.5, 1027.4, 1028, 1028.2, 1029, 1029.6, 1029.7, 1030, 1030.4, 
    1031, 1031.5, 1032, 1032.2, 1032.7, 1033.3, 1033.7, 1034, 1034.1, 1034.2, 
    1034.5, 1034.6, 1034.6, 1034.7, 1034.7, 1034.8, 1034.9, 1034.8, 1034.5, 
    1034.5, 1034, 1033.7, 1033.5, 1033.2, 1032.9, 1032.6, 1032.2, 1031.8, 
    1031.7, 1031.4, 1030.9, 1030.4, 1030, 1029.4, 1028.7, 1028.3, 1027.9, 
    1027.3, 1027, 1026.6, 1026.3, 1026.1, 1025.9, 1025.4, 1025, 1024.5, 1024, 
    1023.3, 1022.8, 1022.2, 1021.7, 1021.1, 1020.6, 1020.1, 1019.7, 1019.1, 
    1018.4, 1018.1, 1017.5, 1017.1, 1016.5, 1015.8, 1015.3, 1015, 1014.6, 
    1014.4, 1014.3, 1013.8, 1013.5, 1013.2, 1012.8, 1012.5, 1012.2, 1012.1, 
    1012, 1012, 1011.9, 1012.2, 1012.1, 1012.3, 1012.4, 1012.1, 1011.8, 
    1011.9, 1011.9, 1011.8, 1012, 1012.2, 1012.8, 1013.3, 1013.9, 1014.1, 
    1014.2, 1014.9, 1015.4, 1015.9, 1016.3, 1016.4, 1016.7, 1017.4, 1017.5, 
    1017.8, 1018.3, 1018.6, 1018.5, 1018.4, 1018.7, 1018.9, 1018.9, 1018.8, 
    1019.1, 1019.2, 1019.2, 1019.5, 1019.8, 1019.8, 1019.8, 1020.2, 1020.5, 
    1020.8, 1020.8, 1021, 1021.4, 1021.2, 1021.4, 1021.5, 1021.8, 1021.7, 
    1021.7, 1021.4, 1021.4, 1021.1, 1021, 1021.1, 1020.7, 1020.7, 1020.7, 
    1021.1, 1021.4, 1021.7, 1021.8, 1021.7, 1021.5, 1021.2, 1021, 1020.8, 
    1020.6, 1020.5, 1020.3, 1020.2, 1020.1, 1020.1, 1019.6, 1019.3, 1019.1, 
    1018.7, 1018.3, 1017.8, 1017.5, 1017.3, 1017.2, 1017.2, 1016.8, 1016.2, 
    1015.8, 1015.5, 1015.1, 1014.3, 1013.6, 1013.2, 1012.7, 1012.4, 1012, 
    1011.5, 1010.7, 1009.9, 1008.6, 1007.4, 1006.2, 1005.3, 1004.2, 1003.4, 
    1002.7, 1002.2, 1001.8, 1001.8, 1001.6, 1001.5, 1001.5, 1001.3, 1001.2, 
    1001.1, 1000.9, 1000.7, 1000.6, 1000.9, 1001.1, 1001.3, 1001.4, 1001.5, 
    1001.3, 1001.4, 1001.5, 1001.6, 1001.5, 1001.5, 1001.8, 1002, 1002.4, 
    1002.9, 1003.3, 1003.6, 1003.6, 1003.6, 1003.7, 1003.7, 1003.6, 1003.7, 
    1003.9, 1004.1, 1004.2, 1004, 1004, 1004, 1004, 1004, 1004.2, 1004.5, 
    1004.6, 1005, 1004.9, 1005.3, 1005.8, 1006, 1006.3, 1006.5, 1006.7, 1007, 
    1007.1, 1007.1, 1007.4, 1007.8, 1008, 1008.1, 1008.5, 1008.8, 1008.9, 
    1009.1, 1009.2, 1009.2, 1009.3, 1009.5, 1009.3, 1009.3, 1009.3, 1009.3, 
    1009.3, 1009.2, 1009.4, 1009.1, 1008.8, 1008.5, 1008.4, 1008.1, 1007.8, 
    1007.4, 1007.6, 1007.3, 1007.1, 1007.2, 1007, 1006.9, 1006.6, 1006.6, 
    1006.6, 1006.3, 1006.2, 1006, 1005.8, 1005.8, 1005.7, 1005.7, 1005.7, 
    1005.6, 1005.4, 1005.4, 1005.6, 1005.8, 1005.4, 1005.2, 1004.6, 1004.2, 
    1004, 1003.6, 1003.5, 1003.1, 1002.9, 1002.7, 1002.5, 1002.2, 1001.9, 
    1001.6, 1001.3, 1001.2, 1001, 1000.9, 1000.9, 1000.6, 1000.5, 1000.4, 
    1000.1, 999.8, 999.4, 999.2, 998.9, 998.9, 999.1, 999.3, 999, 998.7, 
    998.4, 998.1, 998.1, 997.9, 997.6, 997.3, 997, 996.8, 996.7, 996.6, 
    996.6, 996.5, 996.4, 996.1, 996, 995.8, 995.1, 994.7, 994.4, 994.1, 
    993.5, 993.1, 992.8, 992, 991.4, 991.2, 990.9, 990.7, 990.2, 989.9, 990, 
    989.5, 989.4, 989, 988.8, 988.4, 987.6, 987.3, 986.5, 985.9, 985.7, 
    985.5, 984.7, 984.3, 984.1, 983.8, 983.5, 983.5, 983.6, 984, 984.6, 
    985.3, 986.1, 987.2, 988, 988.9, 989.6, 990, 990.5, 990.6, 990.7, 991.1, 
    991.5, 992.2, 992.5, 993.1, 993.9, 994.7, 995.3, 995.8, 996.1, 996.5, 
    996.8, 996.7, 997.2, 997.6, 998, 998.3, 999.1, 999.8, 1000.3, 1001.3, 
    1002.1, 1002.8, 1003.6, 1004.2, 1004.2, 1004.4, 1004.7, 1005.7, 1005.8, 
    1006, 1006.4, 1006.5, 1006.8, 1007.3, 1007.6, 1007.7, 1007.7, 1007.7, 
    1007.6, 1007.8, 1007.8, 1007.6, 1007.4, 1007.4, 1007.7, 1007.4, 1006.9, 
    1006.8, 1006.6, 1005.9, 1005, 1004.7, 1004.2, 1003.4, 1003.3, 1002.7, 
    1002.6, 1003.3, 1003.3, 1002.7, 1002.8, 1003, 1003.7, 1004.3, 1004.7, 
    1004.8, 1005.7, 1006.1, 1006.3, 1006.4, 1006.3, 1006.1, 1005.9, 1005.7, 
    1005.4, 1005, 1004.8, 1004.4, 1004.3, 1004.2, 1004.1, 1003.8, 1003.5, 
    1003.3, 1003.2, 1003, 1002.7, 1002.6, 1002.4, 1002.6, 1002.6, 1002.7, 
    1002.7, 1002.6, 1002.5, 1002.3, 1002.2, 1002, 1002, 1001.9, 1001.7, 
    1001.7, 1001.7, 1001.7, 1001.6, 1001.4, 1001.1, 1000.8, 1000.5, 1000.3, 
    1000.1, 1000, 999.7, 999.5, 999.4, 999.3, 999.6, 999.6, 999.6, 999.7, 
    999.5, 999.5, 999.3, 999.5, 999.5, 999.4, 999.6, 1000, 999.9, 1000, 
    1000.1, 1000.3, 1000.4, 1000.7, 1000.9, 1001.3, 1001.7, 1002.2, 1002.7, 
    1003.4, 1004, 1004.6, 1005.3, 1005.8, 1006.4, 1007, 1007.3, 1007.7, 
    1008.3, 1009.1, 1009.5, 1010, 1010.6, 1011.2, 1011.7, 1012.2, 1012.6, 
    1013.1, 1013.2, 1013.3, 1013.3, 1013.8, 1014, 1014.4, 1015.2, 1015.8, 
    1016.3, 1017.1, 1017.2, 1017.5, 1017.7, 1018, 1018.4, 1018.7, 1018.8, 
    1019, 1019.3, 1019.2, 1019.4, 1019.3, 1019.2, 1019.4, 1019.2, 1018.9, 
    1019, 1019.2, 1019.1, 1019.3, 1019.4, 1019.5, 1019.4, 1019.2, 1019.3, 
    1019.1, 1018.8, 1018.5, 1018.2, 1018.1, 1017.9, 1017.7, 1017.5, 1017.2, 
    1017.1, 1016.7, 1016.3, 1016, 1015.4, 1014.9, 1014.6, 1014.4, 1013.9, 
    1013.8, 1013.4, 1013.2, 1012.9, 1012.3, 1011.6, 1011.4, 1010.9, 1010.8, 
    1010.6, 1010.4, 1010.3, 1010.1, 1010.1, 1009.9, 1009.5, 1009.2, 1008.8, 
    1008.4, 1007.8, 1007.3, 1007.1, 1006.8, 1007.1, 1006.8, 1006.3, 1006.6, 
    1006.2, 1006, 1005.8, 1005.7, 1005.6, 1005.1, 1004.8, 1004.8, 1004.6, 
    1004.6, 1004.6, 1004.4, 1004.3, 1004.1, 1003.7, 1003.4, 1003, 1002.7, 
    1002.6, 1002.3, 1002.2, 1002.1, 1001.9, 1001.6, 1001.3, 1001, 1000.7, 
    1000.3, 1000.1, 999.8, 999.3, 998.8, 998.6, 998.3, 998, 997.4, 997.1, 
    996.6, 996.3, 995.8, 995.5, 995.2, 994.7, 994.5, 994.4, 994.2, 994.2, 
    994, 994.1, 994.1, 994, 993.6, 993.3, 993.1, 993.1, 992.9, 992.9, 992.7, 
    992.8, 992.8, 992.6, 992.6, 992.3, 991.9, 991.6, 991.5, 991.2, 990.6, 
    991.1, 990.9, 990.9, 990.9, 990.8, 990.7, 990.3, 990.7, 991.1, 991.3, 
    991.4, 991.7, 991.8, 991.9, 992.6, 993.2, 993.2, 993, 992.8, 992.5, 
    992.6, 992.7, 993, 993.4, 994.1, 994.8, 995.5, 996.3, 997.1, 997.8, 
    998.4, 999.2, 1000, 1000.7, 1001.5, 1002.4, 1003.3, 1004.4, 1005.5, 
    1006.4, 1007.4, 1008.3, 1009.1, 1009.9, 1010.6, 1011, 1011.7, 1012.1, 
    1012.8, 1013.7, 1014.3, 1015.2, 1015.8, 1016.5, 1016.9, 1017.2, 1017.5, 
    1017.7, 1018, 1017.9, 1017.4, 1017.2, 1016.9, 1016.3, 1015.9, 1015.6, 
    1015.1, 1014.5, 1014.1, 1013.8, 1013.5, 1013.6, 1013.6, 1013.6, 1013.5, 
    1013.6, 1013.5, 1013.6, 1013.3, 1013.2, 1013.2, 1013, 1013, 1013, 1012.9, 
    1012.8, 1012.6, 1012.4, 1012.2, 1012.4, 1012.5, 1012.6, 1013.2, 1013.4, 
    1013.5, 1013.9, 1014.3, 1014.6, 1014.6, 1015.1, 1015.6, 1015.7, 1015.9, 
    1016.4, 1016.8, 1017.4, 1017.8, 1018.2, 1018.7, 1019, 1019.3, 1019.8, 
    1019.9, 1020, 1020.3, 1020.3, 1020.4, 1020.7, 1020.7, 1020.9, 1021.3, 
    1021.7, 1022.1, 1022.3, 1022.3, 1022.2, 1022.2, 1022.2, 1022.1, 1021.9, 
    1021.8, 1021, 1020.3, 1020, 1019.8, 1019.5, 1018.9, 1018.2, 1017.5, 
    1016.9, 1016.1, 1015.3, 1014.7, 1014.1, 1013.5, 1013.2, 1012.7, 1012.3, 
    1011.8, 1011.2, 1010.5, 1009.9, 1009.4, 1008.7, 1007.7, 1006.8, 1005.9, 
    1004.3, 1003.2, 1001.9, 1000.8, 999.7, 998.5, 997.1, 995.2, 993.8, 992.5, 
    992.1, 992.1, 993, 993.2, 993, 993, 992.9, 992.9, 994.2, 994.3, 994.7, 
    995.2, 993.6, 993.9, 994.4, 994.7, 995, 995.1, 995.5, 996, 996.4, 996.7, 
    997.4, 998.1, 998.9, 999.9, 1000.7, 1001.6, 1002.4, 1003.3, 1004.3, 
    1004.6, 1005.2, 1005.7, 1006.2, 1006.7, 1007.1, 1007.5, 1007.7, 1007.8, 
    1007.4, 1006.8, 1006.5, 1006.3, 1006.3, 1006.6, 1007, 1007.4, 1007.8, 
    1008.1, 1008.6, 1009.2, 1010.7, 1009.3, 1009.6, 1009.7, 1009.6, 1009.3, 
    1008.9, 1008.2, 1007.7, 1007.4, 1006.9, 1006.6, 1006.1, 1005.5, 1004.9, 
    1004.3, 1003.4, 1002.1, 1000.9, 999.7, 998.7, 997.6, 996.6, 995.3, 994.2, 
    992.6, 990.9, 989.8, 988.9, 987.7, 986.4, 984.9, 983.4, 982.5, 981.6, 
    980.7, 980.3, 980.3, 980.1, 979.7, 979.3, 979.6, 979, 978.5, 978.3, 
    978.1, 978.1, 977.6, 978.2, 978.1, 977.6, 977.2, 976.9, 977.2, 977.2, 
    977.1, 977.1, 977.5, 977.8, 977.9, 977.8, 977.7, 978.3, 977.8, 978, 
    977.9, 978.2, 978.7, 979.3, 979.7, 980.4, 981.1, 981.6, 981.9, 982.5, 
    982.6, 983.5, 983.6, 983.8, 983.9, 984.4, 984.8, 985.1, 985.5, 985.7, 
    986.1, 986.1, 986.2, 986.2, 986.1, 985.9, 985.8, 985.8, 985.9, 986.2, 
    986.2, 986, 986.1, 986, 986.1, 986.2, 986.3, 986.2, 986.1, 986.1, 986.2, 
    986.4, 986.4, 986.6, 986.8, 986.8, 987.1, 987.2, 987.3, 987.4, 987.9, 
    988.5, 989, 989.8, 990.1, 990.7, 991.1, 991.8, 992.4, 992.9, 993.8, 
    994.3, 994.7, 995.3, 995.8, 996.2, 996.8, 997.1, 997.4, 997.7, 998.1, 
    998.3, 998.5, 998.6, 998.4, 998.3, 998.1, 998.1, 998.3, 998.2, 998, 
    997.9, 997.8, 997.5, 997, 996.4, 996, 995.9, 995.9, 995.9, 996.2, 996.3, 
    996.6, 996.9, 997.1, 997.7, 998.4, 999, 999.7, 1000.4, 1001.3, 1002.4, 
    1003, 1003.8, 1004.5, 1005.1, 1005.8, 1006.3, 1006.7, 1006.9, 1007.1, 
    1007.4, 1007.6, 1007.9, 1008.3, 1009, 1009.1, 1009.1, 1009.3, 1009.3, 
    1009, 1008.3, 1008, 1007.8, 1007.8, 1007.7, 1007.1, 1006.8, 1006.2, 
    1005.7, 1005, 1004.4, 1004, 1004, 1003.9, 1003.7, 1003.7, 1003.7, 1003.7, 
    1003.6, 1003.7, 1003.7, 1003.9, 1003.8, 1003.9, 1004, 1004, 1004.1, 
    1004.4, 1004.8, 1005.3, 1005.8, 1005.9, 1005.6, 1005.5, 1005.7, 1005.9, 
    1005.8, 1005.6, 1005.5, 1005.6, 1005.7, 1005.7, 1005.9, 1006, 1006, 
    1006.1, 1006.1, 1006.2, 1006.1, 1006.1, 1006.1, 1006.6, 1006.7, 1006.9, 
    1006.9, 1006.9, 1007.2, 1007.1, 1007.2, 1007.2, 1007.1, 1007.1, 1007.2, 
    1007.2, 1007.4, 1007.6, 1007.7, 1007.7, 1007.6, 1007.6, 1007.5, 1007.6, 
    1007.5, 1007.8, 1007.9, 1008.1, 1008.2, 1008.4, 1008.3, 1008.5, 1008.6, 
    1008.8, 1008.8, 1008.9, 1008.7, 1008.6, 1008.5, 1008.6, 1008.6, 1008.9, 
    1009, 1008.5, 1008.1, 1008.1, 1007.6, 1007.4, 1007, 1006.5, 1006.4, 
    1005.9, 1005.5, 1005.3, 1005.1, 1005.2, 1004.9, 1005, 1004.4, 1004.6, 
    1004.4, 1004.3, 1004, 1004, 1003.8, 1003.6, 1003.7, 1003.5, 1003.1, 
    1002.6, 1002.5, 1002.2, 1001.9, 1001.4, 1001.5, 1001.7, 1001.8, 1002.3, 
    1002.8, 1003.2, 1003.5, 1003.4, 1003.4, 1003.1, 1003.1, 1003, 1003, 
    1002.9, 1003.1, 1003.3, 1003.2, 1003.1, 1002.9, 1002.8, 1003, 1002.9, 
    1003, 1003.2, 1003.3, 1003.3, 1003.5, 1003.8, 1004, 1004.2, 1004.3, 
    1004.4, 1004.6, 1005, 1004.9, 1005, 1005.3, 1005.4, 1005.7, 1005.9, 
    1005.8, 1005.8, 1005.7, 1005.6, 1005.7, 1005.5, 1005.2, 1005, 1004.7, 
    1004.6, 1004.4, 1004, 1003.4, 1002.9, 1002.5, 1001.9, 1001.3, 1000.8, 
    1000, 999.4, 998.5, 997.8, 997, 996.4, 995.8, 995.1, 994.3, 993.4, 992.4, 
    991.6, 990.6, 990, 989.4, 989, 988.8, 988.6, 988.5, 988.4, 988.2, 987.9, 
    988, 988.1, 988.1, 988.2, 988.4, 988.6, 988.8, 989, 989, 989.2, 989.2, 
    989.2, 989.3, 989.3, 989.5, 989.6, 990.1, 990.3, 990.7, 991.1, 991.2, 
    991.6, 992, 992.3, 992.6, 992.9, 993.3, 993.6, 994.1, 994.4, 994.7, 
    995.2, 995.3, 995.7, 995.9, 996.3, 996.7, 997, 997.4, 997.6, 997.9, 
    998.3, 998.6, 998.8, 998.8, 998.7, 998.7, 998.4, 998, 997.8, 997.6, 
    997.7, 997.6, 997.5, 997.6, 997.7, 997.5, 997.6, 997.5, 997.5, 997.7, 
    997.9, 998, 998.1, 998.3, 998.5, 998.7, 999, 999.1, 999.4, 999.5, 999.8, 
    1000.1, 1000.6, 1001.1, 1001.8, 1002.7, 1003.6, 1004.4, 1005.1, 1005.9, 
    1006.7, 1007.3, 1008.1, 1008.7, 1009.3, 1009.8, 1010.2, 1010.4, 1010.3, 
    1010.1, 1009.7, 1009.9, 1009.5, 1009.7, 1010.2, 1011.1, 1012.1, 1013.3, 
    1014.2, 1015.2, 1016.6, 1017.4, 1017.8, 1018.2, 1018.5, 1018.7, 1018.8, 
    1018.2, 1018.1, 1016.9, 1016.4, 1016, 1015.2, 1014.7, 1014, 1013.6, 
    1013.4, 1013.4, 1013.5, 1013.8, 1014.2, 1014.8, 1015.7, 1016.5, 1017.4, 
    1018.4, 1019.5, 1020, 1020.2, 1021.5, 1022, 1022.2, 1022.4, 1022.3, 
    1022.3, 1022.4, 1022.3, 1022.3, 1021.4, 1020.8, 1020.2, 1019.1, 1018.6, 
    1017.2, 1015.9, 1014.7, 1013.4, 1011.9, 1009.8, 1008.4, 1007.9, 1007.5, 
    1007.6, 1007.9, 1007.8, 1007.5, 1007.3, 1007.3, 1007.3, 1006.9, 1006.6, 
    1006.4, 1006.7, 1006.6, 1006.6, 1006.7, 1005.9, 1005.3, 1004.9, 1004.4, 
    1004.5, 1004.8, 1005.4, 1005.8, 1006.5, 1006.9, 1007.3, 1007.9, 1008.2, 
    1008.8, 1009.4, 1009.9, 1010.7, 1011.1, 1012.1, 1012.5, 1013.3, 1013.5, 
    1013.7, 1014.1, 1014.5, 1014.5, 1015, 1014.7, 1014.8, 1015.4, 1015.5, 
    1016, 1016, 1015.8, 1016.2, 1016.1, 1016.4, 1016.5, 1016.7, 1016.5, 
    1016.4, 1016.7, 1016.9, 1017.1, 1017.1, 1017.1, 1017.2, 1016.9, 1016.8, 
    1016.6, 1016.6, 1016.5, 1016.4, 1016.6, 1016.9, 1016.9, 1017, 1016.6, 
    1016.4, 1016.6, 1016.7, 1016.6, 1016.4, 1016.1, 1015.9, 1015.7, 1015.7, 
    1015.8, 1015.9, 1015.6, 1015.4, 1015.3, 1015.1, 1014.9, 1015, 1015, 
    1014.5, 1014.6, 1014.8, 1015.3, 1015.2, 1014.9, 1014.3, 1014.1, 1014, 
    1013.7, 1013.3, 1012.6, 1011.7, 1010.9, 1010.3, 1009.7, 1009.2, 1008.7, 
    1007.8, 1007.4, 1006.9, 1006.3, 1005.8, 1005.2, 1004.8, 1004.7, 1004.6, 
    1004.2, 1003.8, 1004, 1004, 1004.1, 1004.1, 1004.4, 1004.7, 1004.6, 
    1004.3, 1004.2, 1004.7, 1004.9, 1005.3, 1005.4, 1005.4, 1005.6, 1005.8, 
    1006, 1006.1, 1006.3, 1006.3, 1006.3, 1006.4, 1006.7, 1007.1, 1007.3, 
    1007.3, 1007, 1007, 1007.1, 1007.2, 1007.1, 1007.1, 1007, 1007.1, 1007.3, 
    1007.3, 1007.1, 1007.1, 1007, 1006.9, 1006.9, 1006.7, 1006.4, 1005.8, 
    1005.6, 1005.3, 1005, 1004.8, 1004.5, 1004.2, 1003.6, 1003.3, 1002.8, 
    1002, 1001.5, 1000.8, 1000.1, 999.4, 998.8, 998, 997.1, 996.4, 995.7, 
    995.3, 995.2, 995, 994.9, 995, 995.3, 995.4, 995.7, 996.3, 996.5, 996.7, 
    997.2, 997.7, 998, 998.3, 998.3, 998.5, 998.7, 999.3, 999.6, 1000, 
    1000.4, 1000.8, 1001.2, 1001.5, 1001.9, 1002.3, 1002.5, 1002.9, 1003.3, 
    1003.7, 1004, 1004.5, 1004.9, 1005.5, 1005.8, 1006.1, 1006.5, 1007.1, 
    1007.4, 1007.8, 1008, 1008.7, 1009.1, 1009.9, 1010.6, 1011.2, 1011.6, 
    1012.1, 1012.4, 1012.8, 1013.1, 1013.5, 1013.8, 1014.2, 1014.8, 1015.2, 
    1016, 1016.4, 1017, 1017.4, 1017.7, 1017.8, 1018.1, 1018.4, 1018.8, 
    1019.3, 1019.8, 1020.1, 1020.2, 1020.5, 1020.9, 1021.1, 1021.2, 1021.2, 
    1021.4, 1021.3, 1021.4, 1021.4, 1021.7, 1021.9, 1022, 1022.2, 1021.7, 
    1021.3, 1021.2, 1021.2, 1020.9, 1020.7, 1020.6, 1020.8, 1020.8, 1020.6, 
    1020.7, 1020.7, 1020.5, 1020.4, 1020.1, 1019.6, 1019, 1018.7, 1017.9, 
    1017.5, 1017.1, 1016.6, 1016, 1015.8, 1015.6, 1015.3, 1014.9, 1014.4, 
    1014, 1013.7, 1013.2, 1012.7, 1012.5, 1012.1, 1011.7, 1011, 1010.3, 
    1009.6, 1008.7, 1008, 1007.1, 1006.3, 1005.6, 1005.1, 1004.4, 1003.6, 
    1002.5, 1001.5, 1000.7, 999.7, 999, 998.1, 997.3, 996.5, 995.8, 995.2, 
    994.6, 994.2, 993.8, 993, 992.8, 992.6, 992.5, 992.6, 992.5, 992.6, 993, 
    993.3, 993.5, 993.8, 993.8, 994.1, 994.1, 994, 993.6, 993.1, 992.6, 
    992.3, 992.3, 992.4, 992.2, 992.3, 992.3, 992.5, 992.8, 993.1, 993.5, 
    994.1, 994.4, 994.9, 995.2, 995.6, 996, 996.1, 996.4, 996.5, 996.5, 
    996.7, 996.9, 997, 997.2, 997.3, 997.6, 997.7, 998.2, 998.6, 999, 999.4, 
    999.6, 1000, 999.9, 1000.2, 1000.8, 1001, 1001.3, 1001.6, 1002, 1002.4, 
    1002.6, 1002.4, 1002.1, 1002, 1002.3, 1002.2, 1002.3, 1002.1, 1002, 1002, 
    1002, 1002, 1001.9, 1002, 1002, 1001.8, 1001.8, 1001.7, 1001.7, 1001.6, 
    1001.7, 1001.9, 1002.2, 1002.2, 1002.2, 1002.1, 1002.5, 1002.6, 1002.8, 
    1003.1, 1003.5, 1003.7, 1003.7, 1004, 1004.3, 1004.4, 1004.3, 1004.7, 
    1004.8, 1004.9, 1004.9, 1005.1, 1005.2, 1005.4, 1005.7, 1006, 1006.2, 
    1006.1, 1006.3, 1006.7, 1007, 1007.3, 1007.6, 1007.8, 1008.1, 1008.3, 
    1008.2, 1008.1, 1008.2, 1008.5, 1008.8, 1008.6, 1008, 1008.1, 1007.9, 
    1008, 1007.9, 1007.9, 1007.8, 1007.6, 1007.3, 1007.1, 1006.8, 1006.2, 
    1005.7, 1004.9, 1004.1, 1003.2, 1002.1, 1000.9, 999.6, 998.5, 997.3, 
    995.9, 994.2, 992.9, 991, 989.5, 987.9, 987, 985.8, 984.6, 983.3, 982.1, 
    981.2, 979.9, 978.7, 977.8, 976.6, 975, 974.4, 973.9, 974.1, 974.3, 
    974.8, 975.2, 975.7, 976.3, 976.7, 977.3, 977.3, 978.9, 979.6, 980.2, 
    981.1, 981.9, 983, 983.9, 984.9, 985.6, 986.3, 987.4, 988.3, 989, 989.7, 
    990.3, 991, 991.4, 992, 992.5, 993.1, 993.6, 993.9, 994, 994.2, 994.3, 
    994.3, 994.3, 994, 993.5, 993, 992.6, 992.2, 992.1, 991.8, 991.4, 991, 
    990.7, 990.4, 989.9, 989.8, 990, 990.2, 990.3, 990.5, 991, 991.5, 992.2, 
    993, 994, 994.9, 995.7, 996.6, 997.7, 998.9, 999.9, 1001, 1001.9, 1003.2, 
    1004.3, 1005.3, 1006.2, 1007.3, 1008, 1008.3, 1008.3, 1008.5, 1008.6, 
    1008.6, 1008.6, 1008.3, 1007.9, 1007.7, 1007.5, 1006.8, 1006, 1005.5, 
    1005, 1004.7, 1004.7, 1004.8, 1004.6, 1004.9, 1005.1, 1005.4, 1005.4, 
    1004.9, 1004.8, 1004.5, 1004.2, 1003.7, 1003.3, 1002.9, 1002.4, 1001.9, 
    1001.3, 1000.7, 1000.1, 999.6, 999, 998.9, 999.1, 999.3, 1000, 1000.7, 
    1001.8, 1002.8, 1003.9, 1004.4, 1005.6, 1006.6, 1007.6, 1009, 1010.2, 
    1011, 1012.4, 1013.4, 1014.4, 1015.3, 1016.2, 1016.9, 1017.6, 1018.1, 
    1018.3, 1018.7, 1018.8, 1019, 1019.4, 1019.6, 1019.6, 1019.7, 1019.7, 
    1019.7, 1019.8, 1019.7, 1019.8, 1019.6, 1019.2, 1019.2, 1019.2, 1019.1, 
    1018.8, 1018.3, 1018.2, 1017.8, 1017.7, 1017.2, 1016.4, 1016.5, 1016.5, 
    1016.5, 1016.7, 1016.9, 1017, 1017.3, 1017.6, 1018.1, 1018.3, 1018.7, 
    1019.4, 1019.9, 1020.4, 1020.8, 1021.7, 1022.2, 1022.5, 1023, 1023.7, 
    1024.2, 1024.6, 1024.8, 1024.9, 1025.2, 1025.3, 1025.4, 1025.7, 1026, 
    1026, 1025.9, 1025.8, 1025.7, 1025.5, 1025.2, 1025, 1024.6, 1024.6, 
    1024.5, 1024.2, 1024, 1024, 1023.9, 1023.7, 1023.4, 1023.2, 1023, 1022.9, 
    1022.6, 1022.5, 1022.6, 1022.8, 1022.9, 1022.9, 1022.9, 1023, 1023, 1023, 
    1022.9, 1022.9, 1022.9, 1022.9, 1023, 1023, 1022.9, 1022.7, 1022.7, 
    1022.5, 1022.6, 1022.4, 1021.5, 1021.1, 1021.5, 1021.3, 1021.2, 1021, 
    1020.8, 1020.5, 1020.1, 1019.7, 1019.3, 1018.9, 1018.6, 1018.2, 1017.4, 
    1017.3, 1017, 1016.7, 1016.5, 1016.5, 1016.3, 1016.4, 1016.5, 1016.3, 
    1016.2, 1016.2, 1016.2, 1016.4, 1016.6, 1016.9, 1017.4, 1017.9, 1018.2, 
    1018.7, 1018.9, 1019.1, 1019.3, 1019.7, 1019.9, 1020.4, 1021, 1021.5, 
    1021.9, 1022.5, 1022.7, 1023.2, 1023.9, 1024.2, 1024.5, 1024.6, 1024.7, 
    1024.9, 1025.2, 1025.4, 1025.3, 1025.4, 1025.4, 1025.3, 1025, 1024.7, 
    1024.2, 1023.6, 1023.2, 1022.5, 1022, 1021.7, 1021.3, 1021.2, 1021.3, 
    1021.4, 1021.3, 1021.1, 1021.3, 1021.2, 1021, 1021, 1021, 1021.3, 1021.5, 
    1021.2, 1020.9, 1020.7, 1020.7, 1020.5, 1020.4, 1020.2, 1020.1, 1020.1, 
    1020.1, 1020.2, 1020.1, 1020.1, 1019.9, 1020, 1019.9, 1019.7, 1019.6, 
    1019.4, 1019.2, 1019, 1018.9, 1018.8, 1018.7, 1018.8, 1018.3, 1018.2, 
    1018.2, 1018, 1017.8, 1018, 1018, 1018, 1018.2, 1018.1, 1018.3, 1018.2, 
    1018.5, 1018.4, 1018.4, 1018.6, 1018.8, 1019.2, 1019.3, 1019.4, 1019.6, 
    1020.1, 1020.3, 1020.6, 1020.8, 1021, 1021.3, 1021.5, 1021.9, 1022.2, 
    1022.4, 1022.7, 1022.8, 1023.2, 1023.6, 1023.6, 1024, 1024.2, 1024.4, 
    1024.6, 1024.6, 1024.8, 1024.9, 1025, 1025.1, 1025.2, 1025.3, 1025.4, 
    1025.6, 1025.6, 1025.5, 1025.4, 1025.5, 1025.2, 1025.2, 1025, 1024.9, 
    1025, 1025, 1024.9, 1024.7, 1024.5, 1024.3, 1024.3, 1024, 1023.7, 1023.7, 
    1023.5, 1023.4, 1023.3, 1023.2, 1023, 1022.9, 1022.7, 1022.6, 1022.5, 
    1022.2, 1022.1, 1022, 1022.1, 1022.1, 1022, 1022, 1022.1, 1022.3, 1022.3, 
    1022.4, 1022.5, 1022.6, 1022.7, 1022.7, 1022.9, 1022.8, 1022.8, 1023.1, 
    1023.3, 1023.3, 1023.3, 1023.1, 1023, 1023.2, 1023.1, 1023, 1023.2, 
    1023.2, 1023.2, 1023.4, 1023.3, 1023.4, 1023.4, 1023.4, 1023.4, 1023.7, 
    1023.8, 1023.7, 1023.6, 1023.6, 1023.6, 1023.6, 1023.8, 1024.1, 1024.3, 
    1024.8, 1024.9, 1025.1, 1025.4, 1025.7, 1025.9, 1026.1, 1026.3, 1026.3, 
    1026.6, 1026.9, 1026.9, 1026.7, 1026.5, 1026.6, 1026.8, 1027, 1027, 1027, 
    1027, 1026.8, 1026.7, 1026.2, 1025.9, 1025.6, 1025.5, 1025, 1024.5, 
    1024.2, 1023.8, 1023.4, 1023.1, 1022.8, 1022.5, 1022.2, 1021.7, 1021.2, 
    1020.8, 1020.3, 1019.9, 1019.4, 1018.8, 1018.2, 1017.5, 1016.7, 1016.2, 
    1015.4, 1014.6, 1014.2, 1013.7, 1013.4, 1013.1, 1012.8, 1012.9, 1013.6, 
    1013.8, 1014.2, 1014.5, 1014.7, 1014.8, 1014.8, 1014.6, 1014.3, 1014.3, 
    1014.1, 1013.8, 1013.5, 1013, 1012.6, 1012.1, 1011.8, 1011.2, 1010.8, 
    1010.2, 1009.6, 1009.1, 1008.9, 1008.7, 1008.6, 1008.4, 1008.2, 1008.1, 
    1008.1, 1008, 1007.8, 1007.6, 1007.4, 1007.3, 1007.2, 1007.3, 1007.3, 
    1007.5, 1007.4, 1007.6, 1007.5, 1007.6, 1007.6, 1007.6, 1007.5, 1007.3, 
    1007.4, 1007.4, 1007.6, 1007.8, 1007.7, 1007.5, 1007.4, 1007.3, 1006.9, 
    1007, 1007.1, 1007.1, 1007.1, 1007.2, 1007.4, 1007.3, 1007.4, 1007.3, 
    1007.4, 1007.4, 1007.5, 1007.3, 1007.2, 1006.9, 1006.9, 1006.9, 1007, 
    1007, 1006.9, 1006.6, 1006.7, 1006.6, 1006.6, 1006.6, 1006.4, 1006.3, 
    1006.2, 1006.3, 1006.4, 1006.7, 1006.7, 1006.9, 1006.9, 1007.1, 1007.1, 
    1007.1, 1007.1, 1007.2, 1007.2, 1007.2, 1007.5, 1007.7, 1007.9, 1008.2, 
    1008.5, 1008.6, 1008.9, 1008.9, 1009, 1009.2, 1009.2, 1009.4, 1009.6, 
    1009.9, 1010.1, 1010.2, 1010.2, 1010.3, 1010.2, 1010.2, 1010.1, 1009.8, 
    1009.9, 1009.9, 1009.9, 1009.9, 1010, 1010.2, 1010.3, 1010.3, 1010.4, 
    1010.3, 1010.4, 1010.5, 1010.7, 1011, 1011.2, 1011.4, 1011.7, 1011.8, 
    1011.9, 1012.1, 1012.1, 1012.3, 1012.5, 1012.4, 1012.6, 1012.7, 1012.9, 
    1013.2, 1013.5, 1013.7, 1014, 1014, 1014.1, 1014.2, 1014.3, 1014.3, 
    1014.5, 1014.6, 1014.7, 1014.9, 1014.9, 1015.1, 1015.2, 1015.1, 1015.1, 
    1014.9, 1014.8, 1014.9, 1014.7, 1014.6, 1014.6, 1014.6, 1014.4, 1014.3, 
    1014.2, 1014.4, 1014.3, 1014.1, 1013.5, 1013.2, 1012.6, 1012.3, 1011.6, 
    1011.2, 1010.8, 1010.2, 1009.6, 1009.6, 1009.3, 1009.2, 1009, 1008.6, 
    1008.3, 1008, 1007.7, 1007.2, 1006.8, 1006.3, 1005.8, 1005.2, 1004.4, 
    1003.4, 1002.3, 1001.2, 1000.1, 999.2, 998.2, 997.2, 996.4, 995.7, 995.3, 
    994.9, 994.7, 994.3, 994, 993.2, 993.9, 994.1, 995.2, 996.5, 997.1, 
    997.1, 997.4, 998.1, 998.2, 998, 998.4, 998.5, 998.9, 999, 999.2, 999.5, 
    1000, 1000.6, 1001, 1001.7, 1002.3, 1003, 1003.9, 1004.6, 1005.1, 1005.9, 
    1006.9, 1007.8, 1008.6, 1009.3, 1010, 1010.8, 1011.4, 1011.9, 1012.2, 
    1012.7, 1013.1, 1013.5, 1014.2, 1014.7, 1015.2, 1015.4, 1015.7, 1015.8, 
    1015.9, 1016, 1015.8, 1015.6, 1015.4, 1015.3, 1015.3, 1015, 1014.9, 
    1014.7, 1014.4, 1014.1, 1013.9, 1013.6, 1013.3, 1012.9, 1012.7, 1012.6, 
    1012.6, 1012.4, 1012.4, 1012.4, 1012.6, 1012.4, 1012.4, 1012.2, 1011.9, 
    1011.7, 1011.6, 1011.6, 1011.7, 1011.8, 1011.6, 1011.4, 1011.4, 1011.4, 
    1011.2, 1010.9, 1011.1, 1011.4, 1011.2, 1011, 1011.1, 1011.1, 1010.8, 
    1010.4, 1009.8, 1009.5, 1009.1, 1009.1, 1008.7, 1008.1, 1007.5, 1007.1, 
    1007.1, 1007, 1007, 1007.6, 1007.8, 1008.3, 1008.9, 1009.5, 1009.9, 
    1010.3, 1011, 1011.6, 1012.3, 1013, 1013.7, 1014.4, 1014.9, 1015.6, 
    1015.9, 1016.3, 1016.5, 1017, 1017.2, 1017.6, 1017.9, 1018.5, 1018.9, 
    1019.5, 1020, 1020.3, 1020.8, 1021, 1021.2, 1021.5, 1021.8, 1022.1, 
    1022.6, 1023, 1023.5, 1024, 1024.1, 1024.4, 1024.7, 1024.8, 1025.1, 
    1024.8, 1025.1, 1025.2, 1025.4, 1025.4, 1025.7, 1026.1, 1026.3, 1026.4, 
    1026.3, 1026.4, 1026.3, 1026.1, 1025.9, 1025.7, 1025.7, 1025.7, 1025.8, 
    1025.7, 1025.6, 1025.6, 1025.6, 1025.4, 1025.4, 1025.4, 1025.5, 1025.6, 
    1025.8, 1026, 1026.3, 1026.4, 1026.5, 1026.7, 1027, 1027.3, 1027.6, 
    1027.8, 1028, 1028.2, 1028.5, 1028.8, 1029.2, 1029.7, 1030.1, 1030.4, 
    1030.8, 1031.1, 1031.3, 1031.4, 1031.7, 1031.9, 1032.2, 1032.4, 1032.7, 
    1032.9, 1033.1, 1033.5, 1033.7, 1033.7, 1033.7, 1034, 1033.9, 1033.9, 
    1034, 1034.3, 1034.3, 1034.6, 1034.9, 1034.8, 1034.7, 1035, 1034.9, 
    1034.8, 1034.8, 1034.9, 1035, 1034.9, 1035, 1035.1, 1034.9, 1034.9, 
    1034.8, 1034.8, 1034.4, 1034, 1033.8, 1033.5, 1033.2, 1033, 1032.8, 
    1032.6, 1032.2, 1032, 1032, 1031.8, 1031.6, 1031.5, 1031.2, 1030.9, 
    1030.8, 1030.8, 1030.8, 1030.5, 1030.8, 1030.4, 1030.1, 1029.6, 1029, 
    1028.5, 1028, 1027.5, 1027, 1027.1, 1027.4, 1027.4, 1027.3, 1027.4, 
    1027.3, 1027.1, 1027.2, 1027, 1026.9, 1026.8, 1026.7, 1026.2, 1025.9, 
    1025.6, 1025.4, 1025.1, 1025, 1024.5, 1024, 1023.5, 1023.3, 1023.1, 
    1022.9, 1022.9, 1022.7, 1022.5, 1022.6, 1022.7, 1022.4, 1022.3, 1022.2, 
    1022.1, 1022.3, 1022.3, 1022.5, 1022.9, 1023.2, 1023.2, 1023.3, 1023.3, 
    1023.2, 1022.7, 1022.6, 1022.5, 1022.2, 1022, 1021.8, 1021.5, 1021.3, 
    1020.9, 1020.8, 1020.5, 1020.1, 1020, 1019.8, 1019.5, 1019.1, 1019.1, 
    1019, 1018.9, 1018.7, 1018.5, 1018.3, 1017.8, 1017.6, 1017.1, 1016.8, 
    1016.4, 1015.8, 1015.5, 1015.2, 1015.1, 1014.8, 1014.6, 1014.4, 1014.4, 
    1014.2, 1014, 1013.8, 1013.8, 1014, 1014.1, 1014, 1014.2, 1014.2, 1014.2, 
    1014.3, 1014.2, 1014.3, 1014.4, 1014.5, 1014.6, 1014.6, 1014.4, 1014.5, 
    1014.8, 1014.9, 1015, 1015.1, 1015.3, 1015.2, 1015.4, 1015.4, 1015.5, 
    1015.5, 1015.7, 1015.8, 1016.4, 1016.8, 1016.9, 1017.2, 1017.4, 1017.6, 
    1017.8, 1017.7, 1017.8, 1017.7, 1018, 1018.1, 1018.2, 1018.3, 1018.3, 
    1018.3, 1018.4, 1018.4, 1018.5, 1018.2, 1018.2, 1018, 1017.8, 1017.7, 
    1017.7, 1017.9, 1017.4, 1017.2, 1016.8, 1016.6, 1016.3, 1016, 1015.7, 
    1015.5, 1015.4, 1015.1, 1014.9, 1014.8, 1014.6, 1014.2, 1013.9, 1013.8, 
    1013.8, 1013.7, 1013.6, 1013.7, 1014.1, 1014.5, 1015.2, 1015.5, 1016, 
    1016.4, 1017, 1017.5, 1018, 1018.4, 1018.9, 1019.4, 1019.9, 1020.2, 
    1020.6, 1021.1, 1021.9, 1022.1, 1022.6, 1023, 1023.2, 1023.4, 1023.5, 
    1023.9, 1024.3, 1024.7, 1025, 1025.2, 1025.4, 1025.7, 1025.8, 1025.8, 
    1025.8, 1025.8, 1025.6, 1025.4, 1025.1, 1025, 1025, 1024.8, 1024.6, 
    1024.6, 1024.4, 1024.1, 1024, 1023.7, 1023.3, 1023.1, 1022.8, 1022.5, 
    1022.2, 1021.8, 1021.7, 1021.4, 1021.2, 1021, 1020.7, 1020.4, 1020.4, 
    1020.1, 1019.8, 1019.5, 1019.5, 1019.4, 1019.4, 1019.1, 1019.1, 1018.9, 
    1018.6, 1018.7, 1018.4, 1018.3, 1018.3, 1018.1, 1018.1, 1018.2, 1018, 
    1017.8, 1017.9, 1018.1, 1018.1, 1018, 1017.7, 1017.7, 1017.6, 1017.7, 
    1017.9, 1018.1, 1018.2, 1018.2, 1018.4, 1018.5, 1018.5, 1018.6, 1018.6, 
    1018.6, 1018.5, 1018.7, 1018.6, 1018.6, 1018.4, 1018.4, 1018.2, 1018, 
    1017.6, 1017.5, 1017.4, 1016.9, 1016.7, 1016.6, 1016.5, 1016.3, 1016, 
    1015.9, 1015.9, 1015.9, 1015.8, 1015.6, 1015.7, 1015.4, 1015.5, 1015.3, 
    1015.3, 1015.6, 1015.7, 1015.8, 1016, 1016.3, 1016.4, 1016.7, 1016.7, 
    1016.8, 1017.1, 1017.4, 1017.6, 1018.2, 1018.7, 1019, 1019.1, 1019.3, 
    1019.6, 1020, 1020.1, 1020.4, 1020.5, 1020.9, 1021.2, 1021.5, 1021.8, 
    1021.9, 1022, 1022.1, 1022.2, 1022.3, 1022.2, 1022.1, 1022, 1021.9, 
    1021.9, 1022.1, 1021.7, 1021.3, 1021, 1020.6, 1020.6, 1020.2, 1019.7, 
    1019.4, 1018.9, 1018.6, 1018.3, 1017.8, 1017.6, 1017.3, 1016.9, 1016.7, 
    1016.5, 1016.4, 1016, 1015.6, 1015.5, 1015.5, 1015.7, 1015.9, 1015.8, 
    1015.9, 1015.8, 1015.9, 1016, 1015.8, 1015.8, 1015.6, 1015.7, 1015.7, 
    1015.8, 1015.9, 1015.9, 1015.6, 1015.5, 1015.4, 1015.3, 1015.1, 1014.8, 
    1014.6, 1014.2, 1014.1, 1014.2, 1014, 1014, 1013.9, 1013.8, 1013.5, 
    1013.4, 1013.5, 1013.6, 1013.6, 1013.6, 1013.9, 1014.1, 1014.3, 1014.5, 
    1014.7, 1014.9, 1015, 1015.2, 1015.1, 1015.3, 1015.5, 1015.7, 1015.9, 
    1016.1, 1016.5, 1016.3, 1016.3, 1016.3, 1016.4, 1016.3, 1016.3, 1016.1, 
    1015.9, 1015.6, 1015.3, 1015, 1014.8, 1014.1, 1013.7, 1013.4, 1012.8, 
    1012.2, 1011.5, 1011.3, 1010.8, 1010.1, 1009.7, 1009.2, 1009, 1008.4, 
    1007.8, 1007.4, 1007.2, 1006.6, 1006.4, 1006.2, 1006.1, 1005.9, 1005.7, 
    1005.5, 1004.9, 1004.1, 1003.7, 1003.2, 1003.5, 1004.3, 1004.5, 1005, 
    1004.8, 1004.5, 1004.2, 1004.3, 1004.2, 1004.9, 1005.4, 1005.7, 1005.8, 
    1006.1, 1006.4, 1007.1, 1007.5, 1007.6, 1008.5, 1009.1, 1009.6, 1010.2, 
    1010.7, 1011.4, 1011.4, 1012.2, 1012.7, 1013.1, 1013.3, 1013.7, 1014.1, 
    1014.9, 1015, 1015.9, 1015.5, 1015.8, 1016, 1016.3, 1016.1, 1016, 1015.9, 
    1015.8, 1015.5, 1015.2, 1014.9, 1014.5, 1014.1, 1013.6, 1013.1, 1012.6, 
    1011.9, 1011.4, 1011, 1010.6, 1009.8, 1009.1, 1008.7, 1008.1, 1007.7, 
    1007.2, 1006.9, 1006.8, 1006.6, 1006.4, 1006.4, 1006.5, 1006.5, 1006.7, 
    1006.9, 1007.4, 1007.6, 1007.9, 1008.3, 1008.7, 1009.1, 1009.1, 1009.3, 
    1009.3, 1009.3, 1009.3, 1009.6, 1009.8, 1010, 1010.2, 1010.5, 1010.7, 
    1010.9, 1010.9, 1011.2, 1011.3, 1011.6, 1011.6, 1011.6, 1011.9, 1012.3, 
    1012.8, 1013.1, 1013.6, 1013.7, 1013.9, 1013.7, 1013.9, 1013.9, 1013.9, 
    1013.8, 1013.8, 1014.1, 1013.8, 1013.6, 1013.7, 1013.9, 1013.7, 1013.7, 
    1013.6, 1013.6, 1013.6, 1013.6, 1013.9, 1014.1, 1014.3, 1014.6, 1014.9, 
    1015.1, 1015.3, 1015.9, 1015.9, 1016.4, 1016.8, 1016.9, 1017.2, 1017.4, 
    1017.9, 1018.2, 1018.2, 1018.2, 1018.5, 1018.8, 1018.8, 1018.9, 1019.1, 
    1019.4, 1019.3, 1019.5, 1019.5, 1019.6, 1019.4, 1019.4, 1019.2, 1019.1, 
    1019, 1019, 1019, 1018.9, 1018.7, 1018.7, 1018.5, 1018.3, 1018.2, 1018, 
    1017.8, 1017.8, 1017.8, 1017.8, 1017.8, 1017.6, 1017.5, 1017.7, 1017.7, 
    1017.8, 1017.9, 1017.9, 1017.9, 1018.1, 1018.3, 1018.4, 1018.6, 1018.8, 
    1019, 1019.2, 1019.4, 1019.8, 1020, 1020.3, 1020.6, 1020.8, 1021.1, 
    1021.5, 1021.8, 1022.2, 1022.4, 1022.5, 1022.8, 1022.8, 1022.9, 1022.9, 
    1023, 1023, 1023.2, 1023.5, 1023.7, 1023.6, 1023.7, 1023.8, 1023.9, 1024, 
    1023.9, 1024, 1024, 1024.2, 1024.3, 1024.5, 1024.6, 1024.7, 1024.7, 
    1024.9, 1024.8, 1025, 1024.8, 1024.8, 1024.8, 1024.7, 1024.8, 1024.8, 
    1024.8, 1024.8, 1024.8, 1024.8, 1024.8, 1024.8, 1024.8, 1024.8, 1024.7, 
    1024.7, 1024.7, 1024.9, 1025.1, 1025.1, 1025.1, 1025, 1025, 1025, 1024.8, 
    1024.6, 1024.7, 1024.7, 1024.6, 1024.4, 1024.2, 1024.1, 1024, 1023.7, 
    1023.6, 1023.3, 1023.3, 1023.1, 1022.8, 1022.5, 1022.3, 1022.3, 1022, 
    1021.8, 1021.5, 1021.3, 1021.2, 1021, 1021, 1020.7, 1020.5, 1020.3, 
    1020.3, 1019.8, 1019.5, 1019.4, 1019.1, 1018.9, 1018.7, 1018.5, 1018.3, 
    1018.3, 1018, 1017.8, 1017.5, 1017.4, 1017.3, 1017, 1016.8, 1016.7, 
    1016.8, 1016.8, 1016.8, 1016.8, 1016.8, 1016.8, 1016.7, 1016.7, 1016.7, 
    1016.6, 1016.6, 1016.6, 1016.5, 1016.6, 1016.8, 1016.6, 1016.8, 1016.7, 
    1016.9, 1016.9, 1016.9, 1017, 1017.2, 1017.2, 1017.2, 1017.1, 1017, 
    1017.1, 1017, 1016.9, 1016.9, 1017.1, 1017.1, 1017.1, 1017.2, 1017.1, 
    1017.1, 1017.1, 1017, 1017.1, 1017.1, 1017.1, 1017, 1017, 1017, 1017, 
    1016.9, 1016.9, 1016.7, 1016.6, 1016.3, 1016.1, 1015.6, 1015.3, 1015, 
    1014.8, 1014.5, 1014.3, 1014, 1013.6, 1013.2, 1013, 1012.8, 1012.5, 
    1012.2, 1011.8, 1011.5, 1011.3, 1011.1, 1010.7, 1010.5, 1010.5, 1010.4, 
    1010.2, 1009.9, 1009.6, 1009.4, 1009.3, 1009.2, 1009, 1008.8, 1008.7, 
    1008.5, 1008.4, 1008.1, 1007.9, 1007.8, 1007.8, 1007.5, 1007.3, 1007.4, 
    1007.4, 1007.5, 1007.4, 1007.4, 1007.4, 1007.5, 1007.7, 1007.8, 1007.8, 
    1007.7, 1007.5, 1007.6, 1007.7, 1007.9, 1007.9, 1008, 1008.1, 1008.2, 
    1008.4, 1008.4, 1008.7, 1008.9, 1009.1, 1009.3, 1009.5, 1009.8, 1010, 
    1010.1, 1010.5, 1010.8, 1011, 1011.2, 1011.6, 1012, 1012.4, 1012.6, 
    1013.2, 1013.7, 1014, 1014.4, 1014.7, 1014.7, 1014.9, 1015.5, 1015.9, 
    1016.1, 1016, 1016.3, 1016.3, 1016.7, 1016.7, 1017, 1017.2, 1017.3, 
    1017.4, 1017.4, 1017.3, 1017.3, 1017.3, 1017.1, 1017.2, 1017.1, 1017, 
    1017, 1016.9, 1016.8, 1016.5, 1016.4, 1016.2, 1016.2, 1016, 1015.9, 
    1016.1, 1016.4, 1016.4, 1016.6, 1016.6, 1016.7, 1016.7, 1016.7, 1016.8, 
    1016.6, 1016.7, 1016.6, 1016.4, 1016.4, 1016.6, 1016.5, 1016.3, 1016.2, 
    1016.1, 1016.2, 1015.9, 1015.8, 1015.8, 1015.8, 1015.9, 1015.8, 1016.1, 
    1016.3, 1016.5, 1016.5, 1016.6, 1016.7, 1016.7, 1016.9, 1016.9, 1016.8, 
    1017, 1017.3, 1017.5, 1017.6, 1017.9, 1018, 1018.2, 1018.4, 1018.3, 
    1018.3, 1018.3, 1018.3, 1018.6, 1018.8, 1018.9, 1019.1, 1019.3, 1019.1, 
    1019.2, 1019.2, 1019.2, 1019.1, 1019.1, 1019.1, 1019.1, 1019.4, 1019.4, 
    1019.4, 1019.4, 1019.3, 1019.1, 1019.3, 1019.4, 1019, 1019.1, 1019, 
    1018.9, 1018.8, 1019, 1019, 1019.2, 1019.3, 1019.3, 1019.4, 1019.5, 
    1019.6, 1019.7, 1019.9, 1020.1, 1020.3, 1020.5, 1021.1, 1021.4, 1021.8, 
    1021.9, 1022.2, 1022.5, 1022.8, 1023, 1023.5, 1023.9, 1024.3, 1024.8, 
    1025.1, 1025.2, 1025.5, 1025.5, 1025.5, 1025.7, 1025.7, 1025.8, 1025.9, 
    1026, 1026.1, 1026.3, 1026.5, 1026.7, 1026.9, 1027.2, 1027.4, 1027.4, 
    1027.4, 1027.3, 1027.4, 1027.7, 1027.9, 1028.2, 1028.5, 1028.3, 1028.4, 
    1028.5, 1028.4, 1028.5, 1028.4, 1028.3, 1028.2, 1028.2, 1028.1, 1028.5, 
    1028.4, 1028.3, 1028.3, 1028, 1027.7, 1027.2, 1027, 1026.5, 1026.2, 
    1025.6, 1025.3, 1025, 1024.8, 1024.4, 1024.1, 1023.8, 1023.2, 1022.8, 
    1022.6, 1022.1, 1022, 1021.5, 1021.2, 1021.3, 1020.6, 1020, 1019.7, 
    1019.1, 1018.3, 1017.6, 1016.8, 1016.2, 1015.5, 1014.8, 1014.3, 1013.4, 
    1012.6, 1011.9, 1011.5, 1011.1, 1010.8, 1010.4, 1010, 1009.6, 1009.4, 
    1009.4, 1009.3, 1009.6, 1009.8, 1009.9, 1010.4, 1010.5, 1010.5, 1010.7, 
    1010.7, 1010.8, 1010.8, 1010.6, 1010.6, 1010.6, 1010.1, 1009.8, 1009.3, 
    1008.9, 1008.3, 1007.8, 1007.5, 1007.1, 1006.8, 1006.4, 1006.2, 1006, 
    1006.3, 1006.3, 1006.6, 1007.1, 1007.3, 1007.8, 1008.2, 1008.2, 1008.9, 
    1009.3, 1009.8, 1010.5, 1010.9, 1011.6, 1011.7, 1012.1, 1012.5, 1012.9, 
    1013.1, 1013.5, 1013.6, 1014, 1014.3, 1014.8, 1015.1, 1015.6, 1015.9, 
    1016.2, 1016.5, 1016.7, 1016.7, 1016.7, 1016.8, 1017, 1017.2, 1017.5, 
    1017.9, 1018, 1018, 1018.3, 1018.3, 1018.4, 1018.5, 1018.4, 1018.5, 
    1018.8, 1019, 1019.1, 1019.2, 1019.6, 1019.8, 1019.8, 1019.9, 1019.9, 
    1019.8, 1019.9, 1019.8, 1019.7, 1019.7, 1019.9, 1020.2, 1020.4, 1020.5, 
    1020.6, 1020.5, 1020.3, 1020.4, 1020.3, 1020.4, 1020.5, 1020.6, 1020.7, 
    1021, 1021.1, 1021.3, 1021.3, 1021.7, 1021.8, 1021.8, 1021.8, 1021.8, 
    1021.7, 1021.9, 1022.1, 1022.3, 1022.5, 1022.4, 1022.4, 1022.4, 1022.3, 
    1022.2, 1022, 1021.9, 1022, 1022, 1021.9, 1021.9, 1021.8, 1021.9, 1021.7, 
    1021.1, 1020.8, 1020.1, 1019.4, 1019, 1018.6, 1018.5, 1018.4, 1017.9, 
    1017.3, 1017.1, 1017, 1016.7, 1016.2, 1015.6, 1015.1, 1015, 1014.7, 
    1014.3, 1014.1, 1013.8, 1013.6, 1013.6, 1013.8, 1013.7, 1013.4, 1013.4, 
    1013.1, 1013.2, 1013.2, 1013.2, 1013.3, 1013.3, 1013.5, 1013.5, 1013.7, 
    1013.6, 1013.5, 1013.6, 1013.6, 1013.6, 1013.7, 1014, 1014.3, 1014.6, 
    1014.7, 1015, 1015.1, 1015.3, 1015.6, 1015.9, 1015.9, 1016.1, 1016.4, 
    1016.7, 1017.1, 1017.3, 1017.6, 1017.5, 1017.5, 1017.5, 1017.5, 1017.6, 
    1017.8, 1017.8, 1018, 1018.3, 1018.8, 1018.9, 1019, 1019.3, 1019.6, 
    1019.8, 1019.8, 1019.8, 1019.8, 1020, 1019.8, 1019.8, 1019.8, 1019.3, 
    1019.1, 1018.8, 1018.5, 1017.7, 1017, 1016.2, 1016, 1015.9, 1016, 1016.2, 
    1016.4, 1016.3, 1016, 1016, 1015.9, 1015.6, 1015.5, 1015.1, 1014.9, 
    1014.5, 1014.3, 1014.4, 1014.5, 1014.4, 1014.5, 1014.6, 1014.8, 1014.9, 
    1014.9, 1015.1, 1015.3, 1015.4, 1015.6, 1016, 1016.1, 1016.3, 1016.3, 
    1016, 1015.9, 1015.8, 1015.8, 1015.5, 1015.1, 1015.1, 1014.9, 1014.8, 
    1014.8, 1014.8, 1015, 1015, 1015.2, 1015.1, 1015.4, 1015.8, 1016, 1016.2, 
    1016.6, 1017, 1017.5, 1017.8, 1018, 1018.2, 1018.5, 1018.9, 1019.2, 
    1019.4, 1019.5, 1019.8, 1020, 1020.2, 1020.4, 1020.6, 1020.7, 1020.6, 
    1020.4, 1020, 1019.6, 1019.1, 1018.8, 1018.2, 1017.9, 1017.5, 1017, 
    1016.5, 1015.9, 1015.4, 1014.8, 1014.3, 1013.7, 1013.1, 1012.4, 1012.2, 
    1011.8, 1011.5, 1011, 1010.5, 1010.2, 1009.7, 1009.4, 1009.1, 1008.9, 
    1008.7, 1008.6, 1008.5, 1008.2, 1008.2, 1008.1, 1007.9, 1007.7, 1007.7, 
    1007.3, 1006.9, 1006.5, 1005.9, 1005.3, 1004.9, 1004.9, 1004.8, 1004.7, 
    1004.4, 1004.2, 1004.3, 1004.4, 1004.3, 1004.3, 1004.7, 1004.7, 1005.1, 
    1005.2, 1005.9, 1006.5, 1007, 1007.5, 1008.1, 1008.9, 1009.6, 1010.2, 
    1010.7, 1011.1, 1011.3, 1011.8, 1012, 1012.1, 1012, 1012.4, 1012.2, 1012, 
    1011.7, 1011.4, 1011.3, 1011, 1010.7, 1010.6, 1010.4, 1010.1, 1009.9, 
    1009.7, 1009.6, 1009.5, 1009.3, 1009.1, 1009, 1008.9, 1008.7, 1008.6, 
    1008.6, 1008.7, 1008.8, 1008.8, 1008.9, 1009.1, 1009.2, 1009.4, 1009.4, 
    1009.3, 1009.3, 1009.4, 1009.8, 1010, 1010.2, 1010.4, 1010.5, 1010.6, 
    1010.4, 1010.6, 1010.6, 1010.6, 1010.6, 1010.7, 1010.8, 1011, 1011.1, 
    1011.4, 1011.7, 1011.8, 1011.6, 1011.4, 1011.4, 1011.5, 1011.6, 1011.5, 
    1011.7, 1011.6, 1011.7, 1011.6, 1011.5, 1011.5, 1011.4, 1011.4, 1011.4, 
    1011.4, 1011.5, 1011.7, 1011.9, 1012.1, 1012.4, 1012.7, 1012.8, 1013, 
    1013, 1013, 1013.2, 1013.4, 1013.5, 1013.6, 1013.8, 1014, 1014.3, 1014.4, 
    1014.5, 1014.7, 1014.6, 1014.6, 1014.6, 1014.5, 1014.5, 1014.7, 1014.8, 
    1014.9, 1014.9, 1015.1, 1014.9, 1014.9, 1014.8, 1014.6, 1014.6, 1014.3, 
    1014.2, 1014.1, 1014.2, 1014.2, 1014.2, 1014.2, 1014.3, 1014, 1014, 
    1013.9, 1013.8, 1013.7, 1013.6, 1013.4, 1013.5, 1013.3, 1013.2, 1013.1, 
    1012.7, 1012.3, 1011.9, 1011.6, 1011.2, 1010.9, 1010.1, 1009.4, 1009, 
    1008.8, 1008.5, 1008.2, 1008, 1007.6, 1007.2, 1006.9, 1006.3, 1005.8, 
    1005.3, 1004.9, 1004.4, 1004, 1003.7, 1003.2, 1002.8, 1002.5, 1002.1, 
    1001.6, 1001.3, 1001.1, 1000.6, 1000.4, 1000.2, 1000, 999.8, 999.9, 
    999.9, 1000.1, 999.8, 999.7, 999.6, 999.6, 999.8, 999.8, 999.9, 1000, 
    1000.1, 1000.2, 1000.5, 1000.6, 1000.8, 1000.9, 1001, 1001.1, 1001.3, 
    1001.5, 1001.8, 1001.9, 1002.1, 1002.5, 1002.7, 1002.9, 1003.1, 1003.5, 
    1003.6, 1004, 1004.3, 1004.4, 1005.1, 1005.6, 1006.1, 1006.3, 1006.9, 
    1007.8, 1008.3, 1008.8, 1009.2, 1009.7, 1010, 1010.5, 1010.9, 1011.3, 
    1011.8, 1012.3, 1012.6, 1012.7, 1012.7, 1012.8, 1012.7, 1012.7, 1012.7, 
    1012.6, 1012.7, 1013.1, 1013.4, 1013.5, 1013.6, 1013.7, 1013.9, 1014, 
    1014.1, 1014.1, 1013.6, 1013.8, 1014, 1014.3, 1014.6, 1014.8, 1015, 
    1015.1, 1015.3, 1015.3, 1015.3, 1015.3, 1016.2, 1016.3, 1015.9, 1015.9, 
    1016.4, 1015.9, 1015.8, 1016.5, 1016.7, 1016.6, 1016.6, 1016.6, 1016.8, 
    1017, 1017.2, 1017.4, 1017.7, 1018.1, 1018.3, 1018.4, 1018.5, 1018.6, 
    1018.8, 1018.9, 1019.3, 1019.5, 1018.5, 1018.7, 1018.8, 1019.2, 1019.3, 
    1019.4, 1019.4, 1019.2, 1019.1, 1019.2, 1019.2, 1019, 1019, 1019.1, 
    1019.2, 1019.2, 1018.9, 1018.9, 1018.9, 1018.9, 1018.7, 1018.6, 1018.5, 
    1018.4, 1018.4, 1018.6, 1018.7, 1018.9, 1018.8, 1018.5, 1018.4, 1018, 
    1017.7, 1017.4, 1017.3, 1017.6, 1017.9, 1018, 1018.2, 1018.3, 1018.5, 
    1018.6, 1018.7, 1018.7, 1018.8, 1019.1, 1019.5, 1019.9, 1020.2, 1020.5, 
    1020.7, 1021, 1021, 1021, 1021, 1021, 1020.9, 1020.7, 1020.5, 1020.4, 
    1020.6, 1020.5, 1020.4, 1020.3, 1021, 1020.9, 1019.6, 1019.3, 1019, 
    1018.7, 1018.5, 1018.4, 1018.4, 1018.3, 1018.1, 1017.8, 1017.6, 1017.4, 
    1017.3, 1017.1, 1016.9, 1016.7, 1016.7, 1016.7, 1016.8, 1016.7, 1016.6, 
    1016.7, 1016.7, 1016.9, 1017, 1017.2, 1017.7, 1017.6, 1017.8, 1018.1, 
    1018.3, 1019.1, 1019.4, 1019.7, 1019.9, 1020.3, 1020.7, 1021, 1021.3, 
    1021.5, 1021.4, 1021.5, 1020.9, 1021.1, 1021.3, 1021.5, 1021.3, 1021, 
    1020.9, 1020.8, 1020.7, 1020.6, 1020.4, 1020.3, 1020, 1020, 1019.8, 
    1019.5, 1019.4, 1019.2, 1019, 1018.6, 1018.1, 1017.8, 1017.5, 1017.3, 
    1017.3, 1017.2, 1017.2, 1017.2, 1017.2, 1016.6, 1016.5, 1016.3, 1016.1, 
    1015.9, 1015.9, 1015.8, 1015.6, 1015.5, 1015, 1014.8, 1014.7, 1014.8, 
    1014.5, 1014.2, 1013.9, 1013.6, 1013.5, 1013.5, 1013.3, 1013.2, 1013.2, 
    1013.1, 1012.9, 1012.5, 1012.2, 1012.1, 1012, 1011.7, 1011.7, 1011.6, 
    1011.5, 1011.4, 1011.6, 1011.3, 1011, 1011, 1010.9, 1010.7, 1010.5, 
    1010.2, 1010.2, 1010.1, 1010.2, 1010.2, 1010, 1009.6, 1009.3, 1010.9, 
    1010.8, 1010.6, 1010.2, 1009.9, 1009.7, 1008.1, 1008.1, 1008.1, 1007.7, 
    1007.7, 1007.5, 1007.3, 1007.1, 1007, 1006.8, 1006.8, 1006.7, 1006.7, 
    1006.7, 1006.5, 1006.8, 1006.8, 1006.8, 1006.8, 1006.9, 1007, 1007, 
    1006.9, 1006.9, 1006.9, 1007.1, 1007.1, 1007.1, 1007.1, 1007.1, 1007, 
    1007, 1007.2, 1007.3, 1007.4, 1007.4, 1007.6, 1007.9, 1007.9, 1007.8, 
    1007.8, 1007.6, 1007.6, 1007.6, 1007.7, 1007.7, 1007.8, 1007.9, 1008, 
    1008, 1008.3, 1008.5, 1008.6, 1008.7, 1008.7, 1008.9, 1009, 1009.2, 
    1009.4, 1009.7, 1009.9, 1010.1, 1010.2, 1010.1, 1010.3, 1010.6, 1010.5, 
    1010.9, 1011.2, 1011.4, 1011.7, 1011.8, 1011.8, 1011.6, 1011.6, 1011.6, 
    1011.9, 1011.9, 1011.7, 1011.5, 1011.5, 1011.4, 1011.2, 1011.3, 1011.3, 
    1011.3, 1011.6, 1011.6, 1011.4, 1011.8, 1011.5, 1011.3, 1011.3, 1010.9, 
    1010.6, 1010.4, 1010.5, 1010.4, 1010.1, 1010, 1009.7, 1009.6, 1009.6, 
    1009.6, 1009.6, 1009.7, 1009.4, 1009.4, 1009.3, 1009.3, 1009.2, 1009.2, 
    1009.1, 1008.8, 1008.6, 1008.6, 1008.5, 1008.3, 1008.3, 1007.9, 1007.8, 
    1007.8, 1007.7, 1008, 1008, 1007.8, 1007.7, 1007.6, 1007.4, 1007.4, 
    1008.3, 1008.1, 1008.2, 1008.3, 1008.5, 1008.8, 1009.2, 1009.6, 1008.6, 
    1008.7, 1008.8, 1009, 1009.3, 1009.6, 1009.9, 1010.2, 1010.4, 1010.6, 
    1010.9, 1011.3, 1011.5, 1011.9, 1011.9, 1011.9, 1012.4, 1013, 1013.3, 
    1014.8, 1015, 1015.3, 1015.6, 1015.6, 1014.7, 1014.7, 1014.6, 1014.6, 
    1014.5, 1014.5, 1014.5, 1014.4, 1014.4, 1014.2, 1014.1, 1013.8, 1013.6, 
    1013.7, 1013.5, 1013.3, 1012.9, 1012.9, 1013, 1013, 1012.9, 1012.9, 
    1012.8, 1012.9, 1012.8, 1012.4, 1012, 1013, 1012.5, 1012.1, 1011.1, 1011, 
    1011.6, 1010.7, 1010.6, 1010.4, 1010, 1009.7, 1009.5, 1010, 1009.9, 
    1008.8, 1008.8, 1008.9, 1008.8, 1008.8, 1008.9, 1008.9, 1008.7, 1008.5, 
    1008, 1007.8, 1007.2, 1007, 1006.9, 1006.9, 1007, 1007, 1006.7, 1006.5, 
    1006.5, 1006.5, 1007.2, 1007.1, 1007, 1006.7, 1006.9, 1007.1, 1006.9, 
    1006.8, 1006.7, 1006.6, 1006.7, 1006.9, 1006.8, 1007, 1007.2, 1007.5, 
    1007.9, 1008.1, 1008.3, 1008.4, 1008.5, 1008.7, 1008.6, 1008.7, 1008.9, 
    1010.7, 1010.9, 1010.3, 1010.6, 1011, 1010.3, 1010.6, 1010.9, 1011.2, 
    1011.4, 1011.5, 1011.8, 1012, 1012, 1012.2, 1012.4, 1012.6, 1012.7, 
    1012.9, 1013.1, 1013.3, 1013.4, 1013.6, 1014, 1014.2, 1014.4, 1014.9, 
    1015.2, 1015.6, 1015.9, 1016.2, 1016.4, 1016.8, 1017.1, 1017.2, 1017.2, 
    1017.2, 1017.5, 1017.7, 1017.9, 1018, 1018.2, 1018.3, 1018.5, 1018.6, 
    1018.6, 1018.4, 1018.4, 1018.4, 1018.4, 1018.5, 1018.6, 1018.8, 1019.1, 
    1018.9, 1018.9, 1019.1, 1019, 1018.9, 1018.8, 1018.7, 1018.6, 1018.5, 
    1018.6, 1018.7, 1018.7, 1018.6, 1018.6, 1018.5, 1018.3, 1018.1, 1017.8, 
    1017.5, 1017.4, 1017.3, 1017.4, 1017.4, 1017.4, 1017.4, 1018.3, 1018, 
    1017.2, 1017, 1016.8, 1016.6, 1016.4, 1016.2, 1016, 1015.9, 1015.7, 
    1015.5, 1015.2, 1014.9, 1014.7, 1014.3, 1013.9, 1013.4, 1013.1, 1012.8, 
    1012.3, 1011.8, 1011.3, 1010.9, 1010.5, 1010.2, 1010, 1009.2, 1008.9, 
    1008.8, 1008.1, 1007.9, 1007.7, 1007.4, 1006.9, 1006.8, 1006.7, 1006.3, 
    1006.1, 1005.9, 1005.6, 1005.3, 1005.6, 1005.7, 1005.5, 1005.3, 1005.1, 
    1004.8, 1004.9, 1004.7, 1004.8, 1004.9, 1004.9, 1005.2, 1005.6, 1006.3, 
    1006.7, 1006.9, 1007.1, 1007.3, 1007.5, 1007.8, 1007.8, 1008, 1008.2, 
    1008.6, 1009, 1009.4, 1009.9, 1010.6, 1011.4, 1011.8, 1012.4, 1013.2, 
    1013.6, 1013.9, 1014.3, 1014.5, 1014.6, 1014.5, 1014.5, 1014.4, 1014.4, 
    1014.1, 1013.8, 1013.1, 1012.4, 1011.8, 1010.9, 1010, 1009.2, 1008.2, 
    1007.6, 1007.5, 1006.4, 1006.9, 1007.3, 1007.7, 1008.1, 1008.5, 1008.6, 
    1009, 1009, 1009.4, 1009.7, 1010.3, 1010.5, 1010.6, 1010.6, 1010.8, 
    1010.8, 1010.8, 1010.7, 1010.8, 1010.6, 1010.4, 1010.1, 1010, 1010.1, 
    1010.2, 1010.2, 1010.1, 1010.3, 1010.2, 1010.2, 1010.5, 1010.4, 1010.5, 
    1010.9, 1011.1, 1011.2, 1011.4, 1011.7, 1011.9, 1012, 1012.2, 1012.1, 
    1012.3, 1012.2, 1012.4, 1012.5, 1012.6, 1012.6, 1013, 1013, 1013.1, 
    1013.1, 1012.9, 1012.7, 1012.6, 1012.5, 1012.3, 1012.3, 1012.2, 1012.2, 
    1012.4, 1012.3, 1012.2, 1012, 1011.5, 1011.1, 1011, 1011.1, 1010.7, 
    1010.6, 1010.5, 1010.4, 1010.2, 1010, 1009.9, 1009.9, 1009.8, 1009.8, 
    1009.5, 1009.5, 1009.4, 1009.2, 1009.1, 1009, 1009, 1009.1, 1009.1, 1009, 
    1008.9, 1008.8, 1008.7, 1008.6, 1009.1, 1009, 1008.9, 1008.7, 1008.7, 
    1008.8, 1008.7, 1008.5, 1007.6, 1007.5, 1007.5, 1007.4, 1007.4, 1007.5, 
    1007.7, 1007.9, 1008.3, 1008.5, 1009.4, 1009.6, 1009.8, 1009.9, 1010, 
    1010.2, 1010.3, 1009.3, 1009.5, 1009.9, 1010.1, 1010.3, 1010.5, 1010.6, 
    1010.8, 1010.9, 1011.1, 1011.2, 1011.2, 1011.4, 1011.5, 1011.8, 1012, 
    1012, 1012, 1011.8, 1011.6, 1011.9, 1011.6, 1011.3, 1011.3, 1010.8, 
    1010.5, 1010.2, 1009.9, 1009.8, 1009.5, 1008.9, 1008.3, 1007.6, 1007, 
    1006.5, 1005.8, 1005.6, 1005.2, 1004.8, 1004.5, 1003.9, 1003.1, 1002.4, 
    1001.7, 1001.1, 1000.3, 999.7, 999.4, 999.5, 999, 998.9, 998.9, 999.2, 
    999.3, 999.5, 999.8, 1000.6, 1001.2, 1002, 1003.4, 1004.3, 1005.4, 
    1006.5, 1007, 1007.8, 1008.3, 1009.3, 1010, 1010.5, 1011, 1011.4, 1012, 
    1012.6, 1013.1, 1013.2, 1013.8, 1014, 1014.2, 1014.2, 1014, 1014, 1014.1, 
    1013.9, 1013.9, 1013.8, 1013.6, 1013.3, 1013.3, 1012.9, 1012.6, 1012.1, 
    1011.4, 1011, 1010.6, 1010, 1009.3, 1008.5, 1007.9, 1006.9, 1006.1, 
    1005.2, 1004, 1002.8, 1001.6, 1000.5, 999.7, 999.2, 998.8, 998.5, 998.3, 
    998.1, 998, 997.9, 997.8, 997.8, 997.8, 997.7, 997.9, 998.2, 998.4, 
    998.6, 998.8, 999.4, 999.6, 999.6, 999.6, 999.7, 999.8, 1000, 1000.2, 
    1000.3, 1000.3, 1000.1, 1000.2, 1000.3, 1000.3, 1000.2, 1000.1, 1000, 
    999.9, 999.7, 999.7, 999.7, 999.7, 999.7, 999.7, 1000.4, 1000.5, 1000.5, 
    1000.4, 1000.3, 1000, 998.6, 998.3, 998, 997.7, 997.4, 997.3, 996.8, 
    996.8, 996.8, 996.9, 997.1, 997.4, 997.8, 998.4, 998.8, 999.2, 999.6, 
    1000.2, 1000.8, 1001.5, 1003.7, 1003.5, 1004.4, 1005.2, 1006, 1006.8, 
    1007.2, 1007.9, 1008.2, 1008.7, 1009, 1009.4, 1009.7, 1010, 1010.1, 
    1010.2, 1010.2, 1009.6, 1008.7, 1008.2, 1007.1, 1007.4, 1006.7, 1006, 
    1005.2, 1004.1, 1002.7, 1001.6, 1000.6, 999.2, 997.9, 997.5, 995.3, 994, 
    992, 990.4, 988.4, 986.5, 984.5, 983, 982.5, 982.4, 982.3, 982.2, 982.1, 
    982.3, 982.5, 983.3, 983.9, 984.7, 985.4, 986.7, 987.9, 989.4, 990.9, 
    991.8, 993.6, 996, 997.8, 999.6, 1000.9, 1002.1, 1003, 1003.7, 1004.5, 
    1005.1, 1005.9, 1006.8, 1007.3, 1008.2, 1008.9, 1009.5, 1010.2, 1011.2, 
    1011.9, 1011.9, 1012.7, 1013.1, 1013.6, 1014.6, 1015.1, 1016.2, 1016.5, 
    1016.7, 1017.3, 1017.5, 1017.7, 1017.7, 1017.8, 1017.6, 1017.5, 1017.4, 
    1017.2, 1017, 1016.6, 1016.2, 1015.9, 1015.3, 1014.4, 1013.6, 1013.1, 
    1012.3, 1011.6, 1011.3, 1010.9, 1010.4, 1009.9, 1009.2, 1008.6, 1007.8, 
    1006.9, 1006.4, 1005.7, 1005.2, 1005.1, 1004.9, 1004.7, 1004.5, 1003.9, 
    1003, 1002.2, 1001.4, 1000.7, 999.8, 999.8, 999.3, 999.2, 999, 999, 999, 
    998.5, 998.9, 999.5, 999, 998.7, 998.8, 999.2, 999.6, 1000, 1000.4, 
    1000.8, 1000.5, 1001.3, 1001.8, 1001.7, 1001.5, 1001.4, 1001.3, 1001.1, 
    1001.1, 1001.1, 1001.3, 1001.7, 1002, 1002.3, 1002.4, 1002.1, 1002.1, 
    1001.5, 1001.3, 1005.2, 1005.2, 1005.2, 1005.2, 1005, 1004.6, 1000.7, 
    1000.4, 1000.1, 999.8, 999.5, 999.3, 999.1, 998.9, 998.6, 998.5, 998.8, 
    999, 999.3, 999.7, 999.8, 999.8, 1000.1, 1000.2, 1000.6, 1000.7, 1001, 
    1001.6, 1001.8, 1001.9, 1002.1, 1002.3, 1002.6, 1002.9, 1003.2, 1003.5, 
    1003.8, 1004.3, 1004.5, 1004.8, 1005, 1005.1, 1005.7, 1005.9, 1006.1, 
    1007, 1007.6, 1008, 1008.3, 1008.5, 1008.6, 1008.5, 1008.6, 1009, 1009.2, 
    1009.6, 1010, 1010.6, 1010.8, 1010.9, 1011.8, 1011.7, 1011.9, 1012.3, 
    1012.8, 1013.2, 1013, 1013.7, 1014.1, 1014.5, 1015.1, 1015.6, 1015.9, 
    1016.4, 1016.9, 1017.2, 1017.7, 1018.2, 1018.8, 1019.4, 1019.9, 1021.7, 
    1021.9, 1021.9, 1021.4, 1021.8, 1022, 1021.7, 1022.1, 1022.4, 1022.4, 
    1022.6, 1022.5, 1022.6, 1022.6, 1022.3, 1022.1, 1022, 1022, 1021.4, 
    1021.2, 1021, 1020.8, 1020.8, 1020.6, 1020.2, 1019.8, 1019.8, 1019.4, 
    1019.3, 1019.3, 1019.5, 1019.7, 1019.8, 1020, 1020.1, 1020.3, 1020.4, 
    1020.1, 1020, 1019.9, 1019.8, 1019.6, 1019.4, 1019.4, 1019.4, 1019.3, 
    1019.1, 1018.9, 1018.6, 1018.3, 1018, 1017.8, 1017.5, 1017.2, 1016.9, 
    1016.9, 1016.8, 1016.8, 1016.7, 1016.4, 1016, 1015.2, 1014.7, 1013.9, 
    1013.7, 1013.5, 1012.8, 1012.5, 1012.1, 1011.9, 1011.6, 1011.4, 1010.5, 
    1010, 1009.4, 1009.1, 1008.8, 1008.3, 1007.8, 1007.4, 1007.2, 1007.1, 
    1006.7, 1006.2, 1005.5, 1005.2, 1004.7, 1004, 1003.2, 1002.4, 1001.7, 
    1000.8, 1000.1, 999.2, 998.4, 997.5, 996.5, 996.5, 994.4, 993.3, 992.6, 
    991.6, 990.6, 990, 989.2, 988.5, 988.2, 987.9, 987.5, 987.1, 987, 986.5, 
    986, 985.8, 985.6, 985.5, 985.3, 985.1, 985, 984.8, 984.7, 984.7, 985, 
    985.4, 985.8, 986.2, 986.4, 986.9, 987, 987.1, 987.8, 988.7, 989.2, 
    989.5, 989.9, 991.2, 990.7, 991.2, 991.7, 992.2, 992.6, 993, 993.3, 
    993.6, 994.1, 994.5, 994.6, 994.9, 995.1, 995.2, 995.4, 995.5, 995.8, 
    996.1, 996.9, 996.8, 997.1, 997, 997.2, 997.3, 997.7, 997.8, 997.9, 
    997.9, 998.2, 999.1, 998.8, 999.1, 999.2, 999.2, 999.5, 999.7, 999.9, 
    1000.2, 1000.6, 1001.1, 1001.5, 1002, 1002.4, 1002.9, 1003.4, 1004, 
    1004.5, 1005.1, 1005.5, 1005.9, 1006.4, 1007, 1007.5, 1008, 1008.7, 
    1009.4, 1009.8, 1010.5, 1011.2, 1011.8, 1012.7, 1013, 1013.3, 1013.5, 
    1013.3, 1013.4, 1013.3, 1012.9, 1012.7, 1012.7, 1013, 1014.8, 1014.1, 
    1014.6, 1014.8, 1015.1, 1015.4, 1015.7, 1016.1, 1016.1, 1016.2, 1016.3, 
    1017.6, 1017.6, 1017.4, 1017.5, 1017, 1016.3, 1016.2, 1015.8, 1015.4, 
    1015, 1014.5, 1014.1, 1013.1, 1012.6, 1011.9, 1011, 1010.2, 1009.3, 
    1008.5, 1007.6, 1006.7, 1005.7, 1004.7, 1003.6, 1002.5, 1001.5, 1000.9, 
    1000.5, 1000.4, 1000.7, 1001, 1000.9, 1001.3, 1001.8, 1002.3, 1002.6, 
    1002.9, 1003.2, 1004.6, 1003.9, 1004.3, 1004.8, 1006.2, 1006.2, 1007, 
    1007.9, 1008.7, 1009.5, 1011, 1011, 1011.8, 1012.6, 1013.4, 1014.1, 
    1014.7, 1015.7, 1016.3, 1016.8, 1017.2, 1017.7, 1017.9, 1017.6, 1017.4, 
    1017.5, 1017.4, 1017.3, 1017.4, 1017.5, 1017.5, 1016.9, 1016.2, 1015.9, 
    1015.5, 1014.8, 1014, 1013.5, 1012.7, 1012.9, 1013.3, 1012.9, 1013, 
    1012.9, 1012.7, 1012.8, 1012.5, 1012.9, 1012.7, 1012.8, 1012.9, 1013.1, 
    1013.3, 1013.6, 1013.8, 1013.9, 1014.6, 1015.4, 1016, 1016.5, 1017.5, 
    1017.6, 1017.7, 1018.1, 1018.3, 1018.4, 1018.3, 1018, 1016.9, 1016.4, 
    1015.1, 1013.4, 1012.5, 1011.9, 1011.7, 1012.4, 1013.6, 1014.5, 1015.7, 
    1016.9, 1018.1, 1019.1, 1019.9, 1020.9, 1021.9, 1022.8, 1023.3, 1024.2, 
    1024.9, 1025.9, 1026.7, 1027.4, 1028, 1028.3, 1028.6, 1029, 1029.6, 
    1030.3, 1030.7, 1031.3, 1031.9, 1032.5, 1032.8, 1033.1, 1033.5, 1033.9, 
    1034, 1033.8, 1033.8, 1034.2, 1034.6, 1034.9, 1035.2, 1035.4, 1035.6, 
    1035.9, 1036.3, 1036.6, 1036.7, 1036.6, 1037, 1037.1, 1036.9, 1037.7, 
    1037.5, 1036.8, 1037, 1037.1, 1037.1, 1037.1, 1036.9, 1036.9, 1036.7, 
    1036.5, 1036.5, 1036.5, 1036.4, 1036.5, 1036.3, 1036, 1035.9, 1035.8, 
    1035.5, 1035.3, 1035.2, 1034.9, 1034.6, 1034.2, 1034, 1033.8, 1033.4, 
    1033.1, 1032.8, 1032.3, 1031.7, 1031.2, 1030.8, 1031.2, 1030, 1029.7, 
    1029.4, 1029, 1028.6, 1028.3, 1027.8, 1027.2, 1026.7, 1026.1, 1025.6, 
    1025.2, 1024.9, 1024.9, 1024.6, 1023.8, 1023.4, 1023, 1022.6, 1022, 
    1021.3, 1020.8, 1020.3, 1020, 1020, 1019.9, 1019.6, 1019.5, 1019.6, 
    1019.6, 1019.4, 1019.1, 1019.2, 1019.2, 1019, 1019.3, 1019.5, 1019.7, 
    1019.7, 1020.1, 1020.4, 1020.4, 1020.2, 1020.1, 1020.1, 1019.9, 1019.8, 
    1019.9, 1019.9, 1019.7, 1019.7, 1019.7, 1019.7, 1019.5, 1019.5, 1019.3, 
    1019.2, 1019, 1019, 1018.9, 1018.9, 1018.7, 1018.5, 1018.4, 1018.1, 
    1017.6, 1017.3, 1017.3, 1016.7, 1016.3, 1016, 1015.6, 1015.4, 1014.9, 
    1014.6, 1014.2, 1014.1, 1014.2, 1014, 1014.1, 1014, 1014.3, 1014.5, 
    1014.7, 1014.9, 1015.3, 1015.6, 1015.8, 1015.8, 1016, 1016.3, 1016.3, 
    1016.3, 1016.2, 1016.2, 1016.1, 1016, 1016.1, 1016.4, 1016.5, 1016.7, 
    1016.9, 1017.2, 1017.3, 1017.6, 1017.7, 1018, 1018.3, 1018.5, 1018.7, 
    1018.9, 1019.1, 1019.2, 1019.4, 1019.3, 1019.3, 1019.2, 1019.4, 1019.2, 
    1019.2, 1019.2, 1019.2, 1019.4, 1019.6, 1019.7, 1019.8, 1019.8, 1019.8, 
    1019.8, 1019.8, 1019.9, 1020.1, 1020.3, 1020.5, 1020.7, 1021.4, 1022, 
    1022.7, 1023.2, 1023.4, 1023.6, 1023.9, 1024.1, 1024.1, 1024.1, 1024.2, 
    1024.4, 1024.3, 1024.4, 1024.4, 1024.2, 1023.9, 1023.7, 1023.4, 1023, 
    1022.6, 1022.5, 1022.4, 1022, 1021.5, 1022.3, 1022, 1020.5, 1020.1, 
    1019.8, 1019.5, 1019, 1018.7, 1018.5, 1018.2, 1018, 1017.9, 1017.6, 
    1017.3, 1017.1, 1016.9, 1016.3, 1016.1, 1015.8, 1015.5, 1015.4, 1015, 
    1015.6, 1014.3, 1013.9, 1013.6, 1013, 1012.7, 1012.2, 1012, 1011.9, 
    1011.7, 1011.6, 1011.7, 1011.9, 1012.3, 1012.5, 1012.8, 1013.2, 1013.7, 
    1013.9, 1014.1, 1014.3, 1014, 1014.8, 1015.1, 1015.4, 1015.7, 1015.9, 
    1016, 1016.2, 1016.5, 1016.7, 1016.9, 1017, 1018.6, 1017.5, 1017.7, 1018, 
    1018.2, 1018.6, 1018.8, 1019, 1019.2, 1019.3, 1019.3, 1020.6, 1020.6, 
    1021.1, 1020.9, 1020.4, 1020, 1019.8, 1018.2, 1018, 1017.8, 1017.6, 
    1017.1, 1016.6, 1016.3, 1016.1, 1015.8, 1015.9, 1015.7, 1015.7, 1015.6, 
    1015.5, 1015.3, 1015.3, 1015.3, 1015.3, 1017.5, 1016.9, 1017, 1016.9, 
    1015.2, 1015.3, 1015.3, 1015.2, 1015.1, 1014.8, 1014.6, 1014.5, 1014.4, 
    1014.4, 1014.3, 1014.3, 1014.7, 1015, 1015.1, 1015.2, 1015.2, 1015.3, 
    1015.5, 1015.5, 1015.6, 1015.7, 1015.8, 1016, 1016.1, 1016.3, 1016.5, 
    1016.5, 1016.3, 1016.1, 1016.4, 1016.4, 1016.3, 1016.1, 1016.4, 1016.7, 
    1016.9, 1017.2, 1017.4, 1017.7, 1017.8, 1017.6, 1019, 1017.2, 1017, 
    1016.6, 1018.4, 1018.1, 1015.9, 1015.6, 1015.6, 1015.2, 1014.9, 1014.5, 
    1013.9, 1013.7, 1013.3, 1012.9, 1012.6, 1013.1, 1012.9, 1012, 1011.8, 
    1011.5, 1011.1, 1010.5, 1010.1, 1009.7, 1009.2, 1008.8, 1008.5, 1009.4, 
    1009.1, 1008.8, 1008.7, 1008.3, 1008, 1007.6, 1006.4, 1006.2, 1006, 
    1005.7, 1005.2, 1005.8, 1005.9, 1006.2, 1006.7, 1007.1, 1007.1, 1007, 
    1007, 1007, 1007, 1007.2, 1007.1, 1006.9, 1006.6, 1006.6, 1006.1, 1006.9, 
    1006.6, 1004.7, 1004.2, 1003.7, 1003.5, 1003.2, 1003, 1003.1, 1003.5, 
    1003.5, 1003.4, 1003.2, 1003, 1003, 1004.1, 1003.1, 1003.2, 1003.4, 
    1003.4, 1003.5, 1003.7, 1003.6, 1003.3, 1003.1, 1003, 1002.3, 1002.4, 
    1001.7, 1001.4, 1001.9, 1002, 1002, 1002.1, 1002.2, 1002.3, 1002.7, 
    1002.8, 1003.2, 1003.6, 1004, 1004.1, 1004.8, 1005, 1005.2, 1005.3, 
    1005.4, 1005.4, 1005.4, 1004.8, 1004.2, 1003.6, 1003.1, 1002.3, 1001.6, 
    1001.1, 1000.6, 1000.1, 1000.1, 999.4, 999.1, 998.8, 998.4, 998.2, 997.8, 
    997.5, 998.4, 997, 996.6, 996.2, 995.8, 995.3, 995, 994.9, 994.6, 994.2, 
    994, 995.3, 993.8, 993.6, 993.5, 993.4, 993.4, 993.4, 993.8, 994.1, 
    994.2, 994.3, 996.2, 996.6, 996.6, 995.4, 995.8, 996.4, 996.8, 997.3, 
    997.8, 998.3, 999, 999.5, 999.9, 1000.2, 1000.9, 1001.7, 1002.5, 1003.2, 
    1003.7, 1004.3, 1004.6, 1005.1, 1005.3, 1005.5, 1006, 1006.1, 1006.7, 
    1007.2, 1007.5, 1008.1, 1008.3, 1009.2, 1009.3, 1009.5, 1008.6, 1008.6, 
    1008.5, 1008.4, 1008.3, 1008.6, 1008.9, 1009, 1009.3, 1009.3, 1009.6, 
    1009.7, 1009.7, 1010.1, 1010.1, 1010, 1010.2, 1010.4, 1010.6, 1010.7, 
    1010.9, 1011.3, 1011.6, 1011.8, 1012, 1012.1, 1012.3, 1012.7, 1013.2, 
    1013.6, 1014.1, 1014.7, 1015.3, 1015.5, 1015.9, 1016.1, 1016.4, 1016.6, 
    1016.7, 1016.8, 1017.1, 1017.2, 1017.4, 1017.7, 1017.9, 1017.9, 1017.9, 
    1018.1, 1018.1, 1018.1, 1018.1, 1018.1, 1018.3, 1018.3, 1018.6, 1018.7, 
    1018.6, 1018.5, 1018.5, 1018.2, 1017.9, 1017.5, 1017.2, 1016.9, 1016.7, 
    1016.4, 1016.3, 1016.1, 1015.6, 1015.2, 1014.9, 1014.5, 1014.2, 1013.9, 
    1013.6, 1013.4, 1013.2, 1013.2, 1013.1, 1012.8, 1012.4, 1012.5, 1012.1, 
    1011.8, 1011.6, 1011.1, 1010.6, 1010.3, 1009.9, 1009.7, 1009.4, 1009.1, 
    1008.7, 1008.4, 1007.8, 1007.4, 1007, 1006.6, 1006.2, 1005.9, 1005.6, 
    1005.1, 1005.1, 1004.9, 1004.8, 1004.5, 1004.2, 1003.8, 1003.6, 1003.6, 
    1003.6, 1003.4, 1003.3, 1003.4, 1003.3, 1003.2, 1002.9, 1002.8, 1002.7, 
    1002.5, 1002.5, 1002.4, 1002.3, 1002.3, 1002.6, 1002.6, 1002.8, 1002.7, 
    1002.9, 1002.8, 1003, 1003.2, 1003.3, 1003.4, 1003.6, 1003.8, 1004.4, 
    1004.9, 1005.3, 1005.6, 1005.9, 1006.1, 1006.1, 1006.1, 1006.3, 1006.5, 
    1006.8, 1006.8, 1006.5, 1006.7, 1006.6, 1006.6, 1006.4, 1006.2, 1006, 
    1006, 1005.7, 1005.3, 1005.3, 1005, 1004.7, 1004.1, 1003.8, 1003.3, 
    1002.8, 1002.4, 1001.9, 1001.4, 1001, 1000.3, 1000, 999.9, 999.6, 999.7, 
    999.8, 1000, 1000.1, 999.9, 1000.2, 1000.3, 1000.4, 1001, 1001.7, 1002.1, 
    1002.8, 1003.6, 1004.1, 1004.6, 1005.3, 1006.2, 1006.6, 1007, 1007.4, 
    1007.5, 1008, 1008.2, 1008.6, 1008.9, 1009.1, 1009.6, 1009.6, 1010, 
    1009.9, 1009.9, 1010.1, 1010.1, 1009.9, 1009.8, 1009.7, 1009.4, 1009.1, 
    1008.5, 1007.7, 1006.8, 1006.5, 1006.2, 1005.6, 1004.9, 1004.5, 1004.2, 
    1003.5, 1002.9, 1002.4, 1001.9, 1001.2, 1000.6, 999.9, 999, 997.7, 996.5, 
    995.5, 994.6, 993.4, 992.7, 991.9, 990.8, 989.7, 988.5, 987.6, 986.9, 
    986, 985.4, 984.5, 983.9, 984.1, 984.2, 984.1, 985.3, 986.2, 986.9, 
    987.3, 988.1, 988.8, 989.4, 990, 990.1, 990.4, 991.4, 992.1, 992.9, 
    993.8, 994.5, 995.2, 995.8, 996.9, 997.8, 998.5, 999.2, 1000.3, 1001, 
    1001.3, 1001.9, 1002.4, 1003, 1002.9, 1002.9, 1003.3, 1003.5, 1003.7, 
    1003.8, 1003.7, 1003.8, 1004.1, 1004.3, 1004.5, 1004.8, 1004.9, 1005.1, 
    1005.2, 1005.4, 1005.5, 1005.9, 1006.2, 1006.6, 1007.1, 1007.6, 1008.2, 
    1008.9, 1009.4, 1009.9, 1010.4, 1010.8, 1011.2, 1011.5, 1011.7, 1011.5, 
    1011.5, 1011.7, 1011.8, 1012, 1011.9, 1012, 1012, 1012.2, 1012.5, 1012.9, 
    1013.3, 1013.6, 1014.3, 1014.9, 1015.4, 1016, 1016.2, 1016.4, 1016.6, 
    1017, 1017.3, 1017.6, 1018, 1018.4, 1018.7, 1018.9, 1019.4, 1020, 1020.3, 
    1020.4, 1020.7, 1021.1, 1021.5, 1022, 1022.5, 1023.2, 1023.7, 1024.3, 
    1024.8, 1025.2, 1025.5, 1025.7, 1026.1, 1026.4, 1026.7, 1027, 1026.9, 
    1027.1, 1027.1, 1027.5, 1027.6, 1027.8, 1027.8, 1027.5, 1027.9, 1027.7, 
    1028, 1028.2, 1028.3, 1028.6, 1028.9, 1029.4, 1029.9, 1030.1, 1030.3, 
    1030.2, 1030.5, 1030.6, 1030.6, 1030.8, 1031.2, 1031.4, 1031.8, 1032, 
    1032.4, 1032.6, 1032.7, 1032.8, 1032.8, 1032.7, 1032.8, 1032.7, 1032.7, 
    1032.8, 1032.5, 1032.1, 1032, 1031.9, 1031.3, 1030.7, 1030.2, 1029.8, 
    1029, 1028.4, 1027.6, 1026.6, 1025.5, 1024.5, 1023.4, 1022, 1020.5, 
    1018.9, 1017, 1015.3, 1013.3, 1011.8, 1011, 1009.5, 1007.7, 1006.9, 
    1005.8, 1005.8, 1005.6, 1005.7, 1005.3, 1005.3, 1005.8, 1007, 1007.5, 
    1007.9, 1008.8, 1009.3, 1009.7, 1010.3, 1011.3, 1011.9, 1012.2, 1012.6, 
    1013.4, 1013.8, 1014.2, 1015, 1015.4, 1015.4, 1015.3, 1015.4, 1015.5, 
    1015.3, 1014.7, 1014.7, 1014.7, 1014.5, 1014.1, 1013.9, 1013.7, 1013.1, 
    1012.5, 1011.3, 1010.1, 1009.6, 1008.6, 1007.5, 1006.1, 1004.9, 1003.4, 
    1002.4, 1001.2, 1000.6, 1000.1, 999.5, 999.5, 999.6, 999.8, 999.7, 999.9, 
    1000, 1000.3, 1000.8, 1000.7, 1001.1, 1001.1, 1001.1, 1001, 1001.2, 
    1001.1, 1001.1, 1001.1, 1001.5, 1001.9, 1001.7, 1002, 1002.4, 1002.7, 
    1003, 1003.3, 1003.3, 1003.9, 1004.1, 1004.5, 1005.1, 1005.4, 1005.8, 
    1006.2, 1006.2, 1006.5, 1006.5, 1006.4, 1006.6, 1006.4, 1006.1, 1006.2, 
    1006.4, 1006.7, 1007, 1007.3, 1008.3, 1009, 1010.2, 1011.3, 1012.3, 
    1013.3, 1014.8, 1015.7, 1016.7, 1017.6, 1018.6, 1018.9, 1019.9, 1020.4, 
    1021.1, 1021, 1021.3, 1021.5, 1021.1, 1021.3, 1020.8, 1020.6, 1019.9, 
    1020.1, 1019.8, 1018.9, 1018.4, 1017.7, 1016.9, 1016, 1015.6, 1015.5, 
    1015.3, 1014.9, 1014.3, 1014.2, 1013.6, 1013.3, 1012.6, 1011.7, 1011.1, 
    1010.4, 1009.9, 1009, 1008.7, 1007.9, 1007.7, 1008.1, 1008, 1008.9, 
    1009.6, 1009.7, 1009.9, 1010.4, 1010.6, 1011.1, 1011.3, 1011.7, 1011.9, 
    1012.5, 1012.8, 1013, 1013.1, 1013.1, 1012.7, 1012.8, 1012.5, 1012.2, 
    1011.6, 1011.4, 1011.3, 1011.1, 1011.4, 1010.9, 1010.5, 1010.4, 1011.2, 
    1010.9, 1011.1, 1011.4, 1011.6, 1012, 1011.8, 1011.7, 1011.6, 1011.3, 
    1011.2, 1010.8, 1010.3, 1010.4, 1010.5, 1010.1, 1009.9, 1009.9, 1009.8, 
    1009.3, 1009.2, 1008.5, 1008.4, 1007.4, 1006.2, 1005.2, 1004.2, 1003.3, 
    1002.1, 1000.8, 999.6, 999.1, 998.1, 999.2, 1000.3, 1001.1, 1002.2, 
    1003.3, 1004.9, 1006.4, 1006, 1006.7, 1007.6, 1008.5, 1008.6, 1008.9, 
    1009.2, 1009.3, 1009.5, 1009.2, 1008.8, 1008.5, 1008, 1007.9, 1008.2, 
    1008, 1007.9, 1007.9, 1007.5, 1007.5, 1007.5, 1007.6, 1007.7, 1007.7, 
    1007.8, 1007.9, 1008.2, 1008.7, 1009, 1008.9, 1008.7, 1009.1, 1009.1, 
    1009.2, 1009.2, 1009, 1009.2, 1009.3, 1009.1, 1009.1, 1009.2, 1009.3, 
    1009.2, 1009.2, 1008.8, 1008.5, 1007.8, 1007.4, 1007.4, 1007.5, 1006.8, 
    1006.6, 1006.1, 1005.4, 1005.3, 1004.7, 1003.8, 1002.8, 1002.2, 1001.9, 
    1001.7, 1001.3, 1001.1, 1000.7, 1000.8, 1000.6, 1000.1, 999.2, 998.4, 
    997.7, 996.9, 996.3, 995.8, 995.6, 995.5, 994.8, 993.8, 993.1, 992.7, 
    992.1, 991.7, 991.7, 992.2, 992.7, 993.1, 993.9, 994.8, 995.5, 996.4, 
    997, 997.5, 997.6, 997.8, 997.9, 998, 997.4, 997.4, 996.8, 996.7, 996.2, 
    995.8, 995.9, 996.9, 998.1, 999.4, 1001.1, 1002.4, 1004.2, 1006, 1008.2, 
    1010.6, 1013.1, 1015.1, 1016.9, 1018.6, 1020, 1021.1, 1022.3, 1023.1, 
    1024, 1024.6, 1025.4, 1026.1, 1027, 1027.3, 1028.1, 1028.3, 1028.7, 
    1028.8, 1028.8, 1029.2, 1029.5, 1029.8, 1030.1, 1030.3, 1030.3, 1030.5, 
    1030.8, 1030.9, 1031.1, 1031, 1030.9, 1031.1, 1031.1, 1031.3, 1031.3, 
    1031.4, 1031.4, 1031.4, 1031.2, 1031.1, 1031.1, 1030.9, 1030.8, 1030.6, 
    1030, 1029.8, 1029.2, 1028.8, 1028.3, 1027.9, 1027.5, 1027.1, 1026.9, 
    1026.5, 1026.1, 1025.5, 1025.2, 1024.9, 1024.8, 1024.7, 1024.4, 1024.2, 
    1024.1, 1023.7, 1023.3, 1023, 1022.3, 1022.1, 1022.1, 1021.5, 1021.5, 
    1022.3, 1022, 1021.2, 1021.2, 1020.9, 1020.3, 1020.1, 1019.6, 1018.9, 
    1018.2, 1018, 1018.1, 1018.1, 1017.6, 1017.7, 1017.2, 1016.6, 1015.9, 
    1015.6, 1015.2, 1014.7, 1014.1, 1013.7, 1013.5, 1013.3, 1013, 1012.8, 
    1013, 1012.3, 1011.5, 1011.4, 1011.1, 1010.6, 1010.6, 1010.4, 1010.2, 
    1009.9, 1009.9, 1010.4, 1010.3, 1010.2, 1010.4, 1010.5, 1010.8, 1011, 
    1011.5, 1010.8, 1011, 1011.6, 1012.4, 1013, 1013.6, 1013.9, 1014.4, 
    1015.4, 1016, 1016.4, 1017.2, 1017.1, 1017.1, 1017.6, 1017.7, 1017.8, 
    1017.8, 1017.8, 1017.7, 1017.6, 1017.6, 1017.2, 1016.9, 1016.5, 1016.2, 
    1015.9, 1015.5, 1015.3, 1015, 1014.5, 1014, 1013.2, 1012.6, 1011.7, 
    1010.7, 1009.9, 1009.2, 1007.8, 1007, 1006.4, 1005.2, 1003.8, 1002.6, 
    1001.4, 1000.2, 998.9, 998, 996.4, 995.2, 994.2, 993.1, 992.3, 991.2, 
    990.4, 989.6, 988.8, 987.6, 986.6, 985.7, 984.8, 984.6, 983.4, 982.4, 
    982.1, 981.6, 981, 980.1, 979.6, 978.8, 978.3, 977.8, 977.2, 976.2, 
    975.7, 975.3, 974.6, 974.1, 973.8, 973.3, 973, 972.4, 971.6, 971.5, 
    971.5, 971.3, 971.9, 972.1, 972.2, 972.5, 973.2, 973.6, 974.2, 975.1, 
    975.2, 976.3, 976.7, 977.8, 978.7, 979.7, 980.4, 981.4, 982.1, 982.9, 
    983.2, 983.2, 983.6, 984.2, 985.1, 985.1, 985.4, 985.7, 986.2, 986.8, 
    987.3, 987.4, 987.2, 987.7, 987.7, 988, 988.1, 987.9, 988.2, 988.6, 
    988.7, 988.9, 989, 988.8, 988.8, 988.9, 988.7, 988.6, 988.4, 988.3, 
    988.4, 988.4, 988.5, 988.7, 988.8, 988.7, 988.7, 988.7, 988.8, 989.1, 
    989.2, 989.2, 989.6, 990, 990.1, 990.2, 990.3, 990.5, 990.4, 990.4, 
    990.1, 990.1, 990.2, 990.3, 990.6, 991.1, 991.6, 992.1, 992.5, 992.5, 
    992.7, 992.7, 992.7, 993, 993.3, 993.2, 993.3, 993.6, 993.6, 993.4, 
    993.1, 993.1, 992.7, 992, 991.6, 991.1, 990.6, 990, 989.8, 989.1, 988.4, 
    987.6, 986.4, 985.6, 984.7, 984, 982.7, 981.4, 979.9, 978.6, 978.4, 978, 
    977.8, 976.8, 976.4, 975.9, 975.2, 975.2, 974.9, 974.8, 974.7, 974.7, 
    974.7, 974.8, 974.9, 975, 975.1, 975, 974.8, 975.2, 975.2, 975, 975.1, 
    975.1, 975.2, 975, 974.9, 975, 974.8, 974.5, 974.4, 974.5, 974.7, 974.7, 
    974.6, 974.5, 974.9, 975.4, 975.7, 976.3, 977, 977.8, 978.6, 979.3, 
    979.9, 980.4, 980.9, 981.6, 982.2, 982.7, 983.2, 983.4, 983.6, 983.8, 
    984, 984, 984.3, 984.6, 985.1, 985.2, 985.7, 986.5, 987, 987.3, 987.4, 
    987.7, 988.1, 988.1, 988.1, 988.2, 988.1, 988, 988, 988.1, 988.1, 987.7, 
    987.7, 987.6, 987.6, 987.2, 987, 986.9, 986.8, 986.9, 986.6, 986.5, 
    986.3, 986.2, 986, 985.8, 985.7, 985.3, 985.1, 984.9, 984.5, 984.3, 
    983.9, 983.8, 983.4, 983.3, 983.3, 983.3, 983.1, 983.2, 983.1, 983, 983, 
    983, 983.1, 983.1, 982.9, 982.7, 982.7, 982.6, 982.8, 982.9, 982.9, 
    983.3, 983.5, 983.8, 984.2, 984.6, 985, 985.7, 986.4, 986.9, 987.2, 
    987.3, 987.6, 987.9, 988.4, 988.6, 989.2, 990.2, 991.1, 991.6, 992.2, 
    992.5, 993.1, 993.4, 993.9, 994.4, 995.2, 995.3, 995.9, 996.4, 996.7, 
    997.2, 997.5, 997.4, 997.9, 998, 998.2, 998.4, 998.6, 998.6, 998.9, 
    998.9, 999.1, 998.8, 998.7, 998.6, 998.1, 997.9, 997.8, 997.2, 996.8, 
    996.5, 996.4, 995.8, 995.6, 995.2, 994.6, 993.8, 993.4, 992.8, 992.4, 
    991.9, 991.6, 991.4, 991.7, 992.1, 993.1, 993.5, 994, 994.1, 994.2, 
    994.4, 994.5, 994.8, 994.9, 994.7, 994.4, 994.6, 994.7, 994.8, 995.1, 
    995.5, 995.6, 995.9, 996, 996.2, 996.5, 996.9, 997.3, 998, 998.6, 999.4, 
    999.5, 999.7, 1000.1, 1000.6, 1001, 1001.3, 1001.7, 1002.1, 1002.3, 
    1002.9, 1003.3, 1003.5, 1003.9, 1004.2, 1004.6, 1004.8, 1004.9, 1005.2, 
    1005.1, 1005.3, 1005.6, 1005.9, 1005.9, 1006.3, 1006.1, 1006.2, 1006.2, 
    1006.2, 1006.5, 1006.5, 1006.6, 1006.4, 1006.2, 1006.2, 1006.3, 1006.2, 
    1006.1, 1006.1, 1006.2, 1005.9, 1005.8, 1005.7, 1005.5, 1005.4, 1005.6, 
    1005.9, 1006, 1005.8, 1005.5, 1005.4, 1005.2, 1005.3, 1005.3, 1005.5, 
    1005.5, 1005.5, 1005.5, 1005.7, 1005.4, 1005.3, 1005.2, 1005.6, 1005.5, 
    1005.8, 1005.7, 1005.6, 1005.8, 1005.8, 1005.8, 1006.2, 1006.4, 1006.6, 
    1006.3, 1006.3, 1006.4, 1006.5, 1006.4, 1006.6, 1006.5, 1006.7, 1006.9, 
    1007, 1007.1, 1007.3, 1007.2, 1007.4, 1007.3, 1007.4, 1007.4, 1007.3, 
    1007.2, 1007.2, 1007.6, 1007.7, 1008.1, 1008.2, 1008.4, 1008.6, 1008.7, 
    1008.8, 1009, 1009.1, 1009.2, 1009.3, 1009.4, 1009.4, 1010, 1010.4, 
    1010.5, 1010.9, 1011.2, 1011.5, 1011.8, 1011.9, 1012, 1012, 1012.6, 
    1012.9, 1013.5, 1013.9, 1014.1, 1014.7, 1015, 1015.3, 1015.7, 1015.9, 
    1016.2, 1016.2, 1016.5, 1016.6, 1017, 1017.4, 1017.4, 1017.3, 1017.6, 
    1017.9, 1017.8, 1018, 1018.5, 1018.5, 1018.5, 1018.9, 1019.3, 1019.3, 
    1019.7, 1020, 1020.2, 1020.4, 1020.7, 1020.8, 1020.9, 1021.1, 1021.3, 
    1021.7, 1021.9, 1022.2, 1022.2, 1022.5, 1022.8, 1022.6, 1022.9, 1023, 
    1023, 1022.8, 1022.7, 1022.9, 1022.9, 1022.8, 1022.7, 1022.3, 1021.9, 
    1021.5, 1021.3, 1021.3, 1020.9, 1020.6, 1020.2, 1019.9, 1019.8, 1019.5, 
    1019, 1018.4, 1018, 1017.7, 1017.1, 1016.2, 1015.3, 1014.8, 1014, 1013.2, 
    1012.7, 1012.3, 1012, 1011.4, 1010.6, 1010.1, 1009.5, 1009.1, 1008.2, 
    1007.8, 1006.9, 1006.2, 1005.7, 1004.9, 1003.9, 1003.1, 1002.5, 1001.7, 
    1000.9, 1000, 1000, 999, 998.8, 999.4, 999.8, 1000.2, 1000.4, 1000.7, 
    1000.2, 1000.3, 1000.8, 1001.1, 1000.7, 1000.6, 1000.4, 1000.4, 1000.4, 
    1000.4, 1000.1, 999.7, 999.2, 998, 997.1, 996, 995.1, 993, 991.5, 989.9, 
    988.8, 987.9, 987, 985.2, 984, 982.1, 981, 979.5, 978.7, 977.7, 977.4, 
    976.7, 976.3, 976.1, 976.1, 976.6, 977.2, 977.7, 978.4, 978.6, 978.7, 
    979, 979.7, 980.8, 981.6, 982.5, 982.8, 983.5, 983.7, 984.3, 984.8, 
    985.2, 985.5, 985.7, 985.9, 986.3, 986.4, 986.5, 986.6, 986.6, 986.5, 
    986.5, 986.4, 986.1, 985.7, 985.7, 985.7, 985.7, 985.6, 985.5, 985.1, 
    984.8, 984.4, 984.2, 983.8, 983.5, 983, 982.7, 982.5, 982.1, 981.8, 
    981.6, 981.2, 980.8, 980.7, 980.6, 980.2, 980, 979.5, 979.3, 979.2, 
    979.3, 979.3, 979.2, 979.1, 979, 978.8, 978.8, 979, 979.2, 979.1, 979.4, 
    979.7, 980.1, 980.9, 981.7, 982.3, 983, 983.7, 984.5, 985.2, 986.3, 
    987.4, 988.4, 989.9, 991.1, 992.4, 993.3, 994.3, 995.4, 996.4, 997.6, 
    998.5, 999.3, 1000.2, 1000.7, 1001.4, 1002.4, 1003.2, 1004.1, 1004.8, 
    1005.4, 1006.2, 1007, 1007.8, 1008.3, 1009, 1009.7, 1010.4, 1011.1, 
    1011.9, 1012.3, 1012.8, 1013.4, 1013.9, 1014.4, 1014.8, 1015.1, 1015.6, 
    1016, 1016.5, 1016.9, 1017.3, 1017.8, 1018.3, 1018.5, 1018.8, 1019.2, 
    1019.2, 1019.4, 1019.5, 1019.6, 1020, 1020.3, 1020.2, 1020.3, 1020.2, 
    1020.4, 1020.4, 1020.3, 1020.1, 1020.3, 1019.9, 1019.4, 1019.5, 1019.1, 
    1018.7, 1018.3, 1018.1, 1017.3, 1016.7, 1016.1, 1015, 1014.2, 1012.8, 
    1011.6, 1010.9, 1010.1, 1009.1, 1008.1, 1007.3, 1006.4, 1005.3, 1004.1, 
    1003.1, 1002.5, 1001.6, 1000.8, 1000.5, 1000, 999.3, 998.7, 998.2, 997.6, 
    997.2, 996.7, 996.4, 995.8, 995.4, 995.1, 994.9, 994.4, 994.4, 994.3, 
    993.6, 993.3, 992.6, 991.7, 990.9, 990.7, 990.4, 990.4, 990.6, 991, 
    991.5, 992.4, 993.2, 993.4, 994.1, 994.3, 994.9, 995.3, 995.6, 996, 
    996.2, 996, 996.3, 996.6, 996.5, 996.4, 996.7, 996.9, 996.7, 996.8, 
    996.9, 996.8, 996.7, 996.1, 995.4, 995.4, 995.4, 995.1, 994.7, 994.5, 
    994.5, 994.1, 995.2, 995.9, 996.4, 996.8, 997.6, 997.9, 998.2, 999.1, 
    999.7, 999.9, 1000.1, 1000.5, 1001, 1001.8, 1002.1, 1002.9, 1003.4, 
    1003.9, 1004.5, 1004.7, 1005.1, 1005.5, 1005.7, 1005.9, 1006.1, 1006.3, 
    1006.4, 1006.5, 1006.2, 1006.3, 1006.1, 1005.9, 1005.8, 1005.5, 1005.4, 
    1005.4, 1005.4, 1005.2, 1005.2, 1005.4, 1005.5, 1005.8, 1005.6, 1005.6, 
    1005.9, 1005.9, 1006, 1006.1, 1006.2, 1006.8, 1007.1, 1007.3, 1007.6, 
    1007.7, 1008.2, 1008.3, 1008.5, 1008.8, 1008.9, 1009.2, 1009.5, 1009.7, 
    1009.9, 1009.9, 1010, 1010.2, 1010.5, 1010.5, 1010.7, 1010.7, 1010.5, 
    1010.2, 1010.2, 1010.1, 1010.2, 1010.2, 1010.3, 1010.2, 1009.9, 1009.6, 
    1009.2, 1008.9, 1008.7, 1008.5, 1008.2, 1008, 1007.7, 1007.3, 1006.9, 
    1006.4, 1005.9, 1005.3, 1004.9, 1004.2, 1003.7, 1003.3, 1002.9, 1002.6, 
    1002.6, 1002.9, 1003.3, 1003.5, 1003.8, 1004.6, 1004.9, 1005.4, 1005.2, 
    1005.3, 1004.9, 1004.9, 1004.8, 1005, 1005, 1005.2, 1005.4, 1005.2, 
    1005.2, 1005.1, 1005, 1005, 1004.5, 1004.3, 1004.6, 1005.3, 1005, 1005.1, 
    1005.4, 1005.4, 1005.6, 1005.8, 1005.9, 1005.8, 1005.7, 1005.7, 1005.8, 
    1005.9, 1005.9, 1006, 1006, 1006.1, 1006.2, 1006.1, 1006.1, 1005.9, 
    1005.7, 1005.8, 1005.6, 1005.7, 1005.6, 1005.4, 1005.4, 1005.5, 1005.3, 
    1005.4, 1005.6, 1005.7, 1005.9, 1006.5, 1007, 1007.5, 1008, 1008.4, 
    1008.7, 1009.2, 1009.3, 1009.5, 1009.6, 1009.7, 1009.7, 1009.9, 1010.3, 
    1010.6, 1010.8, 1011, 1011.1, 1011, 1010.8, 1011, 1010.9, 1010.8, 1010.9, 
    1011.2, 1010.8, 1011, 1011.2, 1011.4, 1011.6, 1011.7, 1011.9, 1012.2, 
    1012.3, 1012.3, 1012.5, 1012.7, 1013.1, 1013.5, 1014, 1014.3, 1014.6, 
    1014.9, 1015, 1015.2, 1015.4, 1015.6, 1015.9, 1016, 1016.4, 1016.9, 
    1017.3, 1017.8, 1017.9, 1017.9, 1017.9, 1018.1, 1018, 1017.8, 1017.6, 
    1017.5, 1017.2, 1016.6, 1016.1, 1015.1, 1014.5, 1013.3, 1012.1, 1011.4, 
    1010.9, 1010.4, 1010.3, 1010.4, 1011, 1011.8, 1013.1, 1013.2, 1014.3, 
    1014.6, 1014.8, 1014.3, 1013.9, 1013.2, 1012.2, 1010.9, 1009.8, 1008.6, 
    1007.2, 1006, 1004.6, 1003.5, 1002.4, 1001.3, 1000.4, 1000.5, 1000, 
    999.9, 1000.2, 1000.7, 1001, 1001.5, 1001.9, 1001.7, 1001.9, 1002.2, 
    1002.4, 1002.8, 1002.3, 1003.7, 1004.7, 1005.3, 1006.2, 1007.2, 1008.1, 
    1009.1, 1009.7, 1010.4, 1011.6, 1012.4, 1013.1, 1013.8, 1014.6, 1015.3, 
    1015.9, 1016.6, 1017.3, 1017.8, 1018.3, 1018.5, 1019.1, 1019.4, 1019.9, 
    1020.3, 1020.7, 1020.8, 1020.8, 1020.8, 1020.7, 1020.1, 1019.5, 1018.5, 
    1017.4, 1016.2, 1015.3, 1013.9, 1012.1, 1010.3, 1008.5, 1007.5, 1007, 
    1006.1, 1005.7, 1005.1, 1004.1, 1003.5, 1002.6, 1002, 1002.4, 1002.5, 
    1003, 1003, 1003.1, 1002.7, 1002.3, 1002.1, 1002.3, 1002.1, 1002.4, 
    1002.4, 1001.8, 1001.8, 1002, 1001.7, 1001.7, 1001.7, 1001.6, 1002, 
    1001.9, 1002, 1002.4, 1002.6, 1002.7, 1002.8, 1003, 1003.4, 1003.8, 
    1002.6, 1002.5, 1002.6, 1002.9, 1003, 1002.9, 1002.7, 1002.6, 1002.5, 
    1002.2, 1002.1, 1002.1, 1001.7, 1001.3, 1001.1, 1000.9, 1000.8, 1001, 
    1001, 1000.9, 1001.2, 1001.4, 1001.9, 1002.2, 1002.3, 1002.2, 1002.5, 
    1002.9, 1003.2, 1003.4, 1003.9, 1004.3, 1004.5, 1004.8, 1005.2, 1005.5, 
    1005.7, 1006, 1006.2, 1006.3, 1006.7, 1006.9, 1007.2, 1007.6, 1008.2, 
    1008.5, 1008.7, 1009, 1009.1, 1009.4, 1009.4, 1009.4, 1009, 1009.2, 
    1009.1, 1009, 1008.9, 1008.6, 1008.8, 1008.2, 1008.2, 1008, 1007.5, 
    1007.4, 1007.4, 1007, 1006.9, 1007, 1006.7, 1007, 1006.9, 1007, 1006.7, 
    1007.1, 1007.1, 1007.5, 1008, 1008.3, 1008.2, 1008.6, 1008.8, 1008.8, 
    1009.1, 1009.6, 1009.4, 1009.9, 1009.8, 1009.7, 1010.1, 1010.5, 1010.5, 
    1011.2, 1011, 1011.6, 1012.1, 1012, 1012.1, 1012.4, 1012.5, 1013.2, 
    1013.2, 1013.3, 1013.2, 1012.9, 1013, 1013.6, 1013.8, 1013.8, 1013.7, 
    1013.6, 1014, 1014.1, 1014.5, 1014.4, 1014.6, 1015.1, 1015.3, 1015.7, 
    1016.1, 1016.2, 1016.2, 1016.3, 1016.2, 1016.4, 1016.1, 1015.5, 1015.1, 
    1015, 1014.9, 1014.5, 1014.7, 1014.6, 1014.2, 1013.8, 1013.5, 1013, 1013, 
    1012.9, 1012.7, 1012.7, 1013.1, 1013.3, 1013.7, 1013.6, 1013.8, 1014, 
    1013.9, 1014.1, 1014.3, 1014.4, 1014.5, 1014.6, 1014.8, 1015.1, 1015.4, 
    1015.4, 1015.5, 1016, 1016, 1016.1, 1016.4, 1016.5, 1016.7, 1017.1, 
    1017.7, 1017.7, 1017.7, 1018.1, 1017.8, 1017.7, 1017.8, 1018.1, 1018.1, 
    1017.9, 1017.8, 1017.8, 1017.7, 1018.2, 1018.2, 1018.3, 1018.2, 1018.2, 
    1018.2, 1018.2, 1018.2, 1018.4, 1018.4, 1018.6, 1018.8, 1019.2, 1019.4, 
    1019.5, 1019.7, 1019.9, 1020, 1020.2, 1020.5, 1020.5, 1020.7, 1020.8, 
    1021.1, 1021.3, 1021.8, 1021.8, 1021.5, 1021.7, 1021.5, 1021.2, 1021.3, 
    1021.2, 1021.4, 1021.7, 1021.8, 1022.2, 1022.3, 1022.5, 1022.7, 1022.7, 
    1022.8, 1022.8, 1023.1, 1023.6, 1023.5, 1023.7, 1023.8, 1023.7, 1024.1, 
    1024.3, 1024.2, 1024.2, 1024.3, 1024.3, 1024.4, 1024.8, 1025, 1025.5, 
    1025.9, 1026.3, 1026.5, 1026.3, 1026.3, 1026.5, 1026.6, 1027, 1026.9, 
    1026.8, 1026.7, 1026.1, 1026.3, 1026, 1025.6, 1025.3, 1024.9, 1024.6, 
    1024.1, 1023.3, 1022.5, 1022.1, 1021.5, 1020.9, 1020.3, 1019.7, 1019.2, 
    1018.4, 1017.7, 1017.1, 1016.1, 1015.7, 1015.1, 1014.7, 1013.8, 1012.9, 
    1012.5, 1012.1, 1011.5, 1011, 1010, 1009.2, 1008.6, 1008.1, 1007.2, 
    1006.8, 1006.3, 1005.7, 1005.3, 1004.4, 1003.6, 1002.4, 1001.3, 1000, 
    998.6, 997.1, 995.5, 994, 991.9, 990, 988.6, 987, 985.1, 983.6, 981.8, 
    979.6, 977.3, 975.1, 972.8, 970.9, 968.9, 967.5, 966.3, 965.8, 965.7, 
    966.2, 966.7, 967.3, 967.4, 967.7, 968.7, 969.6, 970.9, 972.5, 974.9, 
    976.6, 978.4, 980.5, 982.1, 983.6, 984.8, 985.8, 986.7, 987.3, 987.5, 
    988, 988.5, 988.8, 989.1, 991, 991.2, 989.8, 990, 989.9, 989.9, 989.9, 
    989.6, 989.7, 989.6, 989.4, 989.1, 989, 987.9, 987.5, 987.3, 987, 986.8, 
    986.4, 986.2, 986.2, 986.2, 986.2, 986.1, 985.9, 986, 986.2, 986.4, 
    986.8, 987.3, 987.2, 987.4, 987.9, 988.5, 989, 989.8, 990.4, 990.8, 991, 
    990.8, 990.8, 991, 991.2, 991.6, 992, 992, 992.3, 992.3, 992.3, 992.4, 
    992.5, 992.9, 992.9, 992.8, 992.6, 992.7, 992.8, 993.1, 993.3, 993.8, 
    993.9, 993.5, 992.9, 992.6, 992.2, 991.9, 992.6, 991.2, 990.8, 989.8, 
    989.1, 988.7, 987.9, 987.2, 986.3, 985.4, 984.4, 983.9, 983.8, 983.4, 
    982.8, 982.2, 982.1, 982.4, 982.6, 982.7, 982.6, 982.9, 983.2, 983.4, 
    983.5, 983.8, 984.2, 984.8, 985.6, 986.2, 986.6, 987, 987.2, 987.2, 
    987.6, 987.9, 988, 987.9, 988, 988.1, 988.2, 988.5, 988.5, 988.5, 988.2, 
    988.2, 988, 987.7, 987.9, 987.9, 987.7, 987.3, 987, 987, 986.8, 986.5, 
    986.4, 986.1, 985.8, 985.7, 985.4, 985.7, 985.5, 985.6, 985.7, 985.8, 
    985.7, 985.7, 985.8, 986, 986.2, 986.4, 986.5, 986.5, 986.6, 987.2, 
    987.6, 988, 988.3, 988.3, 988.7, 989.1, 989.6, 990, 990.4, 990.6, 991, 
    991.4, 991.7, 992, 992.4, 992.6, 992.9, 993.2, 993.6, 993.8, 994.2, 
    994.6, 995, 995.8, 996.5, 997.2, 997.7, 998.5, 999.2, 999.9, 1000.7, 
    1001.5, 1002, 1002.6, 1003.5, 1004.6, 1005.5, 1006.2, 1007, 1007.3, 
    1007.8, 1008, 1008.6, 1008.7, 1008.9, 1009.1, 1009.3, 1010, 1010.2, 
    1010.2, 1010.7, 1011.3, 1011.6, 1011.9, 1012.6, 1013.4, 1013.7, 1014.6, 
    1015, 1015.8, 1016.3, 1016.9, 1017.1, 1017.3, 1017.8, 1017.7, 1017.3, 
    1017.3, 1016.4, 1015.2, 1013.9, 1012.6, 1010.6, 1008.6, 1006.8, 1004.4, 
    1002.1, 999.5, 996.7, 994.2, 991.6, 988.7, 986.8, 985.2, 984.4, 983.8, 
    983.6, 983.6, 983.3, 983, 982.8, 982.7, 982.4, 982.2, 981.8, 981.5, 
    981.3, 981.2, 981, 981.3, 981.5, 981.6, 981.5, 980.7, 980.3, 979.8, 
    980.7, 980.9, 981.7, 983.1, 983.7, 984.4, 984.4, 984.7, 984.6, 984.2, 
    984.1, 983.7, 983.5, 983.8, 983.3, 983.2, 982.8, 982.3, 981.5, 981, 
    980.1, 980.3, 980.1, 980.3, 980.7, 981.2, 982, 982.3, 982.4, 982.6, 
    982.8, 983, 983.3, 983.9, 984.1, 984.8, 985, 985.4, 986.1, 986.5, 986.9, 
    987.7, 988, 988.5, 988.9, 989.2, 989.3, 989.2, 989.5, 989.8, 990.1, 
    990.4, 990.6, 990.9, 991, 990.8, 990.9, 991, 991.1, 991.4, 991.6, 991.6, 
    991.8, 992.2, 992.8, 993.1, 992.7, 992.8, 993.1, 993.1, 993, 992.8, 993, 
    993.2, 993.4, 993.2, 993.2, 993.3, 993.3, 993.1, 993.2, 993.6, 993.6, 
    993.9, 993.8, 994.1, 994.5, 994.7, 994.7, 994.6, 994.5, 994.4, 994.1, 
    993.5, 993.2, 993, 992.9, 992.7, 992.6, 992.4, 992.2, 992.1, 991.8, 
    991.5, 991.3, 991.1, 991.1, 991.1, 990.9, 990.7, 990.9, 990.9, 990.7, 
    990.6, 990.5, 990.3, 990.3, 990.1, 990, 989.9, 989.7, 989.8, 989.8, 
    989.6, 989.2, 988.9, 988.5, 988.5, 988.2, 987.8, 987.9, 987.8, 987.6, 
    987.7, 987.7, 987.6, 987.8, 988.2, 988.2, 988, 988.2, 988.6, 988.8, 
    989.3, 989.6, 990, 990.4, 990.9, 991, 991.6, 992.1, 992.5, 992.8, 993.6, 
    994.3, 994.7, 995.4, 995.8, 996.5, 997.1, 997.6, 998.1, 998.2, 998.6, 
    998.9, 999.1, 999.6, 1000, 1000.3, 1000.8, 1001.4, 1001.8, 1002.2, 
    1002.3, 1002.5, 1002.8, 1003.1, 1003.4, 1003.3, 1003.5, 1003.9, 1004.2, 
    1004.3, 1004.7, 1004.5, 1004.4, 1004.3, 1003.7, 1004, 1003.8, 1003.7, 
    1003.8, 1003.2, 1002.8, 1002.7, 1002.6, 1002.1, 1001, 1000, 998.7, 998.3, 
    997.6, 996.9, 996.8, 996.8, 996.6, 996.4, 996.4, 995.9, 995.3, 995.1, 
    995.1, 995, 994.8, 994.7, 995, 995.6, 995.9, 996.2, 996.6, 997.4, 998, 
    998.7, 999.3, 999.9, 1000.4, 1001, 1001.5, 1002.4, 1003.1, 1004.1, 
    1005.2, 1006, 1006.8, 1007.6, 1008.2, 1009, 1009.6, 1010.1, 1011, 1011.3, 
    1011.7, 1012.6, 1013.1, 1013.6, 1013.7, 1013.9, 1014.1, 1013.8, 1013.7, 
    1013.6, 1013.7, 1013.6, 1013.5, 1013.6, 1014, 1013.3, 1012.1, 1011.9, 
    1012.3, 1011.8, 1011, 1010.8, 1010, 1009.7, 1009, 1008.4, 1008.1, 1007.5, 
    1006.9, 1006.7, 1006.3, 1005.4, 1005, 1004.6, 1004, 1003.8, 1003.7, 
    1003.5, 1003.6, 1003.1, 1002.9, 1002.8, 1002.4, 1002, 1001.8, 1001.6, 
    1001.2, 1000.6, 1000.7, 1000.1, 1000.1, 999.6, 998.9, 998.6, 998.7, 
    998.3, 997.9, 997.1, 996.8, 996.7, 996.7, 996.7, 996.4, 996.2, 995.8, 
    996.1, 995.7, 995.7, 995.4, 995.7, 995.1, 994.7, 995, 995.4, 995.8, 
    995.9, 995.8, 996.1, 996.1, 996.1, 996.1, 995.9, 995.9, 995.9, 996.3, 
    996.5, 996.8, 996.8, 996.6, 996.6, 996.4, 996, 995.9, 995.5, 995.1, 
    994.8, 994, 994.3, 993.2, 992.9, 992.4, 991.9, 991.4, 991, 990.8, 990.9, 
    990.9, 991.2, 991.6, 992.1, 992.3, 993, 993.3, 993.8, 994.2, 994.4, 995, 
    995.7, 996.4, 997.1, 997.9, 998.4, 998.7, 999.3, 999.8, 1001.2, 1001.7, 
    1002.1, 1002.4, 1002.7, 1003.4, 1003.8, 1003.9, 1004, 1004.1, 1004.1, 
    1003.9, 1003.9, 1004, 1003.9, 1003.5, 1003.1, 1003.4, 1003, 1002.6, 
    1002.3, 1002, 1001.7, 1000.8, 1000.4, 999.9, 999.3, 999, 998.7, 998.8, 
    998.6, 998.4, 998.2, 998.3, 998.8, 998.8, 998.7, 999.1, 999.2, 999.2, 
    999.4, 999.2, 999, 999, 998.8, 998.3, 997.6, 996.6, 995.8, 995.4, 994.6, 
    993.5, 992.8, 991.7, 991.2, 990.5, 989.6, 989.2, 988.6, 987.5, 986.9, 
    986.3, 985.7, 985.2, 984.9, 985, 984.4, 984, 983.5, 983.1, 982.8, 982.4, 
    982, 981.6, 981, 980.5, 979.7, 979.4, 979, 978.8, 978.3, 977.7, 976.8, 
    975.1, 973.7, 972.4, 971, 968.9, 966.9, 969.6, 967.7, 966.5, 965, 963.3, 
    961.8, 960.6, 959.4, 958.2, 956.9, 955.8, 954.8, 953.6, 952.6, 952, 
    951.8, 951.6, 951.6, 951.9, 952.4, 952.9, 952.9, 952.8, 952.7, 955.1, 
    955, 955, 954.9, 955.1, 955.2, 955.4, 955.7, 956.1, 956.3, 956.7, 957, 
    958.9, 959.4, 960, 960.6, 961.5, 962.1, 962.8, 963.7, 964.6, 965.5, 
    966.4, 967.4, 968.7, 969.4, 970.2, 971.2, 971.9, 972.8, 973.7, 974.4, 
    975.2, 975.8, 976.3, 977, 977.6, 978.4, 979, 980.8, 981.7, 982.3, 983.3, 
    984.4, 985.4, 986.2, 986.9, 986.4, 987.1, 988.1, 989.1, 990.2, 991, 
    991.6, 992.4, 993.3, 994.2, 994.8, 995.6, 995.2, 996, 996.7, 997.7, 
    998.7, 999.6, 1000.3, 1001, 1001.7, 1002.1, 1002.5, 1002.4, 1002.8, 1003, 
    1003.5, 1003.8, 1003.5, 1003.6, 1003.4, 1003.1, 1003, 1002.5, 1002.1, 
    1001.5, 1001.9, 1000.8, 1000.2, 999.5, 998.3, 996.3, 994.4, 992.9, 991.1, 
    989, 987.3, 986.1, 986.2, 985.9, 986.4, 987.6, 989.2, 990.8, 992.6, 
    994.5, 996.4, 998.6, 999.3, 1001.7, 1002.3, 1003.2, 1004.6, 1005.2, 
    1005.2, 1005, 1004.6, 1003.6, 1002.7, 1001.9, 1001.4, 1000.7, 1000.6, 
    1000.3, 1000, 1000, 1000.5, 1001.2, 1002.3, 1003.7, 1005.8, 1008, 1009.5, 
    1011.3, 1014.5, 1015.7, 1016.6, 1018.3, 1019, 1019.2, 1019.4, 1020, 
    1019.8, 1019.7, 1018.6, 1018, 1016.8, 1015.3, 1013.5, 1011.9, 1009.9, 
    1008.2, 1006.3, 1004.4, 1002, 1000.5, 998.6, 997.6, 996.8, 996.1, 995.8, 
    995.4, 994.9, 994.2, 993.2, 991.1, 988.4, 985.6, 981.9, 979.4, 977.7, 
    980.7, 981.6, 981.4, 981.8, 982.7, 984.6, 986.7, 989.2, 992.3, 996.8, 
    1000, 1002.2, 1004.9, 1007.1, 1009.4, 1011.4, _, 1014.6, _, 1015.5, 
    1016.4, 1016.1, 1015.8, 1014.4, 1015, 1015, 1014.6, 1014.5, 1014.3, 
    1014.1, 1014, 1013.6, 1013.6, 1013.8, _, 1013.5, 1014.2, 1014.8, 1015.2, 
    1015.8, 1016.5, 1016.7, 1017, 1016.8, 1016.7, 1016.9, 1016.9, 1017.2, 
    1017.5, 1017.9, 1018.2, 1018.4, 1018.9, 1020, 1019, 1019, 1019, 1019, 
    1019.2, 1019.2, 1019.2, 1019.2, 1019.5, 1019.4, 1019.2, 1018.8, 1018.7, 
    1018.6, 1018.4, 1018, 1017.8, 1017.9, 1018.2, 1018.6, 1018.7, 1019.1, 
    1019.3, 1019.4, 1019.6, 1019.6, 1019.8, 1021.8, 1021.9, 1020.4, 1020.8, 
    1021, 1021.7, 1022.2, 1022.5, 1022.4, 1022.7, 1022.9, 1022.9, 1023.1, 
    1023.6, 1023.6, 1023.3, 1023.5, 1023.7, 1023.9, 1023.8, 1023.9, 1025.2, 
    1024.1, 1024.4, 1023.9, 1024.3, 1024.5, 1024.7, 1024.9, 1025.7, 1025.9, 
    1025.7, 1025.5, 1025.4, 1025.4, 1025, 1024.8, 1024.6, 1024.7, 1024.5, 
    1024.2, 1024.1, 1023.9, 1024.2, 1024, 1022.9, 1022.8, 1022.4, 1021.9, 
    1021.7, 1021.4, 1021.1, 1021, 1020.7, 1020.6, 1019.9, 1019.4, 1018.8, 
    1018, 1017.7, 1016.9, 1016.2, 1015.4, 1014.8, 1014.4, 1015.3, 1012.7, 
    1014.4, 1011.3, 1011, 1010.5, 1009.7, 1012, 1011.6, 1008.7, 1008.6, 
    1011.1, 1010.9, 1010.8, 1008.6, 1008.7, 1008.8, 1009.1, 1009.2, 1009.3, 
    1009.3, 1011.7, 1010, 1010.1, 1012.1, 1010.8, 1011.2, 1011.6, 1013.4, 
    1012.1, 1012.1, 1013.9, 1012.8, 1013.2, 1015.2, 1013.9, 1015.7, 1014.7, 
    1015, 1015.2, 1015.4, 1015.7, 1016.1, 1016.4, 1016.5, 1016.2, 1017.4, 
    1016.7, 1017.1, 1017.1, 1017.9, 1017.1, 1017.2, 1017.2, 1017.2, 1017.2, 
    1017.3, 1017, 1016.8, 1016.8, 1016.8, 1016.6, 1016.6, 1016.6, 1016.6, 
    1016.4, 1016.2, 1016.1, 1015.9, 1015.7, 1015.7, 1015.6, 1015.5, 1015.4, 
    1015.1, 1014.4, 1014.5, 1014.2, 1014.2, 1014.1, 1014.4, 1013.9, 1013.5, 
    1012.8, 1012.3, 1012, 1011.7, 1011.1, 1010, 1009.2, 1008.2, 1007.8, 
    1007.1, 1006.4, 1005.8, 1005.3, 1006.4, 1004.9, 1004.3, 1003.4, 1002.4, 
    1001.6, 1001, 1000.9, 1000.9, 1000.5, 1000.2, 999.6, 999.2, 999.4, 999.6, 
    999.9, 1000.1, 1000.2, 1000.8, 1001.1, 1001.4, 1001.4, 1001.9, 1001.5, 
    1001.8, 1001.2, 1000.4, 1000.1, 999.5, 999, 998.3, 997.9, 997.5, 997.1, 
    996.6, 996.2, 994.5, 994.1, 993.2, 992.2, 991.5, 990.9, 990.7, 990.3, 
    989.9, 989.5, 989.3, 989.2, 989.1, 989, 988.9, 988.9, 989.9, 988.8, 989, 
    989.2, 989.3, 989.6, 989.8, 990, 990.2, 990.5, 990.7, 991.4, 992, 992.5, 
    993.1, 993.6, 994.3, 994.9, 995.4, 995.8, 996, 996.2, 996.5, 996.5, 
    996.5, 996.8, 997.1, 997.4, 998.4, 998.9, 999.1, 999, 998.9, 999, 998.9, 
    998.5, 998.3, 1000.4, 1000.1, 1000.6, 1000.9, 1000.8, 1000.8, 1000.4, 
    1000, 999.7, 999, 998.1, 998.1, 999, 998.3, 998, 997.5, 997, 996.8, 
    996.3, 995.9, 994.9, 994.6, 994.3, 994.2, 993.6, 993.1, 992.1, 992, 
    992.4, 991.7, 991.9, 992.5, 991.4, 991.3, 993.6, 993.8, 993.3, 992.9, 
    994.4, 994.3, 995.3, 995, 995.6, 995.8, 997, 997.5, 997.6, 998.4, 998.9, 
    999.1, 999.5, 1000, 1000.5, 1000.8, 1001.4, 1002.3, 1001.8, 1002, 1002, 
    1002.3, 1002.6, 1002.9, 1003, 1002.7, 1002.9, 1002.8, 1002.6, 1002.2, 
    1002.1, 1002.3, 1002.2, 1001.7, 1001.3, 1001.3, 1001.4, 1001.9, 1001.7, 
    1000.9, 1001.3, 1001.5, 1001.7, 1002.1, 1002.2, 1002.2, 1002.8, 1002.7, 
    1003.5, 1004.1, 1004.9, 1005.2, 1005.9, 1006.6, 1006.9, 1007.8, 1008.6, 
    1009.3, 1010.3, 1010.9, 1011.8, 1012.5, 1013.2, 1013.5, 1014.7, 1015.2, 
    1015.8, 1016.2, 1017, 1017, 1017.6, 1018.5, 1018.7, 1019.3, 1019.6, 
    1019.9, 1019.9, 1020, 1020.2, 1020.6, 1021, 1021.3, 1021.7, 1021.7, 1022, 
    1022.4, 1022.7, 1023.1, 1023.4, 1023.7, 1024.2, 1024.4, 1024.3, 1024.4, 
    1024.5, 1024.5, 1024.8, 1025, 1025.4, 1026, 1026.2, 1026.3, 1026.4, 
    1026.2, 1026.5, 1026.5, 1026.9, 1027, 1027.2, 1027, 1027.7, 1026.8, 
    1026.6, 1027.6, 1025.9, 1025.6, 1025.8, 1025.9, 1026, 1025.4, 1025.1, 
    1024.8, 1024.6, 1024, 1023.4, 1023.2, 1022.6, 1022.5, 1021.9, 1020.9, 
    1020.7, 1020.5, 1019.6, 1019, 1017.7, 1018.1, 1015.9, 1015.1, 1014, 
    1013.1, 1012.3, 1011.5, 1012.4, 1009.9, 1009.4, 1008.6, 1007.7, 1006.8, 
    1006.1, 1005.4, 1004.2, 1003.5, 1002.6, 1002, 1001.7, 1001.1, 1000.4, 
    999.7, 999, 998.4, 997.9, 998.9, 996.8, 996.4, 997.1, 995.7, 995.3, 
    994.8, 994.4, 993.5, 992.5, 991.9, 991, 990.4, 989.6, 989.3, 988.9, 
    988.5, 988.2, 988, 987.8, 987.5, 988.1, 987.9, 988, 988.6, 988.3, 988.4, 
    988.9, 989.5, 990.1, 990.5, 991.1, 991.6, 992.2, 992.8, 993.3, 993.8, 
    994.3, 994.8, 995.4, 995.7, 996, 996.2, 996.3, 996.6, 996.5, 997.3, 
    997.6, 996.8, 997.1, 997.1, 997, 997, 998, 996.9, 996.9, 996.8, 996.9, 
    997, 997.2, 997.3, 997.3, 997.1, 996.9, 996.7, 996.6, 996.5, 996.4, 
    996.4, 995.9, 995.4, 995, 994.6, 994.1, 993.5, 993.4, 992.8, 992.1, 992, 
    991.7, 991.6, 991.6, 991.7, 991.6, 991.8, 992, 992.1, 992.4, 992.7, 993, 
    993.4, 994.1, 994.6, 994.9, 995.4, 996.8, 997.2, 997.7, 997.8, 998.3, 
    998.6, 999.1, 999.5, 1000, 1000.2, 1000.9, 1001.1, 1001.4, 1001.4, 
    1001.4, 1001.6, 1001.7, 1002.1, 1002.3, 1002.3, 1002.4, 1002.6, 1002.4, 
    1002.6, 1002.5, 1002.5, 1002.5, 1002.4, 1002.6, 1002.5, 1002.6, 1002.6, 
    1002.3, 1002.4, 1002.5, 1002.2, 1002.1, 1001.9, 1001.7, 1001.7, 1001.7, 
    1001.4, 1001.1, 1000.7, 1000.6, 1000.3, 1000, 999.6, 999.4, 999.2, 999, 
    998.8, 998.3, 998.2, 997.8, 997.3, 997.2, 996.3, 995.8, 995.2, 994.9, 
    994.8, 994.7, 994.8, 994.9, 996.7, 997.1, 997.8, 998.5, 999.3, 999.8, 
    1000.3, 1000.8, 1001.2, 1001.6, 1001.9, 1002.3, 1002.5, 1002.7, 1003.1, 
    1003.2, 1003.4, 1003.6, 1003.6, 1003.7, 1003.7, 1003.6, 1003.8, 1003.8, 
    1003.6, 1003.4, 1003.5, 1003.4, 1003, 1002.8, 1002.7, 1000, 999.5, 999.1, 
    998.7, 998, 997.4, 996.5, 995.7, 994.7, 993.6, 994, 993.8, 994.2, 994.7, 
    995.6, 996.3, 997.2, 998.6, 1000.1, 1001.2, 1002.6, 1004.2, 1005.4, 
    1006.5, 1007.6, 1008.3, 1008.6, 1009.1, 1009.6, 1010.1, 1010.6, 1010.7, 
    1010.3, 1009.4, 1008.2, 1007.6, 1006.5, 1005.3, 1003.6, 1002.4, 1001.5, 
    1000.8, 1000.1, 999, 998.1, 997.1, 996.1, 995.4, 994.7, 994.1, 993.5, 
    993.1, 993.1, 993.1, 993.5, 993.9, 994.3, 995, 995.9, 996.8, 997.6, 
    998.3, 999.1, 999.6, 1000.5, 1001.3, 1002, 1002.8, 1003.5, 1004, 1004.8, 
    1005.6, 1006.2, 1006.9, 1007.2, 1007.6, 1007.8, 1008, 1008.1, 1008.2, 
    1008.2, 1007.9, 1007.6, 1007.4, 1007.2, 1007.1, 1006.7, 1006.5, 1006.6, 
    1006.8, 1007.1, 1007.5, 1007.7, 1008.3, 1008.6, 1009, 1009.4, 1010, 
    1010.7, 1011.1, 1011.4, 1011.9, 1012.4, 1012.5, 1013.1, 1013, 1012.9, 
    1013.1, 1013.2, 1013.2, 1013, 1013.2, 1013, 1012.7, 1012.4, 1011.9, 
    1011.4, 1010.1, 1008.4, 1007.8, 1006.7, 1006, 1005.4, 1004.9, 1004.4, 
    1003.9, 1003.3, 1003.2, 1003.5, 1003.3, 1003.1, 1003.4, 1003.3, 1003.2, 
    1003.1, 1003.1, 1003.3, 1003.4, 1003.9, 1003.8, 1003.7, 1003.4, 1003.1, 
    1003.1, 1002.7, 1002.7, 1002.3, 1002.4, 1002.5, 1001.9, 1002, 1002.2, 
    1003.3, 1003.7, 1004.3, 1004.5, 1004.8, 1007.1, 1008.3, 1008.9, 1009.8, 
    1010.2, 1011, 1012, 1012.9, 1013.9, 1015.1, 1018.2, 1019.3, 1020.4, 1021, 
    1022.1, 1024.3, 1025, 1026.1, 1026.3, 1027, 1027.4, 1027.5, 1027.4, 
    1026.9, 1026.7, 1026.1, 1025.8, 1025.2, 1024.9, 1024.6, 1024.3, 1024.4, 
    1023.9, 1024.2, 1023.9, 1023.4, 1022.7, 1022, 1020.1, 1019.7, 1019.1, 
    1018.9, 1018.2, 1018.6, 1018.7, 1019, 1019.5, 1020.1, 1020.1, 1019.9, 
    1019.7, 1019.2, 1019.6, 1019.7, 1019.6, 1019.6, 1019.8, 1019.5, 1019.5, 
    1019.5, 1019.3, 1018.6, 1018.4, 1018.3, 1017.9, 1018, 1017.7, 1017.3, 
    1016.7, 1017, 1016.9, 1016.8, 1017.1, 1017.1, 1017, 1016.7, 1016.4, 
    1016.6, 1016.6, 1017, 1016.9, 1017.1, 1017.1, 1017.2, 1017.2, 1017.3, 
    1017.3, 1017.3, 1017.4, 1017.6, 1017.8, 1018.2, 1018.2, 1018, 1018.3, 
    1018.5, 1018.8, 1018.8, 1018.9, 1019, 1018.7, 1018.7, 1018.6, 1018.7, 
    1018.6, 1018.3, 1018.3, 1018.1, 1018.1, 1018.1, 1018, 1018.1, 1018.1, 
    1018.1, 1018, 1018.1, 1018.1, 1018.3, 1018.5, 1018.8, 1018.9, 1019, 1019, 
    1019, 1018.9, 1018.9, 1018.9, 1019.2, 1019.3, 1019.4, 1018.8, 1019, 1019, 
    1019, 1018.9, 1018.8, 1018.8, 1018.8, 1018.7, 1018.6, 1018.4, 1018.5, 
    1018.5, 1018.5, 1018.4, 1018.5, 1018.5, 1018.3, 1018.2, 1018, 1018, 1018, 
    1017.9, 1017.9, 1017.7, 1017.5, 1017.3, 1017.2, 1017, 1016.7, 1016.4, 
    1016.3, 1016, 1015.3, 1012.2, 1012.5, 1012.6, 1012.5, 1012.5, 1012.7, 
    1012.9, 1013, 1013.3, 1013.3, 1013.3, 1013.5, 1013.7, 1013.9, 1014, 
    1014.4, 1014.4, 1014.5, 1014.8, 1015, 1015.2, 1015.6, 1016, 1016.3, 
    1016.7, 1016.9, 1017, 1017.2, 1017.3, 1017.1, 1016.9, 1017, 1016.9, 
    1016.8, 1016.4, 1016.2, 1016.1, 1016.4, 1016.4, 1016.4, 1016.4, 1016.5, 
    1016.5, 1016.6, 1016.7, 1016.3, 1016.3, 1016.4, 1016.5, 1016.1, 1016.1, 
    1016.1, 1016.2, 1016.2, 1016.2, 1016.1, 1016, 1016, 1015.5, 1015.3, 
    1015.3, 1015.4, 1015.2, 1015.2, 1014.8, 1014.7, 1014.6, 1014.5, 1014.5, 
    1014.3, 1014.4, 1014.4, 1014.2, 1014.2, 1014.4, 1014.6, 1014.7, 1014.7, 
    1014.8, 1015.1, 1015.1, 1015.4, 1015.5, 1015.9, 1016, 1016, 1016.3, 
    1016.5, 1016.6, 1016.9, 1017.3, 1017.5, 1017.3, 1017.6, 1017.9, 1018.2, 
    1018.6, 1018.9, 1019, 1019, 1019.1, 1019.1, 1019.3, 1019.6, 1019.7, 
    1019.7, 1019.6, 1019.4, 1019.4, 1019.3, 1019.2, 1019, 1019.2, 1019, 1019, 
    1018.7, 1018.5, 1018.3, 1018.1, 1018, 1017.9, 1017, 1016.6, 1016.4, 
    1016.2, 1016.1, 1015.9, 1015.6, 1015.3, 1015.1, 1014.7, 1014.4, 1014.1, 
    1013.8, 1013.7, 1013.3, 1013.2, 1013, 1012.8, 1012.7, 1012.4, 1012.1, 
    1011.5, 1011.1, 1010.7, 1010.3, 1010, 1009.7, 1009.4, 1009, 1008.7, 
    1008.4, 1007.4, 1007.1, 1006.8, 1006.8, 1006.6, 1006.5, 1006.4, 1006.4, 
    1006.4, 1006.3, 1006.2, 1006.2, 1006.1, 1005.7, 1005.5, 1005.5, 1005.8, 
    1005.9, 1006, 1005.9, 1006.1, 1006, 1006, 1006.1, 1006.3, 1006.5, 1006.7, 
    1007.1, 1007.3, 1007.6, 1007.8, 1008, 1008.1, 1008.3, 1008.2, 1008.3, 
    1008.4, 1008.6, 1008.8, 1009, 1009.2, 1009.2, 1009.2, 1009.5, 1009.7, 
    1009.8, 1009.8, 1009.9, 1010.1, 1010.2, 1010.6, 1010.9, 1011, 1011.1, 
    1011.3, 1011.6, 1011.8, 1012, 1012.1, 1012.4, 1012.8, 1014.1, 1014.1, 
    1014.5, 1014.8, 1015.2, 1015.3, 1015.5, 1015.6, 1016, 1016.4, 1016.6, 
    1017.1, 1017.4, 1017.5, 1017.8, 1017.9, 1018.1, 1018.2, 1018.1, 1018.2, 
    1018.2, 1018.3, 1018.4, 1018.4, 1018.4, 1018.2, 1017.6, 1017.4, 1017.2, 
    1017.1, 1017.2, 1017.2, 1017.2, 1017.2, 1017, 1016.9, 1016.8, 1016.6, 
    1016.3, 1016.2, 1016.1, 1015.7, 1015.5, 1015.4, 1015.2, 1014.9, 1014.5, 
    1014.3, 1014.3, 1014.2, 1014.1, 1013.7, 1013.5, 1013.2, 1012.7, 1012.3, 
    1012.2, 1011.9, 1011.5, 1011.4, 1011, 1010.8, 1010.7, 1010.8, 1010.7, 
    1010.7, 1010.2, 1010.1, 1010.3, 1010.5, 1010.8, 1011.1, 1011.2, 1011.5, 
    1011.7, 1012.2, 1012.5, 1012.9, 1013.2, 1013.5, 1013.8, 1014.1, 1014.4, 
    1014.6, 1014.8, 1014.8, 1015, 1015.1, 1015.3, 1015.6, 1015.8, 1016, 
    1016.3, 1016.3, 1016.3, 1016.2, 1016.1, 1016.3, 1016.3, 1016.3, 1016.5, 
    1016.4, 1016.5, 1016.4, 1016.1, 1015.9, 1015.7, 1015.6, 1015.5, 1015.4, 
    1015.2, 1015.1, 1015, 1014.8, 1014.7, 1014.3, 1014.1, 1014, 1013.8, 
    1013.8, 1013.6, 1013.4, 1013.4, 1013.3, 1013.5, 1013.6, 1013.4, 1013.4, 
    1013.4, 1013.3, 1013.3, 1013.2, 1013.5, 1013.6, 1013.6, 1013.5, 1013.1, 
    1013.1, 1012.7, 1012, 1011.8, 1011.8, 1011.7, 1011.3, 1010.9, 1010.6, 
    1010.3, 1009.8, 1009.2, 1009.2, 1009, 1008.9, 1008.6, 1008.5, 1008.3, 
    1007.9, 1007.3, 1007.1, 1006.4, 1006.1, 1005.7, 1005.3, 1005, 1004.7, 
    1004.4, 1004.2, 1003.8, 1003.5, 1003.1, 1002.7, 1002.2, 1001.7, 1001, 
    1000.6, 1000, 999.5, 999.2, 998.1, 997.5, 997.3, 997.1, 997, 996.6, 
    996.3, 996.3, 996.3, 996.4, 996.5, 996.8, 997, 997, 997.2, 997.3, 997.2, 
    997.3, 997.5, 997.6, 998, 998.6, 998.7, 999, 999.4, 999.2, 999.5, 999.5, 
    999.8, 999.8, 1000.2, 1000.6, 1000.9, 1001.2, 1001.6, 1001.9, 1002.2, 
    1002.5, 1002.8, 1003, 1004.8, 1005.2, 1005.5, 1006, 1007, 1007.3, 1009.3, 
    1009.4, 1009.5, 1009.7, 1010, 1010.2, 1010.3, 1010.3, 1010.9, 1011.1, 
    1011.3, 1011.3, 1011.4, 1011.8, 1012.1, 1012.4, 1012.7, 1012.9, 1013, 
    1013.5, 1013.7, 1013.8, 1014.1, 1014.2, 1014.2, 1014.7, 1015.3, 1015.7, 
    1015.8, 1016, 1016.2, 1016.4, 1016.7, 1017.3, 1017.5, 1018.3, 1018.5, 
    1019, 1019.2, 1019.4, 1019.7, 1020, 1020, 1020.2, 1020.2, 1020.6, 1020.9, 
    1021.2, 1021.4, 1021.5, 1022, 1022, 1021.9, 1021.9, 1022, 1022, 1022, 
    1022, 1021.9, 1022, 1021.9, 1021.7, 1021.5, 1021.2, 1020.9, 1020.7, 
    1020.5, 1020.3, 1019.9, 1019.8, 1019.8, 1019.6, 1019.4, 1019.2, 1018.8, 
    1018.5, 1018.2, 1018, 1017.8, 1017.7, 1017.5, 1017.3, 1017, 1016.8, 
    1016.6, 1016.4, 1016.2, 1015.9, 1015.8, 1015.6, 1015.3, 1015.3, 1015.1, 
    1014.8, 1014.6, 1014.5, 1014.2, 1014.1, 1013.7, 1013.4, 1013, 1013.1, 
    1013.4, 1013.5, 1013.6, 1013.7, 1013.6, 1013.4, 1013.3, 1013.1, 1013, 
    1013, 1012.8, 1012.8, 1012.6, 1012.5, 1012.6, 1012.6, 1012.4, 1012.1, 
    1011.9, 1011.8, 1011.5, 1011.3, 1011.3, 1011.3, 1011.3, 1011.2, 1011.3, 
    1011.5, 1011.5, 1011.4, 1011.4, 1011.5, 1011.5, 1011.3, 1011.4, 1011.4, 
    1011.6, 1011.5, 1012.2, 1012.4, 1012.4, 1012.7, 1013, 1012.9, 1013.3, 
    1013.3, 1013.6, 1013.7, 1014, 1014.3, 1014.5, 1014.9, 1015.1, 1015.5, 
    1015.9, 1016.2, 1016.6, 1016.9, 1016.6, 1017.2, 1017.4, 1017.7, 1017.6, 
    1017.9, 1018.5, 1018.6, 1018.8, 1018.8, 1018.7, 1018.7, 1018.7, 1018.6, 
    1018.7, 1018.6, 1018.4, 1018.2, 1017.9, 1017.7, 1018.1, 1017.7, 1017.3, 
    1017.1, 1016.8, 1016.5, 1016.2, 1015.5, 1015.3, 1015.1, 1015.1, 1014.5, 
    1014.1, 1013.8, 1013.6, 1013.6, 1013.1, 1012.6, 1012.4, 1012.2, 1011.7, 
    1011.3, 1011.1, 1010.8, 1010.8, 1010.3, 1009.8, 1009.6, 1008.9, 1009.8, 
    1008.1, 1007.8, 1007.1, 1006.4, 1006, 1005.4, 1004.6, 1003.8, 1003.3, 
    1002.3, 1001.9, 1001.3, 1001, 1000.2, 999.8, 999.4, 999.1, 998.7, 998.5, 
    997.8, 998, 998, 997.7, 997.6, 997.6, 997.4, 997.3, 997.4, 997.1, 996.9, 
    996.7, 996.4, 996.3, 995.8, 995.9, 996.1, 995.8, 995.5, 995.6, 995.4, 
    995.8, 996, 996.1, 996.2, 995.7, 996.4, 996.3, 996.2, 995.9, 995.1, 995, 
    995.8, 996, 996.3, 996, 996.4, 996.3, 996.2, 995.9, 996.1, 996.4, 996.6, 
    996.9, 997.4, 997.6, 997.9, 998.2, 998.6, 998.8, 999.2, 999.4, 999.9, 
    1000.2, 1000.9, 1001.2, 1001.5, 1002, 1002.3, 1002.7, 1003, 1003.4, 
    1003.6, 1003.9, 1003.9, 1004.5, 1004.8, 1005.2, 1005.3, 1005.7, 1005.9, 
    1006.1, 1006.4, 1006.6, 1006.5, 1006.6, 1006.6, 1006.8, 1006.8, 1006.8, 
    1006.9, 1006.9, 1007.1, 1007.2, 1007, 1007, 1006.9, 1006.9, 1006.9, 
    1007.1, 1007.4, 1007.6, 1007.8, 1007.9, 1008, 1008.1, 1008, 1007.9, 
    1007.9, 1007.7, 1007.5, 1007.4, 1007.4, 1007.4, 1007.2, 1007, 1006.9, 
    1006.6, 1006.4, 1006.2, 1005.9, 1005.4, 1005.1, 1005, 1004.8, 1004.7, 
    1004.5, 1004.1, 1004.1, 1003.8, 1003.3, 1003.1, 1002.9, 1002.7, 1002.7, 
    1002.5, 1002.3, 1002.1, 1002.2, 1002.1, 1001.9, 1001.7, 1001.5, 1001.4, 
    1001.3, 1001.1, 1001, 1000.9, 1000.9, 1001.1, 1001.1, 1000.9, 1000.8, 
    1000.7, 1000.4, 1000.4, 1000.1, 1000, 999.8, 999.5, 999.2, 998.9, 998.8, 
    998.8, 998.7, 998.6, 998.5, 998.8, 998.9, 999.1, 999.1, 999.2, 999.5, 
    999.7, 1000.1, 1000.2, 1000.5, 1000.8, 1001.2, 1001.6, 1001.8, 1002, 
    1002.1, 1002.2, 1002.5, 1002.8, 1002.9, 1003.1, 1003, 1003.4, 1003.2, 
    1003, 1002.9, 1003, 1003, 1002.7, 1002.2, 1002.5, 1002.5, 1002.5, 1002.3, 
    1002, 1001.1, 1000.3, 999.5, 998.7, 997.2, 996.3, 996.2, 995.5, 996, 996, 
    995.7, 995.4, 995.6, 995, 994.5, 994.5, 995.1, 994.3, 994.2, 994.5, 995, 
    994.7, 995.3, 995.3, 994.5, 994, 993.6, 994.1, 993.6, 994, 994.4, 994.1, 
    994.8, 995.3, 995.4, 995.8, 995.6, 995.8, 995.7, 995.7, 996.1, 996.4, 
    996, 996.2, 995.8, 996.1, 996.5, 996.9, 997, 997.3, 997.4, 997.6, 998, 
    998, 998.3, 998.7, 998.7, 999.1, 999.5, 999.4, 999.5, 999.6, 999.7, 1000, 
    1000.2, 1000.4, 1000.2, 1000.3, 1000.4, 1001.2, 1001.6, 1002.3, 1002.9, 
    1003.4, 1004, 1004.3, 1004.8, 1005.3, 1005.6, 1006.2, 1006.4, 1006.6, 
    1006.8, 1007.1, 1007.2, 1007.8, 1008.3, 1008.5, 1009.1, 1009.6, 1009.8, 
    1010.2, 1010.7, 1011.1, 1011.4, 1011.6, 1011.6, 1011.6, 1011.6, 1011.5, 
    1011.4, 1011.2, 1011, 1010.7, 1010.6, 1010.4, 1010.3, 1010.3, 1010.1, 
    1009.9, 1009.9, 1009.7, 1009.6, 1009.4, 1009.3, 1009.3, 1009.4, 1009.3, 
    1009.1, 1009, 1009, 1008.9, 1008.8, 1008.5, 1008.3, 1008.2, 1008.1, 1008, 
    1008, 1007.9, 1007.7, 1007.6, 1007.5, 1007.3, 1007.3, 1007.2, 1007, 
    1006.8, 1006.6, 1006.5, 1006.3, 1006.4, 1006.4, 1006.4, 1006.2, 1006, 
    1005.9, 1005.6, 1005.3, 1005.1, 1005, 1005, 1004.9, 1004.9, 1004.9, 
    1004.8, 1004.9, 1004.9, 1004.8, 1004.9, 1005, 1005.1, 1005.3, 1005.6, 
    1005.8, 1006.1, 1006.3, 1006.6, 1006.9, 1006.9, 1007.1, 1007.3, 1007.5, 
    1007.6, 1007.8, 1008.1, 1008.3, 1008.5, 1008.8, 1008.9, 1009.2, 1009.3, 
    1009.5, 1009.7, 1009.9, 1010.1, 1010.3, 1010.6, 1010.8, 1011, 1011.2, 
    1011.3, 1011.3, 1011.3, 1011.5, 1011.6, 1011.5, 1011.6, 1011.7, 1011.9, 
    1012, 1012, 1012.1, 1012.3, 1012.5, 1012.6, 1012.6, 1012.5, 1012.4, 
    1012.4, 1012.5, 1012.5, 1012.5, 1012.6, 1012.7, 1012.6, 1012.6, 1012.6, 
    1012.5, 1012.6, 1012.6, 1012.8, 1013, 1013.2, 1013.4, 1013.6, 1013.8, 
    1014, 1014.2, 1014.3, 1014.7, 1014.7, 1015.1, 1015.2, 1015.5, 1015.9, 
    1016.3, 1016.5, 1016.8, 1017.3, 1017.6, 1017.7, 1018.1, 1018.2, 1018.4, 
    1018.7, 1019.2, 1019.5, 1020, 1020.2, 1020.4, 1020.6, 1020.9, 1020.9, 
    1021, 1021.1, 1021.1, 1021.3, 1021.5, 1021.4, 1021.4, 1021.4, 1021.5, 
    1021.5, 1021.8, 1021.9, 1021.7, 1021.4, 1021.4, 1021.3, 1021.4, 1021.7, 
    1022, 1022, 1022.1, 1022.3, 1022.1, 1022.3, 1022.2, 1022.1, 1022, 1022, 
    1022, 1022, 1021.9, 1022, 1021.8, 1021.7, 1021.4, 1021.1, 1020.7, 1020.5, 
    1020.6, 1020.5, 1020.5, 1020.5, 1020.4, 1020.4, 1020.4, 1020.6, 1020.4, 
    1020.1, 1020, 1019.8, 1019.5, 1019.5, 1019.4, 1019.2, 1019.2, 1019.1, 
    1019, 1018.7, 1018.5, 1018.4, 1018.4, 1018.2, 1018.2, 1018, 1017.9, 
    1017.9, 1017.9, 1017.8, 1017.5, 1017.3, 1017.1, 1017.2, 1017, 1016.6, 
    1016.3, 1016.3, 1016.2, 1016, 1015.9, 1015.8, 1015.6, 1015.5, 1015.4, 
    1015.1, 1015, 1014.8, 1014.4, 1014.2, 1014.4, 1014.2, 1014.2, 1014.3, 
    1014.3, 1014.2, 1014.2, 1014, 1014.1, 1013.9, 1014, 1014.1, 1014.2, 1014, 
    1014.2, 1014, 1013.6, 1013.7, 1013.8, 1013.6, 1013.6, 1013.5, 1013.3, 
    1013.2, 1013.1, 1012.7, 1012.6, 1012.5, 1012.4, 1012.1, 1012, 1012, 
    1011.8, 1011.5, 1011.4, 1011.1, 1011.2, 1011.1, 1011.1, 1011.1, 1011, 
    1011, 1010.9, 1010.9, 1010.9, 1011, 1011.1, 1011.3, 1011.6, 1011.8, 1012, 
    1012.2, 1012.5, 1012.9, 1013.2, 1013.5, 1013.6, 1013.9, 1014.1, 1014.4, 
    1014.7, 1014.9, 1015.4, 1015.6, 1016, 1016.3, 1016.5, 1016.7, 1017, 
    1017.1, 1017.2, 1017.2, 1017.3, 1017.6, 1017.7, 1017.9, 1017.8, 1017.8, 
    1017.7, 1017.6, 1017.5, 1017.6, 1017.5, 1017.5, 1017.7, 1017.6, 1017.8, 
    1017.8, 1017.9, 1018, 1018, 1017.9, 1017.8, 1017.6, 1017.5, 1017.3, 
    1017.2, 1017.1, 1017.2, 1017.3, 1017.4, 1017.1, 1016.8, 1016.7, 1016.8, 
    1016.7, 1016.9, 1016.9, 1017, 1017.3, 1017.8, 1018, 1018.1, 1018.2, 
    1018.5, 1018.5, 1018.8, 1018.8, 1018.9, 1018.9, 1018.9, 1018.9, 1019.1, 
    1019.4, 1019.4, 1019.5, 1019.7, 1019.8, 1019.8, 1019.8, 1019.9, 1020, 
    1020.3, 1020.2, 1020.3, 1020.4, 1020.5, 1020.3, 1020, 1019.7, 1019.5, 
    1019, 1018.6, 1018.5, 1018.5, 1018.2, 1018, 1017.8, 1017.6, 1017.3, 
    1017.2, 1016.8, 1016.5, 1016.1, 1015.9, 1015.6, 1015.4, 1015.4, 1015.2, 
    1015, 1015, 1014.6, 1014.3, 1014.3, 1014.1, 1014.2, 1014.1, 1014.2, 
    1014.4, 1014.7, 1014.7, 1015, 1015.2, 1015.2, 1015.3, 1015.3, 1015.6, 
    1015.8, 1016.1, 1016.1, 1016.6, 1016.8, 1017.2, 1017.5, 1017.8, 1017.9, 
    1018.2, 1018.7, 1019, 1019, 1019.1, 1019.4, 1019.7, 1020.1, 1020.3, 
    1020.6, 1020.6, 1020.7, 1020.7, 1020.8, 1020.7, 1020.7, 1020.7, 1020.7, 
    1020.9, 1021.1, 1021.5, 1021.5, 1021.8, 1022, 1022, 1022.2, 1022.4, 
    1022.6, 1022.7, 1022.9, 1022.9, 1023, 1023.1, 1023.1, 1023.2, 1023.3, 
    1023.7, 1023.8, 1023.8, 1024, 1024, 1024.4, 1024.6, 1024.9, 1025.2, 
    1025.3, 1025.5, 1025.7, 1025.9, 1025.9, 1026.2, 1026.3, 1026.4, 1026.6, 
    1026.5, 1026.5, 1026.6, 1026.7, 1026.7, 1026.8, 1026.9, 1027, 1026.9, 
    1026.7, 1026.7, 1026.6, 1026.4, 1026.2, 1026.1, 1025.9, 1026.1, 1026, 
    1025.7, 1025.2, 1025.2, 1025, 1025, 1024.4, 1024.3, 1024.2, 1024.2, 
    1024.1, 1024, 1023.6, 1023.5, 1023.4, 1022.8, 1022.5, 1022.1, 1021.3, 
    1020.8, 1020.3, 1020, 1019.7, 1019.5, 1019.4, 1019.3, 1018.9, 1019, 
    1018.8, 1018.7, 1018.8, 1018.5, 1018.9, 1018.9, 1019, 1019.3, 1019.4, 
    1019.5, 1019.7, 1020, 1020.1, 1020.2, 1020.7, 1020.8, 1020.8, 1021.4, 
    1021.9, 1021.9, 1022.3, 1022.6, 1022.7, 1022.6, 1022.7, 1022.5, 1022.6, 
    1022.7, 1022.7, 1022.8, 1022.7, 1022.8, 1022.8, 1022.9, 1023, 1022.9, 
    1022.8, 1023, 1023.1, 1023.2, 1023.1, 1023.1, 1022.9, 1022.9, 1022.8, 
    1022.7, 1022.7, 1022.6, 1022.7, 1022.5, 1022.5, 1022.2, 1022.4, 1022.2, 
    1022.2, 1022.4, 1022.2, 1022.1, 1022.2, 1022.1, 1021.9, 1021.8, 1021.4, 
    1021.5, 1021.7, 1021.9, 1021.8, 1021.4, 1021.3, 1021.2, 1021.2, 1021, 
    1020.8, 1020.8, 1020.8, 1020.9, 1021.1, 1021, 1021.2, 1021.3, 1021.3, 
    1021.1, 1020.9, 1021, 1021.3, 1021.8, 1021.9, 1022, 1022.1, 1022.2, 
    1022.3, 1022.3, 1022.5, 1022.6, 1022.6, 1022.5, 1022.7, 1022.9, 1023.1, 
    1023.3, 1023.5, 1023.6, 1023.7, 1023.7, 1023.7, 1023.7, 1023.7, 1023.7, 
    1023.7, 1023.7, 1023.7, 1023.7, 1023.9, 1023.9, 1023.7, 1023.6, 1023.5, 
    1023.4, 1023.4, 1023.4, 1023.3, 1023.3, 1023.3, 1023.1, 1022.9, 1022.7, 
    1022.6, 1022.5, 1022.4, 1022.3, 1022, 1021.7, 1021.3, 1021.1, 1020.8, 
    1020.6, 1020.5, 1020.2, 1020, 1019.8, 1019.6, 1019.3, 1018.9, 1018.7, 
    1018.6, 1018.1, 1017.8, 1017.5, 1017.4, 1017.2, 1016.9, 1016.6, 1016.3, 
    1016, 1015.9, 1015.6, 1015.3, 1015.2, 1014.9, 1014.8, 1014.5, 1014.3, 
    1014.2, 1014.2, 1014.2, 1014.1, 1014, 1013.9, 1013.8, 1013.6, 1013.4, 
    1013.3, 1013.3, 1013.4, 1013.4, 1013.3, 1013.3, 1013.1, 1012.9, 1012.5, 
    1012.1, 1011.9, 1011.4, 1011.6, 1011.6, 1011.5, 1011.2, 1011, 1010.7, 
    1010.4, 1010, 1009.1, 1008.3, 1007.6, 1007.3, 1007.2, 1007.1, 1007.6, 
    1007.2, 1008.2, 1008.4, 1008.9, 1009, 1009.3, 1009.1, 1009.5, 1009.4, 
    1009.8, 1009.5, 1009.5, 1009.2, 1009.6, 1010.4, 1010.6, 1010.9, 1010.7, 
    1011, 1011.1, 1011.4, 1012, 1012.1, 1012.6, 1012.5, 1012.7, 1012.8, 
    1012.6, 1012.8, 1013, 1013.1, 1013.4, 1013.6, 1013.9, 1013.9, 1014, 
    1013.9, 1014, 1013.9, 1013.9, 1013.9, 1013.9, 1013.9, 1014, 1014.2, 
    1014.4, 1014.5, 1014.6, 1014.8, 1014.8, 1015, 1015.2, 1015.3, 1015.1, 
    1014.8, 1014.8, 1014.4, 1014.3, 1013.9, 1013.8, 1013.7, 1013.7, 1013.8, 
    1013.7, 1014, 1013.9, 1013.8, 1013.6, 1013.9, 1014, 1014, 1014, 1014.3, 
    1014.4, 1014.6, 1014.8, 1014.9, 1014.9, 1014.9, 1014.8, 1014.8, 1015, 
    1015.4, 1015.5, 1015.6, 1015.8, 1016, 1016, 1016.3, 1016.1, 1016.1, 
    1016.2, 1016.3, 1016.4, 1016.3, 1016.4, 1016.7, 1016.8, 1016.8, 1016.6, 
    1016.6, 1016.7, 1016.5, 1016.4, 1016.4, 1016.4, 1016.7, 1016.8, 1016.9, 
    1017, 1017, 1016.9, 1016.9, 1016.8, 1016.6, 1016.7, 1016.6, 1016.3, 
    1016.2, 1016.2, 1016.2, 1016.2, 1016.2, 1016.2, 1016.1, 1016.1, 1015.9, 
    1015.7, 1015.4, 1015.3, 1015.2, 1014.9, 1014.8, 1014.8, 1014.8, 1014.8, 
    1014.9, 1014.9, 1014.7, 1014.7, 1014.6, 1014.7, 1014.6, 1014.7, 1014.7, 
    1014.7, 1014.7, 1014.8, 1014.7, 1014.7, 1014.4, 1014.2, 1014, 1013.9, 
    1014, 1013.7, 1013.6, 1013.3, 1013.2, 1012.6, 1012.4, 1012.1, 1011.7, 
    1011.1, 1011, 1010.5, 1010.5, 1010.1, 1009.6, 1009.1, 1008.8, 1008.6, 
    1008.3, 1007.7, 1007, 1006.6, 1006, 1006.4, 1005.8, 1005.6, 1005.3, 
    1005.1, 1005.2, 1004.9, 1004.6, 1004.4, 1004.1, 1003.9, 1003.8, 1003.5, 
    1004, 1004, 1003.8, 1003.7, 1003.6, 1003.5, 1003.4, 1003.4, 1003.1, 
    1003.1, 1003.1, 1003, 1002.7, 1002.7, 1002.7, 1002.7, 1002.7, 1002.7, 
    1002.6, 1002.7, 1002.7, 1002.8, 1002.9, 1003, 1003.4, 1003.5, 1003.6, 
    1003.8, 1004, 1004.2, 1004.5, 1004.8, 1005.2, 1005.3, 1005.7, 1006, 
    1006.2, 1006.6, 1007, 1007.3, 1007.7, 1008.1, 1008.4, 1008.9, 1009.4, 
    1009.7, 1010.1, 1010.7, 1011.3, 1011.8, 1012.3, 1012.8, 1013.5, 1014, 
    1014.4, 1014.8, 1015.3, 1015.8, 1016.1, 1016.4, 1016.8, 1017.3, 1017.6, 
    1017.9, 1018.2, 1018.5, 1018.9, 1019.2, 1019.4, 1019.7, 1019.9, 1020.1, 
    1020.3, 1020.6, 1021, 1021.2, 1021.2, 1021.3, 1021.3, 1021.2, 1021.3, 
    1021.4, 1021.4, 1021.7, 1021.8, 1021.9, 1021.9, 1021.9, 1021.9, 1021.7, 
    1021.7, 1021.3, 1021, 1020.9, 1020.8, 1020.7, 1020.4, 1020.4, 1019.9, 
    1019.5, 1019.8, 1019.5, 1019.3, 1019.4, 1018.8, 1018.5, 1018.3, 1018, 
    1017.7, 1017.1, 1016.9, 1016.1, 1015.2, 1015, 1015.3, 1015.3, 1014.5, 
    1013.8, 1013.4, 1013.2, 1013, 1012.7, 1012.6, 1012.7, 1012.3, 1012.8, 
    1012.8, 1012.9, 1013.1, 1013.3, 1013.6, 1013.5, 1013.8, 1013.8, 1014, 
    1014.2, 1014.4, 1014.5, 1014.6, 1014.8, 1014.9, 1015.3, 1015.7, 1016, 
    1016.4, 1016.7, 1016.9, 1017.1, 1017.5, 1017.8, 1018.1, 1018.4, 1018.7, 
    1019, 1019.2, 1019.4, 1019.8, 1020, 1020.2, 1020.3, 1020.2, 1020.4, 
    1020.5, 1020.5, 1020.5, 1020.4, 1020.5, 1020.7, 1020.9, 1020.9, 1021.1, 
    1021.2, 1021.2, 1021, 1021, 1021.1, 1020.9, 1020.8, 1020.6, 1020.3, 
    1020.2, 1020.4, 1020.3, 1020.2, 1019.8, 1019.9, 1019.7, 1019.5, 1019.5, 
    1019.5, 1019.1, 1019.2, 1019.7, 1019.8, 1019.9, 1020.1, 1020.4, 1020.4, 
    1020.6, 1020.4, 1020.3, 1020.4, 1020.7, 1021, 1021.1, 1021.2, 1021.2, 
    1021.3, 1021.5, 1021.5, 1021.5, 1021.7, 1021.4, 1021.3, 1021.2, 1021.4, 
    1021.7, 1022, 1022.1, 1022.1, 1021.9, 1021.8, 1021.5, 1021.5, 1021.3, 
    1021.2, 1020.9, 1020.8, 1020.8, 1020.9, 1020.8, 1020.9, 1020.8, 1020.8, 
    1020.6, 1020.2, 1019.7, 1019.6, 1019.5, 1019.5, 1019.7, 1019.7, 1019.7, 
    1019.5, 1019.3, 1019.1, 1018.9, 1018.8, 1019, 1018.8, 1018.7, 1018.8, 
    1018.8, 1018.9, 1019, 1019, 1019, 1019.2, 1019.3, 1019.4, 1019.5, 1019.7, 
    1020.2, 1020.5, 1020.7, 1021, 1021.2, 1021.3, 1021.5, 1021.8, 1021.9, 
    1022.1, 1022.2, 1022.4, 1022.5, 1022.6, 1022.9, 1023, 1023, 1023.1, 1023, 
    1023, 1023, 1023, 1022.9, 1022.7, 1022.4, 1022.2, 1022.1, 1021.9, 1021.3, 
    1021.3, 1021, 1020.7, 1020.3, 1019.9, 1019.8, 1019.2, 1018.7, 1018.1, 
    1017.9, 1017.8, 1017.4, 1017, 1016.7, 1015.6, 1015.4, 1014.7, 1014.2, 
    1013.8, 1013.5, 1013.3, 1013.2, 1013.1, 1012.9, 1012.7, 1012.5, 1012.5, 
    1012.3, 1012.2, 1011.9, 1011.7, 1011.5, 1011.4, 1011.1, 1010.9, 1010.9, 
    1010.7, 1010.5, 1010.5, 1010.2, 1010.2, 1010.1, 1010.1, 1010, 1010, 1010, 
    1010.1, 1010.3, 1010.1, 1010.1, 1010.2, 1010.2, 1010.2, 1010.2, 1010.1, 
    1010.2, 1010.3, 1010.3, 1010.6, 1010.8, 1011, 1011.1, 1011.3, 1011.4, 
    1011.2, 1011.4, 1011.5, 1011.5, 1011.5, 1011.7, 1011.8, 1011.9, 1011.9, 
    1011.9, 1012, 1012.1, 1011.9, 1011.7, 1011.5, 1011.7, 1011.8, 1011.8, 
    1011.7, 1011.7, 1011.8, 1011.7, 1011.5, 1011.4, 1011.2, 1011.2, 1011.1, 
    1010.9, 1010.9, 1011, 1011, 1010.9, 1011.1, 1011.1, 1011.1, 1011.2, 
    1011.1, 1011.2, 1011.1, 1011.2, 1011.3, 1011.3, 1011.3, 1011.6, 1011.7, 
    1011.8, 1011.9, 1011.8, 1011.8, 1011.8, 1011.8, 1011.8, 1012, 1012.2, 
    1012.4, 1012.7, 1012.9, 1013, 1013.1, 1013.4, 1013.5, 1013.7, 1013.8, 
    1013.9, 1014.1, 1014.2, 1014.4, 1014.7, 1014.8, 1014.9, 1015.1, 1015.1, 
    1015.1, 1015.1, 1015.1, 1015, 1015.1, 1015.1, 1015.1, 1015.2, 1015.2, 
    1015.2, 1015, 1015.2, 1015.2, 1015, 1014.8, 1014.9, 1015.1, 1015, 1015, 
    1014.9, 1014.8, 1014.8, 1014.6, 1014.3, 1014.1, 1014.2, 1014.2, 1014.4, 
    1014.5, 1014.6, 1014.6, 1014.6, 1014.6, 1014.5, 1014.3, 1014.1, 1014, 
    1013.8, 1013.6, 1013.4, 1013.2, 1013.1, 1012.9, 1012.9, 1012.7, 1012.5, 
    1012.2, 1011.9, 1011.6, 1011.2, 1010.9, 1010.8, 1010.7, 1010.7, 1010.6, 
    1010.4, 1010.2, 1010.2, 1010.1, 1010.1, 1010.3, 1010.2, 1010.1, 1010.2, 
    1010.3, 1010.4, 1010.3, 1010.5, 1010.6, 1010.8, 1011.1, 1011.4, 1011.6, 
    1011.9, 1012.2, 1012.5, 1013, 1013.4, 1014, 1014.7, 1015.3, 1015.8, 
    1016.5, 1017, 1017.5, 1017.9, 1018.2, 1018.6, 1019.3, 1019.7, 1020.4, 
    1021.2, 1021.9, 1022.2, 1022.7, 1023.2, 1023.6, 1023.9, 1024.1, 1024.4, 
    1024.6, 1025.1, 1025.4, 1025.6, 1025.9, 1026.3, 1026.3, 1026.1, 1026.2, 
    1026.4, 1026.5, 1026.8, 1026.8, 1027.2, 1027.4, 1027.7, 1027.9, 1028, 
    1028, 1028.1, 1028.1, 1028.1, 1028, 1027.9, 1027.6, 1027.4, 1027.3, 
    1027.1, 1027.2, 1026.9, 1026.6, 1026, 1025.7, 1025.7, 1025.5, 1025.1, 
    1025, 1025, 1025, 1024.9, 1024.6, 1024.6, 1024.2, 1023.8, 1023.4, 1022.9, 
    1022.5, 1021.9, 1021.5, 1021, 1020.5, 1020.2, 1020.1, 1019.7, 1019.6, 
    1019.1, 1018.8, 1018.4, 1017.7, 1016.9, 1016.1, 1015.8, 1015.3, 1015.2, 
    1014.9, 1014.8, 1014.3, 1014.1, 1013.4, 1013.3, 1013.3, 1013.2, 1012.8, 
    1012.8, 1013, 1012.9, 1012.7, 1013.2, 1013.2, 1013, 1013.2, 1013.1, 
    1012.8, 1012.6, 1012.4, 1012.4, 1012.3, 1012.4, 1012.3, 1012.3, 1012.6, 
    1012.6, 1012.5, 1012.4, 1012.4, 1012.6, 1012.8, 1012.9, 1013.1, 1013.1, 
    1013, 1013, 1013.2, 1012.3, 1011.5, 1010.8, 1010.2, 1010.5, 1010.4, 
    1010.7, 1010.5, 1010.6, 1011.1, 1011.1, 1011.3, 1011.6, 1011.8, 1011.8, 
    1012, 1012, 1012, 1012.3, 1012.6, 1012.7, 1012.7, 1012.5, 1012.4, 1012.3, 
    1012.6, 1012.4, 1012.5, 1012.6, 1012.6, 1012.8, 1013.2, 1013.4, 1013.6, 
    1013.8, 1014.2, 1014.8, 1015.4, 1015.7, 1016.2, 1016.8, 1017.3, 1018, 
    1018.2, 1018.7, 1019.1, 1019.4, 1019.8, 1020.3, 1020.5, 1020.8, 1021.2, 
    1021.5, 1022, 1022.6, 1022.9, 1023.1, 1023.5, 1023.6, 1024, 1024.2, 
    1024.3, 1024.5, 1024.6, 1024.8, 1025.2, 1025.6, 1025.7, 1026.1, 1026.3, 
    1026.3, 1026.6, 1026.8, 1026.8, 1026.8, 1026.8, 1027, 1026.9, 1027.2, 
    1027.2, 1027.1, 1027.2, 1027.1, 1026.7, 1026.4, 1026, 1025.8, 1025.1, 
    1024.7, 1023.8, 1023.5, 1023.2, 1022, 1021.1, 1020.3, 1019.4, 1018.5, 
    1017.8, 1016.8, 1015.9, 1015.3, 1015, 1014.9, 1014.8, 1014.6, 1014.3, 
    1014.2, 1014.2, 1014.1, 1013.9, 1014.2, 1014.2, 1014.1, 1014.2, 1014.3, 
    1014.5, 1014.5, 1014.8, 1014.8, 1014.8, 1014.9, 1015.1, 1015, 1015, 
    1015.2, 1015.3, 1015.6, 1015.9, 1016.1, 1016.3, 1016.6, 1016.7, 1016.8, 
    1016.9, 1017.3, 1017.3, 1017.5, 1017.6, 1017.8, 1017.9, 1018.3, 1018.2, 
    1018.2, 1018.1, 1018.2, 1018.4, 1018.4, 1018.5, 1018.3, 1018.5, 1018.8, 
    1018.8, 1018.8, 1019.1, 1019.2, 1019.1, 1019.1, 1019.2, 1019.2, 1019.1, 
    1019.1, 1019, 1019, 1019, 1018.9, 1018.9, 1018.9, 1018.9, 1018.7, 1018.5, 
    1018.4, 1018.2, 1017.9, 1017.7, 1017.5, 1017.4, 1017.2, 1017.1, 1016.9, 
    1016.7, 1016.7, 1016.7, 1016.7, 1016.5, 1016.4, 1016.4, 1016.5, 1016.5, 
    1016.7, 1016.9, 1016.9, 1017.2, 1017.3, 1017.2, 1017.2, 1017.3, 1017.4, 
    1017.5, 1017.5, 1017.7, 1017.9, 1018, 1018.1, 1018.2, 1018.2, 1018.1, 
    1018, 1017.9, 1017.8, 1017.9, 1018.2, 1018.1, 1018.3, 1018.5, 1018.7, 
    1018.4, 1018.2, 1018.2, 1018, 1018, 1018, 1017.8, 1017.9, 1017.8, 1017.6, 
    1017.2, 1017.4, 1017.2, 1016.6, 1016.2, 1015.7, 1015, 1014.5, 1014.2, 
    1014.2, 1013.6, 1013.2, 1012.5, 1012.1, 1012, 1011.8, 1011.2, 1010.5, 
    1010.5, 1010.4, 1010, 1009.9, 1009.6, 1009.4, 1009, 1008.9, 1008.8, 
    1008.8, 1008.8, 1009.2, 1009.1, 1009.1, 1009.3, 1009.4, 1009.8, 1009.9, 
    1010, 1010.3, 1010.2, 1010.4, 1010.3, 1010.2, 1010.1, 1009.9, 1009.8, 
    1009.7, 1009.8, 1009.5, 1009.3, 1009.2, 1009, 1008.8, 1008.7, 1008.4, 
    1008, 1008.1, 1008.1, 1008.1, 1008, 1007.8, 1007.6, 1007.3, 1007.3, 
    1007.2, 1007.4, 1007.5, 1007.3, 1007.2, 1007.7, 1007.8, 1007.8, 1008.2, 
    1008.4, 1008.8, 1009.1, 1009.1, 1009.5, 1009.8, 1010.2, 1010.8, 1011, 
    1011.9, 1012, 1012.4, 1013.3, 1013.7, 1014.3, 1014.9, 1015.3, 1015.6, 
    1016.3, 1016.5, 1016.7, 1017, 1017.5, 1017.8, 1018.3, 1018.4, 1018.8, 
    1019, 1019.3, 1019.7, 1019.9, 1020.2, 1020.4, 1020.6, 1020.6, 1020.6, 
    1020.7, 1020.7, 1020.7, 1020.6, 1020.5, 1020.2, 1020.1, 1019.8, 1019.6, 
    1019.4, 1019.5, 1019.3, 1019.1, 1018.8, 1018.6, 1018.2, 1018, 1017.6, 
    1017, 1016.6, 1016.3, 1015.9, 1015.3, 1014.9, 1014.6, 1014.1, 1013.8, 
    1013.4, 1013.2, 1012.8, 1012.2, 1011.8, 1011.4, 1011.3, 1011.1, 1010.9, 
    1010.8, 1010.6, 1010.5, 1010.3, 1010.3, 1010.4, 1010.1, 1010, 1009.7, 
    1009.8, 1009.9, 1010, 1009.5, 1009.6, 1009.6, 1009.3, 1008.9, 1008.4, 
    1008, 1007.6, 1007.3, 1007.2, 1006.9, 1006.6, 1006.4, 1006.2, 1006.1, 
    1006.1, 1006, 1005.8, 1005.7, 1005.6, 1005.7, 1005.7, 1005.8, 1006, 
    1006.2, 1006.3, 1006.4, 1006.6, 1006.8, 1007, 1007.1, 1007.4, 1007.8, 
    1008.1, 1008.6, 1009, 1009.2, 1009.5, 1009.8, 1010, 1010.3, 1010.4, 
    1010.6, 1010.7, 1010.9, 1011.1, 1011.3, 1011.3, 1011.4, 1011.4, 1011.3, 
    1011.2, 1011.3, 1011.2, 1011, 1011, 1010.9, 1010.8, 1010.9, 1010.8, 
    1010.7, 1010.6, 1010.4, 1010.2, 1010, 1010, 1009.9, 1009.6, 1009.4, 
    1009.1, 1009, 1008.5, 1008, 1007.4, 1007.1, 1006.8, 1006.4, 1005.7, 
    1005.4, 1004.7, 1003.9, 1003.1, 1002.4, 1002, 1000.8, 999.8, 998.6, 
    997.8, 997.2, 997.2, 997.4, 997.7, 998.2, 998.9, 999.2, 999.7, 1000.1, 
    1000.3, 1000.6, 1001, 1001.2, 1001.1, 1001.5, 1002, 1002.4, 1002.4, 
    1002.6, 1003, 1003.4, 1003.5, 1003.5, 1003.4, 1003.8, 1003.9, 1004, 
    1004.1, 1004.5, 1004.8, 1005.2, 1005.3, 1005.4, 1005.7, 1005.8, 1006.1, 
    1006.1, 1005.9, 1006.3, 1006.6, 1006.9, 1007.4, 1008.2, 1008.7, 1009.3, 
    1009.9, 1010.7, 1011.2, 1011.7, 1012.1, 1012.3, 1012.6, 1012.9, 1012.5, 
    1013.3, 1013, 1012.7, 1012.8, 1012.2, 1011.6, 1010.8, 1010.4, 1009.7, 
    1009.1, 1008.8, 1008.7, 1008.7, 1008.6, 1008.6, 1008.7, 1008.9, 1009.1, 
    1009.2, 1008.9, 1008.9, 1009.1, 1009.4, 1009.4, 1009.8, 1010.1, 1010.1, 
    1010.1, 1009.9, 1009.8, 1009.5, 1009, 1008.5, 1008.2, 1007.4, 1007.2, 
    1006.8, 1006.2, 1005.2, 1004.6, 1004.3, 1004.1, 1004.2, 1004.6, 1004.5, 
    1005.2, 1005.5, 1006.7, 1007.1, 1007.8, 1008.3, 1008.7, 1009.2, 1009.8, 
    1010.5, 1011.3, 1012.3, 1012.9, 1013.6, 1014, 1014.2, 1014.3, 1014.5, 
    1014.9, 1014.7, 1014.5, 1014.2, 1014.2, 1014, 1013.8, 1013.6, 1013.3, 
    1013.1, 1013, 1012.9, 1012.7, 1012.5, 1012.7, 1013.4, 1013.6, 1013.9, 
    1014, 1014.7, 1015.1, 1015.5, 1015.4, 1016, 1016.2, 1016.4, 1016.8, 
    1016.9, 1016.9, 1017, 1017.2, 1017.3, 1017.2, 1017.4, 1017.2, 1017.1, 
    1016.9, 1016.7, 1016.3, 1015.9, 1015.5, 1014.9, 1014.5, 1013.9, 1013.6, 
    1013.5, 1013.1, 1012.7, 1012.1, 1011.6, 1011.3, 1011.1, 1010.9, 1010.7, 
    1010.7, 1010.5, 1010.6, 1010.9, 1011, 1011.1, 1011.3, 1011.4, 1011.9, 
    1012.2, 1012.7, 1013.6, 1014, 1014.5, 1015.1, 1015.7, 1016.3, 1016.6, 
    1017.3, 1017.5, 1017.8, 1018, 1018.2, 1018.3, 1018.7, 1018.9, 1019.1, 
    1019.1, 1019.2, 1019.3, 1019.1, 1019.1, 1018.8, 1018.6, 1018.4, 1018.4, 
    1018.5, 1018.3, 1018.1, 1017.9, 1017.8, 1017.5, 1017.4, 1017.1, 1016.7, 
    1016.6, 1016.3, 1015.9, 1015.3, 1014.9, 1014.7, 1014.4, 1013.9, 1013.5, 
    1013.3, 1013, 1012.9, 1012.6, 1012.7, 1012.5, 1012.5, 1012.6, 1012.7, 
    1013, 1013, 1013, 1013.2, 1013.5, 1013.5, 1013.6, 1013.9, 1013.9, 1014, 
    1014, 1014.2, 1014.3, 1014.4, 1014.6, 1014.6, 1015, 1015, 1014.9, 1015, 
    1015.2, 1015, 1014.9, 1014.9, 1015, 1015.1, 1015.2, 1015.4, 1015.5, 
    1015.3, 1015.1, 1014.9, 1014.5, 1014.2, 1014.4, 1014.3, 1014.4, 1014.4, 
    1014.3, 1013.9, 1013.7, 1013.4, 1013.4, 1013.5, 1013.5, 1013.6, 1013.8, 
    1014.2, 1014.3, 1014.3, 1014.1, 1014.1, 1014.2, 1014.1, 1014, 1014, 
    1013.6, 1013.3, 1013.3, 1013.5, 1013.5, 1013.2, 1013.4, 1013.4, 1013.5, 
    1013.4, 1013.2, 1013, 1012.9, 1012.9, 1012.8, 1012.8, 1012.8, 1012.9, 
    1012.9, 1013, 1013.1, 1013.1, 1013.2, 1013.3, 1013.1, 1013.4, 1013.9, 
    1014.3, 1014.7, 1014.9, 1015.3, 1015.8, 1016.2, 1016.6, 1016.6, 1016.6, 
    1016.8, 1016.8, 1017.3, 1017.9, 1018.4, 1018.6, 1019, 1019.1, 1019, 
    1018.8, 1018.8, 1018.7, 1018.5, 1018.3, 1018, 1017.8, 1017.6, 1017.2, 
    1016.8, 1016.3, 1015.9, 1015.3, 1014.7, 1014.3, 1013.9, 1013.5, 1012.9, 
    1012.7, 1012.7, 1012.1, 1011.9, 1011.6, 1011.2, 1010.7, 1010.3, 1010.2, 
    1009.9, 1009.7, 1010, 1010.2, 1010, 1010, 1009.7, 1009.7, 1009.7, 1009.8, 
    1009.8, 1009.8, 1010.1, 1010.5, 1010.6, 1010.5, 1010.6, 1010.7, 1011.1, 
    1011.4, 1011.5, 1011.6, 1011.6, 1011.8, 1011.8, 1012.2, 1012.3, 1012.5, 
    1012.6, 1012.6, 1012.5, 1012.5, 1012.4, 1012.4, 1012.4, 1012.5, 1012.7, 
    1012.8, 1012.7, 1012.8, 1012.9, 1012.9, 1012.9, 1012.9, 1012.8, 1012.8, 
    1012.7, 1012.8, 1012.7, 1012.7, 1012.6, 1012.6, 1012.8, 1012.8, 1012.7, 
    1012.7, 1012.7, 1012.6, 1012.6, 1012.6, 1012.7, 1013, 1013, 1013.3, 
    1013.6, 1013.7, 1013.9, 1013.9, 1014.1, 1014.3, 1014.4, 1014.6, 1014.9, 
    1015.3, 1015.3, 1015.6, 1015.9, 1016.1, 1016.4, 1016.5, 1016.7, 1017, 
    1017.3, 1017.6, 1017.9, 1018.1, 1018.6, 1019.2, 1019.5, 1019.9, 1020.3, 
    1020.5, 1020.7, 1021, 1021.4, 1021.9, 1022.4, 1022.9, 1023.1, 1023.4, 
    1023.5, 1023.9, 1024.1, 1024.4, 1024.7, 1024.9, 1025.3, 1025.7, 1025.9, 
    1026.1, 1026.5, 1026.9, 1027.2, 1027.4, 1027.7, 1027.9, 1028.1, 1028.2, 
    1028.5, 1028.5, 1028.5, 1028.3, 1027.9, 1027.8, 1027.7, 1027.7, 1027.3, 
    1026.7, 1026.1, 1025.4, 1024.7, 1023.8, 1023.1, 1022.1, 1021.2, 1020.4, 
    1019.5, 1018.4, 1017.4, 1016.5, 1015.3, 1014.3, 1013.1, 1012, 1011.1, 
    1010.6, 1010, 1009.5, 1009.3, 1008.8, 1008.1, 1007.3, 1006.4, 1005.3, 
    1004.4, 1003.1, 1002.4, 1001.1, 999.8, 998.1, 996.3, 994.3, 991.8, 988.7, 
    985.3, 981.8, 978.8, 975.3, 972.3, 970.2, 967.9, 966.6, 966.1, 966.1, 
    965.9, 965.9, 966.2, 966.3, 967, 967.8, 968.8, 970.1, 971.5, 973.1, 
    974.9, 976.6, 978.2, 979.4, 980.9, 982.4, 983.5, 984.5, 985.6, 986.7, 
    987.8, 988.5, 989.4, 990.2, 990.7, 991.3, 991.8, 992, 992.6, 993.1, 
    993.5, 994, 994.1, 994.6, 995, 995.4, 995.6, 995.7, 995.9, 996.1, 996.2, 
    996.5, 996.7, 996.7, 996.6, 996.7, 997, 997, 997, 997.3, 997, 997.1, 
    997.2, 997.3, 997.2, 997.3, 997.3, 997.6, 997.9, 998, 998.2, 998.5, 
    998.7, 998.8, 998.9, 999.2, 999.4, 999.4, 999.7, 999.7, 1000, 1000.2, 
    1000.3, 1000.6, 1000.9, 1001.1, 1001.4, 1001.7, 1001.9, 1002.3, 1002.7, 
    1003.1, 1003.5, 1004, 1004.5, 1004.7, 1005, 1005.3, 1005.6, 1005.8, 
    1006.1, 1006.3, 1006.4, 1006.6, 1006.8, 1007.3, 1007.4, 1007.6, 1008, 
    1008.3, 1008.7, 1008.7, 1008.9, 1009.4, 1009.6, 1010.1, 1010.7, 1011.1, 
    1011.5, 1011.9, 1012.4, 1012.9, 1013.3, 1013.7, 1014.1, 1014.6, 1014.9, 
    1015.5, 1016.1, 1016.6, 1017, 1017.5, 1018.1, 1018.7, 1019.2, 1019.9, 
    1020.4, 1021, 1021.5, 1022.2, 1022.7, 1023.2, 1023.7, 1024.4, 1025.2, 
    1025.4, 1025.5, 1025.7, 1026.3, 1026.3, 1026.7, 1026.9, 1027.3, 1027.4, 
    1027.6, 1027.7, 1027.9, 1028, 1027.5, 1027.5, 1027.3, 1027.1, 1027.1, 
    1027.2, 1027.3, 1027.4, 1027.5, 1027.6, 1027.6, 1027.8, 1028.2, 1028, 
    1028, 1028.3, 1028.5, 1028.8, 1029, 1029, 1029.1, 1029, 1029.2, 1029.6, 
    1029.6, 1029.6, 1029.9, 1030.1, 1030.6, 1030.8, 1031.3, 1031.7, 1031.6, 
    1031.7, 1031.8, 1032, 1032.1, 1032.2, 1031.9, 1031.9, 1031.8, 1031.8, 
    1032.1, 1032, 1031.7, 1031.3, 1031.2, 1031.1, 1031, 1030.9, 1030.8, 
    1030.6, 1030.5, 1030.5, 1030.5, 1030.4, 1030.3, 1030.1, 1029.8, 1029.5, 
    1029.4, 1029.1, 1028.7, 1028.6, 1028.7, 1028.3, 1028.2, 1028, 1027.9, 
    1027.7, 1027.3, 1027.1, 1026.7, 1026.3, 1025.7, 1025.4, 1025.5, 1025.5, 
    1025.5, 1025.5, 1025.2, 1025, 1025.1, 1025.2, 1025.1, 1024.7, 1024.6, 
    1024.2, 1023.8, 1023.5, 1023.3, 1022.8, 1022.5, 1022.3, 1021.8, 1021.3, 
    1020.9, 1020.5, 1020.2, 1019.9, 1019.5, 1019.2, 1018.8, 1018.5, 1018, 
    1017.4, 1016.8, 1016.2, 1015.6, 1015, 1014, 1013.2, 1012.4, 1011.6, 
    1010.8, 1010.5, 1009.9, 1009.4, 1009.4, 1009.1, 1008.8, 1008.4, 1008, 
    1007.7, 1007.3, 1006.9, 1006.7, 1006.3, 1005.7, 1005.3, 1005, 1004.5, 
    1004.3, 1004.1, 1003.7, 1003.6, 1003.5, 1003.4, 1003.4, 1003.5, 1003.4, 
    1003.6, 1003.9, 1004.2, 1004.5, 1004.9, 1005.3, 1005.6, 1006, 1006.4, 
    1006.8, 1007.2, 1007.4, 1007.6, 1007.8, 1007.8, 1008.1, 1008.2, 1008.4, 
    1008.6, 1008.7, 1008.7, 1008.7, 1008.8, 1008.9, 1008.9, 1008.9, 1009, 
    1009, 1009.1, 1009.1, 1009.3, 1009.3, 1009.5, 1009.6, 1009.9, 1010.2, 
    1010.5, 1010.6, 1011, 1011.1, 1011.2, 1011.2, 1011.6, 1011.8, 1012, 
    1012.3, 1012.6, 1012.7, 1012.6, 1012.7, 1012.4, 1011.9, 1011.6, 1011.2, 
    1010.6, 1009.9, 1009.6, 1008.9, 1008.5, 1007.9, 1007.2, 1006.4, 1005.7, 
    1005.3, 1005.1, 1004.6, 1004.6, 1004.5, 1004.2, 1004, 1003.5, 1003.3, 
    1003.1, 1002.7, 1001.8, 1000.9, 1000.6, 999.9, 998.6, 997.3, 995.9, 
    995.1, 994.1, 992.9, 991.7, 990.6, 989.6, 988.7, 987.6, 986.5, 985.3, 
    984.5, 983.7, 983.1, 982.5, 981.7, 981.1, 981.1, 981.4, 981.3, 981.8, 
    982.5, 983, 983.7, 984.6, 985.4, 986.2, 987, 987.7, 988.2, 989, 989.7, 
    990.2, 991, 991.6, 992.2, 992.9, 993.6, 994.4, 995, 995.6, 996.1, 996.9, 
    997.5, 998.1, 998.7, 999.3, 999.9, 1000.7, 1001.5, 1002.2, 1002.9, 
    1003.4, 1003.8, 1004.3, 1004.9, 1005.2, 1005.1, 1005.6, 1005.6, 1005.9, 
    1006.4, 1006.3, 1006.5, 1006.5, 1006.7, 1006.6, 1006.5, 1006.9, 1006.5, 
    1006.4, 1006.4, 1006.2, 1006, 1005.6, 1005.1, 1004.6, 1003.8, 1003.1, 
    1002.1, 1001.4, 1000.5, 999.9, 999, 998.5, 998, 997.3, 996.4, 995.5, 
    995.4, 995, 994.6, 994.1, 993.8, 993.1, 992.9, 992.5, 992.2, 992.2, 
    992.2, 991.9, 992, 992.6, 992.6, 992.9, 993.1, 993.3, 993.9, 994.9, 
    995.7, 996.1, 997, 997.6, 998.7, 999.5, 1000.6, 1001.5, 1002.3, 1003.4, 
    1004.3, 1005.1, 1005.8, 1006.6, 1007.1, 1007.4, 1007.8, 1007.9, 1008.3, 
    1008.4, 1008.6, 1008.4, 1008.3, 1008, 1007.7, 1007.4, 1007.2, 1007, 
    1006.8, 1006.3, 1005.7, 1005.2, 1004.9, 1004.7, 1004.3, 1003.9, 1003.5, 
    1003, 1002.6, 1001.9, 1001.4, 1000.9, 1000.7, 1000.4, 1000, 999.7, 999.3, 
    998.8, 998.4, 998.3, 998, 997.4, 996.9, 996.4, 996.2, 996.3, 996.1, 
    995.8, 995.3, 995.4, 995.5, 995.6, 995.7, 995.5, 995.3, 995.3, 995.2, 
    995.3, 995.1, 995.1, 995, 994.8, 994.9, 994.8, 994.8, 994.8, 994.9, 995, 
    995, 994.9, 995.1, 995, 995.1, 995.4, 995.3, 995.4, 995.3, 995.1, 995.1, 
    994.7, 994.6, 994.1, 993.9, 993.9, 993.6, 993.3, 993.3, 992.5, 992.1, 
    992, 991.7, 991, 990.7, 990.7, 990.3, 990.1, 990.4, 990.3, 990, 989.8, 
    989.1, 988.4, 987.5, 986.5, 985.3, 984.3, 983.4, 982.5, 981.5, 980.6, 
    980.1, 980, 979.1, 978.3, 977.7, 977.4, 977, 976.5, 976.2, 976.2, 976.3, 
    976.9, 977, 977.7, 978.3, 978.9, 979.8, 980.4, 981.2, 982.1, 983.1, 
    983.9, 984.9, 985.6, 986.6, 987.7, 988.5, 989.4, 990.3, 991, 991.6, 
    992.4, 992.9, 993.6, 994.6, 995.4, 996.4, 997.4, 998.1, 998.6, 999.3, 
    1000.1, 1001.1, 1001.8, 1002.5, 1003, 1003.8, 1004.5, 1005, 1005.7, 
    1006.2, 1006.7, 1007, 1007.4, 1007.7, 1007.7, 1008, 1008.1, 1008.4, 
    1008.6, 1008.9, 1009.1, 1009.3, 1009.4, 1009.4, 1009.3, 1009.2, 1009.3, 
    1009.4, 1009.5, 1009.7, 1009.8, 1010.3, 1010.5, 1010.8, 1011.3, 1011.9, 
    1012.4, 1012.8, 1013.2, 1013.6, 1014.4, 1015.2, 1015.7, 1016, 1016.5, 
    1017.1, 1017.9, 1018.4, 1018.9, 1019.3, 1019.8, 1020.2, 1020.4, 1020.4, 
    1020.9, 1021, 1021.4, 1021.5, 1021.4, 1021.2, 1020.7, 1020.2, 1019.8, 
    1019.6, 1019.3, 1019.3, 1019.2, 1019.1, 1018.9, 1019, 1018.8, 1018.7, 
    1018.4, 1018.3, 1018.2, 1018.2, 1017.7, 1017.5, 1016.9, 1016.1, 1015.7, 
    1014.8, 1014.1, 1013.3, 1012.6, 1012.1, 1011.4, 1010.5, 1009.4, 1008.7, 
    1008.3, 1008.3, 1008.3, 1008.3, 1008.3, 1008.2, 1008.3, 1008.9, 1009.1, 
    1009.3, 1009.2, 1009, 1009.2, 1008.5, 1008.4, 1008.4, 1008.4, 1008.1, 
    1007.8, 1007.4, 1007, 1006.7, 1006.6, 1006.9, 1007.1, 1007.2, 1007.4, 
    1007, 1006.7, 1006.4, 1005.9, 1005.1, 1004.4, 1003.1, 1002.4, 1001, 
    1000.4, 999.1, 997.1, 995.7, 994.8, 993.4, 991.9, 990.8, 989.7, 988.5, 
    987.2, 986.6, 985.8, 985.2, 984.8, 984.5, 984, 983.9, 983.9, 984, 983.8, 
    983.9, 983.9, 983.9, 984.1, 984.4, 984.5, 984.6, 984.6, 984.8, 985.3, 
    985.7, 985.6, 985.6, 985.6, 986, 986.4, 986.9, 986.9, 987.2, 987.7, 
    988.3, 988.5, 988.8, 989.3, 990, 990.4, 991.2, 991.9, 992.5, 993.1, 
    993.9, 994.4, 994.9, 995.3, 995.8, 995.9, 996.2, 996.5, 996.7, 997, 
    997.4, 997.7, 997.6, 997.4, 997.4, 997.2, 997.4, 997.4, 997.2, 996.8, 
    996.7, 996.6, 996.5, 996.2, 996.3, 996.3, 996.5, 996.5, 996.5, 996.8, 
    996.9, 997, 997.5, 998, 998.5, 998.8, 999.3, 999.8, 1000.7, 1001.1, 
    1001.8, 1002.1, 1002.5, 1003.1, 1003.8, 1004.3, 1004.8, 1005.4, 1006.1, 
    1006.8, 1007.4, 1008.1, 1008.4, 1008.8, 1009.5, 1010, 1010.7, 1011.2, 
    1011.8, 1012.4, 1012.9, 1013.6, 1013.7, 1014.5, 1015.1, 1015.5, 1015.8, 
    1016.1, 1016.3, 1016.8, 1017.1, 1017.2, 1017.7, 1018.1, 1018.2, 1018, 
    1018.3, 1018.5, 1018.5, 1018.4, 1018.4, 1018.3, 1018.4, 1018.1, 1017.9, 
    1017.8, 1017.8, 1017.1, 1017, 1016.5, 1016.1, 1015.7, 1015.5, 1015.3, 
    1015.1, 1014.7, 1014.6, 1014.4, 1013.8, 1013.3, 1012.6, 1012.2, 1011.6, 
    1011.1, 1010.9, 1010.9, 1010.7, 1010.4, 1009.7, 1009.3, 1009.2, 1008.7, 
    1008.3, 1007.6, 1007, 1006.5, 1006.1, 1005.6, 1004.9, 1005.1, 1004.7, 
    1003.7, 1002.8, 1001.6, 1000.8, 1000.1, 999.2, 998.5, 997.8, 997, 996.2, 
    995.3, 994.4, 993.6, 993.1, 992.4, 991.9, 991.6, 991.2, 990.8, 990.9, 
    990.8, 990.9, 990.8, 990.6, 990.5, 990.4, 990.8, 990.7, 990.4, 990.3, 
    990.2, 990.5, 990.9, 991.1, 991.7, 992.3, 992.5, 992.5, 992.7, 992.9, 
    993.2, 993.5, 993.4, 993.5, 993.9, 994.1, 994.4, 994.2, 993.9, 993.6, 
    993.5, 993.3, 993, 993, 992.9, 992.8, 992.9, 993, 993.2, 992.7, 993.2, 
    992.9, 992.3, 992.9, 992.7, 991.9, 991.8, 991.5, 992.1, 992.6, 992.8, 
    993.1, 993.6, 994.6, 994.8, 995.2, 995.7, 996.1, 997.2, 998, 998.8, 
    999.4, 1000.4, 1001.1, 1001.3, 1002.1, 1002.6, 1003.2, 1003.8, 1004.6, 
    1005.1, 1005.6, 1006.2, 1006.9, 1007.6, 1008.1, 1008.5, 1008.9, 1009.2, 
    1009.9, 1010.4, 1010.8, 1011.4, 1011.8, 1012.5, 1013.5, 1014, 1014.8, 
    1015.5, 1015.9, 1016.4, 1017, 1017.4, 1017.7, 1018.5, 1018.9, 1019.5, 
    1020.1, 1020.5, 1020.8, 1021, 1021.3, 1021.9, 1022.1, 1022.2, 1022.2, 
    1022.4, 1022.2, 1022.3, 1022.5, 1022.3, 1022.5, 1022.4, 1021.9, 1021.5, 
    1021.2, 1020.7, 1020.6, 1020.3, 1020.1, 1019.8, 1019.6, 1019.1, 1018.8, 
    1018.5, 1018.2, 1017, 1016.1, 1015.5, 1015.1, 1013.9, 1013.7, 1013.2, 
    1012.7, 1012.3, 1011.7, 1011.3, 1010.7, 1010.3, 1009.8, 1009.1, 1008.5, 
    1007.3, 1006.5, 1006, 1005.3, 1004.2, 1003.7, 1002.6, 1001.5, 1000.6, 
    999.2, 997.9, 996.3, 995, 994.2, 993.3, 992.4, 991.8, 991.3, 990.8, 
    990.3, 990, 990.1, 990.3, 990.3, 990.2, 990.2, 990.1, 990.1, 990.2, 
    990.5, 990.2, 990.2, 990.1, 990.2, 990, 990.2, 990.1, 990.5, 990.7, 
    990.7, 990.5, 990.7, 990.7, 990.4, 990.2, 990, 989.9, 989.9, 990, 989.9, 
    990.1, 990.3, 990.5, 990.8, 991, 991, 991.3, 991.4, 991.4, 991.5, 991.5, 
    991.8, 992.1, 992.3, 992.4, 992.4, 992.3, 992.3, 992.4, 992.6, 992.8, 
    993, 993.3, 993.9, 994.3, 994.9, 995.4, 996, 996.3, 996.5, 996.9, 997.3, 
    997.4, 997.8, 998.4, 998.7, 999.2, 999.6, 1000.3, 1000.5, 1000.6, 1001, 
    1001.2, 1001.6, 1001.7, 1001.7, 1001.9, 1002, 1001.9, 1002.2, 1002.1, 
    1001.8, 1001.8, 1001.6, 1001.6, 1001.4, 1001.3, 1001, 1000.9, 1000.9, 
    1000.9, 1000.7, 1000.7, 1000.3, 999.9, 999.4, 999, 998.5, 998, 997.4, 
    997.1, 996.8, 996.4, 996.1, 996.1, 995.7, 995.4, 995.2, 995.3, 995.2, 
    995.1, 994.8, 994.6, 994.8, 994.5, 994.6, 994.6, 994.6, 994.6, 994.7, 
    994.7, 995, 994.9, 995.1, 995.1, 995.4, 995.6, 996, 996.3, 996.5, 996.7, 
    996.8, 996.9, 997.1, 997.3, 997.5, 998.1, 998.5, 998.9, 999.3, 999.6, 
    999.7, 999.6, 999.9, 1000, 1000.2, 1000.6, 1000.3, 1000.5, 1000, 999.9, 
    999.9, 999.6, 999.2, 998.5, 997.6, 996.9, 995.7, 994, 992.9, 991.9, 
    990.9, 989.9, 988.7, 987.8, 987.8, 987.6, 987.9, 988.7, 989.5, 990.4, 
    991, 991.6, 992.1, 992.3, 992.2, 992, 991.9, 992, 992, 991.9, 992.1, 
    992.5, 992.7, 992.7, 993.4, 993.9, 994.3, 994.7, 994.7, 995.1, 995.2, 
    995.4, 995.6, 995.7, 996.4, 996.5, 996.6, 996.5, 997.2, 997.3, 997.9, 
    997.9, 998, 998.1, 998.1, 998.6, 998.6, 998.6, 999.3, 999.1, 999, 999.3, 
    999.3, 999.3, 999, 999.5, 999.5, 999.2, 998.7, 998.6, 998.4, 998.7, 
    998.8, 999, 999, 999, 999, 998.5, 998.6, 998.5, 998.2, 998.2, 998.2, 998, 
    998, 998.2, 998, 997.8, 997.3, 997.4, 997.1, 996.8, 996.6, 996.3, 996.1, 
    995.8, 995.6, 995.3, 994.8, 994.3, 994, 993.5, 993.1, 992.6, 992.2, 
    991.7, 991.2, 990.9, 990.1, 989.8, 989.4, 988.9, 988.5, 988.1, 987.7, 
    987.3, 986.5, 985.8, 985.5, 985.3, 985, 985.3, 984.8, 984.6, 984.3, 984, 
    983.8, 984, 983.9, 983.9, 984.6, 984.6, 984.8, 985, 985.1, 985.6, 985.9, 
    986.4, 986.8, 987.4, 987.9, 988.4, 988.6, 989, 989.4, 989.3, 989.6, 
    989.6, 990, 990.1, 990.7, 990.6, 990.7, 990.8, 990.9, 991.5, 991.9, 
    992.2, 992.4, 992.5, 992.5, 992.3, 992.4, 992.4, 992.4, 992.1, 991.9, 
    991.9, 991.8, 991.9, 991.6, 991.2, 990.9, 990.5, 990.1, 989.6, 989.3, 
    988.9, 989, 989.7, 989, 989.9, 989.8, 990, 990.1, 989.8, 990.1, 990.2, 
    990.4, 990.6, 990.4, 990.4, 990.6, 991, 991.3, 991.7, 991.8, 991.9, 992, 
    992, 992, 992.4, 992.6, 992.9, 993.2, 993, 993, 992.8, 992.7, 992.9, 
    993.3, 993.8, 994.3, 994.8, 995.5, 995.7, 996.1, 996.3, 996.2, 996.2, 
    996.1, 996, 995.8, 996.1, 996.3, 996.5, 996.9, 997.5, 997.9, 998.3, 
    998.9, 999, 999.1, 999.6, 999.9, 1000.2, 1000.3, 1000.6, 1000.9, 1001.4, 
    1001.5, 1001.8, 1002, 1002.3, 1002.5, 1002.5, 1002.6, 1002.6, 1002.7, 
    1002.6, 1002.7, 1002.8, 1002.8, 1002.6, 1002.3, 1002.1, 1001.6, 1001, 
    1000.6, 1000.2, 999.8, 999.2, 998.5, 997.8, 997.1, 996.4, 995.7, 995.1, 
    994.6, 994.1, 993.2, 992.4, 991.7, 991, 990.2, 989.7, 989.1, 988.4, 
    987.7, 987.3, 986.7, 986.2, 986, 985.4, 985.1, 984.7, 984.4, 984.4, 
    984.2, 983.7, 983.4, 983, 982.9, 982.5, 982.5, 982.3, 981.8, 981.8, 
    981.5, 981.2, 981, 981.2, 981.1, 981.4, 981.2, 981.2, 981.1, 980.7, 
    980.9, 980.8, 980.6, 980.7, 980.6, 980.5, 980.3, 980.1, 979.8, 979.6, 
    979.2, 978.8, 978.4, 978.2, 977.7, 976.7, 975.8, 975.3, 975.1, 975.2, 
    975.9, 976.4, 976.6, 976.6, 977.2, 978.2, 979.1, 979.1, 979.8, 979.9, 
    980.3, 980.6, 980.9, 981.3, 981.7, 982.1, 982.2, 982.8, 983.3, 983.5, 
    983.8, 984.1, 983.9, 984, 984.2, 984.1, 984.7, 985, 985.5, 986.1, 986.8, 
    987.5, 987.8, 988.3, 988.9, 989.4, 989.9, 990.6, 991, 991.6, 992, 992.6, 
    993.5, 994.4, 995.1, 995.6, 996.4, 997, 997.7, 998.5, 999.2, 999.5, 
    1000.5, 1001.2, 1001.9, 1002.4, 1003.4, 1004.3, 1005.1, 1005.6, 1006.4, 
    1007, 1007.4, 1007.9, 1008.4, 1008.9, 1009.2, 1010, 1010.4, 1010.7, 
    1011.1, 1011.2, 1011.4, 1011.3, 1011.1, 1010.9, 1010.7, 1010.6, 1010.4, 
    1010.2, 1010, 1009.5, 1009.2, 1008.8, 1008.2, 1008, 1007.8, 1007.4, 1007, 
    1006.9, 1006.8, 1006.6, 1006.8, 1006.8, 1006.8, 1006.8, 1006.5, 1006.5, 
    1006.2, 1006.2, 1005.8, 1005.5, 1005.3, 1005.3, 1005.2, 1004.8, 1004.7, 
    1004.3, 1004.1, 1003.5, 1002.8, 1001.9, 1001, 1000, 999.1, 998.2, 997.3, 
    996.1, 994.9, 994.3, 993.2, 992.2, 992, 991.8, 991.9, 992, 991.7, 991.8, 
    992, 992.7, 993.1, 993.5, 993.5, 993.8, 993.9, 993.9, 994.1, 994.1, 
    994.6, 994.8, 995.1, 995.6, 995.8, 995.4, 996, 996.2, 996.4, 996.7, 
    996.6, 996.6, 997.1, 997.4, 997.6, 998, 998.3, 998.1, 998.4, 998.8, 
    998.8, 998.8, 998.9, 999.2, 999.2, 999.6, 1000.1, 1000.4, 1000.7, 1000.7, 
    1000.9, 1001, 1001.2, 1001, 1000.7, 1001, 1001.2, 1001.2, 1001.1, 1001.2, 
    1001.2, 1001.2, 1001, 1000.8, 1000.8, 1000.5, 1000.4, 1000.2, 1000.3, 
    1000.6, 1000.7, 1000.7, 1000.7, 1000.7, 1000.5, 1000.7, 1000.7, 1000.6, 
    1000.4, 1000.3, 1000.2, 1000.3, 1000.3, 1000.1, 999.9, 999.7, 999.6, 
    999.7, 999.6, 999.5, 999.4, 999.3, 999.3, 999.1, 999.1, 998.8, 998.8, 
    998.7, 998.3, 998.4, 998.5, 998.5, 998.7, 999, 999.1, 999.5, 1000.1, 
    1000.5, 1000.9, 1000.9, 1001.4, 1001.9, 1002.6, 1003.2, 1003.7, 1004, 
    1004.4, 1005, 1005.3, 1005.3, 1005.5, 1005.4, 1006, 1006.3, 1006.7, 
    1007.3, 1007.8, 1008.5, 1009.1, 1009.7, 1010.4, 1011.2, 1012.6, 1012.8, 
    1013.6, 1013.9, 1014.9, 1015.5, 1016, 1016.6, 1017.1, 1017.6, 1018.2, 
    1018.7, 1019, 1019.3, 1019.6, 1020.2, 1020.2, 1020.4, 1020.5, 1020.5, 
    1020.7, 1020.8, 1021.1, 1021.1, 1021.2, 1021.1, 1021, 1020.9, 1020.5, 
    1020.4, 1020.2, 1019.8, 1019.5, 1019.6, 1019.4, 1019, 1018.4, 1017.6, 
    1017.3, 1016.5, 1015.9, 1015.4, 1014.2, 1013.5, 1012.3, 1011.6, 1011, 
    1010.1, 1009.2, 1007.9, 1006.9, 1005.8, 1004.1, 1002.9, 1001.6, 1000.6, 
    999.3, 998.4, 997, 996.4, 995.1, 993.2, 991.7, 990.2, 988.7, 987.2, 
    985.6, 984.3, 983.1, 982.4, 981.5, 980, 978.9, 977.8, 977.3, 976.2, 
    975.1, 974.8, 974.6, 973.8, 973.2, 971.8, 970.6, 972.5, 972.8, 973.6, 
    974.3, 974.1, 973.7, 973.3, 972.7, 973.2, 972.8, 972.1, 972.3, 971.8, 
    971.8, 971.8, 972.4, 972.1, 971.5, 971.3, 971.1, 970.5, 970.3, 970.7, 
    970.9, 970.9, 970.7, 970.6, 970.7, 970.7, 970.4, 970.2, 970.2, 969.6, 
    969.8, 969.8, 969.5, 969.3, 968.9, 968.9, 968.8, 968.7, 968.5, 968.3, 
    968.2, 968.2, 968.4, 968.6, 968.8, 968.9, 969.1, 969.2, 969.3, 969.6, 
    969.9, 970.2, 970.5, 970.9, 971.5, 972.1, 972.9, 973.5, 974, 974.7, 
    975.4, 976.2, 976.9, 977.8, 978.8, 980, 981.2, 982.5, 983.5, 984.5, 
    985.3, 986.4, 987.1, 987.7, 988.3, 988.4, 989.1, 989.6, 990.1, 990.7, 
    991, 991.1, 991.2, 991.5, 992.1, 992, 991.9, 991.5, 991.1, 991, 990.9, 
    990.3, 990.1, 989.6, 989.1, 988.6, 988, 987.3, 986.2, 985.4, 984.7, 
    983.8, 983.6, 983.7, 983.7, 983.4, 983.2, 983, 982.8, 982.3, 982, 981.6, 
    981, 980.5, 980.2, 980.1, 979.8, 979.5, 979.1, 978.8, 978.6, 978.5, 978, 
    977.6, 977.3, 977, 976.6, 976.4, 976.1, 975.7, 975.3, 975.6, 975.6, 
    975.6, 975.6, 975.7, 975.6, 975.7, 976.1, 976.4, 976.8, 977.3, 977.3, 
    977, 977, 977.2, 977.6, 978.1, 978.4, 978.5, 979.2, 979.4, 980.2, 980.7, 
    981.1, 981.7, 982.4, 983.2, 983.8, 984.1, 984.4, 985.1, 985.6, 986, 
    986.8, 987.2, 988, 988.7, 989, 989.2, 989.6, 989.8, 990.4, 991.1, 991.6, 
    992.3, 993, 993.8, 994.7, 995.3, 996, 996.8, 997.6, 998.5, 999.2, 999.9, 
    1000.4, 1001.3, 1002, 1002.8, 1003.8, 1004.6, 1005.5, 1006.4, 1006.6, 
    1007.2, 1007.7, 1007.8, 1008.1, 1008.1, 1006.7, 1005.2, 1004.8, 1004.4, 
    1004.1, 1004, 1004.3, 1004.4, 1004.8, 1005.2, 1006.2, 1007.3, 1008.6, 
    1009.7, 1010.3, 1011.8, 1012.7, 1013.7, 1014.6, 1014.8, 1014.7, 1015.1, 
    1015.3, 1015.5, 1016.2, 1016.3, 1016.2, 1016.4, 1016.4, 1015.9, 1015.5, 
    1014.9, 1014.3, 1013.7, 1013.6, 1013.6, 1012.8, 1012.3, 1011.9, 1011.4, 
    1010.7, 1009.8, 1008.4, 1007.5, 1007.2, 1006.2, 1005.4, 1004.8, 1004.1, 
    1003.7, 1003.4, 1002.5, 1001.4, 1000.3, 999.5, 998.4, 997.1, 996.8, 997, 
    997.1, 997.4, 997.7, 999, 999.9, 1000.9, 1001.5, 1002.3, 1002.4, 1002.8, 
    1002.8, 1002.4, 1002.8, 1002.6, 1002.7, 1002.6, 1002.5, 1001.4, 1000.5, 
    999.4, 998.2, 996.6, 996.2, 994.6, 994.8, 994.9, 995.7, 996, 996.4, 
    996.7, 996.9, 997, 997.9, 998.9, 1000.1, 1001.2, 1002.3, 1003.5, 1004.7, 
    1005.8, 1006.8, 1007.6, 1008.1, 1008.9, 1008.4, 1008.4, 1008.4, 1008.4, 
    1008.3, 1008.1, 1007.3, 1006.8, 1006.2, 1005.1, 1003.9, 1003.2, 1002.8, 
    1003.3, 1003.1, 1003.4, 1004.3, 1004.6, 1005.7, 1006.7, 1007, 1007.3, 
    1007.6, 1007.2, 1006.7, 1006.1, 1006.2, 1005.3, 1003.9, 1003.5, 1003.3, 
    1003.3, 1003.6, 1005.1, 1006.7, 1008.5, 1010.4, 1012, 1013.9, 1015.6, 
    1017.1, 1018.9, 1020.6, 1021.4, 1021.3, 1020.9, 1020.2, 1020.1, 1018.9, 
    1018, 1017.4, 1016.9, 1015.8, 1015.3, 1014.6, 1014, 1013.2, 1012.5, 
    1012.3, 1011.6, 1012, 1013, 1012.9, 1013.4, 1013.5, 1013.7, 1014.1, 
    1014.4, 1014.1, 1014.4, 1014.3, 1014.1, 1014, 1014.2, 1014.5, 1014.7, 
    1015, 1015.3, 1015.2, 1015.3, 1015.6, 1016.1, 1016, 1016.3, 1016.8, 1017, 
    1017.3, 1017.8, 1018.2, 1018.8, 1019.2, 1019.6, 1020, 1020.5, 1020.9, 
    1021.1, 1021.4, 1021.7, 1022.1, 1022.2, 1022.5, 1022.7, 1022.7, 1022.7, 
    1022.4, 1022.4, 1022.5, 1022.5, 1022.3, 1022.1, 1022, 1021.9, 1021.7, 
    1021.5, 1021.3, 1020.9, 1020.8, 1020.5, 1020.3, 1020.3, 1019.9, 1019.4, 
    1019.3, 1019.3, 1019.5, 1019.4, 1019.3, 1019.2, 1019.1, 1019, 1019, 
    1019.2, 1019.4, 1019.5, 1019.8, 1020, 1020.3, 1020.5, 1020.6, 1020.8, 
    1020.9, 1021.1, 1021.3, 1021.4, 1021.5, 1021.7, 1022.1, 1022.3, 1022.7, 
    1023, 1023.2, 1023.3, 1023.2, 1023.4, 1023.4, 1023.3, 1023.4, 1023.3, 
    1023.3, 1023.4, 1023.4, 1022.9, 1022.6, 1022.4, 1022, 1021.9, 1021.4, 
    1021, 1020.6, 1020, 1019.7, 1019.5, 1019.5, 1019.6, 1019.4, 1019.3, 
    1019.3, 1019.3, 1019.4, 1019.4, 1019.5, 1019.5, 1019.7, 1020, 1020.2, 
    1020.4, 1020.5, 1020.7, 1020.7, 1020.9, 1021, 1021.2, 1021.3, 1021.5, 
    1021.5, 1021.7, 1021.9, 1021.9, 1021.8, 1021.8, 1021.9, 1021.9, 1021.7, 
    1021.8, 1021.7, 1021.7, 1021.7, 1021.7, 1021.9, 1022, 1022, 1021.9, 
    1021.9, 1022.1, 1022.1, 1022, 1021.8, 1021.7, 1021.9, 1022.2, 1022.5, 
    1022.8, 1022.8, 1022.7, 1022.9, 1022.8, 1022.7, 1022.6, 1022.9, 1023, 
    1023.2, 1023.4, 1023.9, 1024.3, 1024.5, 1024.8, 1024.9, 1024.9, 1025.2, 
    1025.4, 1025.6, 1025.9, 1026.3, 1026.9, 1027.5, 1027.9, 1028.3, 1028.7, 
    1029.2, 1029.6, 1029.9, 1030.2, 1030.5, 1030.9, 1031.3, 1031.7, 1032.3, 
    1032.5, 1032.7, 1033, 1033, 1033.3, 1033.5, 1033.8, 1033.8, 1033.7, 
    1033.8, 1034, 1034.2, 1034.1, 1034.2, 1034, 1033.8, 1033.7, 1033.4, 1033, 
    1032.5, 1032.4, 1031.7, 1031.3, 1030.9, 1030.3, 1029.8, 1029.1, 1028.3, 
    1027.6, 1026.9, 1026.1, 1025.5, 1024.7, 1024, 1023.7, 1023.4, 1023.3, 
    1022.9, 1022.5, 1022, 1021.5, 1020.9, 1020.5, 1020.2, 1019.8, 1019.2, 
    1018.6, 1018.1, 1017.6, 1016.8, 1015.9, 1015.4, 1014.5, 1013.8, 1012.8, 
    1011.7, 1010.5, 1009.7, 1009.3, 1009.1, 1009.4, 1009.3, 1008.9, 1008.5, 
    1008.6, 1008.7, 1008.9, 1009.1, 1009.4, 1009.5, 1009.9, 1010.3, 1010.7, 
    1011.4, 1011.6, 1011.9, 1012.1, 1012.5, 1013, 1013, 1013.2, 1013.5, 
    1013.6, 1014, 1014.4, 1014.7, 1014.8, 1014.6, 1014.6, 1014.9, 1015.1, 
    1015, 1015, 1015.2, 1015, 1015.2, 1015.2, 1015.3, 1015.4, 1015.3, 1015.3, 
    1015.2, 1015.2, 1015.2, 1015.1, 1015.1, 1015.3, 1015.9, 1016.5, 1016.6, 
    1016.6, 1017, 1017.3, 1017.1, 1017.4, 1017.2, 1017.2, 1017.3, 1017.3, 
    1017.7, 1018.1, 1018.6, 1019, 1019.2, 1019.1, 1019.1, 1019.1, 1019.3, 
    1019.2, 1019.2, 1018.7, 1018.7, 1018.8, 1018.6, 1018.7, 1018.2, 1017.9, 
    1017.6, 1017.2, 1017, 1016.6, 1016.1, 1015.9, 1015.7, 1015.3, 1014.7, 
    1014.2, 1013.5, 1013.2, 1012.6, 1012.1, 1011.8, 1011.7, 1011.7, 1011.3, 
    1011.2, 1011.2, 1011.3, 1011.1, 1011.5, 1011.6, 1011.7, 1011.8, 1011.8, 
    1012, 1011.8, 1011.7, 1011.8, 1011.8, 1011.8, 1011.7, 1011.7, 1011.5, 
    1011.4, 1011.4, 1011.1, 1010.9, 1011, 1010.8, 1010.7, 1010.7, 1010.6, 
    1010.5, 1010.2, 1010.2, 1009.9, 1009.7, 1009.5, 1009.2, 1009.1, 1008.8, 
    1008.7, 1008.5, 1008, 1007.8, 1007.6, 1007.4, 1007.1, 1006.8, 1006.5, 
    1006.5, 1006.4, 1006.2, 1006.2, 1006.5, 1006.5, 1006.3, 1006, 1005.8, 
    1005.9, 1006.3, 1006.5, 1006.5, 1006.5, 1006.9, 1007.2, 1007.2, 1007.4, 
    1007.5, 1007.6, 1007.6, 1007.7, 1007.6, 1007.3, 1007, 1007, 1006.9, 
    1006.8, 1006.7, 1006.1, 1005.5, 1004.5, 1004.3, 1004.1, 1003.8, 1003, 
    1002.7, 1002.3, 1001.9, 1001.6, 1001.3, 1000.8, 1000.3, 1000.2, 999.7, 
    999.7, 999.6, 999.4, 999.3, 999.4, 999.5, 1000.1, 1000.4, 1000.5, 1000.7, 
    1000.8, 1001, 1001.2, 1001.2, 1001, 1000.9, 1000.8, 1001, 1001.1, 1000.9, 
    1001, 1001.2, 1001.3, 1001.6, 1001.9, 1002.5, 1002.7, 1003.1, 1003.7, 
    1003.9, 1004.8, 1005.6, 1006, 1006.5, 1006.8, 1006.9, 1007.4, 1007.6, 
    1008.1, 1008.5, 1008.5, 1009, 1008.8, 1009.4, 1009.4, 1009.4, 1009.5, 
    1009.6, 1009.5, 1009.7, 1009.2, 1008.9, 1008.7, 1008.6, 1008.6, 1008.6, 
    1008.5, 1008.6, 1008.8, 1008.6, 1008.5, 1008.6, 1008.7, 1008.6, 1008.5, 
    1008.7, 1009.1, 1009, 1009.2, 1009.5, 1009.6, 1009.9, 1010, 1009.9, 
    1009.8, 1009.7, 1009.8, 1009.9, 1010.4, 1010.9, 1011.4, 1011.5, 1011.7, 
    1011.9, 1012.3, 1012.6, 1012.7, 1013, 1012.7, 1012.7, 1012.8, 1012.7, 
    1012.4, 1011.9, 1011.2, 1010.6, 1010, 1009.1, 1008.6, 1007.9, 1007, 
    1006.3, 1006.1, 1005.4, 1004.8, 1004.4, 1004.1, 1003.5, 1002.8, 1002.1, 
    1001.3, 1000.6, 999.8, 999.5, 998.8, 998.3, 997.6, 996.9, 996.2, 995.5, 
    995, 994.4, 993.6, 993.1, 992.5, 991.9, 991.6, 991.5, 991.1, 990.7, 
    990.5, 990.2, 989.5, 989.2, 988.9, 988.6, 988.1, 987.8, 987.8, 987.5, 
    987.3, 987.2, 986.9, 986.8, 986.4, 986.1, 985.7, 985.2, 985, 984.7, 
    985.2, 984.7, 984.3, 983.8, 983.4, 983.2, 983.1, 983.2, 982.8, 982.9, 
    982.7, 982.3, 982.1, 981.8, 981.3, 980.9, 980.5, 980, 979.6, 979.2, 
    979.1, 979, 978.9, 979.1, 979.3, 979.5, 979.5, 979.5, 979.7, 979.4, 
    979.1, 979.2, 979.4, 979.3, 979.3, 979.5, 979.7, 979.6, 979.5, 979.8, 
    979.5, 979.6, 979.5, 979.9, 980.4, 980.9, 980.9, 981.3, 982.1, 982.8, 
    983.8, 984.2, 984.7, 985.2, 985.4, 986, 986.5, 987.4, 987.5, 987.9, 
    988.3, 988.6, 988.7, 989.1, 989.5, 989.5, 989.6, 990, 989.8, 989.5, 
    989.6, 989.7, 990.2, 990.5, 990.3, 990.4, 990.1, 989.7, 989.5, 989.7, 
    989.9, 990, 989.9, 990.2, 990.2, 990.4, 990.3, 990.8, 990.1, 990.9, 
    991.2, 991.2, 991.3, 991.8, 991.9, 992.2, 992.4, 992.8, 992.5, 993.1, 
    993, 993, 992.9, 992.9, 992.6, 992.9, 993, 993, 993.6, 994.2, 994, 994.5, 
    994.9, 994.6, 994.5, 994.7, 995.5, 995.2, 995.2, 995.5, 994.8, 995.1, 
    995.6, 996.4, 996.7, 997.2, 997.5, 998.3, 998.8, 998.6, 998.8, 999.1, 
    999.7, 1000, 1000.1, 1000.4, 1000.8, 1001.1, 1001.1, 1001.3, 1002, 
    1002.2, 1002.2, 1002.6, 1003.1, 1003.5, 1003.8, 1003.7, 1004.5, 1005.1, 
    1005.4, 1005.4, 1005.3, 1005.5, 1005.6, 1005.9, 1006.9, 1006.9, 1007.1, 
    1008.1, 1009, 1009.6, 1009.7, 1010.3, 1010.9, 1011.5, 1011.6, 1011.7, 
    1012.2, 1012.1, 1012.6, 1012.7, 1013.2, 1013.5, 1013.7, 1014, 1014.3, 
    1014.1, 1013.8, 1013.6, 1013.5, 1013.6, 1013.5, 1013.1, 1012.7, 1012.5, 
    1012.2, 1011.8, 1011.4, 1010.8, 1010.2, 1009.9, 1009.8, 1009.7, 1009.4, 
    1009, 1008.6, 1008.2, 1007.8, 1007.6, 1007.3, 1006.8, 1006.4, 1006.4, 
    1006.2, 1006, 1005.8, 1005.8, 1005.4, 1005.3, 1005.3, 1005.3, 1005.2, 
    1005, 1004.9, 1004.8, 1005.1, 1005.1, 1005.3, 1005.4, 1005.3, 1005, 
    1005.2, 1005, 1004.9, 1004.8, 1004.9, 1004.9, 1005.2, 1005.1, 1004.9, 
    1004.9, 1004.7, 1004.5, 1004.5, 1004.5, 1004.4, 1004.3, 1004.3, 1004.5, 
    1004.6, 1004.4, 1004.2, 1004.1, 1003.9, 1003.8, 1003.5, 1003.3, 1003.1, 
    1002.9, 1003, 1002.7, 1002.8, 1002.6, 1002.3, 1001.9, 1001.6, 1001.2, 
    1000.9, 1000.7, 1000.3, 1000.1, 999.7, 999.6, 999.5, 999.3, 999.1, 998.7, 
    998.1, 997.7, 997.4, 997.3, 997, 996.5, 996.2, 995.9, 995.6, 995.2, 
    994.2, 993.1, 992.5, 991.8, 990.9, 990.3, 989.5, 988.7, 988.9, 987.6, 
    987.7, 987.6, 987.7, 986.9, 986.8, 986.2, 985.8, 985.5, 985.2, 985.2, 
    984.9, 985.1, 985.1, 985.1, 985.2, 985.7, 985.9, 985.8, 986.1, 986.6, 
    986.6, 986.9, 987, 987.1, 987.4, 987.6, 988.2, 988.3, 988.4, 988.4, 
    988.7, 988.9, 989.1, 989.1, 989.2, 989.4, 989.6, 989.8, 990, 990.1, 
    990.2, 990.6, 990.9, 991.1, 991.2, 991.2, 991.4, 991.7, 992.2, 992.5, 
    992.7, 992.9, 993.1, 993.3, 993.4, 993.6, 993.9, 994.1, 994.3, 994.5, 
    994.8, 995, 995.4, 995.5, 996.2, 996.7, 997.1, 997.6, 997.9, 998.3, 999, 
    999.8, 1000.5, 1001.3, 1001.9, 1002.4, 1003, 1003.4, 1003.8, 1004.2, 
    1004.4, 1004.6, 1004.7, 1004.8, 1004.9, 1005.3, 1005.4, 1005.5, 1005.5, 
    1005.5, 1005.6, 1005.8, 1005.8, 1005.8, 1005.9, 1005.8, 1006.4, 1006.6, 
    1006.7, 1006.8, 1006.9, 1006.9, 1006.9, 1006.8, 1006.3, 1005.9, 1005.4, 
    1005, 1004.7, 1004.3, 1004.3, 1004.5, 1004.6, 1004.7, 1004.8, 1005.4, 
    1005.5, 1005.8, 1006.1, 1006.6, 1007.3, 1007.8, 1008.3, 1008.5, 1008.5, 
    1008.7, 1009, 1009, 1009.1, 1009, 1009, 1009.1, 1009.3, 1009.7, 1009, 
    1009.1, 1008.4, 1007.7, 1007, 1007, 1006.7, 1006.3, 1006, 1005.8, 1005.6, 
    1005.6, 1005.8, 1006.1, 1006.4, 1006.6, 1006.9, 1007.1, 1007.4, 1007.4, 
    1007.4, 1007.7, 1007.9, 1007.8, 1007.5, 1007.3, 1007.1, 1006.9, 1006.8, 
    1006.6, 1006.5, 1006.2, 1006.1, 1006.1, 1006.2, 1006.3, 1006.3, 1006.5, 
    1006.7, 1006.8, 1006.7, 1006.8, 1006.9, 1007, 1007, 1007.3, 1007.6, 
    1007.5, 1007.8, 1008, 1007.9, 1007.9, 1007.7, 1007.3, 1006.7, 1006.4, 
    1006, 1005.7, 1005.4, 1004.8, 1004.5, 1004.4, 1003.7, 1002.9, 1002.4, 
    1002.3, 1001.8, 1001.2, 1000.8, 1000.6, 1000.5, 1000.6, 1000.8, 1000.8, 
    1000.9, 1000.9, 1001.4, 1001.5, 1001.7, 1001.9, 1002.2, 1002.7, 1003.2, 
    1003.5, 1003.8, 1004.1, 1004.1, 1003.9, 1003.6, 1003.1, 1002.8, 1002.3, 
    1001.7, 1001.7, 1001.7, 1001.5, 1001, 1000.4, 999.6, 998.8, 998.2, 997.4, 
    996.6, 995.8, 995.6, 995.3, 995.2, 994.8, 994.4, 994, 993.5, 992.7, 
    992.3, 991.8, 991.8, 991.3, 990.9, 990.6, 990.5, 990.5, 990.2, 989.9, 
    989.8, 989.7, 989.5, 989.3, 989.2, 988.8, 989.1, 989.6, 989.8, 990.3, 
    990.8, 991.4, 991.5, 991.7, 992.1, 992.5, 993.1, 993.6, 994.2, 994.8, 
    995.4, 996.3, 996.9, 997.5, 998, 998.4, 998.8, 999.4, 999.7, 1000.2, 
    1000.3, 1000.5, 1000.9, 1001.1, 1001.2, 1001.4, 1001.6, 1001.3, 1001.3, 
    1001.1, 1000.9, 1000.4, 1000, 999.9, 999.3, 998.9, 998.8, 998.4, 998.3, 
    997.8, 997.2, 996.6, 996.8, 996.9, 997.1, 997.1, 996.9, 997.3, 997.5, 
    998, 998.3, 998.3, 998.5, 999.3, 999.7, 1000.2, 1000.8, 1001.5, 1001.9, 
    1002.4, 1003, 1003.5, 1003.8, 1004.3, 1004.7, 1005.2, 1005.6, 1005.9, 
    1006.1, 1006.3, 1006.7, 1007.2, 1007.1, 1007.1, 1007.1, 1006.5, 1006.5, 
    1006.7, 1007.3, 1007.4, 1007.8, 1008.2, 1008.4, 1008.9, 1009.4, 1009.9, 
    1010.5, 1011.2, 1011.9, 1012.4, 1012.9, 1013.3, 1013.5, 1013.9, 1014.4, 
    1014.9, 1015.3, 1015.4, 1015.2, 1015.5, 1015.8, 1016, 1016, 1015.8, 
    1015.8, 1017.1, 1015.8, 1015.9, 1015.9, 1015.8, 1015.8, 1015.6, 1015.4, 
    1015.5, 1015.2, 1014.8, 1014.7, 1015, 1014.9, 1014.7, 1014.8, 1014.6, 
    1014.3, 1014, 1014, 1013.8, 1013.8, 1014, 1014, 1014, 1014.2, 1014.3, 
    1014.1, 1014, 1014, 1013.8, 1013.9, 1014, 1013.9, 1014, 1014.1, 1014.5, 
    1014.3, 1014.4, 1014.8, 1015, 1015.1, 1014.9, 1014.6, 1014.7, 1014.8, 
    1014.7, 1014.8, 1015, 1015, 1014.8, 1014.5, 1014.3, 1014, 1013.5, 1013.1, 
    1012.9, 1012.8, 1012.4, 1012.1, 1011.8, 1011.8, 1011.7, 1011.3, 1010.9, 
    1010.6, 1010.4, 1010.2, 1010, 1009.6, 1009.1, 1008.9, 1008.8, 1008.4, 
    1008.3, 1008.1, 1007.8, 1007.6, 1007.4, 1007.3, 1007.2, 1007.1, 1007, 
    1007, 1006.9, 1007, 1007.1, 1007.1, 1007, 1007, 1006.8, 1006.7, 1006.6, 
    1006.6, 1006.4, 1006.4, 1006.3, 1006.3, 1006.3, 1006.3, 1005.9, 1005.8, 
    1005.5, 1005.3, 1005.2, 1005, 1004.7, 1004.6, 1004.4, 1004.5, 1004.4, 
    1004.5, 1004.4, 1004.5, 1004.5, 1004.4, 1004.3, 1004.3, 1004.1, 1003.9, 
    1003.7, 1003.2, 1002.9, 1002.7, 1002.3, 1002.2, 1001.8, 1001.5, 1001.5, 
    1001.1, 1001.1, 1000.9, 1000.7, 1000.7, 1000.9, 1001.2, 1001.2, 1001.5, 
    1001.6, 1001.6, 1001.5, 1001.6, 1001.8, 1001.5, 1001.2, 1000.8, 1000.4, 
    999.9, 999.4, 998.7, 997.9, 996.9, 995.8, 995, 994.7, 993.9, 993.6, 
    993.4, 993.6, 994.3, 994.8, 995.2, 995, 994.9, 995.3, 995.2, 995.5, 
    995.8, 996, 996.4, 996.6, 997.2, 997.8, 998.2, 998.5, 998.6, 998.6, 
    998.6, 998.6, 998.7, 998.6, 998.9, 999.2, 999.5, 999.7, 1000, 999.9, 
    999.9, 999.9, 1000, 1000, 1000.1, 1000.3, 1000.7, 1000.8, 1001, 1001.3, 
    1001.3, 1001.2, 1001.6, 1001.7, 1001.8, 1002, 1002.3, 1002.4, 1002.3, 
    1002.7, 1002.9, 1002.9, 1003.1, 1002.9, 1002.7, 1002.7, 1002.6, 1002.7, 
    1002.4, 1002.1, 1002.1, 1002.1, 1002.2, 1002.2, 1002.1, 1001.9, 1001.7, 
    1001.5, 1001.4, 1001.4, 1001.1, 1001.3, 1000.8, 1000.9, 1000.8, 1000.8, 
    1000.8, 1001.1, 1001.7, 1002.1, 1002.3, 1002.8, 1003.2, 1003.8, 1004.2, 
    1004.6, 1004.9, 1004.8, 1004.9, 1005.1, 1005, 1005.2, 1005.2, 1005.4, 
    1005.6, 1005.7, 1006, 1006.1, 1006.6, 1006.6, 1006.8, 1007.1, 1007.2, 
    1007.5, 1007.8, 1008, 1008.3, 1008.6, 1009, 1009.4, 1009.7, 1010.1, 
    1010.3, 1010.4, 1010.4, 1010.5, 1010.4, 1010.7, 1010.7, 1010.7, 1010.9, 
    1011, 1011.4, 1011.3, 1011, 1011, 1011, 1010.8, 1010.8, 1010.8, 1010.8, 
    1010.9, 1010.8, 1010.8, 1011, 1011, 1011, 1011, 1011.2, 1011.4, 1011.6, 
    1011.8, 1012.1, 1012.3, 1012.5, 1012.8, 1013.1, 1013.3, 1013.4, 1013.5, 
    1013.6, 1014, 1014, 1014.4, 1014.6, 1014.8, 1015.1, 1015.3, 1015.5, 
    1015.8, 1015.9, 1015.7, 1015.7, 1015.7, 1015.7, 1015.6, 1015.6, 1015.5, 
    1015.7, 1015.8, 1015.7, 1015.8, 1015.5, 1015.3, 1015.2, 1015, 1015.1, 
    1015.1, 1015.1, 1014.8, 1014.6, 1014.3, 1014.1, 1014, 1014, 1014, 1014.1, 
    1014, 1014, 1013.8, 1014.1, 1013.9, 1014, 1014.1, 1014.3, 1014.5, 1014.7, 
    1014.6, 1014.6, 1014.7, 1014.5, 1014.3, 1014.4, 1014.3, 1014, 1013.7, 
    1013.4, 1013.1, 1012.9, 1013.1, 1013, 1012.6, 1012.3, 1011.8, 1011.5, 
    1011.4, 1011.1, 1010.8, 1010.4, 1010.6, 1009.9, 1009.4, 1008.6, 1007.5, 
    1006.9, 1006.1, 1005.1, 1004.1, 1003.7, 1003.2, 1003, 1002.8, 1003.5, 
    1003.8, 1004.1, 1004.3, 1004.8, 1005.1, 1005.4, 1005.1, 1005, 1005.2, 
    1005.2, 1005.2, 1005.3, 1005, 1005.3, 1005, 1005, 1004.6, 1004.7, 1004.7, 
    1004.4, 1003.8, 1003.6, 1003.1, 1002.6, 1002.1, 1001.5, 1000.4, 999, 
    997.2, 995.4, 993.9, 992.4, 991.6, 992.1, 992.2, 992.3, 992.5, 992.2, 
    991.7, 991.7, 991.6, 991, 990.6, 991.1, 991.4, 993.3, 995.7, 997.3, 
    999.5, 1001.2, 1003.1, 1004.4, 1005.8, 1006.8, 1007.2, 1007.3, 1007.4, 
    1007, 1006.6, 1004.9, 1003.4, 1001.8, 999.3, 996.5, 993.8, 990.4, 987.4, 
    985, 982.6, 981, 979.7, 978.9, 978.7, 979, 979.6, 980.5, 981.7, 982.9, 
    984.6, 986.4, 988.4, 990.6, 992.5, 994.5, 996, 997.2, 998.5, 999.4, 
    1000.6, 1002, 1002.7, 1003.9, 1004.7, 1005.5, 1005.8, 1006.2, 1006.1, 
    1006.4, 1006.5, 1006.7, 1007.2, 1007.4, 1007.9, 1007.9, 1008.5, 1008.8, 
    1008.8, 1008.7, 1008.9, 1008.9, 1009.2, 1009.6, 1009.9, 1010.2, 1010.5, 
    1011.5, 1012.2, 1012.7, 1013.3, 1013.6, 1014.2, 1014.8, 1015, 1015.2, 
    1015.5, 1015.7, 1016.1, 1016.3, 1016.7, 1017.3, 1017.6, 1017.8, 1017.8, 
    1018, 1018.1, 1018, 1018.1, 1017.9, 1018.1, 1018.3, 1018.3, 1018.5, 
    1018.7, 1018.6, 1018.5, 1018.2, 1018.1, 1017.8, 1017.8, 1017.3, 1017, 
    1016.9, 1017, 1016.6, 1017.3, 1016.9, 1016.8, 1016.5, 1016.2, 1015.9, 
    1015.1, 1015.2, 1015.1, 1015.1, 1014.9, 1014.8, 1014.8, 1014.5, 1014.1, 
    1013.9, 1013.6, 1013.3, 1012.9, 1012.7, 1012.5, 1012.3, 1012.1, 1012.1, 
    1012, 1011.8, 1011.5, 1011.5, 1011.8, 1011.6, 1011.6, 1011.3, 1011.1, 
    1011.2, 1011.3, 1011.4, 1011.3, 1011.3, 1011.3, 1011.2, 1011.3, 1011.6, 
    1011.2, 1011.2, 1011.4, 1011.8, 1012, 1012.2, 1012.3, 1012.3, 1012.2, 
    1012.3, 1012.1, 1012.2, 1012, 1012, 1011.8, 1011.7, 1011.5, 1011.5, 
    1011.5, 1011.3, 1010.8, 1010.4, 1010.3, 1010.1, 1009.8, 1009.7, 1009.4, 
    1009.2, 1009.3, 1009.1, 1009, 1008.8, 1008.5, 1008.2, 1008, 1008, 1007.7, 
    1007.5, 1007.5, 1007.3, 1007.1, 1007.2, 1007, 1006.9, 1006.8, 1006.6, 
    1006.5, 1006.4, 1006.3, 1006.3, 1006.3, 1006.4, 1006.4, 1006.5, 1006.8, 
    1006.8, 1007, 1007.3, 1007.3, 1007.7, 1007.6, 1008, 1008.2, 1008.3, 
    1008.6, 1008.9, 1009, 1009.2, 1009.4, 1009.3, 1009.4, 1009.6, 1009.6, 
    1009.7, 1009.7, 1010, 1010.1, 1010.4, 1010.5, 1010.6, 1010.9, 1011, 
    1011.2, 1011, 1010.9, 1010.9, 1010.6, 1010.4, 1010.2, 1010, 1010.1, 
    1009.9, 1009.7, 1009.3, 1009.2, 1009, 1008.7, 1008.6, 1008.5, 1008.5, 
    1008.5, 1008.5, 1008.4, 1008.4, 1008.1, 1008, 1008, 1008, 1007.9, 1007.8, 
    1007.8, 1007.8, 1007.8, 1007.5, 1007.4, 1007.3, 1007.1, 1007.2, 1007, 
    1006.8, 1006.6, 1006.6, 1006.3, 1006, 1005.8, 1005.8, 1005.6, 1005.4, 
    1005.4, 1005.4, 1005.2, 1005.3, 1005.2, 1005.1, 1005.2, 1005.4, 1005.6, 
    1005.6, 1005.5, 1005.5, 1005.5, 1005.5, 1005.4, 1005.3, 1005.1, 1005, 
    1004.8, 1004.6, 1004.5, 1004.3, 1004.2, 1003.8, 1003.5, 1003.2, 1002.8, 
    1002.3, 1001.8, 1001.7, 1001.4, 1000.8, 1000.4, 999.8, 999.5, 998.7, 
    997.9, 997.5, 997.1, 996.4, 995.8, 995, 994.5, 993.8, 993.2, 992.6, 
    992.1, 990.9, 989.8, 989.1, 987.4, 986.2, 985, 984.1, 983.3, 982.6, 
    981.7, 981.2, 980.6, 979.8, 979.2, 978.3, 977.5, 976.8, 976.5, 975.9, 
    975.3, 974.9, 974.4, 973.8, 973.3, 973, 973.1, 973.1, 973, 973.4, 973.7, 
    974.1, 974.8, 975.7, 976.7, 977.8, 978.9, 980.1, 981.2, 982.2, 983.1, 
    983.7, 984.1, 984.8, 985.5, 986.4, 987.3, 987.8, 988.3, 988.7, 989.1, 
    989.5, 989.7, 989.8, 990.1, 990.3, 990.4, 990.8, 990.7, 991, 990.9, 991, 
    991.1, 991.3, 991.5, 991.5, 991.6, 991.9, 992.4, 992.3, 992.8, 992.9, 
    993, 993.1, 993.3, 993.3, 993.3, 993.4, 993.2, 993.2, 993.4, 993.4, 
    993.3, 993.6, 994, 994, 994.3, 994.5, 994.6, 995.1, 995.3, 995.8, 996.3, 
    996.6, 997, 997.5, 998.1, 998.7, 999, 999.7, 1000.1, 1000.9, 1001.2, 
    1001.5, 1002, 1002.5, 1003.1, 1003.8, 1004.3, 1005.1, 1005.7, 1006.2, 
    1006.5, 1006.8, 1007.3, 1007.8, 1008.2, 1008.7, 1009.3, 1009.8, 1010.2, 
    1010.6, 1010.8, 1011.4, 1011.6, 1011.8, 1012.4, 1012.8, 1013.2, 1013.4, 
    1014, 1014.2, 1014.2, 1014.4, 1014.8, 1014.8, 1015.1, 1015.2, 1015.3, 
    1015.3, 1015.5, 1015.7, 1015.8, 1016, 1016.2, 1016.3, 1016.5, 1016.4, 
    1016.5, 1016.7, 1016.8, 1016.9, 1016.9, 1016.9, 1017.1, 1017.2, 1017.2, 
    1017, 1017, 1016.9, 1016.9, 1017, 1017, 1017.1, 1017.3, 1017.5, 1017.5, 
    1017.7, 1017.7, 1017.6, 1017.4, 1017.3, 1017, 1017, 1017.1, 1017.1, 
    1017.4, 1017.4, 1017.5, 1017.7, 1017.8, 1017.8, 1017.6, 1017.6, 1017.5, 
    1017.3, 1017.4, 1017.4, 1017.4, 1017.7, 1018, 1018.3, 1018.2, 1018.4, 
    1018.5, 1018.5, 1018.6, 1018.6, 1018.7, 1018.7, 1018.9, 1019.1, 1019.1, 
    1019.1, 1019, 1018.7, 1018.5, 1018.4, 1018.3, 1018.1, 1018.1, 1018.1, 
    1018.1, 1018, 1018, 1018, 1017.9, 1017.7, 1017.6, 1017.3, 1017, 1016.7, 
    1016.6, 1016.5, 1016.5, 1016.4, 1016.4, 1016.4, 1016.2, 1015.9, 1015.6, 
    1015.2, 1015.2, 1015.1, 1015.1, 1015, 1015, 1015.1, 1015.2, 1015.2, 
    1015.1, 1015, 1014.7, 1014.7, 1014.7, 1014.7, 1014.7, 1014.7, 1014.6, 
    1014.5, 1014.7, 1014.8, 1014.9, 1015.1, 1015.3, 1015.4, 1015.6, 1015.8, 
    1016.2, 1016.4, 1016.6, 1016.8, 1016.9, 1017.1, 1017.2, 1017.3, 1017.3, 
    1017.2, 1017.1, 1017.1, 1017.3, 1017.3, 1017.3, 1017.4, 1017.4, 1017.5, 
    1017.5, 1017.3, 1017, 1017.1, 1017.1, 1017.1, 1017, 1017, 1017, 1016.9, 
    1017, 1016.9, 1016.6, 1016.5, 1016.3, 1016.1, 1016.1, 1016.1, 1015.9, 
    1015.9, 1015.7, 1015.5, 1015.6, 1015.4, 1015.3, 1014.8, 1014.4, 1014.2, 
    1013.8, 1013.6, 1013.3, 1013.2, 1012.9, 1012.5, 1012.3, 1012.2, 1012.1, 
    1011.9, 1011.9, 1011.8, 1012.1, 1012.4, 1012.6, 1013, 1013.5, 1013.9, 
    1014.1, 1014, 1014.2, 1014.8, 1014.8, 1015.2, 1015.4, 1015.7, 1015.9, 
    1016.4, 1016.5, 1016.6, 1017, 1017.1, 1016.9, 1017.2, 1017.6, 1017.6, 
    1018, 1017.8, 1018, 1018, 1018.3, 1018.5, 1018.7, 1018.7, 1018.8, 1019.1, 
    1019.2, 1019.4, 1019.5, 1019.7, 1019.2, 1019.4, 1019.6, 1020, 1020.1, 
    1019.8, 1020.1, 1020.1, 1020.2, 1020.1, 1019.9, 1019.8, 1019.9, 1019.9, 
    1020.1, 1020.6, 1020.5, 1021, 1020.9, 1021.3, 1021.8, 1021.9, 1022.1, 
    1022, 1021.9, 1022, 1021.8, 1021.9, 1022.1, 1022.2, 1022.1, 1022, 1022.2, 
    1022, 1021.8, 1021.4, 1021.2, 1021, 1020.8, 1020.9, 1020.7, 1020.3, 1020, 
    1019.6, 1019.2, 1018.6, 1018.5, 1017.6, 1017.2, 1016.7, 1016, 1015.5, 
    1015, 1014.2, 1013.9, 1013.6, 1012.9, 1012.5, 1012.2, 1012.1, 1011.8, 
    1011.7, 1011.5, 1011.4, 1011.4, 1011.3, 1011.2, 1011.2, 1011.1, 1011.2, 
    1011.1, 1010.9, 1010.8, 1010.6, 1010.3, 1011.1, 1011.1, 1011.3, 1011.3, 
    1011.9, 1011.9, 1011.8, 1012.1, 1012.2, 1012.4, 1012.3, 1012.3, 1012.7, 
    1012.6, 1012.8, 1013.3, 1013.1, 1013.2, 1013.4, 1013.1, 1013.3, 1013.3, 
    1013.5, 1013.3, 1013.6, 1013.8, 1014, 1013.9, 1014.2, 1014.4, 1014.3, 
    1014.4, 1014.2, 1014.2, 1014.2, 1014.3, 1014.5, 1014.6, 1014.6, 1014.6, 
    1014.6, 1014.6, 1014.7, 1014.9, 1014.7, 1014.8, 1014.8, 1015, 1015.1, 
    1015.2, 1015.3, 1015.4, 1015.4, 1015.4, 1015.5, 1015.3, 1015.4, 1015.6, 
    1015.7, 1015.8, 1016, 1016, 1015.9, 1015.6, 1015.6, 1015.6, 1015.5, 
    1015.2, 1015, 1014.8, 1014.6, 1014.5, 1014.5, 1014, 1014.1, 1013.8, 
    1013.5, 1013.4, 1013.1, 1013, 1012.7, 1012.5, 1012.2, 1012, 1011.8, 
    1011.5, 1011.6, 1011.5, 1011.3, 1011, 1010.8, 1010.6, 1010.5, 1010.1, 
    1010, 1009.9, 1009.7, 1009.4, 1009.1, 1008.9, 1008.7, 1008.5, 1008.2, 
    1008, 1007.8, 1007.7, 1007.8, 1007.5, 1007.6, 1007.7, 1007.9, 1008, 
    1008.1, 1008.3, 1008.5, 1008.6, 1008.7, 1008.9, 1009, 1009, 1009.3, 
    1009.4, 1009.7, 1010.1, 1010.3, 1010.5, 1010.5, 1010.6, 1010.7, 1010.9, 
    1010.9, 1011, 1011, 1011.1, 1011.1, 1011.3, 1011.3, 1011.3, 1011.4, 
    1011.2, 1011.2, 1011.3, 1011.3, 1011.3, 1011.3, 1011.5, 1011.6, 1011.8, 
    1012.1, 1012.2, 1012.2, 1012.3, 1012.4, 1012.4, 1012.5, 1012.6, 1012.7, 
    1012.9, 1013.2, 1013.4, 1013.5, 1013.7, 1013.9, 1014, 1014.1, 1014.4, 
    1014.6, 1014.9, 1015.3, 1015.4, 1015.7, 1015.8, 1015.9, 1016.2, 1016.4, 
    1016.3, 1016.3, 1016.2, 1016.2, 1016.1, 1015.9, 1015.9, 1015.7, 1015.4, 
    1015.2, 1014.9, 1014.7, 1014.5, 1014.4, 1014.2, 1014.2, 1014.1, 1014.2, 
    1014.1, 1014.1, 1014, 1013.7, 1013.8, 1013.7, 1013.6, 1013.4, 1013.1, 
    1013.2, 1013.3, 1013.3, 1013.3, 1013.2, 1013.3, 1013.2, 1013.2, 1013, 
    1012.9, 1012.6, 1012.5, 1012.5, 1012.5, 1012.4, 1012.4, 1012.2, 1012, 
    1011.9, 1011.6, 1011.6, 1011.5, 1011.5, 1011.7, 1011.7, 1011.9, 1012.2, 
    1012.6, 1012.7, 1013, 1013.2, 1013.3, 1013.5, 1013.9, 1014.4, 1014.6, 
    1015.1, 1015.7, 1016.3, 1016.7, 1017.1, 1017.7, 1018.2, 1018.6, 1019.1, 
    1019.5, 1019.7, 1020.1, 1020.4, 1020.9, 1021.4, 1021.8, 1022.2, 1022.6, 
    1022.9, 1023.2, 1023.3, 1023.5, 1023.6, 1023.9, 1024.3, 1024.6, 1024.9, 
    1025.4, 1025.9, 1026.4, 1026.9, 1027.3, 1027.5, 1027.8, 1028.3, 1028.6, 
    1029, 1029.6, 1030.2, 1030.7, 1031.1, 1031.6, 1032, 1032.3, 1032.7, 
    1033.1, 1033.5, 1033.9, 1034.4, 1034.9, 1035.4, 1035.7, 1035.9, 1036.1, 
    1036, 1036.2, 1035.8, 1035.8, 1036.2, 1036.1, 1036.1, 1036, 1036, 1035.8, 
    1036, 1035.5, 1035.6, 1035.8, 1035.3, 1034.9, 1034.7, 1034.7, 1034.7, 
    1035, 1035.1, 1035, 1035, 1034.8, 1035, 1034.8, 1034.5, 1034.4, 1034.1, 
    1034.1, 1033.8, 1033.7, 1033.6, 1033.7, 1033.6, 1033.2, 1032.9, 1032.6, 
    1032.1, 1031.6, 1031.2, 1031, 1030.9, 1030.8, 1030.6, 1030.3, 1030.1, 
    1030.2, 1030.3, 1030.1, 1030.2, 1030.2, 1030.4, 1030.7, 1031.2, 1031.7, 
    1032, 1032.5, 1033.1, 1033.5, 1033.7, 1034, 1034.3, 1034.6, 1034.8, 
    1035.2, 1035.5, 1035.7, 1035.9, 1036.1, 1036.2, 1036.5, 1036.7, 1036.8, 
    1036.7, 1036.3, 1036.2, 1035.9, 1035.7, 1035.5, 1035.5, 1035.2, 1035.1, 
    1034.9, 1034.8, 1034.5, 1034.3, 1034.1, 1033.8, 1033.7, 1033.4, 1033.1, 
    1032.9, 1032.7, 1032.2, 1031.8, 1031.3, 1031.1, 1030.6, 1030, 1029.4, 
    1028.6, 1028.1, 1027.8, 1027.4, 1026.8, 1026.3, 1026, 1025.4, 1024.9, 
    1024.5, 1024.1, 1023.5, 1022.8, 1022.3, 1021.9, 1021.3, 1021.3, 1021.3, 
    1021, 1021, 1020.7, 1020.4, 1020.3, 1020.1, 1019.9, 1019.8, 1019.6, 
    1019.5, 1019.5, 1019.4, 1019.5, 1019.7, 1019.8, 1019.7, 1019.6, 1019.3, 
    1019.1, 1019.2, 1019.3, 1019.3, 1019.6, 1019.8, 1019.8, 1019.9, 1019.7, 
    1019.8, 1019.8, 1019.7, 1019.6, 1019.4, 1019.5, 1019.6, 1019.7, 1020, 
    1020.1, 1020.3, 1020.3, 1020.3, 1020.2, 1020.4, 1020.6, 1020.8, 1021.2, 
    1021.7, 1022.2, 1022.4, 1022.6, 1022.9, 1023.2, 1023.4, 1023.5, 1023.5, 
    1023.6, 1023.9, 1024.1, 1024.3, 1024.6, 1024.7, 1024.9, 1024.8, 1024.8, 
    1024.8, 1024.9, 1024.8, 1024.5, 1024.5, 1024.7, 1024.8, 1024.7, 1024.5, 
    1024.4, 1024.3, 1024.2, 1023.8, 1023.4, 1023, 1023, 1022.6, 1022.3, 
    1022.2, 1022, 1021.9, 1021.5, 1021.3, 1021.2, 1021, 1020.8, 1020.6, 
    1020.5, 1020.8, 1021, 1021.4, 1021.7, 1021.9, 1022, 1022.2, 1022.3, 
    1022.5, 1022.5, 1022.8, 1022.9, 1022.9, 1023, 1022.9, 1023, 1023.1, 
    1022.9, 1022.7, 1022.6, 1022.2, 1021.9, 1021.5, 1021.3, 1021.3, 1021.2, 
    1021.2, 1021.4, 1021.1, 1021.1, 1021, 1020.8, 1020.7, 1020.5, 1020.2, 
    1019.9, 1019.7, 1019.4, 1019.1, 1019.1, 1019.1, 1018.9, 1018.8, 1018.5, 
    1018.3, 1018.1, 1018.1, 1018, 1017.8, 1017.9, 1017.8, 1017.7, 1017.6, 
    1017.5, 1017.6, 1017.5, 1017.1, 1016.7, 1016.5, 1016.2, 1016.1, 1016, 
    1015.7, 1015.6, 1015.4, 1015, 1014.7, 1014.5, 1014.4, 1014.3, 1014.1, 
    1014.1, 1014.1, 1014, 1014.3, 1014.4, 1014.7, 1014.8, 1015, 1015.3, 
    1015.4, 1015.5, 1015.5, 1015.7, 1016.2, 1016.2, 1016.5, 1016.9, 1017.2, 
    1017.5, 1017.9, 1018.1, 1018.3, 1018.4, 1018.5, 1018.7, 1019, 1019.2, 
    1019.4, 1019.5, 1019.7, 1019.7, 1019.8, 1019.9, 1019.8, 1019.9, 1019.7, 
    1019.5, 1019.5, 1019.2, 1019.2, 1019.3, 1019.2, 1019.2, 1019, 1019, 
    1018.9, 1018.8, 1018.6, 1018.8, 1018.8, 1018.9, 1018.9, 1019, 1019, 
    1018.9, 1019, 1019, 1018.9, 1018.6, 1018.4, 1018, 1018.2, 1018.1, 1018, 
    1017.4, 1017.1, 1017.2, 1017.1, 1017, 1017, 1016.6, 1016.2, 1015.7, 
    1015.3, 1015.1, 1014.6, 1014.5, 1014.2, 1013.5, 1012.6, 1012.3, 1011.7, 
    1011.3, 1011.3, 1011, 1010.8, 1010.7, 1010.4, 1010.4, 1010.2, 1009.3, 
    1008.5, 1008.1, 1007.3, 1006.8, 1006.6, 1005.9, 1006, 1005.9, 1006.1, 
    1006.3, 1006.7, 1007.1, 1007.6, 1008.3, 1009, 1009.4, 1009.9, 1010.5, 
    1011, 1011.2, 1011.7, 1012.1, 1012.4, 1012.8, 1013.4, 1013.6, 1013.9, 
    1014.1, 1014.1, 1014.2, 1014.5, 1014.7, 1014.8, 1014.9, 1015.2, 1015.3, 
    1015.3, 1015.4, 1015.5, 1015.3, 1015.2, 1015.2, 1014.9, 1014.7, 1014.4, 
    1014.4, 1014.2, 1014.2, 1013.9, 1013.8, 1013.4, 1013.1, 1012.4, 1012.1, 
    1011.4, 1010.9, 1010.3, 1010.1, 1009.9, 1009.4, 1008.8, 1008.2, 1007.7, 
    1007.2, 1006.6, 1005.7, 1005.3, 1004.7, 1003.9, 1003.2, 1002.5, 1002, 
    1001.5, 1001.1, 1000.6, 1000.2, 999.9, 999.9, 999.7, 999.5, 999.3, 999.1, 
    999.1, 999.1, 999.2, 999.1, 999, 998.9, 998.9, 998.8, 998.9, 999, 999.1, 
    999.1, 999.2, 999.3, 999.3, 999.4, 999.3, 999.2, 999.2, 999.3, 999.3, 
    999.5, 999.8, 999.9, 1000.2, 1000.4, 1000.5, 1000.4, 1000.5, 1000.4, 
    1000.4, 1000.4, 1000.3, 1000.4, 1000.4, 1000.5, 1000.5, 1000.4, 1000.3, 
    1000.2, 1000, 999.7, 999.4, 999.3, 999.5, 999.5, 999.7, 999.9, 1000, 
    1000.1, 999.9, 999.6, 999.3, 999.3, 998.8, 998.7, 998.6, 998.4, 998.3, 
    998, 997.7, 997.5, 997.4, 997.3, 997, 996.5, 996.2, 995.3, 995.5, 996, 
    996.1, 996.3, 996.8, 996.8, 997.1, 997.2, 997.1, 997, 997, 997, 997, 
    996.9, 996.9, 997.1, 997, 996.8, 997, 997, 996.9, 997, 997.3, 997.8, 
    998.3, 998.4, 998.7, 999.1, 999.6, 999.9, 1000.3, 1000.7, 1001, 1001.3, 
    1001.6, 1001.9, 1002.3, 1002.7, 1002.9, 1003.3, 1003.8, 1004.1, 1004.3, 
    1004.5, 1004.8, 1005, 1005.2, 1005.5, 1005.7, 1006.1, 1006.4, 1006.7, 
    1007, 1007.4, 1007.7, 1008.1, 1008.5, 1008.9, 1009.3, 1009.6, 1010.2, 
    1010.6, 1010.9, 1011.7, 1012.2, 1012.8, 1013.2, 1013.5, 1014, 1014.2, 
    1014.4, 1014.7, 1014.7, 1014.9, 1015.2, 1015.3, 1015.2, 1015.5, 1015.9, 
    1016.3, 1016.6, 1016.7, 1017, 1017.2, 1017.4, 1017.8, 1018, 1018.3, 
    1018.6, 1018.9, 1019.1, 1019.3, 1019.5, 1019.6, 1019.7, 1019.8, 1019.9, 
    1020.2, 1020.3, 1020.4, 1020.5, 1020.5, 1020.1, 1019.9, 1019.5, 1019.2, 
    1018.9, 1018.7, 1018.6, 1018.2, 1018, 1017.8, 1017.6, 1017.4, 1016.9, 
    1016.5, 1016.3, 1015.8, 1015.7, 1015.8, 1015.8, 1015.9, 1016, 1016.1, 
    1016.2, 1016.3, 1016.1, 1016.1, 1015.8, 1015.8, 1015.6, 1015.5, 1015.7, 
    1015.8, 1015.9, 1015.9, 1015.6, 1015.7, 1015.6, 1015.6, 1015.5, 1015.5, 
    1015.4, 1015.4, 1015.6, 1015.5, 1015.4, 1015.3, 1015.3, 1015.3, 1015.3, 
    1015.2, 1015.1, 1015, 1015.2, 1015.1, 1015.3, 1015.4, 1015.5, 1015.5, 
    1015.5, 1015.7, 1015.8, 1016, 1016.2, 1016.1, 1016.2, 1016.4, 1016.5, 
    1016.7, 1016.9, 1016.9, 1016.9, 1017, 1017.2, 1017.3, 1017.2, 1017.2, 
    1017.2, 1017.2, 1017.2, 1017, 1016.9, 1016.9, 1017, 1016.9, 1016.9, 
    1016.8, 1016.7, 1016.2, 1015.8, 1015.4, 1015.1, 1014.9, 1014.7, 1014.3, 
    1013.9, 1013.6, 1013.3, 1012.9, 1012.6, 1012.4, 1012.1, 1011.7, 1011.4, 
    1011.2, 1011.1, 1011.1, 1011.1, 1010.6, 1010.4, 1010, 1009.8, 1009.3, 
    1008.6, 1007.7, 1007.2, 1006.1, 1005.3, 1004.8, 1004.3, 1004.3, 1004.9, 
    1005.2, 1005.2, 1005.2, 1005.2, 1005.6, 1005.7, 1005.9, 1006, 1006.2, 
    1006.4, 1006.4, 1006.4, 1006.3, 1006.5, 1006.2, 1006, 1006.1, 1006.2, 
    1006.9, 1007.5, 1008.4, 1009.5, 1010.4, 1011.6, 1012.6, 1013.9, 1014.5, 
    1015.6, 1016.2, 1017.5, 1018.5, 1019.6, 1020.7, 1021.7, 1022.6, 1023.8, 
    1024.9, 1025.1, 1025.7, 1026.7, 1027.2, 1027.7, 1028.3, 1028.9, 1029.5, 
    1030.2, 1030.6, 1030.9, 1031.3, 1031.7, 1032, 1032.1, 1032.2, 1032.4, 
    1032.6, 1032.8, 1032.8, 1032.9, 1033, 1032.9, 1032.8, 1032.6, 1032.3, 
    1032.2, 1031.9, 1031.5, 1031.4, 1031.2, 1030.9, 1030.7, 1030.4, 1030, 
    1029.6, 1029.3, 1028.7, 1028.2, 1027.8, 1027.2, 1026.7, 1026.3, 1025.8, 
    1025.2, 1024.7, 1024.1, 1023.4, 1022.8, 1022.2, 1021.5, 1021.1, 1020.4, 
    1019.9, 1019.4, 1018.9, 1018.4, 1018.1, 1017.7, 1017.5, 1017.2, 1016.9, 
    1016.4, 1016.2, 1015.9, 1015.8, 1015.7, 1015.5, 1015.5, 1015.5, 1015.4, 
    1015.4, 1015.4, 1015.6, 1015.9, 1016.2, 1016.6, 1017.2, 1017.9, 1018.7, 
    1019.2, 1019.6, 1020.2, 1020.7, 1021, 1021.4, 1021.2, 1021.4, 1021.3, 
    1021.5, 1021.3, 1021.3, 1021.3, 1020.8, 1020.4, 1020, 1019.6, 1018.9, 
    1018.3, 1017.7, 1017.2, 1016.4, 1016.1, 1015.8, 1015, 1014.4, 1013.8, 
    1013.2, 1012.6, 1012.3, 1012.1, 1011.7, 1012, 1011.8, 1012.2, 1012.2, 
    1012.4, 1012.6, 1012.5, 1012.8, 1013.2, 1013.4, 1013.3, 1013.5, 1013.9, 
    1014.1, 1014.4, 1014.6, 1014.9, 1015, 1015.2, 1015.4, 1015.3, 1015.6, 
    1015.5, 1015.3, 1015.7, 1015.6, 1015.3, 1015.6, 1015.7, 1015.3, 1015.5, 
    1015.7, 1015.6, 1015.7, 1015.6, 1015.5, 1015.7, 1015.7, 1015.8, 1015.9, 
    1016.5, 1017, 1017.3, 1017.5, 1017.7, 1018, 1018.2, 1018.6, 1018.9, 
    1019.3, 1019.9, 1020.3, 1020.7, 1020.9, 1021.1, 1021.4, 1021.5, 1021.7, 
    1021.7, 1021.8, 1022, 1022.2, 1022.6, 1022.6, 1022.6, 1022.8, 1023, 
    1023.2, 1023.1, 1022.9, 1022.7, 1022.5, 1022.3, 1022.2, 1022.1, 1021.9, 
    1021.4, 1021.2, 1021.1, 1020.8, 1020.6, 1020.1, 1019.8, 1019.6, 1019.3, 
    1019.2, 1019, 1018.9, 1018.5, 1018.4, 1018.2, 1017.7, 1017.6, 1017.5, 
    1017.2, 1016.8, 1016.5, 1016.3, 1016.2, 1015.8, 1015.7, 1015.6, 1015.4, 
    1015.1, 1014.9, 1014.7, 1014.4, 1014.2, 1014.1, 1014, 1013.9, 1013.8, 
    1013.6, 1013.6, 1013.4, 1013.4, 1013.2, 1013.1, 1013, 1013, 1013.1, 
    1013.2, 1013.2, 1013.4, 1013.5, 1013.8, 1014, 1014.1, 1014.1, 1014.2, 
    1014.2, 1014.1, 1014.3, 1014.5, 1014.8, 1015.3, 1015.5, 1015.6, 1015.7, 
    1015.7, 1015.5, 1015.6, 1015.6, 1015.6, 1015.7, 1015.8, 1015.8, 1015.6, 
    1015.5, 1015.4, 1015.1, 1015, 1014.9, 1014.7, 1014.5, 1014.5, 1014.5, 
    1014.6, 1014.4, 1014.3, 1014.2, 1014.5, 1014.5, 1014, 1014, 1014, 1014, 
    1013.9, 1013.7, 1013.9, 1014.1, 1014.1, 1014.1, 1014, 1013.8, 1013.7, 
    1013.4, 1013.2, 1012.9, 1012.6, 1012.3, 1011.9, 1011.6, 1011.2, 1010.8, 
    1010.4, 1009.8, 1009.4, 1009.1, 1008.7, 1008.2, 1007.9, 1007.6, 1007, 
    1006.7, 1006.3, 1006.2, 1006.2, 1006.2, 1006.3, 1006.5, 1006.5, 1006.4, 
    1006.5, 1006.8, 1007.1, 1007.3, 1007.6, 1007.9, 1008.3, 1008.4, 1008.6, 
    1008.5, 1008.6, 1008.8, 1008.9, 1009, 1009.3, 1009.5, 1009.7, 1010.1, 
    1010.2, 1010.3, 1010.4, 1010.4, 1010.5, 1010.4, 1010.4, 1010.4, 1010.5, 
    1010.7, 1010.7, 1010.7, 1010.7, 1010.7, 1010.7, 1010.7, 1010.9, 1010.8, 
    1010.8, 1011.1, 1011.3, 1011.4, 1011.6, 1011.7, 1011.8, 1012.2, 1012.4, 
    1012.4, 1012.5, 1012.6, 1012.7, 1013, 1013.4, 1013.6, 1013.8, 1014, 
    1014.4, 1014.5, 1014.6, 1014.6, 1015, 1015.3, 1015.5, 1015.7, 1016, 
    1016.4, 1016.6, 1016.9, 1017, 1017.3, 1017.5, 1017.6, 1017.7, 1018.1, 
    1018, 1018.3, 1018.4, 1018.8, 1018.7, 1018.7, 1018.7, 1018.9, 1018.9, 
    1018.9, 1018.9, 1019, 1018.7, 1018.3, 1018.3, 1018, 1017.9, 1017.7, 
    1017.5, 1017.1, 1016.7, 1015.8, 1015.2, 1015.1, 1014.8, 1014, 1013.2, 
    1012.1, 1011.8, 1011.3, 1010.3, 1009.5, 1008.7, 1007.9, 1007.4, 1006.5, 
    1006.4, 1006.1, 1005.9, 1005.8, 1005.6, 1005.9, 1005.6, 1005.3, 1005.2, 
    1004.7, 1004.5, 1004.4, 1004.4, 1004.1, 1004.1, 1004.1, 1004.3, 1004.5, 
    1005, 1004.9, 1005.1, 1005.2, 1005.2, 1005.3, 1005.5, 1005.7, 1006.1, 
    1006.4, 1006.6, 1006.8, 1006.7, 1006.8, 1006.9, 1007.1, 1007.4, 1007.6, 
    1007.7, 1007.7, 1008, 1008, 1008.2, 1008.5, 1008.6, 1008.7, 1008.9, 1009, 
    1009.3, 1009.4, 1009.7, 1009.6, 1009.7, 1010.3, 1010.8, 1010.7, 1010.6, 
    1010.4, 1010.3, 1009.8, 1009.5, 1009.2, 1009, 1008.8, 1008.7, 1008.6, 
    1008.6, 1008.5, 1008.3, 1008.2, 1008, 1007.8, 1007.6, 1007.5, 1007.4, 
    1007.3, 1007.3, 1007.2, 1007.4, 1007.3, 1007.3, 1007.2, 1007, 1006.8, 
    1006.5, 1006.2, 1006.2, 1006, 1005.9, 1005.8, 1005.7, 1005.7, 1005.5, 
    1005.5, 1005.5, 1005.5, 1005.5, 1005.2, 1005.2, 1005.1, 1005, 1005, 1005, 
    1004.9, 1004.6, 1004.7, 1004.3, 1004.3, 1004.3, 1004.2, 1004, 1004.1, 
    1004.2, 1004.2, 1004.4, 1004.6, 1004.9, 1005.3, 1005.7, 1006, 1006, 
    1006.2, 1006, 1006.4, 1006.6, 1006.7, 1007, 1007.1, 1007.1, 1007.3, 
    1007.5, 1007.5, 1007.5, 1007.7, 1007.9, 1008.1, 1008.3, 1008.6, 1008.6, 
    1008.8, 1008.8, 1008.9, 1008.9, 1009.1, 1009.1, 1009, 1008.7, 1008.4, 
    1008.4, 1008.4, 1008.4, 1008.2, 1008.3, 1008.3, 1008.1, 1008, 1007.9, 
    1007.7, 1007.5, 1007.6, 1007.6, 1007.7, 1007.3, 1007.4, 1007.3, 1007.5, 
    1007.5, 1007.3, 1007.3, 1007.1, 1007, 1006.8, 1006.5, 1006.5, 1006.3, 
    1006.2, 1005.9, 1005.6, 1005.4, 1005.2, 1005, 1004.9, 1005, 1004.7, 
    1004.8, 1004.9, 1005.3, 1005.8, 1005.9, 1006.3, 1006.5, 1006.4, 1006.8, 
    1006.9, 1007.1, 1007.3, 1007.5, 1007.7, 1008, 1007.8, 1007.9, 1007.8, 
    1007.8, 1007.8, 1007.8, 1007.7, 1007.6, 1007.7, 1007.6, 1007.9, 1008.1, 
    1008.4, 1008.5, 1008.9, 1008.9, 1009.2, 1009.5, 1009.6, 1009.7, 1010, 
    1010.3, 1010.8, 1011.2, 1011.4, 1011.8, 1012, 1012.3, 1012.6, 1012.8, 
    1012.9, 1013.1, 1013.5, 1013.9, 1014.2, 1014.6, 1014.8, 1015.1, 1015.4, 
    1015.6, 1015.7, 1015.8, 1015.8, 1016, 1016.1, 1016.2, 1016.2, 1016.3, 
    1016.5, 1016.4, 1016.5, 1016.4, 1016.2, 1016.1, 1016.2, 1015.9, 1015.7, 
    1015.5, 1015.5, 1015.6, 1015.3, 1015.2, 1015.1, 1014.9, 1014.3, 1013.9, 
    1013.7, 1013.3, 1012.9, 1012.7, 1012.6, 1012.3, 1011.7, 1011.4, 1011.3, 
    1010.9, 1010.6, 1010.2, 1009.8, 1009.4, 1009.2, 1009.2, 1009.4, 1009.7, 
    1009.9, 1010.2, 1010.1, 1010.1, 1010.2, 1010.2, 1010.4, 1010.5, 1010.7, 
    1010.9, 1011.1, 1011.4, 1011.5, 1011.6, 1011.5, 1011.6, 1011.4, 1011.5, 
    1011.3, 1011.4, 1011.6, 1011.4, 1011.5, 1011.6, 1011.5, 1011.6, 1011.5, 
    1011.7, 1011.6, 1011.6, 1011.6, 1011.7, 1011.8, 1011.9, 1012.1, 1012.4, 
    1012.7, 1012.8, 1012.9, 1013.1, 1013.2, 1013.5, 1013.8, 1013.8, 1014, 
    1014.2, 1014.5, 1014.6, 1014.8, 1015.1, 1015.1, 1015.2, 1015.2, 1015.4, 
    1015.5, 1015.6, 1015.9, 1015.8, 1016, 1016.1, 1016.2, 1016.4, 1016.4, 
    1016.5, 1016.6, 1016.6, 1016.4, 1016.3, 1016.3, 1016.4, 1016.5, 1016.3, 
    1016.4, 1016.4, 1016.1, 1016.1, 1015.9, 1015.6, 1015.4, 1015, 1014.8, 
    1014.8, 1014.6, 1014.7, 1014.7, 1014.4, 1014.2, 1014, 1013.8, 1013.7, 
    1013.7, 1013.7, 1013.7, 1013.7, 1013.6, 1013.7, 1013.8, 1013.8, 1013.8, 
    1013.7, 1013.5, 1013.5, 1013.5, 1013.3, 1013.3, 1013.5, 1013.4, 1013.4, 
    1013.3, 1013.2, 1013.1, 1013, 1012.9, 1012.5, 1012.2, 1012.1, 1011.7, 
    1011.4, 1010.9, 1010.9, 1010.6, 1010.3, 1010, 1009.7, 1009.5, 1009.2, 
    1008.9, 1008.8, 1008.5, 1008.5, 1008.3, 1008.5, 1008.5, 1008.4, 1008.2, 
    1008, 1007.6, 1007, 1006.5, 1006.4, 1006, 1005.5, 1005.2, 1004.6, 1004.1, 
    1003.5, 1003.1, 1002.5, 1002, 1001.5, 1000.2, 999.7, 999.1, 998, 996.6, 
    995, 993.1, 991.7, 992.1, 990.2, 990.8, 991.1, 991, 990.5, 990.4, 991, 
    991.5, 992.2, 993.2, 994.5, 995.5, 996.5, 997.3, 998.2, 999.3, 999.9, 
    1000.8, 1001.6, 1002.4, 1003.1, 1004.1, 1004.9, 1005.4, 1006, 1006.7, 
    1007, 1007.5, 1008.2, 1008.6, 1009.3, 1010, 1010.9, 1011.5, 1012.1, 
    1012.8, 1013.5, 1013.8, 1014.3, 1014.7, 1015, 1015.5, 1015.9, 1016.3, 
    1017, 1017.4, 1017.7, 1017.9, 1018.1, 1018.5, 1018.7, 1018.5, 1018.5, 
    1018.7, 1018.9, 1019.1, 1019.3, 1019.3, 1019.4, 1019.4, 1019.3, 1019.1, 
    1019.3, 1019.2, 1019.2, 1019, 1019.2, 1019.4, 1019.4, 1019.3, 1019, 
    1018.9, 1019, 1018.9, 1018.7, 1018.4, 1018.2, 1018.2, 1018.5, 1018.2, 
    1018.2, 1018.3, 1018.5, 1018.4, 1018.5, 1018.4, 1018, 1017.9, 1018, 
    1018.2, 1018.3, 1018.5, 1018.5, 1018.7, 1018.8, 1018.9, 1019.1, 1018.9, 
    1019, 1019.2, 1019.4, 1019.7, 1020.1, 1020.3, 1020.6, 1020.9, 1021.2, 
    1021.4, 1021.8, 1021.7, 1021.7, 1021.8, 1021.9, 1022.1, 1022.5, 1022.5, 
    1022.6, 1022.5, 1022.6, 1022.4, 1022.6, 1022.5, 1022.5, 1022.3, 1022, 
    1022.1, 1022, 1022, 1021.8, 1021.7, 1021.8, 1021.7, 1021.4, 1021.3, 1021, 
    1020.4, 1020.1, 1020, 1019.8, 1019.6, 1019.4, 1019.3, 1019.1, 1018.9, 
    1018.7, 1018.4, 1018.3, 1017.8, 1017.5, 1017.4, 1017.4, 1017.6, 1017.3, 
    1017.5, 1017.2, 1016.9, 1016.8, 1016.6, 1016.3, 1016.1, 1016, 1015.7, 
    1015.7, 1015.3, 1015.2, 1015.6, 1015.6, 1015.6, 1015.5, 1015, 1014.8, 
    1014.4, 1013.9, 1013.8, 1014.1, 1013.7, 1013.8, 1013.4, 1013.2, 1012.8, 
    1012.4, 1011.8, 1011.2, 1011.2, 1011.1, 1010.9, 1010.9, 1011.1, 1011.3, 
    1010.8, 1010.7, 1010.6, 1010.7, 1010.5, 1010.3, 1010, 1010.2, 1010.3, 
    1010.5, 1011.1, 1011.3, 1011.7, 1011.7, 1011.7, 1011.8, 1011.5, 1011.4, 
    1011.2, 1011, 1010.9, 1010.8, 1010.7, 1010.6, 1010, 1009.7, 1009.9, 
    1009.2, 1009, 1009.1, 1009.1, 1009.1, 1009.3, 1009.5, 1009.6, 1009.7, 
    1010.1, 1010.1, 1010.4, 1010.7, 1010.8, 1010.6, 1010.2, 1010.1, 1010.3, 
    1010.5, 1010.3, 1010.1, 1010.1, 1010.1, 1009.7, 1009.4, 1009, 1008.8, 
    1008.8, 1008.9, 1008.8, 1008.3, 1008, 1007.8, 1007.8, 1007.7, 1007.6, 
    1007.5, 1007.3, 1007.2, 1007, 1007.1, 1007.3, 1007.3, 1007.3, 1007.4, 
    1007.5, 1007.5, 1007.4, 1007.5, 1007.4, 1007.3, 1007.2, 1007.1, 1007.2, 
    1007.1, 1007.2, 1007.3, 1007.3, 1007.5, 1007.5, 1007.4, 1007.4, 1007.6, 
    1007.6, 1007.5, 1007.5, 1007.5, 1007.6, 1007.6, 1007.6, 1007.5, 1007.5, 
    1007.7, 1007.6, 1007.5, 1007.3, 1007.2, 1007.4, 1007.2, 1007.3, 1007.4, 
    1007.6, 1007.8, 1007.8, 1007.9, 1008, 1008.1, 1008.1, 1008.3, 1008.4, 
    1008.5, 1008.6, 1009, 1009, 1009.4, 1009.5, 1009.5, 1009.5, 1009.6, 
    1009.5, 1009.5, 1009.5, 1009.7, 1009.7, 1009.7, 1009.7, 1009.9, 1009.7, 
    1009.6, 1009.6, 1009.4, 1009.1, 1009.2, 1009.1, 1009, 1009.1, 1009.1, 
    1009.1, 1008.9, 1008.8, 1008.5, 1008, 1007.6, 1007.6, 1007.4, 1007.1, 
    1007.2, 1007, 1007, 1007, 1006.9, 1006.6, 1006.1, 1005.7, 1005.6, 1005.2, 
    1004.9, 1004.3, 1004.2, 1004.1, 1003.7, 1003.8, 1003.9, 1003.6, 1002.7, 
    1002.1, 1001.1, 1000.3, 999.9, 999.6, 999, 998.9, 998.9, 999.1, 999.4, 
    999.4, 999.5, 999.5, 999.5, 999.6, 999.4, 999.5, 999.5, 999.4, 999.1, 
    998.8, 998.9, 998.9, 998.8, 998.5, 998.4, 998.2, 998.3, 998.3, 998.3, 
    998.3, 998.2, 998.4, 998.7, 998.9, 999.1, 999.3, 999.4, 999.5, 999.9, 
    1000.4, 1000.9, 1001.3, 1001.9, 1002.4, 1002.9, 1003.5, 1004.2, 1004.6, 
    1005.1, 1005.4, 1005.9, 1006.4, 1006.9, 1007.5, 1008.2, 1008.7, 1009.3, 
    1009.9, 1010.3, 1010.7, 1010.9, 1011.2, 1011.7, 1012.4, 1012.9, 1013.3, 
    1013.8, 1014.3, 1014.8, 1015.5, 1015.8, 1016, 1016.2, 1016.4, 1016.5, 
    1016.6, 1017, 1017, 1017.1, 1017.2, 1017.4, 1017.5, 1017.7, 1017.7, 
    1017.5, 1017.6, 1017.7, 1017.8, 1017.9, 1017.9, 1018, 1018.4, 1018.5, 
    1018.5, 1018.3, 1018.4, 1018.2, 1017.9, 1017.9, 1018, 1018.1, 1018.1, 
    1018.2, 1018.2, 1018, 1018.1, 1018.1, 1018, 1017.8, 1017.8, 1017.7, 
    1017.6, 1017.5, 1017.7, 1017.6, 1017.7, 1017.5, 1017.4, 1017.5, 1017.5, 
    1017.1, 1016.9, 1016.5, 1016.5, 1016.2, 1016, 1015.8, 1015.6, 1015.5, 
    1015.2, 1014.9, 1014.3, 1013.9, 1013.5, 1013.3, 1013.2, 1013.3, 1013.6, 
    1014, 1014.1, 1014.3, 1014.3, 1014.7, 1015.1, 1015.5, 1015.8, 1016.1, 
    1016.4, 1016.7, 1017.1, 1017.3, 1017.4, 1017.9, 1018, 1018.3, 1018.5, 
    1018.6, 1018.7, 1018.9, 1019.3, 1019.4, 1019.8, 1020.1, 1020.3, 1020.5, 
    1020.7, 1020.7, 1020.8, 1020.9, 1020.9, 1021.2, 1021.3, 1021.7, 1021.9, 
    1022.2, 1022.3, 1022.4, 1022.6, 1022.7, 1022.7, 1022.8, 1022.7, 1022.7, 
    1022.7, 1022.9, 1023.2, 1023.4, 1023.6, 1023.5, 1023.6, 1023.6, 1023.6, 
    1023.6, 1023.5, 1023.4, 1023.5, 1023.4, 1023.2, 1023.2, 1022.9, 1022.7, 
    1022.7, 1022.5, 1022.4, 1022.2, 1022, 1021.9, 1021.7, 1021.5, 1021.4, 
    1021.8, 1021.8, 1021.5, 1021.4, 1021.3, 1021.4, 1021.3, 1021.2, 1020.9, 
    1020.7, 1020.7, 1020.8, 1020.9, 1020.8, 1020.7, 1020.6, 1020.3, 1019.9, 
    1019.7, 1019.6, 1019.2, 1018.9, 1018.7, 1018.6, 1018.4, 1018.1, 1017.6, 
    1017.4, 1016.9, 1016.7, 1016.4, 1015.9, 1015.6, 1015.2, 1015, 1014.9, 
    1014.8, 1014.6, 1014.5, 1014.4, 1014.2, 1014, 1014.2, 1014.2, 1014.3, 
    1014.2, 1014.2, 1014.2, 1014.3, 1014.3, 1014.3, 1014.5, 1014.4, 1014.4, 
    1014.5, 1014.7, 1014.7, 1014.7, 1014.8, 1015, 1015.2, 1015, 1014.6, 
    1014.2, 1013.8, 1013.4, 1013, 1012.7, 1012.3, 1011.7, 1010.8, 1010.1, 
    1010.2, 1010.2, 1010.3, 1010.5, 1010.5, 1010.5, 1010.6, 1010.6, 1010.6, 
    1010.5, 1010.5, 1010.6, 1010.9, 1011, 1011.1, 1010.9, 1010.8, 1010.6, 
    1010.6, 1010.6, 1010.7, 1010.6, 1010.6, 1010.7, 1010.9, 1010.9, 1011.1, 
    1011.5, 1011.5, 1011.6, 1011.6, 1011.8, 1011.6, 1011.7, 1011.9, 1012, 
    1012.2, 1012.4, 1012.6, 1012.9, 1013, 1013, 1012.9, 1013, 1013.1, 1013.3, 
    1013.6, 1013.7, 1014.2, 1014.5, 1014.6, 1014.8, 1015.1, 1014.9, 1014.9, 
    1015.1, 1015, 1014.8, 1014.8, 1014.9, 1014.9, 1014.9, 1014.9, 1014.8, 
    1014.7, 1014.4, 1014.1, 1013.8, 1013.7, 1013.5, 1013.7, 1013.8, 1014.1, 
    1014.2, 1014, 1014, 1013.8, 1013.7, 1013.5, 1013.2, 1013, 1012.8, 1012.5, 
    1012.4, 1012.3, 1012.2, 1011.9, 1011.7, 1011.4, 1011.2, 1010.9, 1010.6, 
    1010.4, 1010.2, 1010.2, 1010.3, 1010.4, 1010.4, 1010.1, 1009.8, 1009.7, 
    1009.5, 1009.3, 1009, 1008.8, 1008.6, 1008.3, 1008.4, 1008.2, 1008.1, 
    1008.1, 1008, 1007.9, 1007.9, 1007.7, 1007.4, 1007.3, 1007.2, 1007, 
    1007.2, 1007, 1007.1, 1007.1, 1007.1, 1007, 1006.9, 1006.7, 1006.4, 
    1006.3, 1006, 1005.9, 1005.9, 1005.8, 1005.8, 1005.8, 1005.7, 1005.7, 
    1005.5, 1005.2, 1005.1, 1004.6, 1004.4, 1004.4, 1004.2, 1004.2, 1004.2, 
    1004.2, 1004.1, 1003.8, 1003.7, 1003.7, 1003.6, 1003.5, 1003.6, 1003.5, 
    1003.6, 1003.7, 1003.7, 1003.8, 1003.8, 1003.7, 1003.6, 1003.6, 1003.4, 
    1003.3, 1003.2, 1003, 1003, 1002.7, 1002.5, 1002.4, 1002.1, 1001.8, 
    1001.5, 1001.3, 1001.1, 1000.8, 1000.6, 1000.5, 1000.4, 1000.3, 1000.3, 
    1000.2, 1000, 999.8, 999.6, 999.5, 999.5, 999.3, 999.2, 999.1, 999.1, 
    999.2, 999.4, 999.4, 999.4, 999.3, 999.2, 999, 999.1, 998.9, 999, 999.2, 
    999.3, 999.6, 999.9, 1000.2, 1000.5, 1000.8, 1000.9, 1001, 1001.2, 
    1001.9, 1002.1, 1002.3, 1002.7, 1002.9, 1003.1, 1003.2, 1003.2, 1003.3, 
    1003.4, 1003.3, 1003.5, 1003.5, 1003.4, 1003.4, 1003.4, 1003.8, 1003.8, 
    1003.6, 1003.2, 1003.1, 1003, 1003.1, 1003, 1003, 1003, 1002.9, 1002.9, 
    1002.7, 1002.5, 1002.6, 1002.5, 1002.3, 1002.1, 1001.9, 1001.6, 1001.3, 
    1001.2, 1001.3, 1001.2, 1000.9, 1000.9, 1000.8, 1000.6, 1000.5, 1000.8, 
    1000.5, 1000.8, 1000.9, 1001.2, 1001.4, 1001.9, 1002, 1002.5, 1002.7, 
    1003, 1003.3, 1003.6, 1003.9, 1004.2, 1004.4, 1004.7, 1004.9, 1005.1, 
    1005.3, 1005.5, 1005.5, 1005.6, 1005.6, 1005.6, 1005.7, 1006.1, 1006.1, 
    1006.3, 1006.6, 1006.8, 1007.1, 1007.1, 1007.3, 1007.4, 1007.1, 1007.2, 
    1007.2, 1007.1, 1007.1, 1007, 1006.8, 1006.7, 1006.6, 1006.7, 1006.7, 
    1006.4, 1006.3, 1006.1, 1005.9, 1005.6, 1005.4, 1005.4, 1005.2, 1005.2, 
    1005.1, 1005, 1004.9, 1005, 1005, 1005, 1005, 1005, 1005.2, 1005.6, 
    1005.9, 1005.9, 1006.2, 1006.4, 1006.6, 1006.8, 1006.9, 1007, 1007.1, 
    1007, 1007.1, 1007.4, 1007.4, 1007.3, 1007.2, 1007.2, 1007.2, 1006.8, 
    1006.5, 1006.1, 1005.5, 1005.2, 1004.8, 1004.4, 1004.4, 1004, 1003.8, 
    1003.8, 1004, 1004.3, 1004.9, 1005, 1005.8, 1006.3, 1006.8, 1007.1, 
    1007.6, 1007.9, 1008.5, 1009.1, 1009.7, 1010.3, 1010.9, 1011.4, 1011.8, 
    1012.4, 1012.8, 1013, 1013.5, 1013.9, 1014.4, 1014.5, 1014.6, 1014.6, 
    1014.5, 1014.3, 1014.3, 1014.3, 1014.3, 1014.3, 1014.3, 1014.2, 1014.2, 
    1014.2, 1014.3, 1014.4, 1014.4, 1014.4, 1014.6, 1014.9, 1015.3, 1015.5, 
    1015.9, 1015.9, 1016, 1016.5, 1016.7, 1016.7, 1016.5, 1016.5, 1016.4, 
    1016.1, 1016, 1016.2, 1016, 1015.6, 1015.2, 1015, 1014.5, 1013.8, 1012.9, 
    1012.3, 1011.3, 1010, 1009.1, 1008.1, 1007.4, 1006.8, 1006.4, 1005.9, 
    1005.5, 1005.3, 1005, 1004.8, 1005, 1005, 1005.2, 1005.6, 1006, 1006.5, 
    1007.2, 1008, 1009.1, 1009.7, 1010.1, 1011.1, 1011.8, 1012.2, 1012.8, 
    1013.3, 1013.6, 1013.6, 1013.8, 1013.4, 1013.3, 1012.8, 1012.1, 1011.1, 
    1011.5, 1011.3, 1011.1, 1010.9, 1010.7, 1010.7, 1010.8, 1010.7, 1010.4, 
    1010.4, 1010.5, 1010.6, 1011, 1011.3, 1011.8, 1012.5, 1012.9, 1013.4, 
    1013.7, 1013.9, 1013.9, 1013.8, 1013.4, 1013.1, 1012.9, 1012.8, 1012.8, 
    1012.6, 1012.7, 1012.6, 1012.4, 1012.2, 1011.9, 1011.7, 1011.4, 1011.1, 
    1010.7, 1010.3, 1010, 1009.6, 1009.2, 1008.9, 1008.4, 1007.9, 1007.4, 
    1006.9, 1006, 1005.2, 1004.5, 1003.8, 1003.5, 1003, 1002.2, 1001.9, 
    1001.6, 1001, 1000.7, 1000.9, 1001.1, 1001.1, 1000.9, 1001.3, 1001.6, 
    1001.8, 1002, 1002, 1001.8, 1002.3, 1002.4, 1002.4, 1002.8, 1003.1, 
    1003.6, 1003.8, 1004.1, 1004.6, 1005.3, 1005.5, 1005.7, 1006, 1006.3, 
    1006.8, 1007.4, 1007.4, 1007.3, 1007.1, 1007.3, 1007.2, 1007.6, 1007.2, 
    1007, 1006.8, 1006.4, 1005.9, 1005.8, 1006.1, 1006.2, 1006.4, 1006.8, 
    1006.9, 1007.5, 1007.9, 1008.7, 1009.6, 1010.4, 1011.2, 1012.3, 1013.3, 
    1014.3, 1015.2, 1016, 1016.8, 1017.3, 1017.9, 1018.6, 1019.2, 1019.5, 
    1019.8, 1019.9, 1020.1, 1020.3, 1020.5, 1020.7, 1020.7, 1020.6, 1020.7, 
    1021.1, 1021, 1020.5, 1020.4, 1020.2, 1019.9, 1019.5, 1018.9, 1018, 
    1017.4, 1016.8, 1016.3, 1015.7, 1014.9, 1014.2, 1013.7, 1012.9, 1011.8, 
    1010.8, 1010.2, 1009.6, 1008.7, 1007.9, 1007.5, 1006.7, 1005.9, 1005.1, 
    1004.1, 1003.1, 1002.2, 1001.6, 1001.1, 1000.9, 1000.9, 1001.2, 1002, 
    1002.5, 1002.8, 1003.3, 1003.4, 1003.8, 1004.2, 1004.6, 1005.3, 1005.8, 
    1006.4, 1006.8, 1007.6, 1008.3, 1008.6, 1009.1, 1009.5, 1009.7, 1009.9, 
    1009.8, 1009.7, 1009.6, 1009.5, 1009.6, 1009.7, 1010.4, 1010.6, 1010.8, 
    1011, 1011.1, 1010.9, 1011.1, 1011.1, 1011, 1010.8, 1010.8, 1010.6, 
    1010.5, 1010.3, 1009.9, 1009.3, 1008.9, 1008.2, 1007.8, 1007.3, 1006.9, 
    1006.7, 1006.2, 1005.9, 1005.7, 1005.3, 1005.1, 1004.8, 1004.5, 1004.1, 
    1003.5, 1002.9, 1002.1, 1001.5, 1000.9, 1000, 998.9, 998, 997.3, 996.7, 
    996.7, 996.4, 996.2, 995.8, 995.3, 994.5, 993.2, 992.3, 991.2, 990.6, 
    990, 989.4, 988.8, 988.4, 987.5, 986.7, 986.1, 984.9, 984.2, 983.3, 983, 
    982.5, 981.6, 981.3, 980.5, 979.6, 979.3, 979.1, 978.9, 978.9, 979.4, 
    979.8, 980.6, 981, 981.7, 982.3, 982.9, 983.4, 984.3, 985, 985.7, 986.5, 
    987.4, 988.4, 989.5, 990.4, 991, 991.7, 992.4, 993, 993.4, 994, 994.4, 
    994.6, 994.8, 995.2, 995.5, 995.7, 995.7, 995.5, 995.5, 994.9, 994.7, 
    994.2, 994.1, 993.6, 993.5, 993.2, 993, 992.6, 992.3, 991.9, 991.4, 991, 
    990.7, 990.5, 990.5, 990.5, 990.8, 990.8, 991, 991.2, 991.2, 991.2, 
    991.2, 991.2, 991.2, 991.7, 991.7, 991.8, 991.9, 992.1, 992.4, 992.5, 
    992.5, 992.3, 992.3, 992, 991.8, 991.6, 991.7, 991.4, 991.3, 991.1, 
    991.1, 991, 990.8, 990.7, 990.6, 990.7, 990.8, 990.7, 990.8, 990.9, 991, 
    991, 991, 991, 990.9, 991.1, 991.3, 991.3, 991.5, 991.8, 992.2, 992.7, 
    993.2, 994, 994.6, 995.2, 995.7, 996.3, 996.9, 997.8, 998.6, 999.3, 
    999.9, 1000.4, 1001.1, 1001.8, 1002.4, 1002.8, 1003.5, 1004.2, 1004.7, 
    1005, 1005.4, 1005.8, 1006.2, 1006.5, 1006.9, 1007.2, 1007.5, 1007.6, 
    1007.8, 1008.1, 1008.3, 1008.3, 1008.4, 1008.4, 1008.5, 1008.7, 1008.6, 
    1008.5, 1008.6, 1008.6, 1008.7, 1008.8, 1008.7, 1008.6, 1008.7, 1008.9, 
    1009, 1009, 1009, 1009, 1009.1, 1009.3, 1009.5, 1009.7, 1009.8, 1009.8, 
    1010.2, 1010.3, 1010.5, 1010.7, 1011, 1011.2, 1011.3, 1011.5, 1012, 
    1012.2, 1011.4, 1012.7, 1012.9, 1013.1, 1013.4, 1013.7, 1013.6, 1013.5, 
    1013.6, 1013.7, 1013.8, 1014.1, 1013.8, 1013.7, 1013.7, 1013.6, 1013.5, 
    1013.4, 1013.2, 1012.9, 1012.6, 1012.3, 1012.2, 1012.3, 1012, 1011.6, 
    1011.3, 1011.1, 1010.6, 1010.4, 1010.1, 1009.9, 1009.7, 1009.5, 1009.3, 
    1009, 1008.8, 1008.2, 1007.8, 1007.5, 1007.3, 1006.9, 1006.7, 1006.5, 
    1006.2, 1006, 1005.6, 1005.7, 1005.6, 1005.7, 1005.4, 1005.5, 1005.4, 
    1005.7, 1005.9, 1006.2, 1006.6, 1007.1, 1007.6, 1007.9, 1008.4, 1008.9, 
    1009.2, 1009.6, 1010.1, 1010.4, 1010.7, 1011.2, 1011.7, 1012.1, 1012.5, 
    1012.8, 1013.1, 1013.4, 1013.4, 1013.9, 1014.2, 1014.4, 1014.8, 1015.3, 
    1015.7, 1016.1, 1016.3, 1016.5, 1016.7, 1016.6, 1016.9, 1017, 1017, 
    1017.2, 1017.5, 1017.7, 1017.9, 1018.1, 1018.3, 1018.5, 1018.6, 1018.6, 
    1018.7, 1019, 1018.9, 1018.8, 1019.2, 1019.5, 1019.6, 1020, 1019.9, 
    1019.8, 1019.9, 1019.9, 1019.8, 1019.8, 1020.2, 1020.3, 1020.7, 1020.8, 
    1020.8, 1020.7, 1020.6, 1020.7, 1020.7, 1020.6, 1020.4, 1020.2, 1019.9, 
    1019.7, 1019.7, 1019.7, 1019.4, 1019, 1018.8, 1018.6, 1018.4, 1017.9, 
    1017.6, 1017.3, 1017.1, 1017, 1017, 1016.9, 1016.8, 1016.4, 1016.3, 
    1016.1, 1015.6, 1015.1, 1015, 1014.9, 1014.9, 1015, 1015, 1014.5, 1015, 
    1014.6, 1014.4, 1014.6, 1014.8, 1014.8, 1014.7, 1014.7, 1014.6, 1014.7, 
    1015.1, 1015.3, 1014.9, 1015, 1015.4, 1015.3, 1015.4, 1015.5, 1015.4, 
    1015.6, 1015.8, 1016.2, 1016.3, 1016.6, 1016.7, 1016.7, 1016.7, 1016.7, 
    1016.8, 1017, 1016.8, 1016.9, 1016.9, 1017, 1017.2, 1017.3, 1017.1, 
    1016.8, 1016.6, 1016.8, 1016.6, 1016.2, 1015.9, 1015.5, 1015.1, 1014.8, 
    1014.7, 1014.3, 1014, 1013.7, 1012.5, 1011.7, 1011.1, 1009.9, 1008.7, 
    1007.4, 1006.1, 1004.8, 1004, 1003.2, 1002.2, 1001.1, 999.9, 998.7, 998, 
    997.2, 996.3, 995.3, 994.2, 993, 992.1, 991.5, 991, 990.7, 990.8, 990.9, 
    991, 991.3, 991.5, 991.8, 992.5, 992.7, 993.3, 994.3, 995.5, 996.3, 
    997.1, 998.3, 999.5, 1000.9, 1002.1, 1002.9, 1003.8, 1004.6, 1005.8, 
    1006.9, 1008, 1008.8, 1009.5, 1009.9, 1010.7, 1011.4, 1012.3, 1012.8, 
    1013.3, 1014, 1014.8, 1015.3, 1015.8, 1016.3, 1016.6, 1016.9, 1017.1, 
    1017.5, 1017.7, 1017.9, 1018.2, 1018.3, 1018.5, 1018.5, 1018.6, 1018.5, 
    1018.4, 1018, 1018.2, 1018.2, 1018.2, 1018, 1017.7, 1017.4, 1017.1, 
    1016.8, 1016.4, 1016, 1015.3, 1014.1, 1013.9, 1013.7, 1013.2, 1012.3, 
    1011.3, 1010.5, 1009.8, 1008.9, 1008.1, 1007.7, 1007.2, 1006.4, 1006, 
    1005, 1005, 1004.7, 1004.3, 1004.2, 1004.1, 1004.1, 1004.3, 1004.6, 
    1004.8, 1004.8, 1004.8, 1004.8, 1004.7, 1004.5, 1004, 1003.1, 1002.2, 
    1001.2, 1000.2, 998.9, 997.2, 995.5, 994, 991.8, 990.6, 989.9, 988.8, 
    988.2, 988.7, 989.7, 990.2, 991.1, 993, 994.1, 995.7, 997.6, 1000.2, 
    1001.6, 1002.5, 1002.7, 1003.9, 1004.5, 1005.1, 1005.7, 1006, 1006.1, 
    1006.2, 1006.3, 1006.6, 1006.9, 1007.1, 1007.6, 1008.3, 1008.9, 1009.7, 
    1010.4, 1010.8, 1011, 1011.5, 1011.6, 1012, 1012.2, 1012.2, 1012.3, 
    1012.4, 1012.7, 1013.2, 1013.1, 1013.2, 1013.1, 1013.3, 1013.5, 1013.9, 
    1014.2, 1014.7, 1015.3, 1015.6, 1015.6, 1015.5, 1015.1, 1014.7, 1013.7, 
    1012.9, 1011.4, 1009.7, 1007.8, 1006.8, 1006.4, 1007.1, 1007.9, 1008.3, 
    1008.6, 1008.4, 1008.8, 1009.1, 1009.3, 1009.6, 1010.1, 1011.1, 1011.7, 
    1011.8, 1012.1, 1012.4, 1012.6, 1012.5, 1012, 1011.5, 1011, 1010.5, 
    1010.6, 1010.6, 1010.9, 1011.4, 1011.8, 1012.1, 1012.7, 1013.3, 1014.2, 
    1014.9, 1015.6, 1016.2, 1016.8, 1017.4, 1017.7, 1018.4, 1018.7, 1019.1, 
    1019.4, 1019.1, 1019, 1019, 1018.5, 1018.5, 1018, 1017.6, 1017.4, 1017.1, 
    1016.7, 1016.5, 1016.6, 1016.4, 1016.4, 1016.5, 1016.5, 1016.4, 1016.4, 
    1016.7, 1016.9, 1017, 1016.9, 1016.8, 1016.7, 1016.7, 1016.4, 1016.3, 
    1016.4, 1016.5, 1016.5, 1016.7, 1016.8, 1017, 1017, 1017.1, 1017.2, 
    1017.2, 1017, 1016.7, 1016.5, 1016.3, 1016.2, 1016.2, 1016.2, 1016.2, 
    1016.4, 1016.5, 1016.5, 1016.5, 1016.3, 1016.4, 1017.7, 1016.4, 1016.4, 
    1016.4, 1016.7, 1016.9, 1017.1, 1017.1, 1017.4, 1017.4, 1017.4, 1017.6, 
    1017.9, 1018.2, 1018.3, 1018.4, 1018.5, 1018.8, 1019, 1019.2, 1019.3, 
    1019.2, 1019.2, 1019.4, 1019.3, 1019.3, 1019.2, 1019.2, 1019.4, 1019.4, 
    1019.3, 1019.1, 1018.7, 1018.3, 1017.7, 1017.2, 1016.9, 1016.4, 1015.8, 
    1015.2, 1014.4, 1013.7, 1013, 1012.2, 1011.2, 1010.4, 1009.7, 1008.6, 
    1007.9, 1007.6, 1007.2, 1007, 1006.9, 1007.1, 1007.2, 1007.4, 1007.2, 
    1007.1, 1007.1, 1006.8, 1006.6, 1006.2, 1006, 1005.6, 1005.7, 1005.7, 
    1005.4, 1005, 1004.8, 1004.4, 1004.1, 1003.9, 1003.8, 1003.6, 1003.3, 
    1003.3, 1003.4, 1003.5, 1003.7, 1003.6, 1003.6, 1003.5, 1003.5, 1003.6, 
    1003.5, 1003.6, 1003.3, 1003.1, 1003.4, 1003.6, 1003.4, 1003.1, 1003.2, 
    1003.2, 1002.9, 1002.6, 1002.4, 1001.6, 1002.2, 1001.7, 1001.5, 1001.4, 
    1000.9, 1000.4, 1000.1, 999.7, 999.1, 998.3, 997.7, 997.4, 996.6, 996, 
    995.2, 994.3, 993.9, 993.1, 992, 991.4, 1001, 990.5, 990, 989.3, 988.9, 
    988.4, 988.4, 988.1, 988.3, 988.3, 988.6, 988.5, 988.9, 988.8, 988.9, 
    989.1, 989.2, 989.3, 989.6, 989.7, 989.7, 990.1, 990.4, 989.8, 989.8, 
    990, 989.9, 989.7, 989.4, 989.5, 989.7, 989.5, 989.6, 989.4, 989.4, 989, 
    989.3, 989.3, 989.5, 990, 990.4, 990.9, 991, 991.2, 991.1, 991.5, 991.7, 
    991.8, 991.8, 992.1, 992.2, 992.5, 992.8, 993.3, 994.2, 994.8, 995.3, 
    995.8, 996.4, 996.9, 997.5, 998.1, 998.9, 999.4, 1000, 1000.6, 1001.4, 
    1002.4, 1003.3, 1004.2, 1005.1, 1006, 1006.9, 1008, 1009, 1010.2, 1011.2, 
    1012, 1012.8, 1013.7, 1014.1, 1014.3, 1014.3, 1013.9, 1013.9, 1014.5, 
    1014.5, 1015.1, 1015.7, 1016.5, 1017.1, 1018.6, 1019.9, 1021.4, 1022.6, 
    1023.6, 1024.1, 1024.1, 1024.5, 1024.5, 1024.1, 1023.8, 1023.5, 1023.2, 
    1022.8, 1022.2, 1021.2, 1020.1, 1019.4, 1018.9, 1018.6, 1018.1, 1018.2, 
    1017.6, 1016.9, 1015.9, 1015.1, 1014.6, 1013.9, 1012.9, 1011.8, 1010.5, 
    1009, 1007.4, 1006.3, 1005.7, 1005.1, 1004.9, 1005.1, 1005.3, 1005.8, 
    1006.2, 1006.2, 1006.3, 1006.9, 1007.9, 1008.7, 1009.9, 1011.1, 1012.3, 
    1013.6, 1015, 1016.2, 1017.4, 1018.9, 1020.4, 1022.2, 1022.9, 1023.6, 
    1024.7, 1025.5, 1026, 1026.9, 1027.5, 1027.5, 1027.4, 1027.8, 1027.5, 
    1027.5, 1027.2, 1026.9, 1026.4, 1025.3, 1024.3, 1023.2, 1022, 1020.8, 
    1019.5, 1018.3, 1016.9, 1015.6, 1014.8, 1013.4, 1012.1, 1011.3, 1010.7, 
    1010.1, 1009.8, 1010.1, 1011.9, 1012.2, 1012.6, 1012.9, 1012.4, 1012.3, 
    1012.3, 1013.9, 1014.5, 1016.3, 1017.4, 1018.6, 1019.6, 1020.7, 1021.5, 
    1022.6, 1023.4, 1024, 1024.4, 1024.7, 1025, 1025.5, 1026, 1026.6, 1026.7, 
    1026.8, 1027.2, 1027.5, 1027.6, 1027.9, 1028.3, 1028.7, 1028.9, 1029, 
    1029.3, 1029.5, 1029.6, 1029.6, 1029.7, 1029.6, 1029.4, 1028.9, 1029, 
    1028.8, 1028.7, 1028.3, 1027.9, 1027.3, 1026.9, 1026.3, 1025.8, 1025.5, 
    1024.9, 1024.7, 1024.3, 1023.8, 1023.3, 1023.1, 1022.3, 1021.8, 1021.3, 
    1020.9, 1020.1, 1019.5, 1019.3, 1018.6, 1018.5, 1018.2, 1018.3, 1018.3, 
    1018.2, 1017.9, 1017.9, 1018, 1017.7, 1017.7, 1017.8, 1017.8, 1017.7, 
    1017.6, 1017.5, 1017.4, 1017.1, 1016.8, 1016.2, 1015.6, 1015, 1014.2, 
    1013.3, 1012.4, 1012, 1011.3, 1010.8, 1009.8, 1008.9, 1008, 1007.5, 
    1007.2, 1007.3, 1007.4, 1007.6, 1008, 1008.7, 1009.3, 1009.8, 1010.4, 
    1010.9, 1011.5, 1011.9, 1012.6, 1012.8, 1013.1, 1013.3, 1013.8, 1014.1, 
    1014.8, 1015.3, 1015.7, 1016, 1016.3, 1016.5, 1016.6, 1016.7, 1016.8, 
    1017.1, 1017.3, 1017.6, 1017.9, 1018.1, 1018.3, 1018.4, 1018.7, 1018.9, 
    1019.2, 1019.4, 1019.7, 1019.6, 1020, 1020.4, 1020.7, 1020.9, 1021.1, 
    1021.4, 1021.5, 1021.8, 1022.3, 1022.3, 1022.3, 1022.3, 1022.5, 1022.5, 
    1022.5, 1022.5, 1022.4, 1022.5, 1022.3, 1021.9, 1021.2, 1020.6, 1019.7, 
    1018.9, 1018.1, 1017.2, 1016.2, 1015.1, 1014.3, 1013.5, 1012.8, 1012, 
    1011.2, 1010.8, 1010.1, 1009.2, 1008.7, 1008.3, 1007.6, 1006.8, 1006.6, 
    1006, 1005.4, 1005.1, 1004.3, 1003.6, 1002.8, 1001.8, 1001, 1000.5, 
    1000.3, 1001.1, 1001.4, 1002, 1001.8, 1001.7, 1003, 1004.3, 1005.1, 1005, 
    1005.4, 1006.2, 1006.4, 1007.4, 1008.3, 1008.8, 1009.4, 1009.6, 1010.9, 
    1011.9, 1012.7, 1013.6, 1014.2, 1014.6, 1015, 1015.5, 1016, 1016.4, 
    1016.5, 1016.5, 1016.3, 1016.5, 1016.2, 1016.1, 1015.9, 1015.5, 1015.4, 
    1015.3, 1015.3, 1015.3, 1015.5, 1015.7, 1015.8, 1015.6, 1015.7, 1016, 
    1016, 1016, 1016.1, 1016.3, 1016.2, 1016.3, 1016.4, 1016.3, 1016.3, 
    1016.2, 1016.2, 1016.1, 1016, 1015.8, 1015.7, 1016, 1016.1, 1016.2, 
    1016.2, 1016, 1016, 1016, 1016, 1016.3, 1016.3, 1016.3, 1016.6, 1016.8, 
    1016.9, 1016.9, 1016.8, 1016.5, 1016.6, 1016.6, 1016.4, 1016.3, 1016.6, 
    1016.4, 1016.2, 1016.2, 1016.2, 1016.2, 1016.3, 1016.2, 1016.1, 1015.8, 
    1015.8, 1015.7, 1015.4, 1015.4, 1015.3, 1015.3, 1015.4, 1015.4, 1015.3, 
    1015, 1014.9, 1014.7, 1014.7, 1014.6, 1014.4, 1014.4, 1014.6, 1014.5, 
    1014.5, 1014.2, 1014.5, 1014.6, 1014.1, 1014, 1014.1, 1014.1, 1013.9, 
    1013.9, 1014.1, 1014.4, 1014.8, 1015.1, 1015.2, 1014.9, 1014.5, 1014.2, 
    1013.9, 1013.7, 1013.6, 1013.2, 1012.8, 1012.4, 1011.4, 1011.3, 1010.1, 
    1009.8, 1009.5, 1008.4, 1008.3, 1008.2, 1007.9, 1008.1, 1008.2, 1009.2, 
    1009.5, 1010.2, 1010.5, 1011, 1011.8, 1012.3, 1013.4, 1014.2, 1015, 
    1015.5, 1016.5, 1017.3, 1017.9, 1018.2, 1018.2, 1018.2, 1018.6, 1018.6, 
    1018.4, 1018.5, 1018.5, 1019.1, 1019.5, 1020.4, 1021.2, 1022.3, 1023.1, 
    1023.8, 1024.6, 1025.4, 1026.1, 1026.6, 1027, 1027.2, 1027.7, 1028, 
    1028.1, 1028, 1029.3, 1028, 1028, 1028, 1027.9, 1028, 1028.2, 1028.5, 
    1028.6, 1028.6, 1028.5, 1029, 1029.2, 1029, 1028.9, 1029.1, 1029, 1029.1, 
    1029, 1029.3, 1029.7, 1029.5, 1029.8, 1029.8, 1029.4, 1029.4, 1029, 
    1028.6, 1028.4, 1028.1, 1027.6, 1027.4, 1027.3, 1027.2, 1027, 1026.9, 
    1026.3, 1025.8, 1025.5, 1024.9, 1024.2, 1023.5, 1023, 1022.4, 1021.4, 
    1020.7, 1020.1, 1019.5, 1018.8, 1018.2, 1017.4, 1016.8, 1016, 1015.3, 
    1014.7, 1014.1, 1013.6, 1013.2, 1012.8, 1012.4, 1012.1, 1011.7, 1011.3, 
    1010.9, 1010.7, 1010.4, 1010.3, 1010.4, 1010.3, 1010.4, 1010.3, 1010, 
    1009.8, 1009.6, 1009.2, 1009.1, 1009, 1009, 1008.8, 1008.9, 1008.9, 
    1008.7, 1008.6, 1008.4, 1008.4, 1008.3, 1008, 1007.7, 1007.4, 1007, 
    1006.6, 1006.7, 1006.7, 1006.9, 1007.1, 1007.2, 1007.4, 1007.4, 1007.3, 
    1007.5, 1007.6, 1007.8, 1008, 1008.2, 1008.7, 1009.1, 1009.3, 1009.4, 
    1009.7, 1009.9, 1009.7, 1009.6, 1009.7, 1009.5, 1009.1, 1009.1, 1009.1, 
    1009.3, 1009.5, 1009.5, 1009.5, 1009.7, 1010, 1010.2, 1010.3, 1010.5, 
    1010.8, 1011, 1011.5, 1012.1, 1012.5, 1012.5, 1013.1, 1013.3, 1013.4, 
    1014, 1014.6, 1015.4, 1015.7, 1016.9, 1017.3, 1017.6, 1018, 1018.4, 
    1018.6, 1018.9, 1019.5, 1019.8, 1020.9, 1021.4, 1022.1, 1022.7, 1023.4, 
    1024.1, 1024.5, 1025.5, 1026.3, 1026.8, 1027.2, 1027.7, 1027.9, 1028.2, 
    1028.3, 1028.7, 1029, 1029.3, 1029.6, 1030, 1030.4, 1030.9, 1031.1, 
    1031.4, 1031.6, 1031.8, 1032, 1032.3, 1032.4, 1032.7, 1032.8, 1033, 
    1033.2, 1033.2, 1033.4, 1033.4, 1033.5, 1033.3, 1033.2, 1033.3, 1033.5, 
    1033.5, 1033.6, 1033.4, 1033.4, 1033.2, 1033, 1032.8, 1032.5, 1032.3, 
    1032.2, 1032.1, 1032.1, 1032.1, 1032.2, 1032.1, 1032, 1032, 1032.1, 1032, 
    1031.8, 1031.9, 1032, 1032.2, 1032.3, 1032.4, 1032.4, 1032.4, 1032.3, 
    1032.3, 1032, 1031.9, 1031.9, 1031.9, 1031.9, 1031.5, 1031.6, 1031.6, 
    1031.6, 1031.4, 1031.1, 1030.9, 1030.6, 1030.2, 1029.9, 1029.6, 1029.2, 
    1029, 1028.6, 1028.3, 1028.2, 1027.9, 1027.6, 1027.3, 1027, 1026.8, 
    1026.7, 1026.5, 1026.2, 1026.2, 1026.1, 1026, 1026.2, 1026.3, 1026.3, 
    1026.3, 1026.4, 1026.6, 1026.8, 1027, 1026.8, 1027, 1027.3, 1027.5, 
    1027.5, 1027.7, 1027.8, 1028, 1028.1, 1028.3, 1028.4, 1028.4, 1028.4, 
    1028.6, 1028.7, 1029, 1029.3, 1029.4, 1029.4, 1029.5, 1029.5, 1029.5, 
    1029.6, 1029.6, 1029.7, 1029.7, 1029.8, 1029.6, 1029.6, 1029.6, 1029.4, 
    1029.1, 1028.9, 1028.7, 1028.4, 1028.3, 1027.8, 1027.3, 1026.9, 1026.5, 
    1026.3, 1025.9, 1025.4, 1025, 1024.4, 1023.9, 1023.5, 1023, 1022.6, 
    1022.2, 1022.1, 1021.9, 1021.8, 1021.5, 1021.7, 1021.5, 1021.7, 1021.8, 
    1021.9, 1022.1, 1022.4, 1022.6, 1022.9, 1023.3, 1023.4, 1023.3, 1023.4, 
    1023.5, 1023.4, 1023.4, 1023.3, 1023.4, 1023.1, 1022.8, 1022.4, 1022.1, 
    1021.4, 1020.7, 1020, 1019.1, 1018.5, 1017.8, 1017.2, 1016.4, 1015.6, 
    1015.1, 1014.7, 1014.2, 1013.5, 1013, 1012.3, 1011.7, 1010.8, 1010.1, 
    1009.3, 1008.8, 1008, 1007.3, 1006.6, 1005.9, 1005, 1004.3, 1003.5, 
    1002.8, 1001.8, 1001.2, 1000.5, 999.6, 998.7, 997.9, 997, 996.5, 995.8, 
    995.3, 994.6, 993.9, 993.1, 992, 991.2, 990.3, 989.8, 989, 988.7, 987.4, 
    986.6, 986, 985.1, 984.3, 983.8, 983.7, 983.7, 984.5, 985.8, 987.3, 
    989.3, 991.1, 992.3, 993.8, 995.8, 997.3, 998, 999.2, 1000.5, 1001, 
    1001.8, 1002.4, 1002.7, 1003.3, 1003.4, 1003.7, 1004, 1004.2, 1004.6, 
    1005.1, 1005.8, 1006.2, 1006.6, 1007.2, 1007.8, 1008.7, 1009.7, 1010.7, 
    1011.8, 1012.4, 1012.5, 1013.5, 1014.2, 1014.7, 1015.2, 1015.6, 1016, 
    1016.6, 1017.1, 1017.7, 1017.7, 1018, 1018.3, 1018.4, 1018.6, 1019, 
    1019.2, 1019.7, 1020.2, 1020.5, 1021, 1021.2, 1021.5, 1021.7, 1022, 
    1022.1, 1022.1, 1022.2, 1022.1, 1022, 1021.5, 1021.4, 1021.3, 1021.3, 
    1021, 1020.5, 1019.8, 1019.7, 1019.2, 1018.9, 1018.4, 1017.9, 1017.9, 
    1017.9, 1017.7, 1017.3, 1017.1, 1016.7, 1016.1, 1016.1, 1015.8, 1015.5, 
    1014.9, 1014.7, 1014.5, 1014.1, 1013.8, 1013.7, 1013.3, 1012.6, 1012.1, 
    1011.7, 1011.1, 1010.9, 1010.2, 1009.6, 1009.5, 1009.3, 1009, 1008.7, 
    1008.3, 1007.8, 1007.6, 1007.4, 1007.4, 1007.1, 1007, 1006.9, 1006.9, 
    1006.4, 1006.1, 1006, 1005.7, 1005.5, 1005.2, 1005, 1004.6, 1004.2, 
    1003.8, 1003.5, 1003.3, 1003.2, 1002.9, 1002.6, 1002.5, 1002.3, 1001.8, 
    1001.8, 1001.6, 1001.2, 1000.8, 1000.3, 999.7, 999.1, 998.5, 997.6, 
    996.4, 995.6, 994.6, 994, 992.4, 991.8, 990.9, 989.7, 988.3, 986.3, 
    983.6, 981.6, 979.5, 977.4, 975.6, 973.8, 972.6, 971.8, 971.4, 970.9, 
    969.4, 969.1, 968.9, 969.1, 969.7, 970.9, 972, 972.9, 973.8, 974.7, 
    974.8, 975.4, 975.9, 976.5, 977.1, 978.2, 979.2, 980.2, 981.1, 981.9, 
    982.7, 983.6, 983.9, 984.4, 984.9, 985, 985.3, 985.1, 985, 984.6, 984.2, 
    983.3, 982.1, 980.7, 979.9, 979.1, 978.4, 977.9, 977.5, 976.9, 976.2, 
    975.5, 975.4, 974.4, 973.9, 973.7, 973.9, 974.2, 975.1, 978.6, 978.6, 
    981.3, 983.8, 986.3, 988.7, 990.8, 992.5, 993.8, 995.4, 996.9, 997.6, 
    998.8, 1000, 1001, 1001.6, 1002.5, 1003.6, 1004.7, 1005.7, 1006.4, 
    1007.4, 1008.2, 1009.1, 1009.9, 1011, 1011.7, 1012.3, 1012.9, 1013.4, 
    1013.7, 1014, 1014.2, 1014.5, 1014.7, 1015, 1015, 1015.2, 1015.3, 1015.3, 
    1015.4, 1015, 1014.9, 1014.7, 1014.7, 1014.7, 1014.5, 1014.2, 1013.8, 
    1013.5, 1013.3, 1013.4, 1013.2, 1013.2, 1012.5, 1012.1, 1011.6, 1011.2, 
    1010.8, 1010.3, 1009.8, 1009.1, 1009, 1008.8, 1008.4, 1008.2, 1008, 
    1007.6, 1007, 1006.5, 1006, 1005.7, 1005.3, 1004.9, 1004.4, 1004.1, 
    1003.7, 1003.5, 1003.3, 1003.3, 1003, 1003, 1003, 1003.2, 1003.3, 1003.5, 
    1003.4, 1003.3, 1003.5, 1003.3, 1003.4, 1003.6, 1003.8, 1004.5, 1004.8, 
    1005.2, 1005.5, 1006.1, 1006.5, 1006.6, 1006.8, 1007, 1007.4, 1007.4, 
    1008.1, 1008.4, 1008.7, 1009.1, 1009.6, 1010.1, 1010.7, 1011, 1011.3, 
    1011.7, 1012, 1012.3, 1012.8, 1013.1, 1013.4, 1013.7, 1014, 1014.3, 
    1014.3, 1014.3, 1014.3, 1014.5, 1014.6, 1014.7, 1014.8, 1014.9, 1015, 
    1015.3, 1015.8, 1015.9, 1016, 1016.3, 1016.4, 1016.4, 1016.4, 1016.4, 
    1016.4, 1016.4, 1016.6, 1016.9, 1016.8, 1016.9, 1016.6, 1016.5, 1016.6, 
    1016.5, 1016.6, 1016.6, 1016.6, 1016.7, 1016.6, 1016.6, 1016.8, 1017.1, 
    1017, 1017.1, 1017.1, 1017, 1017.2, 1017.1, 1016.9, 1017, 1017.2, 1017.3, 
    1017.3, 1017.3, 1017.4, 1017.6, 1017.8, 1017.6, 1017.6, 1017.5, 1017.4, 
    1017.6, 1017.5, 1017.8, 1018.1, 1018.4, 1018.7, 1019, 1020.2, 1018.9, 
    1019, 1018.9, 1018.8, 1018.8, 1018.7, 1018.8, 1018.9, 1019, 1018.8, 
    1018.8, 1018.6, 1018.2, 1017.9, 1017.7, 1017.4, 1017.1, 1016.8, 1016.6, 
    1016.3, 1016.2, 1016.1, 1015.9, 1015.4, 1015, 1014.6, 1014.5, 1014.5, 
    1014.3, 1014.1, 1014.7, 1015.1, 1015.4, 1015.2, 1014.9, 1014.8, 1015, 
    1015.1, 1015, 1015.3, 1015.3, 1015.4, 1015.4, 1015.6, 1015.7, 1015.9, 
    1015.8, 1015.6, 1016, 1015.9, 1016, 1016.1, 1016.4, 1016.3, 1016.8, 
    1016.8, 1016.8, 1017, 1017.4, 1017.6, 1017.8, 1017.6, 1018.5, 1018.8, 
    1018.9, 1019.3, 1019.5, 1019.7, 1019.8, 1020.1, 1020.3, 1020.4, 1020.3, 
    1020.2, 1019.9, 1019.8, 1019.7, 1019.5, 1019.3, 1019.2, 1019, 1018.5, 
    1017.9, 1017.2, 1016.7, 1016.1, 1015.6, 1015.1, 1014.5, 1013.7, 1013.2, 
    1012.6, 1012.2, 1011.6, 1011, 1010.5, 1009.8, 1009.2, 1008.7, 1007.8, 
    1007.3, 1007, 1006.8, 1006.6, 1006.6, 1006.3, 1006.1, 1005.8, 1005.2, 
    1004.9, 1004.6, 1004.5, 1004.1, 1003.9, 1003.6, 1003.3, 1003.5, 1004.2, 
    1004.5, 1004.5, 1004.9, 1005, 1004.9, 1005.4, 1005.7, 1005.9, 1006.1, 
    1006.4, 1006.4, 1006.5, 1006.7, 1006.4, 1006.7, 1007.3, 1007.8, 1008.4, 
    1008.6, 1008.7, 1008.9, 1009.2, 1009.8, 1010.1, 1010.4, 1011, 1011.1, 
    1011.3, 1011.6, 1012, 1012.3, 1012.3, 1012.5, 1012.9, 1013.3, 1013.8, 
    1014.2, 1014.1, 1014.3, 1014.8, 1015, 1015.3, 1015.5, 1015.6, 1016, 
    1016.4, 1016.7, 1017, 1017.5, 1018, 1018.1, 1018.3, 1018.4, 1018.7, 
    1018.9, 1019.2, 1019.6, 1019.7, 1019.9, 1019.9, 1019.8, 1019.8, 1019.8, 
    1019.7, 1019.7, 1019.5, 1019.1, 1019, 1018.8, 1018.6, 1018.4, 1018.1, 
    1017.9, 1017.5, 1017.1, 1016.7, 1016.2, 1015.9, 1015.5, 1015, 1014.5, 
    1014.1, 1013.6, 1013.2, 1012.6, 1011.9, 1011.4, 1011, 1010.6, 1010.2, 
    1009.9, 1009.6, 1009.6, 1009.6, 1009.7, 1009.6, 1009.3, 1009.1, 1008.9, 
    1008.5, 1008.2, 1008.1, 1007.6, 1007.1, 1007.1, 1006.8, 1006.3, 1005.8, 
    1005.4, 1004.9, 1004.2, 1003.8, 1003.3, 1002.9, 1002.8, 1002.5, 1002.1, 
    1001.5, 1001.2, 1000.8, 1000.4, 999.8, 999.1, 998.5, 998.6, 998.5, 998.9, 
    999.2, 999.4, 999.9, 1000.6, 1001.3, 1001.6, 1002.2, 1002.7, 1003.3, 
    1003.6, 1004.2, 1004.3, 1004.5, 1004.8, 1005, 1005.7, 1006.2, 1007, 
    1007.7, 1008.9, 1010, 1010.8, 1011.4, 1012.1, 1013.1, 1013.4, 1013.6, 
    1013.5, 1013.9, 1014.2, 1014.3, 1014, 1013.9, 1013.5, 1013.2, 1012.9, 
    1012.8, 1012.6, 1012.3, 1011.8, 1011.7, 1011.3, 1010.8, 1010.4, 1010, 
    1009.8, 1009.5, 1009.3, 1009, 1008.9, 1008.8, 1009, 1009.2, 1009.1, 
    1009.1, 1009, 1008.8, 1008.8, 1008.8, 1008.8, 1008.7, 1008.8, 1008.5, 
    1008.7, 1008.6, 1008.4, 1008.2, 1007.7, 1007.5, 1007.3, 1006.8, 1006.5, 
    1006, 1005.4, 1004.9, 1004.7, 1004.4, 1003.8, 1003.3, 1003, 1002.5, 
    1001.7, 1001, 1000.3, 999.8, 999.5, 999.4, 999.1, 999.6, 999.9, 1000.3, 
    1000.6, 1000.9, 1001.3, 1002, 1002.5, 1002.7, 1003.2, 1003.9, 1004.6, 
    1005, 1005.4, 1006.3, 1007, 1007.4, 1008.1, 1008.4, 1008.6, 1009.1, 1010, 
    1010.5, 1011.2, 1011.9, 1012.8, 1013.4, 1014, 1014.6, 1015.1, 1015.2, 
    1015.7, 1015.8, 1016.2, 1016.4, 1016.6, 1017.1, 1017.3, 1017.3, 1017.7, 
    1017.7, 1017.7, 1017.5, 1017.6, 1017.7, 1017.7, 1017.8, 1018.1, 1018, 
    1017.7, 1017.7, 1017.3, 1016.9, 1016.6, 1016.2, 1015.8, 1015.4, 1015.2, 
    1014.7, 1014.4, 1013.9, 1013.4, 1012.9, 1012.4, 1012, 1011.5, 1010.9, 
    1010.3, 1009.9, 1009.7, 1009.4, 1009.2, 1009.2, 1008.9, 1008.8, 1008.7, 
    1008.7, 1008.3, 1008.2, 1007.8, 1007.7, 1007.5, 1007.2, 1007.1, 1007.3, 
    1007.1, 1007, 1007.2, 1007, 1006.9, 1006.7, 1006.3, 1006.2, 1006.5, 
    1006.5, 1006.6, 1006.4, 1006.7, 1006.7, 1006.7, 1006.4, 1006.3, 1006.3, 
    1006.4, 1006.6, 1006.9, 1007.1, 1007.4, 1007.6, 1007.8, 1007.9, 1007.8, 
    1008, 1007.9, 1007.9, 1007.8, 1007.9, 1008.2, 1008.1, 1008.2, 1008.1, 
    1008.2, 1008.1, 1008.4, 1008.5, 1008.5, 1008.5, 1008.4, 1008.6, 1008.8, 
    1008.8, 1008.8, 1008.6, 1008.1, 1007.7, 1007.5, 1007.1, 1007, 1006.7, 
    1006.6, 1006.3, 1006.1, 1006.1, 1006, 1005.8, 1005.7, 1005.5, 1005.2, 
    1005, 1004.8, 1004.5, 1004.1, 1003.7, 1003.5, 1003.3, 1002.7, 1002.4, 
    1002.2, 1001.8, 1001.6, 1001.3, 1001.3, 1000.8, 1000.8, 1000.7, 1000.8, 
    1001.1, 1001.5, 1001.5, 1001.3, 1001, 1000.8, 1000.6, 1000.3, 999.5, 
    998.6, 998.2, 997.8, 997.5, 997, 996.4, 995.8, 995.3, 995, 994.8, 994.5, 
    994.2, 994.2, 994.4, 994.9, 995.4, 996.2, 997, 997.5, 998.4, 999.3, 1000, 
    1000.4, 1000.7, 1000.8, 1001.4, 1002, 1002.3, 1002.2, 1001.7, 1001.9, 
    1001.2, 1000.7, 1000.3, 1000, 999.6, 998.9, 998.3, 998, 997.4, 997.1, 
    996.7, 996.2, 996.1, 995.8, 995.4, 995, 994.7, 994.4, 994.1, 993.8, 
    993.5, 993.2, 992.9, 992.8, 992.8, 992.8, 992.8, 992.8, 992.7, 992.8, 
    992.8, 993, 993, 993.2, 993.3, 993.4, 993.9, 994.2, 994.4, 994.5, 994.7, 
    994.9, 995.5, 996.2, 996.8, 997.6, 998, 998.2, 998.5, 999, 998.1, 997.8, 
    997.1, 996.7, 995.9, 994.6, 993, 991.5, 988.8, 986.8, 984.4, 981, 978.7, 
    975.9, 973.1, 970.5, 968.3, 966.1, 965.2, 966.2, 966.4, 966.9, 967.4, 
    967.9, 968.5, 969, 969.8, 970, 970.9, 972.5, 974.2, 975.2, 976, 977.3, 
    978.7, 979.8, 980.9, 981.4, 981.3, 981.4, 981.4, 981.3, 981.2, 981, 
    980.7, 980.5, 979.8, 978.4, 976.5, 974.5, 971.5, 968.7, 966.3, 964.8, 
    964.7, 965, 964.3, 964, 964.4, 964.8, 964.7, 964.9, 964.8, 963.6, 963.2, 
    963.1, 963.6, 964.1, 964.5, 965.2, 965.5, 966, 966.5, 966.5, 966.9, 
    966.7, 966.5, 966.7, 966.9, 966.7, 967.5, 967.9, 968.2, 968.6, 968.4, 
    968.3, 968.3, 968.1, 967.7, 968.2, 968.1, 968.1, 968.5, 968.7, 968.4, 
    968.4, 968.6, 969, 969.1, 969.3, 969.7, 970, 970.7, 971.2, 971.5, 972.2, 
    972.5, 972.8, 973.1, 973.7, 974.1, 974.2, 974.6, 975, 975.2, 975.4, 
    975.6, 975.8, 975.7, 975.7, 975.7, 975.8, 975.9, 976, 976.1, 976.2, 
    976.8, 977.3, 977.5, 977.7, 977.8, 978.3, 978.8, 979.1, 979.2, 979.4, 
    979.7, 979.9, 980.2, 980.6, 980.9, 981.3, 981.4, 981.7, 981.8, 981.9, 
    982, 982.2, 982.4, 982.4, 982.6, 982.7, 983.1, 983.3, 983.1, 982.9, 
    982.9, 982.9, 982.7, 982.2, 981.8, 981.4, 981.2, 981.4, 981, 980.6, 
    980.3, 980.1, 979.8, 979.4, 979.1, 978.9, 978.8, 978.9, 978.8, 979.1, 
    979.8, 980, 980, 979.8, 979.8, 980.2, 980.3, 981.4, 982.5, 983.8, 985.2, 
    986.8, 988.4, 989.6, 990.8, 992.2, 993.6, 994.6, 996, 997.4, 998.8, 
    999.5, 1000.8, 1002.4, 1003.5, 1004.7, 1005.4, 1006.3, 1007.5, 1008.3, 
    1008.8, 1009, 1009.4, 1009.9, 1010.6, 1011.2, 1011.8, 1012.3, 1012.5, 
    1012.6, 1012.8, 1012.8, 1012.6, 1012.5, 1011.8, 1011, 1009.6, 1008.1, 
    1006.4, 1004.5, 1002.9, 1000.7, 997.8, 995.7, 993.4, 991.4, 989, 986.9, 
    985.3, 983.8, 983.1, 982.3, 982.3, 981.4, 982.1, 981.9, 983, 983.6, 
    984.8, 985.9, 987.2, 988.4, 989.3, 990.1, 990.9, 991.8, 992.1, 992.7, 
    994.1, 994.6, 995.9, 996.9, 997.7, 998.8, 999.5, 1000.4, 1000.7, 1001, 
    1001.3, 1001.6, 1001.7, 1001.3, 1000.9, 1001.3, 1001.4, 1002, 1002.6, 
    1002.5, 1002.6, 1002.4, 1002.8, 1002.3, 1002.6, 1003.2, 1003.7, 1004.4, 
    1005.1, 1005.5, 1005.9, 1006.4, 1006.4, 1006.8, 1007.3, 1007.8, 1008.2, 
    1008.5, 1009.2, 1009.9, 1010.7, 1011.3, 1012.4, 1013, 1014, 1014.7, 
    1015.9, 1016.7, 1017, 1017.6, 1018, 1019, 1019.7, 1020.5, 1021.2, 1021.3, 
    1021.7, 1021.9, 1022.1, 1022.2, 1022.5, 1022.6, 1022.6, 1022.5, 1022.6, 
    1023, 1023, 1023, 1022.9, 1022.6, 1022.5, 1022.5, 1022.5, 1022.5, 1022.4, 
    1022.6, 1022.5, 1022.5, 1022.2, 1021.9, 1021.4, 1021.2, 1020.9, 1020.5, 
    1020, 1019.4, 1019.2, 1019, 1018.8, 1018.8, 1018.4, 1018.2, 1017.6, 
    1017.3, 1017, 1016.5, 1016.3, 1016.1, 1015.7, 1015.7, 1015.2, 1015.3, 
    1015.4, 1015.3, 1015.2, 1015.5, 1015.7, 1015.7, 1015.7, 1015.8, 1016.1, 
    1016.4, 1016.9, 1017.1, 1017.2, 1017.6, 1017.9, 1018.1, 1018.3, 1017.9, 
    1018.4, 1018.2, 1018, 1018.1, 1018.5, 1018.6, 1018.5, 1018.6, 1018.4, 
    1017.9, 1017.5, 1017.3, 1016.9, 1016.5, 1016, 1015.8, 1015.1, 1014.1, 
    1013.7, 1012.9, 1012.1, 1011.2, 1010.7, 1010.4, 1009.6, 1009.2, 1008.9, 
    1008.8, 1008.6, 1008.9, 1008.6, 1007.9, 1007.1, 1006.2, 1005, 1003.5, 
    1001.6, 999.5, 997.9, 997, 995.7, 994.1, 992.4, 991, 989.9, 988.5, 987.8, 
    987.3, 988, 988.7, 988.4, 988.3, 989.1, 989.7, 989.8, 990.1, 990.5, 
    990.6, 990.8, 991.4, 991.5, 991.3, 991.2, 991.1, 990.9, 990.3, 989.8, 
    988.7, 987.9, 986.8, 986, 985.7, 984.6, 984.7, 984.9, 985, 984.8, 985.7, 
    986.1, 986.5, 986.9, 987.1, 987.5, 987.8, 987.7, 988.6, 988.9, 989.4, 
    989.8, 990.1, 990.6, 990.9, 990.9, 991, 991.5, 991.9, 992, 992.3, 992.8, 
    993.6, 993.9, 994.2, 994.2, 994.2, 994.3, 994.3, 994.3, 994.1, 993.9, 
    993.4, 993.3, 993.3, 993.4, 993.4, 993.4, 993.2, 993, 993, 992.9, 992.7, 
    992.7, 993.1, 993.1, 993.1, 993.6, 993.9, 994, 994.3, 994.7, 994.9, 
    994.5, 994.9, 995.3, 995.5, 995.6, 995.7, 996, 996.4, 996.5, 996.5, 
    996.9, 997, 997.1, 997, 997.2, 997, 996.9, 996.8, 997.1, 997, 996.8, 
    996.9, 996.8, 996.8, 996.8, 996.7, 996.5, 996.1, 996.1, 995.8, 995.7, 
    995.9, 995.8, 995.4, 994.9, 994.7, 994.2, 993.6, 993.1, 993, 992.4, 
    992.3, 991.9, 991.5, 991.2, 990.8, 990.2, 989.7, 989.3, 988.6, 988.1, 
    987.5, 987, 986.5, 986.3, 986, 985.7, 985.3, 985, 985, 985.2, 985.3, 
    985.3, 985.5, 985.8, 986, 986.5, 987, 987.5, 987.8, 988.5, 988.7, 989.3, 
    989.6, 990.1, 990.4, 990.6, 991, 991.5, 991.9, 992.5, 992.8, 992.9, 
    993.1, 993.3, 993.2, 993, 993.3, 993.5, 994, 994.4, 994.7, 994.9, 995.3, 
    995.3, 995.3, 995.4, 995.4, 995.4, 995.4, 995.3, 995.4, 995.6, 995.8, 
    995.9, 995.9, 996, 996.2, 995.9, 996.1, 996.1, 996.1, 996.1, 996.1, 
    996.2, 996.1, 996.1, 996.2, 996.3, 996.4, 996, 995.9, 995.7, 995.4, 
    995.4, 995.6, 995.8, 996.1, 996.3, 996.4, 996.4, 996.5, 996.8, 997.1, 
    997.3, 997.3, 997.5, 997.9, 998.3, 998.9, 998.9, 999.3, 999.5, 999.8, 
    1000.4, 1000.7, 1000.9, 1001.2, 1001.7, 1002.2, 1002.5, 1003, 1003.3, 
    1003.8, 1004.2, 1004.7, 1005.3, 1005.5, 1005.2, 1005.5, 1005.7, 1005.8, 
    1005.5, 1006, 1006.2, 1006, 1005.7, 1004.9, 1004.1, 1003.3, 1002.2, 
    1000.7, 999, 997.3, 995.3, 992.9, 990.6, 987.9, 985.7, 983.4, 981.3, 
    979.6, 977.9, 977.7, 977.6, 976.8, 977.3, 976.9, 976.7, 976.1, 975.3, 
    974.2, 973.3, 972.6, 971.6, 970.1, 969, 968.8, 969.7, 969.9, 969.7, 969, 
    969.2, 968.7, 970, 970.2, 970.5, 971.4, 972.5, 974.3, 976.1, 978.4, 
    980.7, 982.9, 984.2, 985.3, 985.6, 985.9, 986.3, 986.1, 985.7, 985, 
    984.4, 983.8, 983.6, 983.6, 983.3, 983.3, 983.1, 983.2, 983.6, 984.1, 
    983.9, 983.6, 983.8, 983.4, 982.9, 982.5, 982, 981.3, 980.4, 979.9, 
    979.4, 978.7, 978.2, 978.1, 978.1, 978.5, 978.7, 979.1, 979.6, 979.8, 
    980.5, 981.4, 981.5, 981.6, 982.1, 982.5, 983, 983.5, 984.2, 984.3, 
    984.5, 984.8, 985.1, 985.1, 984.9, 984.8, 985.4, 986, 986.5, 987.5, 
    988.5, 989.2, 989.7, 990.4, 991, 991.4, 991.9, 992.7, 993.4, 994.1, 
    995.2, 996.6, 997.9, 998.7, 999.2, 999.5, 999.6, 999.8, 999.2, 1000.1, 
    1001.2, 1002, 1002.7, 1003.9, 1004.2, 1004.8, 1005.8, 1006.8, 1007.8, 
    1009, 1009.5, 1010.7, 1011.3, 1011.9, 1012.1, 1012.6, 1013.2, 1013.7, 
    1014, 1014, 1014.1, 1014.3, 1014.3, 1014.1, 1013.9, 1014.1, 1014.3, 
    1014.4, 1014, 1014.1, 1013.8, 1013.6, 1013.4, 1013.1, 1013.1, 1012.8, 
    1012.5, 1012.4, 1012.4, 1012.2, 1011.9, 1011.6, 1011.4, 1011, 1010.7, 
    1010.6, 1010.2, 1009.9, 1009.6, 1009.5, 1009.3, 1009.2, 1008.8, 1008.4, 
    1008.2, 1007.8, 1007.2, 1006.7, 1006.4, 1005.7, 1005, 1004.3, 1003.8, 
    1003.3, 1003, 1002.5, 1001.8, 1000.6, 999.8, 999, 998, 997.1, 996, 994.8, 
    993.9, 992.6, 991.1, 989.8, 989, 987.4, 986.1, 984.8, 983.8, 983.2, 
    983.2, 983.5, 983.7, 984, 984.1, 984.2, 984.1, 984, 983.7, 983.6, 983.5, 
    983.2, 982.9, 982.6, 982.8, 983.4, 983.5, 983.4, 983.6, 984.2, 984.7, 
    984.9, 985.5, 986.4, 987.2, 988.4, 989.4, 990.8, 992.5, 994.1, 995.6, 
    997.2, 998.6, 1000.2, 1001.5, 1003.3, 1004.8, 1006, 1007.5, 1008.7, 
    1009.5, 1010.7, 1011.5, 1012, 1012.5, 1012.5, 1012.7, 1012.8, 1012.8, 
    1013.1, 1013.1, 1013.1, 1013.3, 1013, 1012.6, 1012.4, 1011.6, 1011.4, 
    1010.7, 1010.3, 1009.7, 1009.5, 1009, 1008.5, 1007.7, 1006.7, 1005.9, 
    1004.9, 1004, 1003.6, 1003, 1002.4, 1002.3, 1002.4, 1003.3, 1004.1, 
    1004.6, 1005.3, 1006.1, 1006.7, 1007.3, 1008, 1008.1, 1008.4, 1008.7, 
    1008.9, 1009, 1009.1, 1008.9, 1009, 1009, 1009.1, 1009.1, 1009.1, 1008.8, 
    1008.7, 1008.7, 1009, 1009.2, 1009.4, 1009.3, 1009.1, 1008.5, 1008.1, 
    1007.5, 1006.5, 1006.4, 1005.7, 1004.7, 1004.3, 1004, 1003.6, 1003.2, 
    1002.8, 1002.3, 1001.8, 1000.9, 1000.5, 1000.6, 1000.8, 1000.7, 1000.6, 
    1000.8, 1001.1, 1001, 1001, 1000.9, 1001, 1001.3, 1001.5, 1001.7, 1002.1, 
    1002.8, 1003.2, 1003.6, 1004.2, 1004.5, 1004.9, 1005.3, 1005.7, 1006.1, 
    1006.9, 1007.5, 1007.8, 1008.9, 1009.4, 1009.2, 1010, 1010.5, 1010.9, 
    1010.9, 1011.1, 1011.6, 1012.1, 1013.3, 1013.9, 1014.1, 1014.6, 1015.5, 
    1016.4, 1017.3, 1017.8, 1018.5, 1018.9, 1020, 1020.3, 1020.7, 1020.8, 
    1021.4, 1021.7, 1022.3, 1022.6, 1023, 1023, 1022.7, 1022.8, 1022.9, 
    1022.9, 1022.6, 1022.5, 1022.1, 1022, 1021.9, 1021.5, 1021.2, 1020.7, 
    1020.2, 1019.5, 1018.8, 1018.1, 1017.3, 1016.7, 1016, 1015.2, 1014.4, 
    1013.7, 1012.9, 1012.3, 1011.8, 1011, 1010.7, 1010.2, 1009.6, 1009.1, 
    1008.4, 1008.2, 1008, 1008.1, 1008, 1007.7, 1007.3, 1007.2, 1007.1, 
    1006.8, 1006.4, 1006.1, 1006, 1005.8, 1005.7, 1005.6, 1005.3, 1004.9, 
    1004.6, 1004.5, 1004.4, 1004.2, 1003.8, 1003.3, 1003, 1002.8, 1002.6, 
    1002.4, 1002.1, 1001.7, 1001.7, 1001.5, 1001, 1000.7, 1000.3, 1000, 
    999.8, 999.8, 999.9, 1000, 1000.2, 1000.5, 1000.9, 1001.4, 1001.9, 
    1002.3, 1003, 1003.4, 1004.5, 1005.2, 1006.1, 1006.9, 1007.3, 1007.6, 
    1007.6, 1008.1, 1008.2, 1007.8, 1007.7, 1007.3, 1006.8, 1006.5, 1006.4, 
    1006.1, 1006.2, 1006.2, 1006.4, 1006.4, 1006.3, 1006, 1005.7, 1005.9, 
    1005.7, 1005.6, 1005.9, 1006.4, 1006.7, 1006.7, 1006.4, 1006.2, 1006.3, 
    1006.6, 1006.8, 1006.9, 1007.3, 1007.3, 1007.7, 1007.8, 1008.3, 1008.6, 
    1008.7, 1009.2, 1009.3, 1010.2, 1010.8, 1011.2, 1011.5, 1012, 1012.6, 
    1013.3, 1014.1, 1014.3, 1014.8, 1015.3, 1015.8, 1016, 1016.4, 1016.5, 
    1016.6, 1016.3, 1016.2, 1016, 1015.7, 1015.4, 1014.8, 1014.4, 1014.3, 
    1014.3, 1014.2, 1014, 1013.9, 1014.5, 1015.4, 1016, 1016.6, 1017.3, 
    1017.7, 1017.7, 1018.3, 1018.5, 1019, 1019.6, 1020.5, 1021.4, 1022, 
    1022.2, 1022.9, 1024.4, 1025, 1025.4, 1025.5, 1026, 1026.1, 1026.9, 
    1027.1, 1028.1, 1028.6, 1029.3, 1029.6, 1030, 1030.3, 1030.1, 1029.6, 
    1029.5, 1029.8, 1030.1, 1030.3, 1030.3, 1030.7, 1030.8, 1031.3, 1031.6, 
    1031.5, 1031.9, 1032.4, 1032.3, 1032.1, 1032, 1031.9, 1032.3, 1032.1, 
    1032.3, 1032, 1032.5, 1033, 1032.9, 1032.9, 1032.9, 1033.3, 1033.2, 
    1033.4, 1033.6, 1033.4, 1033.2, 1032.8, 1032.4, 1032.2, 1031.9, 1031.4, 
    1030.9, 1030.6, 1029.9, 1029.2, 1028.6, 1028.2, 1027.5, 1026.9, 1026, 
    1024.7, 1023.6, 1022.3, 1021, 1019.8, 1018.5, 1017, 1015.8, 1014.6, 
    1014.1, 1013.7, 1013.1, 1013, 1013.5, 1013.6, 1014.1, 1014.3, 1014.3, 
    1014.4, 1014, 1013.8, 1013.7, 1013.2, 1012.3, 1011.5, 1010.1, 1008.7, 
    1006.9, 1005.6, 1004.1, 1002.5, 1002.1, 1000.5, 999.2, 997.6, 995.7, 
    994.7, 992.5, 990, 987.8, 985.6, 982.9, 980.6, 979, 978.4, 978.2, 978.4, 
    979, 979.8, 981.2, 983.4, 985.8, 988, 989.6, 991.1, 992.9, 994.2, 994.7, 
    994.8, 995.7, 996.1, 997, 996.9, 996.3, 996.1, 996.3, 996.2, 996.4, 997, 
    998, 999.3, 1000.5, 1001.8, 1003.2, 1005, 1006.6, 1008.1, 1009.2, 1010.9, 
    1012.9, 1014.3, 1016.1, 1017.4, 1018.7, 1020.1, 1021.4, 1022.6, 1023.6, 
    1024.4, 1025.1, 1025.4, 1026.1, 1027, 1027.2, 1026.9, 1026.9, 1027.6, 
    1026.8, 1025.8, 1025, 1024, 1023, 1022.3, 1021.1, 1019.7, 1018.8, 1017.5, 
    1016.6, 1015.5, 1014.6, 1013.8, 1012.5, 1011.4, 1010.3, 1009.4, 1008.7, 
    1007.9, 1007.2, 1006.8, 1006.3, 1006.2, 1006.3, 1006.7, 1007.2, 1007.6, 
    1008.1, 1008.8, 1009.1, 1009.3, 1010.3, 1010.7, 1011.8, 1012.3, 1012.4, 
    1012.3, 1012.6, 1013.1, 1013.2, 1013, 1012.8, 1012.9, 1013.3, 1013.2, 
    1013, 1013.1, 1012.9, 1012.6, 1012.5, 1012.1, 1012, 1012, 1011.9, 1012, 
    1012, 1011.7, 1011.6, 1011.3, 1011.1, 1010.9, 1010.7, 1010.4, 1010.2, 
    1010, 1009.9, 1009.9, 1010, 1010.1, 1010, 1009.9, 1010, 1009.7, 1009.6, 
    1009.5, 1009.3, 1009.4, 1009.4, 1009.4, 1009.5, 1009.4, 1009.3, 1008.9, 
    1008.6, 1008.3, 1008.2, 1008, 1007.5, 1007.1, 1007.2, 1007.1, 1007.1, 
    1006.7, 1006.4, 1005.9, 1005.5, 1005.2, 1004.6, 1004, 1003.6, 1003, 
    1002.3, 1001.8, 1001.2, 1000.3, 999.6, 998.9, 998.1, 997.2, 995.8, 994.6, 
    993.4, 992, 990.7, 989.8, 988.9, 987.4, 985.9, 984, 982.7, 982.3, 982.2, 
    982.5, 982.6, 982.5, 982.6, 982.7, 982.7, 983.1, 983.2, 983, 982.9, 
    982.8, 983.1, 982.5, 982.1, 981.9, 981.4, 980.7, 980.3, 979.3, 978.4, 
    978.4, 978.2, 978.3, 978.6, 978.9, 979.2, 979.8, 979.9, 979.8, 979.7, 
    979.9, 980.1, 980.9, 981.1, 981.8, 982.9, 984, 985.1, 986.8, 988.1, 
    989.8, 991.6, 993, 995.4, 995.5, 996.1, 997.5, 998.3, 999.5, 999.3, 
    999.7, 999.9, 1000.8, 1001.5, 1001.3, 1001.2, 1000.6, 1000.7, 1000.5, 
    999.9, 999.9, 999.5, 999.5, 999.5, 999.5, 999, 998.9, 999.5, 999.6, 999, 
    999.1, 999.3, 999.2, 998.6, 998.7, 998.5, 998.6, 998.4, 998.6, 998.6, 
    998.2, 998.4, 998.6, 998.3, 998.6, 998.3, 998.3, 998.3, 998.2, 998, 
    998.3, 997.9, 997.9, 997.3, 997.2, 996.9, 996.6, 996.3, 996.3, 996.1, 
    996.4, 996.9, 997, 997.4, 997.8, 998.2, 998.8, 999.1, 999.6, 999.8, 
    1000.6, 1000.5, 1001.2, 1001.6, 1002.4, 1002.6, 1003.2, 1003.3, 1003.3, 
    1003.9, 1004.1, 1004.4, 1004.7, 1005, 1005.1, 1005.6, 1005.9, 1006.2, 
    1006.6, 1007.1, 1007.4, 1007.6, 1007.7, 1008.2, 1008.5, 1008.8, 1009.5, 
    1010, 1010.6, 1010.9, 1011.2, 1011.6, 1012, 1012.1, 1012.6, 1013.1, 
    1013.5, 1013.9, 1014.2, 1014.6, 1015, 1015.4, 1015.9, 1016.1, 1016.4, 
    1016.4, 1016.9, 1017.1, 1017.5, 1017.8, 1018.3, 1018.8, 1019.1, 1019.2, 
    1019.4, 1019.6, 1020, 1020.4, 1020.8, 1020.9, 1021.4, 1022, 1022.2, 
    1022.4, 1022.5, 1022.5, 1022.2, 1021.8, 1021.9, 1022, 1022, 1021.7, 
    1021.2, 1021, 1020.9, 1020.6, 1019.8, 1019.5, 1019.1, 1018.7, 1018, 
    1017.6, 1017.1, 1016.6, 1016.4, 1015.9, 1015.2, 1014.5, 1013.9, 1013.4, 
    1012.6, 1012.4, 1012, 1011.8, 1011.4, 1010.9, 1010.4, 1010.4, 1010.4, 
    1010.3, 1010.1, 1009.7, 1009.5, 1009.1, 1008.9, 1009, 1009, 1008.9, 
    1008.7, 1008.5, 1008.8, 1008.7, 1008.8, 1008.7, 1008.5, 1008.3, 1008.1, 
    1007.9, 1008, 1008.3, 1007.7, 1007.5, 1007.4, 1007.4, 1007.5, 1007.7, 
    1007.7, 1007.8, 1007.5, 1007.3, 1007.2, 1007.1, 1007.2, 1007.1, 1007, 
    1007.2, 1007.3, 1007.3, 1007, 1007, 1006.9, 1006.8, 1006.9, 1007, 1007.1, 
    1007, 1007.2, 1007.4, 1007.7, 1008.1, 1008.2, 1008.2, 1008.7, 1009.2, 
    1009.7, 1010.1, 1010.6, 1011.1, 1011.7, 1012.1, 1012.6, 1012.9, 1013.2, 
    1013.7, 1014.1, 1014.2, 1014.5, 1014.6, 1014.6, 1014.9, 1015.2, 1015.4, 
    1015.8, 1016.1, 1015.9, 1016, 1016.2, 1016.3, 1016.2, 1016.2, 1016.1, 
    1015.9, 1015.6, 1015.2, 1015, 1014.9, 1014.3, 1013.6, 1012.8, 1012.4, 
    1012.2, 1011.6, 1011.2, 1010.6, 1010.6, 1010.4, 1010.1, 1010, 1009.8, 
    1009.6, 1009.3, 1009.2, 1008.9, 1008.7, 1008.5, 1008.1, 1007.8, 1007.4, 
    1007.2, 1006.6, 1006.1, 1006, 1005.4, 1005.4, 1005.3, 1005.5, 1005.5, 
    1005.6, 1006, 1006.3, 1007, 1007.6, 1008.2, 1008.8, 1009.8, 1010.9, 
    1011.7, 1012.5, 1013.6, 1014.2, 1014.6, 1015, 1015.5, 1015.9, 1016.2, 
    1016.4, 1016.6, 1016.2, 1016.4, 1015.9, 1015.2, 1014.9, 1014.9, 1014.7, 
    1014.6, 1014.7, 1014.5, 1014.2, 1013.6, 1013.9, 1013.4, 1013, 1012.6, 
    1012.4, 1012.4, 1012.2, 1012.3, 1012.5, 1012.6, 1012.4, 1012.3, 1012.3, 
    1011.9, 1011.5, 1011.2, 1010.7, 1010.2, 1009.9, 1009.6, 1009.5, 1009, 
    1008.5, 1008, 1007.6, 1007.4, 1007.1, 1007, 1007.1, 1007.2, 1007.2, 1007, 
    1006.9, 1006.8, 1006.9, 1006.8, 1006.6, 1006.5, 1006.4, 1006.5, 1006.8, 
    1006.9, 1007.5, 1008.2, 1008.7, 1009.3, 1009.7, 1010, 1010.2, 1010.6, 
    1010.5, 1010.8, 1011, 1011.3, 1011.7, 1011.8, 1011.9, 1012.3, 1012.3, 
    1012.1, 1012.1, 1012.1, 1012.2, 1012.4, 1012.6, 1012.6, 1012.6, 1012.4, 
    1012.4, 1012.4, 1012.3, 1012.1, 1011.8, 1011.4, 1010.8, 1010.3, 1009.9, 
    1009.2, 1008.4, 1007.6, 1006.4, 1005.3, 1003.5, 1001.7, 999.7, 997.4, 
    996.9, 995.8, 995.6, 995.2, 995.2, 994.9, 994.8, 996.1, 997.4, 998.2, 
    999.1, 999.6, 1000.2, 1000.9, 1001.3, 1001.9, 1002.1, 1002.8, 1003, 
    1003.1, 1003.3, 1003, 1002.6, 1002.1, 1001.7, 1001.1, 1000.4, 1000, 
    999.6, 999.3, 999.2, 998.5, 998.6, 998.3, 998.2, 998.1, 997.7, 997.9, 
    998.1, 998.5, 998.9, 999.3, 999.9, 1000.4, 1001.9, 1002.1, 1002.8, 1004, 
    1005.4, 1005.9, 1006.7, 1007.2, 1008.3, 1008.9, 1009.2, 1009.5, 1009.6, 
    1009.6, 1010, 1010.2, 1010.3, 1010, 1009.8, 1009.3, 1008.8, 1007.8, 
    1006.9, 1005.9, 1005, 1004, 1002.6, 1001.3, 1000.2, 999.1, 998.4, 998, 
    997.8, 997.4, 997.1, 996.6, 996, 995.5, 995.1, 994.9, 994.7, 994.5, 
    994.3, 994.1, 993.8, 993.2, 992.6, 991.8, 990.9, 989.6, 988.3, 987, 986, 
    984.9, 984.3, 983.3, 982.2, 981.7, 980.7, 980.1, 979.2, 978.6, 977.9, 
    977, 976.2, 975.5, 975, 974.8, 974.5, 974.5, 974.6, 974.5, 974.4, 974.7, 
    975, 975.5, 975.9, 976.1, 976.4, 977, 978, 978, 978.2, 978.6, 979, 979.4, 
    979.9, 980.4, 980.9, 981.2, 981.6, 981.8, 982.4, 982.7, 983.1, 983.1, 
    983.5, 983.7, 984.1, 984.5, 984.6, 984.5, 984.9, 985.2, 985.3, 984.5, 
    985.1, 985.1, 984.7, 984.7, 984.7, 984.8, 984.9, 984.3, 984.4, 984.3, 
    984.5, 984.8, 984.3, 983.9, 983.6, 983.7, 983.6, 983.3, 983.1, 982.8, 
    982.8, 982.9, 983.3, 983.3, 983.6, 983.7, 983.4, 983.7, 983.4, 983.5, 
    983.5, 983.8, 983.9, 984, 983.9, 984, 984.1, 984.1, 984, 984, 984, 984, 
    983.7, 983.5, 983.6, 983.8, 983.6, 983.5, 983.5, 983.4, 983.3, 983.4, 
    983.2, 983.2, 983.2, 983.1, 983.4, 983.3, 983.6, 983.4, 983.5, 983.4, 
    983.6, 983.9, 984, 984.1, 984.4, 984.8, 984.9, 985.1, 985.2, 985.3, 
    985.5, 985.6, 985.6, 985.4, 985.3, 985.1, 985.1, 985.2, 985.2, 985.3, 
    985.5, 985.9, 986.1, 986.5, 987, 987.3, 987.4, 987.8, 988.2, 988.8, 
    989.4, 989.8, 990.3, 990.9, 991.4, 992.1, 992.6, 992.9, 993.4, 993.6, 
    994.4, 995.2, 995.5, 995.8, 996.5, 996.9, 997.5, 997.8, 998.4, 998.7, 
    999.1, 999.4, 999.5, 999.6, 999.9, 1000, 1000.4, 1000.7, 1000.9, 1001.1, 
    1001, 1001, 1001, 1001.3, 1001.5, 1001.4, 1001.4, 1001.3, 1001.3, 1001.3, 
    1001.2, 1001.1, 1001.1, 1000.8, 1000.4, 1000, 1000, 999.8, 999.5, 999.3, 
    999, 998.8, 998.8, 998.5, 998.2, 997.9, 997.4, 996.9, 996.5, 995.9, 
    995.4, 994.8, 994.7, 993.9, 993.3, 993.1, 992.6, 991.8, 991.4, 991.2, 
    991.2, 991.2, 991.2, 991.5, 991.7, 992.1, 992.4, 992.7, 993, 993.1, 
    993.8, 994.5, 995.3, 996, 997.2, 997.4, 998.3, 998.9, 999.6, 999.6, 1000, 
    1000.2, 1000.2, 1000.2, 1000.2, 1000, 1000, 1000, 999.8, 1000, 1000, 
    999.9, 999.8, 999.4, 999.3, 999.3, 999.7, 999.9, 1000.2, 1000.3, 1000.6, 
    1000.9, 1001.3, 1001.6, 1001.7, 1001.8, 1001.5, 1001.4, 1001, 1000.6, 
    999.9, 999.2, 999.3, 998.2, 997.3, 996.3, 995.4, 993.9, 992.2, 990.7, 
    989.3, 987.6, 986.4, 985.5, 984.6, 983.9, 983.3, 983, 983, 983.3, 983.8, 
    984.4, 984.8, 985.6, 986.8, 987.5, 988.9, 990.8, 992.5, 993.4, 995.7, 
    997.2, 998.1, 998.8, 999.6, 1000, 1000.8, 1001.3, 1001.5, 1002.1, 1002.4, 
    1001.9, 1002.2, 1002.3, 1002.3, 1002.5, 1002.3, 1002.4, 1002.6, 1003, 
    1003.7, 1004.6, 1004.6, 1005.4, 1006.1, 1006.2, 1007.2, 1008.1, 1008.5, 
    1008.6, 1009.1, 1009.7, 1009.9, 1010.4, 1011, 1011.8, 1011.6, 1012, 1012, 
    1012.8, 1012.8, 1013.5, 1014.1, 1014.1, 1014.2, 1014.8, 1014.9, 1014.9, 
    1015.1, 1015, 1014.8, 1014.3, 1014.2, 1014.7, 1014.8, 1015.1, 1015.4, 
    1015.4, 1015.2, 1015.2, 1014.9, 1014.7, 1014.4, 1014.2, 1013.7, 1013.4, 
    1013, 1012.7, 1012.5, 1012.4, 1012.1, 1011.9, 1011.5, 1011.1, 1010.7, 
    1010.5, 1010.3, 1010.4, 1010.6, 1010.7, 1010.6, 1010.7, 1010.4, 1010.4, 
    1010.1, 1009.8, 1009.5, 1009.4, 1009.3, 1009.2, 1009.4, 1009.4, 1009.3, 
    1009.3, 1009.2, 1009.6, 1009.9, 1010.1, 1010.2, 1010.2, 1010.1, 1010, 
    1009.8, 1009.8, 1009.5, 1009.5, 1009.5, 1009.5, 1009.5, 1009.4, 1009.2, 
    1009, 1009, 1009.1, 1009.1, 1009.1, 1008.9, 1009, 1009, 1008.8, 1008.7, 
    1008.4, 1008.3, 1008.3, 1008.3, 1008.1, 1008.4, 1008.3, 1008.3, 1008.5, 
    1008.4, 1008.6, 1009, 1009.1, 1009.4, 1009.6, 1009.8, 1010.1, 1010.2, 
    1010.3, 1010.8, 1011.1, 1011.3, 1011.7, 1011.5, 1011.9, 1012.2, 1012.4, 
    1012.6, 1012.8, 1013.1, 1013.2, 1013.5, 1013.9, 1014.3, 1014.5, 1014.9, 
    1015.1, 1015.3, 1015.1, 1015.2, 1015.3, 1015.2, 1015.2, 1015, 1015, 
    1014.7, 1014.5, 1014.4, 1014.2, 1013.3, 1012.3, 1012, 1011.6, 1011.2, 
    1010.6, 1009.7, 1009, 1008.5, 1008, 1007.6, 1006.9, 1006.2, 1005.3, 
    1004.6, 1004.2, 1003.6, 1003.2, 1002.9, 1002.5, 1002.1, 1002, 1001.6, 
    1001.3, 1001.7, 1001.5, 1001.5, 1001.4, 1002.1, 1002.4, 1003.3, 1004.2, 
    1004.6, 1005.2, 1005.5, 1005.9, 1006.3, 1006.5, 1006.5, 1006.7, 1006.9, 
    1007, 1006.9, 1007.2, 1007.4, 1007.2, 1007.1, 1007.2, 1007.1, 1007.2, 
    1007.3, 1007.6, 1007.8, 1007.8, 1008, 1008.2, 1008, 1007.9, 1007.7, 
    1007.7, 1007.6, 1007.6, 1007.9, 1007.8, 1007.7, 1007.9, 1008.1, 1008.7, 
    1009.2, 1009.4, 1009.7, 1010.1, 1010.4, 1010.6, 1010.4, 1010.2, 1010, 
    1010.1, 1010.2, 1010.2, 1010.2, 1010.3, 1010.1, 1010.1, 1010.1, 1010, 
    1010.1, 1010.2, 1010.5, 1010.5, 1011.2, 1011.3, 1011.3, 1011.4, 1011.7, 
    1011.9, 1012.1, 1012.5, 1012.7, 1013, 1013.5, 1013.2, 1013.3, 1013.4, 
    1013.4, 1013.7, 1013.9, 1014, 1014.2, 1014.4, 1014.6, 1015, 1015.2, 
    1015.4, 1015.6, 1015.7, 1015.6, 1015.7, 1015.9, 1015.8, 1015.9, 1016.1, 
    1016.2, 1016.4, 1016.3, 1016.5, 1016.6, 1016.5, 1016.4, 1016.4, 1016, 
    1015.7, 1015.6, 1015.5, 1015.2, 1015.1, 1015.1, 1015.1, 1015, 1015.1, 
    1015.1, 1014.9, 1014.8, 1014.3, 1014, 1013.8, 1013.4, 1013.3, 1013, 
    1012.8, 1012.9, 1012.7, 1012.3, 1011.8, 1011.4, 1011.1, 1010.9, 1010.9, 
    1011.1, 1011, 1011.1, 1011.2, 1011.1, 1010.9, 1010.9, 1010.5, 1010.4, 
    1010.2, 1009.8, 1009.5, 1009.4, 1008.9, 1008.8, 1008.7, 1008.4, 1008.3, 
    1008, 1007.9, 1008, 1007.9, 1008.1, 1008.3, 1008.5, 1009, 1009.3, 1009.3, 
    1009.3, 1009.4, 1009.9, 1010.1, 1010.3, 1010.5, 1010.8, 1011, 1011.4, 
    1011.6, 1011.9, 1012.2, 1012.6, 1012.9, 1013.1, 1013.3, 1013.8, 1014.1, 
    1014.5, 1014.5, 1015, 1015.3, 1015.7, 1016, 1016.4, 1016.7, 1017.1, 
    1017.3, 1017.6, 1017.9, 1018.2, 1018.1, 1018.4, 1018.6, 1018.9, 1019.4, 
    1019.7, 1019.7, 1019.9, 1020.2, 1020.4, 1020.7, 1020.7, 1020.8, 1021, 
    1021.4, 1022, 1022.2, 1022.4, 1022.6, 1022.8, 1022.9, 1022.9, 1023.1, 
    1023.1, 1023.1, 1023.2, 1023.1, 1023.2, 1023.5, 1023.6, 1023.6, 1023.6, 
    1023.6, 1023.7, 1023.5, 1023.3, 1023.1, 1023, 1023.1, 1023, 1023, 1023.1, 
    1023, 1022.9, 1022.8, 1022.6, 1022.5, 1022.1, 1021.9, 1021.5, 1021.2, 
    1021.2, 1021, 1020.7, 1020.2, 1019.8, 1019.3, 1018.8, 1018.4, 1018.1, 
    1018.2, 1018.9, 1019.6, 1020.4, 1020.8, 1021.3, 1021.7, 1022, 1022.4, 
    1023.2, 1023.3, 1023.7, 1023.6, 1023.7, 1023.9, 1024, 1024.1, 1024.2, 
    1024.3, 1024.5, 1024.4, 1024.5, 1024.8, 1024.9, 1025.2, 1025, 1024.9, 
    1024.8, 1024.9, 1024.8, 1024.9, 1025.1, 1024.7, 1024.5, 1024.5, 1024.3, 
    1024.2, 1023.9, 1024.2, 1024.2, 1024.3, 1024.3, 1024.5, 1024.4, 1024.1, 
    1024.1, 1024.1, 1023.9, 1023.9, 1023.8, 1023.6, 1023.6, 1023.4, 1023.2, 
    1023.1, 1022.9, 1023, 1023, 1022.8, 1022.9, 1022.7, 1022.7, 1022.7, 
    1022.6, 1022.6, 1022.5, 1022.5, 1022.3, 1022.2, 1022.1, 1022.1, 1022, 
    1021.9, 1021.5, 1021.1, 1021.1, 1020.8, 1020.7, 1020.6, 1020.2, 1020.1, 
    1019.9, 1019.7, 1019.7, 1019.4, 1019.2, 1019.1, 1019, 1019.1, 1019.1, 
    1019, 1018.8, 1018.8, 1018.9, 1019.2, 1019.2, 1018.9, 1018.9, 1019.1, 
    1019.2, 1019.3, 1019.3, 1019.4, 1019.7, 1019.6, 1019.4, 1019.4, 1019.4, 
    1019.2, 1019.2, 1019.1, 1019.2, 1019.1, 1018.9, 1019.1, 1019, 1019, 
    1018.9, 1018.7, 1018.4, 1018, 1017.7, 1017.5, 1017.5, 1017.5, 1017.4, 
    1017.2, 1017.1, 1017.1, 1016.9, 1016.7, 1016.4, 1016.1, 1015.9, 1015.7, 
    1015.6, 1015.4, 1015.2, 1015, 1015, 1014.8, 1014.4, 1014.1, 1013.9, 
    1013.5, 1013.4, 1013.3, 1013.2, 1013.4, 1013.6, 1013.6, 1013.5, 1013.1, 
    1013.1, 1012.9, 1012.4, 1012.3, 1012.5, 1012.6, 1013, 1013.4, 1013.7, 
    1013.7, 1013.7, 1013.7, 1013.3, 1013.3, 1013.1, 1012.6, 1012.5, 1012.6, 
    1012.2, 1012.6, 1012.6, 1012.4, 1012.3, 1012.2, 1012.3, 1012.4, 1012.3, 
    1012.7, 1013.5, 1014, 1014.4, 1014.1, 1015.1, 1015.3, 1015.4, 1015.8, 
    1015.9, 1016, 1016.5, 1016.6, 1016.7, 1016.9, 1017.1, 1017.4, 1017.8, 
    1017.9, 1017.8, 1018, 1018, 1017.9, 1017.7, 1017.7, 1017.8, 1018, 1018.1, 
    1018.2, 1018.3, 1018.4, 1018.3, 1018.1, 1017.9, 1018, 1017.8, 1017.6, 
    1017.2, 1017.3, 1017.6, 1017.8, 1018.1, 1017.9, 1017.8, 1017.7, 1017.5, 
    1017.4, 1017.3, 1017.8, 1017.7, 1017.9, 1018.1, 1018.3, 1018.5, 1018.5, 
    1018.6, 1018.3, 1018.4, 1018.2, 1018, 1017.9, 1018, 1017.9, 1017.9, 
    1017.9, 1017.9, 1018.1, 1017.8, 1017.7, 1017.6, 1017.4, 1017.3, 1017.3, 
    1017.3, 1017.2, 1017.3, 1017.4, 1017.2, 1017.1, 1016.9, 1016.6, 1016.3, 
    1016.2, 1016, 1015.7, 1015.6, 1015.5, 1015.4, 1015.3, 1015.1, 1015.1, 
    1015.1, 1014.9, 1014.9, 1015, 1014.9, 1014.8, 1014.7, 1014.8, 1014.9, 
    1015, 1015.1, 1015.1, 1015.3, 1015.4, 1015.6, 1015.6, 1015.8, 1015.7, 
    1015.7, 1015.9, 1016, 1016.2, 1016.3, 1016.4, 1016.4, 1016.3, 1016.3, 
    1016.1, 1016, 1015.7, 1015.5, 1015.3, 1015.1, 1014.5, 1013.7, 1012.9, 
    1012.4, 1011.8, 1011.3, 1011, 1010.5, 1010.2, 1010, 1009.8, 1009.9, 
    1010.1, 1010.2, 1010, 1010.2, 1010.4, 1010.4, 1010.4, 1010.4, 1010.1, 
    1010, 1009.8, 1009.8, 1009.6, 1009.4, 1009.1, 1008.6, 1008.2, 1007.7, 
    1007, 1006.6, 1005.9, 1005.5, 1005.2, 1005, 1004.9, 1005.2, 1005.8, 
    1006.8, 1007.6, 1008.7, 1009.2, 1009.9, 1009.8, 1010.3, 1010.4, 1010.6, 
    1010.8, 1010.8, 1010.7, 1010.6, 1011, 1011, 1011.7, 1012.1, 1012.5, 1013, 
    1013.4, 1013.7, 1014.1, 1014.6, 1014.9, 1015.8, 1016.3, 1017.2, 1018.2, 
    1019.3, 1020.6, 1021.9, 1023, 1023.8, 1025.1, 1026, 1026.7, 1027.1, 
    1027.7, 1028.4, 1028.5, 1028.7, 1028.8, 1028.9, 1029.2, 1029.3, 1029.7, 
    1030.1, 1030.1, 1030.3, 1030.4, 1030.3, 1030, 1029.6, 1029.2, 1029.1, 
    1029, 1028.8, 1028.5, 1028.3, 1028.1, 1027.7, 1027, 1026.7, 1026.5, 
    1026.3, 1025.5, 1024.7, 1024.1, 1023.7, 1023.3, 1023.2, 1022.7, 1022.3, 
    1021.9, 1021.7, 1021.3, 1020.9, 1020.7, 1020.3, 1020.1, 1020, 1020, 
    1020.2, 1020.2, 1020.2, 1020.1, 1020.3, 1020.1, 1020.4, 1020.7, 1021, 
    1021.5, 1022.2, 1022.6, 1023.1, 1023.7, 1024.3, 1024.8, 1025.3, 1025.8, 
    1025.9, 1026.1, 1026.5, 1026.7, 1026.9, 1027, 1027.1, 1027.1, 1027, 
    1027.1, 1027.2, 1027.2, 1026.9, 1026.5, 1026.1, 1025.6, 1025.3, 1024.4, 
    1023.9, 1022.9, 1021.7, 1020.3, 1019, 1017.8, 1016.9, 1015.9, 1015.2, 
    1014.6, 1013.7, 1013.3, 1012.5, 1012.3, 1011.7, 1011.3, 1011.2, 1010.8, 
    1010.6, 1010, 1010.2, 1010.1, 1010.1, 1009.9, 1009.9, 1010.1, 1009.5, 
    1009.9, 1010.5, 1011, 1011.3, 1011.7, 1012.4, 1013.2, 1013.4, 1014.5, 
    1015.5, 1016.1, 1016.7, 1017.6, 1018.1, 1018.9, 1019.9, 1020.4, 1021.1, 
    1021.7, 1022.6, 1023.4, 1024.4, 1025.1, 1025.6, 1026.2, 1026.9, 1027.3, 
    1027.7, 1027.7, 1028, 1028.1, 1028.2, 1028.5, 1028.5, 1028.7, 1028.7, 
    1028.8, 1028.7, 1028.5, 1028.4, 1028, 1027.8, 1027.7, 1027.6, 1027.6, 
    1027.7, 1028.2, 1027.7, 1028.6, 1028.9, 1029.2, 1029.1, 1029.2, 1029.7, 
    1029.7, 1029.7, 1029.9, 1030.3, 1030.2, 1030, 1030.4, 1030.2, 1030.2, 
    1030.4, 1030.5, 1030.6, 1030.4, 1030.5, 1030.7, 1030.9, 1031.1, 1031.2, 
    1031.1, 1031.1, 1031.2, 1031.1, 1031, 1031.3, 1031.4, 1031.9, 1031.8, 
    1032, 1032, 1032.2, 1032.3, 1032.1, 1032.2, 1032.2, 1032.3, 1032.4, 
    1032.5, 1032.3, 1032.7, 1032.7, 1032.8, 1032.8, 1033.1, 1032.9, 1032.7, 
    1032.7, 1032.5, 1032.2, 1032.1, 1032, 1032, 1031.8, 1031.6, 1031.6, 
    1031.3, 1031, 1030.9, 1030.8, 1030.6, 1030.3, 1030.4, 1030.6, 1030.7, 
    1030.8, 1031, 1031.2, 1031.6, 1031.8, 1032.1, 1032.3, 1032.6, 1033, 
    1033.3, 1033.8, 1034, 1034.3, 1034.4, 1034.6, 1034.6, 1034.4, 1034.3, 
    1034.2, 1033.9, 1034.6, 1033.4, 1033.3, 1033.1, 1033.2, 1032.9, 1032.6, 
    1032.3, 1032.2, 1031.9, 1031.6, 1031.3, 1031, 1030.7, 1030.6, 1030.7, 
    1030.6, 1030.3, 1030, 1029.9, 1029.6, 1029.4, 1029.2, 1028.9, 1028.5, 
    1028.5, 1028.5, 1028.6, 1028.7, 1028.6, 1028.6, 1028.5, 1028.4, 1028.4, 
    1028.3, 1028.2, 1028.4, 1028.4, 1028.5, 1028.6, 1028.6, 1028.8, 1028.9, 
    1028.9, 1028.9, 1029.1, 1029, 1028.9, 1028.8, 1029, 1029, 1029, 1029.2, 
    1029.3, 1029.4, 1029.4, 1029.3, 1029.3, 1029.2, 1029.1, 1029, 1029, 
    1029.1, 1029.2, 1029.4, 1029.4, 1029.4, 1029.4, 1029.4, 1029.6, 1029.4, 
    1029.3, 1029.3, 1029.4, 1029.6, 1029.8, 1029.8, 1029.9, 1030.1, 1030.3, 
    1030.4, 1030.4, 1030.6, 1030.6, 1030.6, 1030.6, 1030.7, 1030.7, 1030.9, 
    1031, 1030.9, 1030.7, 1030.7, 1030.8, 1030.8, 1030.8, 1030.7, 1030.6, 
    1030.5, 1030.3, 1030.1, 1029.9, 1029.7, 1029.1, 1028.7, 1028.1, 1027.4, 
    1026.8, 1025.8, 1024.4, 1023.7, 1022.7, 1022, 1021.1, 1020.4, 1019.1, 
    1018.1, 1016.9, 1016.7, 1016.5, 1016.4, 1016.1, 1015.9, 1015.8, 1015.8, 
    1016.2, 1016.2, 1016.6, 1016.7, 1017, 1017.3, 1017.7, 1017.9, 1018.2, 
    1018.4, 1018.7, 1018.9, 1019.1, 1019.3, 1019.4, 1019.5, 1019.7, 1019.7, 
    1019.5, 1019.4, 1019.5, 1019.6, 1019.7, 1020.1, 1020.1, 1020.1, 1020.2, 
    1020.1, 1020, 1020.2, 1020.2, 1020.1, 1020.2, 1020.3, 1020.5, 1020.8, 
    1020.7, 1020.9, 1021, 1021.1, 1020.9, 1021.1, 1021, 1021.1, 1021.1, 
    1021.2, 1021.2, 1021.4, 1021.5, 1021.7, 1021.8, 1021.8, 1021.7, 1021.4, 
    1021.3, 1021.3, 1021.3, 1021.1, 1021, 1021, 1020.9, 1020.8, 1020.7, 
    1020.5, 1020.3, 1020.1, 1019.9, 1019.9, 1019.8, 1019.7, 1019.7, 1019.7, 
    1019.8, 1019.9, 1020, 1020, 1020, 1019.9, 1019.7, 1019.5, 1019.3, 1019.3, 
    1019.4, 1019.4, 1019.5, 1019.4, 1019.2, 1019.2, 1019.2, 1019.3, 1019.2, 
    1019.1, 1019.2, 1019.4, 1019.6, 1019.8, 1019.9, 1019.8, 1019.7, 1019.9, 
    1019.9, 1019.8, 1019.6, 1019.5, 1019.4, 1019.4, 1019.4, 1019.4, 1019.5, 
    1019.2, 1019.1, 1019, 1018.5, 1018.4, 1018.1, 1017.8, 1017.6, 1017.6, 
    1017.5, 1017.7, 1017.6, 1017.5, 1017.2, 1017.1, 1016.6, 1016.3, 1016.2, 
    1016, 1015.7, 1015.5, 1015.3, 1015, 1015.1, 1014.8, 1014.7, 1014.5, 
    1014.4, 1014, 1013.6, 1013.2, 1012.9, 1012.8, 1012.4, 1012, 1011.8, 
    1011.5, 1010.8, 1010.4, 1009.8, 1009.3, 1008.9, 1008.3, 1007.9, 1007.7, 
    1007.7, 1007.7, 1007.9, 1008, 1007.8, 1007.7, 1007.9, 1007.8, 1007.9, 
    1008.2, 1008.1, 1008.1, 1008.4, 1008.8, 1008.8, 1008.7, 1008.9, 1009.1, 
    1009.2, 1009.3, 1009.3, 1009.4, 1009.6, 1010.1, 1010, 1010.3, 1010.3, 
    1010.4, 1010.6, 1010.6, 1010.6, 1010.5, 1010.5, 1010.5, 1010.3, 1010.5, 
    1010.8, 1010.9, 1010.8, 1011.1, 1010.9, 1010.9, 1010.8, 1010.8, 1010.8, 
    1011.1, 1011.1, 1011, 1010.9, 1010.9, 1011.2, 1011.3, 1011.4, 1011.5, 
    1011.5, 1011.4, 1011.6, 1011.6, 1011.6, 1011.8, 1011.9, 1012.1, 1012.2, 
    1012.3, 1012.5, 1012.6, 1012.8, 1012.9, 1013.1, 1013.2, 1013.4, 1013.4, 
    1013.5, 1013.6, 1013.7, 1013.7, 1013.9, 1014, 1014.2, 1014.3, 1014.4, 
    1014.6, 1014.7, 1015.1, 1015.4, 1015.6, 1015.8, 1016, 1016.2, 1016.4, 
    1016.6, 1016.6, 1016.7, 1016.7, 1016.8, 1016.8, 1016.9, 1017, 1017.1, 
    1017.2, 1017.2, 1017.4, 1017.2, 1017.1, 1017, 1017, 1016.8, 1016.8, 
    1016.7, 1016.8, 1016.7, 1016.5, 1016.3, 1016.4, 1016.5, 1016.6, 1016.4, 
    1016.3, 1016.4, 1016.6, 1017, 1017, 1017.4, 1017.8, 1018.2, 1018.5, 
    1018.9, 1019.1, 1019.1, 1019.3, 1019.6, 1020, 1020.2, 1020.5, 1020.6, 
    1021.1, 1021.3, 1021.4, 1021.4, 1021.5, 1021.4, 1021.4, 1021.5, 1021.4, 
    1021.4, 1021.4, 1021.7, 1021.7, 1021.7, 1021.4, 1021.5, 1021.3, 1021.1, 
    1020.8, 1020.8, 1020.8, 1020.9, 1021, 1021.1, 1021.2, 1021.3, 1021.4, 
    1021.3, 1021.3, 1021.3, 1021.2, 1021.1, 1021.2, 1021.4, 1021.3, 1021, 
    1020.7, 1020.2, 1019.6, 1019.2, 1018.9, 1018.2, 1017.7, 1017.3, 1016.5, 
    1016.2, 1015.7, 1015, 1014.6, 1014.1, 1013.1, 1012.2, 1012.6, 1011.8, 
    1011.3, 1010.8, 1011.1, 1011, 1011.1, 1011.1, 1011.1, 1011.4, 1011.5, 
    1012.2, 1012.3, 1012.6, 1012.9, 1013.4, 1013.7, 1014, 1014.3, 1013.9, 
    1013.7, 1013.9, 1013.8, 1013.8, 1014.9, 1015.1, 1015.2, 1014.9, 1016, 
    1016.6, 1016.8, 1017.5, 1017.6, 1017.9, 1018.2, 1018.8, 1019, 1018.9, 
    1019.1, 1019.4, 1019.2, 1019.3, 1019.2, 1019.2, 1019.2, 1019.1, 1019.1, 
    1019.2, 1019.4, 1019.5, 1020.1, 1020.4, 1020.4, 1020.8, 1021.2, 1021.5, 
    1022.5, 1023.3, 1023.8, 1023.9, 1024.3, 1024.8, 1025, 1025.7, 1026.2, 
    1026.4, 1026.9, 1027.3, 1027.6, 1027.9, 1028.2, 1028.3, 1028.8, 1029.1, 
    1029.3, 1029.7, 1030, 1030.1, 1030.2, 1030.3, 1030.3, 1030.2, 1030.2, 
    1030.4, 1030.4, 1030.3, 1030.3, 1030.1, 1030.2, 1030.1, 1030, 1029.8, 
    1029.8, 1029.7, 1029.4, 1029.4, 1029.1, 1028.8, 1028.4, 1028.1, 1027.8, 
    1027.5, 1027.2, 1027, 1026.6, 1026.1, 1025.8, 1025.6, 1025.2, 1024.8, 
    1024.5, 1024.3, 1024.3, 1024.2, 1023.9, 1023.7, 1023.6, 1023.5, 1023.6, 
    1023.5, 1023.4, 1023.4, 1023.4, 1023.3, 1023.2, 1023.1, 1023.3, 1023.4, 
    1023.3, 1023.5, 1023.5, 1023.6, 1023.8, 1023.9, 1023.9, 1024.1, 1024, 
    1024.1, 1024.3, 1024.6, 1024.5, 1024.3, 1024.3, 1024.5, 1024.5, 1024.5, 
    1024.4, 1024.2, 1024.2, 1023.9, 1024, 1023.7, 1023.4, 1023.3, 1023.3, 
    1023, 1022.8, 1022.7, 1022.2, 1022, 1021.7, 1021.7, 1021.4, 1021, 1020.5, 
    1020.3, 1020, 1019.8, 1019.6, 1019.3, 1019.1, 1019, 1018.8, 1018.2, 
    1018.1, 1017.8, 1017.6, 1017.5, 1017.2, 1016.9, 1016.8, 1016.6, 1016.4, 
    1016.6, 1016.3, 1016.5, 1016.5, 1016.3, 1016.8, 1017.1, 1017.1, 1017.3, 
    1017.6, 1017.9, 1018, 1018.2, 1018.5, 1018.9, 1019.3, 1019.4, 1019.8, 
    1020.1, 1020.2, 1020.5, 1020.7, 1020.6, 1020.5, 1020.6, 1020.7, 1020.8, 
    1020.8, 1020.5, 1020.4, 1020.6, 1020.8, 1020.9, 1021.1, 1021.2, 1021.7, 
    1021.9, 1022.2, 1022.4, 1022.8, 1022.9, 1023.1, 1023.4, 1023.8, 1024.3, 
    1024.3, 1024.4, 1024.6, 1025.1, 1025.2, 1025.7, 1026, 1026.3, 1026.4, 
    1026.6, 1026.9, 1027.1, 1027.4, 1027.5, 1027.5, 1027.5, 1027.5, 1027.8, 
    1028.1, 1028.3, 1028.5, 1028.6, 1028.8, 1028.9, 1029.1, 1029.1, 1029.1, 
    1029.3, 1029.3, 1029.4, 1029.6, 1029.2, 1029.2, 1029.3, 1029.2, 1029.2, 
    1029.2, 1029, 1028.7, 1028.4, 1028.3, 1028.3, 1028, 1027.8, 1027.4, 
    1027.4, 1027.4, 1027.3, 1027.1, 1027.1, 1026.9, 1026.9, 1026.9, 1026.9, 
    1026.9, 1026.7, 1026.6, 1026.6, 1026.6, 1026.5, 1026.4, 1026.1, 1025.6, 
    1025.1, 1024.7, 1024.6, 1024.2, 1023.9, 1023.4, 1023, 1022.5, 1022.3, 
    1021.9, 1021.3, 1020.8, 1020.2, 1019.8, 1019.4, 1019.1, 1018.9, 1018.7, 
    1018.3, 1018, 1017.6, 1017.3, 1016.9, 1016.5, 1016.2, 1015.8, 1015.6, 
    1015.2, 1015, 1014.7, 1014.5, 1014.3, 1014, 1013.4, 1013, 1012.6, 1012.2, 
    1011.9, 1011.7, 1011.5, 1011.4, 1011.2, 1011, 1011, 1010.8, 1010.6, 
    1010.5, 1010.2, 1010, 1009.9, 1009.7, 1009.5, 1009.4, 1009.3, 1009.2, 
    1008.8, 1008.7, 1008.6, 1008.6, 1008.3, 1008, 1007.8, 1007.9, 1007.9, 
    1007.8, 1007.5, 1007.4, 1007.4, 1007.2, 1007, 1006.7, 1006.2, 1006, 
    1005.7, 1005.5, 1005.3, 1005, 1004.5, 1004.3, 1004, 1003.8, 1003.5, 
    1003.1, 1002.8, 1002.4, 1002.2, 1002.2, 1001.9, 1001.8, 1001.9, 1001.8, 
    1001.5, 1001.5, 1001.5, 1001.6, 1001.7, 1001.7, 1001.8, 1001.7, 1001.8, 
    1001.8, 1001.9, 1001.8, 1001.8, 1001.8, 1001.8, 1001.6, 1001.4, 1001.3, 
    1001.3, 1001.2, 1001.4, 1001.5, 1001.6, 1001.6, 1001.4, 1001.4, 1001.3, 
    1001.1, 1001.1, 1000.8, 1000.9, 1000.9, 1001, 1001, 1001.1, 1001.3, 
    1001.5, 1001.8, 1002.1, 1002.2, 1002.5, 1002.7, 1003.2, 1003.7, 1004, 
    1004.4, 1004.8, 1005.3, 1005.6, 1005.7, 1006, 1006.3, 1006.6, 1006.9, 
    1007.2, 1007.5, 1007.9, 1008.1, 1008.3, 1008.6, 1008.7, 1008.9, 1009, 
    1008.8, 1009, 1009, 1009.1, 1009, 1009, 1009.2, 1009.2, 1009.2, 1009.2, 
    1009.1, 1008.8, 1008.6, 1008.4, 1008.3, 1008.1, 1007.9, 1008, 1007.8, 
    1007.9, 1007.9, 1007.9, 1007.6, 1007.3, 1007.1, 1006.9, 1006.9, 1007.1, 
    1007.2, 1007.3, 1007.3, 1007.5, 1007.4, 1007.5, 1007.5, 1007.6, 1007.4, 
    1007.3, 1007.3, 1007.3, 1007.4, 1007.4, 1007.5, 1007.5, 1007.6, 1007.5, 
    1007.4, 1007.2, 1007.1, 1006.9, 1006.8, 1007, 1006.9, 1006.9, 1007.2, 
    1007.2, 1007, 1006.9, 1006.9, 1006.7, 1006.7, 1006.7, 1006.6, 1006.5, 
    1006.4, 1006.4, 1006.3, 1006.3, 1006.2, 1006.5, 1006.6, 1006.7, 1006.8, 
    1006.8, 1007, 1007.3, 1007.9, 1008.2, 1008.4, 1008.4, 1008.6, 1008.6, 
    1008.8, 1009, 1009.4, 1009.4, 1009.6, 1009.8, 1009.9, 1010, 1010.2, 
    1010.4, 1010.3, 1010.5, 1010.5, 1010.7, 1010.7, 1010.8, 1011, 1011.1, 
    1011.3, 1011.5, 1011.3, 1011.4, 1011.6, 1011.8, 1011.7, 1011.7, 1011.6, 
    1011.7, 1011.8, 1011.8, 1011.8, 1011.8, 1011.7, 1012, 1012, 1012, 1012, 
    1011.9, 1011.9, 1012, 1012.1, 1012.2, 1012, 1011.9, 1011.8, 1011.8, 
    1011.9, 1011.8, 1011.6, 1011.5, 1011.4, 1011.2, 1011.1, 1011.1, 1011.1, 
    1011.1, 1011.1, 1011, 1011.1, 1011.3, 1011.3, 1011.3, 1011.2, 1011.3, 
    1011.3, 1011.2, 1011.4, 1011.5, 1011.6, 1011.5, 1011.5, 1011.3, 1011.4, 
    1011.4, 1011.2, 1011, 1010.9, 1010.6, 1010.3, 1010.2, 1010.3, 1010.4, 
    1010.3, 1010.3, 1010.3, 1010, 1009.9, 1009.8, 1009.9, 1009.9, 1009.8, 
    1010, 1010, 1009.9, 1009.9, 1009.9, 1009.9, 1009.9, 1009.9, 1009.7, 
    1009.5, 1009.6, 1009.7, 1009.7, 1009.7, 1009.9, 1009.9, 1009.9, 1009.9, 
    1009.6, 1009.5, 1009.4, 1009.4, 1009.3, 1009.1, 1009.3, 1009.3, 1009.3, 
    1009.1, 1009, 1008.6, 1008.6, 1008.6, 1008.5, 1008.3, 1008.1, 1008.1, 
    1007.8, 1007.6, 1007.5, 1007.2, 1007, 1006.8, 1006.4, 1006.1, 1005.7, 
    1005.4, 1005.2, 1005, 1004.9, 1004.7, 1004.5, 1004.3, 1003.9, 1003.7, 
    1003.6, 1003.3, 1003.2, 1003, 1003, 1003, 1002.9, 1002.8, 1002.7, 1002.6, 
    1002.4, 1002.4, 1002.4, 1002.3, 1002.4, 1002.3, 1002.3, 1002.3, 1002.5, 
    1002.5, 1002.5, 1002.6, 1002.5, 1002.4, 1002.4, 1002.6, 1002.6, 1002.3, 
    1002.2, 1002.1, 1002.2, 1002, 1001.8, 1001.7, 1001.4, 1001.2, 1000.7, 
    1000.6, 1000.3, 1000, 999.9, 999.9, 999.7, 999.4, 999.1, 999.1, 998.9, 
    998.6, 998.3, 998.4, 998.3, 998.5, 998.6, 998.8, 998.9, 999.4, 999.6, 
    999.8, 1000.2, 1000.6, 1000.9, 1001.2, 1001.6, 1002.1, 1002.4, 1002.9, 
    1003.5, 1003.9, 1004.3, 1004.8, 1005.3, 1006, 1006.6, 1007.2, 1007.8, 
    1008.5, 1009.1, 1009.9, 1010.6, 1011.2, 1011.9, 1012.4, 1013, 1013.4, 
    1013.7, 1013.9, 1014.3, 1014.6, 1014.8, 1015.3, 1015.6, 1015.9, 1016.1, 
    1016.3, 1016.4, 1016.6, 1016.9, 1017.1, 1017, 1017.2, 1017.7, 1017.9, 
    1018.1, 1018.2, 1018.2, 1018.4, 1018.2, 1018.1, 1018, 1017.7, 1017.6, 
    1017.5, 1017.2, 1017.1, 1017.2, 1017, 1016.8, 1016.6, 1016.3, 1016.1, 
    1015.7, 1015.4, 1015.1, 1014.9, 1014.9, 1014.7, 1014.8, 1014.8, 1014.7, 
    1014.6, 1014.3, 1014.2, 1014, 1013.9, 1013.7, 1013.7, 1013.6, 1013.7, 
    1013.8, 1013.5, 1013.5, 1013.5, 1013.5, 1013.5, 1013.4, 1013.4, 1013.2, 
    1013.2, 1013.2, 1013.1, 1013.3, 1013.4, 1013.4, 1013.4, 1013.4, 1013.3, 
    1012.9, 1012.6, 1012.3, 1012, 1011.9, 1011.7, 1011.6, 1011.8, 1011.7, 
    1011.7, 1011.2, 1010.7, 1010.5, 1009.8, 1009.7, 1009.3, 1008.8, 1008.5, 
    1008.3, 1007.6, 1007, 1006.8, 1006.4, 1006.1, 1005.8, 1005.4, 1005, 
    1004.6, 1004.5, 1004.2, 1003.9, 1003.8, 1003.4, 1003.2, 1002.9, 1002.7, 
    1002.3, 1001.9, 1001.7, 1001.5, 1001.4, 1001.5, 1001.5, 1001.5, 1001.5, 
    1001.4, 1001.4, 1001.2, 1001.4, 1001.5, 1001.5, 1001.6, 1001.8, 1002.1, 
    1002.4, 1002.8, 1003, 1003.3, 1003.5, 1003.8, 1004.2, 1004.3, 1004.5, 
    1004.8, 1005, 1005.4, 1005.7, 1006.3, 1007, 1007.2, 1007.3, 1007.6, 
    1007.8, 1007.9, 1007.9, 1008.2, 1008.2, 1008.6, 1009, 1009.4, 1009.7, 
    1009.9, 1009.8, 1010, 1009.9, 1009.8, 1009.9, 1009.8, 1009.7, 1009.9, 
    1010, 1010.1, 1010.1, 1010.1, 1009.9, 1009.6, 1009.4, 1009.3, 1009.1, 
    1009, 1008.9, 1008.6, 1008.4, 1008.2, 1008, 1007.6, 1007.1, 1006.9, 
    1006.6, 1006.2, 1005.7, 1005.4, 1005, 1004.6, 1004.2, 1004.1, 1003.8, 
    1003.4, 1003, 1002.6, 1002.4, 1002.2, 1001.8, 1001.6, 1001.4, 1001.2, 
    1001.3, 1001.4, 1001.5, 1001.6, 1001.3, 1001.4, 1001.2, 1001.3, 1001.4, 
    1001.5, 1001.7, 1001.9, 1002.2, 1002.7, 1002.9, 1003.4, 1003.7, 1003.9, 
    1004.1, 1004.3, 1004.5, 1004.7, 1004.8, 1005.1, 1005.2, 1005.3, 1005.4, 
    1005.5, 1005.4, 1005.5, 1005.5, 1005.4, 1005.7, 1005.8, 1006.2, 1006.5, 
    1006.7, 1007.1, 1007.5, 1007.6, 1007.8, 1008, 1007.9, 1008.1, 1008.4, 
    1008.6, 1008.8, 1009.1, 1009.2, 1009.3, 1009.3, 1009.3, 1009.3, 1009.4, 
    1009.4, 1009.5, 1009.4, 1009.4, 1009.4, 1009.4, 1009.5, 1009.5, 1009.5, 
    1009.4, 1009.3, 1009.1, 1009, 1009, 1008.8, 1008.6, 1008.5, 1008.3, 
    1008.1, 1008, 1008, 1008.1, 1008, 1007.7, 1007.6, 1007.5, 1007.4, 1007.4, 
    1007.4, 1007.4, 1007.4, 1007.5, 1007.4, 1007.3, 1007.2, 1007.2, 1007, 
    1007, 1006.8, 1006.9, 1006.9, 1007.1, 1007, 1007, 1006.9, 1006.9, 1007, 
    1007, 1007.1, 1007.2, 1007.3, 1007.4, 1007.4, 1007.6, 1007.4, 1007.5, 
    1007.3, 1007.3, 1007.2, 1006.9, 1006.6, 1006.4, 1006.2, 1006, 1005.7, 
    1005.3, 1005.1, 1004.5, 1004.1, 1003.9, 1003.6, 1003.1, 1002.8, 1002.5, 
    1002.2, 1001.7, 1001.6, 1001.3, 1001, 1000.9, 1000.9, 1000.9, 1001, 1001, 
    1000.9, 1000.8, 1000.4, 1000.3, 1001.1, 1001.8, 1002.5, 1003.2, 1003.8, 
    1004.2, 1005, 1005.8, 1006.2, 1007.2, 1007.9, 1008.9, 1009.9, 1010.6, 
    1011.4, 1011.9, 1012, 1012.1, 1012.6, 1012.7, 1013.1, 1013.4, 1013.7, 
    1013.9, 1014, 1014.1, 1014.4, 1014.5, 1014.5, 1014.3, 1014.1, 1013.8, 
    1013.9, 1013.8, 1013.5, 1013, 1012.7, 1012.3, 1012.5, 1011.9, 1011.6, 
    1010.7, 1010.1, 1009.5, 1008.7, 1008.2, 1007.5, 1006.2, 1005.2, 1004.6, 
    1004, 1003.4, 1002.8, 1002.2, 1001.3, 1000.7, 1000.5, 1000.2, 1000.2, 
    1000.3, 1000.3, 1000.2, 1000.6, 1000.9, 1001.1, 1001.1, 1001.2, 1001.1, 
    1001, 1000.6, 1000.2, 1000.5, 1000.3, 1000.7, 1000.9, 1001.4, 1001.6, 
    1002.1, 1002.8, 1002.9, 1003.1, 1003.7, 1004.4, 1005.1, 1005.8, 1006, 
    1006.5, 1007.3, 1007.8, 1008.1, 1008.5, 1008.8, 1008.8, 1009.4, 1009.9, 
    1009.8, 1010.1, 1010.5, 1010.6, 1010.8, 1010.9, 1011, 1010.8, 1011, 
    1010.6, 1010.1, 1009.9, 1009.7, 1009.5, 1009.3, 1009.4, 1009.3, 1009.1, 
    1008.6, 1008.5, 1008.2, 1008, 1008.1, 1007.9, 1008, 1007.8, 1007.8, 
    1007.8, 1007.8, 1008, 1008.2, 1008.5, 1008.5, 1008.7, 1008.9, 1009.3, 
    1009.7, 1010, 1010.4, 1010.7, 1011.1, 1011.2, 1011.3, 1011.3, 1011.4, 
    1011.6, 1011.3, 1011.2, 1010.9, 1010.4, 1009.8, 1009.3, 1008.6, 1007.9, 
    1007.3, 1006.8, 1006.2, 1006.1, 1006.3, 1006.5, 1006.6, 1006.8, 1006.9, 
    1007.1, 1007.5, 1007.7, 1008.2, 1008.6, 1009.1, 1009.2, 1009.4, 1009.7, 
    1010.1, 1010.6, 1011.3, 1011.8, 1012.4, 1013, 1013.8, 1014.5, 1014.9, 
    1015.3, 1015.5, 1015.8, 1016.2, 1016.7, 1017.2, 1017.8, 1018.3, 1018.5, 
    1018.8, 1019.1, 1019.3, 1019.5, 1019.8, 1019.9, 1019.9, 1019.7, 1019.6, 
    1019.8, 1019.8, 1019.9, 1020.1, 1019.8, 1019.4, 1018.8, 1018.3, 1017.9, 
    1017.4, 1017, 1016.7, 1015.9, 1015.7, 1015.4, 1015.2, 1015.4, 1015.9, 
    1016.3, 1016.7, 1016.9, 1017.5, 1017.9, 1018.1, 1018.4, 1018.5, 1019.1, 
    1019.8, 1019.9, 1019.8, 1019.5, 1019.6, 1019.7, 1019.8, 1019.8, 1019.7, 
    1019.7, 1019.6, 1019.6, 1019.5, 1019.6, 1019.3, 1019.3, 1019.2, 1018.9, 
    1018.8, 1018.7, 1018.5, 1018.4, 1018.1, 1017.8, 1017.6, 1017.2, 1016.7, 
    1016, 1015.7, 1015.5, 1014.9, 1014.8, 1014.7, 1014.5, 1014.2, 1013.7, 
    1013.5, 1013.4, 1013.4, 1013.3, 1013.1, 1013, 1012.9, 1013.1, 1013.3, 
    1013.5, 1013.7, 1014, 1014.1, 1014, 1014, 1014, 1014.1, 1014.3, 1014.4, 
    1014.6, 1014.8, 1014.9, 1015.2, 1015.4, 1015.5, 1015.5, 1015.5, 1015.4, 
    1015.3, 1015.2, 1015.1, 1014.9, 1014.6, 1014.3, 1014.2, 1014.1, 1013.7, 
    1013.3, 1013.1, 1012.7, 1012.4, 1011.9, 1011.6, 1011.4, 1011.1, 1011, 
    1010.6, 1010.2, 1010, 1009.7, 1009.2, 1008.8, 1008.7, 1008.5, 1008.4, 
    1008.1, 1007.8, 1007.4, 1007.2, 1007.1, 1006.9, 1006.8, 1006.8, 1006.5, 
    1006.2, 1006.1, 1006.1, 1005.8, 1005.8, 1005.7, 1005.7, 1005.5, 1005.4, 
    1005.3, 1005.2, 1005.1, 1005, 1005.3, 1005.5, 1005.8, 1006.2, 1006.4, 
    1006.8, 1007.2, 1007.6, 1008.1, 1008.4, 1008.8, 1009.2, 1009.3, 1010.2, 
    1010.4, 1010.6, 1010.9, 1011.5, 1011.8, 1011.9, 1012.1, 1012.2, 1012.5, 
    1012.5, 1012.7, 1012.9, 1012.9, 1013.1, 1013.4, 1013.5, 1013.7, 1013.7, 
    1013.9, 1014.1, 1013.9, 1014, 1014.1, 1014, 1014.1, 1014.4, 1014.6, 
    1014.8, 1014.8, 1015, 1014.8, 1014.6, 1014.4, 1014.5, 1014.3, 1014.3, 
    1014.3, 1014.3, 1014.7, 1014.7, 1014.6, 1014.6, 1014.4, 1014.5, 1014.4, 
    1014.2, 1014.2, 1014.4, 1014.5, 1014.4, 1014.5, 1014.6, 1014.3, 1014.2, 
    1013.9, 1013.5, 1013.3, 1013.1, 1012.8, 1012.7, 1012.7, 1012.4, 1012.3, 
    1011.9, 1011.8, 1011.6, 1011.4, 1011.1, 1010.9, 1010.6, 1010.7, 1010.6, 
    1010.8, 1010.9, 1011, 1011, 1010.9, 1010.7, 1010.4, 1010.1, 1010.1, 
    1009.9, 1009.6, 1009.3, 1009.7, 1009.7, 1009.4, 1009.2, 1009.1, 1009.1, 
    1009.1, 1008.8, 1008.5, 1008.4, 1008.3, 1008.5, 1008.3, 1008.6, 1008.6, 
    1008.9, 1008.9, 1008.9, 1009, 1009, 1009.1, 1009.2, 1009.2, 1009.3, 
    1009.3, 1009.7, 1009.8, 1010.1, 1010.1, 1010, 1010, 1009.9, 1010, 1009.9, 
    1010.1, 1010.1, 1010.4, 1010.5, 1010.5, 1010.8, 1011.3, 1011.1, 1010.9, 
    1011, 1011.1, 1011, 1010.9, 1010.8, 1010.9, 1011, 1011, 1011, 1011.1, 
    1011.1, 1010.9, 1010.8, 1010.5, 1010.2, 1010.3, 1010.3, 1010.4, 1010.5, 
    1010.6, 1010.7, 1010.7, 1010.8, 1010.9, 1010.9, 1011, 1011, 1011, 1011.1, 
    1011.1, 1011, 1011.1, 1011.3, 1011.4, 1011.4, 1011.4, 1011.3, 1011.3, 
    1011.1, 1011.1, 1011.1, 1011.3, 1011.5, 1011.6, 1011.8, 1011.9, 1012, 
    1012, 1012.2, 1012.2, 1012.2, 1012.3, 1012.4, 1012.6, 1012.7, 1012.8, 
    1013.2, 1013.5, 1013.7, 1014, 1014.1, 1014.2, 1014.1, 1014.1, 1014.2, 
    1014.4, 1014.5, 1014.5, 1014.6, 1014.7, 1014.8, 1014.9, 1014.7, 1014.7, 
    1014.7, 1014.7, 1014.8, 1015.1, 1015.3, 1015.4, 1015.6, 1015.8, 1015.8, 
    1015.9, 1015.8, 1015.6, 1015.7, 1015.6, 1015.5, 1015.5, 1015.6, 1015.7, 
    1015.9, 1015.8, 1015.8, 1015.8, 1015.9, 1015.8, 1015.6, 1015.5, 1015.5, 
    1015.4, 1015.5, 1015.5, 1015.6, 1015.6, 1015.6, 1015.6, 1015.5, 1015.5, 
    1015.4, 1015.4, 1015.3, 1015.6, 1015.6, 1015.8, 1015.9, 1016.1, 1016.4, 
    1016.5, 1016.6, 1016.6, 1016.6, 1016.6, 1016.8, 1017, 1017.2, 1017.3, 
    1017.7, 1018, 1018.2, 1018.4, 1018.7, 1018.8, 1018.9, 1018.9, 1018.9, 
    1019.1, 1019.4, 1019.8, 1020, 1020.2, 1020.5, 1020.7, 1020.7, 1020.8, 
    1020.7, 1020.7, 1020.7, 1020.9, 1021, 1021, 1021.1, 1021.1, 1021.1, 1021, 
    1020.8, 1020.6, 1020.3, 1019.9, 1019.7, 1019.5, 1019.6, 1019.3, 1019.1, 
    1018.8, 1018.3, 1018.1, 1017.8, 1017.3, 1017, 1016.7, 1016.6, 1016.6, 
    1016.5, 1016.5, 1016.5, 1016.3, 1016.4, 1016.3, 1016.1, 1016, 1015.8, 
    1015.7, 1015.6, 1015.3, 1015.3, 1015.1, 1015, 1015, 1014.8, 1014.7, 
    1014.4, 1014.2, 1014, 1013.7, 1013.5, 1013.3, 1013.3, 1013.3, 1013.1, 
    1013, 1012.7, 1012.2, 1011.9, 1011.7, 1011.4, 1011.3, 1011.2, 1011.3, 
    1011, 1010.9, 1010.6, 1010.4, 1009.9, 1009.3, 1008.9, 1008.4, 1007.9, 
    1007.5, 1007, 1006.6, 1006.2, 1006.2, 1005.9, 1005.6, 1005.2, 1004.8, 
    1004.9, 1004.9, 1004.5, 1004.2, 1003.9, 1003.6, 1003.1, 1003.1, 1003, 
    1002.7, 1002.5, 1002.3, 1002.1, 1002, 1001.9, 1001.9, 1001.6, 1001.6, 
    1001.4, 1001.1, 1000.9, 1000.7, 1000.4, 1000, 999.8, 999.5, 999.4, 999.1, 
    999, 998.8, 998.5, 998.3, 998.1, 997.8, 997.6, 997.4, 996.9, 996.5, 
    996.2, 995.6, 995.3, 995, 994.9, 994.6, 994.4, 994.2, 993.9, 993.8, 
    993.6, 993.5, 993.4, 993.2, 993, 993, 993, 993, 993.2, 993.2, 993.3, 
    993.5, 993.6, 993.8, 994, 994.3, 994.5, 994.7, 994.9, 995.1, 995.4, 
    995.9, 996.1, 996.2, 996.2, 996, 995.9, 996.1, 996, 996, 995.9, 995.8, 
    995.8, 995.8, 995.5, 995.2, 995.2, 995.1, 995, 994.7, 994.8, 995.1, 995, 
    995.1, 995.1, 995.5, 996.3, 997.3, 998.6, 999.8, 1001.4, 1002.6, 1003.6, 
    1004.8, 1005.7, 1006.7, 1007.8, 1008.7, 1009.1, 1009.5, 1009.5, 1009.9, 
    1010, 1010.1, 1010.1, 1010.3, 1010.3, 1010.6, 1010.7, 1010.9, 1011, 
    1011.4, 1011.7, 1011.9, 1012.2, 1012.4, 1012.6, 1012.9, 1013, 1013.3, 
    1013.6, 1013.6, 1013.8, 1014, 1014.1, 1014.3, 1014.3, 1014.2, 1014.4, 
    1014.8, 1014.9, 1015.2, 1015.4, 1015.4, 1015.3, 1015.1, 1015, 1015, 1015, 
    1014.9, 1015, 1015, 1015.1, 1015.2, 1015.1, 1015, 1015.2, 1015, 1014.9, 
    1014.9, 1014.7, 1014.6, 1014.6, 1014.6, 1014.6, 1014.4, 1014.3, 1014.1, 
    1013.7, 1013.5, 1012.9, 1012.8, 1012.6, 1012.3, 1012.3, 1012.3, 1012.1, 
    1012.1, 1011.9, 1011.9, 1011.8, 1011.7, 1011.3, 1010.9, 1010.5, 1010.4, 
    1010.3, 1010.3, 1010.3, 1010.3, 1010, 1010, 1009.8, 1009.8, 1009.4, 
    1009.2, 1009.2, 1008.9, 1008.8, 1008.6, 1008.8, 1008.8, 1008.7, 1008.7, 
    1008.7, 1008.7, 1008.6, 1008.4, 1008.3, 1008.3, 1008.3, 1008.3, 1008.4, 
    1008.5, 1008.7, 1008.7, 1008.7, 1008.8, 1008.6, 1008.4, 1008.2, 1008.1, 
    1008, 1008.3, 1008.5, 1008.9, 1009, 1009.2, 1009.5, 1009.8, 1010.1, 
    1010.4, 1010.4, 1010.8, 1011.1, 1011.3, 1011.8, 1012.2, 1012.7, 1013.2, 
    1013.5, 1013.7, 1013.9, 1014, 1014.2, 1014.4, 1014.6, 1014.9, 1015.2, 
    1015.6, 1016, 1016.1, 1016.5, 1016.7, 1016.7, 1016.6, 1016.8, 1017, 
    1017.2, 1017.1, 1017.2, 1017.5, 1017.7, 1017.8, 1018, 1018.1, 1018, 
    1018.1, 1018.1, 1018, 1018.1, 1018, 1018.1, 1018.4, 1018.3, 1018.4, 
    1018.5, 1018.6, 1018.5, 1018.4, 1018.4, 1018.5, 1018.5, 1018.4, 1018.4, 
    1018.3, 1018.1, 1017.6, 1017.4, 1016.9, 1016.5, 1016, 1015.8, 1015.6, 
    1015.5, 1015, 1014.6, 1014.1, 1013.8, 1013.5, 1013.4, 1013.1, 1012.7, 
    1012.5, 1011.7, 1011.4, 1011, 1010.8, 1010.8, 1010.7, 1010.3, 1009.7, 
    1009.7, 1009.5, 1009.5, 1009, 1008.7, 1008.3, 1008.3, 1008.2, 1008, 
    1007.9, 1007.6, 1007.4, 1007.2, 1006.7, 1006.2, 1006, 1005.7, 1005.5, 
    1005.3, 1005.2, 1005.1, 1004.7, 1004.6, 1004.5, 1004.6, 1004.8, 1004.7, 
    1005, 1005.1, 1005.4, 1005.8, 1006.1, 1006.4, 1006.6, 1007, 1007, 1006.9, 
    1006.8, 1006.9, 1006.9, 1006.8, 1006.5, 1006.3, 1006.3, 1006.5, 1006.6, 
    1006.6, 1006.4, 1006.3, 1006.1, 1006, 1005.6, 1005.2, 1004.8, 1004.5, 
    1004.1, 1003.5, 1002.9, 1002.5, 1001.9, 1001.3, 1000.8, 1000.2, 999.9, 
    999.4, 999.2, 999.1, 998.7, 998.7, 998.6, 998.4, 998.1, 997.9, 997.5, 
    997.5, 997.2, 997.1, 996.9, 996.5, 996.2, 995.9, 995.8, 995.5, 995.4, 
    995.4, 995.3, 995, 994.8, 994.6, 994.6, 994.5, 994.4, 994.5, 994.3, 
    994.2, 994.2, 993.9, 993.5, 993.1, 992.5, 992.2, 991.8, 991.4, 991.2, 
    990.9, 990.4, 990, 989.5, 989.3, 988.9, 988.7, 988.4, 988.3, 988.3, 
    988.5, 988.4, 988.9, 989.3, 989.7, 990, 990.4, 990.8, 991.3, 991.6, 
    991.5, 992, 992.3, 992.6, 992.9, 993.2, 993.5, 994.1, 994.6, 995, 995.2, 
    995.7, 996.2, 996.8, 997.2, 997.9, 998.5, 999.3, 999.8, 1000.6, 1001.4, 
    1001.8, 1002.5, 1002.9, 1003.3, 1003.8, 1004.1, 1004.6, 1004.9, 1005.5, 
    1005.9, 1006, 1006.3, 1006.8, 1006.9, 1007, 1007.2, 1007.2, 1007.3, 
    1007.4, 1007.8, 1007.7, 1007.7, 1007.7, 1007.5, 1007.6, 1007.6, 1007.5, 
    1007.5, 1007.4, 1007.5, 1007.5, 1007.7, 1007.8, 1007.7, 1007.7, 1007.8, 
    1007.8, 1007.8, 1007.8, 1007.8, 1007.9, 1007.8, 1007.8, 1007.7, 1007.8, 
    1007.8, 1007.8, 1007.9, 1007.9, 1007.6, 1007.4, 1007.2, 1007, 1006.8, 
    1006.5, 1006.2, 1005.7, 1005.4, 1005.3, 1004.8, 1003.9, 1002.9, 1001.9, 
    1001.2, 1000.6, 1000.2, 999.7, 999.4, 999.4, 999, 998.4, 998, 997.5, 
    997.1, 996.6, 996.7, 996.7, 997.3, 998.4, 1000.1, 1001, 1001.9, 1003, 
    1003.9, 1004.6, 1005.5, 1006.3, 1007.1, 1008, 1008.9, 1009.7, 1010.7, 
    1011.7, 1012.7, 1013.5, 1014.1, 1014.8, 1015.3, 1015.7, 1016.3, 1016.8, 
    1017.6, 1018.4, 1019, 1019.6, 1020.2, 1020.6, 1020.9, 1020.7, 1020.8, 
    1021.1, 1021.3, 1021.3, 1021.8, 1021.9, 1022.1, 1022.7, 1022.8, 1022.9, 
    1022.9, 1022.9, 1022.6, 1022.6, 1022.6, 1022.4, 1022.3, 1022.6, 1022.6, 
    1022.7, 1022.8, 1022.8, 1022.7, 1022.7, 1022.6, 1022.4, 1022.3, 1022.4, 
    1022, 1022, 1022, 1022.3, 1022.3, 1022.1, 1021.7, 1021.4, 1021.3, 1020.9, 
    1020.5, 1019.9, 1019.6, 1019.4, 1019.1, 1019, 1018.8, 1018.5, 1018, 
    1017.9, 1017.6, 1017.2, 1016.8, 1016.6, 1016.6, 1016.7, 1016.5, 1016.5, 
    1016.1, 1015.7, 1015.4, 1015.2, 1015.1, 1015, 1015, 1014.9, 1014.9, 
    1014.9, 1015.1, 1015.3, 1015.5, 1015.4, 1015.9, 1016.1, 1016.3, 1016.3, 
    1016.5, 1017, 1017.4, 1017.6, 1018, 1018.2, 1018.4, 1018.7, 1018.9, 
    1019.1, 1019.5, 1019.5, 1019.4, 1019.3, 1018.9, 1018.9, 1019, 1019.1, 
    1019.1, 1019.1, 1019, 1019.3, 1019.5, 1019.9, 1019.9, 1020.1, 1020.3, 
    1020.6, 1020.7, 1020.4, 1020.1, 1020.1, 1020.3, 1020.3, 1020.2, 1020, 
    1019.8, 1019.6, 1019.3, 1019.2, 1018.9, 1018.6, 1018.3, 1018.4, 1018.2, 
    1018, 1017.9, 1017.8, 1017.4, 1017.2, 1017, 1017, 1017, 1016.8, 1016.8, 
    1016.4, 1016.3, 1016, 1015.9, 1015.9, 1015.9, 1015.8, 1015.7, 1015.1, 
    1014.9, 1014.8, 1014.9, 1014.7, 1014.5, 1014, 1013.8, 1013.5, 1013.2, 
    1013.2, 1013.2, 1013.2, 1013, 1013, 1012.7, 1012.6, 1012.6, 1012.6, 
    1012.4, 1012.3, 1012.5, 1012.3, 1012.3, 1012, 1012.3, 1012, 1012.4, 
    1012.4, 1011.8, 1011.9, 1011.6, 1011.3, 1011.4, 1011.3, 1011.3, 1011.5, 
    1011.7, 1012.1, 1012.3, 1012.6, 1012.8, 1013.1, 1013.1, 1013.4, 1013.6, 
    1013.8, 1014, 1014, 1014.4, 1014.7, 1015, 1015.6, 1015.6, 1015.6, 1015.8, 
    1015.9, 1016.3, 1016.8, 1017, 1016.9, 1017.3, 1017.7, 1018.1, 1018.4, 
    1018.6, 1018.8, 1019.1, 1019.3, 1019.7, 1020.3, 1020.2, 1020.7, 1021, 
    1021.1, 1021.4, 1021.8, 1022.1, 1022.1, 1022.3, 1022.5, 1022.6, 1022.8, 
    1022.9, 1023.1, 1023.1, 1023, 1023, 1022.9, 1022.6, 1022.7, 1022.5, 
    1022.2, 1022, 1022, 1021.7, 1021.4, 1021, 1020.8, 1020.6, 1020.3, 1020, 
    1019.9, 1019.6, 1019.6, 1019.3, 1019.3, 1019.1, 1018.9, 1018.6, 1018.6, 
    1018.7, 1018.8, 1018.5, 1018.4, 1018, 1017.9, 1017.8, 1017.8, 1017.5, 
    1017.4, 1017.3, 1017.2, 1016.8, 1016.6, 1016.3, 1016, 1015.4, 1015.1, 
    1014.5, 1014.4, 1014, 1013.6, 1013.2, 1012.9, 1012.7, 1012.5, 1011.8, 
    1011.2, 1010.4, 1009.8, 1009.4, 1008.8, 1008.2, 1007.8, 1007.5, 1007.1, 
    1006.9, 1006.7, 1006.6, 1006.6, 1006.7, 1007, 1007.2, 1007.8, 1008.2, 
    1008.7, 1009.4, 1009.6, 1010.2, 1010.6, 1011.1, 1011.7, 1012, 1012.7, 
    1013, 1013.4, 1013.7, 1013.9, 1014, 1014.3, 1014.5, 1014.8, 1015.2, 
    1015.1, 1014.8, 1014.4, 1014.1, 1013.7, 1013.9, 1013.9, 1013.7, 1013.3, 
    1012.8, 1012.3, 1012.1, 1011.8, 1011.5, 1011.5, 1011.3, 1011, 1011.2, 
    1011.5, 1011.7, 1011.9, 1012, 1011.9, 1011.9, 1011.6, 1011.7, 1011.6, 
    1011.4, 1011.6, 1012, 1012.3, 1013.1, 1014.3, 1015.5, 1016.8, 1018.1, 
    1019.5, 1020.5, 1021.8, 1023, 1023.9, 1024.8, 1025.7, 1026.4, 1027, 
    1027.7, 1028.5, 1029.1, 1029.5, 1030, 1030.2, 1030.3, 1030.6, 1030.4, 
    1030.8, 1030.9, 1031, 1031.4, 1031.3, 1031.2, 1031, 1030.8, 1030.4, 
    1030.3, 1030.1, 1030, 1029.9, 1029.8, 1029.8, 1029.9, 1029.8, 1029.8, 
    1029.6, 1029.5, 1029.2, 1029.3, 1029.1, 1029, 1029, 1028.8, 1028.8, 
    1028.7, 1028.8, 1028.7, 1028.4, 1028.1, 1027.6, 1027.2, 1026.8, 1026.4, 
    1026, 1025.7, 1025.2, 1024.7, 1024.3, 1023.6, 1022.9, 1022.4, 1021.8, 
    1021.2, 1020.6, 1019.9, 1019.5, 1018.9, 1018.7, 1018.5, 1018.3, 1018.2, 
    1017.8, 1017.7, 1017.6, 1017.5, 1017.2, 1017.1, 1017.2, 1017.1, 1017, 
    1016.7, 1016.5, 1016.2, 1015.5, 1014.4, 1013.5, 1011.7, 1010.7, 1009.9, 
    1010.1, 1010.1, 1010.4, 1010.6, 1010.4, 1010.4, 1009.7, 1009.1, 1009.1, 
    1008.8, 1008.8, 1009.9, 1010.1, 1011, 1011.8, 1013.1, 1014, 1014.7, 
    1015.8, 1016.6, 1017.4, 1018, 1018.7, 1019.4, 1020.5, 1021.4, 1022.4, 
    1023.5, 1024.5, 1025, 1025.8, 1026.7, 1027.1, 1027.4, 1028, 1028.5, 
    1028.8, 1028.9, 1028.8, 1028.8, 1028.3, 1028.1, 1027.4, 1026.5, 1025.8, 
    1025.6, 1025.5, 1025.2, 1025, 1025.1, 1024.9, 1025.1, 1024.9, 1024.5, 
    1023.7, 1023.3, 1022.3, 1021.1, 1020, 1019.8, 1019, 1018.5, 1019, 1018.4, 
    1018.6, 1018.5, 1018.4, 1018.9, 1019.4, 1019.7, 1019.9, 1020.3, 1020.7, 
    1020.8, 1021.2, 1021.9, 1022.5, 1022.7, 1023, 1023.1, 1023, 1023.1, 
    1023.5, 1023.8, 1023.8, 1024, 1024.1, 1024, 1024.1, 1023.8, 1023.5, 
    1023.2, 1023.5, 1023.8, 1024.1, 1024.3, 1024.9, 1025.3, 1025.5, 1025.9, 
    1025.8, 1025.7, 1025.6, 1025.9, 1025.9, 1025.9, 1026.2, 1026.3, 1026.5, 
    1026.8, 1027, 1027.2, 1027.4, 1027.6, 1027.7, 1027.8, 1027.7, 1027.4, 
    1027.7, 1028.1, 1028.3, 1029, 1029.7, 1029.8, 1029.3, 1029.1, 1029.1, 
    1029, 1029, 1029, 1029.1, 1029.3, 1029.2, 1029.1, 1029.2, 1029.3, 1029.5, 
    1029.5, 1029.6, 1029.7, 1029.4, 1029.6, 1028.9, 1029, 1028.9, 1028.6, 
    1028.3, 1027.9, 1027.4, 1027, 1026.6, 1026.3, 1026.1, 1026, 1026.1, 
    1026.1, 1026.2, 1025.9, 1025.6, 1025.5, 1025.3, 1025.3, 1025.2, 1025.1, 
    1025.4, 1025.5, 1025.7, 1025.9, 1026.4, 1026.7, 1026.7, 1026.4, 1026.7, 
    1026.8, 1026.9, 1026.9, 1026.9, 1027, 1027, 1026.9, 1026.7, 1026.2, 
    1026.1, 1025.5, 1025.3, 1025.1, 1025.1, 1024.5, 1024.3, 1024.1, 1023.5, 
    1023.8, 1023.8, 1023.6, 1023.1, 1022.6, 1022.2, 1022, 1021.4, 1021, 
    1020.9, 1020.8, 1021.1, 1020.7, 1020.3, 1020.3, 1020.1, 1019.8, 1019.3, 
    1018.9, 1018.6, 1018.2, 1017.8, 1017.1, 1016.4, 1015.7, 1015.3, 1014.9, 
    1014.5, 1014, 1013.5, 1012.9, 1012, 1011.3, 1010.6, 1010, 1009.6, 1009.1, 
    1008.7, 1008.1, 1007.8, 1007.8, 1007.3, 1006.4, 1005.4, 1004.8, 1004.9, 
    1005, 1004.8, 1004.3, 1003.4, 1003.4, 1003.6, 1003, 1002.8, 1002.5, 
    1002.3, 1002.1, 1001.9, 1001.8, 1001.5, 1001.4, 1001.3, 1001.1, 1001.1, 
    1001, 1001, 1000.8, 1000.6, 1000.2, 1000, 1000, 999.9, 999.9, 1000.1, 
    999.9, 999.8, 999.8, 999.9, 1000, 1000.1, 1000.1, 1000.4, 1000.7, 1000.9, 
    1001, 1001.1, 1001.5, 1001.7, 1001.9, 1002, 1002.2, 1002, 1002, 1002, 
    1002.1, 1002.2, 1002.5, 1002.8, 1003.1, 1003.2, 1003.6, 1003.5, 1003.6, 
    1003.8, 1004, 1004.2, 1004.4, 1004.8, 1005, 1005.3, 1005.7, 1005.9, 
    1006.4, 1006.8, 1007.1, 1007.5, 1007.8, 1008.2, 1008.4, 1008.6, 1009.1, 
    1009.6, 1010.1, 1010.5, 1010.8, 1011.2, 1011.6, 1011.9, 1012.4, 1012.7, 
    1012.9, 1013.2, 1013.5, 1013.7, 1013.9, 1014.1, 1014.1, 1014.1, 1014.3, 
    1014.3, 1014.3, 1014.4, 1014.5, 1014.6, 1014.7, 1014.9, 1015, 1015.2, 
    1015.3, 1015.4, 1015.4, 1015.7, 1015.7, 1015.8, 1015.8, 1015.7, 1015.9, 
    1015.8, 1015.9, 1016, 1016.1, 1016.1, 1016, 1015.9, 1015.9, 1016, 1015.9, 
    1015.7, 1015.7, 1015.9, 1016.1, 1016.2, 1016.1, 1016.2, 1016.2, 1016.1, 
    1015.9, 1015.7, 1015.8, 1015.7, 1015.6, 1015.6, 1015.6, 1015.8, 1015.6, 
    1015.3, 1015.2, 1015.2, 1015.1, 1015, 1015.1, 1014.8, 1014.8, 1014.7, 
    1014.8, 1015.3, 1015.8, 1016, 1016.3, 1016.5, 1016.8, 1017, 1017.3, 
    1017.3, 1017.5, 1017.7, 1017.8, 1017.8, 1017.8, 1017.7, 1017.7, 1017.6, 
    1017.4, 1017.4, 1017.4, 1017.3, 1017.4, 1017.2, 1017.5, 1017.8, 1018.1, 
    1018.2, 1018.1, 1018.1, 1018.1, 1018.1, 1018.2, 1018.1, 1018.2, 1018.2, 
    1018.3, 1018.5, 1018.5, 1018.3, 1018.2, 1017.9, 1017.9, 1017.9, 1017.8, 
    1017.9, 1018, 1017.8, 1018, 1018.1, 1017.9, 1017.8, 1017.6, 1017.6, 
    1017.5, 1017.3, 1017.2, 1017.3, 1017.2, 1017.2, 1017.1, 1017, 1016.9, 
    1016.9, 1016.6, 1016.3, 1015.9, 1015.8, 1015.6, 1015.5, 1015.5, 1015.4, 
    1015.5, 1015.8, 1016, 1015.9, 1015.7, 1015.6, 1015.5, 1015.4, 1015.2, 
    1015.1, 1015, 1014.9, 1014.7, 1014.5, 1014.4, 1014.2, 1014.3, 1014.4, 
    1014.4, 1014.3, 1014.3, 1014.4, 1014.5, 1014.8, 1015, 1015.3, 1015.3, 
    1015.2, 1014.7, 1014.6, 1014.4, 1014, 1013.8, 1013.8, 1013.4, 1013.4, 
    1013.5, 1013.4, 1013.3, 1013, 1012.8, 1012.4, 1012.3, 1012, 1011.6, 1012, 
    1011.7, 1011.9, 1011.7, 1011.5, 1011.7, 1011.7, 1011.6, 1011.7, 1011.3, 
    1010.9, 1010.7, 1010.9, 1010.5, 1010.6, 1010.7, 1010.9, 1011, 1011.2, 
    1011.3, 1011.6, 1011.7, 1011.8, 1011.5, 1011.8, 1012, 1012.1, 1012.4, 
    1012.4, 1012.6, 1012.5, 1012.3, 1012.3, 1012, 1011.8, 1011.6, 1011.3, 
    1011, 1010.6, 1010.5, 1010.3, 1010.1, 1009.7, 1009.6, 1009.2, 1008.8, 
    1008.1, 1008.1, 1007.9, 1007.7, 1007.6, 1007.5, 1007.6, 1007.5, 1007.5, 
    1007.2, 1007.2, 1007.2, 1007.3, 1007.5, 1007.6, 1007.9, 1008.2, 1008.4, 
    1008.6, 1008.6, 1008.6, 1008.9, 1008.9, 1009.2, 1009.4, 1009.8, 1010.2, 
    1010.7, 1011.1, 1011.6, 1012, 1012.1, 1012.4, 1012.7, 1013, 1013.3, 
    1013.5, 1013.8, 1014, 1014.5, 1014.9, 1015, 1015.2, 1015.5, 1015.8, 
    1016.1, 1016.3, 1016.6, 1016.8, 1017.2, 1017.5, 1017.9, 1018.1, 1018.5, 
    1018.8, 1019.1, 1019.4, 1019.6, 1019.8, 1019.9, 1020, 1020, 1020.1, 
    1020.2, 1020.2, 1020.2, 1020.4, 1020.4, 1020.2, 1020.2, 1020.2, 1020.3, 
    1020.1, 1020.1, 1019.9, 1019.9, 1019.9, 1019.8, 1019.8, 1019.9, 1019.7, 
    1019.5, 1019.4, 1019.1, 1018.5, 1018.1, 1017.6, 1017.1, 1016.6, 1016.3, 
    1015.9, 1015.3, 1014.8, 1014.4, 1014, 1013.9, 1013.5, 1013.5, 1013.3, 
    1013.4, 1013.4, 1013.7, 1013.9, 1014.2, 1014.5, 1014.7, 1015, 1015.2, 
    1015.4, 1015.6, 1016, 1015.9, 1016.3, 1016.3, 1016.6, 1016.8, 1016.8, 
    1017, 1016.9, 1017.1, 1017.1, 1017.2, 1017.4, 1017.3, 1017.6, 1017.8, 
    1017.8, 1017.8, 1017.8, 1018.1, 1018.1, 1018.1, 1018.4, 1018.4, 1018.4, 
    1018.7, 1018.9, 1019, 1019.4, 1019.5, 1019.7, 1019.4, 1019.6, 1019.7, 
    1019.7, 1019.6, 1019.2, 1019, 1018.7, 1018.3, 1018.2, 1017.7, 1017.3, 
    1017, 1016.1, 1015.6, 1015.3, 1014.6, 1014, 1013.4, 1013, 1012.4, 1011.8, 
    1011.8, 1011.4, 1010.7, 1009.9, 1009.9, 1009.6, 1009.4, 1009.3, 1009, 
    1008.4, 1008, 1007.7, 1007.4, 1007.4, 1006.9, 1006.7, 1006.9, 1007.2, 
    1007.4, 1007.9, 1008.4, 1008.7, 1009.2, 1009.8, 1010.3, 1010.6, 1011, 
    1011.5, 1011.8, 1011.6, 1011.7, 1011.6, 1011.4, 1011.5, 1011.5, 1011.2, 
    1011, 1010.5, 1009.9, 1009.7, 1009.1, 1008.6, 1007.9, 1007.6, 1007.2, 
    1007, 1007, 1006.9, 1006.5, 1006.5, 1006.3, 1006.4, 1006.3, 1006.4, 1006, 
    1006.2, 1006.2, 1006.2, 1006.2, 1006.4, 1006.4, 1006.6, 1006.7, 1006.1, 
    1005.8, 1005.9, 1005.7, 1005.3, 1005.2, 1005.5, 1005.5, 1005.4, 1005.3, 
    1004.9, 1004.3, 1004.2, 1004, 1003.9, 1003.1, 1002.4, 1001.5, 1001.2, 
    1000.6, 1000.1, 999.1, 998, 997, 996.2, 995.4, 994.5, 993.9, 992.9, 992, 
    991, 990, 988.9, 988.3, 987.8, 987.1, 986.3, 985.6, 984.9, 984.8, 984.7, 
    984.9, 985, 984.9, 985, 985.2, 985.4, 985.3, 985.4, 985.4, 985.8, 986, 
    986.3, 986.3, 986.5, 986.7, 987.3, 987.4, 987.3, 987.3, 987.5, 988.1, 
    988.5, 988.4, 988.8, 989.2, 989.4, 989.9, 990.2, 990.7, 991.2, 991.7, 
    991.8, 991.5, 991.7, 991.6, 991.3, 991.8, 992, 992.7, 993.2, 993.5, 
    993.5, 993.1, 993.5, 995.2, 993.9, 995.3, 995.3, 996.3, 996.3, 996.3, 
    996.5, 996.9, 996.9, 995.9, 995.1, 995.8, 995.3, 995.3, 995.9, 995.4, 
    995.9, 996.3, 996.9, 996.7, 996.8, 996.3, 996.1, 996, 995.9, 995.8, 
    995.5, 995.6, 995.7, 995.8, 995.8, 996.7, 996.8, 997, 996.9, 996.9, 
    996.9, 996.9, 997.1, 997, 997, 997.1, 996.8, 996.5, 996.5, 996.3, 996.2, 
    996.4, 996.3, 996.3, 996.2, 996.3, 996.6, 996.7, 996.9, 997.2, 997.5, 
    997.6, 997.5, 997.5, 997.4, 997.5, 997.7, 997.7, 997.5, 997.5, 997.4, 
    997.6, 997.7, 997.6, 997.3, 997.2, 997.1, 997, 997, 996.8, 996.8, 996.8, 
    996.9, 996.8, 996.5, 996.3, 995.9, 995.5, 994.9, 994.6, 994.2, 993.9, 
    993.5, 993, 992.5, 991.8, 991.6, 991.3, 990.7, 989.9, 989.6, 989.3, 
    988.8, 988.5, 988.2, 987.8, 987.6, 987.2, 986.2, 986.2, 985.9, 985.6, 
    985.2, 984.8, 984.6, 984.3, 984.1, 983.8, 983.7, 983.5, 983.5, 983.2, 
    982.8, 982.7, 982.7, 982.5, 982.5, 982.6, 982.7, 982.9, 983.1, 983.2, 
    983.2, 983.3, 983.1, 983.1, 983.1, 982.6, 982.6, 982.2, 982.5, 982.5, 
    982.5, 982.5, 982.5, 982.8, 982.9, 983.3, 983.7, 984.2, 984.8, 985.9, 
    987.2, 988.9, 990.1, 991, 991.7, 992.8, 993.9, 994.5, 995.1, 995.5, 
    996.5, 997, 997.5, 997.9, 998.7, 999.2, 999.7, 999.7, 1000.5, 1000.4, 
    1000.6, 1001, 1001.5, 1001.9, 1002.3, 1003.1, 1003.9, 1004.6, 1004.9, 
    1005.5, 1005.8, 1006.4, 1006.9, 1007.5, 1007.6, 1008.1, 1008.6, 1009, 
    1009.5, 1009.8, 1010.1, 1010.3, 1010.7, 1011.2, 1011.5, 1011.8, 1012, 
    1012.4, 1012.8, 1013.2, 1013.5, 1013.8, 1014.3, 1014.4, 1014.7, 1015, 
    1015.3, 1015.8, 1016, 1016.4, 1016.8, 1017.1, 1017.5, 1017.9, 1018, 
    1018.2, 1018.5, 1018.8, 1019.3, 1019.6, 1019.8, 1020.1, 1020.4, 1020.8, 
    1021.2, 1021.8, 1022.2, 1022.2, 1022.6, 1022.7, 1022.8, 1022.8, 1022.7, 
    1022.8, 1022.8, 1022.4, 1022.2, 1022.1, 1021.8, 1021.9, 1021.2, 1020.7, 
    1020.4, 1019.8, 1019.5, 1018.9, 1018.2, 1018.4, 1018, 1017.2, 1016.9, 
    1016.6, 1016.2, 1015.7, 1015.1, 1014.1, 1013.5, 1012.7, 1011.9, 1011.7, 
    1011.7, 1011, 1010.3, 1010.1, 1009.1, 1008.6, 1008, 1007.5, 1006.7, 1006, 
    1006.2, 1006.1, 1005.6, 1005.4, 1005.1, 1004.9, 1004.5, 1004.6, 1004.7, 
    1004.9, 1004.8, 1004.5, 1004.2, 1004.2, 1004.4, 1004, 1004.1, 1003.8, 
    1003.6, 1004.3, 1004.8, 1005.4, 1006, 1006.1, 1005.8, 1005.4, 1005.2, 
    1005, 1005, 1005.3, 1005.4, 1004.7, 1004.5, 1004.6, 1004.3, 1004.3, 
    1003.9, 1003.8, 1003.3, 1003, 1003, 1002.9, 1002.9, 1002.4, 1001.7, 
    1001.4, 1001.2, 1000.5, 1000.5, 999.8, 1000, 1000.2, 1000.1, 1000.2, 
    1000.2, 1000.2, 1000.1, 999.7, 999.4, 999.6, 999.7, 999.9, 1000, 999.9, 
    1000.1, 1000.2, 1000.2, 1000, 1000, 999.9, 999.8, 999.7, 999.9, 1000.3, 
    1000.6, 1000.8, 1001.1, 1000.8, 1000.9, 1001.2, 1001.2, 1001.3, 1001.5, 
    1001.6, 1001.6, 1001.7, 1001.7, 1001.9, 1002.3, 1002.3, 1002.5, 1002.6, 
    1002.8, 1002.8, 1002.9, 1003, 1003.1, 1003.3, 1003.4, 1003.3, 1003.3, 
    1003.6, 1003.7, 1003.8, 1003.7, 1003.7, 1003.9, 1004.1, 1004.2, 1004.5, 
    1004.6, 1004.6, 1004.8, 1005, 1005.2, 1005.3, 1005.4, 1005.7, 1005.8, 
    1006.1, 1006.2, 1006.4, 1006.6, 1006.9, 1006.9, 1006.9, 1007.3, 1007.4, 
    1007.5, 1007.5, 1007.4, 1007.4, 1007.5, 1007.4, 1007.4, 1007.6, 1007.8, 
    1008.2, 1008.5, 1008.5, 1008.8, 1008.8, 1008.8, 1009.4, 1009.7, 1010, 
    1010.3, 1010.7, 1011, 1011.4, 1011.8, 1012, 1012.1, 1012.1, 1012, 1012.3, 
    1012.8, 1013.1, 1013.2, 1013.6, 1013.7, 1014, 1014.1, 1014.2, 1014.2, 
    1014.4, 1014.5, 1014.5, 1014.9, 1015.2, 1015.5, 1015.5, 1015.4, 1015.3, 
    1015.3, 1015.4, 1015.4, 1015.5, 1015.4, 1015.7, 1015.7, 1015.9, 1016, 
    1015.9, 1015.8, 1015.7, 1015.7, 1015.8, 1015.9, 1015.7, 1015.5, 1015.4, 
    1015.2, 1015.2, 1015.1, 1014.9, 1014.8, 1014.7, 1014.6, 1014.3, 1014.5, 
    1014.7, 1014.7, 1014.7, 1015, 1015.1, 1015.2, 1015.4, 1015.4, 1015.4, 
    1015.6, 1015.4, 1015.7, 1015.8, 1016.1, 1016.5, 1017.6, 1017.5, 1018.2, 
    1018.6, 1019.1, 1019.7, 1020, 1020.2, 1020.6, 1020.7, 1020.9, 1021.1, 
    1021.5, 1021.9, 1022.4, 1022.5, 1022.9, 1023, 1023.3, 1023.2, 1023.3, 
    1023.4, 1023.7, 1023.9, 1024.2, 1024.6, 1025, 1025.4, 1025.6, 1026, 1026, 
    1026.3, 1026.2, 1026.1, 1026, 1026.2, 1026.4, 1026.8, 1027.1, 1027.4, 
    1027.5, 1027.7, 1027.8, 1028.2, 1028.4, 1028.5, 1028.4, 1028.8, 1029.6, 
    1030, 1030.3, 1030.5, 1030.8, 1031.1, 1031.6, 1032, 1032.5, 1032.8, 
    1033.3, 1033.5, 1033.9, 1034.5, 1035, 1035.3, 1035.4, 1035.4, 1035.5, 
    1035.7, 1035.8, 1036.2, 1036.5, 1036.8, 1037.4, 1037.7, 1038, 1038.5, 
    1038.3, 1038.2, 1038, 1038, 1037.5, 1037.5, 1037.2, 1037.1, 1037.4, 
    1037.5, 1037.6, 1037.7, 1037.7, 1037.3, 1037.2, 1037, 1036.9, 1036.9, 
    1036.7, 1036.8, 1036.9, 1037.1, 1037.4, 1037.8, 1037.8, 1038, 1038.2, 
    1038.2, 1038.1, 1038.2, 1038.4, 1038.6, 1038.8, 1038.6, 1038.6, 1038.4, 
    1038.3, 1038.1, 1037.8, 1038.1, 1037.9, 1037.3, 1037.2, 1037.1, 1037.3, 
    1037.3, 1037.1, 1036.9, 1036.5, 1036.1, 1036.1, 1036.2, 1035.7, 1035.4, 
    1035.2, 1035.1, 1034.7, 1034.6, 1034.1, 1033.8, 1033.5, 1033.1, 1032.9, 
    1032.7, 1032.5, 1031.8, 1031.7, 1031.6, 1031.4, 1031.3, 1031.2, 1030.7, 
    1030.5, 1030.1, 1029.8, 1029.5, 1029.3, 1029, 1028.9, 1028.5, 1028.3, 
    1027.8, 1027.6, 1027.2, 1026.8, 1026.4, 1026.1, 1025.4, 1025.1, 1024.6, 
    1024, 1023.5, 1023, 1022.7, 1022.6, 1022.3, 1021.7, 1021, 1020.1, 1019.6, 
    1019.1, 1018.6, 1018.3, 1017.8, 1017.4, 1017, 1016.4, 1016, 1015.7, 
    1015.1, 1014.6, 1014, 1013.5, 1012.9, 1012.2, 1011.8, 1011.5, 1011.1, 
    1010.8, 1010.4, 1009.9, 1009.3, 1008.7, 1008.2, 1007.8, 1007.3, 1006.8, 
    1006.4, 1006.1, 1006, 1005.6, 1005.2, 1004.9, 1004.2, 1003.7, 1003.4, 
    1003.1, 1002.8, 1002.9, 1003.1, 1003.2, 1003.7, 1004.1, 1004.5, 1004.6, 
    1005, 1005.2, 1005.6, 1005.8, 1006.1, 1006.4, 1006.8, 1007.2, 1007.6, 
    1008, 1008.2, 1008.3, 1008.7, 1009, 1009.5, 1009.8, 1009.7, 1009.9, 1010, 
    1010.2, 1010.4, 1010.6, 1010.5, 1010.5, 1010.6, 1011.2, 1011.3, 1011.2, 
    1011.4, 1011.7, 1012.4, 1013, 1013, 1013.2, 1013.3, 1013.5, 1013.5, 
    1013.4, 1013.3, 1013.3, 1013.2, 1013.2, 1013, 1012.7, 1012.7, 1013, 1013, 
    1012.9, 1012.7, 1012.7, 1012.7, 1012.8, 1012.9, 1012.9, 1012.9, 1012.9, 
    1012.6, 1012.4, 1012.4, 1012.2, 1011.9, 1011.4, 1011, 1010.5, 1010.2, 
    1010, 1009.6, 1009.2, 1008.6, 1008.5, 1008.4, 1007.8, 1006.6, 1005.8, 
    1004.8, 1003.9, 1003.6, 1003.1, 1002.2, 1001.2, 1000.2, 998.9, 998, 
    997.1, 995.8, 994.6, 993.8, 993.3, 992.7, 992.9, 992.7, 992.6, 992.9, 
    992.9, 992.6, 992.3, 992.2, 991.9, 991.5, 991.2, 990.8, 990.6, 990.3, 
    990.6, 990.4, 990.4, 990.4, 990.4, 990.2, 990.1, 990, 989.9, 990.1, 990, 
    989.7, 989.6, 989.4, 989.3, 989.2, 988.9, 988.3, 988.4, 987.9, 987.4, 
    987.5, 987, 986.7, 986.6, 986.4, 986.5, 986.6, 986.5, 986.4, 986.2, 
    985.9, 985.8, 985.5, 985.5, 985.3, 985.5, 985.6, 985.8, 985.7, 985.5, 
    985.7, 985.6, 986.2, 986.5, 987, 988.2, 988.9, 990, 990.5, 991.3, 992.3, 
    993, 994.3, 995.1, 995.7, 996.2, 996.7, 997.4, 997.7, 998.2, 998.7, 
    999.1, 999.5, 1000, 1000.3, 1001, 1001.2, 1002, 1002.3, 1002.7, 1003, 
    1003.4, 1003.6, 1003.9, 1004.2, 1004.2, 1004.4, 1004.3, 1004.5, 1004.7, 
    1004.6, 1004.8, 1005.1, 1005.4, 1005.4, 1005.5, 1005.6, 1005.9, 1005.8, 
    1005.9, 1006, 1005.9, 1006, 1006.2, 1006.5, 1006.5, 1006.7, 1006.6, 
    1006.6, 1006.5, 1006.4, 1006.3, 1006.2, 1006.1, 1006.1, 1006.2, 1006.3, 
    1006.3, 1006.7, 1006.8, 1007, 1007.3, 1007.5, 1007.8, 1008.1, 1008.4, 
    1008.5, 1008.7, 1008.7, 1008.8, 1009.2, 1009.4, 1009.2, 1009.4, 1009.6, 
    1009.8, 1010.1, 1010, 1010, 1010.5, 1010.4, 1010.7, 1010.8, 1011.1, 
    1011.1, 1011.2, 1011, 1010.9, 1010.8, 1010.8, 1010.7, 1010.7, 1010.8, 
    1010.8, 1011.3, 1011.9, 1012, 1011.9, 1012.5, 1012.9, 1013, 1012.9, 
    1013.4, 1013.6, 1013.8, 1014.2, 1014.8, 1015.2, 1015.3, 1015.6, 1015.7, 
    1016, 1016.2, 1016.6, 1016.9, 1017.5, 1018.1, 1018.5, 1019, 1019.3, 
    1019.4, 1018.9, 1018.9, 1019, 1018.9, 1018.9, 1019.2, 1019.4, 1019.3, 
    1019.4, 1019.7, 1020.2, 1020.4, 1020.1, 1019.8, 1019.5, 1018.9, 1018.5, 
    1018.3, 1018.1, 1017.8, 1017.6, 1017.6, 1017.4, 1017, 1016.6, 1016.2, 
    1015.9, 1015.5, 1015, 1014.8, 1014.5, 1014.3, 1014.1, 1014.1, 1013.9, 
    1013.7, 1013.5, 1013.2, 1012.8, 1012.8, 1012.2, 1012.1, 1012, 1012, 
    1011.8, 1011.8, 1011.9, 1012.2, 1012.2, 1012.5, 1012.5, 1012.5, 1012.5, 
    1012.3, 1012.2, 1011.9, 1011.7, 1011.6, 1011.9, 1011.3, 1010.6, 1009.9, 
    1009.4, 1009.1, 1008.7, 1008.5, 1008.4, 1008.1, 1007.8, 1007.4, 1006.9, 
    1006.4, 1006.2, 1006, 1005.6, 1005.4, 1004.9, 1004.5, 1004.3, 1003.4, 
    1002.9, 1002.4, 1001.9, 1001.3, 1000.6, 1000.2, 999.9, 999.1, 998.9, 
    998.3, 998, 997.5, 997.1, 996.5, 996.4, 996.2, 995.6, 995.2, 994.6, 
    994.3, 994.1, 993.8, 993.4, 993.1, 993.1, 992.9, 992.6, 992.4, 992.4, 
    992.3, 992.3, 992.4, 992.7, 993.1, 993.3, 993.4, 993.5, 993.6, 994, 
    993.8, 994, 993.8, 994.1, 994.1, 994.6, 994.6, 995.2, 995.5, 995.8, 
    995.9, 996.3, 996.2, 996.8, 997.6, 998, 998.2, 998.9, 999.3, 999.3, 
    1000.6, 1000.6, 1001.1, 1001.3, 1001.4, 1001.6, 1001.6, 1001.6, 1001.8, 
    1001.8, 1001.7, 1001.7, 1001.9, 1002, 1002.4, 1002.6, 1002.5, 1002.6, 
    1002.5, 1002.5, 1002.5, 1002.5, 1002.5, 1002.4, 1002.4, 1002.4, 1002.3, 
    1002.5, 1002.5, 1002.4, 1002.3, 1002.2, 1002.1, 1002, 1001.8, 1001.6, 
    1001.5, 1001.5, 1001.5, 1001.4, 1001.2, 1001.1, 1000.8, 1000.8, 1000.7, 
    1000.4, 1000.3, 1000.2, 1000, 999.8, 999.6, 999.3, 999.1, 998.9, 998.7, 
    998.3, 998.3, 998, 998.3, 997.4, 996.9, 996.9, 997.3, 997.4, 997.4, 
    997.5, 997.6, 997.6, 997.6, 997.9, 998.3, 998.8, 999.2, 999.7, 999.9, 
    1000.2, 1000.5, 1000.8, 1001.2, 1001.7, 1002.1, 1002.3, 1002.6, 1002.8, 
    1003, 1003.4, 1003.8, 1004, 1004.5, 1004.9, 1005.3, 1005.5, 1005.5, 
    1005.6, 1005.9, 1006, 1005.6, 1005.4, 1005.2, 1005.2, 1005.3, 1005.4, 
    1005.3, 1004.9, 1004.2, 1003.4, 1002.6, 1001.5, 1000.2, 999.1, 998.5, 
    996.8, 995.7, 994.1, 991.3, 988.8, 985.9, 982.5, 979.5, 975.7, 972.1, 
    969.2, 967.1, 964.9, 962.8, 961, 959.1, 957.9, 957, 956.5, 955.7, 955.3, 
    954.7, 954.4, 954.7, 955.1, 955.6, 956.3, 957.2, 957.8, 958.3, 958.4, 
    958.1, 958.2, 959.1, 960, 960.8, 961.5, 962.2, 962.9, 963.6, 963.7, 
    965.5, 966.2, 966.7, 966.9, 967.3, 967.9, 968.5, 969, 969.8, 970.4, 
    971.1, 971.9, 972.8, 973.5, 974.4, 975.3, 975.9, 976.7, 977.5, 978.2, 
    978.9, 979.5, 980, 980.9, 981.5, 982.4, 983.3, 983.6, 984.3, 985.1, 
    986.1, 986.8, 987.5, 988.1, 988.8, 989.2, 989.5, 989.6, 990.1, 990, 990, 
    989.7, 989.6, 989.6, 989.4, 989.2, 988.9, 988.8, 989, 989.2, 989.5, 
    989.8, 990.2, 990.8, 991.3, 991.7, 992.2, 992.1, 992.3, 992.7, 993.5, 
    994.2, 994.9, 995.7, 996.2, 996.6, 997.5, 998.2, 998.5, 998.9, 999.5, 
    1000.2, 1000.4, 1001.1, 1001.5, 1001.7, 1002.1, 1002.2, 1002.6, 1003.1, 
    1003.1, 1003.2, 1003.5, 1003.5, 1004, 1004, 1004.2, 1004.2, 1004.3, 
    1004.2, 1004.6, 1005, 1005.2, 1005.7, 1005.9, 1006.5, 1006.9, 1007.2, 
    1007.6, 1008.1, 1008.6, 1009.2, 1009.9, 1010.7, 1011.2, 1011.8, 1012.3, 
    1013.2, 1013.7, 1013.9, 1014.3, 1014.6, 1014.8, 1014.7, 1015.1, 1015.5, 
    1016, 1016.4, 1016.6, 1016.8, 1016.9, 1016.5, 1016.9, 1016.8, 1016.8, 
    1017, 1016.9, 1016.8, 1016.6, 1016, 1014.7, 1013.7, 1012.5, 1011.4, 
    1009.8, 1008.5, 1007.4, 1006.4, 1006.2, 1006, 1005.7, 1005.1, 1005, 
    1004.8, 1005.1, 1005.3, 1005, 1004.8, 1005.6, 1006.1, 1006.1, 1006.1, 
    1006.1, 1006, 1005.2, 1005, 1005, 1004.3, 1003.7, 1002.7, 1001.2, 999.3, 
    997.7, 995.8, 993.4, 990.9, 988.4, 985.3, 982.8, 983.8, 985.8, 986.7, 
    986.4, 986.6, 987.5, 987.8, 987.6, 988.2, 988.8, 989, 989.3, 989.8, 
    989.7, 990.3, 991, 991.6, 992.3, 993.1, 994.2, 995.2, 996, 996.6, 997.2, 
    997.9, 998.3, 999, 999.6, 1000, 1000.7, 1001.6, 1002.3, 1003, 1003.7, 
    1004.1, 1004.8, 1005.2, 1005.8, 1006.4, 1006.9, 1007.1, 1007.5, 1008.2, 
    1008.6, 1009, 1009.5, 1009.5, 1009.5, 1009.6, 1009.8, 1009.8, 1009.8, 
    1010, 1010.4, 1010.6, 1010.6, 1010.7, 1010.7, 1010.5, 1010.3, 1010.3, 
    1010.1, 1010.2, 1010, 1009.8, 1009.5, 1009.4, 1009.5, 1009.3, 1009, 
    1008.9, 1008.5, 1008.5, 1008.4, 1008.5, 1008.5, 1008.6, 1008.8, 1008.9, 
    1009.1, 1009.2, 1009.1, 1008.9, 1009, 1009, 1009, 1008.9, 1008.8, 1008.8, 
    1008.6, 1008.4, 1008.5, 1008.3, 1007.9, 1007.7, 1007.7, 1007.5, 1007.1, 
    1006.9, 1006.7, 1006.5, 1006.7, 1006.6, 1006.4, 1006, 1005.7, 1005.4, 
    1005.1, 1004.8, 1005, 1004.7, 1004.7, 1004.8, 1005, 1005, 1005.1, 1005.1, 
    1005.2, 1005.2, 1005, 1005, 1004.8, 1004.6, 1004.7, 1004.9, 1005, 1005.4, 
    1005.7, 1005.7, 1005.9, 1005.9, 1006.1, 1006.1, 1006.2, 1006.3, 1006.4, 
    1006.5, 1006.7, 1006.6, 1006.7, 1006.8, 1006.7, 1006.5, 1006.4, 1006.4, 
    1006.4, 1006.4, 1006.6, 1006.6, 1007, 1007.2, 1007.3, 1007.4, 1007.7, 
    1007.8, 1007.8, 1008, 1008, 1008, 1008.1, 1008.2, 1008.2, 1008.3, 1008.2, 
    1008.3, 1008.3, 1008.2, 1008.2, 1008.1, 1007.9, 1007.8, 1007.8, 1007.7, 
    1007.9, 1008.2, 1008.3, 1008.1, 1008.2, 1008.2, 1007.7, 1008, 1007.9, 
    1007.9, 1008.2, 1008.3, 1008.3, 1008.3, 1008.4, 1008.9, 1008.9, 1008.8, 
    1008.7, 1008.6, 1008.4, 1008.5, 1008.6, 1008.9, 1009.1, 1009.2, 1008.8, 
    1008.8, 1008.3, 1008, 1007.4, 1006.9, 1006.2, 1005.8, 1005.5, 1005.3, 
    1005, 1004.7, 1004.4, 1003.6, 1003.3, 1002.4, 1002.1, 1001.8, 1001.5, 
    1001.3, 1001.3, 1001.5, 1001.7, 1002.7, 1002.8, 1003.3, 1003.2, 1003.1, 
    1002.9, 1003.6, 1003.9, 1004.4, 1004.5, 1004.5, 1004.6, 1004.7, 1004, 
    1003.5, 1003.4, 1003, 1002.4, 1001.8, 1001.2, 1000.9, 1000.6, 999.9, 
    1000, 999.9, 999.5, 998.9, 998.3, 998.2, 998.2, 998.1, 998.1, 998.3, 
    998.1, 998.3, 998.5, 999, 998.7, 998.7, 998.9, 999.5, 999.9, 1000.5, 
    1000.7, 1001, 1001.8, 1002.9, 1003.8, 1004.9, 1005.5, 1006.2, 1007, 
    1007.6, 1008, 1008.3, 1008.9, 1009.5, 1010, 1010.3, 1010.6, 1010.5, 
    1010.7, 1010.9, 1011.4, 1011.4, 1011.5, 1011.6, 1011.7, 1012, 1012, 1012, 
    1012.1, 1012.4, 1012.3, 1012.2, 1012.4, 1012.6, 1012.8, 1012.6, 1012.9, 
    1013.2, 1013.6, 1013.6, 1013.8, 1013.6, 1013.9, 1014, 1013.8, 1014, 
    1014.3, 1014.4, 1014.3, 1014, 1014.1, 1014.2, 1014.3, 1014.5, 1014.7, 
    1014.8, 1014.6, 1014.5, 1014.5, 1014.6, 1014.7, 1014.7, 1014.9, 1015.2, 
    1015.3, 1015.5, 1015.4, 1015.4, 1015.6, 1015.4, 1015.4, 1015.3, 1015.2, 
    1015.3, 1015.3, 1015.5, 1016, 1016.3, 1016.5, 1016.4, 1016.5, 1016.3, 
    1015.9, 1015.7, 1015.2, 1014.9, 1014.3, 1013.7, 1013.4, 1013.1, 1012.6, 
    1012, 1011.5, 1010.8, 1010.3, 1009.4, 1008.9, 1008.4, 1007.9, 1007.3, 
    1006.9, 1007.1, 1007.1, 1007.2, 1007.7, 1008.3, 1008.6, 1009.2, 1009.5, 
    1009.9, 1010.2, 1009.7, 1009.4, 1008.9, 1007.9, 1007.2, 1006, 1004.8, 
    1003.8, 1002.9, 1002, 1000.8, 1000.1, 999.2, 997.8, 996.9, 995.4, 995.1, 
    994.5, 993.1, 992.3, 991.8, 990.9, 990, 989.2, 988.2, 987.4, 987, 987, 
    987.6, 988.5, 989.1, 989.7, 991.3, 991.6, 992.4, 993.1, 993.6, 994.4, 
    994.5, 994.9, 995.3, 995.5, 995.5, 995.3, 994.6, 994.2, 994, 993.8, 
    993.5, 993.6, 993.3, 993.2, 992.6, 992.1, 991.8, 991.7, 991.8, 991.9, 
    991.8, 991.9, 992.3, 992.7, 993.1, 993.5, 993.9, 993.9, 993.8, 994.8, 
    994.9, 995.1, 995.4, 995.8, 996.1, 996.5, 997, 997.4, 997.5, 997.5, 
    997.5, 997.2, 997.2, 997.1, 997.4, 996.2, 996.9, 997.1, 997.3, _, 997.3, 
    997.4, 997.7, 997.8, 998.1, 998.3, 998.5, 997.8, 998.4, 998.9, 999.3, 
    999.5, 1000.1, 1000.6, 1001, 1001.6, 1002.1, 1002.6, 1002.9, 1003.8, 
    1004.5, 1005.3, 1006.2, 1007.2, 1007.8, 1008.3, 1008.7, 1009.4, 1010.1, 
    1010.3, 1010.6, 1010.9, 1011.1, 1011.2, 1011.7, 1012.3, 1012.7, 1012.8, 
    1013.1, 1013.4, 1013, 1012.7, 1012.5, 1012.5, 1012.6, 1012.7, 1012.7, 
    1012.7, 1012.2, 1011.4, 1011.1, 1010.9, 1009.9, 1009.7, 1009.9, 1010.3, 
    1011.2, 1011.9, 1013.1, 1014.1, 1014.7, 1015.2, 1015.6, 1016, 1016.1, 
    1016.2, 1016.4, 1017.3, 1017.5, 1017.6, 1017.7, 1017.9, 1018.1, 1018, 
    1017.9, 1017.9, 1018, 1017.9, 1017.8, 1017.9, 1017.7, 1017.4, 1017.4, 
    1017.5, 1016.9, 1016.5, 1016.2, 1015.9, 1015.3, 1014.8, 1014.5, 1013.6, 
    1012.9, 1012.5, 1012.2, 1011.9, 1011.8, 1011.2, 1010.8, 1010.6, 1010.6, 
    1010.6, 1010.8, 1010.7, 1010.9, 1011.4, 1012, 1012.5, 1012.8, 1013.1, 
    1013.5, 1013.8, 1014.1, 1014.4, 1014.5, 1015.1, 1015.5, 1015.8, 1016.2, 
    1016.4, 1016.4, 1016.3, 1016.3, 1016.3, 1016.3, 1016.3, 1016.3, 1017.4, 
    1017.4, 1017.3, 1017.1, 1017.2, 1017.2, 1016.9, 1016.5, 1016.3, 1015.9, 
    1015.6, 1015.6, 1016, 1016, 1016, 1016.3, 1016.6, 1016.7, 1016.7, 1016.8, 
    1016.9, 1016.6, 1016.4, 1016.6, 1017.2, 1017.2, 1017.2, 1017.2, 1017.3, 
    1017.3, 1017.3, 1017.5, 1017.5, 1017.6, 1017.5, 1017.5, 1017.7, 1018, 
    1018.3, 1018.5, 1018.5, 1018.7, 1018.6, 1018.3, 1017.9, 1017.6, 1017.5, 
    1017.5, 1017.3, 1017.3, 1017.2, 1017, 1016.9, 1016.4, 1016.1, 1015.9, 
    1015.7, 1015.4, 1015, 1014.9, 1014.4, 1014.3, 1014.1, 1013.9, 1013.8, 
    1013.7, 1013.6, 1013.2, 1013.1, 1012.9, 1012.5, 1012.4, 1011.6, 1011.6, 
    1011.8, 1011.7, 1011.5, 1011.5, 1011.3, 1011.2, 1011.2, 1011, 1010.7, 
    1010.5, 1010.6, 1010.5, 1011, 1011.3, 1011.1, 1011.1, 1010.9, 1010.9, 
    1010.7, 1010.9, 1011, 1010.8, 1010.7, 1010.7, 1010.7, 1010.9, 1010.9, 
    1010.8, 1010.8, 1010.8, 1010.6, 1010.3, 1010, 1010.1, 1009, 1009.2, 
    1009.1, 1009.2, 1009, 1008.9, 1009.2, 1009.7, 1009.8, 1010, 1010.4, 
    1010.9, 1010.6, 1010.6, 1010.5, 1010.5, 1011, 1011.4, 1011.8, 1012, 1012, 
    1012, 1012, 1011.8, 1012.5, 1012.5, 1012.7, 1012.7, 1012.9, 1012.7, 
    1012.7, 1012.2, 1011.6, 1011.2, 1010.6, 1010.3, 1009.6, 1009.1, 1008.6, 
    1008.2, 1007.9, 1007.7, 1007.4, 1006.9, 1006.5, 1006.2, 1006, 1005.7, 
    1006.2, 1006.3, 1006.3, 1006.6, 1006.9, 1007.1, 1007.5, 1007.7, 1007.7, 
    1007.8, 1008, 1008.6, 1009.5, 1010.1, 1010.2, 1010.7, 1011.2, 1011.7, 
    1012.2, 1012.4, 1012.6, 1012.8, 1013, 1013.4, 1012.1, 1012.6, 1013.1, 
    1013.5, 1013.7, 1013.9, 1014.2, 1014.6, 1014.6, 1014.6, 1014.7, 1015.1, 
    1015.3, 1015.8, 1016.1, 1016.2, 1016.4, 1016.6, 1016.9, 1017.1, 1017.3, 
    1017.5, 1017.6, 1017.4, 1016.6, 1016.8, 1017, 1017.3, 1017.6, 1018, 
    1018.1, 1018.1, 1017.7, 1017.4, 1017.6, 1018.1, 1017.6, 1017.6, 1017.5, 
    1017.7, 1017.8, 1018, 1018, 1018.2, 1018.5, 1018.5, 1018.3, 1018.2, 
    1017.8, 1018.3, 1018.8, 1019.4, 1019.8, 1019.7, 1019.8, 1020.4, 1021, 
    1021.2, 1021, 1020.9, 1021.7, 1022.2, 1022.7, 1023.4, 1023.9, 1024.2, 
    1024.2, 1024.5, 1025.1, 1025.5, 1025.6, 1025.7, 1025.9, 1026.1, 1026.5, 
    1026.8, 1027.3, 1027.3, 1027.1, 1026.9, 1026.8, 1026.6, 1026.5, 1026.3, 
    1025.8, 1025.6, 1025.5, 1025.5, 1025.1, 1024.8, 1024.4, 1023.9, 1023.2, 
    1022.8, 1022.6, 1022.1, 1021.1, 1021, 1020.7, 1020.3, 1020, 1019.6, 
    1019.2, 1018.9, 1018.5, 1017.6, 1017.1, 1016.5, 1016.4, 1016.2, 1015.9, 
    1015.7, 1015.6, 1015.4, 1015.2, 1014.9, 1014.3, 1014.1, 1014.1, 1014.1, 
    1013.3, 1013.5, 1013.6, 1013.8, 1013.8, 1013.7, 1013.5, 1013.2, 1012.8, 
    1012.7, 1012.2, 1011.7, 1010.9, 1010.5, 1010.2, 1009.4, 1008.5, 1008.2, 
    1007.5, 1006.8, 1006.1, 1005.4, 1004.4, 1003.5, 1001.8, 1000.4, 999.3, 
    999, 998.7, 998.3, 997.8, 997.2, 996.7, 996.6, 996.5, 996.1, 994.4, 
    992.5, 991, 989.3, 987.3, 983.6, 979.6, 976.4, 973.5, 972.5, 973.2, 
    973.4, 973, 973.5, 974.4, 975.3, 976.5, 978.1, 979.8, 981.1, 982.3, 
    983.5, 984.2, 985, 985.9, 986.8, 987.5, 988, 988.6, 989.4, 990.2, 991.3, 
    992.9, 994.6, 996.4, 997.9, 1000.4, 1002.3, 1004.1, 1005.6, 1006.4, 
    1006.8, 1007, 1007.1, 1007, 1006.8, 1007.7, 1009, 1010.8, 1011.4, 1011.6, 
    1011.8, 1012.1, 1011.9, 1011.5, 1010.6, 1009.2, 1007.6, 1006.2, 1005.1, 
    1002.5, 1001.1, 999.3, 997.3, 995.1, 993.3, 992.1, 990.9, 990, 989.1, 
    988.5, 987.8, 988.2, 987.7, 987.3, 986.9, 986.6, 986.3, 986.1, 985.5, 
    985.1, 984.8, 984.9, 985, 985.7, 985.8, 986.2, 986.7, 987.1, 987.8, 
    988.3, 988.8, 989.5, 990, 990.2, 990.5, 991.4, 991.8, 992.1, 992.4, 
    992.5, 992.4, 992.5, 992.5, 992.4, 991.9, 991.5, 991.2, 992.9, 993.2, 
    993.9, 994.3, 994.8, 995.3, 996.1, 996.7, 997.1, 997.1, 997.1, 997.6, 
    997.8, 997.7, 997.5, 997, 996.3, 995.3, 995.4, 995.2, 995.3, 995.2, 
    994.8, 994.6, 994.6, 994.7, 994.2, 993.5, 993, 992.1, 990.7, 988.8, 
    987.4, 986.4, 985.3, 984.7, 984.4, 985, 986.3, 987.8, 989, 990.5, 991.9, 
    992.5, 992.5, 992.6, 992.5, 993, 991.5, 990.3, 991.7, 994.4, 996.8, 998, 
    999.3, 1000.2, 1001.3, 1002.4, 1003.6, 1004.5, 1004.9, 1005.5, 1006.1, 
    1006.6, 1006.9, 1007.2, 1007.6, 1007.9, 1008.2, 1008.7, 1009.1, 1009.4, 
    1009.2, 1009.5, 1009.9, 1010.5, 1010.9, 1011.1, 1011.2, 1011.3, 1011.5, 
    1011.7, 1011.8, 1012, 1012.8, 1013, 1013.4, 1013.6, 1013.7, 1013.9, 
    1014.2, 1014.3, 1014.4, 1014.2, 1014.1, 1014.1, 1013.9, 1013.9, 1014.2, 
    1014.4, 1014.5, 1014.6, 1014.4, 1014.1, 1013.7, 1013.4, 1013.4, 1013.5, 
    1013.4, 1013.5, 1013.5, 1013.4, 1013.3, 1013.3, 1013.3, 1013.4, 1013.6, 
    1013.6, 1013.5, 1013.2, 1013.4, 1013.6, 1014, 1014.3, 1014.6, 1014.8, 
    1014.9, 1015, 1015, 1015, 1015, 1015.2, 1015.7, 1015.7, 1015.6, 1015.4, 
    1015.5, 1015.8, 1015.9, 1016, 1016.1, 1016, 1015.9, 1016, 1016.9, 1017.1, 
    1017.5, 1017.5, 1017.7, 1017.9, 1018, 1018.2, 1018.3, 1018.7, 1018.7, 
    1018.8, 1018.8, 1019.2, 1019.5, 1019.7, 1019.9, 1020.1, 1020.4, 1020.8, 
    1020.8, 1020.6, 1020.5, 1020.6, 1021.7, 1022, 1022.2, 1022.6, 1023, 
    1023.4, 1023.8, 1023.9, 1023.8, 1023.9, 1023.9, 1024.3, 1024.8, 1025, 
    1025.2, 1025.6, 1025.7, 1025.8, 1026, 1026.3, 1026.5, 1026.6, 1026.6, 
    1026.8, 1026.5, 1026.7, 1027, 1027.4, 1027.8, 1028.2, 1028.4, 1028.8, 
    1029.3, 1029.7, 1030.1, 1030.3, 1030.1, 1030.5, 1030.9, 1031.1, 1031.4, 
    1031.6, 1031.6, 1031.8, 1032.1, 1032.1, 1032.1, 1032, 1031.7, 1031.9, 
    1032, 1032.3, 1032.5, 1032.6, 1032.7, 1032.8, 1032.8, 1032.8, 1032.7, 
    1032.7, 1032.3, 1032.2, 1032.1, 1032.2, 1032.2, 1032.1, 1032, 1032, 
    1032.1, 1032, 1031.8, 1031.5, 1032.1, 1032.1, 1032.2, 1032.4, 1032.7, 
    1032.6, 1032.5, 1032.5, 1032.4, 1032.2, 1031.9, 1031.6, 1031.5, 1031.1, 
    1030.8, 1030.6, 1030.4, 1030.1, 1030.1, 1030.1, 1030.1, 1029.9, 1029.6, 
    1029.4, 1030, 1029.9, 1029.9, 1029.9, 1030, 1030.2, 1030.3, 1030.3, 
    1030.5, 1030.6, 1030.7, 1030.9, 1031.7, 1032.2, 1032.3, 1032.1, 1032, 
    1032.2, 1032.6, 1032.9, 1032.6, 1032.3, 1032.2, 1032.3, 1032.2, 1032.1, 
    1032.1, 1032.6, 1032.9, 1033, 1033, 1033.1, 1033, 1033, 1033, 1033.2, 
    1032.9, 1033.3, 1033.6, 1033.9, 1034.1, 1034.2, 1034.6, 1034.7, 1034.7, 
    1034.6, 1034.5, 1034.3, 1034.5, 1034.7, 1035, 1035, 1035.1, 1035.1, 
    1035.1, 1035.3, 1035.3, 1035.5, 1035.4, 1035.6, 1036.7, 1036.9, 1037.2, 
    1037.2, 1036.9, 1037, 1036.9, 1036.6, 1036.5, 1036.1, 1035.6, 1035.1, 
    1034.3, 1034, 1033.8, 1034, 1033.8, 1033.7, 1033.6, 1033.5, 1033.2, 
    1032.9, 1032.7, 1032.5, 1032.7, 1032.5, 1032.4, 1032.6, 1032.8, 1033.4, 
    1034, 1034.7, 1035.5, 1036.1, 1037.1, 1038, 1038.6, 1039.6, 1040.5, 
    1041.2, 1042, 1041.5, 1042.3, 1042.9, 1043, 1043.1, 1043.1, 1043.5, 
    1043.7, 1044, 1044.5, 1044.7, 1044.9, 1044.9, 1044.7, 1043.9, 1043.8, 
    1043.5, 1043, 1042.4, 1042.2, 1041.9, 1041.4, 1040.8, 1040, 1039.3, 1039, 
    1038.7, 1037.8, 1037.3, 1037.2, 1037.2, 1037.7, 1036.7, 1036.1, 1035.9, 
    1035.9, 1035.9, 1036, 1036.5, 1037, 1037.3, 1037.2, 1037.1, 1038.4, 
    1038.8, 1038.6, 1038.7, 1038.6, 1037.7, 1036.7, 1035.8, 1034.4, 1033.7, 
    1032.7, 1032.3, 1032, 1032.2, 1031.6, 1030.7, 1030, 1029.7, 1028.9, 
    1027.7, 1026.6, 1025.6, 1024.5, 1023.7, 1022.3, 1021.2, 1020.4, 1019.6, 
    1018.4, 1016.9, 1015.5, 1013.9, 1012.8, 1012.2, 1011.6, 1011.3, 1014.4, 
    1015, 1015.9, 1016.8, 1017.6, 1019.2, 1021, 1022.6, 1024, 1025, 1026, 
    1027.5, 1027.5, 1028.5, 1029.6, 1030.6, 1030.4, 1031.3, 1032.1, 1032.6, 
    1033.4, 1033.7, 1034.2, 1034.7, 1035.1, 1035.5, 1035.8, 1036.1, 1036.4, 
    1036.8, 1036.7, 1036.4, 1036.2, 1036.1, 1036.2, 1036.1, 1036.1, 1036.2, 
    1036.1, 1036.1, 1036.3, 1036.3, 1036.2, 1036.1, 1035.8, 1035.8, 1036, 
    1035.8, 1035.7, 1035.2, 1035.4, 1035.3, 1035.1, 1035.1, 1034.8, 1034.6, 
    1034.5, 1034.1, 1033.5, 1032.9, 1032.5, 1032.2, 1031.9, 1031.8, 1031.8, 
    1031.7, 1031.6, 1031.3, 1030.9, 1030.6, 1030.2, 1030.2, 1029.7, 1029.3, 
    1029.2, 1029, 1029, 1028.9, 1028.8, 1028.8, 1029, 1028.9, 1028.8, 1028.8, 
    1029.1, 1028.8, 1029, 1029.4, 1029.5, 1029.6, 1029.9, 1029.9, 1030, 
    1030.3, 1030.3, 1030.2, 1030.3, 1030.1, 1030.4, 1030.6, 1030.9, 1031.1, 
    1031.1, 1031.2, 1031.4, 1031.4, 1031.5, 1031.7, 1031.7, 1031.9, 1032.2, 
    1032.4, 1032.8, 1033, 1033, 1033, 1032.9, 1033, 1032.9, 1032.9, 1032.9, 
    1032.7, 1032.9, 1033, 1033.1, 1032.9, 1032.7, 1032.4, 1032.3, 1032.1, 
    1031.9, 1031.8, 1031.8, 1031.9, 1031.9, 1031.9, 1031.8, 1031.8, 1031.6, 
    1031.6, 1031.4, 1031.3, 1031.4, 1031.4, 1031.5, 1031.1, 1031, 1030.9, 
    1030.8, 1030.6, 1030.4, 1030.3, 1030.2, 1030.1, 1030, 1029.8, 1029.5, 
    1029.4, 1029.4, 1029.6, 1029.5, 1029.6, 1029.5, 1029.3, 1029.2, 1029.1, 
    1029, 1028.9, 1028.6, 1028.7, 1028.5, 1028.5, 1028.4, 1028.3, 1028.3, 
    1028, 1027.9, 1028, 1027.8, 1027.7, 1027.8, 1027.8, 1028, 1028.3, 1028.3, 
    1028.3, 1028.3, 1028.3, 1028.3, 1028.4, 1028.3, 1028.2, 1028.2, 1028.3, 
    1028.4, 1028.5, 1028.6, 1028.5, 1028.5, 1028.3, 1028.4, 1028.4, 1028.4, 
    1028.4, 1028.6, 1028.7, 1028.8, 1029.2, 1029.3, 1029.3, 1029.3, 1029.4, 
    1029.4, 1029.6, 1029.6, 1029.6, 1029.6, 1029.7, 1029.9, 1030.1, 1030.3, 
    1030.3, 1030.4, 1030.4, 1030.4, 1030.5, 1030.5, 1030.4, 1030.5, 1030.7, 
    1031, 1031.2, 1031.2, 1031.2, 1031.4, 1031.5, 1031.5, 1031.5, 1031.4, 
    1031.5, 1031.6, 1032, 1032, 1031.9, 1031.9, 1031.9, 1031.7, 1031.6, 
    1031.6, 1031.5, 1031.4, 1031.5, 1031.5, 1031.6, 1031.5, 1031.7, 1031.8, 
    1031.7, 1031.5, 1031.5, 1031.3, 1031.3, 1031.3, 1031.1, 1030.9, 1030.9, 
    1031, 1030.9, 1030.7, 1030.4, 1030.2, 1029.8, 1029.6, 1029.4, 1029.1, 
    1028.8, 1028.3, 1028.1, 1028, 1028.1, 1027.7, 1027.4, 1027, 1026.7, 
    1026.4, 1026.3, 1026, 1025.8, 1025.9, 1026, 1026, 1026.1, 1025.8, 1025.5, 
    1025.3, 1024.9, 1024.7, 1024.5, 1024.5, 1024.4, 1024.4, 1024.3, 1024.5, 
    1024.6, 1024.6, 1024.5, 1024.6, 1024.6, 1024.5, 1024.5, 1024.5, 1024.6, 
    1024.7, 1024.7, 1024.7, 1025.1, 1025.2, 1025.2, 1025.2, 1025, 1025.1, 
    1025.1, 1025.2, 1025.1, 1025.2, 1025.4, 1025.5, 1025.6, 1025.7, 1025.6, 
    1025.7, 1025.8, 1025.6, 1025.7, 1025.8, 1025.8, 1025.8, 1025.9, 1025.8, 
    1025.8, 1026, 1025.8, 1025.7, 1025.8, 1025.9, 1025.6, 1025.5, 1025.7, 
    1025.7, 1025.8, 1026.1, 1026.5, 1026.4, 1026.7, 1026.7, 1026.8, 1027, 
    1027.1, 1027.1, 1027.2, 1027.3, 1027.2, 1027.4, 1027.4, 1027.5, 1027.4, 
    1027.5, 1027.4, 1027.2, 1027.2, 1027.1, 1027, 1027.2, 1027.2, 1027, 
    1026.7, 1026.7, 1026.6, 1026.2, 1026.4, 1026, 1025.6, 1025.2, 1024.8, 
    1024, 1023.7, 1023.6, 1023.2, 1022.9, 1022.5, 1022, 1021.3, 1020.7, 
    1020.4, 1019.8, 1019.4, 1019, 1018.6, 1018.2, 1017.9, 1017.9, 1017.6, 
    1016.7, 1016.3, 1015.8, 1015.1, 1014.2, 1013, 1012.2, 1011.3, 1010.3, 
    1009.3, 1007.9, 1006.5, 1004.9, 1003, 1001.3, 999.3, 997.2, 995.3, 993.3, 
    991.5, 989.8, 988.2, 986.7, 984.9, 983.9, 982.6, 981.9, 981.5, 981.2, 
    981.1, 980.7, 981.4, 982.3, 983.3, 984.5, 986, 987.2, 988.6, 990.7, 
    993.5, 995.6, 996.9, 999.4, 1001.7, 1003.1, 1005, 1006.7, 1008.2, 1009.4, 
    1010.8, 1012.1, 1013.6, 1015, 1016, 1016.6, 1016.9, 1017.8, 1018.6, 1019, 
    1019.2, 1019.7, 1019.9, 1020.1, 1020.4, 1020.7, 1021.1, 1021.2, 1021.8, 
    1022, 1022.2, 1022.4, 1022.2, 1022.4, 1022.3, 1022.3, 1022, 1021.8, 
    1021.3, 1020.9, 1020.6, 1020.5, 1020.2, 1019.7, 1019.2, 1018.7, 1017.8, 
    1017.2, 1016.9, 1016.5, 1016, 1015.8, 1015.4, 1015, 1014.5, 1014.1, 
    1013.5, 1013, 1012.9, 1012.5, 1012.2, 1011.7, 1011.2, 1011.1, 1010.7, 
    1010.5, 1010.3, 1009.8, 1009.2, 1008.9, 1008.7, 1008.4, 1008, 1007.6, 
    1007.6, 1007.6, 1007.2, 1007.3, 1007.4, 1007.6, 1007.6, 1007.6, 1007.9, 
    1008.4, 1008.7, 1009.1, 1009.1, 1009.4, 1009.5, 1009.8, 1010.1, 1010.5, 
    1010.5, 1010.5, 1010.5, 1010.4, 1010.1, 1010, 1009.8, 1009.6, 1009.1, 
    1008.8, 1008.3, 1008, 1007.6, 1007.3, 1007.2, 1007, 1007, 1006.5, 1006.5, 
    1006.3, 1006.5, 1006.5, 1006.6, 1006.7, 1006.9, 1006.9, 1006.9, 1007.1, 
    1007.2, 1007.3, 1007.6, 1007.4, 1007.3, 1007.1, 1007.3, 1007.4, 1007.4, 
    1007.4, 1007.8, 1008, 1008.3, 1008.9, 1009.6, 1010.3, 1010.8, 1011.1, 
    1011.5, 1011.8, 1012, 1012.3, 1012.2, 1012.5, 1012.4, 1012.9, 1013.9, 
    1014.3, 1014.5, 1014.9, 1015.4, 1015.7, 1015.8, 1016, 1016.1, 1015.9, 
    1016.2, 1016.6, 1016.8, 1017.5, 1017.9, 1018.4, 1018.7, 1018.8, 1018.8, 
    1018.9, 1019, 1019, 1019.1, 1019, 1019, 1019, 1019, 1019.1, 1019.6, 
    1019.8, 1020, 1020.1, 1020.4, 1020.4, 1020.2, 1020.1, 1019.8, 1019.7, 
    1019.1, 1018.6, 1018.3, 1017.6, 1017.1, 1016.8, 1015.7, 1015.5, 1015.5, 
    1015.1, 1014.8, 1014.5, 1014.3, 1014.2, 1014.2, 1014.5, 1014.3, 1014.2, 
    1014, 1013.9, 1013.7, 1013.6, 1013.4, 1013.5, 1013.1, 1013.1, 1013.3, 
    1013.2, 1013.2, 1013, 1012.8, 1012.6, 1012.4, 1012.4, 1012.2, 1011.9, 
    1012, 1011.9, 1011.8, 1011.7, 1012, 1011.7, 1012, 1011.8, 1011.4, 1010.9, 
    1010.3, 1009.9, 1009.8, 1009.3, 1008.6, 1008, 1007.5, 1006.8, 1006.1, 
    1005.7, 1005.2, 1005, 1004.8, 1004.8, 1004.7, 1004.9, 1005.3, 1005.7, 
    1006.1, 1006.5, 1006.9, 1007.3, 1007.6, 1008, 1008.3, 1008.6, 1009.1, 
    1009.5, 1009.9, 1010.1, 1010.4, 1010.7, 1011, 1011.1, 1011.3, 1011.5, 
    1011.7, 1011.8, 1012.1, 1012.3, 1012.6, 1012.9, 1013.2, 1013.3, 1013.2, 
    1013.1, 1013, 1013.2, 1012.9, 1013, 1012.9, 1013, 1013, 1013.1, 1013, 
    1013, 1012.7, 1012.7, 1012.4, 1012.3, 1012.1, 1012, 1012, 1011.8, 1011.8, 
    1011.8, 1011.8, 1011.7, 1011.6, 1011.2, 1011.1, 1011, 1010.9, 1010.9, 
    1010.9, 1011.1, 1011.2, 1011.3, 1011.4, 1011.4, 1011.5, 1011.5, 1011.4, 
    1011.6, 1011.7, 1011.7, 1012, 1012.2, 1012.5, 1012.7, 1013, 1013.2, 
    1013.4, 1013.6, 1013.7, 1013.6, 1013.9, 1014.2, 1014.4, 1014.8, 1015.1, 
    1015.6, 1016, 1016.4, 1016.6, 1016.8, 1017.2, 1017.5, 1017.8, 1018.4, 
    1019.2, 1020.1, 1020.6, 1021.2, 1021.9, 1022.2, 1022.7, 1023.2, 1023.5, 
    1023.8, 1024.2, 1024.5, 1024.9, 1025.1, 1025.5, 1026, 1026.4, 1026.5, 
    1026.7, 1026.8, 1027, 1027.4, 1027.5, 1027.9, 1028.4, 1028.6, 1028.6, 
    1029, 1029.1, 1029.3, 1029.3, 1029.2, 1029.3, 1029.2, 1029.3, 1029.5, 
    1029.8, 1029.9, 1030, 1029.9, 1030.2, 1030, 1029.8, 1029.5, 1029.4, 
    1029.5, 1029.2, 1029.3, 1029.2, 1029, 1028.8, 1028.9, 1028.7, 1028.4, 
    1028.3, 1028.1, 1027.8, 1027.9, 1027.4, 1027.1, 1027.1, 1027, 1027, 
    1026.9, 1026.8, 1026.8, 1026.8, 1026.5, 1026.4, 1026, 1026.1, 1025.9, 
    1025.7, 1025.7, 1025.4, 1025.2, 1025.2, 1024.9, 1024.5, 1024.3, 1024.1, 
    1023.9, 1023.7, 1023.4, 1023.2, 1023.3, 1023.2, 1022.9, 1022.6, 1022.5, 
    1022.1, 1021.7, 1021.3, 1020.9, 1020.7, 1020.6, 1020.3, 1020, 1019.8, 
    1019.6, 1019.4, 1019.2, 1018.8, 1018.5, 1018.2, 1017.9, 1017.9, 1017.9, 
    1017.9, 1017.7, 1017.7, 1017.5, 1017.3, 1017.5, 1017.6, 1017.4, 1017.5, 
    1017.4, 1017.5, 1017.6, 1017.5, 1017.8, 1018.1, 1018.1, 1018.2, 1018.3, 
    1018.2, 1018.1, 1018.2, 1018.2, 1018.3, 1018.5, 1018.7, 1018.8, 1018.8, 
    1018.9, 1019.1, 1019.1, 1019.2, 1019.3, 1019.3, 1019.3, 1019.2, 1019.4, 
    1019.4, 1019.2, 1019.3, 1019.2, 1019.3, 1019.4, 1019.4, 1019.3, 1019.2, 
    1019.2, 1019, 1018.9, 1018.8, 1018.8, 1018.7, 1018.6, 1018.4, 1018.4, 
    1018.5, 1018.3, 1018.2, 1018.1, 1018, 1018, 1017.9, 1017.9, 1017.5, 
    1017.4, 1017.1, 1017.1, 1016.9, 1016.9, 1016.7, 1016.5, 1016.2, 1015.9, 
    1015.7, 1015.2, 1015, 1014.7, 1014.4, 1013.9, 1013.5, 1013, 1012.2, 
    1011.5, 1010.7, 1009.9, 1009.4, 1008.6, 1007.4, 1006.1, 1005, 1003.9, 
    1003, 1002.1, 1001.6, 1000.3, 1001.1, 1001.1, 1001.8, 1001.7, 1002.3, 
    1002.8, 1003.2, 1003.6, 1004.4, 1004.9, 1005.8, 1006.4, 1007, 1007.7, 
    1008.6, 1009.4, 1009.7, 1010.2, 1010.8, 1011.2, 1011.6, 1011.9, 1011.9, 
    1012, 1011.9, 1011.7, 1011.6, 1011.6, 1011.7, 1011.1, 1010.6, 1010.8, 
    1010.4, 1010.1, 1009.3, 1009, 1008.8, 1008.3, 1008.2, 1007.7, 1007.2, 
    1006.4, 1005.8, 1004.8, 1004.3, 1004.3, 1004.2, 1004.3, 1004.5, 1005, 
    1005.4, 1006.6, 1007.2, 1008, 1008.3, 1008.8, 1009.1, 1009.2, 1009.8, 
    1010.1, 1009.7, 1010, 1009.9, 1009.4, 1009.6, 1009.1, 1008.4, 1007.4, 
    1006, 1005, 1004.1, 1003.5, 1002.8, 1002.2, 1002, 1001.9, 1002.1, 1002.2, 
    1002.6, 1003, 1003.4, 1003.8, 1004.2, 1004.4, 1004.7, 1005.3, 1005.9, 
    1006.5, 1007.3, 1008.2, 1008.8, 1009.5, 1010.3, 1011.2, 1012, 1012.7, 
    1013.2, 1013.5, 1014, 1014.6, 1015, 1015.4, 1016.1, 1016.6, 1016.7, 
    1017.1, 1017.3, 1017.5, 1017.7, 1018, 1018, 1018.1, 1018.5, 1018.6, 
    1018.6, 1018.4, 1018.2, 1018, 1017.5, 1016.9, 1016.2, 1015.7, 1015.5, 
    1015.8, 1016.4, 1016.8, 1017.1, 1017.8, 1018.1, 1018.5, 1018.7, 1018.9, 
    1018.9, 1018.8, 1018.9, 1019, 1019.1, 1019.2, 1019, 1018.6, 1018.5, 
    1018.3, 1017.8, 1017.3, 1016.7, 1016.1, 1015.6, 1015.6, 1015.2, 1014.7, 
    1014.3, 1013.6, 1013.4, 1013, 1012.8, 1012.5, 1012.4, 1012.2, 1012.1, 
    1012.3, 1012.4, 1012.6, 1012.5, 1012.4, 1012.3, 1012.2, 1012.1, 1011.9, 
    1011.5, 1011.2, 1011.1, 1010.9, 1010.9, 1010.6, 1010.5, 1010.4, 1010.2, 
    1010.3, 1010.4, 1010.7, 1010.7, 1011.4, 1012.2, 1013, 1013.6, 1014.3, 
    1014.9, 1015.5, 1016.1, 1016.7, 1017.3, 1017.7, 1018.3, 1018.6, 1019.3, 
    1020, 1020.6, 1021.2, 1021.5, 1021.5, 1021.5, 1022.2, 1022.6, 1022.9, 
    1023.1, 1023, 1022.9, 1023.4, 1023.7, 1024.3, 1024.4, 1024.9, 1025.3, 
    1025.4, 1025.3, 1025.6, 1025.9, 1026, 1026.3, 1026.5, 1026.9, 1027.5, 
    1027.8, 1028.1, 1028.1, 1028.3, 1028.4, 1028.6, 1028.8, 1029, 1028.8, 
    1028.9, 1028.9, 1028.9, 1028.9, 1028.8, 1028.6, 1028.4, 1028.2, 1027.8, 
    1027.2, 1026.6, 1026.1, 1025.7, 1025.1, 1024.8, 1024.3, 1023.8, 1023.2, 
    1022.7, 1021.9, 1021.4, 1020.7, 1020.3, 1019.7, 1019.1, 1018.5, 1018.1, 
    1017.8, 1017.4, 1016.8, 1016.4, 1015.6, 1014.9, 1014.2, 1013.7, 1013.1, 
    1012.7, 1012.3, 1011.9, 1011.7, 1011.3, 1010.8, 1010.4, 1010, 1009.5, 
    1009, 1008.4, 1007.9, 1007.5, 1007.1, 1006.8, 1006.5, 1006, 1005.2, 
    1005.1, 1005, 1005.2, 1005.4, 1005.7, 1006, 1005.9, 1006, 1006.3, 1006.6, 
    1006.7, 1007.2, 1007.5, 1007.8, 1008.2, 1008.7, 1008.9, 1009.2, 1009.4, 
    1009.6, 1009.9, 1010.1, 1010.3, 1010.3, 1010.5, 1010.3, 1010.6, 1010.5, 
    1010.8, 1010.9, 1011.1, 1011.1, 1011.3, 1011.2, 1011.2, 1011.2, 1010.7, 
    1010.5, 1010.1, 1009.8, 1009.5, 1009, 1008.6, 1008.3, 1008, 1007.6, 
    1007.4, 1007.2, 1007, 1006.5, 1006.3, 1006.4, 1006.5, 1006.7, 1007, 
    1006.9, 1007, 1007.2, 1007.4, 1007.6, 1007.5, 1007.6, 1007.5, 1007.5, 
    1007.5, 1007.4, 1007.7, 1007.6, 1007.7, 1007.7, 1007.6, 1007.4, 1007.1, 
    1006.9, 1006.8, 1006.8, 1006.9, 1006.8, 1006.8, 1006.8, 1006.8, 1006.8, 
    1006.8, 1006.7, 1006.6, 1006.5, 1006.4, 1006.3, 1006.2, 1006.5, 1006.5, 
    1006.6, 1006.6, 1006.8, 1006.9, 1007, 1007.1, 1007.2, 1007.2, 1007.3, 
    1007.5, 1007.6, 1007.8, 1007.9, 1008.2, 1008.4, 1008.5, 1008.8, 1008.9, 
    1009, 1009.2, 1009.3, 1009.6, 1009.9, 1010.1, 1010.4, 1010.6, 1010.8, 
    1011.1, 1011.4, 1011.5, 1011.7, 1011.9, 1012.2, 1012.4, 1012.6, 1013, 
    1013.3, 1013.5, 1013.5, 1013.7, 1014, 1014.1, 1014.2, 1014.2, 1014.3, 
    1014.5, 1014.7, 1014.9, 1015.1, 1015.5, 1015.5, 1015.7, 1015.8, 1015.8, 
    1015.8, 1016, 1016.1, 1016.2, 1016.5, 1016.5, 1016.4, 1016.3, 1016.2, 
    1016.1, 1015.9, 1015.8, 1015.7, 1015.5, 1015.3, 1015, 1014.9, 1014.8, 
    1014.7, 1014.3, 1013.8, 1013.4, 1013, 1012.9, 1012.5, 1012.2, 1012, 
    1011.8, 1011.7, 1011.6, 1011.5, 1011.1, 1010.8, 1010.6, 1010.5, 1010.5, 
    1010.4, 1010.2, 1010.2, 1010.3, 1010.5, 1010.7, 1010.9, 1011, 1011, 
    1011.2, 1011.5, 1011.7, 1011.7, 1011.7, 1011.9, 1012, 1011.9, 1012.1, 
    1012.5, 1012.5, 1012.6, 1012.8, 1012.9, 1012.9, 1012.9, 1012.9, 1013.1, 
    1013.3, 1013.5, 1013.7, 1013.8, 1014, 1014.2, 1014.5, 1014.6, 1014.8, 
    1014.6, 1014.8, 1015, 1015.1, 1015.1, 1015.4, 1015.6, 1015.8, 1015.9, 
    1016.1, 1016.2, 1016.4, 1016.8, 1016.9, 1016.9, 1017.2, 1017.5, 1017.5, 
    1017.8, 1017.9, 1018.1, 1018.5, 1018.7, 1019, 1019.1, 1019, 1018.9, 1019, 
    1019.3, 1019.4, 1019.6, 1019.8, 1019.9, 1019.9, 1020.1, 1020.2, 1020.2, 
    1020.2, 1020.3, 1020.3, 1020.5, 1020.7, 1021, 1021.3, 1021.5, 1021.4, 
    1021.4, 1021.5, 1021, 1020.7, 1020.3, 1020, 1020, 1020, 1019.9, 1019.6, 
    1020.1, 1019.9, 1019.9, 1019.8, 1019.7, 1019.5, 1019.1, 1018.9, 1018.9, 
    1018.7, 1018.4, 1018.1, 1017.7, 1017.7, 1017.4, 1017, 1016.6, 1016.4, 
    1016.1, 1015.9, 1015.7, 1014.9, 1014.3, 1013.8, 1013.6, 1013.3, 1012.9, 
    1012.6, 1011.9, 1011.2, 1011, 1010.4, 1010.1, 1009.8, 1009.8, 1009.3, 
    1009.1, 1009.3, 1009.3, 1009.7, 1009.7, 1009.8, 1009.8, 1009.9, 1010, 
    1010.1, 1010.1, 1009.8, 1009.4, 1009.1, 1008.9, 1008.6, 1007.8, 1007.2, 
    1006.6, 1006.1, 1005.1, 1004.4, 1004.2, 1003.4, 1002.5, 1002, 1001.1, 
    1000, 998.9, 998, 997.2, 997.1, 998.4, 999.1, 999.5, 999.8, 1000.1, 
    1000.3, 1000.5, 1000.6, 1000.4, 1000.3, 999.9, 999.5, 998.6, 998, 997.3, 
    996.7, 996, 994.3, 992.7, 991.6, 991.2, 991, 981, 991.3, 992.2, 993, 
    993.8, 994.6, 995.4, 996, 996.7, 997.4, 998, 998.8, 999.5, 1000.1, 
    1000.8, 1001.3, 1002.2, 1002.7, 1003.2, 1003.5, 1004.1, 1004.1, 1004.2, 
    1004.3, 1004.3, 1004, 1003.7, 1003.6, 1003.7, 1003.9, 1004.2, 1004.2, 
    1004, 1004.2, 1003.9, 1003.4, 1002.9, 1002.6, 1002.4, 1002.3, 1002.2, 
    1002.4, 1002.4, 1002.5, 1002.6, 1003.1, 1003.2, 1003.8, 1004.6, 1005.2, 
    1005.9, 1006.4, 1006.9, 1007.4, 1008, 1008.5, 1009, 1009.1, 1009.3, 1009, 
    1008.9, 1009, 1008.4, 1007.8, 1006.9, 1006, 1005.1, 1004.2, 1003, 1001.8, 
    1000.3, 998.7, 996.9, 995.4, 994.3, 993.2, 992.9, 992.8, 992.8, 993.2, 
    994.1, 995, 996.3, 997.4, 998.7, 999.8, 1001.1, 1002.3, 1003.4, 1004.5, 
    1005.5, 1006.6, 1007.5, 1008.5, 1009.2, 1009.9, 1010.8, 1011.6, 1012, 
    1012.6, 1013, 1013.6, 1013.9, 1014.2, 1014.1, 1014.1, 1014, 1014.2, 
    1014.2, 1014.1, 1013.9, 1014, 1013.9, 1013.5, 1013.3, 1013, 1012.5, 
    1011.7, 1010.6, 1009.6, 1008.2, 1007.2, 1006.6, 1006, 1005.5, 1005.2, 
    1005, 1005.1, 1005.4, 1005.7, 1006, 1006.2, 1006.6, 1007.2, 1007.8, 
    1008.6, 1009.4, 1010.3, 1011, 1011.9, 1012.5, 1013.2, 1013.9, 1014.4, 
    1015.1, 1015.8, 1016.4, 1017.1, 1017.8, 1018.3, 1018.6, 1019, 1019.4, 
    1019.3, 1019.1, 1018.9, 1018.4, 1017.9, 1017.2, 1016.4, 1016, 1015.4, 
    1015, 1014.5, 1014.2, 1014.2, 1014.2, 1013.8, 1014.9, 1015.6, 1016.8, 
    1017.9, 1018.8, 1020, 1020.3, 1021.7, 1022.5, 1023.5, 1024.2, 1024.7, 
    1025, 1025.2, 1025.7, 1026.2, 1026.8, 1026.8, 1026.7, 1026.9, 1027.3, 
    1027.3, 1027.2, 1026.8, 1026.2, 1025.8, 1025.3, 1024.8, 1024.3, 1023.9, 
    1023.4, 1022.9, 1022.4, 1021.8, 1021.1, 1020.4, 1019.5, 1019.1, 1018.7, 
    1018.4, 1017.9, 1017.6, 1017.4, 1017, 1016.5, 1016.3, 1015.8, 1015.2, 
    1014.9, 1014.5, 1014.3, 1014.3, 1013.8, 1014, 1013.8, 1013.5, 1012.9, 
    1012.5, 1012.5, 1011.9, 1011.2, 1010.8, 1011, 1011.2, 1011.2, 1011.2, 
    1011.2, 1011, 1011.1, 1010.9, 1010.7, 1010.7, 1010.3, 1010, 1009.8, 
    1009.5, 1008.9, 1008.4, 1007.6, 1006.7, 1005.8, 1005.3, 1004.4, 1003.7, 
    1002.8, 1001.4, 1000.8, 1000.4, 1000.6, 1000.9, 1001.1, 1000.5, 1000.4, 
    1000.2, 1000.3, 1000.8, 1000.7, 1000.7, 1000.8, 1000.9, 1001, 1000.9, 
    1000.9, 1000.8, 1001, 1000.9, 1000.9, 1000.9, 1001.1, 1001.1, 1001.3, 
    1001.5, 1001.6, 1001.5, 1001.6, 1001.4, 1001.4, 1001.4, 1001.2, 1000.8, 
    1000.6, 1000.4, 1000.3, 1000.1, 1000.1, 999.8, 999.5, 999.3, 999, 998.7, 
    998.5, 998.1, 998, 998, 998.1, 998.1, 998, 998, 997.9, 997.8, 998.1, 
    998.1, 998.3, 998.4, 998.6, 998.5, 998.7, 998.9, 999.1, 999.5, 999.8, 
    1000, 1000.5, 1000.9, 1001.2, 1001.3, 1001.4, 1001.6, 1001.9, 1002.1, 
    1002.3, 1002.1, 1002.2, 1002, 1001.8, 1001.7, 1001.2, 1000.7, 1000.1, 
    999.2, 999, 998.8, 998.4, 998, 997.9, 997.9, 998, 998, 998.3, 998.5, 
    998.9, 999.1, 999.7, 1000.3, 1000.8, 1001.3, 1001.9, 1002.5, 1002.9, 
    1003.4, 1003.8, 1004.2, 1004.6, 1004.8, 1005.4, 1005.8, 1006.1, 1006.4, 
    1006.7, 1006.9, 1007.1, 1007.1, 1007.1, 1007.3, 1007.3, 1007.3, 1007.3, 
    1007.6, 1007.5, 1007.6, 1007.8, 1008, 1008.1, 1008.2, 1008.4, 1008.6, 
    1008.8, 1009.1, 1009.4, 1009.8, 1010.3, 1010.6, 1011.1, 1011.5, 1012, 
    1012.4, 1012.7, 1013.1, 1013.1, 1013.2, 1013.6, 1013.8, 1014, 1014.8, 
    1015.2, 1015.5, 1015.8, 1015.8, 1015.7, 1015.3, 1014.9, 1014.5, 1014, 
    1013.7, 1013.3, 1012.8, 1012, 1011.1, 1010.3, 1009.7, 1008.9, 1008.2, 
    1007.6, 1007.2, 1006.8, 1006.3, 1005.9, 1005.6, 1005.3, 1005.1, 1005.1, 
    1005.1, 1005.1, 1005.3, 1005.6, 1005.8, 1006.1, 1006.5, 1006.9, 1007.1, 
    1007.7, 1008.1, 1008.7, 1009.3, 1010, 1010.2, 1010.5, 1010.6, 1011, 1011, 
    1011.4, 1011.3, 1011, 1010.5, 1010.2, 1009.5, 1008.7, 1007.8, 1007, 
    1006.2, 1005.2, 1004.3, 1003.8, 1003.7, 1003.6, 1003.5, 1003.5, 1003.6, 
    1004, 1004.3, 1004.8, 1005.4, 1006.2, 1006.9, 1007.8, 1008.4, 1009.1, 
    1009.6, 1010.3, 1010.8, 1011.5, 1012.2, 1012.8, 1013.4, 1014, 1014.4, 
    1014.4, 1014.7, 1015, 1015.4, 1015.6, 1015.4, 1015, 1014.5, 1014.2, 
    1014.2, 1014.4, 1014, 1013.8, 1014, 1014.1, 1013.8, 1013.5, 1012.8, 
    1012.1, 1011.5, 1010.6, 1009.9, 1009.4, 1008.7, 1008.2, 1007.8, 1007.4, 
    1007.2, 1007.2, 1007.6, 1007.7, 1008.1, 1008.5, 1008.9, 1009.3, 1009.9, 
    1010.4, 1011, 1011.7, 1012.2, 1012.4, 1012.7, 1013.2, 1013.4, 1013.6, 
    1013.7, 1013.9, 1014, 1014.4, 1014.4, 1014.4, 1014.4, 1014.4, 1014.4, 
    1014.4, 1015.2, 1015.9, 1016.2, 1016.6, 1016.9, 1017.3, 1017.7, 1018.1, 
    1018.5, 1018.8, 1018.6, 1018.4, 1018.5, 1018.6, 1018.6, 1018.7, 1018.8, 
    1018.9, 1019.3, 1019.6, 1019.9, 1020.3, 1020.6, 1020.9, 1021.5, 1022.1, 
    1022.6, 1023, 1023.6, 1024, 1024, 1024.3, 1024.3, 1024.3, 1024.3, 1024.1, 
    1023.7, 1023.5, 1023.2, 1022.8, 1022.4, 1021.9, 1021.4, 1020.8, 1020.3, 
    1019.3, 1018.7, 1017.8, 1016.8, 1015.7, 1014.8, 1013.6, 1012.6, 1011.8, 
    1010.8, 1009.7, 1008.7, 1007.9, 1006.6, 1005.7, 1005, 1004.2, 1003.8, 
    1003.5, 1003.2, 1003, 1003, 1002.8, 1002.7, 1002.9, 1003.1, 1003.1, 
    1003.3, 1003.5, 1003.6, 1003.7, 1003.9, 1004.1, 1004.2, 1004.4, 1004.7, 
    1004.1, 1004.1, 1003.9, 1003.9, 1003.8, 1003.6, 1003.5, 1003.3, 1002.9, 
    1002.6, 1002.3, 1001.9, 1001.7, 1001.5, 1001.1, 1000.8, 1000.7, 1000.5, 
    1000.4, 1000.3, 1000.2, 1000.1, 1000.2, 1000.1, 1000, 999.8, 999.8, 
    999.8, 999.8, 999.8, 999.8, 999.8, 999.5, 999.3, 999.1, 999, 998.9, 
    998.8, 998.5, 998.4, 998.3, 998.1, 998.4, 998.4, 998.4, 998.3, 998.4, 
    998.7, 998.8, 999.1, 999.2, 999.5, 999.8, 1000.1, 1000.6, 1001, 1001.4, 
    1001.8, 1002.2, 1002.9, 1003.4, 1004, 1004.7, 1005.5, 1006.1, 1006.8, 
    1007.5, 1008.4, 1009.1, 1009.8, 1010.4, 1011.1, 1011.8, 1012.1, 1012.5, 
    1012.6, 1012.9, 1013.4, 1013.6, 1013.7, 1014.2, 1014.5, 1014.5, 1014.5, 
    1014.8, 1014.7, 1014.8, 1014.9, 1014.9, 1015, 1014.9, 1014.9, 1014.8, 
    1014.8, 1014.8, 1014.9, 1015, 1014.7, 1014.6, 1014.5, 1014.3, 1013.8, 
    1013.6, 1013.6, 1013.2, 1013.1, 1012.6, 1012.5, 1012.4, 1012.1, 1011.6, 
    1011.4, 1010.8, 1010.5, 1010.6, 1010.3, 1010.1, 1009.7, 1009.5, 1009.6, 
    1009.2, 1008.8, 1008.6, 1008.3, 1008, 1007.8, 1007.3, 1007.1, 1006.7, 
    1006.6, 1006.2, 1006, 1006.1, 1005.8, 1005.2, 1004.7, 1004.5, 1004, 
    1003.4, 1003, 1002.3, 1002, 1001.5, 1001, 1000.2, 999.5, 998.9, 998.5, 
    998.3, 997.8, 997.6, 997.6, 997.3, 997, 997, 997, 997.3, 997.6, 998, 
    998.3, 998.6, 999.2, 999.9, 1000.6, 1001.2, 1001.9, 1002.7, 1003.3, 1004, 
    1004.6, 1004.9, 1005.4, 1006.1, 1006.6, 1007.1, 1007.7, 1008.4, 1008.9, 
    1009.4, 1009.9, 1010.4, 1010.8, 1011.1, 1011.7, 1011.8, 1012.3, 1012.6, 
    1013, 1013.3, 1013.5, 1013.6, 1013.7, 1013.9, 1014, 1014, 1014, 1013.8, 
    1013.9, 1013.9, 1014.1, 1014.1, 1014.1, 1014.2, 1014.2, 1014.1, 1014.1, 
    1014.1, 1014.1, 1014.2, 1014.3, 1014.3, 1014.2, 1014.4, 1014.4, 1014.4, 
    1014.3, 1014.6, 1014.7, 1014.8, 1014.9, 1015.1, 1015.1, 1015.2, 1015.2, 
    1015.1, 1015.3, 1015.3, 1015.3, 1015.4, 1015.5, 1015.3, 1015.1, 1015, 
    1015, 1015, 1014.7, 1014.7, 1014.7, 1014.5, 1014.2, 1014, 1013.7, 1013.2, 
    1013, 1012.6, 1012.4, 1012.2, 1012.2, 1011.7, 1011.3, 1010.7, 1010.2, 
    1010.1, 1009.9, 1009.2, 1008.5, 1007.9, 1007.6, 1007.3, 1007.1, 1006.7, 
    1006.1, 1006, 1005.7, 1005.4, 1004.8, 1004.6, 1004.1, 1003.7, 1003.2, 
    1002.7, 1002.1, 1001.6, 1000.9, 1000.5, 1000.1, 999.7, 999.2, 998.7, 
    998.3, 997.9, 997.6, 997.3, 997.2, 997.1, 997.2, 997.1, 997, 997.1, 
    997.2, 997.3, 997.3, 997.5, 997.6, 997.6, 997.7, 998.1, 998.4, 998.6, 
    998.9, 999.1, 999.6, 999.8, 1000.1, 1000.3, 1000.5, 1000.7, 1001.2, 
    1001.6, 1002, 1002.4, 1002.7, 1003.2, 1003.5, 1003.8, 1004.2, 1004.4, 
    1004.8, 1005.2, 1005.6, 1006.1, 1006.5, 1007, 1007.2, 1007.6, 1007.8, 
    1008.2, 1008.5, 1008.7, 1008.7, 1008.5, 1008.9, 1009, 1009, 1008.9, 
    1008.4, 1007.7, 1007.3, 1006.9, 1005.6, 1004.7, 1003.5, 1003.1, 1002.9, 
    1001.7, 1001.1, 1000.2, 999.9, 1000.1, 1000, 1000.2, 999.7, 999.3, 999.4, 
    999.4, 999.3, 999.2, 998.8, 998.8, 998.6, 998.6, 998.4, 998.1, 997.3, 
    997.3, 997.2, 997.2, 996.9, 996.2, 995.7, 995.2, 994.9, 994.7, 994.4, 
    994.2, 994.1, 993.9, 994.1, 994.5, 995.4, 996.1, 996.9, 997.8, 998.7, 
    999.3, 1000.2, 1000.9, 1001.4, 1002.2, 1002.4, 1002.7, 1003.3, 1003.8, 
    1004.4, 1005, 1005.6, 1006.4, 1006.9, 1007.4, 1008.1, 1008.6, 1009.2, 
    1009.5, 1009.9, 1010.5, 1011, 1011.2, 1011.3, 1011.4, 1011.5, 1011.4, 
    1011.3, 1010.8, 1010.9, 1010.6, 1010.3, 1010, 1009.7, 1009.3, 1008.7, 
    1008.2, 1007.6, 1006.9, 1005.9, 1005.3, 1004.8, 1004.4, 1003.9, 1004, 
    1003.2, 1002.3, 1001.3, 1000.2, 999.4, 998.8, 998.3, 997.3, 996.9, 996.6, 
    996.3, 995.9, 995.6, 995.4, 995.2, 995, 995, 995.1, 995.3, 995.5, 995.9, 
    996.4, 997, 997.7, 998.3, 999, 999.7, 1000.5, 1001.3, 1002, 1002.5, 1003, 
    1003.5, 1004.1, 1004.4, 1004.8, 1005.3, 1005.7, 1006, 1006.2, 1006.6, 
    1006.9, 1007.3, 1007.3, 1007.4, 1007.7, 1008.3, 1008.5, 1008.9, 1009.2, 
    1009.4, 1009.7, 1010, 1010.3, 1010.4, 1010.7, 1010.6, 1010.9, 1011, 
    1011.1, 1011.2, 1011.2, 1011.4, 1011.5, 1011.5, 1011.6, 1011.4, 1011.7, 
    1011.7, 1011.9, 1011.8, 1011.8, 1012, 1012.2, 1012.3, 1012.2, 1012, 1012, 
    1012, 1012, 1011.7, 1011.6, 1011.6, 1011.7, 1011.7, 1011.6, 1011.6, 
    1011.4, 1011.4, 1011.3, 1011.1, 1011, 1010.9, 1010.8, 1010.7, 1011.1, 
    1011.2, 1010.8, 1010.7, 1010.5, 1010.3, 1010, 1009.7, 1009.4, 1008.5, 
    1008.2, 1007.7, 1007.5, 1007, 1006.7, 1006.1, 1005.7, 1005.4, 1005, 
    1004.8, 1004.2, 1003.3, 1003, 1002.6, 1002.1, 1001.5, 1001.2, 1000.9, 
    1000.3, 999.8, 999.3, 999.3, 999, 998.5, 998.2, 998.2, 998.2, 998.3, 
    998.3, 998.2, 998.2, 998.2, 998.2, 998.3, 998.4, 998.4, 998.5, 998.6, 
    998.9, 999, 999.1, 999.3, 999.2, 999, 998.6, 998.3, 998, 997.7, 997.7, 
    997.3, 997, 996.7, 996.4, 995.8, 995.5, 995.2, 994.8, 994.4, 993.8, 
    993.3, 992.9, 992.6, 992.3, 991.8, 991.7, 991.1, 990.7, 990.7, 990.6, 
    990.3, 990.2, 990.2, 990.4, 990.4, 990.8, 991.1, 991.2, 991.4, 991.6, 
    991.9, 992.1, 992.2, 992.6, 992.9, 993.6, 994.5, 995.1, 995.7, 996.3, 
    996.4, 996.8, 997.3, 997.6, 997.9, 998.3, 998.7, 999, 999.6, 1000, 
    1000.4, 1000.7, 1001.1, 1001.4, 1001.7, 1001.9, 1002.2, 1002.4, 1002.5, 
    1002.9, 1003.1, 1003.5, 1003.7, 1003.9, 1004, 1004.1, 1004.2, 1004.2, 
    1004.2, 1004.3, 1004.5, 1004.5, 1004.7, 1005, 1005, 1005, 1005.5, 1005.3, 
    1005.3, 1005.4, 1005.4, 1005.4, 1005.5, 1005.8, 1005.9, 1006.4, 1006.3, 
    1006.6, 1006.9, 1006.9, 1007.1, 1007.2, 1007.2, 1007.3, 1007.5, 1007.6, 
    1008.1, 1008.2, 1008.6, 1008.6, 1009.1, 1009.1, 1009.7, 1010, 1010.3, 
    1010.6, 1010.6, 1010.7, 1010.8, 1011, 1010.9, 1010.8, 1010.8, 1011.1, 
    1011.2, 1011, 1011.1, 1011, 1011.2, 1011.5, 1011.8, 1011.7, 1011.9, 
    1011.8, 1011.8, 1011.7, 1011.4, 1011.1, 1010.9, 1010.5, 1010.2, 1009.9, 
    1009.6, 1009.2, 1008.8, 1008.1, 1007.5, 1006.9, 1006.2, 1005.6, 1004.8, 
    1004.3, 1003.9, 1004.1, 1004.3, 1004.8, 1005.8, 1006.5, 1007.4, 1008, 
    1008.6, 1009.1, 1009.6, 1010.1, 1010.8, 1011.3, 1012, 1012.7, 1013.1, 
    1013.7, 1014.1, 1014.5, 1014.8, 1014.9, 1015.1, 1015.1, 1015.3, 1015.4, 
    1015.4, 1015.7, 1015.5, 1015.4, 1015.4, 1015.6, 1015.4, 1015.4, 1015.2, 
    1015.2, 1015.4, 1015.4, 1015.6, 1015.4, 1015.3, 1015.7, 1015.6, 1015.5, 
    1015.4, 1015.3, 1015.4, 1015.4, 1015.3, 1015.2, 1014.9, 1015, 1015.1, 
    1015.1, 1015.1, 1014.9, 1014.8, 1014.9, 1014.6, 1014.4, 1014.3, 1014.3, 
    1014.4, 1014.2, 1014.3, 1014.2, 1014.1, 1013.8, 1013.9, 1013.9, 1013.9, 
    1013.8, 1013.8, 1013.8, 1013.8, 1013.7, 1013.8, 1013.8, 1013.7, 1013.5, 
    1013.4, 1013.3, 1013.1, 1012.9, 1013.1, 1013.2, 1013.2, 1013.2, 1013.3, 
    1013.3, 1013.3, 1013.4, 1013, 1012.7, 1012.7, 1012.6, 1012.6, 1012.8, 
    1012.9, 1013.1, 1013, 1013.1, 1013.3, 1013.1, 1013.1, 1013.3, 1013.3, 
    1013.5, 1013.5, 1013.8, 1013.9, 1013.9, 1014.1, 1014.1, 1014.3, 1014.3, 
    1014.1, 1014, 1013.7, 1013.7, 1013.6, 1013.5, 1013.4, 1013.5, 1013.3, 
    1013.2, 1013.1, 1012.9, 1012.6, 1012, 1011.6, 1011.5, 1011.5, 1011.2, 
    1011, 1011, 1010.8, 1010.8, 1011, 1011.1, 1011.1, 1010.9, 1010.5, 1010.3, 
    1010, 1009.6, 1009.1, 1008.8, 1008.4, 1007.9, 1007.3, 1006.7, 1006.4, 
    1006, 1005.4, 1004.7, 1004.5, 1004.2, 1003.9, 1003.7, 1003.4, 1003.7, 
    1003.9, 1003.8, 1004, 1003.9, 1004, 1004, 1004.3, 1004.9, 1004.8, 1004.5, 
    1004.4, 1004.6, 1004.9, 1005, 1005.3, 1005.5, 1005.9, 1006.2, 1006.6, 
    1007, 1007.4, 1007.5, 1007.9, 1007.9, 1007.9, 1008, 1007.7, 1007.7, 
    1007.5, 1007.2, 1006.7, 1006.5, 1006.3, 1006.1, 1005.6, 1005.2, 1004.7, 
    1004.1, 1003.4, 1003, 1002.5, 1002, 1002.2, 1002.2, 1002.6, 1002.8, 
    1002.2, 1001.8, 1001.5, 1001, 1000.4, 1000, 999.4, 999.4, 999.1, 999.1, 
    999.6, 999.4, 1000, 1000.3, 1001.2, 1001.6, 1002.5, 1003.3, 1003.9, 
    1004.4, 1005, 1005.6, 1006.4, 1006.9, 1007, 1007, 1006.8, 1006.9, 1007, 
    1007.1, 1007.3, 1007.6, 1007.9, 1008.2, 1008.6, 1008.9, 1009.2, 1009.5, 
    1009.4, 1009.7, 1009.5, 1009.5, 1009.2, 1008.6, 1008.1, 1007.5, 1006.6, 
    1005.5, 1004.9, 1004.1, 1003.4, 1002.9, 1002.5, 1002.5, 1002.3, 1002.4, 
    1002.7, 1003, 1003.1, 1003.4, 1003.8, 1004.1, 1004.3, 1004.6, 1004.7, 
    1005, 1005, 1005.4, 1005.8, 1006.4, 1006.8, 1007.5, 1008, 1008.4, 1008.9, 
    1009.3, 1009.4, 1009.5, 1009.6, 1009.5, 1009.4, 1009.4, 1009.4, 1009.1, 
    1008.7, 1008.5, 1008.2, 1007.5, 1006.9, 1006, 1005.3, 1004.6, 1003.9, 
    1003.7, 1003.3, 1002.8, 1002.6, 1002.4, 1002.2, 1002.3, 1002.4, 1002.6, 
    1003, 1003.4, 1003.8, 1004.3, 1004.9, 1005.1, 1006, 1006.2, 1006.6, 
    1007.1, 1007.3, 1007.4, 1007.6, 1007.7, 1007.8, 1007.8, 1007.8, 1007.8, 
    1007.6, 1007.7, 1007.6, 1007.4, 1007.3, 1006.9, 1006.6, 1006.4, 1006.1, 
    1005.8, 1006, 1006, 1006, 1005.6, 1005.2, 1005.3, 1004.9, 1004.6, 1004.2, 
    1003.7, 1003.7, 1004.1, 1004.2, 1004.6, 1005, 1005.4, 1006, 1006.5, 
    1006.7, 1007, 1007.7, 1008.4, 1008.8, 1009.3, 1009.5, 1010.1, 1010.3, 
    1010.7, 1011.4, 1011.7, 1011.9, 1011.9, 1012.1, 1012.3, 1012.6, 1012.8, 
    1013.1, 1013.1, 1013.4, 1013.5, 1013.6, 1013.7, 1013.9, 1014.2, 1014.4, 
    1014.7, 1014.9, 1015.3, 1015.8, 1016.2, 1016.7, 1017.1, 1017.5, 1017.9, 
    1018.1, 1018.3, 1018.6, 1018.4, 1018.5, 1018.4, 1018.5, 1018.5, 1018.1, 
    1018.1, 1018, 1017.7, 1017.4, 1017.2, 1016.9, 1016.8, 1016.8, 1016.9, 
    1017.3, 1017.4, 1017.3, 1017.4, 1017.6, 1017.8, 1017.4, 1017.4, 1017.2, 
    1016.9, 1016.8, 1016.2, 1015.8, 1015.1, 1014.3, 1013.5, 1013.1, 1012.3, 
    1011.3, 1010.5, 1009.8, 1008.5, 1007.8, 1007, 1006.3, 1005.8, 1005, 1005, 
    1005.1, 1005, 1004.9, 1004.5, 1003.9, 1003.7, 1003.2, 1002.8, 1002.5, 
    1002, 1001.8, 1001.6, 1001.7, 1001.8, 1002, 1002, 1002, 1001.9, 1001.8, 
    1002, 1002.2, 1002.5, 1002.9, 1003.2, 1003.6, 1004.1, 1004.5, 1004.8, 
    1005.1, 1005.4, 1005.8, 1006.2, 1006.4, 1007, 1007.4, 1008, 1008.6, 
    1009.2, 1009.6, 1009.9, 1010.1, 1010.5, 1010.8, 1011.1, 1011.3, 1011.5, 
    1011.6, 1011.7, 1011.5, 1011.4, 1010.9, 1010.7, 1010.3, 1010, 1009.9, 
    1009.5, 1009.1, 1008.8, 1008.6, 1008.4, 1008, 1007.4, 1007, 1006.3, 1006, 
    1005.7, 1005.4, 1005.3, 1005.3, 1005.1, 1004.8, 1004.9, 1004.7, 1004.6, 
    1004.2, 1004.1, 1003.8, 1003.5, 1003.4, 1003.2, 1003, 1002.9, 1003.2, 
    1002.9, 1002.8, 1002.5, 1002.3, 1001.9, 1001.8, 1001.7, 1001.2, 1001.3, 
    1001, 1001, 1000.7, 1000.4, 1000.1, 999.8, 999.5, 999.2, 999.4, 999.5, 
    999.7, 999.8, 1000, 1000.4, 1000.8, 1001.4, 1002.3, 1002.9, 1003.1, 
    1003.5, 1003.8, 1004.2, 1005.1, 1005.6, 1005.9, 1006.5, 1006.8, 1007.4, 
    1007.8, 1008, 1008.1, 1008.2, 1008.5, 1008.5, 1008.6, 1008.4, 1008.2, 
    1007.9, 1007.8, 1007.6, 1007.1, 1006.8, 1006.5, 1005.9, 1005.7, 1005.5, 
    1005.4, 1005.1, 1005, 1005.3, 1005.5, 1005.6, 1005.7, 1005.5, 1005.4, 
    1005.2, 1005.2, 1005.6, 1006.2, 1006.6, 1007.6, 1008.7, 1009.4, 1009.9, 
    1009.9, 1010.4, 1010.7, 1010.9, 1010.8, 1011.1, 1011.1, 1011.5, 1011.6, 
    1011.9, 1012.1, 1012.4, 1012.7, 1012.7, 1012.8, 1012.8, 1013.1, 1012.9, 
    1013.4, 1014.2, 1014.9, 1016, 1016.6, 1016.8, 1017.4, 1017.6, 1017.5, 
    1017.9, 1017.8, 1017.7, 1017.3, 1016.8, 1016.1, 1015.4, 1014.8, 1014.2, 
    1013.7, 1013.5, 1013.6, 1013.4, 1013.4, 1013.7, 1013.9, 1014, 1014.5, 
    1014.5, 1014.8, 1015.4, 1015.5, 1015.8, 1016, 1016.3, 1016.3, 1016.6, 
    1016.6, 1016.6, 1016.8, 1016.9, 1016.7, 1016.5, 1016.5, 1016.4, 1016.5, 
    1016.5, 1016.6, 1016.4, 1016.5, 1016.8, 1017.4, 1017.8, 1017.9, 1018.2, 
    1018.5, 1018.7, 1018.6, 1018.7, 1019.1, 1019.2, 1019.7, 1020.2, 1020.6, 
    1020.7, 1021.1, 1021.4, 1021.8, 1022, 1022.1, 1022.1, 1022.3, 1022.2, 
    1022.1, 1022.1, 1022.2, 1022.3, 1022.3, 1022.3, 1022.5, 1022.4, 1022.4, 
    1022.3, 1021.9, 1021.7, 1021.7, 1021.7, 1021.7, 1021.7, 1021.4, 1021.3, 
    1021.1, 1021.1, 1021, 1020.7, 1020.3, 1020, 1019.8, 1019.8, 1020, 1019.9, 
    1019.7, 1019.6, 1019.2, 1018.9, 1018.8, 1018.4, 1017.8, 1018, 1018.1, 
    1018.6, 1018.7, 1018.7, 1018.8, 1018.6, 1018.6, 1018.6, 1018.6, 1018.6, 
    1018.7, 1018.7, 1018.3, 1018.2, 1018.3, 1018.6, 1018.8, 1018.5, 1018.4, 
    1018.5, 1018.3, 1018, 1017.5, 1017.6, 1017.7, 1017.6, 1017.7, 1017.5, 
    1017.2, 1017.1, 1017.2, 1017.1, 1017, 1017.2, 1017.2, 1017.3, 1017.5, 
    1017.5, 1017.6, 1017.6, 1017.6, 1017.8, 1018.3, 1018.6, 1018.9, 1019.3, 
    1019.6, 1019.6, 1019.9, 1019.9, 1020, 1019.9, 1020, 1020, 1019.9, 1019.9, 
    1020, 1019.8, 1019.7, 1019.5, 1019.3, 1019.3, 1019.2, 1019.2, 1019.2, 
    1018.9, 1018.8, 1018.6, 1018.3, 1018.1, 1017.8, 1017.6, 1017.2, 1016.9, 
    1016.7, 1016.4, 1016.4, 1016.1, 1015.9, 1015.6, 1015.4, 1015.1, 1014.8, 
    1014.5, 1014.1, 1014, 1013.9, 1013.8, 1013.6, 1013.4, 1013.3, 1013.1, 
    1012.7, 1012.6, 1012.3, 1012.2, 1012, 1012, 1012, 1011.9, 1012, 1011.7, 
    1012, 1011.9, 1012, 1012.1, 1012, 1012.1, 1012.3, 1012.6, 1012.9, 1013.2, 
    1013.4, 1013.5, 1013.5, 1013.7, 1013.7, 1013.8, 1013.5, 1013.2, 1013.4, 
    1013.2, 1013.2, 1013.2, 1013.2, 1012.9, 1012.7, 1012.5, 1012.1, 1011.8, 
    1011.2, 1010.4, 1010.2, 1009.8, 1009.7, 1009.4, 1009.1, 1008.8, 1008.5, 
    1008.3, 1008, 1007.5, 1007.2, 1007, 1006.3, 1006.1, 1005.6, 1005.1, 
    1004.9, 1004.1, 1003.6, 1003.3, 1002.1, 1002.4, 1002.1, 1001.7, 1001.5, 
    1001.1, 1000.4, 1000, 999.4, 999.1, 998.6, 998.6, 998.4, 998, 997.7, 
    997.4, 997.3, 997.6, 997.3, 997.9, 998.5, 998.1, 998.4, 999, 999, 999.1, 
    999.5, 999.4, 999.5, 999.8, 1000.1, 1000.4, 1000.7, 1001, 1001.2, 1001.4, 
    1001.5, 1001.6, 1001.8, 1002, 1002.3, 1002.6, 1002.8, 1003.1, 1003.3, 
    1003.4, 1003.5, 1003.5, 1003.7, 1003.7, 1003.6, 1003.7, 1003.9, 1004.1, 
    1004.2, 1004.3, 1004.3, 1004.4, 1004.7, 1004.8, 1004.9, 1004.9, 1005.2, 
    1005.3, 1005.4, 1005.7, 1005.9, 1006.4, 1006.7, 1006.9, 1007.1, 1007.3, 
    1007.7, 1007.7, 1007.8, 1008, 1008.3, 1008.6, 1009, 1009.2, 1009.5, 
    1009.8, 1009.9, 1010.1, 1010.2, 1010.4, 1010.6, 1010.7, 1010.7, 1010.9, 
    1011.2, 1011.5, 1011.6, 1011.8, 1011.8, 1011.9, 1012, 1011.9, 1011.9, 
    1011.6, 1011.7, 1011.8, 1011.7, 1011.9, 1011.7, 1011.6, 1011.5, 1011.4, 
    1011.2, 1010.9, 1010.8, 1010.6, 1010.6, 1010.5, 1010.4, 1010.4, 1010.3, 
    1010, 1010.1, 1010.1, 1009.9, 1009.6, 1009.5, 1009.4, 1009.3, 1009.2, 
    1009.1, 1009.3, 1009.3, 1009.3, 1009.3, 1009.3, 1009.1, 1009, 1008.8, 
    1008.9, 1009.1, 1009.1, 1009.2, 1009.3, 1009.1, 1009.1, 1009.1, 1009.1, 
    1009, 1009.1, 1009, 1008.8, 1008.7, 1008.5, 1008.6, 1008.5, 1008.6, 
    1008.5, 1008.4, 1008.4, 1008.3, 1008.3, 1008.2, 1008.1, 1008.1, 1008, 
    1007.7, 1007.7, 1007.6, 1007.9, 1007.8, 1008, 1008, 1008, 1007.9, 1007.8, 
    1007.7, 1007.7, 1007.7, 1007.9, 1007.9, 1008.1, 1008.1, 1008.2, 1008.1, 
    1008.1, 1008.1, 1008, 1007.9, 1007.8, 1007.8, 1007.9, 1008.1, 1008.2, 
    1008.4, 1008.3, 1008.5, 1008.5, 1008.5, 1008.5, 1008.5, 1008.6, 1008.7, 
    1008.8, 1008.9, 1009.1, 1009.1, 1009.2, 1009.3, 1009.4, 1009.4, 1009.5, 
    1009.7, 1009.8, 1009.8, 1010, 1010.3, 1010.4, 1010.6, 1010.8, 1011.1, 
    1011, 1011.1, 1011.2, 1011.4, 1011.5, 1011.6, 1011.7, 1011.8, 1011.9, 
    1011.7, 1011.6, 1011.5, 1011.4, 1011.5, 1011.1, 1010.9, 1010.7, 1010.9, 
    1010.7, 1010.5, 1010.3, 1010.2, 1009.9, 1009.6, 1009.2, 1008.7, 1008.2, 
    1007.8, 1007.2, 1006.8, 1006.5, 1006.2, 1005.4, 1004.7, 1004.4, 1003.8, 
    1003.1, 1002.6, 1001.8, 1001, 1000, 999.2, 998.4, 997.1, 996, 995.4, 
    994.2, 992.7, 991.4, 989.8, 988.1, 986.7, 985.9, 985.7, 985.1, 984.9, 
    984.6, 984.8, 984.6, 984.5, 984.5, 984.2, 984.3, 984.3, 984.2, 984.5, 
    984.6, 984.6, 984.8, 984.8, 984.8, 984.7, 984.8, 984.8, 984.7, 984.8, 
    984.9, 985, 985, 985.2, 985.2, 985.5, 985.5, 985.7, 985.8, 985.9, 985.9, 
    985.9, 986, 986, 986.1, 986.3, 986.5, 986.6, 986.6, 986.6, 986.7, 986.7, 
    986.6, 986.7, 986.7, 987, 987.2, 987.3, 987.5, 987.6, 987.7, 988, 988.4, 
    988.6, 989.2, 989.5, 989.8, 990.4, 990.9, 991.4, 991.6, 992, 992.5, 
    992.6, 992.8, 992.9, 993.1, 993.9, 994.3, 994.9, 995.1, 995.7, 996, 
    996.4, 996.8, 997.1, 997.6, 998, 998.2, 998.6, 998.8, 999.4, 999.7, 
    999.9, 1000.3, 1000.6, 1000.6, 1000.6, 1000.9, 1001.2, 1001.4, 1001.4, 
    1001.5, 1001.7, 1001.9, 1002.3, 1002.5, 1002.8, 1003.2, 1003.2, 1003.5, 
    1004, 1004.8, 1004.9, 1005.1, 1005.5, 1005.8, 1006.1, 1006.4, 1006.8, 
    1006.9, 1007.1, 1007.3, 1007.4, 1007.8, 1008, 1008.4, 1008.5, 1008.9, 
    1009.2, 1009.5, 1009.6, 1010, 1010.2, 1010, 1010.1, 1010.4, 1010.5, 
    1010.5, 1010.5, 1010.6, 1010.7, 1010.9, 1011, 1010.9, 1010.9, 1010.9, 
    1010.9, 1010.9, 1011, 1011.1, 1011.1, 1011.3, 1011.3, 1011.3, 1011.5, 
    1011.6, 1011.6, 1011.5, 1011.6, 1011.7, 1011.6, 1011.7, 1011.8, 1011.9, 
    1012, 1012, 1011.9, 1011.9, 1011.6, 1011.2, 1010.9, 1010.9, 1010.7, 
    1010.4, 1009.9, 1009.4, 1008.7, 1008.5, 1008.1, 1007.6, 1007.6, 1006.6, 
    1006.3, 1005.5, 1004.8, 1004.3, 1003.6, 1003.1, 1002.7, 1002.2, 1001.7, 
    1001.2, 1000.6, 1000.4, 1000.1, 999.8, 999.6, 999.5, 999.4, 999.5, 999.6, 
    999.7, 1000, 1000.3, 1000.5, 1000.9, 1001.4, 1001.8, 1002.2, 1002.6, 
    1003.1, 1003.7, 1004, 1004.6, 1004.9, 1005.2, 1005.3, 1005.6, 1005.6, 
    1005.8, 1006.1, 1006.3, 1006.4, 1006.4, 1006.5, 1006.6, 1006.7, 1006.8, 
    1006.9, 1007, 1007, 1007.1, 1007.3, 1007.3, 1007.3, 1007.4, 1007.5, 
    1007.7, 1007.9, 1008.2, 1008.3, 1008.5, 1008.8, 1009.1, 1009.5, 1009.9, 
    1010.3, 1010.6, 1011.2, 1011.6, 1011.9, 1012.2, 1012.5, 1012.8, 1013.1, 
    1013.5, 1013.8, 1014, 1014, 1014.1, 1014.1, 1014.2, 1013.9, 1013.7, 
    1013.3, 1013, 1012.6, 1012.4, 1012, 1011.8, 1011.7, 1012.2, 1012.2, 
    1012.2, 1012.2, 1012, 1011.8, 1011.6, 1011.3, 1010.6, 1010, 1009.4, 
    1008.4, 1008.1, 1007.7, 1007.2, 1006.5, 1005.7, 1004.9, 1003.9, 1002.8, 
    1001.9, 1000.8, 999.8, 998.7, 997.2, 996.1, 994.4, 992.4, 990.7, 989.1, 
    987.4, 987.2, 989.1, 990.6, 990.9, 991.7, 991.5, 990.9, 990.8, 990.8, 
    991.7, 991.8, 991.4, 991.8, 992.2, 992.8, 994, 995.3, 996.3, 997.5, 
    998.3, 999, 1000.5, 1002, 1003.3, 1004.5, 1005.2, 1005.5, 1006.7, 1007.2, 
    1008.3, 1009, 1009.8, 1010, 1010.1, 1010.2, 1010.3, 1010.1, 1009.9, 
    1009.9, 1009.7, 1009.4, 1009.5, 1009.7, 1010, 1010.2, 1010.1, 1009.9, 
    1009.6, 1009.5, 1009.5, 1009.1, 1009, 1008.5, 1008.4, 1008.1, 1007.7, 
    1006.9, 1006.3, 1005.5, 1005.2, 1004.6, 1004.1, 1003.9, 1003.8, 1004, 
    1003.9, 1004, 1003.8, 1003.6, 1003.5, 1003.2, 1002.8, 1002.6, 1002.2, 
    1002, 1001.8, 1001.5, 1001.4, 1001.4, 1001.4, 1001.3, 1001, 1000.3, 
    999.8, 999.5, 999.2, 998.4, 997.9, 996.6, 995.4, 994.2, 992.9, 991.9, 
    991.2, 990.8, 990.7, 991, 991.7, 992.3, 993.1, 994.1, 994.9, 996, 996.9, 
    997.9, 998.9, 999.8, 1000.8, 1001.9, 1003, 1004, 1005, 1006.1, 1007, 
    1008, 1009, 1010, 1010.8, 1011.3, 1012.1, 1012.6, 1013.4, 1014.2, 1015, 
    1015.8, 1016.5, 1017, 1017.3, 1017.7, 1018.2, 1018.4, 1018.5, 1018.8, 
    1019, 1019.2, 1019.1, 1019, 1018.6, 1018.3, 1017.7, 1017.1, 1016.4, 
    1015.6, 1014.8, 1014.2, 1013.7, 1013.2, 1012.5, 1011.9, 1011.1, 1010.7, 
    1010.5, 1009.8, 1009.9, 1010.5, 1010.8, 1011.2, 1011.5, 1011.8, 1012, 
    1012.6, 1013.1, 1013.6, 1014, 1014.5, 1015, 1015.4, 1015.9, 1016.5, 
    1017.1, 1017.7, 1018.2, 1018.7, 1019.1, 1019.4, 1019.8, 1020, 1020.3, 
    1020.3, 1020.4, 1020.4, 1019.9, 1019.9, 1019.7, 1019.4, 1018.9, 1018.4, 
    1017.8, 1017.6, 1017.1, 1016.8, 1016.2, 1015.8, 1015.7, 1015.6, 1015.7, 
    1015.6, 1015.7, 1016, 1015.9, 1015.9, 1015.8, 1015.8, 1015.7, 1015.7, 
    1016, 1015.7, 1015.7, 1015.5, 1015.2, 1015.1, 1014.9, 1014.6, 1014.3, 
    1014, 1013.9, 1013.5, 1013.3, 1013.3, 1013.2, 1013.1, 1013.1, 1013.3, 
    1013.3, 1013.2, 1013.4, 1013.4, 1013.4, 1013.7, 1013.8, 1014.1, 1014.4, 
    1014.7, 1015.1, 1015.5, 1015.8, 1016.1, 1016.3, 1016.5, 1016.7, 1016.8, 
    1016.8, 1016.9, 1017, 1016.9, 1016.8, 1016.7, 1017, 1017.3, 1017.3, 
    1017.1, 1016.9, 1016.6, 1016.7, 1016.6, 1016.7, 1016.7, 1016.5, 1016.3, 
    1016.1, 1016.1, 1016.2, 1016.1, 1015.8, 1015.6, 1015.7, 1015.9, 1015.9, 
    1016.1, 1016.1, 1016, 1015.7, 1015.7, 1015.6, 1015.5, 1015.5, 1015.1, 
    1014.8, 1014.8, 1014.6, 1014.2, 1014.2, 1013.8, 1013.6, 1013.2, 1013, 
    1012.8, 1012.5, 1012.1, 1011.7, 1011.4, 1011, 1010.9, 1010.5, 1010.1, 
    1009.9, 1009.8, 1009.5, 1009.2, 1008.9, 1008.8, 1008.5, 1008.1, 1008, 
    1008, 1008.4, 1008.3, 1007.8, 1007.8, 1008.1, 1008, 1008.2, 1008.1, 
    1008.4, 1008.5, 1008.4, 1008.5, 1008.6, 1008.6, 1008.5, 1008.5, 1008.3, 
    1008, 1007.7, 1007.3, 1007.1, 1007, 1006.9, 1006.8, 1006.7, 1006.6, 
    1006.5, 1006.4, 1006.2, 1006, 1005.6, 1005.3, 1005, 1004.7, 1004.5, 
    1004.4, 1004.3, 1004, 1004, 1003.8, 1003.7, 1003.7, 1003.8, 1003.6, 
    1003.8, 1004.3, 1004.6, 1004.9, 1005.3, 1005.4, 1005.7, 1006, 1006.1, 
    1006.2, 1006.2, 1006.3, 1006.3, 1006.5, 1006.7, 1007, 1007, 1007.2, 
    1007.1, 1006.9, 1006.9, 1007.1, 1007.2, 1007.2, 1007.2, 1007.4, 1007.8, 
    1008.3, 1008.8, 1009.2, 1009.2, 1009.4, 1009.7, 1009.9, 1010.2, 1010.5, 
    1010.9, 1011.3, 1011.6, 1012, 1012.4, 1012.6, 1012.8, 1013, 1013.3, 
    1013.4, 1013.6, 1014, 1014.1, 1014.4, 1014.6, 1014.9, 1015, 1015.1, 
    1015.4, 1015.5, 1015.5, 1015.6, 1015.6, 1015.9, 1015.9, 1016.1, 1016.2, 
    1016.2, 1016.4, 1016.3, 1016.1, 1015.9, 1016, 1015.8, 1015.8, 1015.8, 
    1015.9, 1015.5, 1015.4, 1015.2, 1015, 1014.7, 1014.3, 1013.7, 1013.6, 
    1013.4, 1013.1, 1013.1, 1012.9, 1012.8, 1012.8, 1012.7, 1012.6, 1012.3, 
    1012.1, 1012.2, 1012.2, 1012.2, 1012.2, 1012.2, 1012.4, 1012.4, 1012.4, 
    1012.4, 1012.7, 1012.6, 1012.6, 1012.7, 1012.8, 1012.9, 1013.1, 1013.4, 
    1013.6, 1013.9, 1014, 1014.1, 1014.2, 1014.2, 1014.3, 1014.6, 1014.6, 
    1014.8, 1015, 1015.1, 1015, 1015, 1014.9, 1014.8, 1014.9, 1014.7, 1014.6, 
    1014.5, 1014.6, 1014.6, 1014.6, 1014.5, 1014.4, 1014.1, 1014.1, 1013.5, 
    1013.2, 1013.1, 1012.7, 1012.7, 1012.3, 1012.1, 1011.9, 1011.7, 1011.2, 
    1011, 1011, 1010.6, 1010.4, 1010.4, 1010.1, 1009.9, 1009.6, 1009.3, 
    1009.4, 1009.2, 1008.9, 1008.2, 1008.1, 1008.3, 1008.1, 1007.8, 1007.7, 
    1007.3, 1006.9, 1006.6, 1006.3, 1006.2, 1006.5, 1006.4, 1006.3, 1006.4, 
    1006.4, 1005.9, 1005.6, 1005.6, 1005.6, 1005.7, 1005.6, 1005.5, 1005.3, 
    1005.3, 1005.2, 1005.2, 1005.3, 1005.5, 1005.7, 1005.7, 1005.7, 1005.8, 
    1005.6, 1005.1, 1005.1, 1004.8, 1004.5, 1004.7, 1004.9, 1004.7, 1004.3, 
    1004.1, 1004, 1004, 1003.9, 1004.1, 1003.5, 1003.3, 1002.8, 1002.8, 
    1002.3, 1001.7, 1001, 1000.5, 999.8, 998.8, 998.2, 997.5, 996.3, 995, 
    993.5, 992.5, 991.2, 991, 990.2, 989, 987.8, 987.4, 986.4, 985.5, 983.9, 
    982.5, 981.2, 980.8, 980.1, 979.2, 978.9, 978.9, 978.6, 978.2, 978.2, 
    977.9, 977.6, 977.2, 977.3, 977.3, 977.4, 977.3, 977.1, 977.1, 977.1, 
    977, 976.8, 976.8, 976.6, 976.7, 976.9, 977.1, 977.2, 977.2, 977.4, 
    977.7, 977.8, 977.8, 978, 978.2, 978.6, 978.8, 979.1, 979.5, 979.8, 
    980.3, 980.8, 981.1, 981.6, 981.9, 982.3, 982.5, 982.7, 982.7, 982.9, 
    983.2, 983.6, 983.9, 984, 983.9, 984.1, 984.1, 984.2, 984.2, 984.2, 
    984.5, 984.7, 985, 985.3, 985.8, 986.3, 986.6, 986.8, 987.1, 987.5, 
    987.8, 988.1, 988.5, 988.7, 989.1, 989.5, 989.6, 989.9, 990.1, 990.2, 
    990.3, 990.4, 990.4, 990.5, 990.7, 990.9, 991.1, 991.5, 991.9, 992.1, 
    992.3, 992.4, 992.6, 992.7, 993.2, 993.4, 993.8, 993.9, 994.3, 994.5, 
    994.5, 994.6, 994.7, 994.8, 994.9, 995.1, 994.9, 995.2, 995.1, 995, 
    995.2, 995.2, 995.3, 995.3, 995.5, 995.4, 995.5, 995.5, 995.5, 995.5, 
    995.5, 995.3, 995.4, 995.7, 995.7, 995.8, 995.8, 995.7, 996.1, 996.4, 
    996.8, 997.2, 997.6, 997.9, 998.3, 998.5, 999.1, 999.3, 999.5, 999.7, 
    1000.1, 1000.2, 1000.4, 1000.4, 1000.9, 1001.1, 1001.5, 1001.9, 1002.4, 
    1002.4, 1002.5, 1002.7, 1003, 1003.2, 1003.2, 1003.6, 1004.1, 1004.5, 
    1004.8, 1005.1, 1005.7, 1006.3, 1006.7, 1007.1, 1007.6, 1008, 1008.3, 
    1008.8, 1009.1, 1009.4, 1009.7, 1009.8, 1010, 1010.3, 1010.1, 1010, 
    1009.7, 1009.6, 1009.4, 1009, 1008.7, 1008.6, 1008.4, 1008.3, 1008.1, 
    1007.8, 1007.6, 1007.3, 1006.8, 1006.4, 1005.8, 1005.4, 1005.2, 1005.1, 
    1004.8, 1004.8, 1004.5, 1004.6, 1004.4, 1004.3, 1004.2, 1004.2, 1004.2, 
    1004.2, 1004.2, 1004.3, 1004.2, 1004.1, 1004.1, 1004.1, 1004.2, 1004.1, 
    1004.3, 1004.4, 1004.5, 1004.6, 1004.8, 1004.8, 1004.8, 1005.4, 1005.7, 
    1006, 1005.8, 1006, 1006.5, 1006.5, 1006.5, 1006.5, 1006.8, 1006.8, 
    1006.7, 1007, 1007.3, 1007.6, 1007.6, 1007.6, 1007.6, 1007.5, 1007.5, 
    1007.3, 1007.3, 1007, 1006.9, 1006.7, 1006.6, 1006.1, 1005.9, 1005.6, 
    1005.3, 1005.1, 1004.9, 1004.6, 1004.3, 1004.1, 1004.1, 1004.2, 1004.1, 
    1004.1, 1004.1, 1004, 1003.9, 1003.8, 1003.6, 1003.2, 1002.9, 1002.6, 
    1002.2, 1001.6, 1001.4, 1000.9, 1000.3, 1000, 999.1, 998.3, 997.2, 996.4, 
    995.7, 995.1, 994.6, 993.9, 993.1, 992.5, 991.6, 990.8, 990.1, 989.3, 
    988.7, 987.9, 987.3, 986.8, 986.2, 985.7, 985.4, 984.9, 984.9, 984.9, 
    984.7, 984.7, 984.7, 984.6, 984.8, 985.3, 985.8, 986.4, 986.8, 987.4, 
    988, 988.4, 988.8, 988.8, 989.1, 989.4, 989.5, 989.9, 990.2, 990.6, 
    990.9, 990.9, 991.1, 991.3, 991.5, 991.8, 992, 992.2, 992.3, 992.4, 993, 
    993.4, 993.6, 994, 994.3, 994.6, 994.3, 994.1, 994, 994.1, 994, 993.9, 
    993.6, 993.4, 993.3, 992.9, 992.6, 992.2, 991.7, 991.3, 990.9, 990.7, 
    990.3, 990, 989.9, 989.8, 989.8, 989.7, 989.6, 989.4, 989.2, 988.9, 
    988.9, 988.7, 988.6, 988.7, 988.7, 988.6, 988.6, 988.6, 988.4, 988.3, 
    988.2, 988.1, 987.9, 987.6, 987.6, 987.6, 987.8, 988, 988.1, 988.2, 
    988.3, 988.4, 988.5, 988.6, 988.8, 989.1, 989.4, 989.7, 990.1, 990.5, 
    990.9, 991.3, 991.6, 992.2, 992.7, 993.2, 993.8, 994.4, 995.1, 995.5, 
    996.4, 997.2, 997.9, 998.7, 999.4, 1000, 1000.8, 1001.4, 1001.8, 1002.7, 
    1003.4, 1004.1, 1004.9, 1005.6, 1006.3, 1006.8, 1007, 1007.5, 1007.9, 
    1007.9, 1008.2, 1008.7, 1009.1, 1009.8, 1010.5, 1011.2, 1011.9, 1012.4, 
    1012.8, 1013.4, 1014, 1014.5, 1014.9, 1015.2, 1015.6, 1016, 1016.3, 
    1016.6, 1016.9, 1017, 1017, 1016.7, 1016.3, 1016.2, 1016.3, 1016.5, 
    1016.5, 1016.6, 1016.9, 1017.2, 1017.5, 1017.6, 1017.8, 1017.6, 1017.7, 
    1017.7, 1017.6, 1017.6, 1017.4, 1017, 1016.7, 1016.3, 1015.7, 1015.3, 
    1014.8, 1014.2, 1014.2, 1013.4, 1013.1, 1012.3, 1011.6, 1011.2, 1010.6, 
    1009.6, 1008.5, 1007.9, 1007.3, 1006.2, 1005.1, 1004, 1002.7, 1001.2, 
    1000.3, 999, 998, 997, 994.9, 994, 992, 991.4, 990.7, 990.5, 989.6, 989, 
    988.1, 987.6, 986.9, 986.3, 985.6, 985.3, 985.4, 986, 986.6, 987.3, 
    988.7, 989.3, 989.9, 990, 990.4, 991, 990.9, 991, 990.8, 990.9, 990.8, 
    990.5, 990.1, 990, 990, 990.1, 990.1, 990.1, 990.4, 990.6, 990.8, 991, 
    991, 991.1, 991.2, 991.4, 991.3, 991.4, 991.5, 991.5, 991.5, 991.5, 
    991.4, 991.6, 991.4, 991.7, 991.9, 992, 992.2, 992.6, 993.1, 994, 994.5, 
    995.1, 995.5, 995.9, 996.6, 997.2, 997.8, 998.5, 999, 999.6, 1000.2, 
    1000.6, 1001.1, 1001.5, 1001.9, 1002.2, 1002.5, 1002.6, 1002.8, 1003, 
    1003, 1003.2, 1003.3, 1003.5, 1003.5, 1003.4, 1003.3, 1003.3, 1003, 
    1002.6, 1002.4, 1002.1, 1001.6, 1001.4, 1001.1, 1000.8, 1000.4, 1000.3, 
    1000, 999.7, 999.2, 998.9, 998.6, 998.2, 998, 998, 998.2, 998.3, 998.2, 
    998.3, 998.3, 998.4, 998.6, 998.7, 998.9, 999.3, 999.6, 999.8, 1000.2, 
    1000.6, 1001.3, 1001.8, 1002.3, 1002.8, 1003.3, 1003.9, 1004.5, 1004.9, 
    1005.5, 1006.1, 1006.8, 1007.5, 1008.2, 1008.7, 1009.4, 1010.1, 1010.4, 
    1010.7, 1010.8, 1011.1, 1011.4, 1011.4, 1011.5, 1011.9, 1011.8, 1011.6, 
    1011.4, 1011.1, 1010.8, 1010.4, 1009.9, 1009.4, 1009.2, 1009.1, 1008.3, 
    1008, 1007.7, 1007.2, 1006.5, 1005.6, 1004.5, 1003.5, 1002.5, 1001.7, 
    1000.6, 999.7, 998.5, 997.5, 996.7, 995.9, 994.8, 994.1, 993, 991.7, 
    990.8, 990.7, 989.9, 989.3, 988.8, 988.3, 987.7, 987.1, 986.5, 986.4, 
    985.9, 985.1, 984.7, 983.9, 983.4, 982.9, 982.6, 982, 981.6, 981.3, 
    981.2, 980.8, 980.7, 980.6, 980.5, 980.5, 980.5, 981, 981.1, 981.5, 
    981.8, 982.4, 982.8, 983, 983.1, 983.4, 983.9, 984.3, 984.8, 985.1, 
    985.7, 986.6, 987, 987.5, 988.4, 989.4, 990.4, 991, 992.2, 993.3, 994.3, 
    995.3, 996.4, 998, 999.3, 1000.7, 1001.2, 1002, 1002.5, 1003.8, 1004.3, 
    1005.1, 1005.5, 1006.4, 1006.7, 1007.5, 1008, 1008.7, 1008.7, 1009.4, 
    1009.7, 1010.2, 1010.6, 1010.9, 1011.3, 1011.9, 1012.2, 1012.4, 1012.6, 
    1013, 1013.3, 1013.6, 1013.8, 1014.2, 1014.5, 1014.4, 1014.6, 1015.3, 
    1015.3, 1015.8, 1015.9, 1016.1, 1016.2, 1016.4, 1016.7, 1017, 1017.1, 
    1017.6, 1017.9, 1018.4, 1018.4, 1018.8, 1019.4, 1020, 1020.5, 1020.9, 
    1021.1, 1021.4, 1021.7, 1021.9, 1022.3, 1022.6, 1022.9, 1023.3, 1023.6, 
    1024, 1024.2, 1024.5, 1025, 1025.4, 1025.9, 1026.4, 1026.9, 1027.6, 
    1028.3, 1028.9, 1029.2, 1029.5, 1029.9, 1030.1, 1030.7, 1031, 1031, 
    1031.3, 1031.5, 1031.8, 1031.6, 1031.4, 1031.3, 1031.1, 1030.9, 1030.4, 
    1030.3, 1030.1, 1029.5, 1029.2, 1028.3, 1028.5, 1028.3, 1028.1, 1027.5, 
    1027, 1026.7, 1026.1, 1025.8, 1025.6, 1025, 1024.4, 1023.8, 1023.4, 
    1022.9, 1022.1, 1021.8, 1021.1, 1020.4, 1019.6, 1018.9, 1018.4, 1017.9, 
    1017.1, 1016.4, 1016, 1015.4, 1014.8, 1014.2, 1013, 1012.4, 1011.5, 
    1010.6, 1009.9, 1009.1, 1007.8, 1006.9, 1006.2, 1005.5, 1004.9, 1004.2, 
    1003, 1002.2, 1001.4, 1000.7, 1000.2, 999.9, 999.5, 999.5, 999.8, 1000.5, 
    1001.3, 1002.1, 1002.6, 1003.2, 1003.6, 1003.8, 1003.7, 1003.7, 1004, 
    1005, 1006.1, 1007.4, 1008.7, 1009.6, 1010.2, 1011.6, 1013, 1013.5, 
    1014.7, 1015.6, 1016.9, 1018.3, 1019.2, 1020.2, 1021.1, 1021.1, 1021, 
    1021.4, 1021.3, 1020.8, 1020.4, 1020, 1019.5, 1019.1, 1018.7, 1018.3, 
    1017.8, 1017.7, 1017.5, 1016.8, 1016.4, 1015.8, 1015, 1014.3, 1013.7, 
    1013.1, 1012.7, 1012.4, 1012.2, 1012, 1011.6, 1011.2, 1011.1, 1010.8, 
    1010.5, 1010.6, 1010.6, 1010.7, 1010.7, 1010.7, 1010.7, 1010.7, 1010.9, 
    1010.9, 1010.8, 1011.1, 1011.1, 1011.2, 1011.4, 1011.5, 1012, 1012.6, 
    1012.9, 1013.5, 1013.9, 1014.3, 1014.6, 1015, 1015.3, 1015.5, 1015.8, 
    1016, 1016.4, 1016.5, 1016.7, 1017.2, 1017.6, 1017.5, 1017.8, 1018.1, 
    1018.3, 1018.6, 1019, 1019.2, 1019.5, 1019.9, 1020.5, 1020.5, 1020.7, 
    1020.9, 1021.1, 1021.1, 1021.2, 1021.1, 1021.1, 1021.4, 1021.2, 1021.1, 
    1020.9, 1020.6, 1020.4, 1019.7, 1019.4, 1019.1, 1018.3, 1017.8, 1017.5, 
    1017.1, 1016.7, 1016.4, 1016.3, 1016.1, 1015.9, 1016, 1015.4, 1015.2, 
    1014.5, 1014.2, 1014.2, 1014.2, 1013.8, 1013.8, 1013.4, 1013, 1012.6, 
    1012.1, 1011.4, 1010.7, 1010, 1009.2, 1008.3, 1007.3, 1006.8, 1006.7, 
    1006.3, 1005.7, 1005.7, 1005.4, 1005.1, 1004.4, 1003.7, 1003.4, 1002.8, 
    1002, 1001.4, 1001.1, 1000.8, 1000.2, 1000, 999.4, 999, 998.5, 998.2, 
    998.2, 998.2, 998.7, 999.1, 999.5, 999.6, 1000.2, 1000.5, 1000.9, 1001.4, 
    1002.3, 1002.3, 1002.6, 1003.4, 1003.9, 1004.7, 1004.9, 1005.5, 1006, 
    1006.6, 1006.6, 1006.8, 1007.3, 1007.4, 1007.7, 1008, 1008.1, 1008.6, 
    1009.6, 1010.2, 1010.8, 1011.1, 1011.6, 1012.2, 1012.5, 1013.2, 1013.8, 
    1014.4, 1015.4, 1016, 1016.8, 1017.4, 1018.1, 1018.6, 1019.4, 1019.8, 
    1020.3, 1020.7, 1020.6, 1020.8, 1021, 1021.2, 1021.5, 1022.1, 1022.9, 
    1023.6, 1024.2, 1024.7, 1025.1, 1025.3, 1025.4, 1025.6, 1025.9, 1026.5, 
    1026.5, 1026.7, 1026.8, 1027.1, 1027.3, 1027.5, 1027.6, 1027.7, 1028, 
    1028, 1028.1, 1028.6, 1029, 1029.2, 1029.3, 1029.5, 1029.6, 1029.5, 
    1029.6, 1029.8, 1029.2, 1028.9, 1028.9, 1028.7, 1028.6, 1028.6, 1028.5, 
    1028, 1028.1, 1027.8, 1027.6, 1027.4, 1026.9, 1026.3, 1025.7, 1025.4, 
    1025.4, 1024.9, 1024.4, 1024, 1023.7, 1023.2, 1022.5, 1022, 1021.5, 
    1020.8, 1020.3, 1019.7, 1019.2, 1018.8, 1018, 1017.2, 1016.5, 1015.8, 
    1015.1, 1014, 1013.1, 1012.7, 1012.2, 1011.8, 1011.2, 1010.9, 1010.2, 
    1009.7, 1009, 1008.3, 1007.8, 1007.5, 1006.7, 1005.9, 1005.2, 1005, 1005, 
    1004.8, 1004.5, 1004.3, 1004.5, 1004.5, 1004.5, 1004.9, 1005.1, 1005.3, 
    1005, 1005.5, 1005.3, 1005.4, 1005.4, 1005.8, 1006, 1006.2, 1006.1, 
    1006.3, 1006.4, 1006.8, 1006.9, 1007, 1007, 1007.4, 1007.4, 1007.3, 
    1007.5, 1007.5, 1007.7, 1007.7, 1007.5, 1007.3, 1007.3, 1007.4, 1007.2, 
    1007, 1006.9, 1007.1, 1006.9, 1007.1, 1007, 1007.5, 1007.7, 1007.8, 
    1008.1, 1008.5, 1008.8, 1009, 1009.8, 1010, 1010.2, 1010.3, 1010.5, 
    1010.7, 1010.9, 1011.2, 1011.3, 1011.6, 1011.9, 1012.2, 1012.5, 1012.6, 
    1012.6, 1013, 1013.1, 1013.4, 1013.5, 1013.6, 1013.7, 1013.7, 1013.8, 
    1014, 1014.1, 1014.1, 1014.2, 1014.3, 1014.3, 1014.1, 1014, 1013.7, 
    1013.3, 1013.1, 1013, 1012.8, 1012.2, 1011.7, 1011.4, 1010.9, 1010.5, 
    1010.1, 1009.6, 1009.3, 1008.6, 1008.3, 1007.9, 1007.4, 1006.9, 1006.2, 
    1005.6, 1005.2, 1004.6, 1004.2, 1004.1, 1004, 1003.9, 1004.2, 1004.2, 
    1004.7, 1005, 1005.3, 1005.6, 1006.2, 1006.5, 1006.9, 1007.2, 1007.5, 
    1008, 1008.6, 1009.1, 1009.8, 1010.2, 1011.2, 1012, 1012.3, 1012.8, 
    1013.3, 1013.8, 1014.3, 1014.9, 1015.1, 1015.2, 1015.6, 1015.5, 1015.5, 
    1015.5, 1015.6, 1015.6, 1015.5, 1015.4, 1015.7, 1016, 1016.5, 1017.1, 
    1017.7, 1018.6, 1019.4, 1020.5, 1021.8, 1022.7, 1023.5, 1024.6, 1024.9, 
    1025.5, 1026.1, 1027.2, 1028.2, 1029.1, 1029.4, 1030.2, 1031.6, 1031.4, 
    1031.7, 1031.3, 1030.9, 1030, 1029.1, 1028.1, 1026.2, 1024.8, 1023.5, 
    1022.1, 1020.8, 1019.7, 1018.1, 1016.5, 1014.9, 1013.1, 1012.1, 1011.7, 
    1011.5, 1011.7, 1011.5, 1011, 1011, 1010.6, 1009.8, 1009, 1008.4, 1007.2, 
    1006.2, 1004.5, 1003, 1001.2, 999.5, 999, 997.9, 997, 995.8, 995, 995.1, 
    994.9, 996.3, 997, 997.8, 997.9, 998.1, 998.3, 998.7, 998.9, 1000.4, 
    1002, 1003.8, 1005.6, 1008, 1011.1, 1013.8, 1016.8, 1017.8, 1020.7, 
    1022.1, 1023.4, 1024.2, 1025.3, 1025.8, 1026.9, 1027.4, 1028, 1028.8, 
    1029.5, 1029.7, 1029.9, 1029.7, 1029.2, 1028.5, 1027.4, 1027.1, 1026.1, 
    1025, 1023.9, 1022.5, 1021.1, 1019.8, 1018.2, 1018, 1017.7, 1017.5, 
    1017.5, 1017.3, 1017.3, 1018.2, 1018.5, 1019.1, 1019.8, 1020.1, 1020.4, 
    1020.8, 1021, 1021.1, 1021.7, 1021.9, 1021.9, 1021.8, 1022.1, 1022, 
    1021.5, 1021.2, 1020.8, 1020.2, 1019.7, 1019.3, 1018.7, 1017.6, 1016.5, 
    1015.7, 1014.5, 1013.3, 1012.6, 1011.3, 1010, 1008.8, 1007.7, 1006.1, 
    1004.6, 1003.3, 1001.9, 1000.8, 999.8, 998.5, 997.3, 996.3, 995.3, 994.6, 
    994.2, 993.9, 994.2, 994.6, 995.5, 996.6, 997.7, 998.6, 999.9, 1000.7, 
    1001.6, 1002.3, 1003.3, 1004.5, 1005.2, 1006, 1006.3, 1007, 1007.7, 
    1008.4, 1009.1, 1009.3, 1009.8, 1010.3, 1010.5, 1010.6, 1011, 1010.8, 
    1011, 1011.1, 1011.2, 1011.5, 1011.8, 1012.3, 1012.5, 1012.9, 1013.1, 
    1013, 1013, 1013.2, 1013.5, 1014, 1014.1, 1014.5, 1014.6, 1014.6, 1014.7, 
    1014.8, 1015, 1015.1, 1015.2, 1015.3, 1015.5, 1015.8, 1016.2, 1016.3, 
    1016.6, 1016.7, 1016.7, 1016.8, 1016.9, 1016.9, 1017, 1016.8, 1017, 
    1017.1, 1017.3, 1017.4, 1017.6, 1017.4, 1017.5, 1017.6, 1017.8, 1017.9, 
    1017.6, 1017.6, 1017.7, 1017.6, 1017.9, 1018, 1018, 1018, 1017.9, 1017.7, 
    1017.4, 1017, 1016.5, 1016.1, 1015.6, 1015.2, 1014.6, 1014.1, 1013.3, 
    1012.5, 1011.3, 1010.4, 1009.7, 1008.7, 1007.4, 1006.1, 1004.8, 1003.9, 
    1002.6, 1001.8, 1000.6, 1000, 1000.2, 999.9, 999.6, 999.7, 999.3, 998.4, 
    998.2, 998, 997.8, 997.5, 997.1, 996.8, 996.5, 996.1, 995.8, 995.7, 
    995.8, 996.1, 996.5, 996.5, 996.9, 997.1, 997.3, 997.4, 996.9, 996.5, 
    996.1, 994.5, 992.5, 994, 996.4, 997.4, 997.4, 998.1, 999.4, 999.9, 
    999.8, 999.3, 999, 998.9, 999.6, 999.8, 1000.2, 1000.9, 1001.9, 1002.4, 
    1002.6, 1002.4, 1002, 1002.7, 1002.1, 1002.2, 1002.6, 1002.5, 1002.9, 
    1002.1, 1002.4, 1002.4, 1002.5, 1002.4, 1002.4, 1002.5, 1002.4, 1002.5, 
    1002.9, 1003, 1003.4, 1003.4, 1003.5, 1003.9, 1003.6, 1003.9, 1003.9, 
    1003.7, 1003.3, 1003.3, 1003.6, 1004.1, 1004.1, 1004.1, 1004.4, 1004.3, 
    1004.3, 1004.4, 1004.5, 1004.5, 1004.8, 1004.7, 1004.6, 1003.9, 1004.1, 
    1004, 1004, 1003.9, 1003.9, 1003.8, 1003.5, 1003.1, 1003.1, 1002.7, 
    1002.9, 1002.5, 1002.2, 1001.9, 1001.9, 1001.4, 1001.2, 1000.8, 1000.1, 
    999.6, 999, 998.6, 997.9, 997.5, 996.9, 996.7, 996.6, 996.9, 996.9, 997, 
    996.9, 996.7, 996.7, 996.6, 996.6, 996.2, 996.1, 996.2, 996.4, 996.3, 
    996.2, 996.5, 996.3, 996, 995.5, 995.5, 995.5, 995.1, 994.8, 994.6, 
    994.7, 994.7, 994.8, 994.4, 994.1, 993.9, 993.4, 993.2, 992.8, 992.7, 
    992.7, 992.8, 992.4, 992.2, 992.3, 992.1, 992.1, 991.9, 991.8, 991.7, 
    991.4, 991.6, 991.6, 991.7, 991.8, 991.9, 992, 992.1, 992, 992.4, 992.6, 
    992.8, 992.8, 992.8, 992.5, 993, 993, 992.9, 992.7, 992.5, 992.2, 992, 
    992.1, 991.9, 991.6, 991.3, 991.2, 991, 991, 991.1, 991.1, 991, 990.6, 
    990.5, 990.6, 990.5, 990.8, 990.9, 990.9, 990.9, 991.2, 991.6, 992, 
    992.2, 992.4, 992.6, 992.9, 993.2, 993.3, 993.5, 993.8, 994.1, 994.2, 
    994.7, 994.9, 995.1, 995.1, 995.2, 995.3, 995.3, 995.3, 995.2, 994.9, 
    994.7, 994.9, 994.9, 994.4, 993.6, 993.3, 992.9, 992.7, 992.8, 992.2, 
    992, 991.7, 991.6, 991.4, 991.3, 991.1, 990.7, 990.8, 990.9, 990.9, 
    990.9, 990.7, 990.9, 990.9, 991, 991, 991.3, 991.5, 991.4, 991.5, 991.8, 
    991.8, 992.1, 992.2, 992.4, 992.6, 992.9, 993.3, 993.4, 993.8, 994, 
    994.1, 994, 994.1, 994.2, 994.4, 994.6, 994.5, 994.5, 995, 995.7, 995.6, 
    996.1, 996.4, 996.6, 997.1, 997.2, 997.8, 998.2, 998.7, 999.2, 999.9, 
    1000.6, 1001.3, 1001.7, 1001.8, 1002.1, 1002.8, 1003.3, 1003.7, 1003.9, 
    1004.2, 1004.2, 1004.8, 1005.1, 1005.6, 1005.9, 1006.2, 1006.8, 1007.1, 
    1007.5, 1008, 1008.2, 1008.6, 1009, 1009.6, 1010, 1009.8, 1009.4, 1009, 
    1008.4, 1008.2, 1008, 1008.3, 1008.8, 1008.8, 1008.8, 1009.1, 1009.1, 
    1009.2, 1009.2, 1008.7, 1007.9, 1007.2, 1006.3, 1005.6, 1004.7, 1004.1, 
    1003, 1002.2, 1001.2, 1000.1, 999.1, 998.9, 999, 999.3, 1000.4, 1001.6, 
    1002.5, 1003, 1003.6, 1004.5, 1005.4, 1006, 1006.1, 1006.7, 1007.1, 
    1006.9, 1007.3, 1007, 1006.8, 1006.7, 1006.7, 1006.7, 1006.3, 1006, 
    1005.5, 1005.1, 1004.6, 1003.8, 1003.2, 1002.2, 1001.7, 1000.4, 999.5, 
    998.1, 996.5, 994.4, 991.5, 989.1, 987.4, 986.7, 986.7, 986.5, 986.4, 
    986.8, 987.7, 988.8, 989.5, 990.3, 990.7, 990.7, 990.9, 990.8, 990.5, 
    990, 989.4, 989.9, 990.6, 991.3, 992.4, 993, 993.8, 994.8, 996, 997.4, 
    999.1, 1000.1, 1000.7, 1001.6, 1002.6, 1003, 1003.8, 1004, 1004.3, 
    1004.2, 1004.1, 1003.9, 1003.5, 1003, 1002.2, 1001.4, 1000.7, 999.5, 
    998.4, 997.4, 996.4, 995.8, 994.9, 994.4, 994, 993.8, 993.6, 993.8, 
    994.1, 994, 994.2, 994.4, 994.3, 994.5, 994.4, 994.4, 994.4, 994.3, 
    994.2, 993.8, 993.3, 993.5, 994.4, 995.5, 997.1, 998.9, 999.4, 1000.2, 
    1001.4, 1002.3, 1003.4, 1004.1, 1005.3, 1006.2, 1006.8, 1007.6, 1007.9, 
    1008.4, 1008.5, 1008.6, 1008.7, 1008.7, 1008.6, 1008.7, 1009.1, 1009.9, 
    1010.2, 1010.3, 1010.8, 1011.4, 1011.8, 1012, 1012.6, 1013.3, 1014.2, 
    1014.7, 1015.6, 1016.2, 1017.2, 1018, 1018.9, 1019.5, 1020.3, 1020.8, 
    1021, 1021.5, 1022.8, 1023.4, 1023.8, 1024.4, 1024.7, 1025.1, 1025.4, 
    1025.5, 1025.8, 1025.8, 1025.8, 1025.6, 1025.4, 1025.3, 1025, 1024.6, 
    1024.5, 1024.1, 1023.3, 1022.2, 1020.8, 1020.1, 1019.9, 1019.3, 1018.7, 
    1018.3, 1018.2, 1018.2, 1017.7, 1017, 1016.6, 1016.1, 1015.1, 1014.6, 
    1014.3, 1014.2, 1013.9, 1014.1, 1014, 1013.8, 1013.7, 1013.6, 1013.3, 
    1013.3, 1013.1, 1013.4, 1013.9, 1014.2, 1014.5, 1014.6, 1014.5, 1014.9, 
    1015.2, 1015.5, 1015.6, 1015.8, 1015.8, 1015.5, 1015.3, 1015.1, 1014.9, 
    1014.9, 1015, 1014.7, 1014.4, 1014.1, 1013.7, 1013.5, 1013.1, 1012.9, 
    1012.5, 1012.5, 1012.4, 1012, 1012, 1011.9, 1011.6, 1011.5, 1011.1, 
    1010.5, 1010.2, 1010, 1009.8, 1009.5, 1008.9, 1008.6, 1008.4, 1008.2, 
    1007.9, 1007.8, 1007.3, 1007, 1006.7, 1006.2, 1005.7, 1005.1, 1004.5, 
    1003.7, 1003.1, 1002.5, 1001.8, 1001, 1000.2, 999.3, 998.5, 997.5, 996.2, 
    994.3, 992.7, 991.4, 990, 988.9, 988.2, 987, 985.9, 985.1, 984.6, 983.8, 
    983.3, 983.4, 983, 983.5, 984.4, 985.4, 986.9, 988, 989.1, 990.1, 991.3, 
    992.4, 993.2, 994.1, 995, 996, 996.6, 997.4, 998.7, 999.3, 999.9, 1000.1, 
    1000.3, 1000.7, 1001.4, 1001.9, 1002.6, 1003.3, 1003.5, 1004.1, 1004.3, 
    1004.9, 1005.1, 1005.4, 1005.3, 1005.1, 1005.1, 1004.7, 1004, 1003.2, 
    1002.8, 1002.5, 1002, 1001.2, 1000.3, 999.9, 999.3, 998.7, 998.4, 998.1, 
    997.9, 997.6, 997.6, 997.4, 997.5, 997.4, 997.4, 997.6, 997.8, 998, 
    998.3, 998.6, 998.8, 998.8, 999.3, 999.7, 1000, 1000.3, 1000.4, 1000.6, 
    1000.9, 1000.6, 1000.5, 1000.4, 1000.6, 1000.5, 1000.3, 1000.1, 1000.1, 
    1000.1, 1000.1, 999.9, 999.9, 1000.1, 1000.2, 1000.1, 1000.2, 1000.4, 
    1000.9, 1001.2, 1001.3, 1001.4, 1001.3, 1001.9, 1002.1, 1002.3, 1002.3, 
    1002.4, 1002.5, 1002.5, 1002.6, 1003, 1003.5, 1003.7, 1003.7, 1004, 1004, 
    1004.5, 1004.5, 1004.7, 1004.8, 1004.9, 1005.2, 1005.3, 1005.7, 1005.7, 
    1006, 1006, 1006.3, 1006.2, 1006.4, 1006.5, 1006.6, 1006.5, 1006.5, 
    1006.2, 1005.8, 1005.3, 1005.2, 1004.2, 1003.9, 1003.5, 1003.2, 1003.1, 
    1003, 1003, 1003.2, 1003.3, 1004, 1004.2, 1004.2, 1003.9, 1003.2, 1002.5, 
    1001.6, 1000.9, 999.9, 998.9, 998.1, 997.7, 996.8, 995.8, 994.9, 994.1, 
    993.3, 993.2, 993.3, 993.3, 993.8, 994.3, 995.1, 995.9, 996.5, 997.3, 
    997.9, 998.3, 998.6, 999.1, 999.5, 999.7, 999.8, 999.8, 1000.3, 1001.1, 
    1001.8, 1002.5, 1003.2, 1003.9, 1004.7, 1005.4, 1005.9, 1006.5, 1006.5, 
    1006.7, 1006.8, 1007, 1007.2, 1007.3, 1007.4, 1007.3, 1007.2, 1007.1, 
    1007, 1007, 1006.9, 1006.8, 1006.8, 1007.1, 1007.5, 1007.8, 1007.9, 
    1008.3, 1008.5, 1008.6, 1008.6, 1008.3, 1008.1, 1008, 1008.2, 1008.3, 
    1008, 1008, 1007.6, 1007.5, 1007.2, 1006.8, 1006.4, 1005.5, 1004.9, 
    1004.4, 1004, 1003.6, 1003.5, 1003.7, 1003.9, 1004.3, 1004.6, 1005.1, 
    1005.4, 1005.8, 1006.2, 1006.8, 1007.2, 1008, 1008.7, 1009.3, 1009.8, 
    1010.2, 1010.7, 1011, 1011.6, 1012, 1012.6, 1013, 1013.4, 1013.8, 1014.4, 
    1015, 1015.5, 1015.9, 1016.5, 1016.9, 1017.1, 1017.1, 1017.7, 1017.6, 
    1017.8, 1018.2, 1018.1, 1018.1, 1018.1, 1017.8, 1017.6, 1017.5, 1016.9, 
    1016.2, 1015.7, 1015, 1013.9, 1012.7, 1011.5, 1010.2, 1009.1, 1008.2, 
    1007.3, 1006.6, 1005.8, 1005.2, 1004.6, 1004.1, 1003.6, 1003.6, 1003.4, 
    1003.6, 1003.8, 1004, 1004.2, 1004.8, 1005.2, 1005.6, 1006.3, 1006.6, 
    1006.9, 1007.3, 1007.4, 1007.5, 1007.9, 1008.5, 1008.6, 1008.7, 1008.9, 
    1008.7, 1008.8, 1009, 1009.2, 1009.6, 1009.9, 1009.7, 1009.8, 1009.6, 
    1009.7, 1009.5, 1009.2, 1008.7, 1008.2, 1007.9, 1007.7, 1007.5, 1007.2, 
    1006.9, 1006.8, 1007, 1007, 1006.8, 1006.7, 1006.8, 1006.9, 1006.5, 
    1006.1, 1005.9, 1005.3, 1005.2, 1005.2, 1004.8, 1003.8, 1002.8, 1002.9, 
    1002.6, 1001.8, 1001, 1000.3, 1000, 999.8, 1000, 999.3, 999.2, 998.5, 
    998.5, 998.3, 998.5, 998.1, 997.9, 997.9, 997.6, 997.6, 997.6, 997.1, 
    996.8, 996.9, 997.5, 997, 997.1, 997.2, 997.4, 997.4, 997.3, 997.3, 
    997.5, 998, 998.3, 998.4, 998.3, 998.2, 998.8, 998.9, 999.6, 1000.4, 
    1000.7, 1000.9, 1000.9, 1000.8, 1000.8, 1001, 1001.7, 1001.4, 1001.5, 
    1002.4, 1003.2, 1004, 1005, 1005.9, 1006.6, 1007.5, 1008.4, 1009.1, 
    1009.6, 1010.3, 1010.5, 1010.7, 1011.1, 1011.7, 1012.3, 1012.7, 1012.9, 
    1013, 1013.1, 1013.1, 1013.2, 1013, 1012.6, 1012.4, 1012, 1011.2, 1010.8, 
    1010.2, 1009.5, 1008.8, 1008, 1007.5, 1006.7, 1005.7, 1005, 1004, 1003, 
    1002.3, 1001.9, 1001.7, 1001.7, 1001.3, 1000.9, 1000.9, 1001, 1000.8, 
    1000.4, 999.6, 999, 998.6, 997.7, 997.4, 996.1, 994.7, 993.3, 992.2, 
    990.4, 988.7, 987.1, 985.2, 984.8, 983.6, 983, 982.2, 982, 981.5, 980.6, 
    980.6, 981.3, 982.7, 983.7, 984.9, 986.3, 987.4, 988.9, 990.1, 990.5, 
    992.6, 993.3, 995.3, 996.7, 998.1, 997.7, 998.8, 999.7, 1000.3, 1000.5, 
    1000.4, 1001.1, 1001.2, 1001.3, 1001.3, 1001.5, 1002, 1002.1, 1001.9, 
    1002.2, 1002.4, 1002.5, 1002.9, 1002.9, 1002.8, 1002.7, 1002.7, 1002.6, 
    1002, 1001.7, 1001.7, 1001.7, 1001.7, 1001.4, 1001.1, 1000.9, 1000.6, 
    1000.4, 1000.1, 999.9, 999.5, 999.2, 998.7, 998.4, 997.9, 997.6, 997.1, 
    996.9, 996.4, 995.9, 995.6, 995.4, 994.9, 994.8, 994.5, 994.1, 993.6, 
    993.1, 992.8, 992.8, 992.6, 992.5, 992.8, 993.1, 993.5, 993.9, 994.2, 
    994.1, 994.2, 994.7, 995.1, 995.6, 996, 996, 996.4, 996.8, 997.2, 997.4, 
    997.7, 997.8, 998.2, 998.8, 999.1, 999.5, 999.8, 1000, 1000.4, 1000.8, 
    1001, 1001.3, 1001.5, 1001.6, 1001.8, 1002.1, 1002.4, 1002.9, 1002.8, 
    1002.7, 1002.5, 1002.4, 1002.4, 1002.7, 1002.6, 1002.5, 1002.6, 1002.7, 
    1002.7, 1002.8, 1002.9, 1002.9, 1002.9, 1002.9, 1003.1, 1003.1, 1003, 
    1003, 1002.8, 1002.8, 1002.8, 1002.9, 1002.9, 1002.9, 1002.8, 1002.6, 
    1002.7, 1002.8, 1002.5, 1002.5, 1002.6, 1002.5, 1002.5, 1002.7, 1002.6, 
    1002.3, 1002.3, 1002.1, 1001.9, 1001.8, 1001.8, 1001.7, 1001.8, 1001.8, 
    1001.8, 1001.9, 1001.9, 1001.7, 1001.6, 1001.7, 1001.7, 1001.7, 1001.9, 
    1001.9, 1001.8, 1002, 1002.2, 1002.4, 1002.2, 1001.9, 1001.8, 1001.7, 
    1001.7, 1001.8, 1002, 1001.9, 1001.7, 1001.6, 1001.6, 1001.6, 1001.4, 
    1001.2, 1000.8, 1000.6, 1000.5, 1000.3, 1000.1, 999.9, 999.7, 999.7, 
    999.8, 999.9, 999.9, 999.9, 999.8, 999.8, 999.6, 999.6, 999.5, 999.6, 
    999.5, 999.5, 999.5, 999.9, 1000.2, 1000.3, 1000.5, 1000.3, 1000.4, 
    1000.4, 1000.7, 1001.1, 1001.5, 1001.8, 1002.2, 1002.3, 1002.6, 1003.2, 
    1003.5, 1003.9, 1004.3, 1004.6, 1005.1, 1005.4, 1005.8, 1006.2, 1006.8, 
    1007.2, 1007.8, 1008.2, 1008.6, 1008.8, 1009.4, 1009.7, 1010.1, 1010.4, 
    1010.8, 1011.4, 1011.8, 1012.5, 1012.8, 1013, 1013.1, 1013.5, 1013.8, 
    1014.1, 1014.3, 1014.5, 1014.7, 1014.9, 1015.3, 1015.6, 1015.8, 1016.1, 
    1016.4, 1016.4, 1016.7, 1016.8, 1016.8, 1017, 1017.4, 1017.7, 1018.1, 
    1018.4, 1018.6, 1019, 1018.9, 1019, 1019.2, 1019.4, 1019.6, 1019.8, 1020, 
    1019.9, 1019.9, 1020.4, 1020.5, 1020.5, 1020.6, 1020.8, 1021, 1021.2, 
    1021.3, 1021.5, 1022, 1022.4, 1022.6, 1023.1, 1023.2, 1023.5, 1023.6, 
    1023.9, 1024.1, 1024.3, 1024.5, 1024.8, 1025.1, 1025.4, 1025.7, 1026.2, 
    1026.4, 1026.5, 1026.5, 1026.8, 1027, 1027.1, 1027.2, 1027.4, 1027.7, 
    1027.9, 1028.1, 1028.2, 1028.4, 1028.5, 1028.5, 1028.5, 1028.9, 1028.9, 
    1028.8, 1029, 1029, 1029.2, 1029.3, 1029.4, 1029.4, 1029.4, 1029.4, 
    1029.2, 1029.1, 1029.1, 1028.9, 1028.6, 1028.8, 1028.8, 1028.6, 1028.2, 
    1028.1, 1027.7, 1027.6, 1027.6, 1027.2, 1027.4, 1027.1, 1027.1, 1026.7, 
    1026.5, 1026.3, 1026.2, 1025.9, 1025.5, 1025.4, 1025.3, 1025.2, 1024.9, 
    1024.6, 1024.4, 1024.6, 1024.6, 1024.6, 1024.6, 1024.5, 1024.4, 1024.2, 
    1024.3, 1024.3, 1024.2, 1024.1, 1024.1, 1024, 1024, 1023.9, 1023.8, 
    1023.7, 1023.3, 1023, 1022.9, 1022.5, 1022, 1021.8, 1021.4, 1021.2, 
    1020.8, 1020.4, 1019.8, 1019.5, 1018.9, 1018.4, 1018.1, 1017.6, 1017.4, 
    1016.7, 1016.4, 1015.9, 1015.5, 1015.2, 1014.9, 1014.5, 1014.2, 1013.6, 
    1013.2, 1012.8, 1012.4, 1011.9, 1011.6, 1011.3, 1011.3, 1011.3, 1011.6, 
    1011.5, 1011.5, 1011.8, 1011.8, 1012, 1012, 1011.9, 1011.8, 1011.9, 1012, 
    1012.3, 1012.4, 1012.6, 1012.8, 1013, 1013.5, 1013.5, 1013.7, 1014.1, 
    1014.2, 1014.3, 1014.5, 1014.7, 1015, 1015, 1014.6, 1014.9, 1015, 1015, 
    1014.9, 1014.9, 1015.1, 1015.2, 1015.3, 1015.3, 1015.3, 1015.2, 1015.2, 
    1015, 1015, 1015, 1014.8, 1015, 1014.4, 1014.4, 1014.2, 1014.3, 1014.2, 
    1014, 1014, 1013.6, 1013.1, 1013.3, 1013, 1012.9, 1012.7, 1012.5, 1012.3, 
    1012.4, 1012.3, 1012.4, 1012.3, 1012, 1011.8, 1011.5, 1011.2, 1010.9, 
    1010.7, 1010.5, 1010.2, 1010, 1009.9, 1009.5, 1009.1, 1008.7, 1008.2, 
    1007.9, 1007.7, 1006.9, 1006.6, 1006.5, 1006.7, 1007.2, 1007.9, 1008.5, 
    1009, 1009.4, 1009.9, 1010.5, 1010.9, 1011.6, 1012, 1012.6, 1013.1, 
    1013.8, 1014.5, 1015.4, 1015.9, 1016.5, 1017.2, 1017.7, 1018.2, 1018.9, 
    1019.5, 1020.2, 1021, 1021.9, 1022.5, 1023.2, 1023.5, 1023.8, 1024.1, 
    1024.3, 1024.7, 1025.1, 1025.6, 1026, 1026.4, 1026.9, 1027.2, 1027.6, 
    1027.9, 1027.9, 1028, 1028.1, 1028.4, 1028.5, 1028.7, 1029, 1029.1, 
    1029.4, 1029.7, 1029.7, 1029.7, 1029.6, 1029.4, 1029.3, 1029.3, 1029.1, 
    1029, 1029, 1028.9, 1028.8, 1028.7, 1028.6, 1028.4, 1027.8, 1027.3, 
    1026.8, 1026.6, 1026.3, 1025.9, 1025.4, 1025.1, 1024.6, 1024.4, 1024.2, 
    1024, 1024, 1023.9, 1023.7, 1023.4, 1023.3, 1023.2, 1023.3, 1023.6, 
    1023.7, 1023.9, 1024.1, 1024.1, 1023.9, 1023.7, 1023.4, 1023.3, 1023.4, 
    1023.4, 1023.4, 1023.3, 1023.4, 1023.3, 1023.2, 1023.1, 1022.9, 1022.7, 
    1022.4, 1022.2, 1022.2, 1022.1, 1022.1, 1022.2, 1022.1, 1022.1, 1022.2, 
    1022, 1021.7, 1021.5, 1021.2, 1021.1, 1020.9, 1020.9, 1021, 1021.1, 
    1021.3, 1021.2, 1021.2, 1021.3, 1021.2, 1021.4, 1021.3, 1021.2, 1021.3, 
    1021.2, 1021.4, 1021.4, 1021.7, 1021.8, 1021.9, 1022.1, 1022.1, 1021.9, 
    1021.9, 1021.9, 1021.9, 1021.9, 1022, 1022.2, 1022.2, 1022.2, 1022.3, 
    1022.2, 1021.9, 1021.5, 1021.3, 1020.8, 1020.4, 1020.1, 1019.9, 1020.1, 
    1019.8, 1019.6, 1019.1, 1018.9, 1018.3, 1017.8, 1017.2, 1016.6, 1016.1, 
    1015.5, 1014.9, 1014.6, 1014.1, 1013.6, 1013.1, 1012.5, 1011.8, 1011.6, 
    1011.3, 1011, 1010.5, 1010.2, 1010.1, 1010, 1009.8, 1009.6, 1009.5, 
    1009.5, 1009.5, 1009.2, 1008.7, 1008.6, 1008.4, 1008.1, 1008, 1008, 
    1008.1, 1008.1, 1008.1, 1008.3, 1008.3, 1008.4, 1008.1, 1008, 1008.3, 
    1008.3, 1008.6, 1008.7, 1008.6, 1008.7, 1008.6, 1008.4, 1008.3, 1008.4, 
    1008.4, 1008.3, 1008, 1007.8, 1007.9, 1007.8, 1007.6, 1007.4, 1007.1, 
    1006.9, 1006.4, 1006.1, 1006.1, 1005.6, 1005.6, 1005.6, 1005.4, 1005.4, 
    1005.5, 1005.4, 1005.2, 1005, 1004.9, 1004.7, 1004.4, 1004.3, 1004.1, 
    1004.1, 1003.9, 1003.7, 1003.5, 1003.3, 1003.1, 1002.9, 1002.7, 1002.4, 
    1002.1, 1001.8, 1001.8, 1001.9, 1001.9, 1002, 1002.1, 1001.9, 1002, 
    1002.1, 1001.9, 1001.8, 1001.6, 1001.5, 1001.5, 1001.4, 1001.4, 1001.3, 
    1001.3, 1001.5, 1001.4, 1001.3, 1001.6, 1001.7, 1001.7, 1001.8, 1002.1, 
    1002.2, 1002.4, 1002.8, 1003.1, 1003.2, 1003.3, 1003.7, 1004.1, 1004.4, 
    1004.5, 1004.6, 1004.9, 1005, 1005, 1005.5, 1005.5, 1005.9, 1006.1, 
    1005.9, 1006.1, 1006.3, 1006.4, 1006.6, 1006.8, 1006.9, 1006.9, 1007.3, 
    1007.3, 1007.6, 1007.7, 1007.8, 1007.9, 1007.7, 1007.6, 1007.3, 1007, 
    1006.9, 1006.8, 1006.5, 1006.2, 1006, 1005.7, 1005.5, 1005.2, 1005, 
    1004.8, 1004.5, 1004.4, 1004.4, 1004.3, 1004.6, 1004.7, 1004.7, 1004.9, 
    1004.9, 1004.9, 1004.6, 1004.8, 1004.8, 1004.5, 1004.2, 1004.1, 1003.8, 
    1003.7, 1003.5, 1003.1, 1002.7, 1002.3, 1002, 1001.5, 1000.8, 999.9, 
    999.1, 998.4, 998, 997.4, 997, 996.3, 995.7, 995.2, 994.8, 994.5, 994.3, 
    994.3, 994.1, 994.2, 994.3, 994.6, 995.1, 995.5, 996, 996.4, 996.7, 
    997.6, 998.1, 998.7, 999.1, 999.6, 1000.4, 1000.9, 1001.3, 1001.9, 
    1002.3, 1002.6, 1003, 1003.4, 1003.4, 1003.7, 1004, 1004.1, 1004.3, 
    1004.5, 1004.9, 1004.9, 1004.8, 1004.4, 1004.3, 1004.1, 1003.9, 1003.9, 
    1003.8, 1003.9, 1004, 1004.3, 1004.6, 1004.8, 1005.1, 1005.3, 1005.7, 
    1006.2, 1006.9, 1007.6, 1008.2, 1009, 1009.7, 1010.3, 1010.8, 1011.3, 
    1011.6, 1012.1, 1012.6, 1013.2, 1013.8, 1014, 1014.5, 1014.8, 1015.7, 
    1016.1, 1016.7, 1017.1, 1017.6, 1017.9, 1018.1, 1018.2, 1018.4, 1018.4, 
    1018.2, 1018.1, 1018.1, 1018, 1018.2, 1018.2, 1017.8, 1017.6, 1017.3, 
    1016.8, 1016.6, 1016.3, 1016.4, 1016.1, 1015.7, 1015.6, 1015.3, 1015, 
    1014.7, 1014.2, 1013.8, 1013.4, 1012.8, 1012.6, 1012.4, 1012.1, 1012.1, 
    1011.6, 1011.3, 1011, 1010.6, 1010.4, 1009.8, 1009.4, 1008.8, 1008.3, 
    1007.9, 1007.5, 1007.3, 1007.2, 1007.1, 1006.7, 1006.6, 1006.3, 1006.2, 
    1006.1, 1005.9, 1005.8, 1006.1, 1006.2, 1006.2, 1006.4, 1006.7, 1006.7, 
    1006.5, 1006.5, 1006.6, 1006.7, 1006.8, 1006.9, 1007, 1007.2, 1007.3, 
    1007.5, 1007.8, 1007.5, 1007.3, 1007.2, 1006.4, 1006, 1005.3, 1004.7, 
    1004.2, 1003.8, 1003.3, 1003.3, 1003.4, 1003.6, 1003.7, 1003.9, 1004.3, 
    1004.8, 1005.1, 1005.6, 1006.2, 1006.4, 1006.7, 1007, 1006.9, 1006.8, 
    1007.2, 1007, 1006.4, 1005.6, 1004.6, 1003.5, 1001.7, 1000.2, 999.2, 
    998.4, 997.7, 997.4, 996.5, 996, 995.7, 995, 994.6, 993.3, 992, 990.8, 
    989.3, 987.6, 986, 984.5, 983, 982.1, 981.3, 981, 980.9, 980.7, 980.7, 
    980.7, 981, 981.2, 981.6, 982.2, 982.7, 983.3, 984, 985, 985.9, 986.6, 
    987.8, 989.1, 990, 991.1, 992.2, 993, 994, 994.7, 995.2, 995.8, 996.5, 
    996.5, 996.8, 997.2, 997.1, 997.4, 997.2, 997.1, 996.3, 995.6, 995.2, 
    994.7, 993.9, 992.9, 992.9, 992.5, 992.5, 992.6, 993, 993.8, 994.5, 
    995.5, 996.4, 997.4, 999.2, 1000.4, 1001.6, 1003.2, 1005.2, 1007, 1008.1, 
    1009.2, 1010.4, 1011.4, 1012.4, 1013.1, 1013.9, 1014.1, 1014.4, 1015, 
    1015.4, 1015.7, 1016.2, 1016.1, 1016.2, 1016.2, 1016.2, 1015.6, 1015.4, 
    1015.2, 1015, 1015.2, 1015.2, 1015.6, 1015.5, 1015.4, 1015.5, 1015.5, 
    1015.1, 1014.8, 1014.1, 1013.6, 1013.6, 1013.4, 1013.5, 1013.7, 1013.5, 
    1013.1, 1011.7, 1011, 1010.5, 1009.8, 1009, 1007.7, 1006.7, 1006.2, 
    1006.2, 1006.1, 1006, 1005.7, 1005.6, 1005.8, 1005.8, 1005.8, 1006.1, 
    1006.4, 1006.5, 1007.4, 1007.9, 1008.2, 1008.8, 1009.3, 1009.6, 1009.9, 
    1010.3, 1010.5, 1010.5, 1010.1, 1009.9, 1009.9, 1009.8, 1009.5, 1009.6, 
    1009.3, 1009.3, 1009.1, 1009, 1009, 1008.4, 1008.2, 1008.6, 1008.5, 
    1008.7, 1008.9, 1009.4, 1009.4, 1010.1, 1010.6, 1010.6, 1011.1, 1010.9, 
    1010.9, 1011.3, 1011.6, 1011.4, 1011.8, 1011.4, 1011.9, 1012.3, 1012.2, 
    1012.4, 1012.5, 1012.5, 1012.2, 1012.6, 1012.6, 1012.3, 1012.1, 1012.5, 
    1012.3, 1011.9, 1011.6, 1011.1, 1010.6, 1010, 1009.8, 1009.1, 1008.6, 
    1007.7, 1007.1, 1006.5, 1005.7, 1004.6, 1003.4, 1002.4, 1001.9, 1001.8, 
    1001.6, 1001.1, 1000.9, 1000.9, 1000.7, 1001, 1000.8, 1001, 1001.1, 
    1000.4, 1000.3, 1000.2, 1000.2, 999.8, 999.5, 999.3, 999.1, 998.9, 998.9, 
    998.7, 998.7, 998.7, 998.6, 998.6, 998.5, 999.3, 999.5, 999.8, 1000.5, 
    1000.3, 1000.9, 1000.8, 1000.9, 1000.3, 1001.1, 1001.1, 1001.2, 1001.6, 
    1001.7, 1001.7, 1001.9, 1002.3, 1002.4, 1002.3, 1001.5, 1001.6, 1001, 
    1000.8, 1000.2, 999.2, 998.9, 998.4, 997.7, 997.6, 996.9, 996.9, 996.5, 
    996.2, 996.1, 995.8, 995.5, 995.3, 994.9, 994.7, 994.2, 993.8, 993.3, 
    993, 992.7, 992.2, 991.8, 991.9, 991.8, 992, 992.2, 992.4, 992.4, 992.8, 
    993.3, 993.5, 993.4, 993, 993.5, 993.2, 993.3, 993.2, 992.9, 993.3, 
    993.8, 994.5, 995, 995.1, 995.2, 995.5, 995.5, 995.6, 995.6, 996.1, 
    996.2, 996.9, 998.1, 998.7, 1000, 1001.2, 1001.8, 1002.3, 1003.1, 1004.2, 
    1004.6, 1004.6, 1005.1, 1005.5, 1005.7, 1005.6, 1005.7, 1006.2, 1006.6, 
    1006.3, 1007, 1007.3, 1007.3, 1006.9, 1007.4, 1007.5, 1007.7, 1007.8, 
    1007.8, 1008, 1008, 1008.1, 1008.3, 1008.5, 1008.6, 1008.6, 1008.6, 
    1008.7, 1008.6, 1008.7, 1008.8, 1008.7, 1008.9, 1008.8, 1008.7, 1008.5, 
    1008.5, 1008.5, 1008.7, 1008.7, 1009.1, 1009.2, 1009.3, 1009.3, 1009.3, 
    1009.3, 1008.8, 1008.7, 1008.5, 1008.4, 1008, 1007.9, 1007.6, 1007.2, 
    1007, 1006.8, 1006.4, 1006.2, 1005.9, 1005.2, 1004.8, 1004.6, 1004.4, 
    1004, 1004, 1003.4, 1003.4, 1002.9, 1002.6, 1002, 1001.4, 1001.1, 1000.6, 
    1000.2, 1000.2, 1000.2, 999.9, 999.7, 999.8, 999.6, 999.5, 999.6, 999.4, 
    999.3, 999.4, 999.6, 999.6, 999.8, 999.9, 1000.1, 1000.2, 1000.3, 1000.5, 
    1000.6, 1000.7, 1000.9, 1001.1, 1001.1, 1001.4, 1001.8, 1002.1, 1002.5, 
    1002.7, 1002.9, 1003.2, 1003.5, 1003.9, 1004.1, 1004.4, 1004.4, 1004.8, 
    1005.1, 1005.4, 1005.6, 1005.9, 1005.9, 1005.8, 1005.8, 1005.8, 1005.9, 
    1006, 1005.8, 1005.8, 1005.8, 1005.7, 1005.6, 1005.7, 1005.6, 1005.5, 
    1005.1, 1005, 1004.7, 1004.6, 1004.5, 1004.3, 1004.2, 1004, 1004.2, 
    1003.9, 1003.5, 1003.6, 1003.5, 1003.2, 1003.1, 1003.2, 1003.2, 1003.2, 
    1003.6, 1003.5, 1003.5, 1003.3, 1003.4, 1003.2, 1003.1, 1003.2, 1003.1, 
    1003, 1002.9, 1003, 1003.2, 1003.4, 1003.4, 1003.4, 1003.1, 1003, 1002.8, 
    1002.7, 1002.3, 1002.1, 1001.8, 1001.8, 1001.4, 1001.3, 1001.2, 1001.1, 
    1000.8, 1000.5, 1000.5, 1000.2, 1000, 1000, 999.8, 999.8, 999.8, 1000, 
    1000, 999.8, 999.7, 999.4, 999.3, 999.1, 999.1, 999, 998.7, 998.8, 998.6, 
    998.8, 999, 998.9, 998.9, 999, 999.2, 999.1, 998.7, 998.9, 999.3, 999.5, 
    999.8, 999.9, 1000.2, 1000.4, 1000.4, 1000.7, 1000.8, 1001.1, 1001.3, 
    1001.6, 1001.9, 1002.2, 1002.7, 1002.9, 1003.2, 1003.4, 1003.6, 1003.8, 
    1004.3, 1004.3, 1004.3, 1004.3, 1004.5, 1004.7, 1004.8, 1004.9, 1005, 
    1005.2, 1005.3, 1005.3, 1005.4, 1005.4, 1005.6, 1005.7, 1005.8, 1006, 
    1006.2, 1005.8, 1005.7, 1005.7, 1005.7, 1005.8, 1005.5, 1005.5, 1005.2, 
    1005.1, 1004.8, 1004.9, 1004.9, 1004.6, 1004.9, 1004.9, 1004.2, 1004.5, 
    1004.6, 1004.8, 1004.6, 1004.6, 1004.3, 1004.2, 1004.3, 1004.5, 1004.4, 
    1004.4, 1004.5, 1004.2, 1003.6, 1003.2, 1002.6, 1001.9, 1000.2, 999, 
    997.9, 996.7, 995.8, 994.1, 992.2, 991.4, 989.7, 990.2, 991.1, 992, 
    992.6, 994.6, 996.7, 998.6, 1000, 1000.6, 1001.1, 1002.5, 1003, 1003.6, 
    1003.9, 1004.2, 1004.9, 1005.7, 1006.2, 1006.5, 1007.2, 1007.2, 1007, 
    1006.4, 1006, 1005.4, 1004.4, 1003.7, 1003, 1002.7, 1001.4, 1000.5, 
    998.8, 996.9, 995.6, 994.3, 992.9, 991.6, 990.1, 988.9, 987.5, 986.7, 
    985.8, 985.7, 985.4, 985.6, 985.8, 986.3, 987, 987.8, 988.6, 989.4, 
    989.9, 990.4, 990.8, 991.5, 992, 992.2, 992, 992.1, 991.8, 991.6, 991.5, 
    990.9, 990.6, 990.2, 990.2, 990, 989.5, 989.1, 988.6, 988.4, 988.3, 988, 
    987.5, 987, 986.5, 986.3, 985.8, 985.3, 984.5, 983.9, 983.6, 982.7, 982, 
    980.9, 979.8, 979.6, 979.1, 978.9, 978.7, 978.6, 978.7, 978.9, 978.9, 
    979.2, 979.7, 980.2, 980.9, 981.5, 981.5, 982, 982.2, 982.6, 982.5, 
    982.3, 982, 981.6, 980.9, 980.8, 980.4, 980, 979.8, 979.2, 979.1, 979.2, 
    979.2, 978.9, 978.9, 979, 979.2, 979.7, 980, 980.7, 980.9, 981.2, 981.6, 
    982.3, 982.9, 983.5, 984.2, 984.8, 985.5, 986.3, 986.9, 987.5, 988.2, 
    988.9, 989.8, 990.2, 991.1, 991.6, 991.8, 992.3, 992.4, 992.6, 993.2, 
    993.4, 993.8, 993.4, 993.2, 993.6, 993.9, 993.8, 993.3, 992.9, 992.8, 
    992.6, 993.1, 994.5, 995.2, 995.9, 996.3, 997.8, 998.6, 999.1, 1000.2, 
    1001.1, 1001.4, 1002, 1002.7, 1003.4, 1004, 1004.7, 1005.9, 1006.2, 
    1006.9, 1007.2, 1007.6, 1007.5, 1008, 1008.3, 1008, 1007.9, 1007.7, 
    1007.8, 1007.8, 1007.8, 1007.8, 1007.5, 1007.2, 1006.4, 1005.7, 1005.2, 
    1004.6, 1003.9, 1003.3, 1002.7, 1002, 1001.7, 1001.2, 1000.8, 1000.2, 
    999.5, 999.1, 998.5, 998.1, 997.6, 997.1, 996.7, 996.5, 996.2, 995.8, 
    995.4, 994.8, 994.3, 994.4, 994.2, 993.9, 993, 992.6, 992, 991.8, 991.5, 
    990.7, 990.1, 989.7, 988.8, 988.1, 987.4, 986.6, 986.3, 985.8, 985.1, 
    984.6, 984.6, 984.4, 983.8, 983.3, 982.7, 982.1, 981.6, 981, 980.4, 
    979.5, 978.8, 978, 977.2, 976.7, 975.8, 975.5, 976.3, 976.4, 976.3, 976, 
    976.2, 976.3, 976.9, 977.7, 978.5, 978.7, 978.6, 979.2, 979.4, 978.9, 
    980.3, 980.8, 981.5, 982.2, 983.2, 984, 984.5, 985.5, 986.5, 987.3, 
    987.7, 988.6, 989, 989.9, 990.6, 991, 991.2, 991.7, 992, 992.3, 992.3, 
    992.4, 992.3, 992.6, 992.6, 993.2, 993.6, 994.1, 994.3, 994.6, 994.5, 
    994.5, 994.6, 994.4, 994.4, 994.3, 994, 994.4, 994.9, 994.6, 994.4, 
    994.2, 994.5, 994.8, 994.7, 994.6, 994.9, 995.3, 995.1, 995.2, 995, 
    995.2, 995.6, 995.6, 995.6, 996, 996, 996.1, 996.1, 996.3, 996.2, 996.5, 
    996.6, 996.6, 996.8, 996.9, 997.3, 997.5, 997.7, 998, 998.1, 998.2, 998, 
    997.9, 997.8, 998.1, 998, 998.3, 998.6, 999, 999.1, 999.4, 999.4, 999.4, 
    999.8, 999.9, 999.7, 1000, 1000.3, 1000.9, 1001.3, 1001.5, 1001.6, 1002, 
    1002.3, 1002.6, 1003, 1003.2, 1003.5, 1003.9, 1004.1, 1004.6, 1005, 
    1005.4, 1005.6, 1005.8, 1005.9, 1006.3, 1006.3, 1006.4, 1006.5, 1006.8, 
    1007.2, 1007.8, 1007.9, 1008.2, 1008.6, 1008.8, 1009.1, 1009.3, 1009.4, 
    1009.9, 1010.1, 1010.4, 1010.8, 1011.1, 1011.9, 1012.2, 1012.3, 1012.4, 
    1013, 1013.3, 1013.2, 1013.5, 1013.7, 1014, 1014.2, 1014.5, 1015, 1015.1, 
    1015.1, 1015, 1014.8, 1014.1, 1013.5, 1012.2, 1010.8, 1009.7, 1008.3, 
    1006.4, 1005.1, 1003.6, 1001.8, 1000.2, 999.9, 999, 999.3, 999.6, 1000.3, 
    1000.6, 1000.9, 1001.4, 1002, 1002.6, 1003.7, 1004.6, 1005.8, 1006.4, 
    1007.2, 1007.7, 1007.9, 1007.9, 1008.1, 1008.2, 1008.1, 1008, 1006.7, 
    1006.5, 1006, 1005.8, 1005.5, 1005.3, 1005.3, 1005.5, 1006, 1006.4, 
    1007.2, 1007.9, 1008.7, 1009.3, 1010.4, 1012.1, 1013, 1014.3, 1015.8, 
    1017, 1018.2, 1019.4, 1020.1, 1021, 1021.8, 1022.4, 1022.9, 1023.7, 
    1024.4, 1025.3, 1025.7, 1026.3, 1026.8, 1027.2, 1027.6, 1027.8, 1027.9, 
    1028, 1028.1, 1027.9, 1028, 1028, 1028.2, 1028.3, 1028.7, 1029.3, 1029.9, 
    1030, 1030.1, 1030.4, 1030.7, 1031.1, 1031.8, 1032.2, 1032.3, 1032.6, 
    1032.9, 1033, 1033.3, 1033.6, 1033.8, 1034, 1034.1, 1034.1, 1034.2, 1034, 
    1034, 1033.9, 1033.9, 1033.8, 1033.1, 1032.4, 1032, 1031.6, 1031.3, 
    1030.3, 1029.6, 1029.1, 1028.1, 1027.1, 1026, 1025.2, 1024.6, 1024.3, 
    1023.9, 1023.5, 1023.2, 1022.9, 1022.5, 1022.2, 1021.7, 1021.3, 1021, 
    1020.6, 1020.2, 1019.7, 1019.1, 1018.5, 1018.1, 1017.7, 1017.3, 1016.8, 
    1016.1, 1015.8, 1015.2, 1014.9, 1014.6, 1014.3, 1014.1, 1013.9, 1014, 
    1014, 1013.8, 1013.9, 1014, 1014.2, 1014.4, 1014.5, 1014.7, 1015, 1015.5, 
    1015.7, 1016, 1016, 1016.2, 1016.5, 1016.7, 1017.1, 1017.7, 1018.2, 
    1018.9, 1019.6, 1020, 1020.5, 1020.9, 1021.2, 1021.5, 1021.8, 1022, 
    1022.1, 1022.4, 1022.5, 1022.9, 1022.7, 1022.6, 1022.7, 1022.7, 1022.5, 
    1022.3, 1021.9, 1021.7, 1021.4, 1021.1, 1020.8, 1020.3, 1020, 1019.7, 
    1019.5, 1019.1, 1018.5, 1018, 1017.5, 1017.3, 1016.7, 1016.4, 1016.3, 
    1016, 1015.4, 1015.6, 1015.1, 1014.9, 1014.5, 1014.2, 1013.9, 1013.9, 
    1013.5, 1013.5, 1013.9, 1014.1, 1013.9, 1013.9, 1014.1, 1013.8, 1013.7, 
    1013.2, 1013.1, 1012.5, 1012.4, 1012.7, 1012.8, 1012.9, 1012.6, 1012.7, 
    1012.9, 1013.1, 1012.4, 1011.4, 1010.9, 1010, 1009.4, 1008.6, 1007.6, 
    1007.7, 1007.3, 1007.4, 1007.7, 1008.3, 1008.3, 1008.4, 1008.7, 1009, 
    1009.3, 1009.8, 1010.3, 1010.9, 1011.5, 1012, 1012.8, 1014, 1015, 1015.9, 
    1016.9, 1017.9, 1018.8, 1019.4, 1020.3, 1021.2, 1021.4, 1021.7, 1021.8, 
    1021.5, 1021.1, 1020.5, 1019.9, 1019.6, 1019.3, 1018.8, 1018.2, 1017.7, 
    1017, 1016.3, 1016.3, 1015.8, 1015.3, 1015.5, 1015.1, 1014.9, 1015.2, 
    1015.4, 1015.9, 1016.1, 1016.2, 1016.3, 1016.1, 1015.6, 1015, 1014.6, 
    1014.5, 1014, 1013.2, 1012.7, 1012.5, 1012.4, 1012.5, 1012.4, 1012.9, 
    1013.4, 1014.1, 1014.5, 1015.1, 1015.6, 1016.4, 1017.2, 1017.8, 1018.4, 
    1018.9, 1019.1, 1019.3, 1019.2, 1019.3, 1019.1, 1018.7, 1018.3, 1018, 
    1017.4, 1016.8, 1016.7, 1016.4, 1016.3, 1015.7, 1015.4, 1015.2, 1015.2, 
    1014.8, 1014.4, 1014.4, 1014.4, 1014.5, 1014.5, 1014.4, 1014.4, 1014.5, 
    1014.4, 1014.4, 1014.3, 1013.9, 1013.5, 1012.9, 1012.5, 1012.3, 1012.3, 
    1012.6, 1012.3, 1011.8, 1011.6, 1011.8, 1011.6, 1011.3, 1011.1, 1011.1, 
    1011.2, 1011.1, 1010.8, 1010.5, 1010.2, 1009.3, 1008.3, 1007.3, 1006.2, 
    1005.3, 1004.4, 1003.3, 1002.1, 1001.7, 1001.5, 1001.5, 1001.4, 1001.6, 
    1003, 1004.5, 1005.7, 1006.6, 1007.4, 1007.9, 1008.4, 1007.9, 1008.3, 
    1008.5, 1008.3, 1008.1, 1007.5, 1006.5, 1005.7, 1005.2, 1004.1, 1002.9, 
    1002.1, 1001.8, 1001.3, 1001.1, 1000.7, 1000, 999.6, 999.4, 999.3, 999.4, 
    999.3, 999.3, 999.4, 999.7, 1000.3, 1000.7, 1001, 1001.4, 1001.7, 1002.4, 
    1003.6, 1004.4, 1005.3, 1006.1, 1006.8, 1007.6, 1008.5, 1009.3, 1010, 
    1010.8, 1011.5, 1011.8, 1012.2, 1012.6, 1013, 1013.4, 1013.9, 1014.2, 
    1014.4, 1014.3, 1014.4, 1014.3, 1014.2, 1013.8, 1013.3, 1013.2, 1012.9, 
    1012.5, 1011.9, 1011.7, 1011.6, 1011.4, 1011.2, 1010.7, 1010.4, 1010.4, 
    1010.2, 1010.1, 1010.3, 1010.4, 1010.6, 1010.9, 1011.2, 1011.5, 1011.7, 
    1012.1, 1012.5, 1012.8, 1013.2, 1013.6, 1013.9, 1014.4, 1014.7, 1015.2, 
    1015.8, 1016.3, 1016.9, 1017.6, 1018.2, 1018.9, 1019.5, 1020.3, 1020.9, 
    1021.5, 1022.2, 1022.6, 1023.3, 1023.9, 1024, 1024.4, 1024.6, 1024.4, 
    1024.6, 1024.3, 1024.2, 1024, 1024, 1024.4, 1024.5, 1024.6, 1024.7, 
    1024.7, 1024.8, 1024.9, 1025, 1025, 1024.7, 1024.8, 1024.9, 1024.9, 1025, 
    1025, 1025, 1024.7, 1024.7, 1024.3, 1024.1, 1023.6, 1023.1, 1022.9, 
    1022.5, 1022.5, 1022.4, 1022.6, 1022.4, 1022.4, 1022.4, 1022.5, 1022.7, 
    1022.7, 1023, 1023.2, 1023.3, 1023.5, 1024, 1024.6, 1024.9, 1025.3, 
    1025.7, 1026.1, 1026.5, 1026.7, 1026.8, 1027.1, 1027.3, 1027.5, 1027.7, 
    1028.1, 1028, 1028.1, 1028.1, 1027.9, 1027.7, 1027.6, 1027.3, 1027.2, 
    1027.1, 1027.1, 1027.1, 1027.1, 1027, 1026.7, 1026.4, 1026.2, 1026, 
    1025.7, 1025.4, 1025.1, 1024.8, 1024.6, 1024.4, 1024.2, 1023.9, 1023.7, 
    1023.6, 1023.6, 1023.6, 1023.7, 1023.7, 1023.9, 1024.1, 1024.4, 1024.6, 
    1024.9, 1025.2, 1025.4, 1025.5, 1025.9, 1026.2, 1026.1, 1026.1, 1026.3, 
    1026.5, 1026.8, 1026.9, 1027.1, 1027.1, 1027, 1026.9, 1026.9, 1026.4, 
    1026, 1025.5, 1025, 1024.4, 1024.1, 1023.6, 1022.8, 1022.3, 1021.1, 1020, 
    1019.1, 1018.2, 1017.2, 1016.8, 1017, 1017.3, 1018.2, 1019, 1019.1, 
    1019.2, 1020, 1020.4, 1020.9, 1021.1, 1021, 1020.9, 1020.9, 1021.2, 
    1021.1, 1021.3, 1020.9, 1020.7, 1020.4, 1020.4, 1019.7, 1020, 1019.6, 
    1019.4, 1019.1, 1018.4, 1018.4, 1018.3, 1018.4, 1018.4, 1017.9, 1017.7, 
    1017.2, 1016.8, 1016.5, 1016.2, 1016.1, 1016.1, 1016.5, 1016.9, 1017.3, 
    1017.5, 1017.9, 1018.5, 1017.9, 1018.5, 1019.3, 1020.1, 1021, 1021.2, 
    1022.8, 1023.6, 1024.9, 1025.3, 1025.9, 1025.6, 1025.6, 1026.1, 1026.5, 
    1027.3, 1027.1, 1027.4, 1027.5, 1027.3, 1027.1, 1027.2, 1026.9, 1025.9, 
    1024.4, 1023.9, 1022.8, 1021.2, 1019.6, 1018.1, 1017.3, 1015.9, 1014.5, 
    1013.5, 1012.8, 1012.1, 1011.5, 1010.8, 1011.2, 1010.6, 1010.3, 1010.1, 
    1009.9, 1009.9, 1010, 1010.4, 1010.9, 1011.4, 1011.2, 1011.4, 1012, 
    1011.7, 1012.5, 1012.7, 1012.7, 1013.1, 1013.4, 1013.7, 1013.8, 1014.4, 
    1014.7, 1015.2, 1015.5, 1016.3, 1016.9, 1017.6, 1018.1, 1019, 1019.4, 
    1019.9, 1020.4, 1020.7, 1021.2, 1021.3, 1021.7, 1021.8, 1022, 1022.5, 
    1022.8, 1022.5, 1022.9, 1023.2, 1023.5, 1023.4, 1023.4, 1023.3, 1023.4, 
    1023.3, 1023.4, 1023, 1023.1, 1023, 1022.9, 1022.9, 1022.9, 1023.1, 
    1022.9, 1022.6, 1022.4, 1022.2, 1022.1, 1021.7, 1021.7, 1021.2, 1020.8, 
    1020.6, 1020.5, 1020.3, 1020.1, 1020.3, 1020.6, 1020.7, 1020.6, 1020.6, 
    1020.9, 1021, 1021.2, 1021.3, 1021.4, 1021.7, 1021.8, 1021.5, 1021.4, 
    1021.5, 1022, 1022.4, 1022.8, 1022.9, 1023.3, 1023.7, 1023.9, 1024, 
    1024.4, 1024.6, 1024.6, 1024.8, 1025.2, 1025.2, 1025.3, 1025.4, 1025.4, 
    1025.5, 1025.6, 1025.9, 1025.2, 1025.2, 1025.4, 1025.3, 1025.6, 1025.9, 
    1026.2, 1026.4, 1026.8, 1026.6, 1027.1, 1027.4, 1027.3, 1027.4, 1027.4, 
    1027.7, 1027.9, 1028.1, 1028.3, 1028.1, 1028, 1027.9, 1027.8, 1027.5, 
    1027.3, 1027.1, 1026.8, 1026.3, 1026, 1025.7, 1025, 1024.8, 1024.4, 1024, 
    1023.6, 1023.1, 1022.5, 1021.7, 1020.7, 1020.4, 1020.1, 1019.6, 1019.8, 
    1019.7, 1019.7, 1019.4, 1019.4, 1019.4, 1019.5, 1019.7, 1019.8, 1019.9, 
    1020.1, 1020.3, 1020.8, 1021.1, 1022, 1022.8, 1023.4, 1023.9, 1024.4, 
    1024.8, 1025.3, 1025.5, 1025.9, 1026.1, 1026.6, 1027.2, 1027.6, 1027.8, 
    1028.1, 1028.2, 1028.4, 1028.7, 1029, 1029.2, 1029.6, 1029.9, 1030.3, 
    1030.6, 1030.9, 1031, 1031.1, 1031.2, 1031.1, 1031.1, 1031.1, 1031, 1031, 
    1031.2, 1031.2, 1031.2, 1031.2, 1031, 1030.9, 1030.9, 1030.7, 1030.6, 
    1030.5, 1030.6, 1030.7, 1030.8, 1031, 1030.9, 1030.9, 1031.1, 1031.4, 
    1031.3, 1031, 1030.8, 1030.9, 1031.1, 1030.9, 1031.1, 1031.5, 1031.7, 
    1031.5, 1031.7, 1031.6, 1031, 1030.6, 1030.5, 1030.2, 1030, 1029.9, 
    1029.8, 1029.7, 1029.5, 1029.3, 1028.6, 1028, 1027.7, 1027.5, 1026.5, 
    1026, 1025.6, 1025.1, 1024.6, 1024.6, 1024.3, 1023.6, 1023.6, 1022.1, 
    1020.6, 1020, 1019.7, 1018.8, 1017.9, 1018.5, 1017.1, 1017, 1016.6, 
    1016.1, 1015.4, 1014.9, 1014.4, 1014, 1013.5, 1013.1, 1012.6, 1012.3, 
    1012, 1012, 1011.4, 1010.9, 1010.8, 1010, 1009.6, 1009.3, 1008.9, 1008.3, 
    1007.8, 1007.5, 1007.4, 1007.3, 1007.3, 1007, 1007, 1007.1, 1007.1, 
    1007.3, 1007.4, 1007.4, 1007.5, 1007.7, 1008, 1008.2, 1008.5, 1008.7, 
    1008.9, 1009.2, 1009.6, 1010.2, 1010.5, 1010.7, 1010.9, 1011.1, 1011.3, 
    1011.7, 1011.9, 1012.3, 1012.5, 1012.7, 1013.3, 1013.4, 1013.7, 1014, 
    1013.9, 1014.1, 1014.8, 1015.4, 1016, 1016.4, 1016.9, 1017.6, 1018.3, 
    1018.8, 1019.3, 1019.6, 1019.9, 1020.3, 1020.7, 1021.3, 1021.8, 1022.1, 
    1022.3, 1022.4, 1022.7, 1022.9, 1023.1, 1023.2, 1023.5, 1023.6, 1023.9, 
    1024, 1024.1, 1024.3, 1024.4, 1024.7, 1024.8, 1025, 1025.3, 1025.2, 
    1025.2, 1025.7, 1025.6, 1025.8, 1025.9, 1026.1, 1026.3, 1026.4, 1026.8, 
    1026.9, 1027.3, 1027.2, 1027.4, 1027.5, 1027.7, 1027.9, 1028.2, 1028.7, 
    1028.8, 1028.9, 1029.1, 1029.1, 1029.3, 1029, 1029.3, 1029.2, 1029.2, 
    1029.4, 1029.6, 1029.7, 1029.8, 1029.6, 1029.5, 1029.5, 1029.4, 1029.5, 
    1029.6, 1029.6, 1029.6, 1029.8, 1029.9, 1030.2, 1030.4, 1030.5, 1030.5, 
    1030.7, 1030.8, 1030.7, 1030.5, 1030.4, 1030.3, 1030.3, 1030.5, 1030.3, 
    1030.4, 1030.2, 1030.2, 1029.9, 1029.8, 1029.7, 1029.7, 1029.7, 1029.8, 
    1029.9, 1030, 1030.1, 1030.4, 1030.3, 1030.3, 1030.4, 1030.4, 1030.4, 
    1030.4, 1030.3, 1030.2, 1030.3, 1030.3, 1030.2, 1030.1, 1030.2, 1030.2, 
    1030.1, 1030, 1029.8, 1029.7, 1029.6, 1029.6, 1029.6, 1029.7, 1029.7, 
    1029.7, 1029.7, 1029.5, 1029.5, 1029.5, 1029.4, 1029.6, 1029.8, 1030, 
    1030.2, 1030.6, 1031, 1031.1, 1031.5, 1031.6, 1031.6, 1031.5, 1031.5, 
    1031.5, 1031.4, 1031.4, 1031.2, 1030.9, 1030.7, 1030.5, 1030.3, 1030, 
    1029.8, 1029.3, 1028.9, 1028.7, 1028.2, 1027.9, 1027.7, 1027.2, 1027.5, 
    1027.2, 1026.9, 1026.9, 1026.3, 1025.9, 1025.5, 1025.3, 1024.9, 1024.5, 
    1024.4, 1023.8, 1023.7, 1023.4, 1022.9, 1022.3, 1021.8, 1021.1, 1020.6, 
    1020.1, 1019.6, 1019.5, 1019, 1018.6, 1018.2, 1017.9, 1017.1, 1017.3, 
    1017.2, 1017, 1016.9, 1016.7, 1016.6, 1016.4, 1016.2, 1016.3, 1016.5, 
    1016.4, 1016.4, 1016.3, 1016.4, 1016.4, 1016.1, 1016.2, 1016.2, 1016.3, 
    1016.6, 1016.9, 1017, 1017.3, 1017.5, 1017.8, 1017.6, 1017.5, 1017.5, 
    1017.2, 1016.9, 1016.7, 1016.6, 1016.1, 1015.9, 1015.5, 1015.3, 1015, 
    1014.7, 1014.6, 1014.4, 1014, 1013.7, 1013.4, 1013.3, 1013, 1013, 1013.2, 
    1013.6, 1013.5, 1013.5, 1013.5, 1013.8, 1013.8, 1014.1, 1014.5, 1014.9, 
    1015.4, 1015.5, 1016.2, 1016.8, 1016.9, 1017, 1017.1, 1017.1, 1017.1, 
    1017.3, 1017.6, 1017.8, 1017.8, 1018, 1018.1, 1018.4, 1018.6, 1018.7, 
    1018.7, 1018.8, 1019, 1019, 1019, 1019.1, 1019.3, 1019, 1019, 1018.9, 
    1018.9, 1018.6, 1018.4, 1018.1, 1017.8, 1017.8, 1017.7, 1017.5, 1017.5, 
    1017.3, 1017.1, 1016.5, 1016.4, 1016, 1015.6, 1015, 1015, 1014.6, 1014.2, 
    1014, 1013.9, 1013.8, 1013.7, 1013.7, 1013.9, 1013.9, 1014, 1014, 1014.1, 
    1014, 1014.1, 1014.2, 1014.3, 1014.5, 1014.7, 1014.9, 1015, 1015.4, 
    1015.7, 1016, 1016.4, 1017, 1017.6, 1018.3, 1018.8, 1019.1, 1019.6, 
    1020.1, 1020.4, 1020.7, 1021, 1021.4, 1021.8, 1022.1, 1022.5, 1022.7, 
    1022.7, 1022.6, 1022.9, 1023.2, 1023.3, 1023.5, 1023.6, 1023, 1022.9, 
    1022.6, 1022.5, 1023.1, 1022.5, 1022.1, 1021.5, 1021.2, 1021.1, 1021, 
    1020.8, 1020.4, 1020, 1019.5, 1019.1, 1018.7, 1018.4, 1018, 1018.2, 
    1017.5, 1016.5, 1016.2, 1016.3, 1017.1, 1019.3, 1016.8, 1016.6, 1016.1, 
    1016.8, 1016.6, 1016.4, 1016.6, 1017.3, 1017.5, 1017.5, 1017.6, 1017.4, 
    1017.6, 1017.9, 1017.9, 1017.9, 1017.7, 1017.6, 1017.6, 1018, 1018, 
    1018.1, 1018, 1017.9, 1017.9, 1017.7, 1017.7, 1017.7, 1018.2, 1018.3, 
    1018.4, 1018.5, 1017.8, 1017.7, 1017.3, 1017, 1016.8, 1016.4, 1016.5, 
    1016.3, 1016, 1015.7, 1015.3, 1015.2, 1014.8, 1014.3, 1014, 1013.6, 1013, 
    1012.7, 1012.5, 1012.7, 1012.5, 1012.4, 1012.4, 1012.3, 1011.9, 1011.6, 
    1011.4, 1011.4, 1011.3, 1011.2, 1011.3, 1011.2, 1011.1, 1011.1, 1011, 
    1010.9, 1011, 1010.8, 1010.6, 1010.6, 1010.3, 1010.4, 1010.3, 1010.3, 
    1010.5, 1010.4, 1010.4, 1010.3, 1010.3, 1010.1, 1009.9, 1009.6, 1009.2, 
    1008.9, 1008.7, 1008.7, 1008.5, 1008.4, 1008.3, 1008.3, 1008.4, 1008.2, 
    1008.3, 1008.3, 1008.3, 1008.5, 1008.5, 1008.7, 1008.8, 1008.8, 1009, 
    1009.2, 1009.1, 1009.2, 1009.3, 1009.2, 1009.2, 1009.3, 1009.4, 1009.4, 
    1009.7, 1009.7, 1009.9, 1010, 1009.9, 1009.9, 1009.8, 1009.9, 1009.9, 
    1010, 1010.3, 1010.3, 1010.5, 1010.7, 1010.6, 1010.8, 1010.6, 1010.4, 
    1010.4, 1010.4, 1010.5, 1010.7, 1010.8, 1010.9, 1011, 1011.1, 1011, 
    1010.8, 1011.1, 1011.2, 1011.1, 1011.1, 1011.2, 1011.3, 1011.5, 1011.6, 
    1011.8, 1011.8, 1011.9, 1012.1, 1012.3, 1012.4, 1012.5, 1012.8, 1013, 
    1013.1, 1013.3, 1013.6, 1013.8, 1014.1, 1014.4, 1014.6, 1014.9, 1014.8, 
    1014.9, 1015, 1015.1, 1015.6, 1015.6, 1016, 1016.3, 1016.3, 1016.7, 
    1016.8, 1016.8, 1016.8, 1016.6, 1016.5, 1016.5, 1016.6, 1016.9, 1017.2, 
    1017.5, 1017.6, 1017.5, 1017.5, 1017.7, 1017.7, 1018.1, 1018.1, 1018.4, 
    1018.4, 1018.7, 1019.1, 1019.2, 1019.6, 1019.7, 1019.9, 1020, 1020.3, 
    1020.5, 1020.7, 1020.9, 1021.3, 1021.8, 1022.2, 1022.4, 1022.5, 1022.8, 
    1022.7, 1023, 1023.1, 1023.1, 1023.2, 1023.5, 1023.6, 1023.6, 1023.6, 
    1023.9, 1023.8, 1023.8, 1023.8, 1023.7, 1023.7, 1023.7, 1023.5, 1023.6, 
    1023.5, 1023.7, 1023.7, 1023.8, 1023.7, 1023.6, 1023.5, 1023.3, 1023, 
    1022.6, 1022.6, 1022.6, 1022.6, 1022.8, 1022.8, 1023.2, 1023, 1022.9, 
    1023.1, 1023.3, 1023.5, 1023.6, 1023.7, 1024, 1024, 1024.3, 1024.7, 
    1024.9, 1025, 1025.1, 1025.1, 1025, 1025.1, 1024.9, 1024.9, 1024.9, 1025, 
    1025, 1025.3, 1025.3, 1025.3, 1025.4, 1025.3, 1025.4, 1025.4, 1025.4, 
    1025.3, 1025.3, 1025.3, 1025.3, 1025.5, 1025.6, 1025.8, 1025.7, 1025.9, 
    1026.1, 1026.1, 1026.1, 1026.3, 1026.4, 1026.9, 1027, 1027.6, 1027.8, 
    1027.9, 1028.1, 1028.1, 1028.2, 1028.1, 1027.7, 1028.1, 1027.7, 1027.9, 
    1027.7, 1027.6, 1027.7, 1027.4, 1027.1, 1027, 1026.3, 1026, 1025.7, 
    1025.1, 1024.8, 1024, 1023.6, 1023.2, 1022.6, 1022.3, 1021.8, 1021, 
    1020.9, 1020.7, 1020.7, 1020.5, 1020.1, 1020.2, 1019.8, 1019.9, 1019.7, 
    1019.3, 1019, 1018.9, 1018.5, 1018, 1018.4, 1018.4, 1018.5, 1018.8, 
    1019.1, 1019.4, 1019.6, 1019.3, 1019.1, 1018.6, 1018.1, 1018, 1017.5, 
    1017.2, 1016.4, 1015.6, 1015.2, 1014.5, 1014.1, 1013.4, 1012.9, 1012.3, 
    1011.6, 1011.2, 1011, 1010.8, 1010.4, 1010.2, 1010.2, 1010.2, 1010.4, 
    1010.6, 1010.8, 1010.8, 1010.6, 1010.8, 1010.8, 1011.1, 1011.2, 1011.4, 
    1011.4, 1011.3, 1011.6, 1011.5, 1011.2, 1010.6, 1010.2, 1010, 1010, 
    1009.9, 1010.6, 1009.9, 1009.9, 1010.1, 1009.8, 1009.5, 1009.4, 1009.1, 
    1009, 1009.1, 1009.2, 1009.3, 1009, 1009, 1008.7, 1008.7, 1008.9, 1008.8, 
    1008.9, 1009, 1008.9, 1008.7, 1008.8, 1008.8, 1008.8, 1008.9, 1008.9, 
    1009.1, 1009.4, 1009.7, 1009.8, 1009.9, 1009.8, 1009.7, 1009.8, 1009.7, 
    1009.7, 1009.6, 1009.5, 1009.4, 1009.3, 1009.1, 1008.9, 1008.8, 1008.7, 
    1008.5, 1008.4, 1008.3, 1008.1, 1007.8, 1008.1, 1008.1, 1008.1, 1008, 
    1008.3, 1008.6, 1008.8, 1008.9, 1008.8, 1008.9, 1009.2, 1009.1, 1009.1, 
    1009, 1008.8, 1008.7, 1008.7, 1008.6, 1008.4, 1008.3, 1008.1, 1007.8, 
    1007.6, 1007.7, 1007.8, 1008.2, 1008.4, 1008.7, 1008.9, 1009, 1009, 
    1009.1, 1009.2, 1009.1, 1009.2, 1009.3, 1009.6, 1010, 1010.2, 1010.3, 
    1010.8, 1011, 1011.3, 1011.4, 1011.5, 1011.7, 1011.9, 1012.2, 1012.6, 
    1012.9, 1013.3, 1013.6, 1013.9, 1014.1, 1014.4, 1014.5, 1014.7, 1014.7, 
    1014.7, 1014.9, 1015.2, 1015.3, 1015.6, 1015.7, 1015.7, 1015.7, 1015.7, 
    1015.6, 1015.5, 1015.3, 1015.1, 1014.9, 1014.8, 1014.8, 1014.9, 1014.6, 
    1014.4, 1014.4, 1014.2, 1014.2, 1014, 1013.9, 1013.8, 1013.7, 1013.7, 
    1013.7, 1013.8, 1013.9, 1013.7, 1013.9, 1014, 1013.8, 1013.7, 1013.6, 
    1013.3, 1013.3, 1013.5, 1013.6, 1013.6, 1013.5, 1013.7, 1013.8, 1013.9, 
    1014, 1014, 1014, 1014, 1014, 1014.1, 1014.1, 1014.4, 1014.6, 1014.8, 
    1014.9, 1015, 1015.1, 1015.1, 1015.3, 1015.3, 1015.4, 1015.7, 1015.9, 
    1016.2, 1016.4, 1016.6, 1016.8, 1016.8, 1017, 1017.1, 1016.9, 1017, 1017, 
    1017.1, 1017, 1017.3, 1017.3, 1017.1, 1017.1, 1016.9, 1016.8, 1016.5, 
    1016.2, 1015.9, 1015.6, 1015.2, 1015.1, 1014.8, 1014.5, 1014.3, 1013.8, 
    1013.7, 1013.4, 1013, 1012.5, 1012.1, 1011.9, 1011.6, 1011.4, 1011.1, 
    1010.9, 1010.7, 1010.2, 1010, 1009.6, 1009.3, 1008.9, 1008.5, 1008.2, 
    1008.2, 1008.1, 1007.7, 1007.7, 1007.6, 1007.4, 1007.2, 1007, 1006.8, 
    1006.4, 1006.3, 1006.3, 1006.2, 1006.1, 1006.1, 1006.1, 1006, 1006.1, 
    1005.7, 1005.6, 1005.2, 1004.9, 1004.7, 1004.7, 1004.4, 1004, 1003.7, 
    1003.5, 1003, 1002.7, 1002.1, 1001.5, 1001, 1000.3, 999.6, 998.9, 998.3, 
    997.8, 997.2, 996.5, 996, 995.6, 995, 994.7, 994.3, 994, 993.9, 994.2, 
    994.5, 994.7, 995.2, 995.6, 995.7, 996, 996.4, 996.7, 996.7, 996.9, 
    996.8, 996.8, 997, 997.1, 997.2, 997.9, 998.2, 998.5, 998.8, 999.4, 1000, 
    1000.7, 1001, 1001.6, 1001.9, 1002.4, 1002.9, 1003.1, 1003.4, 1003.7, 
    1003.9, 1003.8, 1004.2, 1004.4, 1004.4, 1004.3, 1004.5, 1004.4, 1004.3, 
    1004.3, 1003.7, 1003.6, 1003.8, 1003.5, 1003.3, 1003.8, 1004.4, 1004.2, 
    1004.2, 1004.5, 1004.7, 1005, 1005.2, 1005.5, 1005.6, 1006, 1006.4, 
    1006.5, 1006.5, 1007.1, 1008, 1008.6, 1009.3, 1009.8, 1010, 1010.7, 
    1010.9, 1010.9, 1011.6, 1011.9, 1012.5, 1012.7, 1012.9, 1013.1, 1012.9, 
    1012.7, 1012.5, 1012.1, 1012.1, 1012.1, 1011.3, 1010.3, 1009.7, 1009, 
    1008.7, 1008.2, 1007.2, 1006.9, 1006.4, 1005.9, 1005.7, 1005.8, 1005.4, 
    1005, 1004.5, 1004.1, 1004.5, 1004.2, 1004, 1004.3, 1004.6, 1004.8, 
    1005.1, 1005.7, 1006, 1006, 1005.8, 1005.8, 1005.9, 1005.6, 1005.3, 
    1004.9, 1004.1, 1004.6, 1005, 1005, 1004.8, 1005, 1004.7, 1005, 1005.2, 
    1005.1, 1004.9, 1005.2, 1005.3, 1005.8, 1006.7, 1007.4, 1007.5, 1007.7, 
    1007.9, 1008.1, 1008.3, 1008.8, 1009.1, 1009.4, 1009.6, 1009.7, 1010.3, 
    1010.9, 1011.2, 1011.9, 1012.3, 1012.9, 1013.4, 1013.7, 1014.1, 1014.5, 
    1014.7, 1015.1, 1015.6, 1016, 1016.2, 1016.6, 1016.8, 1017.1, 1017.4, 
    1017.5, 1017.8, 1018.1, 1018.4, 1018.5, 1018.6, 1018.9, 1018.9, 1019.2, 
    1019.2, 1019.4, 1019.6, 1019.9, 1020, 1019.9, 1020.2, 1020, 1019.9, 
    1019.9, 1019.9, 1019.9, 1019.5, 1020, 1020, 1019.8, 1019.6, 1018.9, 
    1018.4, 1018, 1018, 1018, 1017.6, 1017.2, 1016.7, 1016.5, 1016.3, 1016.1, 
    1016.6, 1016.4, 1016.4, 1015.9, 1015.8, 1016.3, 1015.8, 1016.3, 1016.5, 
    1016.9, 1017.2, 1017.7, 1018.1, 1018.3, 1018.2, 1018.1, 1018.2, 1018.6, 
    1018.7, 1018.7, 1018.9, 1019.1, 1019.5, 1019.8, 1019.9, 1020.1, 1020.5, 
    1020.7, 1020.6, 1020.8, 1021.2, 1021.5, 1021.3, 1021.2, 1021.5, 1021.9, 
    1022.3, 1022.7, 1023, 1023.2, 1023.4, 1023.5, 1023.8, 1023.8, 1023.8, 
    1023.8, 1023.7, 1023.8, 1024, 1024.2, 1024.4, 1024.4, 1024.6, 1024.6, 
    1024.6, 1024.5, 1024.4, 1024.5, 1024.6, 1024.5, 1024.6, 1024.5, 1024.3, 
    1024.2, 1023.8, 1023.7, 1023.5, 1023.3, 1023.2, 1023.1, 1023.1, 1023.2, 
    1023.1, 1023, 1022.9, 1022.9, 1022.5, 1022.4, 1022.5, 1022.5, 1022.5, 
    1022.5, 1022.3, 1022.4, 1022.5, 1022.5, 1022.4, 1022.2, 1022, 1021.8, 
    1021.8, 1021.4, 1024.1, 1021.4, 1021.5, 1021.2, 1021, 1020.6, 1020.3, 
    1020.1, 1019.8, 1019.5, 1019.3, 1018.7, 1018.4, 1018.1, 1017.9, 1017.6, 
    1017.2, 1017, 1016.5, 1016.1, 1015.9, 1015.4, 1015.1, 1014.8, 1014.6, 
    1014.6, 1014.6, 1014.5, 1014.3, 1014.2, 1014, 1013.8, 1013.6, 1013.7, 
    1013.5, 1013.6, 1013.5, 1013.4, 1013.5, 1013.4, 1013.2, 1013.2, 1013.2, 
    1013.1, 1013.1, 1013.1, 1013, 1012.9, 1013.1, 1013.3, 1013.3, 1013.4, 
    1013.3, 1013.5, 1013.5, 1013.5, 1013.3, 1013.4, 1013.3, 1013.1, 1013.1, 
    1013.2, 1013.3, 1013.3, 1013.3, 1013.3, 1013.3, 1013.3, 1013.4, 1013.2, 
    1013.2, 1013.1, 1013.1, 1012.8, 1013, 1013.3, 1013.4, 1013.4, 1013.6, 
    1013.7, 1013.8, 1013.9, 1014.1, 1014.1, 1014.2, 1014.4, 1014.5, 1014.7, 
    1014.8, 1014.7, 1014.7, 1014.6, 1014.5, 1014.7, 1014.6, 1014.5, 1014.7, 
    1015, 1015.5, 1015.5, 1015.5, 1015.5, 1015.6, 1015.3, 1015.1, 1015.1, 
    1015.2, 1015.1, 1014.9, 1015, 1014.9, 1015, 1015.1, 1015.1, 1015.3, 
    1015.3, 1015.2, 1015.3, 1015.3, 1015.3, 1015.2, 1015.3, 1015.7, 1015.8, 
    1015.8, 1015.6, 1015.5, 1015.5, 1015.7, 1015.9, 1015.9, 1016, 1016, 
    1016.2, 1016.4, 1016.5, 1016.5, 1016.5, 1016.6, 1016.6, 1016.6, 1016.6, 
    1016.7, 1016.7, 1016.7, 1016.9, 1017, 1017.1, 1017.1, 1017.1, 1017.1, 
    1017.3, 1017.2, 1017.2, 1017.3, 1017.3, 1017.3, 1017.5, 1017.6, 1017.8, 
    1018.1, 1018.2, 1018.2, 1018.4, 1018.5, 1018.6, 1018.7, 1018.9, 1018.9, 
    1019.1, 1019.5, 1019.9, 1020, 1014.4, 1019.9, 1020.1, 1020.3, 1020.5, 
    1020.8, 1021.2, 1021.3, 1021.5, 1021.8, 1022.2, 1022.5, 1022.5, 1022.6, 
    1022.6, 1022.5, 1022.5, 1022.3, 1022.2, 1022, 1021.8, 1021.4, 1021.2, 
    1021.2, 1020.6, 1020.3, 1019.9, 1019.5, 1018.7, 1018.2, 1017.6, 1016.6, 
    1015.8, 1015.1, 1014.1, 1013.6, 1013, 1012.1, 1011.2, 1010.1, 1009.4, 
    1008.3, 1007.5, 1007, 1006.4, 1006, 1005.8, 1005.9, 1005.8, 1005.8, 
    1005.8, 1006, 1006.5, 1007.2, 1008, 1008.5, 1009, 1009.6, 1010.2, 1011.3, 
    1011.9, 1012.4, 1012.9, 1013.4, 1013.6, 1013.7, 1013.9, 1014.2, 1014.5, 
    1014.7, 1014.8, 1014.8, 1015.1, 1015.1, 1015, 1014.8, 1014.7, 1014.8, 
    1014.7, 1014.5, 1014.5, 1014.5, 1014.1, 1014.1, 1014.1, 1014, 1013.6, 
    1013.2, 1012.9, 1012.9, 1012.8, 1012.6, 1012.7, 1012.7, 1012.6, 1012.5, 
    1012.7, 1012.5, 1012.3, 1012.1, 1012.1, 1012, 1011.7, 1011.5, 1011.5, 
    1011.4, 1011.6, 1011.8, 1012.1, 1012.1, 1012.3, 1012.2, 1012.5, 1012.6, 
    1012.5, 1012.3, 1012.4, 1012.5, 1012.5, 1012.5, 1012.7, 1012.5, 1012.5, 
    1012.2, 1012, 1012, 1011.7, 1011.7, 1011.6, 1011.7, 1011.7, 1011.6, 
    1011.9, 1011.6, 1011.4, 1011.4, 1011.4, 1011.2, 1011, 1010.9, 1010.9, 
    1011, 1011, 1011.2, 1011.3, 1011, 1010.9, 1010.8, 1010.3, 1010.3, 1010.4, 
    1010.4, 1010.4, 1010.4, 1010.7, 1011.1, 1011.3, 1011.3, 1011.6, 1011.8, 
    1011.8, 1012, 1012.4, 1012.6, 1012.9, 1013.4, 1014, 1014.2, 1014.5, 
    1014.6, 1015, 1015.2, 1015.2, 1015.4, 1015.6, 1015.6, 1016.1, 1016.3, 
    1016.6, 1016.6, 1016.7, 1016.8, 1016.6, 1016.6, 1016.7, 1016.6, 1016.5, 
    1016.6, 1016.4, 1016.5, 1016.7, 1016.8, 1016.7, 1016.4, 1016.1, 1016, 
    1016.2, 1016.4, 1016.6, 1016.9, 1017.3, 1017.4, 1017.7, 1017.9, 1018.4, 
    1019.1, 1019.8, 1020, 1020, 1020, 1020.2, 1020.3, 1020.6, 1020.8, 1021.2, 
    1021.3, 1021.5, 1021.7, 1021.7, 1021.5, 1021.7, 1021.9, 1022.2, 1022.3, 
    1022.5, 1022.9, 1022.8, 1023, 1023.1, 1023.2, 1023.2, 1023.2, 1023.1, 
    1023.1, 1023.2, 1023.4, 1023.5, 1023.7, 1023.9, 1024, 1024.1, 1024.2, 
    1024, 1024.2, 1024.2, 1024.3, 1024.5, 1024.7, 1025.1, 1025.6, 1026, 
    1026.6, 1027, 1027.3, 1027.8, 1028.1, 1028.3, 1028.5, 1029, 1029.5, 
    1029.7, 1030.2, 1030.8, 1031.1, 1031.2, 1031.4, 1031.9, 1031.9, 1032.2, 
    1032.3, 1032.4, 1032.8, 1032.9, 1033.2, 1033.4, 1033.6, 1033.8, 1033.8, 
    1033.7, 1033.8, 1033.7, 1033.6, 1033.5, 1033.3, 1033.2, 1033.3, 1033.5, 
    1033.4, 1033.3, 1033.3, 1033.3, 1033.1, 1033, 1033.1, 1033.1, 1033.1, 
    1033.1, 1033.2, 1033.4, 1033.6, 1033.7, 1034.1, 1034.2, 1034.1, 1034.1, 
    1034.1, 1034.1, 1034.2, 1034.2, 1034.1, 1034.1, 1034.1, 1033.9, 1033.8, 
    1033.7, 1033.6, 1033.2, 1033.3, 1033.2, 1032.8, 1032.6, 1032.4, 1032.3, 
    1032.1, 1031.9, 1031.5, 1030.9, 1030.4, 1030.1, 1029.5, 1029.1, 1028.8, 
    1028.5, 1028.2, 1027.7, 1027.6, 1027.3, 1026.9, 1026.5, 1026.2, 1026.1, 
    1025.7, 1025.7, 1025.5, 1025.3, 1025.1, 1024.6, 1024.5, 1024.2, 1024, 
    1023.6, 1023.3, 1022.9, 1022.6, 1022.2, 1022, 1022, 1021.8, 1021.5, 
    1021.5, 1021.4, 1021.3, 1021, 1020.8, 1020.8, 1020.7, 1021.2, 1021.5, 
    1021.9, 1022.2, 1022.7, 1023.1, 1023.3, 1023.5, 1023.8, 1023.9, 1024.1, 
    1024.1, 1024.2, 1024.5, 1024.5, 1024.5, 1024.6, 1024.7, 1024.5, 1024.7, 
    1024.6, 1024.5, 1024.3, 1024, 1023.8, 1023.7, 1023.2, 1023.1, 1023.2, 
    1023.2, 1023, 1022.9, 1022.9, 1022.7, 1022.5, 1022.4, 1022.3, 1022.1, 
    1022.2, 1022.2, 1022, 1022, 1021.9, 1021.8, 1021.7, 1021.5, 1021.3, 
    1021.4, 1021.3, 1021.2, 1021.2, 1021.2, 1021.4, 1021.4, 1021.5, 1021.5, 
    1021.5, 1021.4, 1021.4, 1021.4, 1021.3, 1021.3, 1021.3, 1021.2, 1021.1, 
    1021.1, 1021, 1020.8, 1020.8, 1020.7, 1020.7, 1020.4, 1020.7, 1020.6, 
    1020.7, 1020.7, 1020.9, 1020.9, 1020.7, 1020.8, 1020.7, 1020.5, 1020.3, 
    1020.2, 1020.2, 1020.2, 1020, 1019.8, 1019.8, 1019.8, 1019.6, 1019.4, 
    1019.1, 1018.9, 1018.8, 1018.5, 1018.4, 1018.4, 1018.3, 1018.3, 1018.4, 
    1018.7, 1018.8, 1018.9, 1018.9, 1019, 1019.2, 1019.2, 1019.2, 1019.2, 
    1019.3, 1019.3, 1019.3, 1019.4, 1019.4, 1019.2, 1019.4, 1019.3, 1019.4, 
    1019.2, 1019.3, 1019.3, 1019.3, 1019.2, 1019.3, 1019.4, 1019.4, 1019.3, 
    1019.1, 1019, 1018.8, 1018.5, 1018.3, 1018.1, 1017.9, 1017.7, 1017.5, 
    1017.4, 1017.2, 1017, 1016.8, 1016.6, 1016.4, 1016.6, 1016.6, 1016.6, 
    1016.7, 1017.1, 1017.4, 1017.4, 1017.6, 1017.7, 1017.8, 1017.7, 1017.8, 
    1017.6, 1017.7, 1017.8, 1017.9, 1018, 1018.2, 1018.3, 1018.4, 1018.3, 
    1018.1, 1017.9, 1017.9, 1017.8, 1017.6, 1017.4, 1017.4, 1017.4, 1017.4, 
    1017.4, 1017.4, 1017.4, 1017.4, 1017.2, 1017.2, 1017.2, 1017.3, 1017.2, 
    1017.4, 1017.3, 1017.3, 1017.5, 1017.5, 1017.5, 1017.6, 1017.5, 1017.5, 
    1017.6, 1017.6, 1017.6, 1017.6, 1017.8, 1017.7, 1017.9, 1018, 1018.1, 
    1018.2, 1018.2, 1018.1, 1018, 1017.9, 1017.8, 1017.8, 1017.9, 1017.9, 
    1018.1, 1018.3, 1018.3, 1018.4, 1018.5, 1018.7, 1018.7, 1018.6, 1018.4, 
    1018.4, 1018.6, 1018.7, 1019, 1019, 1019, 1019, 1019, 1019, 1018.8, 
    1018.7, 1018.7, 1018.8, 1018.8, 1018.8, 1018.6, 1018.8, 1018.7, 1018.8, 
    1018.7, 1018.5, 1018.4, 1018.2, 1018.5, 1018.5, 1018.9, 1018.8, 1019, 
    1018.6, 1018.7, 1018.7, 1018.7, 1018.6, 1018.5, 1018.4, 1018.1, 1017.8, 
    1017.7, 1017.6, 1017.6, 1017.4, 1017.1, 1016.8, 1016.5, 1016.3, 1016.2, 
    1016.2, 1016.1, 1016, 1016.1, 1016.2, 1016, 1016.1, 1016.1, 1016.2, 1016, 
    1015.9, 1015.6, 1015.5, 1015.3, 1015.2, 1015, 1015, 1015, 1014.8, 1014.7, 
    1014.6, 1014.2, 1014.1, 1014, 1013.8, 1013.8, 1013.6, 1013.4, 1013.6, 
    1013.1, 1013.2, 1013.2, 1013, 1012.5, 1012.4, 1011.9, 1011.7, 1011.4, 
    1011.1, 1010.8, 1010.6, 1010.3, 1010.1, 1009.8, 1009.3, 1008.9, 1008.6, 
    1007.9, 1007.4, 1006.8, 1006.1, 1006, 1006, 1005.2, 1005, 1004.1, 1003.2, 
    1002.9, 1002.5, 1002.1, 1002.1, 1002, 1002, 1001.8, 1001.7, 1001.6, 
    1001.4, 1001.1, 1000.8, 1000.5, 1000.4, 1000.2, 999.7, 999.5, 999.2, 
    998.9, 998.7, 998.7, 998.5, 998.3, 998.3, 998.2, 998.1, 997.9, 997.8, 
    997.8, 997.7, 997.5, 997.6, 997.4, 997.1, 997, 996.9, 997, 996.9, 997, 
    997.1, 997.2, 997.4, 997.6, 997.9, 998.1, 998.5, 998.6, 998.8, 998.8, 
    998.9, 998.9, 998.8, 999, 999.1, 999.2, 999.3, 999.4, 999.4, 999.4, 
    999.2, 998.8, 998.5, 998.2, 998.1, 998.1, 998.1, 998.2, 998.3, 998.7, 
    998.8, 998.9, 999.2, 999.4, 999.5, 1000, 1000.2, 1000.6, 1000.6, 1001, 
    1001.4, 1001.7, 1002, 1002.3, 1002.6, 1002.8, 1002.8, 1003.1, 1003.4, 
    1003.8, 1004, 1004.1, 1004.4, 1004.9, 1005.2, 1005.5, 1005.7, 1005.9, 
    1006, 1006.2, 1006.4, 1006.6, 1006.9, 1007, 1007.2, 1007.4, 1007.6, 
    1007.8, 1007.9, 1008.1, 1008.2, 1008.5, 1008.5, 1008.6, 1008.8, 1009, 
    1009.1, 1009.3, 1009.4, 1009.5, 1009.5, 1009.5, 1009.7, 1009.7, 1009.6, 
    1009.8, 1010, 1010, 1009.8, 1009.8, 1009.8, 1009.6, 1009.8, 1009.9, 
    1009.7, 1009.6, 1009.6, 1009.4, 1009.1, 1009.1, 1009, 1008.8, 1008.5, 
    1008.2, 1007.9, 1007.5, 1007.3, 1006.9, 1006.5, 1006.1, 1005.4, 1004.9, 
    1004.2, 1003.6, 1003.3, 1002.7, 1002.3, 1002, 1001.8, 1001.4, 1001.3, 
    1001.4, 1001.2, 1001.2, 1001.6, 1001.5, 1001.7, 1002.2, 1002.6, 1002.9, 
    1003.4, 1004.1, 1004.8, 1005.2, 1005.8, 1006.4, 1007, 1007.7, 1008.4, 
    1008.8, 1009.7, 1010.1, 1010.4, 1011.1, 1011.6, 1011.8, 1012.4, 1012.9, 
    1013.4, 1013.8, 1014.2, 1014.6, 1015, 1015.2, 1015.3, 1015.4, 1015.5, 
    1015.7, 1015.8, 1015.9, 1016.1, 1016.2, 1016.2, 1016.2, 1016.3, 1016.4, 
    1016.3, 1016.2, 1016.3, 1016.3, 1016.5, 1016.5, 1016.7, 1016.8, 1017, 
    1017.1, 1017, 1017, 1017.2, 1016.5, 1017.1, 1017.5, 1017.7, 1017.8, 1018, 
    1018.5, 1018.4, 1018.5, 1018.5, 1018.5, 1018.6, 1018.8, 1018.9, 1019.2, 
    1019.3, 1019.5, 1019.4, 1019.5, 1019.6, 1019.5, 1019.7, 1017.2, 1018.3, 
    1018.7, 1019.1, 1019.3, 1019.8, 1020, 1020, 1019.9, 1019.8, 1019.8, 
    1019.7, 1019.5, 1019.3, 1019, 1018.6, 1018.4, 1018.3, 1018.2, 1018.1, 
    1017.9, 1017.9, 1017.9, 1017.6, 1017.4, 1017.3, 1017.2, 1017, 1018.8, 
    1017, 1017, 1016.8, 1016.9, 1016.8, 1016.8, 1016.8, 1016.7, 1016.6, 
    1016.6, 1016.8, 1016.9, 1017, 1017.7, 1018, 1018.2, 1018.4, 1018.6, 
    1018.7, 1019, 1019.2, 1019.6, 1016.8, 1017.3, 1019.9, 1020.3, 1020.8, 
    1021.1, 1021.5, 1021.8, 1021.8, 1021.9, 1021.7, 1021.7, 1021.8, 1021.9, 
    1022, 1021.8, 1021.7, 1021.8, 1020.5, 1020.1, 1020.6, 1021.2, 1021.7, 
    1022, 1021.8, 1019.3, 1018.5, 1018.4, 1017.7, 1017.5, 1016.7, 1015.7, 
    1015.3, 1014.8, 1014.3, 1013.2, 1012.6, 1011.9, 1011.1, 1011, 1010.6, 
    1010, 1009.6, 1009.3, 1008.8, 1008.5, 1008.2, 1008.1, 1018.7, 1013.7, 
    1007.7, 1007.6, 1007.6, 1007.6, 1008, 1008.4, 1008.6, 1008.7, 1008.6, 
    1008.4, 1008.1, 1007.9, 1008, 1008.3, 1008.7, 1008.9, 1009.2, 1009.6, 
    1009.9, 1009.9, 1010.1, 1010.1, 1010.5, 1010.6, 1010.6, 1010.7, 1010.8, 
    1010.6, 1010.5, 1010.5, 1010, 1010, 1009.6, 1009, 1008.7, 1008.2, 1007.5, 
    1007.2, 1006.6, 1006.4, 1006, 1005.8, 1005.4, 1005.2, 1005, 1004.6, 
    1004.5, 1004.4, 1004.2, 1004.6, 1004.5, 1004.2, 1004.4, 1004.4, 1004, 
    1003.6, 1003.6, 1003.5, 1003.3, 1003.3, 1003.4, 1003.4, 1003.2, 1002.9, 
    1002.8, 1003.5, 1003.6, 1003.9, 1003.8, 1003.9, 1003.5, 1004.2, 1004.3, 
    1004.8, 1005.1, 1005.4, 1005.8, 1006.2, 1006.2, 1006.6, 1006.8, 1006.9, 
    1007, 1007.1, 1007.6, 1007.9, 1007.9, 1008, 1008.1, 1008, 1008, 1007.9, 
    1008, 1007.9, 1007.7, 1007.2, 1007.4, 1007.8, 1007.6, 1007.5, 1007.4, 
    1007.4, 1007.3, 1007.2, 1007.1, 1007.1, 1007.1, 1007.1, 1007.4, 1007.4, 
    1007.3, 1007.3, 1007.9, 1007.8, 1007.4, 1007.4, 1007.4, 1007.3, 1007.1, 
    1007.2, 1007, 1007.4, 1007.3, 1007.3, 1006.6, 1006.7, 1006.5, 1006.4, 
    1006.3, 1006.6, 1006.3, 1006.1, 1006.1, 1006.4, 1007.1, 1006.4, 1006.7, 
    1006.2, 1006.3, 1006, 1005.7, 1005.4, 1005.1, 1004.9, 1004.7, 1004.5, 
    1004.4, 1003.5 ;

 wind_speed_10m = 3.6, 3.7, 3.6, 3.6, 3.5, 3.7, 4.7, 5.5, 3.9, 4.3, 4.1, 3.9, 
    4, 4, 3.8, 3.9, 4.2, 4.1, 3.3, 3, 4.6, 4.4, 4.5, 5.1, 5.7, 5, 4.2, 3.4, 
    3.9, 4.7, 5.4, 5.7, 4.3, 4.5, 5, 5.1, 4.9, 4.6, 4.7, 5.2, 5.1, 4.7, 4.5, 
    4.2, 4.8, 4.8, 4.8, 4.7, 4.7, 4.7, 4.6, 4.4, 4.2, 4.1, 4.4, 4.1, 3.2, 
    3.2, 3.2, 3.9, 3.5, 3.6, 3.5, 3.4, 3.3, 3, 3.1, 3.1, 2.6, 2.5, 2.4, 1.5, 
    2.2, 2.6, 2.4, 0.6, 1.4, 1.1, 0.3, 0.3, 0.6, 0.7, 1.9, 1.8, 0.8, 0.5, 1, 
    1, 1.3, 0.2, 0.2, 0.7, 0.7, 0.4, 1.3, 0.7, 0, 0.5, 0.3, 1.3, 4.9, 1.2, 1, 
    5.3, 5.4, 5.8, 5, 5.6, 3.7, 5.9, 5.6, 4.3, 2.7, 0.2, 0.4, 2.1, 0.8, 1.1, 
    0.8, 0.5, 1.2, 0.7, 1.1, 3.8, 3.2, 3.8, 4.7, 3.8, 1, 0.6, 4.7, 1.2, 0.4, 
    1, 0.5, 0.9, 1.4, 1.3, 0.6, 2.2, 1.8, 1, 1.9, 0.1, 1.2, 4.8, 4.7, 0.4, 
    1.4, 2.1, 2.6, 2.3, 3.1, 1.9, 2.1, 0.7, 2.3, 3.9, 3.6, 3.4, 3.5, 3.6, 
    3.4, 3.4, _, _, 0.5, 0.8, 1.4, 1.7, 0.1, 1.4, _, 1.5, 0.6, 0.6, 0.9, 2, 
    1, 1.9, 0.7, 0.9, 2.7, 1.6, 1, 1.5, 1.7, 0.5, 2, 1.1, 0.6, 1.5, 1, 4.4, 
    2.1, 2.3, 1.5, 1.6, 1.3, 1.6, 1.5, 6.7, 6.8, 6, 6.2, 8.5, 8.5, 5.5, 5.6, 
    7.1, 7.7, 7.7, 7.5, 6.7, 6.9, 6.7, 8.2, 8.1, 8.3, 7.6, 7.4, 7.2, 8, 7.6, 
    8.2, 8, 5.8, 2.8, 5.6, 6.2, 5.9, 7.8, 6.3, 6.8, 7, 6.2, 5.3, 6.7, 6, 6.4, 
    7.2, 6.1, 5.9, 6.8, 6.7, 6.5, 3.4, 5.4, 4.9, 3.5, 2.1, 3.3, 7.3, 6.6, 
    7.1, 6.8, 6.8, 6.9, 6.9, 7.5, 8.6, 8.3, 7.7, 7.5, 5, 2.6, 4.8, 4.5, 1.5, 
    1.4, 4.6, 3.5, 4.1, 4.5, 5.6, 4.7, 2, 1.2, 3.9, 2.6, 0.7, 0.7, 4.3, 5.5, 
    5, 3.9, 4.1, 5.5, 5, 5.1, 4.4, 4.4, 3.9, 3.2, 1, 4.6, 5, 4.8, 4.7, 4.9, 
    4.1, 3.4, 4.6, 4.7, 3.6, 4.8, 6.3, 5.2, 4.7, 4.5, 4.4, 4.9, 4.9, 2.4, 
    0.9, 0.9, 0.5, 0.4, 0.8, 0.4, 4.2, 2, 1.2, 1, 1.7, 1.2, 2.1, 1.5, 0.8, 
    0.4, 3.5, 2.1, 3.9, 4.5, 3.8, 6.4, 6.2, 4.5, 4.6, 3.6, 4.2, 2.9, 5.3, 
    5.7, 5.1, 4.6, 3.9, 3.7, 4.9, 4.3, 3.8, 0.9, 0.8, 0.5, 0.8, 1, 0.9, 0.9, 
    0.7, 1.8, 1, 1.3, 3.9, 0.9, 1, 0.2, 1.3, 0.3, 0.5, 0, 0.6, 1, 0.8, 0.8, 
    1.2, 1, 0.3, 1.2, 0.9, 0.3, 0.7, 1.5, 1.7, 3.3, 0, 0.4, 1.1, 0.7, 0.5, 
    0.4, 1.1, 1.4, 1.1, 1.2, 0.7, 1.6, 1.2, 0.7, 0.8, 0.5, 1.4, 0.5, 2.6, 
    0.8, 0.5, 1.5, 1, 1, 0.5, 2.9, 0.2, 0.5, 0.9, 0.8, 0.9, 0.1, 1.3, 0.5, 
    0.2, 2.4, 1.2, 1.5, 0.5, 0.2, 0.6, 0.1, 0.5, 0.7, 0.6, 0.2, 0.5, 0.7, 
    0.5, 0.5, 0.5, 0.5, 0.8, 1.1, 1.2, 0.8, 1, 0.6, 0.7, 0.9, 0.8, 0.6, 0.6, 
    0.5, 0.1, 0.2, 0.7, 0.9, 0.5, 0.8, 0.3, 1.6, 0.1, 0.3, 0.1, 1.2, 0.2, 
    0.4, 0.3, 0.9, 0.1, 1, 2.1, 0.6, 1.8, 2.6, 0.8, 0.7, 0.6, 3.3, 2.9, 0.6, 
    0, 0.6, 0.6, 0.5, 0.5, 0.9, 0.1, 0.3, 0.3, 0.9, 0.5, 0.4, 0.8, 1.6, 0.3, 
    3.4, 6.1, 7.4, 4.8, 4.7, 2.5, 2.4, 1.7, 1.9, 2, 1.3, 1.1, 1.4, 0.9, 2.1, 
    1.3, 1, 1.3, 0.4, 0.3, 0.8, 0.6, 0.6, 0.3, 0.8, 0.6, 0.2, 0.8, 0.8, 0.4, 
    0.8, 0.1, 1.1, 1.4, 0.5, 0.8, 2.6, 0.4, 0.9, 1.3, 0.7, 0.3, 1.1, 0.4, 
    0.8, 0.7, 1.1, 5.2, 6.5, 6.1, 5.6, 6.8, 7.5, 7.6, 5.9, 6, 7.1, 5.7, 5, 
    4.5, 2.7, 0.7, 5.5, 2.1, 0.3, 0.2, 6.1, 5.4, 0.8, 1.1, 1.3, 1.3, _, 1.3, 
    0.9, 1.4, 1.4, 0.6, 0.6, 0.1, 0.8, 0.5, 0.1, 0.1, 0.5, 0.5, 1.2, 0.7, 
    1.1, 0.8, 1.5, 1.8, 1.5, 2.8, 2.4, 1, 1.3, 2.6, 1.7, 0.6, 0.6, 0.3, 0.6, 
    1.1, 2.7, 2.1, 0.7, 1.2, 1.6, 2.9, 0.9, 1, 0.3, 0.8, 0.8, 0.2, 0.3, 1.6, 
    1.4, 0.7, 0.5, 0.3, 0.2, 1, 0.8, 1.6, 0.5, 1, 0.9, 0.4, 0.4, 0.9, 0.4, 
    0.3, 1.7, 0.4, 1.5, 0.5, 1.8, 1.2, 0.9, 0.3, 0.9, 1.4, 0.8, 0.6, 0.4, 
    0.8, 0.9, 0.4, 0.9, 0.5, 0.3, 0.4, 0.4, 0.6, 0.9, 0.8, 1.8, 0.5, 0.7, 0, 
    0.6, 0.5, 0.3, 0.5, 0.5, 0.4, 0.7, 0, 0.2, 0.3, 0.5, 0.7, 0.8, 0.8, 0.8, 
    0.4, 0.5, 0, 1.3, 0.6, 1.2, 0.6, 0.9, 0.6, 0.5, 1, 0.6, 0.9, 1.1, 0.6, 
    0.7, 1.1, 1.4, 0.7, 1.1, 2.2, 0.7, 1.2, 0.4, 1, 3.2, 1.7, 0.6, 1.7, 0.3, 
    0.9, 0.3, 0.4, 3.4, 0.3, 0.6, 1.2, 0, 1.4, 1.7, 1.8, 0.3, 0.2, 0.2, 0.1, 
    3.6, 4.7, 5.5, 5.6, 7.6, 9.8, 9.8, 9.7, 7.9, 6.5, 8.5, 6.9, 7.4, 7.8, 8, 
    8.1, 6.7, 8.1, 6.6, 4.5, 7.1, 3.7, 0.5, 1.4, 0.3, 1.4, 1.1, 0.9, 0.7, 
    0.2, 1.2, 0.6, 0.5, 0.6, 0.5, 0.2, 0.4, 0.9, 0.7, 1.3, 1.5, 1.1, 1.6, 
    1.7, 1.6, 0.9, 2.2, 0.3, 0.6, 1.5, 3.3, 2.2, 2.7, 8.3, 3.9, 1.7, 0.2, 
    0.3, 0.1, 0, 0, 1.7, 6.6, 4.6, 3.9, 4.9, 6.7, 5.4, 2.1, 6.7, 2.7, 0.5, 
    1.2, 0.9, 4, 1.3, 1.6, 2.5, 3.8, 0.4, 1.3, 2.4, 1.4, 0.8, 0.2, 0.2, 0.7, 
    1, 0.7, 0.6, 0.9, 0.6, 0.1, 1.4, 2.1, 1.9, 1.5, 1.1, 0.8, 0.2, 0.7, 0.1, 
    3.1, 0.4, 0.4, 1.1, 0.8, 0.6, 1.3, 0.9, 1.2, 1.8, 2.2, 2.6, 1, 1.2, 0.2, 
    1.2, 6.6, 6.4, 4.6, 4.3, 4.8, 5.5, 4.5, 10.7, 7, 4.9, 6.7, 5.6, 3.4, 5.4, 
    8.5, 7.2, 6.3, 6, 6.2, 5.3, 3.5, 5.6, 3.2, 7, 6.1, 5.4, 4.7, 5.7, 4.1, 
    2.9, 2.7, 1.8, 8, 2.4, 6.8, 6.1, 2.4, 5.4, 1.7, 1.1, 0.9, 0.8, 0.8, 0.3, 
    0.5, 0.5, 0.7, 1.5, 1, 1.4, 1, 1.8, 2.4, 1.3, 2.4, 2.1, 0.3, 0.5, 0.4, 
    0.8, 0.5, 0.3, 0.9, 1.1, 0.9, 1.1, 1.1, 0.4, 0.4, 1.5, 5.8, 6.1, 5.6, 6, 
    4.1, 4.4, 0.9, 2.2, 3.9, 6.4, 3.9, 3.3, 1.7, 3.3, 2, 1.1, 3.4, 2.7, 2.5, 
    3.2, 2.1, 1.1, 0.9, 0.8, 1, 2.1, 1.9, 2.6, 2.8, 1.8, 1, 1.4, 1.1, 1.2, 
    1.4, 0.8, 0.6, 3.9, 2.6, 0.8, 2.3, 1.2, 1.1, 0.4, 1, 5.7, 4.9, 5.4, 5, 
    5.2, 2.6, 2.8, 5.8, 7.8, 6.7, 7.8, 6.2, 6.4, 5.2, 3.5, 1.2, 3.6, 4.7, 
    3.9, 3.6, 3.9, 2.7, 1.7, 1.1, 0.7, 0.8, 1.3, 1.8, 1.5, 2, 2.2, 2.3, 2.5, 
    2, 1.4, 1.1, 1.1, 1.1, 0.2, 0.3, 1, 2.7, 3.9, 1, 0.5, 0.6, 0.4, 0.8, 1.4, 
    0.5, 0.9, 1.1, 0.2, 0.7, 0.2, 1, 0.8, 2.3, 0.6, 1.1, 0.1, 0.7, 0.5, 0.9, 
    1.3, 1.9, 2.1, 1.2, 3.7, 4.5, 2.6, 1.9, 2.5, 2.4, 2.5, 2.7, 1.2, 3.3, 
    2.4, 1.3, 1.5, 1.1, 2.1, 2, 3.4, 4.9, 4.3, 2.6, 2.2, 2.4, 2.3, 3, 2, 1.6, 
    1.7, 0.7, 0.7, 0.7, 0.6, 3.9, 0.7, 1.7, 1.1, 2.7, 2.9, 0.9, 1.4, 1.6, 1, 
    0.5, 3, 4.5, 6.2, 7.2, 8.8, 11.1, 11.2, 8.8, 6.3, 7.5, 7, 7.2, 9.6, 9.4, 
    9.1, 11, 10.9, 13, 13.5, _, _, 14.5, 14.9, 16.3, 15.3, 17, 17.6, 16.1, 
    15.2, 15.1, 14.4, 12, 12.6, 13.3, 14, 12.9, 13.5, 13.5, 13.1, 12.3, 11.3, 
    11.7, 11.2, 10.7, 10.7, 10.1, 9.6, 8.1, 9.5, 9.9, 8.5, 8.1, 6.8, 8.2, 
    8.3, 8.8, 8.3, 7.9, 8.8, 8.3, 8.1, 8.6, 7.5, 7.7, 6.5, 5.2, 2.6, 6.2, 
    5.6, 0.3, 0.5, 0.8, 3.2, 7, 7.3, 6.4, 6.3, 6.6, 6.3, 5.6, 6.5, 6.9, 6.8, 
    5.1, 4, 2.7, 4.9, 5.7, 5.4, 5.3, 4.5, 3.3, 3.9, 2, 3.6, 0.7, 0.2, 0.4, 
    0.2, 0.2, 0.7, 0.9, 0.1, 0.6, 1.1, 1.8, 0.9, 5.5, 7.2, 8.7, 5.9, 4.9, 6, 
    6.9, 4.9, 6, 5.6, 5.2, 4.1, 1.9, 0.2, 0.4, 0.5, 0.4, 0.9, 0.7, 1.7, 0.9, 
    1.2, 0.5, 1.7, 0.3, 0.2, 0.4, 0.8, 0.5, 1.5, 0, 1.3, 1.1, 0.6, 0.6, 0.1, 
    0.7, 1.6, 1.2, 1.3, 1.4, 0.2, 0.3, 1.2, 0.1, 0.4, 1.1, 0.4, 2, 3.7, 3.8, 
    2.6, 2.4, 3.8, 5.4, 7, 13.9, 13.7, 1, 1, 2, 2, 2, 3.3, 0.2, 0.9, 0.3, 
    0.7, 0.3, 0.8, 0.2, 0, 0, 0.6, 0.6, 0.4, 0.4, 4, 5, 6.7, 6.2, 5.9, 5.6, 
    5.1, 3.6, 4.7, 1.8, 1.5, 3.4, 5.6, 5.6, 5, 4.8, 3.4, 4.6, 3.2, 3.1, 2.9, 
    2.4, 2.6, 2.5, 0.9, 2.2, 2.3, 1.3, 0.1, 0.4, 1.3, 1.1, 0.4, 2.4, 0.8, 
    0.7, 0.5, 0.7, 0.4, 1.5, 0.9, 0.8, 0.9, 0.7, 1.3, 3, 1.7, 3, 3.7, 1.2, 
    2.5, 3, 2, 1.8, 1.8, 1.9, 1.8, 0.6, 0.3, 0.8, 1.1, 1.6, 1, 1.5, 0.4, 0.4, 
    0.2, 1, 1.5, 0.7, 0.8, 1.9, 0.6, 0.1, 0.9, 1.8, 3.4, 3.8, 3.3, 0.9, 3.8, 
    0.3, 0.2, 0.8, 4.9, 5.7, 6.2, 7.5, 4.8, 7, 7.6, 5.4, 5, 6.3, 6.5, 8.3, 9, 
    7.3, 6.7, 8.8, 7.6, 5.6, 5.9, 4.5, 8.6, 6.4, 4.4, 5.8, 6.5, 1.9, 5.2, 5, 
    3.1, 7, 6.5, 4.5, 4.8, 4, 5.2, 0.1, 0.2, 3.3, 1.1, 1.1, 2.8, 3.1, 1.3, 
    1.5, 0.4, 1, 0.9, 0.8, 2, 0.9, 1.4, 0.9, 2, 2.4, 3.9, 2.5, 2.2, 2.7, 2.3, 
    1.6, 2.6, 3.1, 2.7, 2.7, 1.9, 2.5, 1.7, 6, 2.8, 1.7, 4, 1.3, 1, 0.9, 0.7, 
    1.5, 0.6, 2.2, 0.7, 1.9, 1.7, 0.9, 1.2, 0.4, 1.3, 0.7, 0.9, 1.6, 0.6, 
    0.9, 0.8, 1.8, 0.7, 0.8, 0.8, 0.7, 0.3, 0.7, 0.7, 0.8, 1.1, 0.9, 0.7, 
    0.1, 0.3, 0.4, 0.6, 0.4, 0.2, 0.8, 0.1, 0.2, 3.2, 0.5, 0.7, 0.3, 1, 1.1, 
    1.2, 0.3, 0.5, 0.3, 1.2, 0.8, 1.1, 1.2, 1.6, 0.7, 0.7, 0.9, 1.4, 1.5, 
    2.1, 0.3, 6.5, 7, 7.1, 6.7, 6.6, 3.9, 6.1, 3.1, 1.3, 0.8, 0.6, 1.5, 4.8, 
    3.7, 2.5, 3, 3.4, 3.2, 2, 1.8, 1.7, 2.5, 1.6, 0.9, 2.6, 0.6, 1.9, 1.2, 
    0.6, 0.4, 0.3, 0.5, 0.7, 0.4, 1.8, 2.4, 4, 4.1, 1.3, 0.6, 0.8, 1.1, 5, 
    2.6, 4.7, 4.9, 5.2, 4.9, 3.5, 6.1, 4.7, 2.4, 1.3, 1.8, 1.2, 1, 0.5, 1.2, 
    0.6, 0.5, 0.7, 0.6, 2.1, 1.1, 0.9, 0.5, 0.6, 1.4, 0.1, 0.5, 0.6, 0.4, 
    0.3, 0.1, 0.8, 0.2, 1, 0.6, 1.9, 2, 1, 0.3, 0.2, 0.4, 0.6, 0.3, 1.3, 1.3, 
    1.3, 0.3, 0.9, 0.4, 0.1, 0, 0.1, 1, 0.8, 0.1, 1.8, 0.8, 0.6, 0.4, 0.3, 
    1.9, 2.9, 0.3, 0.8, 0.9, 0.7, 3.9, 3.5, 2.6, 6.7, 5.7, 4.9, 2.5, 0.4, 
    5.4, 3.7, 2.7, 6.5, 7.6, 7.1, 6.3, 7.5, 8.5, 4.9, 5, 7.5, 2.1, 6.6, 2.9, 
    3.2, 0.2, 1.7, 1, 2.3, 2.2, 2.6, 1.2, 1.2, 1.1, 1.9, 1.7, 2.6, 1.9, 1.3, 
    1.9, 0.4, 0.8, 1, 1.5, 0.9, 0.9, 2.2, 3.9, 1.6, 2, 2.6, 2.7, 3.1, 4.7, 
    1.1, 4.8, 1.8, 1.3, 0.6, 1.3, 1.4, 1.4, 3.6, 4.3, 5.8, 6.3, 5.1, 2, 1.6, 
    4.6, 4.3, 3.3, 3.5, 4, 4.3, 4.5, 3.6, 3.6, 2.3, 3.4, 0.6, 1.9, 1.3, 1.2, 
    0.7, 1.4, 1.7, 2.1, 0.8, 2.2, 0.8, 1.8, 2.1, 0.4, 2, 0.1, 1.7, 0.5, 1.5, 
    0.8, 1.4, 1.3, 0.9, 0.5, 0.9, 0.6, 0.5, 1.5, 2.2, 1.5, 0.4, 2.1, 1.7, 
    0.7, 2.1, 1.9, 1.6, 1.8, 1.7, 0.7, 1, 2.1, 0.6, 0.2, 0.9, 0.7, 1.9, 0.8, 
    1.4, 1.9, 1.1, 1.7, 2.3, 1.6, 0.9, 2.9, 2.7, 2.2, 1.8, 2.4, 1.7, 2.2, 
    1.6, 2.6, 0.8, 1.4, 1.5, 2.1, 0.3, 0.9, 0.7, 1.1, 1.7, 0.3, 1.4, 1.5, 
    0.7, 0.4, 0.9, 1, 1.2, 0.6, 0.7, 0.5, 0.5, 0.1, 0.5, 0.7, 0.7, 0.4, 0.7, 
    1.2, 0.5, 0.4, 0.6, 0.8, 0.1, 0.7, 0.5, 0.6, 0.3, 1.2, 0.7, 0.6, 0.5, 
    0.4, 0, 0.2, 0.6, 0.4, 0, 0.7, 0.8, 0.2, 0.4, 0.7, 0.9, 0.7, 1, 0.5, 0.1, 
    0.7, 0.5, 0.5, 0.1, 0.4, 0.5, 0.7, 0.2, 0.2, 0.5, 0.5, 0.9, 1.1, 0.2, 
    0.2, 0.5, 0.4, 0.6, 0.1, 0.1, 0.7, 0.2, 0.1, 0.5, 0.2, 0.4, 0, 1.7, 1.5, 
    0.6, 0.9, 0.9, 0.1, 1.5, 0.5, 0.6, 0.5, 1.7, 1.6, 0.4, 0.3, 2.3, 2.4, 1, 
    0.6, 0.6, 1, 2.8, 0.9, 0.7, 0.7, 0.9, 1.6, 1.3, 1.4, 1.1, 1.5, 2.2, 1.4, 
    0.5, 0.7, 1.7, 1.6, 1.4, 0.7, 3.2, 1.1, 4.9, 2.2, 4.4, 1.7, 5.5, 6.7, 
    5.2, 5.1, 5.5, 4.6, 5.2, 5, 3.8, 5.4, 4.8, 3.8, 3.9, 5.4, 4.3, 3.3, 3.5, 
    0.6, 0.8, 1.5, 0.3, 0.8, 0.9, 0.4, 0.5, 1, 0.6, 1.2, 0.7, 2.5, 2.3, 2.2, 
    1.9, 0.2, 0.9, 1.5, 0.3, 0.3, 0.2, 0.3, 1.1, 0.5, 0.1, 0.9, 0.6, 0.3, 
    0.9, 0.8, 0.1, 0, 0.9, 0.2, 0.5, 0.2, 0.4, 0.2, 0.1, 0.1, 0.8, 0.4, 0.1, 
    0.2, 0.4, 0.2, 0.5, 0.5, 0.2, 0.8, 0.4, 0.1, 0.4, 0.2, 0.5, 0.7, 0.1, 
    0.5, 0.1, 0.4, 0.3, 0.6, 0.6, 1.3, 0, 0.4, 0.4, 0.3, 0.3, 0.3, 0.6, 1.3, 
    0.8, 0.6, 0.7, 0.4, 1.5, 0.7, 0.3, 1.8, 0.4, 5.4, 4.3, 2.8, 1, 1.1, 3.1, 
    2.2, 1, 1.9, 1.8, 1.4, 0.8, 1.6, 1, 1.1, 1.4, 0.6, 1, 0.5, 0.6, 0.3, 0.4, 
    1.2, 1, 0.4, 0.9, 0.8, 0.8, 1.5, 1.2, 0.6, 1.6, 0.7, 0.4, 0.3, 0.7, 0.4, 
    0.9, 0.2, 0.4, 0.1, 0.6, 0.1, 1, 0.2, 0.2, 1.2, 0.4, 0.1, 0.5, 0.4, 0.7, 
    0.7, 1.3, 0.5, 1.3, 0.5, 0.8, 0.8, 0.7, 0.9, 1.2, 1.7, 1.4, 0.3, 0.8, 
    0.4, 0.6, 0.9, 1, 1.2, 0.3, 1.3, 0.7, 2.3, 0, 0.7, 1, 0, 1, 3.4, 0.7, 
    1.4, 1.5, 0.7, 0.6, 0.9, 0.6, 1.1, 0.4, 0, 0.5, 0.7, 0.2, 0.9, 0.2, 0.9, 
    0.5, 0.8, 1.2, 1.4, 0.1, 0.7, 0.1, 0.4, 0.2, 0.5, 1.2, 0.3, 1.1, 0.9, 
    0.1, 0.1, 0.2, 0.1, 0.6, 0.9, 5, 5.2, 4.6, 4.9, 3.3, 2.2, 2.5, 2.3, 0, 
    0.5, 3.2, 5.1, 3.7, 3.7, 2.4, 1.3, 0.1, 2.2, 2.1, 2.1, 6.1, 5.8, 4.9, 
    4.6, 1.6, 1, 0.4, 0.7, 3, 0.6, 0, 0.7, 1.4, 1.1, 1.5, 2.1, 0.9, 0.3, 0.6, 
    0.1, 0.5, 0.7, 0, 0.3, 0.9, 0.1, 0.1, 0.7, 4, 3.8, 2.4, 3.1, 1.1, 2.1, 
    0.6, 1.5, 0.2, 3.5, 3.5, 4.2, 1.4, 0.8, 0.2, 0.2, 0.4, 0.8, 2.4, 1.4, 
    0.8, 0.9, 0.6, 0.8, 0.4, 0.8, 6.1, 4.1, 5.4, 5.4, 4.5, 4.1, 5.5, 4.5, 
    2.8, 5.1, 4, 4.2, 3.7, 3.7, 4.4, 4, 0.8, 0.3, 1.1, 1, 0.2, 1.2, 0.7, 1.5, 
    0, 0.6, 0.8, 0.5, 0.9, 0.1, 0.5, 0.2, 0.3, 0.7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 0, 0, 0, 0, 1.7, 1.8, 2, 1, 3.8, 2.2, 4.1, 6.1, 1.9, 3.8, 
    8.1, 1.9, 2.4, 1.7, 1.1, 0.8, 1, 1.6, 0.8, 1.4, 0.6, 1.5, 0.9, 0.5, 0.9, 
    0.6, 0.2, 1.9, 3.1, 0.3, 0.3, 0.5, 0.7, 0.4, 1.2, 0.8, 3.6, 0.4, 0.8, 
    0.3, 1.7, 0.8, 0, 0, 0.7, 1.2, 0.5, 0.9, 0.6, 0.2, 0.5, 0.4, 0.2, 0.7, 
    0.2, 1, 1.2, 0.4, 0.2, 0.2, 0.1, 0.5, 0.3, 0.3, 1, 0.6, 0.8, 0.5, 0.8, 
    2.3, 2.8, 5.2, 5, 5.2, 4.1, 4.3, 4.7, 1, 4.8, 2.7, 2.3, 1.7, 1.4, 1.2, 
    0.3, 0.6, 0.3, 0.2, 0.4, 0.3, 1.6, 0.3, 0.8, 0.8, 0.1, 0.5, 0.7, 0.1, 
    1.1, 3.3, 2.1, 3.7, 2.6, 2.3, 1.1, 1.9, 0.1, 0.7, 0.7, 1, 0.4, 0, 0.6, 
    0.2, 0.1, 0.3, 2.3, 1.1, 3.3, 5.4, 4.8, 3.7, 3.7, 5, 5.2, 4.9, 4.2, 3.6, 
    2.4, 3.9, 3.4, 4, 5.2, 1.9, 2.2, 3, 2.7, 3.9, 2.8, 3.6, 1.2, 0.5, 2.8, 
    0.8, 0.9, 0.2, 0.6, 1.4, 0.6, 1.3, 0.9, 1.6, 1.5, 1.4, 0.5, 0.2, 0.7, 
    1.1, 0.4, 0.7, 1, 1.2, 2, 0.2, 0.8, 1.7, 0.1, 1.4, 1.5, 1.9, 4, 4.6, 4.7, 
    4.1, 7.8, 7.6, 5.8, 3.9, 4.1, 4.2, 4.7, 3.3, 3.2, 4.6, 3.4, 3, 5.8, 0.4, 
    4.4, 0.7, 1.1, 0.8, 0.3, 0.9, 1, 1.3, 0.6, 0.5, 0.3, 0.8, 0.4, 0.5, 0.7, 
    0.8, 0.6, 0.7, 1, 0, 0.1, 1, 0.7, 0.4, 0.5, 2.7, 0.7, 0.9, 0.5, 1.7, 1.3, 
    0.8, 0.6, 0.5, 0.3, 0.4, 0.6, 0.5, 0.6, 0.9, 0.5, 1.3, 0.7, 0.9, 0.6, 
    0.8, 0.1, 1, 0, 0.8, 0.8, 0.9, 0.2, 0.4, 5.1, 7.5, 7, 7.1, 6.8, 6.4, 5.4, 
    3.8, 2.7, 5.8, 5, 2.8, 1.9, 1.4, 1.2, 1.1, 1.4, 0.6, 1.7, 1.2, 0.6, 0.6, 
    0.7, 0.6, 2.2, 0.2, 0.7, 0.7, 0.3, 0.9, 0.9, 0.3, 0.4, 0.3, 0.6, 0.5, 
    0.3, 0.2, 0.7, 0.5, 0.6, 0.9, 1.2, 0.6, 1.1, 0.5, 0.5, 2, 1.5, 3.3, 7, 
    7.4, 7.7, 8.6, 8.1, 7.9, 7.9, 8.1, 7.9, 7.9, 7.4, 5.5, 6.5, 5.9, 4.3, 
    4.5, 2.7, 4.8, 1.3, 1.6, 2.2, 1.5, 1.8, 1.2, 1.1, 1, 0.9, 0.9, 0.2, 0.7, 
    0.6, 0, 0, 0.5, 0.1, 0.3, 0.6, 1.3, 0.7, 0.9, 0.5, 0.9, 0.5, 0.2, 1, 0.7, 
    0.2, 0.2, 1, 1.4, 0.1, 1.3, 0.5, 0.5, 0.1, 0.2, 0, 0.8, 0, 0.7, 0.9, 1.3, 
    1.6, 0, 1, 0.8, 0.7, 0.9, 1, 0, 0.7, 0.4, 1.4, 0.5, 0.5, 0.3, 0.2, 1, 
    0.9, 0.8, 1, 1.6, 0.4, 0.6, 3.4, 5.9, 2.4, 0.4, 1.3, 0.6, 0.4, 1.2, 1.5, 
    0.4, 0.6, 0.7, 0.5, 1.3, 0.7, 0.9, 0.5, 1.6, 0.6, 3.5, 3.5, 2, 1.9, 3.4, 
    3.2, 3.7, 1.7, 2.3, 0.9, 0.8, 1.3, 0.3, 0.6, 1.5, 0.4, 1.1, 1.3, 2.6, 
    2.6, 1.3, 1.4, 2.3, 0.5, 0.3, 1.1, 1.2, 1.9, 1.3, 1.6, 1.4, 9.8, 5.4, 
    3.7, 1.8, 4.5, 5.7, 4.2, 8.8, 8.4, 5.4, 4.3, 4.1, 3.1, 1.8, 2.2, 5.6, 6, 
    4.9, 5.9, 5.4, 1.7, 3.3, 2.7, 5.4, 6.2, 5.7, 6.3, 4.5, 2.8, 2.8, 3.4, 
    1.9, 1.1, 1.5, 1.4, 2.1, 0.5, 1, 1, 0.8, 1, 1, 2.3, 1.5, 1.3, 1.1, 1.6, 
    0.7, 1.2, 0.2, 0.8, 1.1, 0.9, 0.2, 1.1, 0.1, 0.4, 0.8, 0, 0.5, 0, 0.4, 
    0.2, 0.2, 0.3, 0.5, 0.3, 0.2, 0.2, 0.3, 0.2, 0.1, 0.9, 0.2, 0.8, 0.2, 
    0.7, 0.1, 1.2, 0.7, 0.2, 0.5, 0.3, 0.4, 0.3, 0.6, 0.8, 0.2, 0.2, 0.5, 0, 
    0.8, 0.2, 1.2, 4.5, 1.4, 0.6, 1.2, 0.5, 0.9, 0.5, 0.8, 0.6, 0.4, 0.7, 
    2.4, 1.3, 1.4, 1.1, 4.5, 2, 0.8, 1.7, 9.1, 9.6, 5.4, 2.6, 4, 4, 4.1, 4.1, 
    3.4, 3.2, 3.9, 3.6, 5.1, 7.1, 1.3, 7.8, 2.9, 1.3, 0.5, 0.5, 2.4, 7.1, 
    4.6, 3.3, 1.2, 1.6, 0.1, 1.6, 1, 0.4, 0.8, 0.6, 0.1, 1.4, 0.8, 0.7, 0.7, 
    0.9, 0.4, 0.9, 1, 1, 1.1, 0.9, 1.6, 0.2, 0.7, 0.7, 0.4, 1.4, 0.9, 1.3, 3, 
    0.6, 1.6, 2.4, 7.1, 3.6, 0.5, 3.9, 5.7, 4.4, 4.5, 4.5, 1.9, 2.7, 3.1, 
    0.6, 1.4, 1.9, 1.6, 0.7, 0.7, 1.1, 2.5, 0.6, 0.7, 0.7, 0.2, 0.8, 1.6, 
    0.9, 0.5, 0.6, 0.1, 0.2, 0.5, 0.1, 0.5, 0.5, 0, 0, 0.6, 0, 0.8, 0.9, 0.4, 
    0.2, 1, 1, 0.6, 0.7, 2, 1.2, 3, 2.2, 2, 1.9, 0.4, 1.9, 1.4, 1.6, 0.3, 
    0.2, 0.7, 0.7, 0.4, 0.7, 0.2, 0.8, 0.1, 0.2, 0, 0.6, 0.4, 0.2, 0.4, 0.9, 
    0.3, 0.9, 2.2, 0.8, 0.2, 0.1, 0.5, 0.4, 0.3, 1.2, 1, 1.7, 1.4, 1.5, 0.9, 
    1.2, 0.5, 0.4, 0.2, 0.7, 0.9, 0.5, 0.2, 0.5, 0.3, 0.5, 2.8, 0.4, 0.2, 
    0.6, 0.4, 0.4, 1.1, 0.7, 0.5, 0.3, 0.3, 1.1, 0.4, 0.1, 0.4, 0.5, 1.2, 
    0.7, 1.3, 1, 1.5, 1.4, 0.7, 0.5, 0.7, 0.9, 0.5, 2.3, 0.4, 0.9, 1.5, 0.4, 
    0.6, 0.2, 0.9, 1, 1.4, 1.3, 0.3, 1.4, 1.1, 0.2, 2.4, 4.8, 4.8, 1, 2, 5, 
    5, 5.1, 7, 6.9, 8.6, 8.1, 6.7, 7.4, 6.9, 6.3, 5.1, 3.7, 5.7, 4.2, 3, 4.8, 
    4.3, 4.1, 2.9, 5.4, 3.1, 6, 8.2, 7.1, 1.9, 4.4, 5.6, 3, 2.4, 4.4, 3.4, 
    1.2, 0.7, 0.5, 1, 1.9, 1.2, 3.3, 2.1, 2, 0.9, 1.2, 0.4, 0.5, 0.3, 0.7, 
    0.3, 0.5, 0.8, 0.2, 0.5, 0.1, 1.3, 0.2, 0.1, 0.3, 0.2, 0.5, 0.8, 0.4, 
    1.1, 1.2, 0.6, 0.2, 0.3, 0.5, 0.6, 0.2, 0.8, 0.3, 0.6, 0.2, 2, 0.4, 0.5, 
    1, 0, 0.3, 0.6, 0.1, 1.3, 0.2, 0.2, 0.3, 0, 0.6, 0, 0.5, 0.5, 0.3, 0, 
    0.5, 0.5, 0.3, 1.1, 1.5, 1.7, 1.8, 0.2, 0.2, 0.2, 0.6, 1.1, 0.6, 0.6, 
    0.9, 0.1, 0.6, 1.3, 0.9, 1.3, 0.8, 1.4, 1.5, 1, 1.4, 0.4, 1, 0.8, 1.3, 
    1.3, 2.5, 2.1, 2.8, 6.5, 10.2, 3.2, 2.7, 2.1, 8.3, 7.1, 8.5, 3, 4.9, 7.3, 
    6.8, 3.5, 5.2, 4.9, 2, 1.7, 1.1, 0.6, 2.9, 3.8, 1.8, 4.3, 5.1, 6.5, 2.2, 
    0.8, 2.5, 2.6, 2.2, 4, 2.1, 2.1, 4, 2, 1, 1.3, 0.6, 0.6, 0.4, 0.3, 0.4, 
    0.2, 1.4, 0.9, 0.5, 0.4, 1, 1.5, 1, 0.1, 0.5, 0.3, 0.7, 0.1, 0.1, 0.1, 
    0.1, 0, 0, 0.4, 0.2, 1, 0.2, 0.6, 0.5, 0.2, 0.9, 1.5, 2.5, 3, 0.5, 2.3, 
    1.3, 1.8, 2.5, 3.5, 4, 2.6, 1.7, 3.7, 2.4, 2.5, 1.7, 2.4, 2.9, 2.2, 2.1, 
    1.6, 2.3, 1.6, 2.1, 5, 4, 8.2, 8.2, 9.9, 9.8, 9.7, 10, 11.8, 8.1, 7.4, 
    7.4, 5.1, 7.8, 8.8, 5.8, 6.9, 6.6, 4.9, 5.3, 6.8, 7.2, 8.4, 10.2, 7.1, 
    7.7, 7.1, 7, 5.6, 4.2, 4.2, 4.2, 3.5, 0.2, 6.6, 5.1, 5.6, 4.5, 5.3, 5.5, 
    4.6, 5.4, 4.7, 0.6, 0.7, 1.5, 0.9, 1.1, 1.5, 0.4, 1.1, 0.9, 1.6, 0.3, 
    0.9, 1.1, 1.9, 0.8, 0.4, 1.5, 0.5, 1, 1.2, 0.1, 0.2, 0.9, 0.1, 0.3, 0, 
    0.3, 0.1, 1.2, 0.9, 1.6, 1.9, 1.9, 2.2, 0.7, 0.8, 0.2, 0.4, 0.9, 0.2, 
    4.5, 5.2, 4.4, 2.2, 1.1, 1.8, 1.6, 0.7, 0.1, 0.3, 0.1, 1.6, 1.6, 3.7, 
    1.4, 1.3, 0.7, 1.9, 0.6, 0.8, 0.9, 0.9, 0.7, 1.3, 1.2, 1, 0.5, 1, 0.6, 
    0.1, 0.3, 0.3, 0.2, 0.2, 0.6, 0.8, 0.4, 0, 0, 0, 0, 0.5, 0, 0.7, 0.4, 
    0.6, 0.8, 1.2, 0, 0.1, 0.6, 0.7, 0.3, 1.1, 1, 0.3, 0.3, 0.5, 0.3, 0.5, 
    0.6, 1.2, 0.3, 1, 0.5, 0.5, 0.4, 0.6, 0, 0.4, 0.1, 0.9, 0.7, 0.1, 0.7, 
    1.3, 0.3, 0.7, 0.2, 0.1, 2.6, 1.5, 1.3, 2, 2.1, 2.5, 0.6, 0.1, 0, 0.4, 
    0.7, 0.7, 0.3, 0.9, 0.6, 0.4, 1.1, 1.1, 0.6, 0.2, 1.8, 0.2, 0.5, 0.6, 1, 
    0.3, 0.9, 0.5, 1, 0.9, 0.7, 1.6, 3, 1.4, 2.5, 2, 1.8, 2.6, 1.5, 3.2, 2.5, 
    6.7, 7.5, 8, 6.7, 7.5, 8, 7.2, 4.4, 7, 9.5, 8.2, 4.9, 6.4, 6.7, 7, 1, 
    7.1, 2.2, 2.3, 7.5, 7.5, 8.7, 3.1, 3.4, 5.3, 6.5, 11.6, 10.2, 10.2, 9.5, 
    7, 2.2, 2, 2, 6.7, 1.4, 6.6, 2.2, 1.3, 2.8, 2.5, 1.7, 4.8, 0.9, 6.1, 3.5, 
    1.8, 3, 0.7, 3.7, 0.5, 4, 1.8, 2.5, 6.5, 7.5, 6.2, 5.3, 5, 5.9, 6.1, 7.7, 
    7.5, 8.1, 8, 9, 7.3, 5.7, 5.1, 1.6, 2.7, 1.6, 3.3, 2.8, 4.1, 1.2, 1.4, 
    4.6, 0.6, 1, 1.3, 1.9, 1.9, 3.8, 4.8, 1.2, 0.3, 0.8, 3.7, 0.9, 1.7, 2.9, 
    2.6, 1.1, 0.5, 0.6, 1.7, 3.7, 3, 4.7, 2.3, 5, 8.1, 7.1, 5.9, 2.9, 2.9, 
    2.3, 0.9, 1.3, 1, 0.6, 0.8, 0.8, 0.2, 0.3, 0.5, 2.1, 2.3, 3.3, 2.9, 3.2, 
    2.4, 2.7, 1.9, 1.6, 0.3, 0.8, 0.2, 0.7, 0.5, 0.3, 0.6, 0.2, 0.1, 0.2, 
    0.3, 0.1, 0.4, 0.6, 0.2, 0.1, 0.4, 1.4, 0.1, 0.4, 0.5, 1.3, 1.3, 1.2, 
    1.8, 1.1, 0.7, 3.8, 3.1, 3.7, 3.9, 0.8, 1.7, 1.3, 3.1, 1.4, 1.1, 1, 1.1, 
    1, 0.9, 0.5, 0.5, 0.8, 0.3, 0.6, 0.9, 0.2, 0.3, 0.4, 0.8, 1.1, 1.9, 0.6, 
    0.3, 0.1, 0, 0.3, 0.7, 0, 0.3, 0.3, 0, 0, 0.5, 1, 0.5, 0.3, 0.2, 0.1, 
    0.2, 0.7, 0, 0.5, 0.7, 0.3, 1.1, 0.1, 0.5, 0.1, 1, 1.5, 0.7, 0.8, 0.7, 0, 
    0.3, 0.3, 0.1, 0.2, 0.7, 0, 0.1, 0.5, 0.7, 0.9, 0.7, 0, 0.1, 0.5, 0.1, 0, 
    0.8, 0.6, 0.4, 0, 0, 0.4, 0.2, 0, 0.4, 0.2, 0, 1.1, 0.9, 0.4, 0.5, 0, 
    0.9, 0.4, 0.2, 0.2, 0.4, 0.8, 1, 0.4, 2.6, 0.9, 0.8, 0.8, 1, 0.9, 0.3, 
    0.7, 0.9, 1.2, 0, 1.3, 1.5, 1.5, 0.4, 0.5, 0.3, 0.2, 2.1, 0, 1.7, 0.2, 
    0.2, 0.2, 0.4, 1, 0.9, 0.2, 0.4, 0.3, 0.2, 0.3, 0.5, 0.6, 0.1, 0.2, 0.2, 
    0.7, 1, 0.1, 0.4, 0.5, 1.2, 1, 1.1, 0.4, 0.7, 0.1, 0.6, 0.2, 0.4, 0.6, 
    1.5, 2.8, 1.3, 0.6, 1.4, 1.5, 1, 1.2, 2.4, 3.5, 2.9, 1.6, 2.2, 2.4, 1.9, 
    0.7, 2.4, 1.6, 1.9, 1.2, 1.3, 1.4, 1.7, 1.1, 1.2, 1, 1.4, 0.9, 1, 1.2, 
    1.1, 0.9, 0.8, 1.6, 0.8, 0.9, 2.1, 0.7, 0.5, 0.1, 2, 0.7, 0.8, 0.4, 0.1, 
    0.5, 0.2, 0.2, 0.1, 0.3, 0.4, 0, 0.3, 0, 1, 0.5, 0.3, 1.1, 0.9, 0.8, 0.5, 
    1.2, 1.3, 1.6, 0.2, 0.1, 0.1, 0.2, 0.3, 0.5, 0.4, 0.2, 0, 0.5, 0, 0.5, 
    0.1, 0.1, 1.2, 0, 1.6, 1.2, 0.8, 0.2, 1.8, 0.6, 0.2, 1.4, 0.5, 0.4, 0.4, 
    0, 0.4, 0, 0.1, 0.9, 0.2, 0.3, 0.3, 0.1, 0.3, 0.1, 1.4, 0.3, 0, 0.4, 0, 
    1.4, 0.2, 0.7, 4.3, 5.2, 7.4, 7.4, 7.4, 8.4, 11.4, 10.1, 8.6, 7.5, 4.2, 
    1.8, 1.9, 1.5, 1.5, 0.7, 5.3, 0.8, 2.2, 3.6, 1.5, 0.7, 1.5, 3.5, 1.1, 
    1.4, 1.1, 0.7, 1.3, 3.5, 1.4, 1.7, 1.2, 1.5, 1.4, 1.1, 1.2, 2, 1, 0.8, 2, 
    2.2, 0.1, 0.4, 0.3, 0.8, 0.4, 0.8, 0.8, 2.3, 0.4, 0.1, 0.4, 0.6, 0.1, 
    0.5, 2.9, 1.8, 2.2, 1.7, 1.3, 2.2, 1.2, 1.5, 2.3, 2.3, 1.4, 0.9, 0.3, 
    1.1, 1.2, 0.6, 0.4, 0.9, 0.2, 0, 2.8, 0.2, 0.5, 0.3, 0.5, 0.4, 0.6, 0.4, 
    0.2, 0.2, 0.1, 0, 0.3, 0.2, 0.7, 0.7, 0.1, 0.8, 0.7, 1.4, 0.6, 0.4, 0.2, 
    0.6, 0, 1.2, 0.3, 0.2, 1, 0.2, 0.8, 0.8, 0, 0.1, 0.4, 0.5, 0.3, 0.2, 0.5, 
    0.3, 0.4, 0.1, 0.1, 0.2, 0.2, 0, 0.1, 0.4, 0, 0.3, 0.1, 1.2, 2.5, 3.5, 
    0.9, 0.4, 0.9, 2.8, 1.6, 1.7, 1.7, 1.5, 0.2, 0.8, 0.4, 1.5, 0.6, 0.4, 
    0.1, 0.6, 0.8, 0.4, 2, 1.2, 0.5, 1, 1.1, 1.2, 1.5, 2.7, 1.4, 2.3, 0.8, 
    2.8, 3.3, 3.4, 5.9, 2.3, 0.9, 1.5, 2.6, 1.1, 1.7, 0.9, 3.8, 1.5, 2, 1.8, 
    2, 1.2, 0.9, 1, 1.1, 0.4, 0.7, 1.6, 0.6, 2, 1.2, 0.9, 1.2, 1.4, 1.6, 1.3, 
    1, 0.3, 0.2, 0.6, 0.3, 1.3, 0.5, 0.5, 0.9, 0.7, 1.2, 1.1, 1, 0.3, 0.7, 
    0.1, 0.5, 1.1, 0, 0.9, 0.1, 0.1, 1, 0.5, 0.1, 0.5, 4.2, 0.8, 5.1, 7.3, 
    4.4, 7.1, 5.5, 4.5, 4.6, 5.4, 5.6, 7.4, 5.7, 5.5, 7.2, 7, 5.2, 3.6, 3, 
    4.6, 5.3, 2.5, 2.5, 3.2, 1.7, 1.4, 1.3, 0.5, 0.6, 1.3, 0.3, 0.5, 0.7, 1, 
    0.7, 0.2, 0.2, 0.2, 0.7, 0.1, 1, 1.5, 0.1, 0.3, 0.7, 0.6, 0.3, 0, 0.1, 
    0.4, 0.9, 0.1, 0.1, 0, 0.1, 0.1, 0.5, 0.8, 0.7, 0, 0, 1, 0, 0.9, 0.5, 
    2.4, 0.7, 1, 2, 1.3, 0.6, 0.4, 2, 2.1, 1.9, 2, 2.5, 2.8, 2.9, 2.6, 2.6, 
    2.5, 2.3, 2.7, 2.4, 0.8, 1.7, 0.2, 1.3, 0.4, 0.8, 0.6, 0.3, 0.2, 0.8, 
    0.3, 0, 0.4, 0.3, 1.1, 0.6, 0.3, 0.3, 1.8, 1.3, 0.7, 2.8, 2.4, 2.4, 0.8, 
    1.5, 2.1, 3.2, 5, 5.2, 4.3, 5.2, 2.5, 5.4, 2.2, 3.9, 1, 1.1, 0.3, 2.6, 
    4.1, 1.3, 0.2, 1, 1.1, 1, 1.7, 1.8, 1.8, 2.3, 2.2, 2.3, 1.3, 2.4, 2.3, 2, 
    2.6, 1.4, 1.6, 1.8, 0.1, 0.1, 0.3, 0.8, 1.5, 1.3, 1, 1.6, 2.2, 3.5, 1.8, 
    2.7, 2.2, 0.9, 1.1, 1.2, 5.1, 5.5, 5.2, 5.3, 3.4, 6.6, 6, 4.5, 3.1, 2.2, 
    3.4, 0.4, 2.1, 0.6, 1.3, 1.8, 1.1, 1.6, 2.1, 2.3, 0.1, 2.1, 1.5, 1, 2.1, 
    1.5, 1.4, 0.7, 0.7, 3.3, 5.5, 4.8, 3.5, 3, 3.4, 3.6, 3.3, 3.2, 1.4, 0.8, 
    2.6, 1.8, 0.5, 0, 2.3, 1.8, 2.5, 2.5, 2.3, 2.2, 1.9, 1.1, 0.3, 0.2, 0.4, 
    0.4, 0.1, 0, 0.8, 1.6, 0.8, 1.1, 0.7, 0.6, 1, 1, 1.3, 1.7, 1.5, 1.2, 2.4, 
    2.7, 1.9, 0.9, 1.2, 0.3, 1.3, 1.1, 0.1, 2.1, 1.9, 2, 0.2, 0.1, 0.8, 0.4, 
    1.2, 0.4, 0.9, 0.1, 0.7, 0.9, 1.9, 1.5, 1.5, 1.5, 1.1, 4, 4.4, 3.3, 2.6, 
    3.7, 3.3, 2.7, 2.6, 3.3, 0.4, 0.3, 0.2, 0.3, 0.7, 0.4, 0, 0.1, 0.4, 0.5, 
    1.9, 1.7, 1.7, 1.8, 0.5, 0.2, 0.9, 1.3, 1, 1.4, 1.2, 0.5, 0.1, 0.3, 1.1, 
    0.4, 0.5, 0.4, 1.3, 0, 0.8, 2, 1.1, 0.2, 1.6, 1.8, 1.1, 1.7, 1.3, 0.8, 
    1.4, 0.8, 1.1, 2.3, 0.9, 1.7, 0.8, 1.1, 1.5, 2, 0.8, 2, 2.5, 2.4, 1.7, 
    1.2, 0.9, 1.5, 2.5, 2.6, 2.1, 1.6, 0.6, 0.2, 0.8, 1.5, 1.7, 0.5, 1.1, 
    0.5, 1.7, 1.5, 2.2, 2, 1.5, 0.6, 0.7, 1.2, 2.3, 2.7, 1.5, 1.9, 2, 1.6, 
    1.5, 1, 0.6, 1.6, 1.6, 1.3, 1.6, 1.8, 1.7, 1.8, 2.3, 1.5, 0.9, 0.2, 1.3, 
    0.2, 0.3, 2.5, 2.2, 2.2, 1, 2.4, 1.6, 2.5, 1.3, 0.4, 1.3, 0.5, 1.3, 1.2, 
    1.6, 1.3, 0.6, 1.1, 2.3, 1.6, 0.9, 0.7, 3.2, 1.3, 0.2, 1.8, 1.2, 1.6, 
    0.3, 2.2, 1.1, 0.7, 0.3, 0.3, 0.6, 4.7, 6.4, 7.3, 6, 5.8, 6.4, 5.5, 6.1, 
    6.7, 5.6, 5, 5.5, 4.4, 1.5, 0.8, 3, 1.4, 1.2, 2.6, 2.4, 0.5, 0.2, 0.3, 1, 
    1, 0.7, 1.3, 0.5, 1.6, 0.8, 1.1, 0.5, 3.4, 1.6, 2.8, 3.1, 0.4, 0.5, 1.2, 
    0.5, 1.3, 1.2, 1.5, 1.3, 1.5, 3.3, 3.1, 2.9, 2.9, 2.5, 1.6, 1.7, 1.1, 3, 
    2.7, 3.2, 3.3, 3.7, 3.5, 3.1, 2, 1.5, 2.3, 1.4, 1.5, 4, 3.6, 3.4, 0.4, 
    1.1, 4, 0.4, 1.2, 0.7, 0.7, 1, 1.2, 2.8, 2, 2.8, 0.9, 1.1, 0.6, 0.9, 0.2, 
    0.2, 0.1, 0.8, 0.9, 1.4, 1.1, 0.3, 0.2, 0.2, 0.2, 2, 1.3, 0.9, 0.9, 0.9, 
    0.8, 2.1, 2.3, 1.9, 2.8, 1.4, 2.1, 1.9, 2.3, 2.2, 1.5, 1.4, 1.5, 0.9, 
    1.1, 2.3, 1.2, 2, 3.6, 3.7, 3.5, 4, 3.6, 3.9, 3.6, 2.5, 4.4, 3, 3.4, 2.7, 
    1.3, 2.5, 3.2, 2.4, 3, 0.6, 0, 1.1, 0.7, 0.7, 0.2, 0.5, 0.7, 0.6, 0.5, 
    1.6, 2.8, 2.1, 1.2, 2.8, 0, 1.7, 1.1, 0.6, 0.5, 0.1, 0.8, 0.6, 0.3, 1, 
    1.1, 0, 1, 1, 0.5, 0.3, 0, 0.1, 0.1, 0.7, 0.1, 0.3, 3.4, 4.3, 6.2, 7, 
    9.8, 8, 9, 10.1, 10.8, 9.5, 8.4, 8.5, 8.3, 8.2, 8.2, 8.2, 7.8, 8, 7.8, 
    6.7, 6.3, 6, 6.8, 6.8, 3.1, 5.3, 3.2, 3.3, 1.3, 3.7, 3.7, 2.9, 1, 1.6, 
    0.2, 0.8, 0.1, 0, 0.2, 0.9, 0.5, 0.8, 1.4, 2.7, 1, 0.4, 1.4, 1.1, 1.1, 
    1.1, 1.8, 0.8, 0.5, 0.2, 0.2, 0.3, 0, 0.1, 0.3, 0.6, 0.2, 1.1, 0.7, 1.5, 
    0.9, 1.2, 0.9, 0.9, 1.4, 1.7, 1, 1.7, 1.3, 0.1, 1.1, 0.9, 1, 0.2, 0.7, 
    0.3, 1.5, 0.5, 0.4, 0.8, 0.4, 1.5, 1.9, 2.2, 2.3, 2.1, 1.5, 1.1, 0.9, 
    0.7, 1.1, 1.4, 0.5, 0.3, 0.6, 2.9, 0.2, 0.3, 2.1, 0.9, 2.7, 2.9, 1.6, 
    6.3, 5.2, 4.6, 4.2, 4.6, 4.3, 4.9, 5.1, 3.9, 2.4, 3.2, 1.6, 1.2, 1.7, 
    2.7, 1.3, 1.1, 0.5, 0.3, 0.3, 0.2, 0.9, 0.7, 0.4, 0, 0.9, 1, 2.5, 1.9, 
    1.2, 2.7, 2.6, 0.1, 0.4, 0, 0.9, 0.3, 1, 0, 0, 1.2, 0.6, 0.2, 1.2, 0.4, 
    0.5, 0.2, 0, 1.3, 2.4, 0.2, 0.5, 0.3, 1.2, 0.7, 1, 0.2, 1, 0.3, 0.8, 0.9, 
    0.9, 1.5, 0.3, 2.8, 0.3, 0.1, 0, 2.2, 2.2, 1.7, 0.6, 2, 0.6, 1.9, 0.8, 
    1.8, 0.8, 1, 0.4, 1.2, 0.7, 1.9, 2.3, 2.5, 2.8, 3.7, 2, 1.6, 0.1, 0, 0.8, 
    0.6, 0, 0.6, 0.1, 1, 1.4, 0.5, 0.5, 0.9, 1.2, 1.1, 0.8, 1, 0.7, 0.8, 1.1, 
    4.3, 0.7, 0.3, 1.1, 0.4, 0.7, 0.2, 0.2, 0.6, 0.1, 0.5, 0.3, 0.3, 0.8, 
    1.4, 3.5, 6.2, 1.9, 1.3, 0.9, 0.4, 0.3, 1.3, 0.3, 1.4, 0.4, 1, 3.6, 4.6, 
    0.6, 1.6, 4.5, 4, 5.1, 6.7, 6.5, 5.4, 4.1, 5.9, 8, 4.9, 6.5, 6.3, 7.1, 
    6.3, 6.6, 6.8, 4.8, 5.8, 4.3, 5.9, 6, 5.6, 3.7, 0.2, 0.1, 0.1, 0.5, 1.6, 
    0.6, 0.8, 6, 3.9, 5.5, 3.4, 5.7, 5.8, 6.8, 5.2, 7.7, 6.5, 6, 5.9, 6.1, 
    6.4, 3.1, 4.6, 2.8, 3, 3.5, 3.2, 2.9, 3, 3.2, 2.7, 4.7, 3.4, 1.9, 1.5, 
    2.2, 1.5, 4.2, 4.9, 5.9, 4.5, 1.5, 1.7, 3.4, 3, 2.4, 3.9, 3.2, 2.4, 0.5, 
    0.9, 1.7, 0, 2.3, 5.6, 5.2, 4.9, 6, 6.2, 5.3, 6.6, 7.5, 4.3, 6.1, 3.9, 
    5.6, 1.2, 2.9, 2.9, 2.7, 3, 0.1, 2.3, 2.5, 2.5, 3.2, 3.4, 3.7, 4.6, 3.8, 
    3.4, 4.9, 4, 3.9, 4.9, 4.9, 4.2, 3.6, 5, 4.1, 5.1, 4.6, 4.8, 4.2, 5.5, 
    3.1, 2.9, 2.5, 3.5, 4.5, 3.4, 4.6, 3.9, 3.1, 4, 3.3, 2.7, 3.3, 3.2, 2.3, 
    0.4, 2.9, 1.4, 3.6, 3.5, 2.9, 3, 2.1, 4.2, 4.9, 5.7, 6.7, 3.3, 5.6, 3.3, 
    2.5, 3, 1.8, 1.9, 1.1, 2, 2.9, 2.1, 2.9, 3.1, 4.1, 4.5, 5.1, 4.6, 5.6, 
    5.4, 4.4, 5.4, 2.2, 0.8, 3.4, 0.4, 0.7, 1.7, 0.8, 0.3, 1.6, 2.4, 2.2, 
    1.6, 2.1, 1.6, 1.6, 2.6, 2.2, 3.5, 3.6, 4.6, 4.1, 4.1, 4.2, 5.2, 3.9, 
    3.9, 3.2, 3.9, 4, 4.8, 4.6, 4, 4.3, 3.8, 2.6, 1.5, 1.4, 3.6, 3, 1.8, 2.6, 
    2.7, 5.3, 7.2, 6.8, 6.7, 4.6, 7, 7.4, 2.3, 6.2, 5.9, 0.7, 2.6, 1.7, 2.6, 
    3.2, 2.7, 3, 2.9, 4.4, 4.3, 3.7, 6, 6.2, 7.2, 6.5, 7.2, 6.5, 7.3, 6.7, 
    5.8, 4.8, 5.3, 5.7, 5.4, 5.6, 5.6, 5.8, 6, 5.1, 5.8, 5.9, 6.2, 4.9, 3.7, 
    5.3, 4.6, 5.4, 4.8, 4.5, 5.8, 6.5, 7, 6.6, 5.3, 4.8, 5.2, 4.8, 2.7, 0.8, 
    1.7, 0.8, 1.7, 3.1, 5.7, 5.4, 4.1, 1, 2.8, 4.9, 1.1, 3.6, 2.7, 3.4, 3.2, 
    1.8, 2.8, 2.8, 2.2, 3.4, 2, 1.7, 0.8, 0.5, 1.7, 1.9, 0.7, 2.4, 2.3, 3.4, 
    4, 5.3, 5.4, 5.9, 4.5, 5.3, 4.3, 4.4, 3.4, 3.7, 4.5, 4.9, 5.5, 5.1, 5, 
    5.3, 4.5, 5.3, 4.1, 3.8, 4.3, 4.3, 4.6, 4.4, 5.4, 4.6, 5.2, 5.6, 5.1, 
    5.5, 6.1, 6.5, 4.7, 4.1, 4.4, 4.1, 4.4, 4.4, 4.7, 5.5, 5.1, 4.8, 4.5, 
    3.1, 3.9, 4.3, 3.3, 2, 1.5, 1.6, 0.3, 2, 3.7, 1.3, 1.4, 0.5, 4.3, 3.9, 4, 
    4.7, 4.8, 5.3, 5.9, 5.2, 4.6, 3, 1.6, 0.6, 2.2, 0.4, 1.4, 0.1, 0.3, 0.5, 
    0.4, 3.7, 4.1, 3.5, 3.3, 2.8, 1.4, 2.2, 0.4, 1.6, 1.7, 4.1, 1.1, 1.4, 
    0.8, 1, 1.7, 1.2, 0.4, 0.2, 0.2, 1.7, 1.5, 1.4, 0.6, 1.2, 1, 1.7, 2.6, 
    1.9, 2, 1.6, 3.4, 1.1, 1.8, 1.6, 1, 0.6, 1.6, 0.8, 0.3, 1, 0.6, 0.4, 1, 
    0.4, 1, 1.7, 1.3, 1.4, 1.7, 1.3, 1.9, 1.4, 0.7, 1.6, 4, 2.7, 1.3, 0.1, 
    1.2, 0.2, 0.3, 0.9, 0.8, 1.1, 1.8, 0.2, 2.7, 1.2, 1.4, 1.2, 1.6, 2.4, 
    4.3, 3.2, 3, 2.9, 4.7, 2.3, 1.8, 2.7, 2.9, 2.5, 0.6, 0.3, 0.8, 0.2, 0.5, 
    1, 1, 1.2, 0.7, 0.5, 1.7, 2.3, 3, 1.3, 1.2, 1.1, 4.4, 5.3, 5.8, 3.9, 5, 
    4.2, 4, 4.9, 3.5, 5.4, 4.6, 4.4, 5.4, 6.5, 5.5, 5.9, 6.7, 5, 4.7, 5.5, 
    3.9, 3.3, 3.8, 2.9, 5.2, 4.5, 3.6, 3.3, 3.4, 3.6, 3.7, 3.3, 2.6, 1.8, 
    1.8, 1.4, 2.9, 1.5, 1.1, 0.2, 2.7, 2.3, 2.3, 1.9, 3.2, 3.9, 2.9, 2.9, 
    2.2, 2.6, 2.4, 2.5, 2.9, 3.1, 2.6, 3.1, 1.4, 0.4, 3.1, 1.4, 2.5, 1.5, 
    2.7, 3.4, 3.9, 4, 3.5, 2.5, 2.1, 1.7, 1.9, 0.4, 0, 1.2, 0.6, 6.3, 4.9, 
    5.2, 5.8, 4.7, 3.5, 0.5, 1.1, 1.2, 3.4, 4.4, 3.1, 4.2, 2.4, 3.5, 3.8, 
    4.4, 4.4, 5.5, 5.8, 4.9, 4.9, 4, 4.7, 3.3, 5.8, 4.5, 5, 4.7, 3.8, 3.7, 4, 
    1.4, 0.8, 2.9, 4.1, 1.3, 3.8, 6.4, 5, 5.2, 3.7, 2.7, 3.4, 2.5, 2.8, 2.6, 
    1.4, 2.2, 2.6, 0.5, 0.5, 0.9, 1.7, 0.5, 0.8, 0.7, 0.1, 0.5, 0.9, 0.2, 
    0.3, 0.6, 1.2, 0.6, 2.4, 2.1, 2.4, 2.9, 1.5, 2.2, 1.5, 3.6, 3.3, 1.7, 
    1.1, 0.2, 0.7, 0.7, 0.3, 1.1, 1.3, 2.2, 0.8, 1.9, 0.6, 0.2, 0.7, 1.2, 
    0.7, 0.7, 1.4, 2, 1.7, 4.4, 0.7, 1.7, 2.8, 8, 7.4, 5.8, 5.3, 4.6, 4.1, 
    2.1, 0, 1.9, 0.1, 1.1, 1.1, 1.3, 0.4, 0.3, 0.1, 0.3, 1.4, 0.3, 1.1, 1, 
    1.8, 0, 1.6, 1.9, 1, 0.8, 0.6, 4.7, 3.5, 4.8, 3.1, 0.1, 0, 1.5, 0.5, 1.1, 
    1, 0.9, 1.9, 1.5, 0.8, 1.5, 0.3, 1.6, 0.9, 1.3, 1.7, 0.3, 2.2, 0.5, 0, 
    0.2, 0.4, 0.5, 1.3, 0.7, 0.7, 0.1, 0.5, 0.2, 0.8, 2, 1.1, 1.9, 3.9, 4.5, 
    3.9, 4.9, 4, 2.7, 5.6, 1.7, 3.4, 2.1, 2.3, 1.6, 0.3, 5.5, 3.3, 3.7, 1.5, 
    1.7, 0.7, 2.7, 0.3, 0.5, 1.4, 1.7, 2, 3.1, 2.4, 2.7, 3.7, 4.7, 3.4, 2.9, 
    1.6, 1.3, 0.7, 1.5, 1.4, 1.6, 0.8, 0.4, 0.6, 0.9, 1.8, 1.2, 2, 1.6, 1.6, 
    0.4, 0.5, 2.3, 0.8, 2.1, 1.2, 0.3, 0.4, 1.2, 1.8, 0.9, 1.7, 0.1, 0.4, 
    0.7, 0.8, 0.7, 0.6, 0.6, 0.9, 0, 0.2, 2.2, 2.2, 2.1, 1.5, 1.4, 0.6, 5.3, 
    0.2, 1.9, 3.3, 4.3, 1.4, 0.9, 2.5, 2.5, 0, 0.2, 0, 0.5, 0.3, 0.9, 0.6, 
    2.8, 1.2, 0.4, 3.6, 2.6, 1.7, 0.8, 2.8, 3.3, 0.3, 0.5, 0.9, 2.4, 3.1, 
    2.1, 3, 1.5, 0.7, 1.7, 1.1, 1.3, 0.7, 0.2, 0.9, 0.8, 0.7, 1.3, 1.7, 1.7, 
    1.7, 2.1, 2, 2, 1, 1.5, 2.1, 2.1, 1.8, 1.5, 1.4, 0.8, 0.8, 1.7, 1, 1.2, 
    0.4, 0.4, 0.2, 0.7, 3, 0.7, 0.9, 1.5, 2, 2.2, 3.4, 2.6, 4.6, 3.7, 4.3, 4, 
    4.3, 4, 5.2, 5.4, 5.2, 4.7, 3.9, 3, 3.2, 2.1, 0.9, 2.3, 2.1, 1, 0.4, 4.6, 
    3.5, 4.7, 5, 2.7, 2.1, 2.4, 5.1, 5.1, 6.5, 3.5, 2.3, 4.3, 2.2, 2.6, 2.5, 
    4.8, 5, 2.1, 1.7, 3.6, 2, 1.1, 2.2, 1.4, 7, 5.7, 0.8, 0.9, 4.1, 4.2, 2, 
    3.8, 2.4, 0.8, 0.3, 0.3, 0.2, 0, 0.2, 0, 0.4, 0.7, 0.4, 0.6, 3, 2.3, 3.1, 
    3.1, 2.9, 2.8, 3.2, 0.4, 1, 0.9, 2.6, 0.5, 0.7, 0, 0.7, 0.4, 0.7, 0.1, 
    0.8, 0.6, 0.2, 1.4, 0.1, 1.7, 3.7, 3.9, 4.4, 4.9, 0.5, 4.8, 4.2, 1.2, 
    4.4, 1.3, 1.3, 1.4, 1.8, 2, 0.5, 0.5, 0.9, 0.8, 0.3, 0.2, 1.8, 0.3, 2, 
    2.8, 4.2, 5.1, 3.2, 6.7, 6.2, 3, 6.8, 3.3, 3.8, 2.6, 2.7, 2.3, 5, 2.5, 
    4.6, 5.1, 5.8, 5.7, 3.2, 2, 4.4, 2.2, 4.9, 2.2, 1.6, 3.3, 1.5, 2.1, 0.8, 
    1.8, 1.1, 5.8, 2.6, 1.9, 2.9, 1.1, 2.5, 2.5, 4.4, 5.4, 5.2, 4.1, 2.4, 
    3.3, 3.6, 3.8, 4.5, 3.6, 3.5, 4.2, 0.9, 2.3, 2.7, 2.1, 1, 1.8, 4.4, 1.6, 
    4.2, 0.4, 2.4, 0.6, 1.3, 3.6, 1.6, 0.4, 0.7, 1.3, 0.7, 1.5, 2.1, 2.9, 
    2.1, 3.5, 3.1, 2.6, 2.4, 2.7, 2.4, 2.5, 1.9, 2.1, 0.6, 0.8, 1, 0.4, 0, 
    0.2, 0, 0.7, 0.1, 0, 0.6, 0.6, 1.4, 0.7, 1.1, 1.7, 1.7, 1.9, 2.2, 2.1, 
    2.4, 1.5, 1.8, 1.7, 1.7, 1.1, 1.4, 1.5, 1.5, 1.1, 0.8, 0.6, 0.5, 0.5, 
    0.7, 1, 2, 1.3, 1, 1.7, 1.8, 3.3, 0.7, 1.7, 5, 1, 6, 4.2, 4.5, 4.7, 3, 2, 
    2.1, 2.9, 4.1, 5.4, 5.4, 4.5, 5, 6.8, 7, 3.7, 5.2, 5.9, 4.2, 1.1, 1.2, 
    1.9, 1.2, 2.2, 2.1, 1.9, 2.1, 1.5, 1.1, 1.4, 2.3, 1.2, 1, 0.8, 1.1, 0.9, 
    0.4, 0.1, 1.7, 1.3, 2.3, 4.1, 3.1, 3.5, 4.4, 3.6, 2.6, 5.4, 5.4, 4.5, 
    5.3, 5, 4.7, 6, 4, 3.6, 2.6, 2.4, 3, 4.3, 4.9, 4.8, 4.3, 2.8, 1.7, 2.3, 
    7.5, 6.5, 5.5, 8, 6, 7.8, 5.4, 4.8, 5.6, 3.8, 3.2, 5.2, 4.1, 3.7, 3.1, 
    3.4, 2.8, 2.5, 1.4, 3.8, 3.6, 2.8, 1.5, 2.6, 2.2, 2.3, 2.9, 2.1, 2.6, 
    2.1, 1.5, 2.5, 2.2, 2.1, 2.4, 1.7, 0.7, 2.9, 1.7, 1, 1.9, 2.4, 1.4, 1.6, 
    2, 1.5, 2.9, 2.9, 3.1, 3.9, 2.3, 0.6, 3.2, 2.6, 2.1, 2.1, 1.9, 1.5, 1.4, 
    1.2, 0.9, 0.3, 0, 0.3, 0, 2.6, 0.2, 0.5, 3.1, 1.5, 3, 3.7, 4, 3.7, 2.6, 
    3.1, 2.9, 3, 2.5, 5, 4.8, 2.8, 3.3, 1.7, 3.4, 3.1, 0.7, 0.5, 3.1, 3.2, 
    1.8, 1.4, 1.2, 1, 1.1, 1.7, 2, 2, 2.1, 2.2, 1.2, 1.1, 0.4, 1.2, 2.2, 1, 
    0.4, 1.3, 0.5, 1, 2, 2.8, 2.7, 2.1, 2, 2.7, 1.9, 1.4, 2.3, 1, 2.2, 1.5, 
    3, 2.7, 1.8, 2.6, 3.6, 1.8, 3.9, 3.6, 3.4, 2.9, 2.8, 2.8, 2.5, 3.2, 1.6, 
    2.7, 3.1, 2.5, 2.3, 0.8, 1.6, 1.7, 1.9, 1.7, 1.9, 1.6, 1.2, 1, 0.7, 0.6, 
    0, 0.1, 0.3, 0, 0.6, 1.4, 0.2, 0.3, 0.3, 0.8, 3.1, 0.4, 1.4, 2.5, 3.5, 
    1.7, 1.8, 2.6, 3.1, 1.5, 1.8, 2.8, 0.5, 1.7, 0.8, 1.6, 1.1, 1.9, 0.5, 
    0.4, 1.9, 1, 0.2, 0, 1.8, 1.5, 1.5, 0.2, 1.7, 0.2, 1.3, 0.5, 1.5, 1.5, 
    1.3, 1.7, 1.5, 2, 1.4, 0.2, 0.4, 1.5, 1, 1.7, 1.2, 1.3, 0.5, 0.5, 1.3, 
    0.3, 0.1, 0.8, 0.5, 1.1, 0, 1.2, 0.4, 0.8, 1.2, 1.4, 1, 0.7, 0.6, 1.2, 
    1.9, 0.9, 1.2, 1.3, 0.8, 1, 1.9, 0.9, 1.4, 0.9, 0.1, 0.4, 0.9, 0.8, 1.2, 
    3.2, 1, 2, 2.1, 0.1, 1, 1, 0.7, 0.3, 0.1, 0.3, 0.8, 1.3, 1, 0.1, 0.4, 
    0.6, 0.8, 0.2, 1.2, 0.1, 0.1, 0, 1.2, 0.6, 0, 1.5, 1.1, 1.6, 1.1, 0.9, 
    0.2, 0, 1.2, 1.5, 2.6, 2.2, 1.8, 0.9, 1, 1, 0.6, 0.4, 0.6, 0.8, 1, 0.7, 
    2, 2.6, 3.1, 1.5, 1.6, 1.5, 1.5, 1.9, 2.3, 1.9, 1.6, 0.8, 1.6, 1.3, 1.4, 
    0.4, 1.7, 0.4, 0.9, 2.5, 1.8, 1.8, 1.8, 1.8, 2, 2.3, 1.6, 1.5, 1.8, 1.9, 
    1.1, 1.6, 1.5, 1.9, 2.1, 1.4, 1.1, 1.9, 1.8, 2.7, 3.8, 1.8, 0.9, 1, 3, 
    0.8, 1.1, 1.2, 1.2, 2.5, 2.8, 3.1, 2.7, 2.4, 2, 1.2, 1.7, 0.1, 2.3, 1.5, 
    0.7, 0.9, 0.4, 0.4, 1.2, 1.1, 0.4, 1, 0.9, 0.4, 0.1, 0.8, 1.4, 1.4, 1.4, 
    1.8, 1.8, 1.9, 2, 1.6, 1.5, 0.8, 1.9, 0.2, 0, 0.3, 0.1, 1.4, 0.3, 0.5, 
    0.2, 0.8, 0, 1, 0.2, 0, 1.5, 0.5, 0.3, 2.7, 0.5, 1.3, 1.3, 0.2, 0, 2.3, 
    3.2, 2.6, 1.5, 1.6, 0.7, 0.6, 0.9, 0.1, 1, 0.6, 1.9, 0.9, 1, 0.5, 0.8, 
    1.6, 1.6, 1.1, 0.6, 1.3, 3.2, 2.9, 0.8, 1, 0.6, 0.3, 0.1, 0.1, 0, 1, 1, 
    0.9, 1, 0.9, 1, 0.8, 2.3, 2.3, 3.9, 3.4, 3.7, 2.6, 1.6, 0.9, 1.6, 1.9, 
    1.9, 2, 1.1, 0.6, 1.7, 4.8, 4, 4.1, 3.9, 4, 4.1, 6, 2.5, 1.5, 3.9, 3.4, 
    4.6, 3.9, 5.2, 3.8, 4.4, 3.2, 6.6, 3.2, 2.2, 3.8, 1.7, 0.4, 2.7, 1, 2, 
    0.1, 0.8, 1.1, 0, 2.5, 3.3, 4.3, 5.4, 5.4, 4.2, 5.5, 5.2, 4.1, 3.6, 4, 
    4.3, 3.8, 4.9, 5.3, 5.2, 3.9, 1.5, 1.4, 2.7, 4.2, 3.7, 2.9, 3, 3.4, 3.7, 
    0.8, 1.1, 0.7, 2.5, 1.1, 0.6, 1.7, 2.1, 1.8, 0.6, 1.3, 1.2, 0.6, 1.3, 
    0.2, 1.8, 1.5, 1.9, 2, 1.3, 1.5, 1.4, 1.5, 2.1, 1.9, 0.5, 0.5, 0.4, 0.6, 
    2.1, 2.8, 0.9, 2, 0.7, 2.2, 2, 3.1, 3, 1.1, 0.9, 0.9, 0.7, 2.7, 0.7, 2.6, 
    2.1, 1.6, 0.8, 1.5, 1, 1.8, 3, 1, 2.9, 0.1, 2.4, 2.5, 3.4, 2.5, 1.7, 2, 
    2.3, 0.9, 6.1, 5.1, 5.8, 6.7, 4.1, 3.9, 2.5, 3.2, 4.1, 1.4, 1, 1.8, 0.8, 
    0.2, 1, 0.2, 0, 0.5, 0.4, 1.2, 1.6, 0.3, 0.1, 0.6, 0.5, 0.1, 0, 0, 1.1, 
    0.5, 0.8, 0.9, 1.3, 0.2, 0.6, 0.1, 0.2, 0.1, 0.1, 3.9, 0.3, 0.7, 0, 0.8, 
    0.8, 1, 0, 1.1, 1.6, 0.8, 0.2, 0, 0.5, 0.6, 2.3, 1.1, 0.1, 0.7, 1, 0, 
    0.7, 0.3, 0.3, 0.8, 0.8, 0.9, 3.8, 2.8, 3.3, 3.2, 2.4, 3.3, 2, 1.8, 0.4, 
    1.5, 2.1, 2.3, 3.7, 6.3, 5.1, 3.9, 6.6, 6.7, 7.6, 7.3, 6, 8.1, 7.8, 6.5, 
    4.6, 2.9, 1.4, 3, 0.6, 0.1, 0.4, 0.7, 1.4, 1.1, 0.4, 1, 1.2, 0.2, 0.5, 
    0.7, 1.8, 1.1, 1.7, 0.6, 1.7, 1.1, 2.9, 4.5, 1, 0.9, 1.5, 0.1, 3.1, 2.2, 
    0.8, 0.8, 1.6, 0.3, 0.3, 0.3, 1.1, 1.4, 0.6, 0.3, 0.9, 0.8, 0.9, 0.5, 
    1.4, 3.4, 4.5, 4, 0.8, 1.4, 3.9, 3.1, 3.9, 3.3, 4.6, 3.8, 3.9, 3.1, 1.4, 
    1.9, 0, 0.9, 0.9, 0.3, 0.2, 5.2, 0.9, 0.8, 0.9, 2, 2.7, 4.2, 4, 1.4, 1.2, 
    0.6, 1, 0.1, 0, 0.3, 0.6, 0.5, 0.4, 0.2, 0.4, 0.3, 0.6, 1.3, 1.6, 1.3, 
    1.7, 1.7, 1.8, 2.5, 1.9, 1, 0.9, 2.5, 2.1, 2, 1.8, 0.7, 0.9, 1.5, 0.6, 
    0.6, 1.6, 0.6, 0.1, 0.8, 1.6, 1.4, 1.6, 1.6, 4.3, 2, 3.9, 4.6, 3.4, 1.6, 
    1.1, 0.5, 0.7, 1.8, 2.1, 1.3, 2, 0.5, 0.5, 0.6, 0.7, 0.6, 0.4, 0.6, 0.6, 
    0.1, 1.3, 1.7, 1.9, 1.6, 0.7, 1, 1.3, 1.8, 2.4, 2.9, 2.5, 1.3, 1.9, 0.8, 
    1.2, 1.5, 1.2, 2.6, 0.5, 0.8, 1.4, 2.7, 2.4, 1.7, 2.9, 2.3, 1, 1.2, 1.2, 
    2.9, 2.1, 1.4, 0.8, 1.3, 1.6, 1.9, 0.1, 0.9, 0.5, 0.2, 1.2, 0.9, 0.6, 
    0.5, 1.3, 0.5, 1.7, 0.7, 0.3, 1.1, 7.9, 1.2, 0.4, 0.6, 0.9, 6.9, 7.9, 
    6.4, 8.3, 7.4, 6.9, 7.4, 7.3, 7.6, 6.5, 6.3, 5.1, 5, 5.3, 4.9, 6.2, 6, 
    5.6, 5, 3.2, 4.1, 3.8, 3.7, 4.4, 4.4, 4.8, 3.5, 3.7, 3.7, 3.6, 4.2, 4.2, 
    3.4, 3.4, 4.1, 4.5, 3.1, 3.1, 0.5, 0.2, 0.5, 2.2, 3, 2.9, 5, 3.4, 4.1, 
    4.4, 3.7, 4.4, 4.6, 5, 4.9, 3.5, 3.5, 3.7, 2.8, 3.7, 1.9, 3.3, 2.6, 1.4, 
    2.4, 2.4, 2.3, 2.5, 1.9, 3.1, 2.7, 2.3, 2.1, 5.7, 2.9, 3.4, 3.6, 4.1, 
    3.9, 2.6, 2.1, 1.6, 3.1, 5.3, 2.1, 2.2, 0.9, 2.2, 1.5, 1.6, 2.4, 2.5, 
    1.5, 3.3, 2.3, 6.3, 3.1, 3.7, 5.5, 1.9, 2.2, 0.9, 0.4, 0.3, 2.8, 1.1, 4, 
    5.2, 4.6, 4.7, 4, 2.6, 3.8, 3.3, 2.9, 3.5, 1, 3.5, 3.6, 3.8, 1.7, 1.1, 
    2.3, 4.2, 3.5, 3.8, 4.7, 0.9, 0.6, 0.5, 0.1, 0, 1.5, 0.6, 0.8, 1, 1.3, 
    0.8, 0, 0, 0.3, 0.3, 1.4, 1, 1.4, 1.6, 1.6, 1.6, 1.5, 1.5, 1.2, 1.2, 1.1, 
    1.6, 1.8, 2.1, 0.1, 2, 2.6, 1.7, 1.3, 2.1, 1.8, 0.4, 1.3, 1.3, 1.4, 0.9, 
    1.8, 1.8, 1.2, 1.9, 1.9, 1.7, 0.4, 1.1, 0.2, 0.1, 0.3, 0.7, 1.1, 1.3, 
    1.6, 0.3, 0, 0.1, 1.7, 2.3, 3.8, 2.7, 1.6, 0.9, 0.6, 0.8, 0.4, 1.4, 1.8, 
    0.4, 0.5, 0.7, 0.5, 0.8, 4.4, 2.8, 4.7, 0.9, 4, 1.9, 2.9, 0.6, 0.2, 0, 
    0.9, 5.2, 1.4, 1.4, 2.5, 3.4, 3.9, 2.4, 0.7, 0.8, 2.2, 0.8, 0.9, 1.6, 
    3.5, 0.5, 6, 0.9, 0.8, 2.5, 3.2, 2.4, 2.7, 2.5, 3.7, 2.6, 5.6, 2.5, 4.4, 
    3.2, 4, 2.6, 3.8, 3, 4, 3.5, 2.7, 3.6, 4, 3.3, 3, 3.8, 3.7, 4.8, 3.7, 4, 
    7, 6.4, 6.1, 6.1, 6.4, 6.1, 6.4, 7.1, 5.1, 4.8, 4.6, 4.9, 3.9, 4.2, 4, 
    7.4, 6.1, 5, 3.3, 3.3, 4.5, 6, 5.4, 4.9, 5.1, 6.2, 4.4, 6.2, 4.7, 4.5, 
    5.3, 4.2, 3.5, 2.4, 2.9, 2.1, 0.3, 0.7, 1.2, 0.7, 0.6, 1.6, 1, 2.3, 1.5, 
    0.6, 0.1, 0.6, 1, 0.2, 1, 1.8, 2.1, 0.7, 2.3, 3.7, 2.7, 2.7, 3, 3.6, 2.9, 
    4.2, 4.2, 4.7, 4, 3.7, 3.1, 2.1, 1.2, 0.5, 0, 0, 0.1, 3.6, 0.1, 0.1, 1.3, 
    0.8, 1.1, 2.3, 3.6, 4.1, 5.5, 4.9, 2.6, 1.1, 3.2, 4.1, 1.2, 0.3, 0.6, 
    2.2, 2.2, 0.2, 0.2, 0.6, 0.5, 0.3, 2.9, 3.8, 3.6, 3.4, 4.9, 5.8, 6.2, 
    6.1, 5.3, 6.2, 5.6, 2.6, 0.7, 1.4, 2.5, 0.9, 1.9, 2.6, 1.8, 1.7, 1.2, 
    1.2, 0.7, 2.4, 0.6, 1.8, 2.1, 2.3, 2.2, 2, 1.6, 1.4, 1.1, 0.5, 0.4, 0.2, 
    0.6, 0.9, 1.2, 1.9, 1, 0.8, 0.2, 3.2, 0.1, 1, 0.9, 0.8, 2.9, 3, 0.3, 2.2, 
    0.6, 1.7, 2.1, 1.5, 1.2, 5, 1.7, 1.4, 0.9, 1.1, 0.4, 0.2, 1.4, 0.8, 0.5, 
    4.4, 2.8, 4.5, 4.7, 5.5, 4.9, 7.4, 5, 5.8, 7.2, 7.2, 7.7, 8.2, 6.5, 4.3, 
    6.3, 3.3, 4, 2, 2.1, 0.3, 1.9, 1.4, 2, 0.9, 1, 2.8, 2.7, 6.3, 3.2, 5.6, 
    3.3, 1.8, 2.5, 2.9, 2.2, 0.6, 0.8, 1.4, 0.3, 0.9, 0.8, 3.3, 2.6, 0.9, 
    2.2, 0.5, 2.4, 1.8, 0.4, 0.4, 0.4, 0.1, 0.1, 0.6, 0.4, 0.6, 0.2, 0.5, 
    0.2, 0.1, 0.6, 0.1, 0.3, 0.1, 0.6, 0, 0, 0.6, 0.2, 0.2, 0, 0.7, 0, 0.1, 
    1, 0.8, 0, 1.6, 0.4, 0.1, 0.1, 0.3, 0.9, 0.9, 0.7, 0.3, 0.8, 0.4, 0.1, 
    0.1, 0.4, 1.5, 0.3, 3.4, 1.3, 1.1, 1.2, 0.6, 0.4, 3.5, 1, 3.4, 1, 0, 0.1, 
    0, 1.1, 0.5, 2.8, 0.3, 0.5, 1.1, 1.6, 1, 1, 0.2, 3.1, 0.1, 0.8, 0.9, 0.6, 
    2.6, 0.3, 2.4, 0, 0, 0.4, 0.2, 0.1, 0.1, 0.1, 1, 0.3, 1.4, 0.3, 0.1, 1.2, 
    1, 0.9, 1.4, 0.3, 0.3, 1, 0, 0.1, 0.3, 0.6, 0.5, 0.3, 4, 0.9, 0.7, 0.9, 
    0.8, 0.6, 0.2, 0.3, 0, 1.1, 0.8, 0.2, 0.8, 0.4, 0.6, 0.6, 0.4, 0.1, 0.4, 
    0.3, 1.4, 0.6, 3.1, 3.1, 0.4, 0.2, 0.6, 0.6, 0.4, 4.1, 2.2, 5.4, 4.4, 
    5.3, 5.3, 4.1, 4.7, 4.5, 1.8, 1.6, 1.3, 0.9, 0.8, 2.5, 0.4, 2, 0.8, 3.4, 
    5, 5.3, 5.4, 5, 4.7, 5.2, 4.4, 5.8, 6.9, 5.7, 4.4, 5.7, 6.7, 6.1, 6, 5.4, 
    5.6, 7.1, 6.6, 6.4, 6.3, 7.1, 7.4, 8.2, 7.7, 7.7, 7.2, 1.1, 1.7, 2.1, 
    2.9, 4, 2.5, 2, 0.8, 1.8, 1.5, 0.1, 1.7, 0.2, 0.9, 1, 4.3, 1.3, 2.1, 0.9, 
    2.4, 2.5, 1, 1, 0.6, 0.2, 1.6, 0.8, 0.6, 0.6, 0.1, 1.1, 0.3, 0.2, 0.7, 
    0.3, 0, 0.1, 0, 0.2, 0.1, 0.6, 2.3, 0.1, 0, 0.2, 0, 0.5, 0.7, 0.1, 0, 
    0.6, 2, 1.3, 1, 1.6, 0.3, 0.7, 0.1, 1.1, 0.6, 0.6, 1.2, 0.4, 0.2, 0, 0.4, 
    0.7, 0.2, 0.9, 0.4, 1.1, 0.8, 1, 0.6, 1, 1, 3.1, 0.7, 0.4, 0.9, 0.9, 0.3, 
    0.1, 0.6, 0.1, 0.6, 0, 0, 0, 0, 0, 0, 0.2, 0.4, 0.1, 0.4, 0.1, 0.5, 0.7, 
    0.9, 0.3, 0.4, 1.2, 0.2, 0.1, 0, 0.6, 0.3, 0, 0.3, 0.7, 0.5, 0.3, 0.4, 
    1.2, 3.2, 0.7, 0.1, 0.3, 0.9, 0, 1.1, 1.2, 1.7, 1.8, 0.9, 0.1, 0.4, 1.2, 
    0.2, 0.9, 0.8, 0.5, 4.1, 0.2, 0, 0.7, 0.4, 0.9, 0.6, 0, 4.1, 4.4, 4.3, 
    4.2, 4.3, 3.9, 4.4, 3.9, 4, 4.3, 4.4, 4.2, 3.9, 4.3, 4.4, 4.4, 4.8, 4.5, 
    5.4, 5, 4.9, 5.1, 5.3, 5.1, 4.7, 4, 0.8, 2.1, 1.5, 0.9, 0.4, 0.6, 0.4, 
    1.6, 1.2, 0.4, 0.6, 4.8, 0.9, 0.7, 1.4, 1.1, 0, 1, 0.1, 0.8, 5.6, 0.4, 
    1.4, 0.4, 0.7, 6.8, 1.5, 1.7, 0.5, 0.6, 2.9, 1.5, 1.3, 0.3, 1.9, 1.5, 
    1.8, 0.7, 1.1, 1.6, 0.8, 1.5, 5.2, 2.4, 1.3, 1.3, 0.8, 1.9, 1.4, 3.5, 
    1.2, 4.2, 3.2, 4.5, 3.2, 3.5, 4.6, 3.1, 4.5, 2.4, 4, 2.4, 2.6, 3.1, 1.6, 
    1.9, 2.9, 2.5, 0.7, 2.3, 6.2, 2, 0.7, 1.8, 0, 4.5, 4.2, 4.9, 3.7, 4.2, 
    3.7, 4.8, 3.1, 6.8, 6.3, 5.2, 5.3, 4.9, 4.9, 4.9, 4.9, 2.3, 4.4, 2.9, 
    3.1, 4.4, 3.9, 3.5, 4.5, 4.7, 2.3, 2.7, 2.5, 4, 4.5, 3.8, 2, 3.6, 1.4, 
    1.2, 0.6, 1, 0.7, 0.5, 1.1, 1.1, 0.5, 1.3, 1, 0.8, 1.2, 0.9, 0.4, 1.5, 
    1.7, 0.7, 0.4, 0.9, 0.9, 3.4, 0.9, 2, 1.8, 7.7, 4.9, 3.2, 5, 2.9, 4.8, 
    5.7, 6.6, 2.7, 2.1, 1.7, 1.1, 1.7, 2.5, 1, 1, 0.6, 1, 0.6, 2.9, 1.7, 2.9, 
    4.2, 3.8, 4.1, 4.3, 3.7, 5, 6.7, 5.7, 6, 6.7, 7.4, 6.6, 8.6, 7, 7.4, 8.3, 
    8.1, 6.4, 6.6, 7.4, 5.9, 9, 8.5, 7.7, 8.3, 5.6, 8.6, 8.3, 7.5, 7.7, 8, 
    8.2, 7.2, 5.9, 6.9, 7.5, 6.4, 6.4, 5, 5.6, 4, 4.4, 4.9, 4.1, 3.5, 4, 5, 
    2.8, 1.7, 3.3, 0.6, 3.2, 2.6, 0.7, 1.1, 0.9, 3.7, 3.8, 0.3, 0.1, 0.5, 
    0.3, 1.9, 3.1, 3.4, 2.8, 3.7, 3.8, 3.5, 3.4, 3.6, 3.7, 3.5, 2.4, 2.8, 
    3.2, 4.2, 2.1, 2.5, 2.8, 2.4, 1.2, 0.8, 1.2, 0.3, 0.6, 1, 0.6, 1.1, 0.6, 
    2.7, 5.5, 2.6, 3.2, 3.2, 4.5, 6.4, 3.9, 3.4, 2.9, 4.8, 0.6, 0.7, 0.7, 
    0.9, 0.2, 0.2, 0.6, 0.6, 2.3, 2.5, 0.4, 0.8, 0.6, 2.7, 1.3, 0.8, 0.6, 
    0.6, 0.6, 1.1, 1.1, 2.2, 1.8, 1.2, 4.4, 6.9, 3.2, 2.7, 4.9, 5.8, 5.6, 
    8.3, 3.1, 2.3, 4.6, 4.3, 4, 3.3, 3.6, 4.5, 2.2, 2.5, 0.9, 1, 0.4, 1.4, 1, 
    1.8, 2.3, 1, 2.4, 1.3, 3.1, 0.6, 0.9, 0.6, 1.3, 0.5, 0.5, 0.9, 2.2, 0.7, 
    1.1, 1, 1.6, 1.1, 1.3, 1.4, 0.6, 1.1, 0.5, 0.7, 1.5, 0.7, 1.3, 0.7, 1.9, 
    1, 0.3, 0.8, 1.6, 2, 0.5, 1.1, 0.7, 0.3, 1, 1.5, 0.1, 0.9, 0.6, 1, 2.1, 
    0.8, 1.1, 1.3, 1.2, 0.8, 1.5, 0.3, 4.3, 8.2, 7.1, 8, 8.9, 7.7, 8.5, 8.7, 
    7.1, 7, 7.8, 8.4, 7.9, 4.6, 2.6, 3.6, 3.5, 3.1, 2.3, 3, 3.1, 2.6, 3.4, 
    1.2, 3.4, 0.8, 1.4, 0.4, 0.7, 0.4, 1.3, 0.9, 0.8, 1.2, 1.1, 1.3, 0.4, 
    1.1, 0.9, 0.6, 0.5, 1, 0.1, 0.8, 1.5, 0.5, 1.4, 0, 0.6, 0.8, 1.4, 1.2, 
    0.1, 1, 1.3, 1.3, 0.6, 0.6, 3.7, 3, 2, 2.2, 3.5, 2.8, 2.1, 2.9, 0.3, 5, 
    5, 4.7, 4.7, 5.4, 4.3, 3.4, 2.2, 3.9, 1.3, 1, 1.8, 3.2, 1.5, 2.1, 3.7, 
    6.4, 6.4, 7.9, 7.3, 5.5, 2.6, 7, 6.4, 6.3, 7.5, 5.9, 8.5, 7.5, 7.4, 5.9, 
    6.9, 6.4, 1.6, 2.6, 1.5, 3.6, 4.1, 4.5, 1.4, 1.4, 1.2, 1.1, 0.4, 0.5, 
    0.3, 0.7, 0.7, 0.3, 0.6, 2, 0.7, 1.5, 1.2, 0.7, 0.6, 0.3, 0.7, 0.7, 0.6, 
    1.4, 1, 0.3, 0.8, 0.3, 0.7, 0.8, 0.5, 0.7, 3, 0.9, 1.6, 1.4, 1, 0.6, 2.3, 
    1, 1.4, 0.6, 0.1, 1.2, 0.3, 1, 1.9, 1.3, 1, 0.8, 0.9, 1, 0.6, 0.8, 0.6, 
    1.1, 0.6, 0.8, 0.8, 1.3, 0.8, 1, 0.5, 0.1, 0.7, 0.9, 1.3, 1.8, 1.7, 1.2, 
    1.7, 2.8, 1.2, 0.5, 0.5, 1.2, 0.8, 0.5, 0.4, 0.4, 1.2, 1.7, 2.9, 1.9, 
    0.5, 3, 0.2, 0.2, 0.1, 0.8, 1, 0.1, 2, 2.3, 0.2, 1.2, 1.3, 0.7, 1.4, 0.7, 
    1.4, 0.7, 1.4, 0.3, 0.3, 0.1, 0.8, 1.4, 1, 1.7, 5.4, 6.7, 6.2, 3.3, 1.2, 
    2, 3.5, 1.6, 1.3, 0.6, 0.2, 0.8, 0.6, 1.1, 0.3, 1, 0.9, 0.9, 0.9, 2.7, 
    2.2, 1, 2.7, 3.2, 1.5, 1.9, 4, 1.8, 3.8, 3.9, 3.5, 0.9, 2.7, 2.6, 3, 3.6, 
    3.6, 3.6, 2.6, 2.7, 2.2, 3.6, 2.8, 0.4, 2.6, 3.3, 0.7, 2.5, 0.6, 0.4, 
    1.1, 2.2, 2.3, 1.8, 0.9, 1.4, 3.8, 4, 4.1, 1.4, 2.8, 2.5, 3.8, 2.4, 3.2, 
    1.3, 1.1, 2.3, 3.5, 0.2, 0.8, 1.1, 0.5, 0.8, 0.5, 0.6, 0.3, 1, 1.1, 0.8, 
    1.3, 0.8, 1.7, 1.1, 1.4, 1.5, 0.7, 1.3, 2.5, 1.7, 0.1, 1.5, 1.2, 0.8, 1, 
    1.1, 1.2, 1.5, 0.9, 0.3, 1.9, 0.1, 0.9, 1.3, 0.8, 1.1, 1.8, 0.1, 1.5, 
    1.4, 1.2, 0.9, 0.8, 0.2, 1, 0, 0.2, 0.4, 0.7, 2.6, 0.6, 0.7, 0, 0.2, 0.7, 
    0.2, 0.2, 0.1, 0.8, 0.7, 1.1, 0.7, 1.3, 0.9, 1.4, 1.6, 3.4, 2.3, 3, 2.8, 
    3.4, 3, 3.5, 3.7, 5, 2.6, 5.6, 7.1, 3.8, 5.8, 4.9, 6.4, 5.7, 5.2, 5.7, 6, 
    5.1, 4.7, 4.5, 4.2, 3.7, 0.8, 0.9, 0.2, 1, 0.8, 1, 2.3, 1.1, 1.9, 1.6, 
    1.5, 1.9, 0.4, 0.8, 0.9, 1.8, 3.9, 2.9, 1.2, 1.1, 1.6, 1.8, 1.5, 1.4, 
    1.1, 0.5, 0.7, 0.5, 1, 0.5, 0.7, 0.8, 0.2, 0.5, 0.8, 0.3, 0.4, 0.6, 0.9, 
    1.1, 0.7, 0.8, 0.4, 0.6, 0.8, 0, 0.6, 0.7, 1.1, 0.1, 1.2, 1.2, 1, 0.7, 
    1.7, 0.5, 1.8, 2.1, 1.6, 0.6, 2.1, 1.4, 1.3, 2, 1.6, 1.8, 1.5, 1.8, 5.3, 
    8, 8, 6.4, 3.1, 4.4, 3.1, 1.4, 1.3, 1.3, 1.8, 1.7, 2.2, 1.7, 2.1, 4.6, 
    3.9, 3.7, 3.5, 3.3, 0.8, 1.5, 2.4, 1.6, 3.6, 2.7, 4.1, 6.3, 3.3, 4.5, 
    1.9, 2.1, 2.1, 3.5, 3.1, 2.9, 3.3, 2.8, 4.9, 4.7, 3.8, 4, 4.4, 5, 5.2, 
    5.3, 4.5, 3.8, 2.5, 1.5, 1.2, 2.8, 1.7, 1.7, 0.9, 0.9, 0.7, 0.6, 0.7, 
    1.2, 1.1, 1.2, 0.9, 1.3, 3.6, 5.6, 5.6, 5.6, 6.7, 6.2, 7.5, 9.1, 9, 8.9, 
    8.5, 8.3, 10.1, 12.1, 12, 11.9, 11.7, 11.5, 9.8, 9.4, 7, 2.2, 3.5, 1.2, 
    5.5, 5, 6.1, 3.6, 1.8, 1.5, 2, 0.8, 2.8, 5.6, 7.1, 4.5, 4.3, 5.6, 5.4, 
    2.2, 1.7, 3.5, 3.2, 4.3, 5.2, 5.2, 5, 5, 5.7, 4.5, 3.8, 3.7, 3.6, 3.6, 
    3.8, 2.8, 2.8, 1.5, 2.9, 3.6, 3.7, 4.1, 4.3, 3.6, 3.7, 4.1, 3.4, 2.7, 
    3.8, 3.2, 3.4, 0.8, 1.8, 0.7, 0.7, 0.3, 1.4, 1.2, 0.5, 1.1, 1.4, 3.3, 
    2.3, 0.8, 2.4, 0.7, 2.8, 3.7, 3, 2.9, 4.4, 4.2, 0.9, 3.5, 3.5, 3.6, 3.5, 
    1.5, 1.2, 0.8, 1.6, 0.7, 0.8, 0.9, 1.7, 0.7, 0.8, 0.8, 1.8, 2.1, 2.7, 
    2.8, 2.9, 3, 2, 1.7, 1.3, 1, 2.1, 1.3, 1.6, 2.6, 0.9, 1.6, 0.8, 2.4, 1.8, 
    0.9, 1.5, 1.4, 1.8, 1.7, 0.9, 1.4, 0.9, 1.5, 1.6, 2, 0.8, 1.7, 2.1, 1.1, 
    0.3, 0, 1, 0.3, 0.5, 1.3, 0.8, 1.4, 0.5, 0.1, 0.7, 1.3, 0.4, 0.6, 1.4, 
    1.5, 1.5, 1.6, 2, 3.9, 2, 4.9, 5.6, 1, 0.9, 5.4, 0.7, 2.6, 1.4, 1.2, 0.9, 
    4.3, 3.4, 4.5, 4.4, 4, 3.3, 3.9, 3.7, 4.2, 3.6, 3.1, 2.5, 4.1, 3.8, 2.6, 
    2.6, 1.3, 1.8, 1.4, 0.4, 0.9, 0.3, 0.2, 0.6, 0.7, 1, 1.2, 0.4, 1, 0.2, 
    0.9, 1.4, 1.2, 2.8, 2.5, 2.8, 0.6, 3.2, 2, 2.3, 2.4, 1.7, 5, 4.9, 4, 5.3, 
    2.9, 1.6, 2.6, 3.2, 2.5, 2.9, 2.6, 2.2, 1.4, 0.1, 0.1, 2.2, 1, 2.2, 0.7, 
    2.2, 2.4, 1.3, 0.8, 1, 0.5, 3.1, 1, 1.7, 1.4, 2.9, 3.1, 2.1, 0.6, 1.3, 
    0.6, 0, 1.5, 1.9, 2.1, 1.7, 1.5, 1.5, 1.4, 7.9, 10.4, 9.7, 10.4, 7.3, 
    4.9, 1.1, 0.9, 1.2, 0.1, 0.2, 0.8, 0.7, 0.2, 0.6, 8.4, 9.4, 10, 10.1, 
    10.3, 11.3, 10.7, 11.7, 11.6, 11.4, 11.1, 10.6, 11.6, 11.1, 10.6, 11.3, 
    10.8, 9.4, 7.6, 8.2, 8.1, 7.4, 7.7, 8.6, 8.2, 8.1, 7.2, 6, 4.1, 2.8, 2.7, 
    0.9, 1.9, 3.7, 4.4, 4.6, 3.9, 3.6, 3.6, 2.5, 2.2, 1.8, 1.1, 0.7, 0.2, 
    0.3, 1.9, 1.4, 1.2, 0.9, 1.4, 1.3, 1.7, 1.3, 1.1, 2.1, 2.5, 1.7, 1.6, 
    1.2, 2.4, 1.3, 1.9, 2.1, 1.1, 1.8, 1.5, 2.2, 1.7, 0.9, 0.5, 0.6, 0.7, 
    1.5, 0.7, 1.5, 1.5, 1.8, 0.6, 0.7, 0.9, 1.4, 0.2, 0.4, 2.5, 2.4, 3.3, 
    4.7, 4.8, 3.7, 2.9, 2.9, 3.3, 4, 3.2, 2.6, 5.2, 6.1, 6, 5.2, 5.9, 6, 7.1, 
    5.5, 5.6, 1.9, 2.7, 0.6, 1.3, 2, 0.4, 0.5, 1.1, 0.6, 0.6, 0.8, 1.2, 0.8, 
    1, 0.9, 1.9, 2.1, 1.1, 0.6, 0.8, 1, 0.2, 1.8, 2.1, 3.3, 0.4, 3, 0.5, 0.7, 
    0.5, 0.6, 0.7, 2.6, 2.1, 1.8, 0.3, 1.5, 1.3, 1.3, 1.4, 1, 1.1, 1.6, 1.8, 
    1.7, 0.8, 1.5, 1.4, 1.1, 1.4, 1.4, 3.6, 4.4, 7.5, 8.9, 10.8, 11.1, 11.2, 
    11.5, 10.6, 9.9, 10.2, 9.1, 10.1, 9.2, 10.1, 10.1, 10.2, 11, 9.5, 9.4, 
    7.9, 9.7, 10.6, 7.2, 5.3, 5.6, 5, 4.5, 3.3, 7.3, 8, 8.9, 6.5, 5.8, 5.5, 
    3.5, 1.3, 1.4, 1.5, 1.6, 0.6, 1.5, 0.4, 0.3, 1.8, 2, 2.1, 2.7, 1.8, 3.4, 
    2.1, 1.6, 0.8, 1, 1.1, 2, 2.5, 2.4, 2.5, 3, 2.5, 1.6, 4.2, 7, 8.4, 8.9, 
    8.7, 8.8, 8.9, 8.3, 7.4, 7.9, 8.3, 7.6, 7.5, 6.4, 6.2, 5.3, 5.8, 6.4, 
    5.1, 2.4, 2.1, 0.5, 3.3, 2.8, 2, 1.7, 2.7, 0.8, 1.6, 2.3, 2, 1.7, 0.9, 
    1.3, 1.7, 1.6, 0.6, 1.1, 0.9, 0.8, 0.8, 1.8, 2.9, 1.4, 0.8, 1.3, 1.8, 
    1.1, 2.4, 2.6, 1.9, 0.7, 1.1, 1.2, 1.2, 0.9, 0.3, 0.5, 0.7, 1.2, 0.9, 
    0.7, 0.8, 0.5, 0.2, 0.6, 0.8, 0.4, 0.8, 0.8, 0.9, 1.5, 1.2, 1.6, 0.7, 
    0.8, 0.8, 0.9, 1.2, 1.6, 0.5, 1.9, 1, 1, 0.4, 1.4, 1, 0.6, 0.9, 1.2, 1.2, 
    0.7, 0.7, 1.6, 0.8, 1.3, 0.6, 0.6, 1.4, 0.9, 0.4, 1.1, 0.6, 1, 1.1, 0.6, 
    1.6, 0.5, 0.8, 2.4, 2.9, 3, 2.5, 2.7, 0.8, 0.1, 1, 0.9, 1.7, 2.9, 3.6, 
    1.9, 2.1, 0.5, 0.4, 2.7, 4.3, 4.9, 3.6, 3.1, 3.8, 4.3, 3.5, 4.3, 4.8, 
    3.3, 2.7, 2.7, 1.8, 1.9, 7.2, 2.7, 4.1, 5.8, 8.8, 8.3, 3.3, 6.2, 6.4, 
    4.6, 0.4, 1.4, 2.2, 2.9, 4.1, 2.2, 3, 2.5, 3.5, 3.4, 3.2, 3.3, 0.4, 1, 
    0.7, 0.7, 1.2, 3.7, 4, 4.3, 0.7, 2.2, 2.3, 1.6, 0.9, 0.5, 1, 0.8, 1.5, 
    0.6, 1.5, 2, 1.1, 1.2, 2.2, 1.1, 0.5, 0.6, 0.5, 0.4, 1.1, 0.5, 0.2, 0.8, 
    0.7, 0.3, 0.8, 0.6, 1.6, 1.2, 0.8, 0.2, 0.9, 1, 0.6, 1.4, 0.5, 0.1, 1.3, 
    0.8, 0.7, 0.6, 0.9, 0.6, 0.8, 0.1, 1, 0.9, 1.4, 4.5, 3.7, 2.9, 5.6, 1.8, 
    4.8, 4.5, 2.9, 4.1, 2.9, 3.7, 1.9, 2.1, 0.8, 0.7, 1.3, 0.7, 0.9, 0.5, 
    0.4, 0.6, 0.4, 0.7, 2.2, 0.8, 1.6, 0.9, 1.2, 1, 0.9, 1.8, 2.3, 1.9, 4.8, 
    6.8, 3.9, 3, 2, 3.7, 6.8, 1.5, 1.8, 4.4, 6.8, 5.2, 7.3, 6.2, 4, 2.1, 1.4, 
    2.3, 0.6, 1, 1.1, 1.8, 2, 2.3, 2.6, 1, 0.3, 1, 6, 4, 6.4, 6.9, 4.2, 4.3, 
    4.2, 4.7, 1.3, 0.7, 0.8, 0.6, 1.4, 0.6, 0.4, 1.9, 2.2, 2.4, 0.8, 1.4, 
    0.6, 0.7, 2.1, 0.9, 0.6, 0.8, 0.7, 1.3, 2.9, 1.1, 0.7, 1.6, 2.3, 4.3, 
    2.6, 1.8, 1.2, 1.1, 1.7, 1, 1.5, 0.9, 1, 0.9, 1.7, 2.3, 1.1, 1.4, 0.4, 
    1.4, 0.6, 0.4, 1.4, 0.4, 0.9, 1, 0.2, 0.8, 0.7, 2.1, 0.8, 1.2, 0.7, 0.4, 
    0.8, 1, 1.7, 1.1, 0.8, 1.1, 0.3, 1.1, 1.6, 0.3, 0.5, 0.3, 0.3, 0.9, 0.5, 
    0.7, 0.6, 1.6, 1.1, 0.9, 0.7, 1.2, 0.4, 0.3, 0.3, 0.5, 0.5, 1.4, 0.7, 
    0.8, 1.1, 0.9, 0.3, 0.7, 1.2, 1.5, 0.6, 0.6, 4.9, 5.1, 7, 5.8, 7.2, 6.8, 
    5.2, 5.4, 1.7, 3.3, 3.5, 3.5, 4.5, 8.3, 6.9, 5.1, 3.9, 2.3, 2.2, 6.3, 
    8.5, 4.7, 5.6, 8.9, 7.9, 4.9, 4, 4.4, 4.6, 6.7, 9.6, 10.4, 9.4, 9.9, 8.7, 
    8.3, 7.6, 7.6, 8.8, 6.6, 7.3, 7.3, 8, 7.7, 6.6, 8.8, 8.8, 9, 7.4, 7.7, 
    7.4, 5.7, 6.8, 3.1, 1.3, 3, 3.1, 1.3, 1, 1, 0.4, 0.1, 0.6, 0, 0.1, 3, 
    1.6, 3.5, 2.7, 0.9, 0.6, 1.3, 0.6, 1.8, 2.3, 2.5, 0.2, 0.7, 1.9, 1.2, 
    1.4, 0.9, 0.7, 3.1, 4.3, 2.9, 3.3, 4.3, 3.1, 3.1, 5.5, 6.9, 2.6, 2.3, 
    2.2, 3, 5.4, 2.8, 3, 5.1, 2.7, 1.7, 1.2, 1.9, 0.8, 2.1, 0.3, 0.9, 1.3, 
    1.6, 0.8, 0.7, 1.5, 1.4, 1.5, 1.7, 1.7, 1.1, 0.5, 0.3, 3.5, 4, 3.9, 4.5, 
    7.6, 3, 1.2, 1.9, 1, 1.1, 2, 2.1, 1.1, 1.2, 3.7, 4.5, 4.9, 6, 4.7, 7.5, 
    6.5, 6.6, 8, 8, 8.1, 8, 7.4, 7.6, 8.1, 4.7, 2.9, 2.4, 2.5, 0.9, 1.2, 6.7, 
    5.8, 6.7, 5.7, 5.8, 4.2, 0.2, 1.9, 5.4, 6, 6, 5.9, 5.6, 5.5, 4.3, 5.4, 
    7.4, 6.9, 4.3, 5.1, 4.5, 3.7, 3.7, 2.9, 2.5, 1.6, 2, 1.2, 1.4, 2.2, 1.3, 
    0.2, 0.2, 0.9, 1.7, 0.5, 1.5, 0.8, 0.4, 0.5, 0.4, 0.4, 1, 0.9, 1.4, 1.3, 
    0.9, 0.9, 0.9, 0.7, 0.9, 1.7, 0.9, 0.1, 0.4, 0.4, 1.1, 0.5, 3.5, 1.1, 
    1.4, 1, 0.6, 0.3, 0.7, 0.6, 1.4, 0.8, 0.5, 0.6, 0.6, 0.8, 1, 0.8, 0.2, 
    2.7, 0.9, 0.7, 0.8, 0.4, 0.3, 1.6, 0.9, 0.7, 0.9, 1.5, 1.7, 1.6, 1.3, 
    0.2, 1.3, 1.8, 1.2, 1.2, 1.2, 1.1, 1.1, 1.5, 1.1, 0.4, 1, 2.6, 1.7, 2.1, 
    1.4, 1.4, 0.8, 1.2, 1.4, 1.3, 1.8, 1.8, 1.3, 3.1, 0.5, 2, 1.8, 1.7, 1.4, 
    1, 0.7, 5.3, 5.5, 5, 2.3, 4.2, 5, 7.3, 6.8, 6.2, 7.8, 9.4, 11.1, 6.6, 
    6.2, 8.4, 7.9, 8.3, 8.7, 8, 8.5, 9.6, 9.9, 9.7, 9.2, 7.3, 7.9, 8.3, 8, 
    7.6, 8, 7, 7.7, 7.9, 9.3, 8.9, 7.8, 8.5, 8.3, 8.5, 9.1, 8.2, 6.1, 5.7, 7, 
    7.7, 5.5, 5.3, 5.1, 5.6, 8.2, 7.5, 5.9, 4, 4.7, 3.2, 3.7, 4.5, 3.4, 4.6, 
    5.4, 3.1, 6.1, 3.8, 4.2, 7.3, 7.1, 6.5, 7.9, 10.6, 9.6, 8.4, 9, 10.6, 
    8.7, 9.9, 10.3, 9.3, 8.8, 8, 8.9, 7.5, 7.9, 8.7, 9.9, 9.4, 9.7, 10, 9.3, 
    9, 9.3, 9, 10, 9.3, 8.3, 7.5, 7.8, 8.7, 8.5, 7.8, 7.6, 8.1, 6.5, 5.7, 
    6.7, 6.5, 6.5, 7, 8.1, 6.9, 6.7, 6, 7.6, 5.1, 5.3, 7.1, 6.7, 5.6, 6.3, 3, 
    3.8, 3.1, 2, 1.4, 4.9, 5.4, 4.8, 4.3, 4, 4.7, 4.3, 4.7, 2.9, 4.3, 3.6, 
    3.2, 3.2, 3.8, 1.1, 0.8, 1, 1, 4.5, 4.3, 5, 5.5, 5.3, 7, 4.7, 5.4, 6.1, 
    5, 6.3, 5.2, 5.2, 5.5, 6.9, 6.5, 7.2, 5.8, 4.8, 4.9, 3.4, 3.2, 3.5, 2.9, 
    1.4, 1.5, 0.6, 1.3, 1.3, 0.5, 0.7, 1.1, 0.2, 1.5, 0.8, 1.5, 2.1, 1.4, 
    0.3, 1.5, 0.5, 0.8, 0.2, 0.4, 0.2, 0, 1, 0.7, 0.7, 0.3, 0.4, 0.4, 0.4, 
    1.1, 1.5, 0.8, 1.7, 0.3, 1, 0.4, 0.1, 0.5, 0.2, 0.6, 1, 1, 1, 0.4, 0.1, 
    0.2, 0.4, 0.9, 0.3, 0.6, 2.7, 2.8, 2.2, 0.8, 2.8, 0.2, 0.5, 1.2, 0.1, 
    0.2, 0.6, 2.2, 0, 0.8, 0.1, 0.7, 1.8, 2, 1.2, 0.8, 2, 1.1, 0.2, 1.2, 1.1, 
    0.8, 1.9, 0.1, 0.9, 0.3, 0.4, 0.5, 3.2, 1.3, 1.8, 0.9, 3.2, 4.4, 4.1, 
    4.5, 3, 2, 1.3, 3, 3.7, 3.4, 0.5, 1.6, 2, 0, 0.9, 1, 2, 2.2, 1.6, 0.4, 
    0.2, 0.6, 1.3, 0.8, 0.6, 0.3, 0.5, 1.1, 0.9, 0.6, 0.6, 1.6, 1.9, 1, 1.2, 
    1.8, 0.8, 0.6, 0.1, 0.9, 0.1, 1.7, 1, 1.2, 1, 0.3, 1, 1.5, 0.4, 0.9, 0.6, 
    3, 4.9, 4.9, 5.2, 5.2, 5.2, 4.6, 4.7, 5.1, 5.3, 5.7, 5.5, 5.6, 7.1, 7.8, 
    6.6, 6.8, 6.7, 6.9, 7.1, 5.9, 7.4, 8.5, 7.8, 5.7, 3.1, 0.8, 1, 5, 1.7, 
    2.9, 0.6, 1.6, 0.8, 0.8, 1.5, 2, 1.3, 3.3, 0.8, 2, 5.1, 4, 2.8, 1.1, 1.8, 
    1.5, 1.3, 1.9, 1.6, 1.6, 2.1, 2.6, 1.6, 1.8, 1.5, 2.4, 1.8, 0.9, 0.3, 1, 
    2.4, 0.8, 0.5, 0.4, 0.5, 0.1, 0.3, 0.2, 0.1, 0.3, 1.5, 0, 0.3, 0.4, 0.4, 
    0.7, 0.1, 0.1, 0.8, 0.2, 0.3, 0.7, 1.4, 0.5, 1.3, 0.1, 0.2, 0.6, 1.7, 
    0.6, 0.5, 0.1, 0.4, 0.1, 0.5, 0.6, 0.6, 0.1, 0.1, 0, 0.2, 0.2, 0.1, 0.6, 
    0.3, 0.8, 0.1, 0.2, 0.7, 0.8, 0.1, 0.4, 0.6, 0.7, 0.3, 0.8, 0.9, 0.1, 
    1.6, 0.3, 1.5, 0.7, 0.7, 1.8, 0.2, 0.6, 1.3, 0.8, 1, 0.6, 1.2, 0, 0.3, 
    0.8, 0.7, 0.5, 0.3, 1.1, 0.1, 1, 1.4, 3.1, 5.1, 5.4, 5.5, 5.1, 2.2, 3.6, 
    3.5, 2.5, 3.1, 2.4, 3.4, 0.3, 1.1, 0.6, 0.9, 0.1, 1.6, 2, 2, 0.9, 0.3, 
    0.1, 0.1, 0, 0.5, 0.9, 1.6, 0.9, 1, 1, 0.3, 0.5, 1, 0.8, 0.9, 0.9, 0.8, 
    0.4, 0.3, 0.3, 0.4, 0.5, 0.5, 0.5, 0.2, 0, 2.1, 3.2, 3.4, 4, 1.8, 0.6, 
    0.8, 0.4, 0.1, 0.5, 0.7, 0.6, 0.3, 0.3, 0.3, 0.1, 0.3, 0.8, 1.1, 0.7, 
    0.9, 0.1, 0.1, 0.3, 0.8, 0.4, 0.6, 0.7, 0.2, 0.2, 0.7, 1.3, 0.3, 1.1, 
    0.6, 0.2, 0.4, 0.1, 0.2, 0.1, 0.2, 0.3, 0.2, 0.6, 1.1, 2.4, 0.5, 1.7, 
    3.6, 4.5, 4.7, 1, 0.7, 1.6, 1.5, 0.7, 0.7, 0.3, 0.4, 0.5, 2.1, 0.7, 0.3, 
    0.6, 0.3, 1.3, 0.6, 0.8, 0.7, 0.4, 0.6, 1.4, 1.7, 1, 0.6, 0.1, 0.2, 0.6, 
    0.5, 0, 0.5, 0.6, 0.7, 0.7, 0.2, 0.6, 0.4, 1, 0.4, 0.6, 1.2, 0.2, 0, 0.2, 
    0.2, 0.3, 0.3, 0.9, 0.4, 0.4, 0.5, 0.2, 0.7, 4.1, 3, 2.3, 3.1, 3.7, 4, 
    4.6, 4.5, 5.3, 3.6, 4.5, 3.7, 4.8, 3.7, 4.8, 3.8, 2.8, 1.4, 2.6, 2.2, 
    4.3, 4.5, 6, 8.7, 6.5, 9, 6.8, 4, 4.1, 4.1, 6.1, 3.7, 3.3, 3.8, 4.6, 1.5, 
    3.3, 3.4, 3.4, 2.9, 1.9, 3.5, 4, 3.2, 4, 5.9, 7.6, 4.9, 6.3, 7.1, 5.5, 
    9.1, 8.7, 6.6, 10.5, 8.8, 7.3, 8.3, 7.4, 4.1, 7.5, 5.7, 4.5, 3.2, 2.8, 
    0.6, 0.8, 0.8, 0.5, 0.3, 0.6, 0.7, 0.7, 1.3, 0.5, 0.4, 0.1, 0.3, 1.1, 
    1.1, 1.2, 0.7, 0.3, 0.6, 1.4, 1.2, 1, 1.5, 0.5, 1.3, 0.4, 0.3, 0.4, 3.1, 
    1.3, 0.6, 0.2, 0.8, 0, 0.3, 0.3, 0, 0.2, 0.3, 0.3, 0.4, 0.1, 0.9, 0.2, 0, 
    0, 0, 0, 0, 4.5, 0.7, 4.5, 4.2, 4.6, 4.6, 5.6, 4.5, 3.4, 4.9, 3.6, 4.7, 
    3.8, 3.6, 1.2, 0.2, 1, 1.3, 1.2, 1.5, 1.6, 0.9, 1.8, 0.6, 1.2, 1, 1.3, 
    1.9, 1.5, 1, 0.2, 0.3, 1.9, 0.1, 0.5, 1.5, 0.8, 0.6, 0.1, 0.5, 0.2, 0.4, 
    1, 0.3, 0.3, 0, 0, 0, 0, 0, 4.1, 5.5, 4.8, 5.2, 5.2, 4, 2.3, 1.1, 1.4, 
    2.7, 2.2, 1.5, 2.2, 3.5, 0.9, 2.5, 1.3, 2.5, 2, 0.9, 2.1, 1.9, 1.4, 1, 
    0.4, 0.1, 0.5, 1.1, 0.4, 1.2, 0.8, 0.5, 0.1, 0.5, 0.1, 0.3, 0.8, 1, 1.1, 
    0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.7, 0, 0, 0.6, 5.4, 6.7, 6.9, 5.8, 5.2, 4.6, 1.8, 6.7, 7.3, 
    6.1, 3.5, 2.2, 1.6, 1.6, 1, 0.9, 1.9, 1.7, 0.8, 1.5, 0.9, 0.3, 1.8, 0.8, 
    2.5, 1.5, 1.3, 3, 1.2, 1.1, 0.4, 1, 0.3, 0.5, 1, 0.5, 0.4, 0.8, 0.4, 0.4, 
    0.3, 0.6, 0.3, 1.2, 0.9, 0.5, 1, 0.4, 1.4, 1.6, 1.1, 0.8, 0.9, 1.2, 2, 
    0.4, 0.8, 0.6, 1.3, 0.4, 0.9, 0.1, 1.2, 1, 0.8, 0.7, 1.6, 0.2, 1, 1, 0.2, 
    1.3, 1.9, 1.4, 0.2, 1.1, 0.6, 1, 1, 1, 1, 1.3, 0.7, 1, 1.2, 0.2, 0.4, 
    0.9, 1.2, 0.9, 0.1, 0.5, 1.1, 0.8, 0.5, 0.3, 0.4, 0.9, 0.7, 0.6, 1.5, 
    1.8, 0.6, 0.7, 1.2, 0.3, 0.7, 0.3, 0.8, 1.1, 1.6, 3.2, 3.5, 3.5, 3.4, 
    0.4, 0.4, 2, 0.6, 0.1, 1.1, 0.5, 0.1, 1.1, 1.1, 0.6, 0.8, 0.3, 2, 0.7, 
    0.8, 1, 0.6, 1.3, 0.8, 4.4, 6.3, 5.7, 5, 4.2, 0.9, 0.6, 2.2, 0.3, 0.1, 
    0.7, 0.3, 0.2, 0.7, 0.1, 0, 0, 1.6, 1.6, 0.5, 0.1, 0.6, 0.4, 1.2, 1.5, 
    0.2, 0.3, 0.9, 0.2, 0.6, 0.3, 1.7, 0.9, 0.7, 0.5, 0.3, 1.2, 1.2, 1.2, 
    2.9, 1.6, 4.7, 5.3, 4.3, 6, 5.6, 6.3, 4.3, 4.5, 2.4, 0.9, 5.8, 6.4, 6.3, 
    7.1, 7.1, 8.6, 8.4, 7.7, 7.1, 9.8, 9.3, 10.6, 10.6, 10.2, 9.6, 9.1, 8.3, 
    7.7, 6.2, 6.6, 6.4, 6.6, 4, 2, 0.5, 2.5, 0.1, 0.3, 0.3, 0.1, 1, 0.4, 0.3, 
    0.5, 0.9, 0.2, 0.4, 0.7, 0.8, 0.8, 0.7, 0.2, 0.1, 0.5, 0.7, 0.6, 0.4, 
    1.1, 0.5, 0.5, 1.5, 0.8, 1.5, 0.4, 0.3, 1, 1.7, 0.8, 1, 1.4, 0.7, 1.6, 
    1.9, 1.2, 0.3, 0.6, 0.4, 0.4, 0.4, 1.1, 0.7, 0.4, 1.5, 0.9, 0.9, 0.2, 
    0.2, 0.2, 0.9, 1.4, 0.4, 1.4, 5.7, 6.6, 5.8, 4.4, 5, 5, 5.7, 5.6, 6.1, 
    4.6, 5.6, 4.5, 3.8, 3.6, 4.6, 4.6, 5.5, 4.3, 2.1, 3.7, 2.1, 1.5, 4.8, 
    5.3, 6.8, 5, 4.9, 4.3, 4.7, 4.4, 4.3, 4.3, 5.5, 6, 8.1, 8.3, 9, 8, 4.6, 
    3.4, 1.5, 1.3, 4.7, 4.8, 6.2, 5.8, 6.1, 5.3, 5.4, 5.5, 5.9, 3.8, 1.6, 
    0.7, 3.5, 5, 5.5, 3.5, 3, 5, 4.1, 2.2, 4.7, 3.6, 3.9, 5.7, 6.2, 6.3, 6.3, 
    4.7, 3.6, 3.6, 2.9, 2.9, 2.5, 4.3, 2.7, 3, 1.4, 0.7, 0.7, 1.2, 0.1, 1.4, 
    3.9, 5.7, 6.3, 4.9, 2.7, 3.7, 4.9, 4.9, 4.5, 6.3, 5.6, 5.8, 5.3, 5.5, 
    4.6, 5.6, 5.5, 3.2, 4, 1.1, 3.8, 1.3, 4.2, 3.9, 2.8, 0.8, 1, 1.3, 1.1, 
    1.3, 0.6, 1.7, 0.1, 1.6, 1.5, 1.6, 0.5, 0.2, 0.6, 1, 0.1, 0.2, 0.1, 1.7, 
    1.1, 0.5, 1.1, 0.9, 1.5, 2.5, 1.1, 1.8, 1.3, 2.2, 1.2, 1.3, 2.4, 2.1, 2, 
    1.6, 1.9, 4.7, 1.6, 1.7, 2.7, 0.9, 0.9, 0.8, 1.8, 1.2, 1.5, 1.7, 1.1, 3, 
    1.5, 5.7, 2.2, 2.8, 5, 3.6, 4.1, 3.2, 1.3, 2.1, 3, 5.3, 3.9, 4.4, 5.3, 
    7.2, 5.6, 6.8, 8.2, 8.3, 7.7, 10.3, 8.5, 7, 7.6, 10.2, 8.1, 8.1, 9.6, 
    10.1, 10.5, 10.5, 10.3, 10, 8, 7.1, 7.3, 6.4, 5.9, 3.6, 6.7, 8.1, 10.2, 
    10.3, 9.9, 9, 9.5, 8.7, 7.9, 8.5, 8, 6.6, 5.2, 5.9, 4.6, 5, 5.5, 5.6, 
    6.6, 5.3, 4.5, 2.8, 1.3, 4.4, 5.4, 5.1, 5.5, 3.3, 3.2, 3, 3, 1.7, 1.5, 
    1.7, 1.6, 3.7, 5, 4.5, 3.7, 4.1, 3.5, 1.7, 3.9, 0.6, 1.9, 0.3, 0.7, 0.4, 
    0.3, 1, 1.1, 0.6, 0.6, 0.5, 0.7, 0.9, 0.6, 1.2, 0.8, 1.3, 0.8, 0.2, 0.4, 
    0.8, 2.5, 4, 5, 5, 3.7, 2.4, 0.3, 0.4, 0.8, 1.7, 1.9, 4.4, 4.7, 5.2, 8.2, 
    7.3, 4.1, 5, 5.7, 6.2, 6.1, 7.7, 5.7, 7.7, 7, 8.1, 7.5, 8.8, 6.8, 6.1, 
    6.2, 6.8, 5.9, 5.9, 6.4, 5.4, 4.9, 6.1, 4.5, 4, 3.1, 3.5, 3, 1.1, 2.6, 
    1.9, 0.4, 0.8, 2.1, 0.4, 0.8, 0.6, 2.4, 1.4, 1.1, 0.9, 0.2, 0.8, 1, 0.7, 
    0.7, 1, 1, 0.7, 1, 1.7, 1.8, 1.7, 1.2, 0.3, 1, 1.2, 1.4, 1.4, 1.5, 1.1, 
    1.1, 0.7, 0.8, 0.6, 4, 3.5, 4, 3.8, 4, 3.5, 6, 6, 4.5, 4.6, 3.3, 4.5, 
    3.6, 3.5, 3.5, 3.1, 2.8, 4.1, 3.6, 2.8, 2.1, 3.5, 1, 3.2, 4.2, 3.1, 3.5, 
    5, 3.8, 5, 4.5, 3.7, 4.3, 4.1, 3, 3.9, 2.8, 3.5, 2.9, 1.9, 0.3, 0.4, 0.8, 
    0.3, 0.3, 0.9, 0.6, 0.7, 1.1, 0.2, 0.9, 0.3, 0.8, 1, 1, 0.9, 1, 0.2, 1.4, 
    0.8, 0.6, 0.7, 1.1, 0.1, 0.9, 1.1, 1.1, 0.6, 0.7, 0.9, 1.2, 1.3, 0.7, 
    1.3, 1.4, 1.3, 0.9, 1.7, 5.3, 3.6, 4.5, 4.4, 0.8, 5.1, 5, 4.7, 4.8, 3.2, 
    2.6, 4.5, 4, 5, 4, 3.4, 5.6, 5.2, 5, 5.8, 6.8, 7.4, 7.4, 8, 8.6, 10.2, 
    3.2, 7.4, 8.9, 9.5, 6.7, 7.5, 8.8, 5.5, 3.5, 2.5, 3.5, 4.2, 4.2, 6.2, 
    6.3, 5.2, 5.9, 6.3, 4.8, 4.5, 5.4, 2.8, 3.6, 2.5, 3, 1.3, 0.1, 0.6, 0.3, 
    0.3, 1, 0.4, 0, 1, 0.5, 0.1, 0.7, 0.8, 0.3, 0.2, 1.2, 1.5, 0.3, 3.1, 6, 
    5.8, 5.1, 4.3, 4.6, 4.1, 4, 3.6, 1.5, 1.7, 2, 0.4, 0.6, 0.8, 1, 0.2, 2.3, 
    0.4, 3.2, 4.4, 5.5, 2.7, 3.8, 4, 4.6, 3.4, 1.9, 0.1, 0.2, 0.2, 0.1, 0.9, 
    1.4, 0.4, 0, 1, 1, 0.1, 1.3, 0.9, 2.7, 1.9, 2.5, 1.4, 1.7, 3.9, 3.6, 3.7, 
    4, 2.7, 1.7, 1.5, 2.4, 1.1, 1.4, 2.1, 3, 2.9, 1.2, 2.1, 1, 1.5, 1.3, 3.5, 
    3.6, 1, 1.2, 1.2, 1.5, 1.5, 0.4, 0.2, 0.4, 0.5, 0.8, 0.3, 0.8, 0.8, 0.8, 
    0.7, 1.7, 0.8, 2.7, 0.9, 1, 0.6, 0.1, 0.7, 0.4, 0, 0.5, 0.4, 0.3, 0.4, 0, 
    0.2, 1.5, 1.6, 1.1, 1.2, 2.2, 0.5, 1.3, 0.5, 0.3, 0.7, 1, 1.1, 2.1, 1.1, 
    2.5, 1, 3.7, 2.8, 1.7, 2.7, 3, 7.7, 3, 3.6, 2.5, 4.3, 4.9, 3.2, 3.3, 3.4, 
    5.6, 6.8, 7.2, 8.6, 8.7, 8.2, 6.4, 3.6, 0.9, 0.6, 0.7, 1.2, 1.8, 0.9, 
    0.7, 0.5, 0.5, 0.6, 0.7, 0.4, 0.6, 0.5, 1.4, 0.4, 0.9, 0.4, 0.2, 0.6, 1, 
    2, 1.4, 2.2, 3, 4, 0.4, 1.5, 0.9, 0.2, 4.4, 4.5, 2.6, 0.9, 0.9, 0.2, 0.2, 
    0.2, 1.9, 0.9, 0.8, 1.3, 2.3, 0.6, 0.2, 1.4, 1, 0.2, 0.7, 1.1, 2.2, 5.5, 
    1.8, 7.6, 7.6, 9, 8.6, 8.9, 8.2, 8.1, 8.2, 7.9, 8.7, 7.1, 5.9, 8.4, 8.2, 
    9.3, 8.2, 8.6, 7.5, 4.2, 1, 1.2, 0.9, 1, 1, 2.4, 5.1, 7.3, 8.7, 9.4, 8.1, 
    6.7, 7.1, 7.6, 7.6, 7.2, 5.1, 7.1, 6, 4.7, 4, 6.6, 6.9, 6.9, 2.8, 7.7, 
    7.6, 7.4, 4.3, 2.3, 3.1, 3.6, 2, 0.5, 0.8, 1.4, 1.2, 1.3, 1.6, 0.3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.1, 5, 5.1, 5.2, 6.1, 4.2, 3.4, 4.3, 
    5, 4.9, 4.4, 6.2, 5.6, 5.3, 4.3, 4.2, 4.2, 4.2, 4, 0.8, 2.2, 2.1, 2.3, 
    3.9, 3.1, 2.7, 1, 1.8, 1.1, 1.7, 0.1, 0.2, 0.1, 0.4, 0.1, 1.3, 0.4, 0.3, 
    0.4, 0.2, 0.3, 0.3, 0.6, 1.1, 0, 0.1, 1.7, 0.9, 0.5, 0.2, 1, 0, 0.1, 1, 
    0.4, 0.6, 0.8, 0.3, 0.2, 0.9, 0.1, 3.8, 3.8, 3.8, 3.7, 2.9, 0.7, 0.9, 
    1.2, 3.2, 4.6, 4.6, 5.1, 6.2, 5.1, 2.2, 1.2, 1.2, 1.1, 0.8, 1.3, 1.2, 
    0.8, 1.1, 0.6, 0.7, 1.1, 1.5, 0.5, 0, 0.5, 1.1, 1, 1.4, 1.5, 0.6, 0.1, 
    0.9, 0.7, 0.8, 0.6, 0.5, 0.6, 1.1, 1.2, 0.4, 0.7, 0.6, 0.5, 0.7, 0.8, 
    0.9, 0.9, 0.5, 0.6, 0.2, 0.3, 0.2, 0.6, 0.4, 0.3, 0.3, 0.4, 0.1, 0.8, 
    0.1, 1.7, 0.4, 0.8, 0.9, 0.1, 0.2, 0.5, 0.5, 0.6, 0.4, 1, 1, 0.9, 0.4, 
    0.7, 0.7, 1.4, 0.9, 2.2, 1.2, 1, 1.2, 1, 0.6, 1, 1.3, 0.3, 0.8, 0.4, 0.1, 
    1, 0.4, 0.4, 1.3, 0.5, 0.8, 0.6, 0.5, 0.1, 0.3, 0.2, 0.2, 0.6, 0.9, 0.4, 
    0.1, 0.4, 0.9, 0.2, 1, 1.2, 1.1, 1.3, 1.6, 0.5, 1.9, 4.8, 1.3, 1.6, 1.5, 
    2, 1.1, 1.2, 1.2, 0.9, 1.6, 2.4, 2.4, 2.3, 3.4, 3.3, 2.6, 2.5, 3, 4, 1.9, 
    3.6, 3.2, 3.3, 2, 2, 3, 1.6, 1.2, 2.2, 2.2, 0.8, 3.7, 4.1, 3, 2.7, 2.1, 
    0.6, 1.5, 2.1, 5.3, 5.2, 2.7, 3.1, 2.2, 1.9, 0.7, 1.1, 2.6, 1.8, 1.4, 
    1.1, 3.6, 3.2, 2.5, 0.5, 0.8, 1, 1.5, 2.4, 2.5, 2.2, 2.6, 1, 0.9, 0.4, 
    0.2, 0.8, 0.6, 1.3, 0.4, 0.1, 0.2, 0.1, 0.5, 0.4, 0.8, 0.5, 0.9, 1, 0.5, 
    0.8, 0.6, 1.5, 0.8, 0.8, 0.4, 0.8, 0.6, 0.4, 0.4, 1.3, 0, 0.6, 0.9, 0.4, 
    1.5, 0.6, 0.5, 0.4, 0.6, 0.1, 0.1, 0.1, 0.4, 0.6, 1.6, 1.1, 0.3, 1.1, 
    0.5, 0.6, 0.4, 0.3, 0.1, 0.5, 0.2, 0.8, 0.5, 0.4, 1.1, 1.5, 1.7, 0.5, 
    0.1, 1.3, 0.2, 1, 0.8, 0.4, 0.2, 0.3, 1, 1.1, 0.5, 0.7, 0.5, 1.2, 0.9, 
    0.3, 2.6, 1, 0.1, 0.5, 0.8, 0.8, 0.8, 0.8, 0.8, 0.4, 0.5, 0.1, 0.9, 0.1, 
    1, 1.4, 1.4, 3, 3.4, 2.8, 4.5, 1.5, 0.5, 0.2, 0.3, 0.4, 0.5, 1.5, 0.6, 
    0.3, 1.1, 0.3, 0.8, 0.5, 2.5, 1.6, 0.2, 0.6, 0.6, 0.3, 0.2, 0.2, 0.2, 
    0.1, 0.2, 0.5, 0, 0.3, 0.5, 0.2, 0.7, 0.1, 1.1, 1, 0.2, 0.6, 0.5, 0.8, 
    3.9, 0.6, 1.2, 2, 5.6, 3.6, 2.1, 0.3, 1.6, 0.9, 0.5, 0.8, 2.6, 4.6, 6.6, 
    4.5, 5.1, 2.8, 1.6, 2, 1.3, 1.7, 1.4, 1.1, 1, 1.1, 1.4, 0.9, 0.3, 0.4, 
    0.3, 0.6, 0.6, 0.6, 0.5, 0.7, 0.5, 0.8, 0.8, 1, 0.5, 1.3, 0.1, 0.6, 0.8, 
    0.6, 1.3, 0.4, 1.9, 1, 1.4, 1, 1.2, 0.3, 0.1, 0.8, 1.5, 1.2, 0.3, 0.9, 
    1.4, 0.2, 2.4, 0.2, 0.3, 0.1, 1, 1.4, 1.2, 0, 0.3, 0.8, 0.9, 0.4, 4.1, 
    3.8, 3.1, 3.3, 4.4, 5.6, 4.6, 4.5, 4.9, 4.6, 7.5, 5.1, 4.6, 4.6, 5.7, 
    7.2, 4.4, 2, 6.3, 2.5, 2.5, 0.6, 2.8, 2.7, 4.1, 1.3, 1.9, 2.7, 4.8, 1.8, 
    1.5, 1.1, 1.7, 1, 0.3, 3, 5, 2.7, 0.8, 0.3, 0.7, 1.3, 0.5, 1.7, 1.2, 1.8, 
    0.9, 1.8, 0.7, 1.1, 2.1, 1.9, 0.6, 0.5, 1.6, 0.4, 2.3, 1.4, 1.4, 2, 0.8, 
    2.2, 4.1, 2.7, 0.6, 2, 3.2, 2.6, 1.1, 3.6, 2.8, 3, 1.2, 2.2, 1.3, 1.2, 3, 
    2.2, 3.1, 2, 1.5, 2.8, 1.9, 0.4, 0.3, 3.8, 5.8, 4, 3.2, 1.7, 1.4, 0.7, 1, 
    0.7, 0.6, 1, 1.1, 0.9, 2.2, 0.7, 0.5, 1.4, 1.4, 2.3, 1.5, 2.1, 0.8, 0.4, 
    1.7, 1.7, 1.4, 1, 2.7, 3.1, 3.9, 3, 2.9, 2.3, 2.1, 1.8, 1.9, 1.5, 1.3, 
    2.2, 3, 1, 0.9, 1.9, 1, 0.5, 0.6, 1.9, 0.6, 1.5, 1.4, 0.8, 0.9, 0.6, 2.7, 
    1.1, 2.7, 1.7, 1.4, 0.6, 0.6, 0.9, 0.7, 0.7, 0.1, 0.6, 0.5, 0.2, 0.9, 
    1.2, 0, 0.7, 0.1, 0.9, 0.2, 0.3, 1.3, 0.8, 0.3, 0.4, 0.6, 0.5, 0.2, 0.4, 
    0, 1.9, 0.6, 0.9, 1.8, 0, 1, 1.3, 0, 0.6, 1.9, 0.5, 2.2, 4.1, 5.1, 1.8, 
    0.9, 1.2, 0.3, 1.2, 1.1, 0.7, 0.8, 0.2, 1.3, 1.7, 0.4, 0.2, 0, 0.2, 1, 
    2.1, 1.9, 1, 0.3, 0.5, 0.2, 1.1, 0.6, 0.6, 0.6, 0.5, 0.5, 0.8, 0.5, 3.3, 
    5.7, 3.7, 2, 3.5, 2, 2.6, 1.8, 1.6, 0.5, 4.5, 3.4, 2.2, 0.9, 2.3, 0.9, 
    1.4, 0.7, 1.3, 2.3, 0.7, 1.7, 0.8, 0.7, 0.2, 0.6, 1.6, 1.5, 0.5, 0.7, 
    0.7, 1, 0.3, 0.5, 0.5, 0.6, 1.8, 0.7, 0.1, 0.3, 0.5, 0.7, 0.4, 0.6, 0.2, 
    0.2, 0.1, 0.2, 0.7, 0.3, 0.5, 1.1, 0.4, 0.8, 1, 0, 0.5, 0.7, 0.2, 0, 0.4, 
    0, 0.2, 1.1, 2.5, 0.3, 0, 0.8, 0.7, 0.2, 0.1, 0.6, 0.8, 0.5, 0, 0.7, 1.8, 
    0.5, 1.1, 0.2, 0, 0.4, 1, 0.1, 0.3, 0.1, 0.6, 1.1, 0.8, 0.3, 0.9, 0.6, 
    0.8, 0.5, 1.2, 0.6, 0.5, 0.7, 0.4, 0.5, 4.9, 4.9, 4.9, 3.4, 3.5, 4, 5.6, 
    4.9, 3.4, 3, 2.8, 2.4, 3.2, 3.9, 6.3, 3.2, 1.9, 1.3, 1.5, 0.3, 0.5, 0.1, 
    0.5, 1.3, 1.4, 2.3, 3.3, 2.6, 0.3, 0.2, 0.1, 1.4, 4.9, 6.1, 3.2, 7.6, 
    7.5, 6.1, 6.1, 7.2, 5.8, 4.1, 2.1, 1.1, 3.1, 0.7, 1.8, 1.9, 0.9, 1.6, 
    1.6, 1, 2, 4.8, 2.9, 2, 1.8, 5, 4.9, 1.4, 2.9, 0.5, 0.9, 0.7, 0.6, 0.6, 
    1.1, 1.1, 0.6, 1.5, 0.3, 0.3, 0.8, 0.5, 1.1, 0.2, 1.2, 0.3, 1.1, 0.8, 0, 
    0.5, 0.1, 1, 0.5, 0.7, 0.7, 0, 0.6, 0.3, 0.3, 0.7, 0.8, 0.1, 0.2, 1, 0.4, 
    0.6, 0.4, 0.5, 0.7, 0.3, 0.9, 0, 0.2, 0, 0, 0.6, 0.1, 0.8, 0.3, 1.2, 1.1, 
    0.2, 2, 1.2, 0.7, 1, 0.5, 0.9, 0.7, 1, 0.8, 1.3, 1.3, 1, 0.3, 2.2, 3.2, 
    2.2, 1.9, 2.1, 0.3, 0.5, 0.3, 0.4, 0.3, 0.1, 0.4, 1.3, 1.5, 1.2, 1, 0.1, 
    1.1, 0.7, 1, 3.5, 3.6, 7.4, 9.1, 7.5, 6, 6.5, 6.3, 3.8, 1.6, 0.8, 0.8, 
    1.9, 6.5, 9.9, 7.9, 6.4, 9.6, 11, 10.5, 10.6, 7.6, 5.5, 3.6, 5.8, 4.2, 
    4.4, 5.1, 3.5, 4.7, 7.2, 2.5, 6.5, 9.3, 5.1, 5.7, 6.4, 6.9, 4.1, 3.4, 
    1.8, 0.3, 0.2, 0.7, 1.3, 1, 0, 2, 0.6, 1.8, 2, 2, 1.9, 2.1, 1.5, 1.7, 
    0.1, 1.9, 2, 0.5, 0.2, 1, 0.1, 1.2, 0.5, 1, 0, 1, 0.4, 0.6, 0.3, 1.7, 
    1.8, 1.9, 0.8, 1.5, 1.8, 1.3, 2.2, 0.2, 1.5, 1, 2.5, 1, 0.3, 0.2, 1.1, 
    0.5, 0.2, 0.9, 0.6, 0.5, 0.7, 1.1, 1.1, 0.3, 0.2, 0.2, 0.7, 0.4, 1.1, 
    0.9, 0.4, 0.4, 2, 1.8, 0.7, 0.3, 0.8, 1.4, 1.3, 1, 0.9, 0.9, 0.5, 0.4, 1, 
    0.7, 0.7, 0.6, 0.8, 0.6, 1.1, 0.9, 0.3, 0.8, 0.9, 0.7, 0.6, 1.4, 0.8, 
    1.1, 1, 3.5, 2.5, 3, 2.6, 3.4, 3.4, 3.9, 6.3, 3, 0.8, 5.6, 4.3, 1.7, 3.4, 
    1.4, 1.4, 1.2, 3.2, 1.2, 3.3, 1.7, 1.7, 0.3, 0.5, 0.2, 0.7, 1.2, 0.4, 
    0.9, 1, 0.4, 0.4, 1.2, 0.8, 0.7, 1.1, 0.2, 0.4, 2.1, 1.4, 2.3, 0.3, 0.4, 
    1.9, 3.7, 1.3, 0.5, 1.1, 0.5, 1.4, 0.7, 0.5, 0.5, 0.7, 0.6, 0.7, 0.3, 
    1.4, 1.7, 2, 1, 3, 1.1, 1.3, 1.8, 1.8, 2.4, 0.9, 0.8, 0.4, 0.4, 0.9, 0.9, 
    0.6, 0.9, 0.4, 0.2, 0.2, 0.3, 0.3, 0.4, 1.4, 0, 0, 0, 0.6, 1, 0.6, 0.9, 
    0.4, 0.2, 0.6, 0.5, 1, 0.9, 1, 1.9, 1.3, 1.1, 1.6, 0.8, 1.6, 0.8, 0.9, 
    0.7, 0.4, 0.3, 1.1, 1.6, 1.6, 0.5, 0.3, 0.3, 0.3, 1, 1.2, 0.2, 0.2, 0.8, 
    0.4, 0.4, 0.3, 0.3, 0.7, 0.6, 1, 1.8, 1.3, 1.2, 0.4, 5.9, 4.6, 4.3, 4.7, 
    2.4, 2.8, 3, 1.4, 1.3, 1.1, 1, 1.6, 0.8, 1.9, 0.8, 1, 0.6, 0.5, 0.1, 0.6, 
    1.2, 1.2, 4.9, 4.7, 4.6, 4.3, 5.4, 4.5, 4.7, 1.2, 5, 1.3, 1.1, 1.8, 2.1, 
    0.6, 0.5, 1.8, 0.4, 0.9, 1.4, 0.9, 0.6, 1, 1.2, 0.7, 0.8, 2, 2.1, 4, 3.7, 
    5.5, 0.8, 0.3, 0.8, 0.5, 0.7, 0.9, 1.5, 1.3, 0.7, 1.5, 0.7, 0.6, 1.6, 
    0.9, 0.9, 1, 0.8, 0.3, 1.2, 1.1, 0.8, 3, 1.4, 4.6, 3, 3.1, 1.1, 3, 1.3, 
    1.1, 1, 1.9, 0.9, 2.6, 1.5, 2.8, 2.9, 1.9, 1.7, 4.7, 3, 3.5, 3, 2.7, 3.1, 
    2.4, 2.6, 4.2, 3.5, 3.2, 3, 3, 2.9, 2.9, 2.4, 3.1, 3.5, 3.3, 3.9, 2.2, 
    1.8, 2.4, 2.5, 3, 3.1, 1.1, 0.6, 0.3, 1.6, 1, 2.8, 1.9, 1.3, 3.5, 2.3, 
    2.3, 2.3, 2.6, 2, 1.8, 0.4, 0.1, 0.3, 1, 0.4, 0.4, 0.1, 0.1, 0.6, 0.5, 
    0.3, 0.7, 0.1, 0.9, 1.2, 1.8, 1.8, 1.5, 1.5, 1.7, 2.6, 1.9, 0.6, 0.2, 
    0.3, 0.3, 0, 0, 0.4, 0.9, 0.5, 0, 0.5, 0.1, 0, 0, 0, 0.1, 0.8, 0, 1.1, 
    0.1, 0.2, 0.5, 0.8, 1.7, 1.6, 0.6, 1, 1.8, 0.1, 1, 1, 0.8, 0.5, 1.2, 0.7, 
    1.6, 1.1, 0.6, 0.7, 0.2, 0.9, 0.3, 0.6, 0.9, 0.8, 2.4, 1, 2.1, 1.3, 0.3, 
    0.1, 1.3, 1.6, 5.1, 4.6, 6.8, 5.2, 3.4, 5.8, 4.4, 0.5, 1.5, 2.2, 1, 1.3, 
    1, 1, 1.8, 1.4, 4.3, 6.2, 6.7, 5.7, 5, 3, 3.9, 4.3, 4.3, 4.1, 4.8, 3.5, 
    2.8, 3.9, 4.3, 3.6, 4.3, 4.9, 4.4, 4.3, 4.9, 4.2, 4.5, 4.1, 4.1, 5.3, 
    4.2, 4.4, 4.6, 5.2, 4.9, 6.6, 6, 6.5, 6.3, 6.3, 4.2, 5.2, 4.7, 4.8, 5.4, 
    3.3, 3, 1.7, 1, 1, 1.1, 1.1, 0.4, 0, 0.5, 1.2, 2, 0.6, 1.6, 0.5, 0.4, 
    0.4, 0.9, 0, 1.2, 1.9, 0.2, 0.1, 1.4, 0, 0.6, 1, 0.8, 0.1, 0.1, 0.6, 0, 
    0, 0.8, 2, 1, 0.8, 1, 1.5, 1.5, 1.8, 1.8, 0.9, 0.7, 1.1, 1.1, 3.9, 6.5, 
    4.6, 5.1, 2.2, 1.9, 1.5, 3.5, 3.8, 3.7, 3.2, 3.3, 2.7, 4.5, 6.5, 6.5, 
    6.7, 6, 6.3, 6.3, 4.9, 5.5, 3.7, 4.8, 5.1, 3.6, 4.5, 3.6, 3.7, 3.7, 3.5, 
    2.5, 1.5, 3.8, 2.4, 3, 3.2, 3.6, 3.3, 2.4, 2.3, 2, 0.4, 0.1, 1.6, 1.6, 0, 
    0.7, 0.8, 1.8, 1.9, 2.9, 3.1, 2.2, 2.3, 2.2, 2, 3.6, 1.2, 1.9, 3.9, 1.6, 
    3.6, 4.2, 4.8, 4.1, 0.6, 1.6, 0.6, 1, 0.3, 1, 2.7, 1.4, 0.7, 2.6, 2, 1.3, 
    1.8, 2.8, 2.3, 3.7, 4.5, 4.9, 2.9, 3.1, 2.5, 3.3, 4.1, 4.4, 5.5, 5.9, 5, 
    3.7, 4.4, 4.3, 1.9, 2.2, 1.9, 4.1, 4.6, 4.5, 4.1, 3.4, 3.7, 4, 4.2, 4, 
    4.2, 4.2, 5.1, 4.7, 4.5, 0.2, 0.1, 0.4, 0.2, 0.2, 0.1, 0.5, 0.9, 1, 1.1, 
    0.8, 1.5, 1.1, 2.7, 1.6, 1.2, 1.6, 1.3, 2.5, 2.8, 3.9, 2.1, 2.5, 2.9, 
    0.2, 1.5, 1.4, 0.3, 0.5, 0.9, 1, 0.3, 0.5, 1.8, 1.3, 1.5, 1.7, 2.6, 2.5, 
    3, 2.5, 1.9, 1.5, 1.7, 1.2, 0.5, 1, 0.8, 1.6, 1.4, 3.4, 3.9, 5, 4.8, 7.3, 
    4.7, 7.2, 6.8, 4.9, 5.3, 5, 6.4, 5.2, 4.3, 3.7, 2.6, 0.6, 1.8, 4.4, 1.7, 
    5.1, 2.6, 0.6, 3.2, 5.5, 3.5, 2.7, 4.6, 4, 4.9, 2.3, 1.4, 1.3, 1.6, 1.6, 
    0.8, 2.4, 2.5, 1.6, 0.8, 1.7, 2, 1, 2, 0.2, 1.1, 0.4, 0.2, 1.6, 0.1, 1.1, 
    1.8, 2.2, 2.6, 1.5, 0.8, 1.8, 1.7, 1.7, 0.5, 0.6, 1.9, 2.3, 1.6, 1.4, 
    0.4, 0.6, 0.3, 1, 0.7, 0, 0.6, 0.1, 0, 0.2, 0.2, 0.5, 0.1, 0.9, 1.3, 0.9, 
    0.6, 0.8, 1, 1.4, 1, 2, 3, 1.2, 1.4, 2.1, 1.4, 0.2, 0.1, 0.7, 0.4, 0.8, 
    1.4, 4.4, 0.7, 3.6, 4, 3.5, 1.9, 4.1, 6, 3.1, 4.9, 5.1, 5.2, 4.3, 4.1, 
    4.4, 5, 2.1, 2.5, 2.8, 1.4, 0.9, 0.8, 0.7, 1.5, 1.1, 0, 1.2, 0.8, 1, 0.8, 
    0.4, 0.5, 0.3, 0.9, 0.8, 0.9, 0.5, 0.4, 0.4, 0.7, 1.1, 0.6, 1.1, 1, 0.6, 
    0.4, 0.1, 0, 1.2, 1.1, 1.8, 0.2, 1.5, 1.4, 2.2, 1.7, 0.3, 0.8, 0.6, 0, 0, 
    0.8, 1.5, 1, 1, 0.1, 0, 0.2, 0, 0.3, 0.1, 0.6, 0.9, 0.7, 0, 0.3, 0.7, 
    1.2, 1.9, 1.6, 0.9, 1.1, 1.3, 1.5, 1.7, 1.4, 3.9, 5.3, 1.4, 0.5, 1.8, 
    0.1, 0.6, 0.5, 0.2, 0.3, 0.4, 0.2, 0.1, 0.7, 0.1, 0.1, 0.9, 1.2, 0.8, 1, 
    0.7, 0.7, 1.1, 0.6, 0.8, 0, 1.1, 1, 0.5, 0.6, 0.7, 0.2, 1.1, 0.7, 0, 0, 
    0.1, 0.1, 1, 0.4, 1.8, 1.2, 1.1, 1.2, 1.4, 1, 2.2, 1.5, 0.9, 0, 1.1, 1.3, 
    1, 0.1, 0.2, 0.6, 3.3, 4.6, 4.4, 3.5, 3, 3.5, 4.7, 6.1, 5.6, 6, 8.3, 6.2, 
    5.6, 7.1, 5.8, 6.6, 8.5, 6.4, 6.5, 6.4, 5.7, 5.3, 5, 3.7, 4.3, 4.5, 4.3, 
    3.6, 4.7, 5.3, 3.4, 4.3, 5, 4.3, 4.3, 3.5, 3.1, 3, 3.1, 2.9, 3.5, 2.5, 
    2.3, 0.6, 1.3, 1.3, 0.4, 0, 0, 0.3, 0, 0.5, 1.1, 0.4, 0.3, 4.5, 3.2, 2.9, 
    3.2, 3.3, 3.1, 3.2, 3.7, 3.4, 4.4, 4.7, 4.4, 3.3, 4.6, 3.8, 3.9, 4.2, 
    4.3, 4.4, 4.1, 4, 4, 3.5, 4.3, 3.5, 3.4, 3.5, 1.1, 0.4, 0.2, 0.1, 1.8, 
    0.2, 0.1, 0, 0.1, 0, 0.3, 0.2, 0.4, 0.2, 0, 0.7, 0.2, 2.3, 0.7, 0.3, 0.5, 
    0.9, 0.6, 1.6, 2.1, 1.4, 0.8, 0.6, 1.4, 1.5, 0.9, 0.8, 0.6, 0.9, 0.8, 
    0.7, 1.1, 0.2, 0.6, 0.6, 0.9, 0.8, 1.2, 2.2, 0.7, 1, 1.3, 1.5, 0.7, 1.4, 
    1.5, 1.3, 1.4, 1, 1.5, 1, 1.4, 1, 0.7, 0.7, 0.9, 0.6, 1.9, 2.8, 1, 1.3, 
    1.1, 0.7, 0.2, 4.1, 3.5, 2.8, 2.1, 0.2, 2, 4.4, 3.7, 3.4, 2.9, 4.1, 3.1, 
    2.6, 3.1, 2.6, 2.1, 1.9, 1.5, 3, 2.8, 2.6, 2.1, 1.7, 2.1, 1.8, 2.1, 3.3, 
    4.6, 5.6, 2.8, 2.8, 2.9, 1.7, 1.1, 1.7, 4, 1.6, 2.9, 3.6, 1.2, 1.5, 1.6, 
    0.2, 0.4, 1.1, 0.9, 1, 0.2, 0.7, 2, 1.8, 1.6, 1.6, 1.5, 2, 2.4, 1.6, 1, 
    0.8, 1.5, 2, 1.2, 1, 0.3, 0.7, 0.1, 0.2, 1.1, 0.5, 0, 0.3, 0.3, 0.8, 0.6, 
    1.7, 1.2, 1.4, 1.3, 1.4, 0.7, 3.2, 1.3, 0.9, 0.5, 2.2, 0.3, 0.4, 0, 0.4, 
    0.9, 0.1, 0, 0.1, 0, 0.3, 0.6, 1.3, 0.6, 0.8, 1.4, 1.2, 1.7, 0.9, 1.7, 
    1.5, 2.5, 1.5, 1.9, 1.4, 0.7, 0.9, 1.2, 3, 2.8, 2.3, 0.6, 3.1, 2.7, 2.9, 
    3.2, 3.1, 2.5, 2.2, 1.2, 1.6, 1.9, 0.9, 1, 1.4, 0.7, 1, 0.3, 1.5, 1.4, 
    0.9, 1.1, 0.8, 0.1, 0.7, 4.6, 3.7, 3.2, 2.5, 1.1, 1.9, 3.8, 3.5, 4.4, 
    6.4, 5.4, 3.7, 3.5, 2.9, 3.4, 3, 3.7, 3.2, 2.5, 3.3, 3.7, 3, 3.5, 2.5, 
    1.8, 1.6, 1.8, 1.3, 1.6, 1.4, 1.4, 1, 0.9, 0.9, 0.9, 0.4, 0.8, 1.1, 1, 
    1.6, 1.1, 1, 0.5, 0.4, 0.3, 0.1, 0, 0.2, 0.3, 0.3, 0.6, 0.5, 0.9, 0.8, 
    0.7, 1.3, 1.1, 2.1, 2.9, 0.8, 1.6, 1.3, 1.5, 1.7, 1.5, 1.3, 1, 2.3, 1.4, 
    0, 0, 1, 0.9, 0.9, 1.5, 2, 4, 2.9, 1.4, 2.3, 3.7, 4.6, 4.1, 3.8, 1.7, 
    1.7, 2.7, 2.8, 1.5, 0.2, 2.2, 0.9, 1.1, 1.7, 1.3, 1.3, 0.6, 1, 2, 1.1, 3, 
    5.9, 5.5, 5.4, 2.1, 2.2, 2.4, 3, 2.7, 2.8, 3.9, 5, 3.3, 5.1, 2.4, 1.1, 
    4.4, 1.1, 2.1, 0, 0.9, 0.3, 2.5, 1.4, 1.7, 1.1, 1.8, 4, 4, 5.7, 5.4, 5.2, 
    4.8, 4.9, 4.5, 3.7, 4.3, 4.3, 4.1, 3.3, 2.7, 4.2, 4.5, 3.3, 5, 3.6, 2, 2, 
    2.2, 2.5, 3.2, 3.5, 5.1, 4.6, 4.9, 8.7, 8.8, 4.8, 2.6, 2.7, 4.6, 5, 5.5, 
    4.8, 5.9, 6.6, 5.6, 5.9, 5.2, 3.3, 2.8, 1.5, 3.5, 2.7, 3.9, 2.8, 1.8, 
    5.4, 2.2, 3.8, 2.7, 4, 5.1, 4.7, 1.2, 2, 3.9, 2.4, 1.6, 2.3, 1.5, 0.8, 
    0.5, 1.1, 2.6, 2.5, 1.2, 2.2, 1.4, 1.9, 2.5, 2.1, 2, 2.2, 2.9, 3.4, 3.9, 
    3.3, 2.6, 2.4, 2.4, 1, 0.6, 1.3, 0.8, 1.3, 2.2, 3.1, 2.7, 1.5, 1.5, 1.1, 
    0.5, 1.6, 0.7, 2, 2.6, 1.7, 2.9, 3.7, 3.3, 2, 3.9, 4.9, 5.1, 5.3, 5.8, 
    5.2, 6, 4.1, 4.1, 4.3, 6.1, 4.4, 4.6, 4.9, 3.2, 4.7, 3.7, 3.4, 6.8, 6.3, 
    8.1, 3.2, 3.6, 5.1, 3.5, 2.4, 3.4, 2, 3.2, 1.2, 3.1, 2.9, 2.5, 3.7, 3.2, 
    3.1, 1.4, 3.8, 3.6, 4.3, 2.8, 5.1, 1.1, 4.1, 6.1, 6.8, 6, 2.1, 1.9, 2.4, 
    1.9, 2.5, 4.6, 2.3, 4.4, 3.7, 4.4, 3, 3.9, 2, 3.1, 3.4, 3.6, 1.5, 3.4, 2, 
    2.9, 2.6, 1.2, 3.6, 2.9, 4.6, 4, 4.7, 4.8, 2.9, 3.1, 3.8, 4.2, 4.3, 3, 
    0.6, 2.3, 3.9, 3.8, 2.1, 1.2, 2.8, 2.8, 3.7, 2.2, 2, 3.1, 3.1, 3.1, 3, 2, 
    2.7, 2.2, 1.5, 1, 1.4, 1.2, 1.1, 1.2, 1.8, 2, 1.6, 1.4, 1.7, 2, 2.2, 2.6, 
    2.4, 2.7, 2.6, 3.2, 3.1, 3.4, 2.8, 3.3, 2.4, 1.7, 1.6, 1.3, 1.3, 1.2, 
    1.4, 0.8, 0.6, 0.9, 1.8, 1, 1.5, 1.8, 2.2, 2.6, 2.8, 2.5, 3.8, 1.2, 1.7, 
    1.5, 1.8, 3.2, 1.7, 0.4, 0.7, 1.6, 2.6, 4.1, 3.5, 4, 4, 4.4, 2.8, 2, 2.6, 
    1.1, 1.5, 2.4, 2.5, 0.8, 0.9, 2, 3.1, 1.4, 2.6, 1.2, 1.5, 1.9, 2.1, 2.1, 
    3.2, 2.4, 1, 0.9, 0.1, 0.9, 1.6, 0.8, 1.2, 1.9, 2.4, 2.5, 2.5, 3.9, 4.9, 
    4.9, 1.9, 1.3, 2.3, 2.2, 0.9, 0, 0.3, 2.6, 2.1, 3.4, 4.1, 4.8, 3, 3, 2.5, 
    1.7, 2.3, 3, 3, 2.7, 2.5, 3, 2.9, 5, 4.3, 4, 3.7, 3.9, 2.1, 1.1, 1.7, 
    0.9, 0.5, 0.7, 1.3, 0.8, 0.2, 0.8, 1, 0.9, 0.7, 1, 1.7, 1.6, 2.2, 1.3, 
    2.1, 2.1, 2.1, 0.5, 0.8, 1.9, 1.1, 1.5, 1.4, 0.9, 0.4, 0.3, 1.7, 1.5, 
    1.5, 0.9, 1.1, 0.9, 0.4, 0.6, 1.6, 0.9, 1.3, 1.6, 2.1, 1.8, 1.7, 1.3, 
    0.9, 0.8, 0.8, 0.5, 0.1, 0, 1.1, 0.4, 0.4, 0.2, 0.2, 0.3, 0.8, 1.3, 0.4, 
    1, 3, 2.1, 2.8, 2.5, 3.2, 4.4, 3.8, 3.5, 3.5, 3.1, 3.2, 2.5, 2.6, 3.7, 
    1.9, 2.6, 2.7, 0.7, 0.9, 1.6, 1.8, 2.7, 3.1, 2, 0.8, 1.5, 1.6, 1.6, 2, 1, 
    1.3, 1.2, 1.5, 1, 0.8, 1.2, 0.7, 0.9, 0.3, 0.7, 1, 0.9, 1.5, 0.9, 0.8, 
    0.6, 1.2, 1.8, 2.6, 0.9, 2.7, 2.6, 4.3, 2, 2.6, 3.1, 3.1, 3.3, 3.8, 3.2, 
    3, 2.4, 2.5, 1, 0.4, 1.8, 1.2, 1.5, 2, 1.6, 1.9, 2.5, 2.4, 2.2, 1.6, 1.4, 
    1.5, 1.8, 1.7, 1.7, 1.6, 1.3, 1.2, 1.9, 2.4, 2.2, 2, 2.8, 1.5, 0.7, 1.5, 
    2, 1.8, 1.5, 0.8, 0.4, 1.4, 1.7, 0.6, 0.8, 0.9, 0.8, 0.3, 0.7, 0.2, 0.4, 
    0.6, 0.2, 0.4, 0.3, 0.6, 0.2, 0, 2.2, 2.7, 2.1, 2.1, 0.8, 0.6, 1.4, 1.4, 
    1, 1.4, 0.6, 1.5, 1.6, 1, 0.8, 0.6, 0.9, 1.1, 1.1, 1.3, 1.7, 1, 0.8, 1, 
    1.1, 0.4, 0.8, 0.6, 1, 1.5, 1.1, 2.4, 2.1, 2.1, 2.2, 2.3, 2.7, 2.4, 2, 
    1.9, 1.7, 1.6, 1.6, 1.1, 2.7, 3.4, 2.7, 1.9, 3.4, 3.4, 2.1, 2.3, 1.8, 
    1.5, 2, 2.6, 3.5, 4.5, 4.1, 4.1, 4.6, 2.9, 2.8, 2.6, 1, 2.4, 1.5, 1.5, 
    1.1, 2.3, 2.4, 1.9, 1.4, 1.6, 0.6, 1.9, 2.1, 2.1, 2.5, 2.4, 2.4, 2.4, 
    2.4, 1.1, 1.9, 1.4, 1.1, 1.4, 0.7, 0.7, 2.4, 1.3, 0.8, 1.3, 3.4, 1.8, 
    0.4, 0.2, 0, 1.2, 3.9, 2.1, 2.8, 2.1, 2.1, 2.6, 1.8, 2.7, 2.2, 2.2, 2.1, 
    1, 2.9, 1.3, 3.2, 2.1, 4.4, 3.2, 2.6, 2.1, 1.1, 1, 1.4, 1.7, 1.2, 0.9, 
    2.1, 1.9, 2.5, 1.3, 1.9, 1.4, 1.8, 2.1, 1.2, 3, 3.3, 2.2, 2.1, 1.7, 1.5, 
    1.3, 0, 0, 0, 0.5, 1.4, 0.7, 1.6, 0.9, 0.1, 1.2, 0.2, 0.1, 1.3, 0.6, 1.2, 
    1, 0.9, 1.1, 0.9, 2.1, 3.4, 0.4, 0.7, 0.9, 0.2, 1.7, 0.6, 0.8, 0.9, 2.7, 
    3.5, 3.2, 3.5, 3.7, 3.1, 3.2, 4.1, 4.6, 3.5, 3.9, 3.7, 3, 2.9, 2.9, 3.8, 
    3.2, 2.2, 2.1, 5, 2.8, 3.1, 1.4, 2, 1.2, 3.1, 1.4, 1.7, 0.8, 1.2, 3, 2.3, 
    2.7, 4.2, 4.2, 4.8, 6.1, 6.4, 4.4, 5.6, 4.3, 4.2, 3.7, 3.7, 3.8, 2.6, 
    3.7, 2.6, 4.8, 5.2, 5, 4.4, 5.1, 4.5, 4.3, 4.2, 4.2, 5.4, 5.7, 4.3, 4.8, 
    4.8, 5.1, 4.2, 4.5, 4.1, 3.8, 4.2, 4, 3.6, 3.3, 2.3, 4.6, 4.8, 7.6, 6.6, 
    6.2, 5.5, 3.7, 3.6, 3.6, 3.8, 3.1, 2.7, 2.1, 2.2, 2, 1.9, 1.1, 1.9, 0.6, 
    0.4, 0, 0.5, 0.3, 2.6, 2.5, 1.8, 2.1, 1.9, 2.3, 2.1, 2.2, 1.9, 2, 2.5, 
    3.1, 2.5, 2.7, 3.4, 3, 2.1, 2.1, 1.5, 1.2, 2.9, 2.2, 1.8, 1.5, 1.5, 1.3, 
    1.3, 1.9, 2.4, 2, 2.4, 2.4, 2.2, 3.2, 2.7, 2.1, 2, 2.1, 0.6, 2.3, 1.7, 
    2.8, 2.6, 2.5, 3.9, 3.1, 1.9, 1.3, 0.6, 2.7, 1.6, 0.9, 1.2, 1.2, 1.3, 
    0.4, 1.4, 1, 1.7, 2.8, 2.5, 2.5, 2.1, 2.9, 1.8, 1.1, 0.2, 0, 0, 2.2, 3, 
    1.8, 2.3, 2.7, 0.9, 1.5, 1.7, 1.2, 2.1, 2.3, 2, 2, 1.5, 0.2, 1.2, 0.6, 
    0.3, 1.9, 4.2, 3.3, 3.7, 4.7, 3.2, 3.3, 3.4, 3.2, 4.2, 4.7, 3, 3.7, 3.8, 
    4.2, 2.4, 2.3, 1.1, 4.2, 1.3, 0.8, 0.6, 1.1, 5.4, 4.4, 4.8, 2.4, 4, 4, 
    3.3, 3.1, 2.3, 2.8, 1.2, 0.8, 1.9, 2.2, 0.5, 3.1, 2.4, 2.5, 0.3, 3.5, 
    3.9, 5, 2.6, 3.1, 4.3, 3.9, 3.6, 2.4, 2.4, 3.1, 2.8, 1.4, 3.6, 3.5, 3.8, 
    3.5, 3.9, 3.9, 3.9, 1.8, 3, 3.2, 3.5, 2.3, 3.3, 2.4, 1.2, 3.6, 2.9, 1.6, 
    2.2, 1.5, 2.9, 2.6, 1, 1.5, 3.3, 2.4, 2.5, 3.2, 2.8, 3, 2.6, 2, 1.7, 2, 
    2.4, 2.5, 2.2, 1.7, 1.5, 1, 1.5, 1.2, 1, 1.9, 0.6, 0.5, 0.1, 0, 0.3, 0.4, 
    0.1, 0.1, 0.1, 1.2, 1.4, 1.1, 1, 1, 0.5, 0.4, 0, 3.7, 3.5, 1.6, 2.7, 3.4, 
    3, 3.4, 2.8, 2.6, 2.8, 0.8, 0.1, 1.1, 1.6, 2.7, 2.9, 1.6, 2, 3.1, 3.4, 
    1.2, 3, 1.5, 2.7, 1.7, 4.3, 3.9, 4.9, 4.9, 5.2, 4.7, 4.2, 3.8, 2.3, 0.7, 
    0.9, 1.7, 1, 0.9, 1.8, 1.7, 1.5, 1.9, 1.6, 1.6, 2.3, 2.4, 2.7, 3.3, 0.9, 
    1.9, 2.1, 0.9, 1, 0.8, 0.1, 1.2, 1, 0.1, 0.4, 0.2, 0.3, 0.2, 0.3, 0.4, 
    0.5, 1.6, 1.1, 1.4, 1.3, 1.8, 3.1, 2.9, 2, 0.3, 0.5, 1.3, 1.3, 1.3, 2.2, 
    2.2, 2, 1.6, 1.7, 2.5, 0.2, 1.1, 4.1, 0.7, 2.5, 3, 3.1, 3.1, 3, 1, 1.6, 
    2.3, 4.3, 0.6, 2.7, 2.4, 1.9, 0.3, 0.4, 0, 0, 0.5, 1.5, 1.4, 2.2, 2, 2.1, 
    2.5, 1.6, 0.5, 1.1, 2.1, 2.2, 1, 1.4, 1.2, 0.9, 1.6, 1.1, 0, 0.1, 0.8, 
    0.2, 0, 0.9, 1.2, 0.8, 0.9, 0.5, 0.9, 1.2, 1.5, 0.6, 1.5, 0.8, 1.6, 1.7, 
    2, 3.2, 2.1, 2.1, 1.1, 2.2, 3.2, 1.2, 0.9, 1.4, 0.2, 0.4, 0.7, 0.8, 0.8, 
    0.9, 0.8, 2.8, 5, 6, 5.6, 2.7, 1.4, 3.3, 2.6, 4.1, 2.1, 0.9, 1, 2.6, 2.5, 
    3.3, 2.9, 3.1, 3.5, 5.4, 5.1, 4.3, 3, 2, 3.8, 3.9, 2.5, 2, 6.1, 5, 5.8, 
    6.3, 3.9, 5.5, 5.3, 5.9, 4, 3.4, 3.1, 3.1, 2.9, 2.6, 0.5, 1.6, 0.7, 1.3, 
    0.5, 2.2, 0.9, 0.6, 1.2, 2.3, 4.6, 3.9, 4.1, 3.5, 2.5, 1, 3.9, 1.3, 1.4, 
    1, 0.7, 0.7, 0.8, 1, 0.7, 0.7, 1, 0, 0.3, 0.6, 0.8, 0, 0.3, 1.6, 1.6, 
    2.2, 0.9, 1.2, 3.1, 3.3, 3.3, 3.3, 3.1, 2.4, 2.1, 1.8, 1.6, 1.4, 0.9, 
    0.8, 1, 1, 0.7, 0.6, 0.2, 1.1, 0.6, 0.8, 1.1, 1, 1.1, 1.2, 1.7, 2.3, 2.3, 
    1.5, 0.6, 1, 1.1, 1.4, 1.8, 1.9, 1.7, 1.6, 1.4, 1.3, 1.4, 1.4, 1.7, 1.2, 
    0.8, 1.8, 2.2, 2.1, 2.6, 2.6, 2.8, 3, 2.9, 2.6, 2.4, 0.2, 0.7, 1.6, 2.3, 
    2.4, 2.3, 2.3, 2.3, 2.2, 2.2, 2, 2, 1.7, 1.5, 3.6, 5.2, 5.2, 5.5, 4.6, 
    4.6, 1, 1.3, 3.4, 3.9, 2.6, 2.7, 1.9, 3, 2.9, 2.5, 2.5, 1.4, 2.1, 3.5, 
    1.9, 2.3, 0.8, 1.4, 2.1, 1.7, 2.4, 2.4, 1.7, 2.8, 2.1, 2.2, 1.2, 0.6, 
    0.5, 0.8, 1.1, 0.9, 1.2, 0.5, 2, 0.8, 0.3, 0.4, 0.8, 0.7, 3, 3.3, 2.9, 
    3.2, 2.5, 2.3, 2.1, 1.2, 1.1, 2, 2.1, 2, 1, 0.9, 1.3, 1.6, 1.4, 0.9, 0.4, 
    0.5, 0.5, 0.6, 0.7, 1.4, 0.6, 1.1, 3.5, 0.9, 0.7, 0.7, 1.2, 1.5, 1.1, 
    1.3, 1.5, 1.7, 1.3, 0.4, 0.2, 0.9, 1.8, 2, 0.3, 0.3, 0, 1.5, 1.9, 2, 1.7, 
    2.6, 1, 1.1, 0.7, 0.6, 0.8, 0.9, 1.4, 1.8, 1.7, 1.7, 1.3, 1, 1.1, 0, 2.2, 
    1.7, 0.3, 0, 0, 0.3, 0.4, 0.8, 0.8, 1.1, 1.8, 1.8, 1.8, 2.8, 2.6, 3.1, 2, 
    2, 1.4, 1.5, 1.2, 1.2, 3, 3.4, 3.8, 3.9, 4, 3.8, 3.6, 3.1, 2.3, 1.2, 3.9, 
    1.7, 2.1, 1.1, 1.6, 3.3, 2.5, 2.4, 3.5, 2.8, 3, 3.6, 2.2, 5.3, 4.8, 3.3, 
    3.1, 2.7, 2.3, 1.7, 0.9, 0.2, 1.7, 1.4, 0.5, 1.8, 1.1, 1.5, 1.4, 2.7, 
    1.6, 1.3, 2, 2.1, 0.9, 0.7, 0.8, 1.1, 0, 0.1, 0.3, 0, 1.9, 1.9, 2.2, 2.3, 
    1.8, 2, 1.8, 1.7, 1.4, 1.7, 1.3, 0.9, 1.5, 1.5, 1.6, 1.4, 2.3, 1.4, 2.1, 
    2.5, 0.4, 0.7, 1, 1.8, 0.5, 1.5, 1, 0.6, 1, 0.8, 0.9, 0.6, 0.6, 0.7, 1.2, 
    1.9, 2, 1.3, 1.1, 1.2, 1.3, 3, 4.6, 6.3, 3.3, 0.2, 1.7, 0.8, 0.7, 2.6, 
    1.6, 1.3, 1.5, 1.2, 2.9, 1.8, 1.7, 1.6, 1.9, 1.9, 6.1, 5.8, 4.8, 2.2, 
    1.7, 3.7, 4.3, 1.5, 2, 1.9, 1.1, 1.5, 0.7, 3, 2.2, 2.7, 3.9, 3.8, 3.8, 
    1.2, 3.9, 1.9, 3.3, 1.8, 1, 2.6, 3.7, 4.6, 2.9, 2.8, 3.7, 4, 2.3, 1.7, 
    2.6, 4, 2.4, 1.4, 0.2, 0.4, 0.4, 1.7, 0.1, 1.1, 0.8, 1.2, 0.8, 0.8, 2.5, 
    2.1, 0.5, 5.7, 6.3, 4.6, 5.8, 0.8, 6.7, 1.2, 0.9, 0.9, 4.5, 4.1, 2.8, 
    1.1, 7.3, 6.9, 6.4, 0.9, 1.5, 4.4, 1.2, 2.6, 5.5, 2.3, 2.2, 2.1, 5.4, 
    5.3, 5.4, 5.5, 5.5, 4.9, 4, 3.2, 2.8, 2.6, 0.9, 0.1, 0.2, 1.3, 0.7, 1.5, 
    1.4, 0.9, 1.4, 1.5, 1.3, 1.9, 1.6, 1.6, 3.7, 3.4, 1.8, 3.2, 3.4, 3.4, 
    3.3, 3.1, 3.3, 3.3, 1.1, 0.4, 3.4, 3.5, 0.5, 3.4, 3.5, 0.6, 3.7, 1.4, 
    1.4, 1.6, 2.5, 3.7, 3.1, 2.6, 0.6, 0.8, 4.1, 4.3, 1.3, 1.6, 0.9, 0.6, 
    1.5, 0.1, 4.1, 4.1, 3.2, 0.1, 0.5, 2.9, 1.7, 1.4, 1.7, 2.4, 2.9, 2.7, 
    2.7, 3.1, 3.6, 4.3, 5.1, 5.9, 6.6, 7, 6.9, 6.1, 5.8, 6, 0.3, 1.1, 0.5, 
    1.3, 4.9, 1, 0.8, 1.4, 3.7, 0.8, 5.6, 5.6, 5.6, 5.6, 5.2, 5.7, 5.8, 5.9, 
    5.5, 6.7, 6.7, 4, 5.1, 6.7, 6.5, 5.9, 3.5, 6.5, 4.6, 4.4, 6, 6.3, 5.5, 
    4.8, 5.7, 4.8, 4.9, 4.8, 4.1, 4.1, 4.4, 4.5, 2.5, 2.5, 4.3, 0.6, 0.8, 
    1.5, 0.6, 0, 3.6, 1.3, 3.2, 2.9, 2.9, 4, 4.2, 4.2, 3.5, 1.3, 1.7, 1.2, 
    0.4, 3.1, 3.1, 2.1, 2.7, 0, 0.3, 0.1, 0.5, 1.5, 0, 0, 1.7, 0.9, 1.4, 1.6, 
    1.7, 1.5, 1.4, 1.5, 1.8, 1.7, 1.8, 2.5, 0.7, 1.2, 0.1, 0.2, 0, 0.1, 0.5, 
    1.2, 2.4, 2.3, 0, 1.8, 2.6, 2.8, 2.1, 1.7, 2.7, 3.1, 1.7, 2, 1.3, 1, 1.7, 
    1.4, 1.5, 0.8, 0.4, 1.6, 1.8, 1.2, 1.2, 2, 0.1, 0.2, 0.4, 0, 0.8, 1, 0.8, 
    1.2, 0.9, 1, 0.6, 0.9, 3.3, 1.2, 0.7, 0, 0.3, 0.6, 0.9, 0.7, 0.8, 1.8, 
    4.6, 0.3, 0.4, 2.5, 1.5, 0.7, 0.3, 0.8, 0.2, 0.7, 0.1, 0.7, 1.2, 1.2, 
    0.9, 4.1, 8, 7.3, 4.8, 5.2, 5.3, 5.4, 5.6, 4.4, 6.3, 6, 5.6, 4.5, 4.7, 
    5.8, 5.6, 5.8, 6.3, 6.9, 6.7, 6.4, 6, 5.7, 4.3, 5.1, 5.6, 6.3, 4.2, 4.3, 
    4.3, 3, 4.9, 4.5, 1.2, 2.6, 2.5, 2.3, 2.8, 3.1, 3.3, 3.5, 2.8, 3.7, 3, 
    1.8, 2.2, 0.9, 3, 4, 3.6, 2.9, 3.3, 0.7, 1.6, 0.1, 1.5, 2.2, 2.6, 1.4, 
    2.6, 3.6, 3.2, 2.8, 1.8, 5, 4.2, 5, 4.2, 6.3, 6.3, 4.8, 5.3, 5.6, 4.8, 6, 
    4.5, 5.2, 3.9, 2.6, 2.8, 3.5, 2.7, 2.3, 2, 0.7, 1.1, 0.4, 0.4, 0.8, 1.9, 
    5.4, 5, 4.9, 4.2, 3.5, 5.2, 3.3, 1.8, 1.8, 1.5, 0.4, 1, 0.4, 0.5, 0, 1.1, 
    0, 0.3, 0.6, 0.6, 0.5, 0.2, 0.2, 1.2, 2.1, 2, 1.6, 2.9, 5.2, 4.5, 5.7, 
    5.9, 6.1, 5.2, 5.6, 6, 7.4, 7.7, 6.6, 6.8, 6.7, 6, 6.3, 6, 6.5, 6.5, 6.5, 
    6.2, 5.8, 6.8, 7.2, 6.4, 5.8, 5.3, 5.1, 5.3, 5.3, 5.2, 5.2, 5.2, 5.1, 
    5.1, 5, 5, 5, 4.9, 4.9, 3.8, 4.4, 5.6, 5.6, 4.6, 4.3, 4.6, 3.2, 3.1, 2.9, 
    2.8, 2.7, 2.5, 2.4, 2.2, 2.1, 0.3, 2, 1.4, 2.5, 3, 2.9, 2.4, 1.7, 1.4, 
    2.5, 0.3, 0.2, 0.5, 0.5, 0.5, 1.9, 1.8, 1.4, 2.3, 2.6, 2.5, 2.7, 2.7, 3, 
    0.5, 0.8, 0.3, 0.4, 1.3, 1.2, 2.4, 1.2, 1.9, 3.9, 4.5, 4.8, 4.1, 0.8, 
    1.1, 0.3, 0.5, 0.3, 2, 1.2, 0.5, 1.6, 1.6, 1.2, 1.6, 2.8, 1.5, 2.9, 9.9, 
    9.3, 9.3, 8.5, 8.6, 10.7, 9.8, 9.3, 9, 8.8, 8.4, 4.6, 6.6, 5.8, 3.1, 3.3, 
    3.1, 1.9, 4.6, 1.9, 2.3, 2.1, 2.6, 1.2, 0.4, 0.8, 0.2, 0.3, 0.4, 0.4, 
    0.9, 1.2, 0, 0.3, 0.7, 0.8, 1, 1.6, 0, 0.4, 0, 1.8, 1.9, 1.2, 1.3, 0.9, 
    0.6, 0.7, 0.8, 2.6, 1.6, 3.2, 0.5, 1.3, 0.8, 1.5, 1.4, 1, 0.8, 1.8, 3.8, 
    1.4, 0.1, 0.3, 0.4, 0.3, 0.5, 0.1, 1.6, 2.2, 2.5, 2.5, 2.4, 2.8, 2.7, 
    0.8, 0.6, 0.4, 0.6, 0.2, 2, 2.4, 1.8, 1.7, 2.2, 1.9, 2.2, 2, 1.8, 0.1, 
    1.1, 1, 0.6, 0.6, 1.1, 1.8, 2.1, 2.4, 2.5, 2.4, 0.9, 0.9, 1, 0.7, 1, 1.9, 
    0.7, 1.4, 0.4, 1.8, 0.9, 0.4, 0.6, 0.1, 1.6, 3, 2.2, 1.6, 4, 3.8, 3.3, 
    3.9, 2.5, 2.2, 2.4, 0.3, 0.8, 0.9, 0.3, 1, 1, 0.9, 1.1, 1, 0.3, 0.6, 0.1, 
    1.8, 5.1, 5.4, 5.4, 0.2, 0.7, 0.8, 2, 1, 1.3, 0.8, 2, 6.4, 7.2, 6.6, 0.8, 
    2, 1.6, 2.2, 1.5, 0.7, 1.1, 3.4, 5.9, 7.5, 7.6, 4.6, 4.1, 4.2, 3.3, 5.5, 
    6.2, 5.9, 8.1, 6.3, 7.6, 6.5, 7.7, 6.9, 5, 7.1, 5.9, 6, 5.4, 6.2, 7.7, 
    5.2, 6.3, 7.1, 4.7, 4.9, 4.1, 4.7, 3.6, 2.2, 2.3, 4.7, 4.8, 1.4, 0.3, 
    2.3, 0.8, 0.1, 1.3, 0.9, 0.4, 0.7, 0.9, 0.2, 0, 0.7, 0.6, 0.3, 2.5, 2.6, 
    2.9, 3.2, 0.3, 1.4, 1.3, 1.2, 2.9, 2, 0.4, 0.5, 0.4, 3.4, 3.8, 0.5, 0.1, 
    0.3, 0.5, 0.7, 1.3, 1.5, 7.7, 5.7, 6.2, 7.1, 2.9, 8.2, 7.2, 10.9, 7.1, 
    8.4, 6.9, 5.3, 4.5, 4.7, 7, 6.6, 5.9, 6.1, 5.5, 5.9, 6.4, 7, 7.5, 5.5, 
    4.9, 10.7, 10.5, 6.7, 5.5, 5.2, 5.4, 3.6, 5.2, 4.1, 4.8, 6.2, 10.8, 10.5, 
    7.6, 5.8, 3.8, 4.3, 4.9, 7.8, 6.3, 7.6, 9.6, 9.5, 9.7, 9.6, 9.6, 9.5, 
    9.5, 10.1, 4, 10.3, 3.3, 4.2, 4, 5.4, 4.6, 4.2, 5, 7.8, 4.6, 4.8, 4.4, 
    4.4, 4.9, 1.5, 3.5, 3.2, 1.8, 4.7, 3.5, 3.6, 3.6, 3.5, 0.9, 3.7, 1.4, 
    3.9, 0.9, 3.7, 3.8, 3.5, 1.4, 3.5, 1.8, 0.5, 3.3, 3.4, 2.3, 1.7, 3.9, 
    4.8, 1.1, 3.8, 1.8, 1.2, 6.5, 4.4, 6.6, 4.7, 4.3, 7.3, 2, 1.7, 2.5, 1.5, 
    3.1, 1.1, 5.7, 5.5, 5.4, 5.5, 5.5, 5.4, 5.3, 2.6, 0.7, 0.6, 0.4, 1.1, 
    1.1, 3, 1.1, 2.2, 1.6, 1.1, 1.5, 1.2, 1.1, 0.9, 1.4, 0.7, 0, 0, 0.2, 2.9, 
    2.9, 2.8, 2.8, 0.3, 0.5, 0.9, 0.7, 3.4, 1.1, 1.7, 1.9, 3.3, 3.6, 0.7, 1, 
    0.7, 1.7, 0.4, 3.8, 3.9, 1.8, 4.7, 4.4, 1.1, 1.4, 1, 1.3, 1.9, 2.8, 3.8, 
    2, 2.6, 1.8, 4.4, 1.8, 1.6, 4.3, 1.9, 3.8, 3.6, 4.1, 1.5, 2.9, 1.9, 3.9, 
    3, 4.7, 4.8, 3.1, 1.3, 4.2, 2, 3.4, 4.1, 2.5, 3.4, 3.4, 3.3, 3.3, 3.7, 
    3.3, 1.2, 1, 2.7, 0.4, 1.3, 1.3, 2.8, 0.4, 0.2, 2.5, 0.6, 4.3, 4.5, 3.9, 
    3.5, 3, 4.4, 4, 1.3, 1.7, 1.2, 0.9, 0.8, 2.7, 2.7, 2.6, 1.3, 1.4, 2.6, 
    4.4, 4.4, 3.8, 3.9, 2.1, 2.7, 2.3, 4.8, 4.9, 3.6, 1.8, 3.3, 3.6, 2, 4.1, 
    1.9, 4, 2, 5, 1.9, 5, 2.5, 2.5, 1.1, 2.9, 4.4, 7.2, 7.3, 6.2, 3.4, 5.7, 
    2.7, 7.3, 7.3, 7.3, 1.7, 6.6, 1.2, 1.5, 6.2, 6.2, 1.1, 0.7, 1, 1.1, 0.2, 
    0.4, 0.5, 0.9, 0.2, 0.9, 4.1, 4.2, 4.2, 3.5, 1.9, 2.4, 3, 2.5, 4.5, 4, 3, 
    4.8, 4.8, 4.8, 0.7, 0.4, 1.2, 3.7, 3.7, 0.5, 0.1, 0.3, 3, 0.5, 0.2, 0.7, 
    0.5, 0.9, 3.1, 0.8, 0.5, 0.5, 3.1, 0.1, 0.2, 0.4, 0.7, 0.6, 1.6, 2.5, 
    1.7, 1.3, 2.9, 2.7, 2.5, 4.1, 2.7, 2.2, 0.6, 4, 2.5, 1, 1.9, 4.8, 4.5, 
    4.1, 4.1, 3.7, 1.7, 1.8, 3.2, 1.5, 2.7, 2.7, 1.8, 1.2, 1.2, 1.4, 0.6, 
    1.1, 1.4, 1.4, 2.6, 1.6, 3.1, 0.5, 0, 1.3, 1.1, 1.3, 1, 1.1, 0.7, 5.8, 
    3.7, 5.8, 6.3, 6, 5.5, 4.9, 3.7, 1.7, 2.9, 2.5, 0.9, 0.7, 0.4, 0.5, 0.5, 
    0.8, 1, 0, 0.9, 0.8, 0.8, 0.4, 1.7, 2.3, 2.5, 0.2, 1.3, 4.9, 1, 1, 1.4, 
    1.7, 0.3, 0.5, 0.4, 1.1, 0.7, 2.6, 2.1, 0.6, 3.1, 1.1, 0.6, 0.6, 1.1, 
    6.3, 4.4, 7, 7.1, 6, 7.8, 7.2, 8.5, 7.9, 9.8, 9.7, 9.4, 9.3, 9.3, 8.1, 
    5.7, 6.5, 3.5, 2.2, 3.2, 1.3, 1.6, 0.4, 4.7, 5.2, 0.7, 5, 5.2, 1.5, 1.8, 
    4, 1.4, 6.7, 4.7, 4.7, 3.6, 3.4, 2.9, 2.9, 2.6, 2.7, 2.6, 2.5, 4, 2, 1.3, 
    1.4, 1.4, 2.2, 1.5, 1.5, 1.2, 4.4, 1.7, 1, 3.7, 2.4, 4.2, 3.2, 4, 4.8, 
    4.8, 4.9, 5.3, 3.8, 6, 3.7, 6.4, 4.8, 4.4, 6.7, 5.3, 6.7, 5.9, 7, 6.5, 
    6.8, 6.6, 4.6, 5.1, 4.1, 4.7, 4, 3.5, 3.5, 3.3, 4.1, 4.1, 1.8, 3.9, 0.7, 
    1.3, 1.1, 1.4, 3, 1.4, 3.7, 1.4, 6.4, 6.3, 5.8, 5.4, 5, 1, 1.4, 0.7, 0.7, 
    1.2, 0.7, 0.7, 0.3, 1.4, 0.6, 1.2, 1.3, 1.3, 0.9, 1.5, 1.8, 1.9, 2.1, 
    0.7, 0.7, 0.6, 1.4, 2, 0, 1.4, 1.8, 2, 1.7, 1.4, 1.2, 0.5, 0.7, 1.3, 0.8, 
    0.3, 0, 0.5, 0.3, 0.8, 0.4, 0.4, 1.9, 2.1, 2.3, 2.4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.8, 0, 0, 0, 0.2, 1.2, 1.1, 1.4, 0.9, 0.2, 0.9, 1.2, 0.6, 0.3, 
    0.6, 1.9, 0.3, 0.2, 0.8, 0.9, 4.8, 0.9, 0.7, 1.2, 1.1, 0, 0.7, 0.7, 0.2, 
    0, 2.4, 0.6, 1.2, 0.6, 1.9, 0.8, 2.2, 0.7, 0.6, 0.4, 2.3, 0.5, 0.1, 0.5, 
    0.7, 0.2, 0.7, 0.2, 1.5, 0.1, 0.6, 0.7, 0.5, 1.9, 1, 0.7, 1.3, 0.6, 1.1, 
    1.6, 1.7, 1.6, 2.5, 1.4, 1.1, 1.4, 0.2, 0.6, 0.6, 0.4, 1.4, 1.2, 0.7, 
    0.6, 0.8, 0.9, 0.9, 0.7, 1.1, 1, 3.2, 3.4, 1.3, 1.4, 0.8, 0.8, 0.8, 1.2, 
    2.7, 2.4, 2.8, 3.6, 3.7, 3.7, 2.2, 1.8, 1.7, 1.3, 1.1, 0.7, 1.2, 1.3, 
    2.1, 2.9, 2.8, 1.4, 2.5, 5.7, 4.7, 6.6, 6.5, 5.9, 4.8, 5.4, 1.9, 1.7, 1, 
    0.7, 2.3, 0.8, 1, 0.6, 1, 0.8, 2.9, 0.9, 0.4, 1.2, 0.5, 0.5, 1, 0.5, 0.9, 
    0.2, 1.9, 2, 1.9, 1.3, 0.2, 0.4, 0.3, 1.4, 0.4, 1, 2.2, 0.7, 0.3, 2.9, 
    1.2, 1.9, 1.5, 4.7, 4.8, 5.4, 5.7, 6.1, 4.6, 4.7, 4.1, 5.6, 4.1, 5.6, 
    5.4, 3.7, 4.8, 5, 4.3, 4.5, 4.8, 4.5, 1.8, 1.6, 1.1, 0.8, 0.2, 1.5, 0.6, 
    6.7, 6.2, 4.1, 2.4, 1.7, 2, 2.8, 2.9, 2.3, 1.6, 1.7, 1.4, 2.5, 2.7, 2.5, 
    1.4, 3, 2.9, 2.7, 2.7, 0.5, 1.4, 1.8, 1.3, 1, 0.7, 0.6, 1, 2.2, 1.5, 1.3, 
    0.5, 2.1, 1.1, 1, 1.3, 1.3, 1.3, 2, 1.8, 2, 1.6, 1.2, 2.4, 1.4, 1.4, 1.5, 
    1.6, 2.5, 2.4, 3.1, 3, 3.1, 3.1, 0.7, 1.2, 1.6, 1.2, 1.1, 1.3, 0.2, 0.4, 
    2.7, 2.3, 1.2, 0.1, 0.3, 0.9, 0.9, 0.4, 0.3, 0.1, 0.5, 1.8, 0.7, 0.2, 1, 
    0.7, 0.8, 0.2, 0.1, 0.5, 1.5, 0.5, 0.6, 0.2, 1.3, 0.9, 0.5, 2.1, 2.7, 
    1.7, 0.4, 0.5, 1.4, 1.3, 1.7, 1.5, 2.2, 2.5, 2.6, 3.1, 1.9, 0.2, 0.3, 
    0.1, 0.1, 0.8, 1.7, 0.9, 1.4, 6.6, 6.6, 6.1, 5.6, 1.8, 0.7, 1.3, 0.6, 
    1.8, 1.1, 1.2, 0.5, 5.8, 5.7, 5.4, 5.3, 5.4, 5, 5.1, 5.5, 6, 0.9, 0.6, 
    1.2, 1.4, 1.3, 1.7, 0.8, 3.4, 1.2, 4.5, 4.2, 0.5, 0.5, 1, 1.7, 0.5, 0.9, 
    1.7, 1.6, 4.5, 4.8, 5, 5, 3.7, 6.7, 5.9, 4.4, 3.6, 1.8, 1.7, 2.5, 2.5, 
    5.8, 1.4, 6.4, 5.8, 5.7, 4.1, 5.2, 5.1, 5.3, 5.1, 6.1, 6.7, 7.2, 8.2, 
    9.1, 9.1, 8.8, 6.6, 6.4, 5.6, 3, 7, 7.4, 1.9, 1.8, 0.6, 1.4, 0.4, 0.6, 
    1.6, 0.4, 0.4, 4.4, 4.9, 4.5, 5.3, 4.8, 4.9, 5.6, 6.7, 7.5, 7.1, 7.6, 
    5.6, 7.9, 6.9, 7.1, 9.1, 8.4, 6.5, 6.9, 7.3, 5.4, 4.7, 4.8, 4.8, 3.7, 
    4.6, 5.1, 2.5, 5, 4.3, 5.1, 5.2, 3.3, 4, 5.8, 6.8, 4.8, 5.7, 4, 4.8, 5.3, 
    5.7, 7.5, 8.1, 7.1, 6.5, 6.9, 6.8, 8.3, 7.9, 9.5, 8.6, 7.6, 6.3, 8.3, 
    6.3, 6.2, 7, 8.7, 8.7, 9, 8.9, 9.1, 9, 10, 9.9, 8.7, 9.5, 8.8, 10.6, 6.2, 
    8.9, 8.5, 7.2, 5.7, 5.5, 5.7, 5.8, 5.6, 8.2, 7.9, 6.7, 7.7, 7.1, 7.3, 
    7.1, 6.7, 4.9, 5.6, 6.7, 6.9, 5.1, 6, 4.4, 5.6, 3.8, 5.5, 4.7, 4.2, 5.4, 
    4.6, 4.1, 2.8, 2.6, 3.2, 3.3, 2.8, 1.9, 1.8, 1.6, 1, 1.5, 1, 0.8, 0.7, 2, 
    0, 0, 0.8, 0.5, 0.6, 0.9, 1.4, 0.8, 0.7, 1, 1.7, 2.2, 0.3, 1.5, 0.2, 1.6, 
    0.9, 0.6, 1.6, 1.3, 0.9, 1, 1.5, 2.4, 0.1, 0.4, 1.1, 0.8, 0.5, 1, 0.1, 
    0.9, 0, 0.6, 0.6, 0, 0.1, 2, 0.2, 0.6, 0.9, 0.9, 1.3, 1.2, 0.4, 1.4, 1.1, 
    0.3, 0.7, 0.7, 0.4, 0.2, 0.2, 0.3, 0.1, 0.2, 1.1, 0.5, 0.8, 0.9, 1.2, 
    1.1, 0.7, 0.7, 0.4, 2.8, 1.3, 2.5, 3, 2.9, 3.1, 5.3, 4.5, 4.2, 3.1, 1.5, 
    1.3, 3.6, 1.1, 1, 0.1, 1.6, 1.9, 3.3, 1.8, 1.9, 2.8, 2.2, 0.9, 2.7, 1.5, 
    2, 1.9, 0.7, 0.7, 2, 0.9, 0.4, 1, 2, 0.8, 1.7, 0.5, 0.6, 0.7, 0.8, 2.6, 
    1, 1.5, 1.3, 0.9, 1.5, 1.5, 3.7, 2, 1.5, 0.7, 0.8, 1.4, 1, 1.7, 1.4, 2, 
    1.8, 1.1, 2.3, 1.9, 1, 1.5, 2, 0.7, 0.8, 1.2, 0, 1.3, 2.6, 1.1, 1.6, 1.1, 
    0.8, 3.5, 0.8, 0.8, 1.6, 0.9, 3.2, 0.7, 1.4, 1.3, 0.4, 0.5, 0.9, 1.4, 
    1.4, 1.3, 2, 2.4, 1.8, 2.3, 1.7, 1.8, 1.8, 1.2, 2.6, 0.9, 0.9, 1.6, 2.1, 
    1.2, 2, 1, 0.6, 1.2, 1.1, 0.5, 0.8, 1.2, 0.9, 5.9, 6, 6.1, 6.3, 6.4, 5.5, 
    6, 4.6, 3, 0.9, 0.9, 1.4, 0.5, 1.2, 3.2, 3.6, 5.5, 1.6, 2, 5.6, 8.6, 7.4, 
    7.8, 6.9, 8.3, 7.3, 7.9, 5.4, 2.6, 4.6, 6.9, 2.9, 2.3, 2.7, 3.7, 5.4, 
    3.1, 3.4, 6.6, 6.4, 8.2, 6.1, 7.8, 7.9, 8.3, 8.8, 9.3, 9.2, 8, 5.6, 9.9, 
    10.3, 7.9, 5.8, 5.7, 6.8, 6.7, 6.4, 9.4, 9.2, 8.4, 8.5, 7.5, 6.9, 7.5, 
    6.7, 7.5, 5.9, 3.8, 2.1, 1.8, 0.9, 2.8, 3.5, 3.1, 1.3, 0.9, 1.6, 1.8, 
    1.5, 0.5, 0.7, 2.7, 1.1, 3.4, 1.9, 3, 2.6, 2.8, 1.9, 1.7, 1.7, 0.8, 2, 
    1.9, 2.7, 0.7, 0.4, 0.9, 1, 0.6, 6.4, 5.6, 2.2, 1.2, 0.5, 1.5, 2.2, 2.6, 
    2.7, 2.8, 1.4, 1.6, 2.3, 1.8, 2.5, 1.6, 1.4, 2.4, 3, 2.2, 0.9, 0.5, 1.2, 
    1.5, 1.8, 1.7, 1.3, 0.5, 0.8, 1.3, 3.6, 1.4, 0.9, 1.9, 1.9, 3.2, 1.8, 
    2.5, 0.3, 2.3, 1.8, 3, 1.9, 3.1, 1.7, 1.3, 0.8, 1.7, 2.5, 1, 1.2, 1.4, 
    0.9, 0.4, 1.9, 1.3, 1.4, 1.5, 1.1, 0.5, 1, 0.7, 1.9, 2.2, 1.4, 1, 1.8, 
    0.9, 1.7, 2, 1.9, 1.8, 1.4, 1.4, 1.2, 1, 1.8, 0.1, 2.1, 2.1, 1.8, 1.5, 
    1.1, 1.6, 1, 1.5, 1.3, 0.8, 1.1, 0.3, 0.4, 0.9, 2.7, 1.5, 6.3, 4.8, 4.9, 
    6.4, 6.7, 7.7, 6.5, 4.8, 4.9, 5.5, 4.7, 4.6, 3.7, 4.2, 6.2, 3.5, 0.8, 
    0.8, 1.2, 3.6, 1.2, 1.1, 2.5, 1.3, 2, 1.6, 0.6, 0.6, 1.5, 1.1, 1.7, 1.4, 
    0.3, 0.8, 1.2, 1.2, 0.6, 2.4, 1.8, 1.3, 1.5, 1.2, 0.4, 3.9, 1.5, 1, 0.1, 
    2.6, 0.6, 1, 0.6, 0.7, 0, 0.7, 1.4, 0.6, 0.3, 0.3, 0.8, 0.1, 2.5, 4.5, 
    3.8, 2.5, 1.9, 1.1, 0.7, 0.6, 1.5, 1.4, 2.4, 2.6, 1.7, 1.5, 0.9, 0.5, 
    0.2, 2, 2.4, 0.6, 0.5, 0.9, 0.6, 0.9, 1.2, 0.4, 0.6, 1, 2.5, 2.8, 0.8, 
    4.4, 0.5, 0.4, 0.2, 0.5, 0.5, 1, 0.9, 0.8, 1.3, 2.3, 6.8, 9.2, 6.9, 5.3, 
    1.7, 1.2, 1.7, 1.1, 0.4, 0.4, 0.8, 1.4, 1.1, 0.8, 1.1, 0.3, 0.8, 0.6, 
    0.8, 1.1, 1.3, 0.8, 0.6, 1.2, 1.5, 1.4, 1.1, 1.4, 2.1, 2.3, 1.4, 4.2, 
    4.5, 2.8, 4, 2.5, 1.5, 1.6, 1.9, 1.3, 2.2, 0.6, 1.8, 1.5, 1, 0, 1.3, 0.1, 
    1.3, 1.5, 2, 0.2, 0.2, 0.7, 1.2, 0.1, 0.3, 1.1, 0.2, 0.6, 0, 0.4, 0.9, 
    1.6, 0.1, 0.4, 0.3, 0.9, 1.6, 3.2, 0.4, 0.7, 6.8, 8.9, 5.7, 5.6, 3.5, 
    3.7, 3.3, 4.1, 2.4, 2, 5.5, 4.8, 4.3, 6.7, 5.9, 5.9, 6.1, 4.1, 3.9, 5.9, 
    5.3, 5.5, 4.2, 5.9, 5.3, 5.4, 6.5, 6.2, 9.4, 6.6, 6.7, 7.4, 8.2, 8.7, 
    7.8, 6, 3.8, 4.9, 4.8, 4.1, 6.9, 5.3, 3.8, 2, 2, 0.8, 0.8, 0.4, 1.3, 0.8, 
    0.8, 1.3, 0.4, 0.5, 0.9, 0.7, 1.6, 1.6, 2.3, 2, 2.2, 2.3, 0, 0.2, 0.5, 
    0.1, 0.5, 0.5, 0.9, 0, 0.7, 0.1, 2.3, 1.4, 0.5, 0.4, 0.4, 0.3, 0.8, 0.5, 
    1.2, 0.1, 1.2, 0.1, 0.8, 0.3, 1.4, 0.4, 1.3, 1, 0.6, 1.4, 0.6, 2, 2.4, 
    3.5, 1.9, 0.7, 2.1, 2.2, 1.5, 0.8, 1.3, 1.8, 0.6, 1.2, 0.3, 0.4, 1, 0.9, 
    0.5, 0.2, 1.3, 0.7, 1.1, 0.7, 0.5, 0.6, 0.9, 1.8, 2.8, 1, 1.3, 1.3, 1.5, 
    2.5, 3, 3.9, 2.5, 2.2, 2.4, 1.2, 5, 1.7, 2.3, 2.1, 1.7, 1.5, 1.5, 2.5, 
    2.2, 0.7, 0.4, 2.3, 2.8, 1, 0.5, 1.1, 2.7, 6.6, 5.5, 7.1, 6.2, 4.8, 3.4, 
    2.2, 0.8, 2.1, 1.9, 2.4, 2.4, 1.4, 1.9, 0.8, 0.5, 0.9, 1, 2.1, 1.4, 2.3, 
    2.6, 0.8, 1.9, 1.1, 2.1, 1.8, 1, 0.3, 1.9, 0.2, 1.2, 0.3, 0.1, 1.8, 0, 
    0.9, 0.8, 0.3, 1.1, 0.7, 2.5, 1, 2.2, 0.6, 0.2, 0.4, 0.1, 0.4, 0.7, 0.7, 
    0.9, 0.2, 0.2, 0.3, 0.4, 0.1, 0.8, 0.3, 0, 0.5, 0.9, 1.3, 0.8, 2.4, 1.5, 
    0.7, 1.9, 1.6, 1.5, 3.8, 7.6, 4.5, 8.2, 7.3, 4.2, 3.9, 5.4, 2.3, 4.9, 
    4.6, 4.6, 5.2, 6.9, 7.9, 9.9, 10.6, 10.2, 10.7, 10.1, 11.6, 12.2, 12.8, 
    13.7, 13.3, 14.1, 12.7, 12.6, 12, 11.5, 11.6, 10.8, 10.6, 10, 11.1, 10.8, 
    10.6, 11.1, 10.9, 8.8, 7.5, 7.4, 10.3, 9.2, 10.6, 6.7, 5.7, 8, 5.1, 7.7, 
    6.7, 7.8, 6, 8.6, 10.5, 8.4, 9.4, 9.9, 5.8, 5.5, 7.9, 7.9, 5.1, 5.9, 5.2, 
    7.3, 4.8, 6.9, 4.7, 4, 2.3, 1.6, 1.1, 1.2, 0.2, 0.2, 0.8, 0.7, 0.6, 1, 
    1.4, 1.1, 0.2, 1.2, 0.3, 0.5, 1, 0.9, 0.9, 1.1, 1.1, 1.1, 3.1, 8.8, 8.7, 
    8.9, 9.5, 10.6, 8, 7.7, 7, 6.9, 8.3, 9.3, 10.1, 9.5, 11.2, 9.9, 10.8, 
    9.5, 9.2, 9.2, 8.5, 8.4, 7.3, 5.2, 3.9, 4.2, 6.1, 2.3, 2, 2.7, 1.6, 2.9, 
    4.3, 3.5, 1.7, 4, 2.9, 5.4, 5.2, 5.4, 2.9, 6.2, 6.2, 7.9, 8.7, 9.4, 5.8, 
    7, 3.9, 2.6, 3.3, 4.6, 8.6, 5.6, 7.4, 7, 6.5, 6.3, 6.1, 4.3, 4.9, 5.5, 
    2.3, 4.4, 5.8, 6.3, 4.6, 4.1, 4.5, 3.3, 5.3, 6.5, 4.6, 6.5, 5.3, 7.7, 
    5.4, 6.8, 7, 7.3, 7.3, 6.2, 7.1, 5.9, 5.9, 6.1, 4.7, 3.7, 3.4, 1, 0.7, 1, 
    1.3, 2, 3.3, 3.5, 3.2, 2.2, 1.9, 1.7, 1.1, 0.5, 0.8, 1.5, 0.5, 2.4, 2.4, 
    0.6, 0.6, 0.6, 1.4, 1.7, 0.8, 0.8, 1.4, 1.5, 1.5, 1.4, 2.1, 0.7, 0.3, 
    0.7, 0.9, 0.9, 1.3, 0.9, 1.3, 0.4, 0.7, 0.5, 0.6, 0.8, 0.7, 0.6, 1.4, 1, 
    1.1, 4.1, 1.6, 4.6, 5.7, 8.4, 7.2, 7.4, 4.3, 4.5, 5, 5.6, 3.1, 4.5, 6.5, 
    6.8, 6.8, 6.7, 6, 8, 9.9, 9, 7.7, 9.1, 6.5, 2.7, 2.3, 0.6, 0.7, 1.7, 1.2, 
    1.1, 1.8, 1.4, 2.7, 2, 1.5, 0.3, 0.6, 0.7, 0.7, 0.8, 0.5, 0.6, 1.1, 1.1, 
    0.7, 1.4, 2.4, 3, 3.3, 4.1, 1.9, 5.2, 3.4, 3.6, 4.5, 3.9, 4.2, 4.4, 4.3, 
    4.9, 4.1, 5.1, 4.7, 4, 3.5, 2.7, 3.4, 3.1, 1.5, 2, 1.6, 0.9, 0.5, 2, 1.4, 
    1, 1.1, 1.1, 0.9, 1, 2.1, 0.6, 0.7, 0.5, 0.1, 1.8, 0.4, 0.1, 0.4, 0.2, 
    0.3, 0.2, 0.3, 1, 0.9, 1, 0.1, 0.9, 0.5, 0.4, 2.1, 1.4, 2.6, 2.6, 3.3, 
    3.3, 3.5, 3.8, 4, 4.4, 3.8, 5.1, 3.5, 4.2, 5.8, 5.5, 4.4, 5.3, 4.5, 5.1, 
    4.1, 3.7, 3.2, 3.3, 3.7, 3.5, 3.9, 2.2, 3.3, 2.1, 1.3, 3.6, 0.5, 0.7, 
    0.2, 0.8, 0.6, 0.1, 4.2, 3.4, 1.8, 3.5, 3.5, 4.7, 4.5, 4.6, 6.1, 5.6, 
    5.7, 4.1, 4.5, 4.7, 3.2, 4.1, 4.4, 3.8, 6.3, 4.9, 4.7, 5.8, 5.4, 1.6, 
    0.5, 1, 0.6, 0.7, 1.1, 1, 1.2, 1.5, 1.3, 2, 0.6, 1.6, 2, 2.1, 1.8, 1.6, 
    0.3, 0.8, 2.3, 0.6, 0.8, 1, 2.9, 2.3, 2.3, 0.8, 3.7, 2.5, 2.4, 1.8, 1, 
    1.9, 1.3, 1, 1.2, 4.8, 3.5, 3.7, 3.7, 4.3, 3.4, 1.5, 1.8, 0.8, 4.9, 5.5, 
    5.2, 2.2, 2.5, 2.7, 2, 0.8, 2.1, 4.7, 4.8, 6.6, 5.8, 8.2, 8.1, 4.8, 4.6, 
    1.4, 1.9, 1.7, 1.8, 1.1, 1.3, 1.2, 1.4, 1.8, 1.2, 2, 1.2, 2.1, 1.1, 0.8, 
    0.8, 1.6, 0.4, 1.4, 0.9, 0.7, 0.7, 0.9, 1.1, 1.2, 0.5, 0.9, 0.4, 0.9, 
    0.9, 1.3, 0.9, 0.5, 0.7, 0.2, 0.7, 1, 0.9, 0.5, 1.2, 0.3, 1.4, 1.5, 0.3, 
    0.1, 0.8, 0.7, 0.4, 0.7, 0.1, 0.7, 0.3, 0.8, 0.4, 0.6, 0.7, 0.7, 0.2, 
    1.4, 1, 1, 0.9, 1.5, 0.8, 1.6, 0.7, 0.5, 1.3, 1.6, 1.1, 2.1, 0.7, 1.3, 
    0.6, 2, 1.7, 2.3, 1.1, 1.9, 1.6, 1.2, 1.4, 1.2, 1.3, 0.7, 1, 1.3, 0.7, 
    1.4, 1.2, 1.6, 2.2, 1, 0.9, 2.8, 0.9, 1.2, 0.5, 0.9, 0.9, 0.8, 1, 2.8, 
    1.2, 2.4, 1.7, 5, 2.8, 1.7, 3.1, 1.3, 1.6, 5.4, 2.2, 1.5, 5.7, 6.2, 6, 
    5.6, 4.6, 2.9, 1.6, 4.4, 2.3, 3.1, 5.6, 5.6, 1.8, 1.6, 1, 0.9, 0.5, 0.6, 
    0.5, 2.1, 2.6, 1.4, 0.5, 2.7, 2.5, 2.1, 2, 5.4, 3, 1.3, 1.2, 4.9, 1.2, 
    1.7, 2.4, 1.8, 3, 0.8, 1, 1, 1.6, 1.9, 1.1, 1.3, 0.8, 0.2, 0.3, 1.2, 1.3, 
    2, 0.9, 1.4, 1.1, 1.5, 1.6, 1.3, 0.9, 0.9, 0.5, 0.5, 1.5, 0.7, 1.3, 1.2, 
    1.6, 1.2, 1.3, 0.3, 0.6, 1, 1, 0.4, 1.1, 1.1, 1.2, 1, 0.8, 0.3, 0.4, 1.7, 
    0.7, 0.8, 0.9, 1.4, 0.8, 1.2, 0.3, 5.6, 8, 8.1, 7.9, 7.2, 6.7, 8.5, 8.8, 
    9.5, 9.1, 10, 9.1, 8.5, 6.5, 7.6, 8.8, 7.8, 5.2, 5.9, 6.1, 4.6, 5, 1, 
    1.1, 2, 2.5, 3.7, 0.8, 1.7, 0.9, 0.8, 1.7, 1.6, 1.9, 0.7, 8.5, 10.8, 8.2, 
    7, 7, 6.8, 9.5, 8.8, 11.6, 10.4, 8.1, 7.9, 5.9, 7.3, 7.3, 7.2, 7.1, 2.6, 
    4.5, 4.9, 3.6, 5.2, 4.4, 4.4, 5.1, 5.1, 5.7, 3.7, 5.3, 2.8, 4.2, 4.8, 
    4.5, 4.6, 4.1, 2.5, 0.6, 0.9, 0.8, 0.2, 1.6, 0.3, 0.2, 1.8, 0.6, 0.1, 
    0.6, 0.6, 0.4, 0.4, 0.6, 0.7, 0.4, 0.2, 0.6, 0.2, 0.5, 0.9, 0.6, 0.5, 
    0.6, 0.8, 0.8, 0.1, 0.9, 1, 0.1, 0.7, 0.4, 0.6, 1.4, 1.2, 0.8, 0.8, 0.8, 
    1.8, 0, 0.2, 0.4, 0.1, 1, 0.9, 3.2, 2.1, 1.1, 0.7, 0, 0.3, 0.4, 0.1, 0.3, 
    0, 0, 0, 0, 0, 0, 0, 0, 3.2, 3.3, 2.9, 2.6, 1.9, 1.4, 2.4, 7.2, 7.5, 3.8, 
    4.5, 4.9, 2, 3.4, 5.6, 5, 4.6, 3.6, 1.3, 1.1, 0.9, 0.9, 0.9, 0.3, 0.5, 
    0.3, 1.2, 2.7, 3.4, 3.5, 0.2, 0.9, 0.2, 1.2, 0.6, 0.5, 0.5, 0.3, 0.5, 
    0.1, 1.1, 0.4, 0.5, 0.3, 0.9, 0.7, 0.8, 0.1, 1, 0.1, 0.7, 0.5, 0.4, 0.3, 
    0.7, 1, 1.1, 0.4, 1.8, 3.2, 2.3, 0.6, 2.4, 0.3, 1.4, 3.2, 1.1, 0.6, 1.1, 
    1.2, 1.4, 1.2, 1.2, 1.2, 0.4, 1.1, 1, 1.6, 1.6, 1.1, 0.1, 0, 5.1, 4.3, 
    3.8, 0.8, 1.7, 1.4, 1.4, 1.7, 0.7, 5.4, 4.3, 5.6, 5.6, 1.8, 6.4, 5.9, 
    5.3, 5.3, 6.7, 4.9, 4.5, 3.2, 1.6, 1.8, 1.8, 0, 1.6, 1.1, 0.5, 0.6, 1.2, 
    1.4, 0.9, 1.6, 0.8, 1.6, 0.9, 0.6, 1, 0.1, 0.1, 0.9, 6.1, 4.3, 6.4, 6, 
    6.8, 7.1, 8.7, 8.3, 7.8, 8, 7.4, 7, 7.1, 8.7, 2, 3.7, 6.1, 6.2, 5.8, 5.7, 
    5.6, 5.1, 4.5, 5.7, 5.7, 5, 5, 4.4, 4.5, 0.2, 1.2, 0.9, 1.1, 0.2, 1.7, 1, 
    2.1, 2, 1.2, 0.1, 0.1, 0.1, 2.6, 0.5, 1, 1, 0.3, 0.2, 0.7, 0.3, 0.6, 0.5, 
    0.1, 1.5, 0.8, 1.1, 3.9, 3.3, 4.5, 4.9, 6.8, 4.9, 8.8, 4, 4.9, 5.7, 4.4, 
    6.3, 4.7, 4.1, 4.2, 4, 3, 1.3, 1.1, 1.5, 1.2, 3, 2.7, 2.4, 3.1, 1.7, 0.1, 
    0.3, 0, 0.8, 0.2, 0.4, 0.2, 0.8, 0.7, 0.2, 0.1, 0.1, 0.5, 0.7, 0.2, 0.3, 
    0.3, 0.7, 0.7, 0.5, 0.2, 0.6, 0.5, 0.9, 0.8, 0.6, 0.4, 1.1, 3.7, 3.8, 
    0.5, 2.8, 3.2, 4.6, 3.5, 7.4, 7.7, 6.1, 5.2, 3.8, 3, 1.8, 0.5, 2.5, 2.1, 
    7.8, 5.8, 5.2, 5.1, 5.6, 5, 5.3, 3.5, 4, 1, 1.8, 3.9, 1.8, 1.6, 2.1, 1.1, 
    1.8, 1.7, 0.8, 0.6, 0.9, 1, 1.1, 1.2, 1.8, 0.6, 1.3, 0.7, 1, 0.3, 0.4, 
    0.7, 0.4, 0.4, 0.4, 0.9, 0.5, 0.4, 0.9, 0.2, 0.8, 0.4, 1.4, 0.8, 0.8, 
    1.2, 1.3, 1.5, 1.9, 2, 1.2, 3.4, 7.6, 6.3, 4.9, 4.2, 2.1, 4.1, 4, 4.9, 
    3.4, 1.8, 0.8, 0.4, 1.3, 1.6, 2, 1.5, 1.1, 1.2, 0.7, 1.2, 2.7, 0.4, 0.8, 
    1.6, 1.2, 1.4, 1.4, 0.8, 1.5, 1.2, 1.2, 0.5, 0.5, 0.3, 0.1, 0.4, 0.6, 
    0.3, 0.5, 0.6, 0.1, 0.4, 0.4, 0.3, 0, 0.7, 0.1, 1, 1.2, 0.3, 0.6, 1.3, 
    0.5, 0.9, 1.1, 0.8, 0.5, 1, 0.4, 0.5, 0, 0.4, 0.5, 0.4, 4.7, 4.4, 5.9, 
    5.8, 5.1, 1.7, 3, 0.3, 0.9, 0.1, 1.2, 1.3, 1.5, 2.9, 2.5, 2.4, 1.5, 1.4, 
    0, 1, 1, 7.2, 5.2, 5, 6, 4.3, 4.6, 5.1, 4.1, 3.1, 4.4, 3.7, 3, 2.6, 2.6, 
    6.1, 3.5, 3.9, 3.3, 2.9, 2.3, 1.9, 3, 2.9, 1.7, 0.7, 0.4, 0.8, 0.3, 0.4, 
    2.8, 0, 0.3, 0.7, 0.3, 0.3, 0.3, 2, 1.4, 0.7, 1, 1, 0.9, 1.1, 2.3, 1.3, 
    1.5, 1.4, 0.9, 0.5, 1.7, 0.8, 1.1, 1.8, 0.1, 1.4, 1.5, 2.7, 2.3, 0.6, 
    0.3, 0, 0, 7.1, 9, 7.8, 7.1, 8.1, 8.8, 8.3, 7.9, 7, 6.8, 7.5, 9.5, 10.1, 
    8.1, 8.7, 11.2, 10.4, 11.7, 10.5, 9.3, 11.6, 4.7, 7.3, 9.7, 8.6, 7.6, 
    7.2, 7, 6, 5.4, 3.6, 6.3, 4.9, 4.9, 2.9, 1.6, 2, 1.7, 1.4, 0.9, 0.8, 1.5, 
    0.6, 0.9, 0.5, 0.5, 1.3, 1, 1.3, 0.6, 0.6, 0.6, 0.6, 0.2, 0.4, 1.7, 0.7, 
    1.4, 0.8, 0.6, 1, 1, 1.6, 2, 2.9, 1.5, 1, 3.3, 4.2, 3.2, 3.2, 2.3, 1.1, 
    2, 4, 2.8, 1.3, 1.1, 1.8, 1.3, 0.4, 0.8, 0, 0.5, 0.3, 0.4, 0.9, 0.6, 1.4, 
    0.4, 1.4, 5.6, 5.9, 6, 6.1, 8.6, 9.3, 7.4, 7.4, 7.6, 8.3, 8.8, 8.2, 9.6, 
    10.7, 9.6, 9.8, 9.8, 9.4, 8, 7.3, 8.4, 6.8, 4.5, 5.6, 7.7, 6.6, 5.7, 9.1, 
    4.7, 3.6, 10.5, 5, 8.8, 4.7, 4.7, 6.8, 4.7, 6, 2.9, 2.5, 3.2, 2, 3.7, 
    2.5, 1.2, 0.9, 1.6, 1.6, 1.3, 1.2, 0.7, 1.1, 1.4, 1.4, 1.9, 1.1, 1.6, 
    0.6, 0.5, 1.5, 1.4, 0.8, 0.9, 0.7, 0.8, 0.2, 0.7, 0.7, 0, 0.2, 0.4, 0.1, 
    0.6, 0.6, 0.4, 0.8, 1, 0.9, 1, 0.5, 1.2, 0.6, 0.1, 1.3, 0.1, 0.3, 1, 0.2, 
    0.7, 1.2, 0.1, 0.1, 0.6, 0.3, 0.2, 0.5, 0.6, 0.6, 0.8, 0.8, 0.3, 0.8, 
    0.2, 0.9, 1.4, 0.9, 1.6, 1, 0.8, 0.4, 2, 1.5, 0.8, 1, 1, 0.6, 0.6, 0.8, 
    1.3, 0.5, 0.1, 0.6, 0.6, 0.8, 0.1, 0.2, 1.2, 0.5, 0.1, 0.5, 0.6, 0.6, 
    1.3, 1.1, 1.1, 0.2, 0.4, 0.3, 0.3, 1.2, 1, 0.5, 0.3, 0.2, 0.8, 0.4, 1.4, 
    1, 0.6, 0.3, 1.2, 0.3, 0.7, 0.7, 0, 0.9, 0.6, 1.6, 1, 1.4, 0.9, 0.8, 1.9, 
    1, 0.8, 0.4, 1.4, 2, 1.7, 1.5, 0.9, 0.7, 0, 0.5, 0.4, 1.7, 1.7, 1.4, 1.4, 
    1.3, 0.6, 0.6, 0.8, 1.2, 1, 0.6, 0.4, 1.5, 0.8, 1.4, 1.7, 0.4, 0.5, 0.3, 
    1.3, 1.2, 0.6, 1.5, 0.5, 0.2, 0.6, 3.5, 0.4, 4.6, 1.2, 4.3, 1.8, 1.8, 
    0.7, 0.5, 0.7, 1.2, 2.2, 2.9, 4.8, 5.9, 6, 6, 5.3, 4.2, 5.5, 4.8, 5, 5.2, 
    5, 3.5, 2.2, 3.7, 1.1, 2.2, 1.7, 2.1, 1.6, 1.6, 0.6, 1.8, 2.5, 3.6, 0.7, 
    3, 3, 2.9, 3.9, 4.6, 2.7, 1.8, 1.5, 0.6, 0.5, 1.7, 4.2, 7.3, 7.5, 3.8, 
    2.5, 3.1, 1.9, 9.5, 8.8, 3.4, 7.7, 6.4, 5.8, 3.2, 4, 3.4, 2.7, 4.3, 5.5, 
    2.9, 3, 4.9, 4.5, 4.1, 4.7, 4.6, 4.7, 4.7, 4.4, 4.1, 4.3, 1.2, 2.4, 2.1, 
    1.7, 1.8, 2.9, 1.3, 2.2, 1.8, 2.5, 7, 0.6, 1.5, 7.5, 2.9, 4.1, 8.8, 3.3, 
    1.9, 8.4, 1.1, 3.7, 8.7, 2.3, 2.4, 10.5, 1.2, 1.7, 2.5, 6.5, 7.8, 7, 7.9, 
    7.7, 3.9, 6.8, 5.8, 6.1, 1.7, 2.1, 3.3, 4.6, 1.8, 4.3, 1.6, 0.9, 1.4, 
    1.3, 1.1, 0.7, 0.7, 3.3, 1.8, 1, 2.7, 1.3, 0.1, 0.1, 0.2, 2, 2, 1.5, 0.7, 
    2.2, 1.6, 1.8, 1, 1.7, 0.2, 1.1, 1.9, 0.9, 0.6, 1.1, 0.4, 0.6, 0.8, 0.5, 
    0.5, 0.6, 0.9, 0.3, 0.1, 3.1, 0.1, 0.8, 1.4, 0.1, 0, 0.7, 0.9, 0.2, 0.3, 
    0.7, 1.4, 1.3, 0.8, 1.4, 1.2, 0.2, 0.5, 0.6, 0.4, 0.7, 0.6, 1.4, 1.2, 
    1.8, 0.8, 2.6, 1.2, 0.8, 0.2, 0.7, 1.8, 1.4, 2.1, 2.3, 2.4, 1, 1.5, 2.5, 
    1.1, 1.6, 0.6, 0.9, 0.4, 0.2, 0.6, 1.1, 0.7, 1.5, 1.1, 0.5, 0.8, 0.6, 
    0.8, 1.4, 0.6, 1, 1, 0.9, 1.1, 0.5, 1.2, 1.3, 1, 1, 1.5, 0.8, 0.7, 0.1, 
    0.9, 1.1, 0.3, 1.2, 0.8, 1.4, 0.5, 0.6, 0.4, 0.5, 0.5, 1, 0.5, 1.4, 1.3, 
    0.3, 0.8, 0.5, 0.5, 0.6, 0.8, 2.4, 0.9, 0.6, 3.1, 2.5, 0.5, 1.4, 0.6, 
    1.4, 0.3, 1.2, 0.2, 0.4, 0.1, 0.3, 0.5, 1.8, 0.5, 0.8, 1.3, 0.5, 1.3, 
    0.7, 1, 0.3, 0.4, 0.8, 1.2, 0.9, 0.8, 1.6, 0.9, 0.2, 0.8, 2.8, 0.6, 1.3, 
    5.4, 9.4, 7.6, 8.9, 9.6, 8.9, 9.5, 9.6, 10, 6.7, 2.2, 3.9, 2.9, 1.1, 1, 
    0.8, 0.8, 0.9, 1.1, 1.4, 1.9, 1.7, 1.4, 0.8, 1.5, 1.5, 5.7, 5.5, 4.1, 1, 
    2.2, 4.1, 1.6, 4.2, 7.9, 8.5, 7.7, 5.4, 6.4, 5.7, 4.4, 3.8, 3.7, 3.3, 
    2.4, 1.4, 0.6, 1, 0.3, 1.1, 1.3, 0.4, 1.3, 1.1, 3.7, 1.1, 2.4, 2.4, 4.3, 
    0.6, 1.4, 1.4, 0.4, 0.7, 10.3, 7.1, 7.1, 4.9, 7.6, 9.3, 7.3, 9.2, 8.7, 
    9.3, 9.2, 9.2, 5.9, 7.4, 4.1, 5.4, 2.7, 3.8, 4.2, 6.4, 5.3, 7, 6.3, 4.5, 
    5, 4.7, 7.1, 3.3, 3.9, 4.2, 7, 5.2, 4, 2.2, 3.8, 5.9, 0.4, 1.1, 0.5, 0.8, 
    0.7, 0.2, 0.9, 0.7, 0.6, 1.7, 1, 1.3, 1.5, 1.2, 1.1, 3, 1.4, 0.9, 1, 1.4, 
    0.7, 0.5, 1.3, 0.7, 1.1, 0.2, 1, 0.3, 0.9, 0.7, 0.4, 0.3, 0.5, 0.6, 0.9, 
    1, 0.8, 1.2, 1.2, 0.9, 0.6, 0.6, 1.2, 1.1, 1, 0.8, 0.7, 1.4, 0.4, 1.2, 
    0.8, 0.8, 0.5, 0.9, 1, 0.5, 0.7, 0.6, 0.3, 1.1, 0.5, 0.2, 1.8, 0.9, 0.5, 
    0.1, 0.2, 0.9, 1, 1.4, 0.4, 0.6, 1, 1, 0.4, 1, 0.5, 1.2, 0.8, 1.2, 1.2, 
    1.3, 0, 0.1, 0.5, 0.8, 1.7, 1.1, 0.8, 0.2, 0.7, 0.7, 0.7, 1.4, 0.4, 0.9, 
    0.5, 0.5, 0.8, 0.2, 0.4, 0.5, 0.5, 0.4, 1.1, 1.1, 0.9, 1, 0.4, 0.4, 0.3, 
    0.8, 1.5, 1.2, 0.3, 0.1, 1.4, 1.1, 6.5, 7.6, 4.7, 5.7, 5.4, 3.7, 7.2, 7, 
    7.8, 6.1, 7.4, 6.5, 7, 6.9, 7, 5.3, 8, 7.5, 6.9, 6.9, 7.2, 5.3, 6.1, 6.5, 
    7.2, 5.9, 5.3, 5.2, 5.8, 4, 1.2, 1, 1.1, 2.5, 0.1, 0.7, 1.9, 1, 0.7, 0.7, 
    0, 1.2, 4.1, 1.4, 2.2, 3.3, 2.1, 2.6, 2.7, 2.6, 1.2, 1.3, 0.7, 0.4, 0.3, 
    0.8, 0.4, 0.3, 0.8, 1.5, 0.1, 1.6, 1, 1.9, 1.3, 1.3, 1.4, 0.9, 0.4, 2.2, 
    1.4, 0.4, 1.6, 0.9, 1.3, 0.6, 0.9, 1, 1.1, 1, 1.4, 0.3, 0.5, 1, 0.9, 0.7, 
    0.5, 1.3, 1.6, 1.4, 0.8, 0.2, 0.9, 1, 1, 0.2, 0.5, 0.4, 1.5, 1.9, 0.5, 
    0.9, 3.9, 6.5, 7.9, 7.4, 6.3, 7.1, 7.9, 7.2, 6.4, 9.7, 9, 8.2, 7.7, 9.4, 
    8.2, 9.6, 10.1, 9.9, 11.2, 11.9, 13.3, 11.9, 9.6, 10.2, 11.4, 11.5, 12.6, 
    11.1, 10.7, 10.9, 10.4, 10.8, 9.5, 8, 10.2, 8, 9.8, 7.9, 9.7, 9.7, 7.6, 
    11, 9.5, 10.2, 10.9, 8.3, 7.7, 7.5, 8.6, 12.1, 10.8, 11.6, 11.2, 7.1, 
    6.3, 7.7, 7.3, 5.3, 2, 0.9, 2, 1.9, 1.6, 1.8, 1.1, 0.3, 0.6, 0, 0.8, 0.1, 
    0, 0.7, 0.7, 0.9, 1.2, 0.5, 0.7, 0.8, 0.9, 0.8, 0.6, 0.1, 0.4, 1.4, 2, 2, 
    1.4, 1.3, 1.5, 1.8, 2, 2.5, 2.8, 2.5, 2.6, 2.1, 2.3, 2.7, 3.2, 2.9, 3.1, 
    3.2, 3.4, 3.4, 3.6, 3.5, 2.5, 2.8, 2.9, 2.9, 2.8, 3.3, 4.9, 4.1, 4.9, 
    6.7, 5.9, 5.3, 4.7, 4.1, 3.2, 3, 2.7, 2.8, 2.9, 2.9, 3.7, 4, 4.1, 5, 6, 
    5.9, 7.7, 7.4, 6.8, 6.2, 6.1, 6.6, 6.6, 6.3, 5.1, 5, 4.4, 3.3, 2.9, 2.7, 
    2.9, 3.7, 4.2, 3.8, 3.5, 4, 4.1, 4.1, 4.6, 4.9, 4.4, 5.4, 5.2, 4.7, 4.5, 
    5.1, 6, 7.3, 7.8, 7.4, 8.1, 7.3, 9, 9.5, 8.9, 7.8, 8, 7.1, 6.7, 6.1, 4.9, 
    4.5, 3.9, 4.3, 3.5, 2.6, 1.5, 2, 5.7, 8.1, 7.4, 7.3, 7, 6.8, 6.4, 4.5, 
    3.9, 2.5, 2.8, 2.8, 2.3, 2.5, 2, 2, 2.2, 2.6, 3, 3, 3.5, 4, 4.1, 4.1, 
    4.4, 5.2, 4.9, 5.2, 5.6, 5.8, 5.7, 5.9, 5.9, 5.1, 4.2, 3.9, 4, 4, 4, 4.1, 
    4, 3.7, 4.1, 3, 3, 3.2, 3.7, 4.1, 3.8, 3.5, 3.3, 3.9, 4.8, 5.4, 5.6, 5.5, 
    5.3, 5.2, 5.2, 5.3, 5.3, 5.3, 5.6, 6, 6.2, 6.2, 5.7, 5.8, 5.8, 5.6, 5.6, 
    5.4, 5.2, 5.1, 5, 4.8, 4.5, 4, 4.1, 3.9, 3.5, 2.9, 2.1, 1.5, 0.9, 1.6, 
    0.6, 1.4, 1.8, 0.8, 1, 2.2, 2.6, 3.2, 3.2, 4.5, 5.1, 6.4, 8.8, 9.7, 9.7, 
    11.1, 11.1, 11.4, 10.2, 7.8, 6.4, 4.4, 2.6, 2.7, 2.9, 2.4, 1.3, 1, 2.6, 
    2.1, 2.1, 2.7, 2.8, 3, 3.2, 2.5, 2.8, 2.6, 3, 2.6, 1.8, 1.6, 1.4, 1.9, 
    2.8, 2.7, 2.6, 2.7, 3.3, 3.6, 3, 3.1, 2.7, 2.2, 1.5, 1.9, 1.6, 2.6, 3.2, 
    2.9, 2.4, 2.7, 3.1, 0.5, 1.3, 0.6, 1.3, 1.6, 2, 3.4, 1.1, 0.1, 2.3, 6.8, 
    8.7, 12.8, 11.8, 16, 14.5, 14.7, 14.9, 14.5, 12.7, 12.1, 7.3, 5.6, 2.5, 
    4.2, 11.6, 11.8, 9, 11, 8.8, 10.7, 9.1, 8.4, 5.7, 7.5, 9.5, 8.6, 5.3, 
    7.8, 7.7, 7.6, 7.4, 7.3, 6.9, 6.4, 6.5, 6.2, 5.5, 4.7, 5.1, 4.2, 3.3, 3, 
    2.1, 1.7, 2.1, 2.6, 2.9, 3.1, 3.4, 3.8, 3.8, 3.7, 3.5, 3.2, 2.9, 2.5, 
    2.2, 2, 1.1, 0.4, 1.3, 0.9, 0.9, 0.4, 1.3, 0.2, 0.6, 1.1, 2.7, 0.7, 0.5, 
    0.4, 0.5, 1.3, 0.5, 0.1, 0.7, 1.7, 0.1, 0.1, 0.7, 1, 0.9, 3.1, 0.4, 1.1, 
    5.4, 4, 4.6, 5.4, 3.8, 3.3, 3.7, 5.8, 7.9, 10.3, 4.7, 4.8, 6.3, 3.3, 9.2, 
    8.7, 6.4, 7.1, 4.1, 2.6, 3.9, 2.1, 1.6, 3.4, 1.8, 6.5, 3, 3.3, 0.8, 3.7, 
    4.7, 7.4, 1.4, 4.2, 2.1, 2.9, 4.2, 4.6, 2.9, 1, 1.6, 1, 0.7, 2.2, 0.6, 
    0.4, 0.1, 0.8, 0.8, 1.1, 1.3, 0.5, 0.2, 2.6, 2.5, 0.6, 0.1, 1.1, 1.1, 
    1.7, 1.1, 0.5, 0.4, 0.4, 0.5, 0.8, 1.7, 0.5, 0.7, 1.4, 0.5, 0.6, 0.9, 
    0.4, 1.8, 1.9, 1, 1.6, 1.3, 1.3, 1.7, 1.5, 2.1, 1.4, 0.5, 2, 2.2, 1.7, 
    1.3, 1.2, 1.2, 0.5, 0.6, 0.1, 1.1, 0.9, 2.1, 3.5, 0.4, 2.3, 4.5, 4, 2.7, 
    1.9, 2.7, 0.9, 0.9, 0.7, 1.2, 1.2, 0.4, 1.7, 0.9, 1.1, 0.4, 0.4, 1.1, 
    0.6, 0.9, 0.9, 0.7, 3.5, 1, 0.4, 1.1, 3.4, 0.3, 0.5, 1, 0.5, 0.3, 0.7, 
    0.7, 1.1, 1, 0.5, 0.1, 0.2, 0.3, 0.8, 0.7, 0.9, 0.5, 0.8, 0.5, 0.3, 0.2, 
    0.9, 0.3, 1.3, 0.5, 0.5, 1.4, 0.5, 1.7, 0.1, 0.6, 1.1, 0.9, 0.2, 0.5, 
    0.5, 0.9, 0.2, 0.6, 0.9, 0.8, 0.7, 0.3, 0.9, 0.6, 3.6, 0.9, 0.8, 0.8, 
    2.1, 3.1, 2.7, 1.2, 0.3, 1.1, 0.3, 6.2, 8.8, 10.3, 11.2, 9.7, 10.8, 11, 
    8.7, 7.5, 7.6, 9.2, 7.6, 5.7, 5.9, 4.7, 5.4, 3, 1.4, 2.5, 1.4, 1.3, 2.2, 
    0.8, 1, 2.8, 2.4, 3.5, 0.6, 0.3, 1.5, 1.6, 1.9, 1.9, 0.6, 0.6, 0.1, 0, 
    0.1, 2, 1.1, 1.3, 1, 0.3, 0, 0, 0, 0.2, 2.2, 1.1, 0.8, 1, 5, 4.1, 3, 2.1, 
    0.9, 1.1, 1.1, 1.2, 0.5, 1.4, 1, 0.6, 0.7, 0.8, 0.7, 1, 0.7, 0.4, 1.4, 
    1.8, 2.6, 3.2, 3.6, 4.4, 4.7, 5, 3.8, 5.3, 4.7, 2.9, 4.4, 4.7, 5.7, 6.1, 
    6.1, 6.3, 8.3, 9.6, 8.5, 9.4, 9.5, 8.6, 8.5, 7.5, 7.4, 7.7, 8.9, 6.4, 
    8.9, 5.7, 5.8, 5.9, 3, 6.4, 5.1, 3.9, 12.6, 11.2, 9.8, 7.5, 7.7, 6.6, 
    6.7, 6.5, 4.5, 4.8, 5.4, 2.2, 5.7, 5.5, 4.7, 0.7, 0.3, 4, 4.9, 4.9, 4.3, 
    5.4, 4.6, 4.2, 4.3, 3.3, 6.1, 5, 3.9, 4.7, 4.6, 9.2, 9.8, 10.6, 9.8, 9.8, 
    7.8, 8.4, 9.5, 9.9, 10.8, 11.7, 12.7, 14.6, 13.4, 11.7, 10.7, 8.4, 11.9, 
    7.7, 7.3, 9.1, 9.2, 6.4, 10.5, 11.3, 8, 9, 11.5, 9.7, 9.5, 10.4, 9.9, 
    9.7, 8.8, 8.6, 11.3, 11, 4.7, 6.5, 5.2, 8.1, 7.4, 3.7, 5, 1.8, 1.8, 2.3, 
    6.5, 6.2, 0.5, 1.4, 1.7, 1.3, 0.4, 1.3, 1.6, 0.5, 0.9, 1, 0.3, 0.5, 0.9, 
    0.5, 0.7, 0.1, 0.5, 0.4, 1.3, 1, 1.2, 0.6, 0.2, 1.7, 1.6, 1.9, 0.5, 2.1, 
    0.4, 0.9, 1.5, 0.4, 1.1, 0.9, 0.9, 0.9, 0.2, 0.8, 0.7, 2.5, 1.3, 0.3, 
    2.1, 0.4, 1, 1.3, 0.6, 0.8, 0.7, 0.7, 3.6, 2.4, 2, 2.2, 3.8, 7.4, 6.9, 
    6.2, 8.7, 7, 8.3, 6.4, 7.2, 7.3, 7.1, 6.4, 4.8, 5.3, 5.2, 2.7, 5.5, 6.9, 
    6.2, 5.2, 6.1, 5.3, 4.7, 3.4, 2.4, 2.9, 3.5, 3.1, 0.6, 1.5, 0.9, 0.8, 
    0.8, 1.5, 0.8, 1.1, 2.3, 1.1, 0.6, 0.9, 1, 0.9, 0.9, 1.7, 1.2, 2.3, 3, 
    3.5, 1.8, 0.7, 0, 0.5, 0.3, 0.9, 0.4, 0.9, 0.9, 3.1, 1, 0.9, 2.8, 0.1, 
    0.8, 1.4, 0.7, 0.1, 1.3, 0.1, 0.7, 0.3, 0.9, 0.4, 0.6, 0.6, 0.7, 1, 0.7, 
    0.4, 0.5, 0.7, 0.3, 0.8, 2, 1.8, 0.2, 1, 0.9, 0.4, 0.1, 2.1, 0.9, 0.7, 
    1.3, 0.7, 0.2, 0.4, 1.2, 1, 2, 0.4, 0.5, 1.3, 3.6, 1.7, 1.7, 1.2, 1.4, 
    1.1, 2.7, 2.2, 2.5, 5.7, 1.6, 3.3, 3.2, 2.1, 2.6, 2, 3.7, 6.4, 2.7, 2.4, 
    4.4, 4.1, 4.1, 4.3, 4, 3, 1.1, 0.2, 1, 0.3, 0.6, 0.7, 0.3, 0.7, 0.6, 0.7, 
    0.2, 0.9, 0.5, 0, 0.7, 0, 1.5, 1.4, 0.2, 0.2, 0.8, 0.8, 0.8, 1.5, 1, 1, 
    0.5, 0.1, 0.8, 0.8, 1, 0.2, 0.6, 1.1, 0.2, 0.9, 0.6, 0.2, 5.1, 3.4, 3.2, 
    1, 2, 2.4, 4.6, 3.6, 3.4, 0.7, 5.8, 5.2, 4.6, 5.5, 5.5, 6, 5.3, 3.7, 0.6, 
    6.6, 6, 3.9, 6.5, 5, 4.7, 4.2, 0.3, 1.8, 1.7, 1.7, 4.4, 4.8, 5.5, 5.3, 
    3.6, 3.4, 4.5, 6.2, 4.7, 4.3, 3.9, 3, 0.7, 0.4, 1.3, 0.6, 3, 1.9, 1.1, 
    0.6, 0.7, 0.5, 0.6, 0.7, 0.3, 0.5, 3.6, 4.3, 6.2, 5.8, 5.4, 1, 2, 0.9, 
    1.6, 1.6, 1, 1, 0.8, 1, 1.6, 4.1, 4.1, 6.7, 4.8, 4.1, 4.8, 5.2, 6.1, 5.7, 
    8.1, 5.3, 4.6, 2.7, 5, 3.3, 2.2, 3.6, 4.2, 4.4, 2.7, 3.8, 2.6, 1.2, 1.5, 
    0.9, 2, 3, 2.6, 1.6, 0.5, 2.3, 0.8, 0.5, 1.2, 0.2, 2.6, 0, 0, 0.9, 0, 0, 
    0.3, 0.9, 1.7, 2.2, 1.4, 2.2, 4.6, 4.4, 3.2, 1.9, 0.5, 0.3, 0.9, 1.3, 1, 
    0.7, 3.8, 2.3, 1.6, 2.6, 4.2, 2.6, 1.6, 0.8, 1.1, 1.1, 0.7, 1.5, 1.5, 
    0.5, 1.3, 0.7, 2.1, 0.2, 1.1, 0.8, 0.3, 1.2, 0.3, 0.7, 0.8, 1.3, 0.8, 
    0.1, 1.4, 1.4, 0.7, 0.9, 1.4, 1.6, 0.3, 1.3, 0.5, 0, 0.7, 0.4, 0.5, 0.7, 
    0.6, 0.3, 1.8, 1.8, 2.3, 1.5, 1.6, 1.8, 0.5, 0.2, 1, 1.3, 0.4, 1, 0.9, 
    0.4, 0.5, 6.4, 6.6, 4.4, 7, 5.9, 5.1, 7.9, 6.7, 8.6, 9.4, 10, 10.4, 10.2, 
    11.3, 12, 10.6, 10.8, 9.2, 10.3, 8.8, 10, 7, 3.9, 2, 3.7, 2, 3.2, 0.8, 
    0.9, 0.5, 0.7, 1.9, 0.9, 0.6, 1.7, 3.4, 1.4, 0.8, 0.5, 0.5, 0.1, 6, 4.9, 
    4, 2.9, 2.5, 1.8, 1, 1.5, 1, 2.9, 3.2, 1.5, 2.9, 1.6, 1.9, 1.6, 2.6, 2.1, 
    6.3, 10, 7.9, 3.2, 4.9, 1.6, 1.7, 1.8, 0.8, 2.5, 2.4, 2.8, 2.6, 1.7, 5, 
    5.2, 2.9, 2.7, 5.2, 1.5, 3.3, 2.3, 2.6, 1.6, 10.1, 8.3, 8.9, 8.4, 4.8, 
    7.8, 5.9, 2.4, 2.4, 4, 4.2, 4.8, 3.1, 1.6, 2.3, 1.9, 4.4, 5.2, 5.4, 4.4, 
    4.6, 5, 6.5, 5.1, 2.5, 1.5, 8.9, 7.7, 2.5, 1.8, 1.9, 1.3, 1, 1.1, 4.1, 
    1.9, 2.8, 2.9, 1, 1.3, 1.9, 1.9, 1.5, 2.4, 1.2, 0.9, 0.6, 0.5, 0.6, 1, 
    0.5, 1.4, 2.1, 2.1, 1.7, 2, 2, 0.4, 0.8, 0.2, 0.6, 0.4, 0.9, 0, 0, 0.3, 
    0.6, 1.4, 0.3, 0.5, 2.1, 1.8, 1.5, 2.4, 1.7, 0.2, 0.2, 0.4, 0.7, 0.1, 0, 
    1.8, 1.1, 0.4, 0.8, 1.8, 2.3, 0.3, 0.6, 0.7, 1.8, 1.5, 1.4, 0.9, 0, 1.2, 
    0.5, 0.1, 0.6, 0.6, 0.3, 1, 0.7, 0.5, 0.2, 0.1, 0.9, 0.6, 1.5, 0.9, 0.4, 
    0.2, 4, 2.5, 2.1, 1.2, 2.2, 1.6, 0.8, 1.5, 0.9, 0.6, 0.1, 0.8, 0.4, 0.4, 
    0.8, 1.4, 0.5, 1.5, 0.4, 0.6, 0.2, 0, 0.7, 0, 0, 1.8, 1.2, 1.4, 1.2, 1.4, 
    0.1, 1.9, 2.1, 0.5, 1, 1.1, 0.8, 0, 0.8, 0.7, 0.5, 0.3, 0.8, 0.3, 0.1, 
    0.2, 1.2, 0.1, 1.5, 1.5, 0.1, 1.3, 0.5, 0.8, 2.4, 5.4, 5.9, 4.2, 4.3, 4, 
    3.6, 4.1, 4.9, 2.5, 1.6, 2.1, 4.2, 3.2, 2.1, 2.3, 1.6, 0.8, 1.8, 1.9, 
    2.9, 3.1, 2.6, 2.2, 0.9, 1.2, 1.4, 1.6, 1.2, 1.7, 1.6, 2.5, 3.6, 4.3, 
    2.7, 2.8, 3.8, 1.8, 5.1, 5.4, 5.5, 6.2, 4.2, 3.9, 3.8, 2.4, 1.1, 1.7, 
    1.8, 1.2, 2, 1.2, 0.4, 1.1, 0.5, 1, 0.9, 5.7, 3.6, 4.2, 4.2, 2.5, 0.3, 
    1.4, 0.2, 0.4, 2.5, 2.7, 1.5, 1.7, 3.7, 3.2, 3.7, 3.2, 2.5, 2.6, 3, 3.5, 
    4.2, 3.8, 4.1, 4.3, 3.6, 3.6, 2.9, 2.7, 1.3, 0.4, 2.2, 2.4, 2, 1.2, 0.7, 
    1.7, 1.2, 1.6, 1, 0.4, 0.6, 0.2, 0.4, 0.3, 0.4, 0.7, 0.6, 0.6, 0.4, 0.4, 
    0.1, 1.7, 2.7, 1.5, 3.3, 3.1, 3.9, 2.5, 3, 2, 2, 1.8, 3.1, 2.6, 3.3, 2.4, 
    2, 2.5, 2, 0.6, 2.2, 2.8, 3, 2, 1, 1.6, 1.5, 0.5, 2.6, 2.4, 2.7, 3.4, 
    3.1, 0.3, 0.5, 0.3, 0.2, 0, 1.4, 0.7, 1.5, 1.7, 1.6, 1.4, 1.3, 1.3, 1.4, 
    1.5, 1.4, 2.5, 1.8, 2.6, 2.4, 2.6, 2.2, 3, 2.5, 2.2, 2.5, 1.4, 1.5, 1.7, 
    1.7, 0.6, 0.7, 1.2, 0.6, 0.3, 0.4, 0.2, 1.6, 0.8, 0.1, 1.4, 1.3, 0.5, 
    0.9, 1.7, 2.1, 1.6, 1.1, 1, 0.9, 0.9, 0.2, 0, 1.5, 1, 0, 0.2, 0.2, 0.2, 
    0.3, 0.3, 0.1, 0, 0.5, 1.4, 1.9, 3.9, 4.5, 5.6, 4.8, 3.8, 2.1, 1.5, 0.6, 
    0.7, 0.5, 1, 1.4, 2.1, 1.1, 5.3, 3.9, 4.1, 4.9, 5.6, 4.5, 3.5, 4.5, 5, 
    2.8, 4.1, 4.2, 2.9, 3.5, 2.7, 1.1, 1.1, 0.8, 0.4, 1.3, 1.3, 0.9, 0.4, 
    0.7, 0, 0.1, 1.1, 1.8, 1.9, 2.4, 0.7, 2.1, 1.1, 2.2, 1.3, 1, 1.6, 2, 1.3, 
    1.1, 1.4, 0.9, 1.6, 1.5, 1.4, 2, 1.7, 0, 0.2, 0.8, 1.4, 1, 0.9, 0.4, 0, 
    0, 0, 0.1, 1.8, 2.5, 2.2, 1.6, 0.2, 0.2, 0.8, 0.6, 0.3, 2.1, 1.5, 0.8, 
    0.8, 0.4, 0.1, 0.3, 2.4, 0.7, 0.5, 0.7, 0.2, 1, 0.1, 0.9, 0.3, 0.5, 0.4, 
    0.1, 0.9, 0.8, 2.2, 1.6, 0.5, 0.9, 1, 0.7, 0.4, 0.8, 1.2, 0.4, 0.2, 0.9, 
    0.2, 0.2, 0.6, 0.3, 0.5, 0.3, 0.4, 0.5, 0.3, 1.1, 1.3, 1.7, 1.3, 1, 1.9, 
    2.6, 1.5, 2.1, 1.9, 4.9, 1.6, 5.1, 4.2, 5.3, 8.1, 7.9, 5.3, 6.5, 3.2, 9, 
    2.8, 5.2, 6.4, 7.6, 9.6, 6, 4.8, 4.2, 2.6, 1.2, 2.3, 2, 4.7, 1.7, 2, 2.1, 
    1, 0.9, 1.4, 2, 1.1, 1.9, 0.6, 0.6, 1, 0.5, 1.1, 0.7, 0.6, 0.1, 0.4, 0.6, 
    1.2, 0.4, 1.2, 1.1, 1.2, 0.1, 1.2, 0.5, 0.4, 0.3, 0, 0, 0.2, 1, 0.7, 0.8, 
    2.1, 1, 1.5, 1.7, 1.1, 1.3, 0.6, 0.4, 0.8, 1.5, 2, 0.1, 0.7, 0.5, 2.1, 
    1.7, 2.1, 1.9, 1.2, 1.1, 0.5, 1.6, 1.4, 1.1, 0.4, 1, 0, 1.7, 0, 0.5, 0.3, 
    0.5, 0.2, 0.4, 0.2, 1.6, 0.5, 0.2, 0, 1.7, 3.3, 2.3, 2.2, 1, 1.5, 1.8, 2, 
    1.1, 1.2, 0.7, 2.2, 1.1, 1.4, 2.6, 2.9, 2.6, 0.5, 1.1, 0.5, 1, 1.1, 0.4, 
    1.2, 1.4, 1.5, 1.3, 1.3, 0.4, 0.7, 1.2, 0.1, 0.2, 0.6, 2.1, 0.4, 0.6, 
    0.1, 0.9, 0.7, 0.5, 0.7, 1.3, 0.3, 1.3, 0.5, 3.1, 4.3, 3.1, 4.6, 3.4, 
    3.3, 2.3, 3.7, 2.4, 2.2, 3.3, 4.3, 3.1, 3.4, 3.7, 4.9, 2.5, 1.6, 0.3, 
    0.2, 0.5, 0.2, 0.4, 2, 1, 0.6, 0.9, 1.5, 0.5, 0.5, 0.2, 0.7, 1.5, 1.2, 
    0.7, 1.1, 2.2, 2.3, 2.6, 0.1, 0.6, 0.9, 0.7, 1.1, 0.4, 0.6, 2.9, 0.2, 
    1.8, 1.8, 1.4, 1.7, 4, 0.4, 2.9, 2.7, 1.6, 2.6, 2.5, 2.2, 0.5, 2.3, 2.4, 
    2.5, 2.2, 0.6, 0.3, 2.8, 0.4, 3, 3, 3.3, 3.7, 2.9, 3.2, 1.3, 1.6, 1.8, 
    5.6, 4.7, 1.2, 1.7, 3.2, 2.1, 4.1, 3.9, 1.3, 2.3, 7.9, 2.4, 2.3, 4.1, 
    1.9, 2.7, 6.7, 6.9, 6.8, 3.2, 4.2, 3.6, 3.2, 2.4, 3.8, 2.9, 4.1, 4.6, 
    4.7, 7.6, 7.3, 5.9, 5.8, 2.8, 3.7, 5.6, 1.9, 4.3, 5.3, 5.6, 2.6, 2.6, 
    1.5, 4.7, 5.7, 3.5, 3.9, 2.1, 3.6, 2.2, 7.7, 2.1, 5.4, 3.3, 3.5, 5.6, 3, 
    5.9, 5, 1.7, 3, 3.5, 5.3, 3.5, 3.8, 4, 5.5, 4.7, 3.9, 6.8, 7, 6.4, 4.3, 
    4.9, 5.7, 1.6, 5.4, 3.7, 10, 10.4, 5.8, 1.6, 5.8, 4.3, 2.1, 6.7, 0.8, 
    1.6, 4.8, 2.8, 4.5, 5.4, 4.8, 4.7, 3.1, 4, 4.5, 5.5, 5, 3.9, 6.9, 3, 5.7, 
    4.6, 2.3, 2.4, 2.5, 4.6, 2.6, 3.2, 2.8, 4.7, 1.5, 2.8, 4.7, 3.4, 2, 0.9, 
    1.9, 2.3, 2.8, 2.6, 2.1, 0.9, 0.8, 1.4, 1.4, 0.8, 2.1, 2.1, 1, 0.1, 0.4, 
    2.2, 0.1, 0.2, 0.7, 0.7, 1.4, 3.7, 3.5, 2.1, 2, 1.3, 2.4, 1.4, 2.1, 1.9, 
    2.3, 2.5, 2.7, 2.4, 2.6, 2.3, 3.1, 1.3, 1.2, 2.9, 2, 2.3, 3.3, 2.3, 1.8, 
    1.1, 0.9, 0.8, 1.2, 0.6, 0.9, 0.9, 3.5, 2.3, 1.9, 2.4, 2.1, 0.9, 1.3, 
    1.6, 0.6, 0.8, 0.6, 0.9, 1, 0.6, 3.2, 4.7, 5.5, 4.9, 3, 2.6, 5.8, 4.4, 3, 
    4.6, 3, 2.4, 3.7, 3.9, 3.1, 2.9, 3.3, 2, 3.3, 4.7, 4.6, 4.4, 4.6, 2.3, 
    5.1, 5.2, 4.4, 4.4, 3.4, 4.9, 3.8, 1.9, 2.4, 1.9, 1.8, 3.1, 2.5, 2, 2.5, 
    3.9, 2.4, 2.1, 3.5, 3.7, 4, 2.6, 1.7, 2.5, 6.4, 5.3, 3.4, 2.9, 4.8, 4.8, 
    5.8, 3.5, 2.6, 10.3, 3.2, 8.4, 5.2, 3.3, 3.8, 3.4, 4, 10.2, 10.9, 11.1, 
    11.8, 5.8, 7.4, 12.6, 9.4, 1.9, 5.1, 7.6, 10.9, 7, 8.3, 6.6, 5.2, 2.8, 
    4.8, 3.3, 2.7, 3.2, 3.5, 8.2, 7.6, 3.5, 5.7, 3.7, 5.6, 3.7, 3, 6, 5.3, 
    5.3, 7.1, 5, 3, 3.6, 3.3, 3.1, 6.6, 3.3, 4.5, 5.3, 4.3, 2.9, 4.3, 4.5, 
    3.9, 5.2, 5.3, 2.4, 3.6, 5.1, 5, 5.6, 4.5, 4.6, 4.6, 5.2, 6.6, 6.4, 5.9, 
    6.1, 7.1, 7.5, 7.2, 6.5, 7.5, 6.4, 6.3, 5, 5.2, 6.1, 3, 2.4, 7.1, 6.4, 
    6.1, 7, 4.5, 6.5, 6, 5.4, 4.9, 4, 0.5, 1.6, 2.1, 1.1, 2.3, 1.1, 2.3, 0.6, 
    1.5, 2.3, 2.2, 0.2, 1.2, 0.9, 0.8, 0.7, 0.7, 0.6, 0.2, 0.8, 0.8, 0.3, 
    1.5, 1.1, 1.2, 1.2, 0.9, 1, 0.9, 1.1, 1.6, 2.6, 3.6, 3.8, 1.4, 1, 0.2, 
    0.4, 0.7, 1.1, 1, 0.3, 1, 1.6, 1.1, 1.3, 1.1, 1.1, 1.3, 1.7, 1.4, 1.3, 
    1.3, 1.9, 1, 3.3, 1.5, 1.8, 1.7, 2.1, 3.3, 0.6, 0.2, 0.1, 0, 0.4, 0.3, 
    0.3, 1.2, 2.6, 1.4, 2.3, 1.8, 2.9, 1.9, 1, 1.5, 0.9, 1.6, 1.8, 1.2, 1, 
    0.9, 0.7, 0.9, 0.5, 0.3, 1, 0.7, 0.8, 0.6, 1, 0.8, 1.6, 1.7, 1.2, 1.5, 
    1.2, 0.7, 1.6, 2, 1.3, 2, 2.3, 1, 1.7, 1.7, 0.8, 0.4, 0.4, 0.5, 1.3, 0.9, 
    1.1, 0.5, 1, 1.4, 1, 1.6, 1.9, 2.1, 2.1, 2, 1.1, 1.3, 1.1, 1.7, 1.8, 2.1, 
    2.6, 2.7, 2.9, 2.9, 2.7, 2.4, 0.6, 2.7, 3, 3.7, 3.1, 2.5, 3.3, 2.8, 2.6, 
    2.9, 2.7, 2.2, 2.4, 2.3, 2.1, 1.8, 2.6, 2.7, 2.6, 3.8, 3.3, 0.6, 1, 1.3, 
    0.7, 1, 1.3, 1.6, 2.9, 2.9, 2.3, 3, 3.4, 2.9, 2.8, 2.5, 2.3, 2.2, 2.3, 
    1.8, 2.4, 1.4, 2.5, 2, 1.8, 1.6, 1.5, 1.1, 2.7, 0.8, 0.9, 0.4, 1.8, 2.6, 
    1.7, 1.4, 1.1, 1.6, 2.4, 1.1, 0.3, 4.2, 1.4, 3.1, 2.9, 3.2, 2.7, 3.8, 
    4.3, 4, 3.9, 2.8, 3.1, 3.4, 2.2, 2.8, 1.3, 1.3, 2.1, 2.3, 4.6, 3.1, 3.8, 
    2.4, 1.9, 1.6, 3.2, 1.2, 1.6, 1.5, 1.4, 2, 1.2, 0.6, 1.3, 1.9, 1.9, 1.1, 
    0.3, 0.9, 1.4, 1.6, 1.5, 2.4, 1.7, 2, 2.8, 2.6, 2.4, 2.9, 3.4, 3.1, 3, 
    3.2, 1.4, 2.7, 1.6, 0.8, 0.7, 0.9, 1.2, 0.9, 0.3, 0.4, 1.6, 2.8, 3.8, 
    4.5, 1.3, 3.3, 3.7, 4, 3.4, 2.7, 2.2, 2.7, 2.7, 2, 0.9, 2.5, 2.6, 2.9, 
    2.9, 2.3, 1.9, 2, 2, 1.9, 0.4, 1.3, 2.2, 0.2, 0.8, 2.7, 1.8, 1.2, 3.6, 
    3.7, 3.4, 2.4, 3.3, 3, 2.7, 3.9, 2.8, 2.8, 3.1, 3.1, 3, 3.4, 2.1, 2.8, 
    2.9, 4.5, 4.2, 4.9, 5.1, 5.1, 5.2, 4.7, 5.3, 5.8, 4.5, 4.6, 4, 3.2, 3, 
    3.8, 4.2, 3.7, 4.5, 4.7, 2.1, 0.8, 1.7, 2.2, 2.1, 2.3, 1.9, 1.5, 0.8, 
    1.8, 0.5, 1.9, 1.7, 1.7, 2.3, 4.2, 1.4, 2.6, 3.4, 1.6, 0.7, 2, 0.5, 0.5, 
    3.2, 0.7, 0.5, 0.6, 1.1, 1, 2.2, 1, 3.6, 3.3, 1.7, 1.2, 1.4, 2.4, 2.3, 
    2.2, 1.4, 2.7, 1.1, 0.7, 3.2, 2.7, 1.9, 3.6, 2.3, 0.4, 3, 3, 3, 5.5, 3.8, 
    4, 4.2, 3.4, 4.3, 4.2, 4.5, 5.1, 5.8, 3.5, 5.6, 3.6, 3.3, 3.2, 3.3, 2.4, 
    3.1, 3.5, 3.3, 4.5, 4.2, 4.1, 4.4, 3.6, 3.6, 3.5, 3.6, 4.3, 5, 4.3, 3.8, 
    4.9, 5.2, 4.1, 3.7, 1.6, 3.9, 4.9, 0.3, 0.5, 0.2, 0.6, 1.7, 2.7, 1, 2, 
    2.4, 2.2, 1.7, 2.9, 3.3, 5, 4.7, 2.2, 3.1, 2.7, 5.1, 4.4, 3.6, 1.1, 4.4, 
    1.4, 0.6, 1.8, 0.2, 0, 0.2, 0.1, 4.2, 2.4, 2.8, 3, 6.1, 6.3, 6.4, 6.6, 
    5.8, 5.8, 2.4, 5.4, 4.3, 3, 0.8, 1.1, 0.5, 2, 1.4, 0.6, 2, 3.3, 1.7, 1, 
    0.6, 2.1, 2.1, 1.4, 1.5, 2.1, 1.4, 1.7, 1.9, 0.8, 2.1, 1.8, 2.1, 1.4, 
    1.7, 1.5, 1.6, 1.6, 1.5, 1.8, 1.9, 1.4, 1.5, 0.9, 1, 1.4, 1.2, 1.1, 2, 
    2.1, 2.4, 3.6, 3.2, 3.7, 5, 7, 6.3, 6.7, 5.8, 5.3, 1.1, 3.2, 3.1, 1.9, 
    1.6, 5.6, 4.8, 1.6, 2, 5.2, 2.1, 4.9, 5.1, 6.5, 7.5, 6.5, 6.2, 5, 3.7, 
    2.9, 2.7, 2.3, 2.4, 3.9, 5.6, 5.5, 2.9, 4.1, 1.8, 1.9, 3.9, 4.7, 1.2, 
    3.1, 4.3, 4.8, 5.8, 3.8, 4.3, 6.2, 4.4, 5.1, 4.1, 2.7, 5.1, 5.1, 4.6, 
    3.3, 2, 2, 2.2, 2.3, 1.1, 0.5, 2.1, 1.7, 2.5, 1, 1.6, 1.5, 2.2, 1.6, 1.4, 
    1.6, 3, 2.8, 2.3, 2.2, 1.7, 1.8, 1.1, 2.4, 1.9, 0.3, 1.6, 1.3, 1, 0.7, 1, 
    0.3, 0.3, 1, 0.1, 0.4, 0.8, 0.3, 0.8, 2, 1.5, 1.5, 2, 2, 2, 0.9, 0.8, 1, 
    1.8, 0.1, 0.6, 0.7, 0, 0, 0.1, 0.5, 1.1, 3.5, 1.9, 2, 1.8, 1.6, 1.6, 1.7, 
    2.2, 1.3, 0.4, 2.1, 1.7, 1.8, 1.8, 2.2, 0.7, 1.6, 1.4, 0.9, 0.3, 0.7, 
    0.4, 0.6, 1, 0.7, 0.3, 1.3, 1, 1.4, 1.3, 1.3, 1.6, 1.9, 2.2, 2.3, 1.9, 
    1.7, 1.8, 0.8, 1, 0.6, 0.6, 0.5, 0.8, 1.6, 0.6, 0.5, 1.1, 0.8, 0.8, 1.3, 
    1, 1.3, 1.8, 1.4, 1.4, 2.1, 1.7, 1.6, 2.2, 1.7, 1.3, 1.6, 0.9, 1, 1.6, 
    0.9, 0, 0.1, 0.3, 1.1, 0.8, 1.4, 2.9, 1.5, 3, 2.2, 2.2, 1.1, 2.6, 0.5, 
    2.8, 2.6, 1.5, 1.5, 1.3, 1.3, 2.1, 3.7, 1.8, 1.2, 1.2, 0.4, 3.2, 1.7, 
    0.6, 1, 0.9, 3.3, 1.8, 2.4, 3.2, 5.7, 2.7, 4.3, 7.2, 3, 6.9, 6.5, 7.3, 
    9.1, 6.8, 2.9, 7.3, 8.4, 8, 2.9, 3.2, 2.1, 1.8, 3.1, 2.5, 5.8, 3, 3.7, 
    4.4, 3.9, 1.2, 3.6, 3.5, 1.7, 4.1, 2, 4.6, 6.8, 5.1, 1.8, 1.8, 3, 3.4, 2, 
    1.8, 2.5, 2.8, 2.5, 1.3, 1.5, 2.7, 2.4, 3.2, 3.1, 4, 2.7, 3.7, 1.6, 2.1, 
    1.3, 2.1, 1.8, 1, 2.9, 2.4, 2, 2, 1.6, 1.6, 2, 4.8, 2.1, 1.5, 3, 2.3, 
    2.5, 2.5, 3.1, 6.2, 3, 5.9, 4.5, 2.6, 3.6, 4.6, 3.3, 2.4, 3.9, 1.9, 3.4, 
    2.3, 3.3, 3.3, 2.4, 3.5, 2.9, 3.1, 4, 3.9, 1.4, 2.8, 4.9, 5.2, 3.6, 3.4, 
    4.2, 2.9, 3.9, 4.8, 5.1, 4.5, 3.1, 3.5, 2.1, 1.2, 0.7, 1.5, 0.8, 0.2, 
    0.1, 0.9, 0.9, 2, 3.1, 2, 1.8, 1.7, 2.3, 1, 2, 2, 2.8, 2, 2.2, 2.8, 2.3, 
    0, 0.2, 0.8, 0, 0.6, 1.5, 2.4, 0.6, 0.4, 0.9, 1.3, 1.1, 2.1, 0.3, 2.2, 
    1.7, 1.4, 2.1, 1.3, 1.2, 0.6, 2.6, 1.9, 1, 0.9, 0.9, 1, 0.7, 0.3, 1.4, 
    0.1, 0.2, 0.8, 1.9, 2.2, 1.6, 2.1, 5.2, 1.9, 2.4, 3.2, 3.7, 6.1, 1, 1.5, 
    2.2, 7.5, 6.9, 2.3, 6, 8, 3.6, 10, 8.2, 5, 7.6, 8.1, 8.5, 3.2, 7.3, 5.5, 
    5.3, 5.7, 3.1, 2.6, 2.1, 2.6, 2.4, 2.6, 2.1, 2.4, 3.3, 2.5, 5.3, 2.1, 
    1.4, 4.7, 2.6, 2.7, 4.1, 1.8, 1, 0.7, 2.1, 0.6, 3.5, 2, 3, 3.2, 2.9, 3.4, 
    1.6, 0.2, 2.8, 0.1, 0.9, 0, 0.3, 0.4, 0.7, 0.4, 0.3, 0, 0.5, 1.2, 1.5, 
    2.6, 3.6, 3.7, 3.8, 3.9, 3.5, 5.4, 3.3, 3.2, 3.2, 1.6, 2.9, 2.8, 2.3, 
    3.3, 1.8, 2.2, 1.8, 0.7, 2.3, 0.8, 1.2, 2.1, 2.6, 0.8, 2.3, 1.5, 2.9, 
    3.2, 2.9, 2.7, 3, 2.9, 2.4, 2.2, 2.2, 1.9, 1.5, 0.8, 2.1, 3.3, 1.6, 0.4, 
    0.5, 0.5, 0.2, 2.5, 3.6, 2.8, 2.6, 2.7, 3.3, 2.2, 3, 2.2, 1.1, 1.3, 2.5, 
    2.3, 2.8, 0.8, 1.2, 0.9, 0.9, 0.1, 1.6, 1.1, 2.3, 4.6, 6.6, 7, 7.5, 4.8, 
    7.6, 3.7, 5.7, 5.5, 6.8, 6.1, 4.3, 7.9, 3.7, 1.3, 5.8, 3.7, 4.7, 4, 4.7, 
    2, 4.6, 4.1, 2.7, 0.1, 2.4, 0.8, 0.1, 0.6, 0.6, 1.2, 0.8, 5, 2.2, 1.8, 
    1.8, 3.6, 1.4, 2.5, 1.9, 0.5, 0.2, 0.1, 1.2, 0.5, 0.1, 0.2, 0.5, 0.2, 
    1.2, 0.5, 0.2, 0.8, 0.3, 0.8, 1.4, 0.8, 1.5, 2.5, 2.8, 3.2, 4.5, 3.7, 
    1.1, 1.4, 4.7, 1.8, 1.4, 0.8, 1.6, 2, 0.9, 1.5, 0.6, 0.8, 1.4, 4.7, 3.8, 
    0.8, 3, 3.4, 5.7, 6, 7, 2.1, 2.2, 4.7, 4.9, 6.3, 5.4, 4, 4.6, 0.3, 1.7, 
    0.5, 0.4, 0.5, 0.5, 0.2, 3.4, 2.6, 4.2, 4.9, 4.6, 5, 5.1, 2.8, 2.9, 6.7, 
    3.4, 2.9, 3.1, 2.7, 1.5, 2.9, 3, 0.9, 0.5, 2.1, 1.3, 0.9, 0.3, 1, 0.3, 
    1.7, 0.9, 0.5, 2.1, 3.4, 6, 4.2, 3.4, 1, 1.2, 2.8, 2.3, 2.1, 0.5, 0.1, 
    1.1, 1.4, 0.8, 1.1, 0.9, 0.7, 0.9, 1.4, 0.5, 1.1, 1.8, 2.2, 1, 1.2, 1.6, 
    3.8, 3.4, 0.2, 1, 3.8, 3.8, 3.4, 3.5, 3.7, 2.6, 1.9, 2.5, 0.3, 2.5, 1.4, 
    2.6, 1.4, 1.9, 2.4, 2, 1.2, 2.8, 1.9, 1.3, 0.8, 0.8, 1.1, 1.5, 0.1, 0.4, 
    1.2, 0.4, 0.7, 1.3, 1.4, 0, 0, 0, 0, 1.3, 1.2, 0.4, 1.2, 0.3, 0.3, 0.5, 
    0.5, 1.2, 2.6, 0.7, 3.5, 2, 3.4, 3.5, 2.6, 3.8, 3.3, 3.4, 1.9, 2.5, 0.7, 
    3.8, 0.9, 0.8, 1.6, 0.5, 0.8, 0.5, 1, 1.4, 2.4, 1.8, 2.5, 2.5, 0.9, 1.2, 
    2.8, 2.5, 1.5, 2.2, 1, 0.7, 1.6, 0.9, 0.5, 0.5, 1.4, 0.6, 1.5, 1, 1.5, 
    3.2, 2.9, 4.1, 3.6, 2.9, 1.4, 5.1, 3.1, 5, 3.4, 3.6, 3.2, 2.4, 2.1, 1.9, 
    2.1, 1.2, 0.6, 1.3, 2.3, 2.1, 1.3, 1.4, 1.5, 1.8, 1.4, 1.8, 2.2, 2.1, 
    2.6, 1.7, 1.8, 1.2, 0.8, 1.1, 2.6, 1.3, 4.2, 4.4, 3.2, 2.8, 2.6, 3, 2.6, 
    2.5, 3.3, 2.7, 3.9, 3.2, 2.5, 1.6, 2.3, 2.8, 2.9, 2.9, 1.7, 1.7, 1.2, 
    0.5, 0.2, 0.3, 0.8, 0.5, 0.5, 0.2, 2, 1, 0.9, 0.9, 1.1, 0.4, 0.3, 1, 1.4, 
    0.8, 0.8, 1.6, 1, 1.2, 1.4, 0.8, 1, 0.9, 1, 0.3, 0.3, 0.8, 1.7, 0.4, 0.5, 
    0.2, 1.2, 1.1, 0.9, 0.8, 2.8, 1.5, 2, 0, 1.1, 0.9, 1.4, 1.3, 1.6, 1.2, 
    2.3, 1.5, 1.3, 1.1, 0.4, 0.7, 0.3, 0, 0.3, 0.3, 0.7, 0.1, 0.2, 1.1, 0.6, 
    1.2, 1.7, 1.4, 2, 1.8, 1.2, 1.9, 1.3, 0.8, 0.2, 0.1, 1.3, 2.3, 1.8, 0.6, 
    0.3, 0.9, 0.2, 0.3, 0.7, 0.8, 0.3, 0.8, 0.5, 0.5, 1.3, 1.4, 1.3, 1.5, 
    1.6, 1.7, 1.8, 1.9, 2.1, 1.9, 1.5, 1.3, 1.2, 1.3, 1.5, 1, 0.2, 1.1, 0.7, 
    0.2, 0.1, 0.9, 0.4, 3.5, 4.9, 3.5, 3, 3.6, 3.1, 3.3, 2.6, 2.8, 2.1, 2.5, 
    2.5, 2.6, 2.2, 1.9, 1.8, 1.9, 1.8, 2.5, 2.1, 1.5, 1.6, 0.3, 1.6, 0.9, 
    3.9, 3.5, 3.5, 2.3, 2.1, 1.7, 1.7, 1.6, 1.3, 1.8, 1.5, 1.3, 0, 0.8, 0.4, 
    0.9, 1.1, 0, 0.1, 1.2, 0.6, 1.3, 1.5, 0.8, 1, 0.9, 0.4, 0.1, 0.4, 0.4, 
    0.4, 0.1, 0.6, 0.8, 0, 0.2, 0, 1.1, 0.4, 0.5, 0.4, 0.1, 0.1, 0, 0.8, 0.1, 
    0.3, 0.4, 0.6, 1.2, 2.1, 1, 0.6, 1.3, 0.1, 1.4, 2, 1.7, 1.3, 0.2, 0.1, 
    1.1, 2.1, 3.4, 1.3, 4, 3.8, 3.3, 1, 2.6, 4.1, 3.9, 6.1, 6.7, 5.3, 4.7, 
    7.4, 6.5, 5, 5.4, 5.7, 4.7, 5.5, 4.9, 2.9, 3.7, 3.3, 2.1, 4.7, 3.3, 1.1, 
    4.4, 8.9, 9, 7.7, 7, 6.9, 7.7, 5.5, 6.3, 5.8, 5.4, 4.9, 4.8, 3, 3.4, 2.5, 
    3.1, 2.3, 2.4, 2.9, 2.9, 2.8, 2.5, 1.7, 1.6, 0.7, 3.4, 2.8, 3.5, 4.1, 
    3.8, 4.5, 4.2, 3.2, 2, 1.9, 1.8, 1.6, 1.3, 1.4, 0.7, 0.7, 1.7, 2.7, 3.8, 
    1.5, 0.3, 1.8, 0.1, 0.9, 1.2, 3.2, 1.5, 1.5, 2.1, 2.2, 1.2, 2.5, 2.2, 
    2.3, 2.4, 3.4, 1.7, 1.3, 2.6, 1.3, 0.9, 0, 0.7, 0.9, 0.3, 0.3, 0.2, 0.2, 
    0.3, 0.3, 0.8, 1.2, 1.4, 1.7, 2.7, 3, 3.4, 3.7, 3.5, 4.7, 4.5, 2.8, 3.9, 
    2.7, 3.7, 3, 1.7, 0.6, 2, 4.2, 3.9, 3.8, 1.7, 3.1, 3.4, 3.4, 2.9, 1.3, 
    0.7, 2, 1.2, 1.8, 1.3, 0.8, 1, 0.8, 0.5, 0.4, 1.4, 1.2, 1.4, 0, 0.3, 0, 
    0.6, 0.6, 0.8, 0.1, 0.7, 0.6, 0, 0.6, 0.7, 1.1, 0.6, 0.2, 0.1, 0.4, 2.1, 
    2, 2.8, 2.4, 1.8, 0.7, 2.2, 0.1, 1.4, 0.1, 0.4, 0.8, 0.1, 0.6, 1.5, 1.2, 
    1.1, 1.7, 1.3, 1.3, 2, 1.8, 1.6, 1.3, 1, 1.6, 1, 1, 0.6, 0.9, 0.2, 0.7, 
    0, 0.4, 0.4, 0.3, 0.2, 0.8, 0.6, 1.8, 1.7, 1.5, 1.7, 2, 2, 2.2, 2, 1.9, 
    1.2, 1.3, 0.9, 1, 0.1, 0.3, 0.7, 1.9, 2.3, 2.6, 2.3, 2.5, 3.2, 2, 1.9, 
    1.1, 0.3, 1.9, 2, 0.4, 0.6, 1.2, 1.9, 2.5, 2.7, 2.3, 2.9, 0.5, 0, 1, 0.9, 
    0.9, 0.1, 0.2, 0, 0.2, 0.3, 1, 1.5, 0.6, 2, 2.7, 2.8, 3.7, 3.7, 3.5, 2.6, 
    3.9, 3.7, 3.6, 2.7, 2.9, 0.1, 0.9, 1.2, 0.3, 3.3, 1, 1.8, 3, 1.8, 0, 0, 
    0, 0, 1.2, 0.1, 0.2, 1.8, 1.4, 5.9, 5.3, 6.2, 3.9, 3.3, 4.1, 2.4, 2.7, 
    3.2, 5.8, 3.4, 3.6, 2.6, 2.5, 3.9, 4.1, 2.3, 2.2, 2.3, 1, 2.1, 1.4, 1.5, 
    2.6, 2.2, 1.8, 2.4, 4.8, 4.1, 6.3, 4.1, 2.6, 2.9, 3.8, 2.9, 2.8, 2.3, 
    4.3, 4.3, 4.9, 5.1, 2.7, 4.1, 3.7, 2.9, 2.4, 3.5, 4.1, 3.6, 3.8, 3.9, 
    3.5, 4.7, 5.7, 6.6, 4.3, 1.4, 6, 6.1, 6.5, 6.3, 6.3, 4.3, 2.2, 3.5, 6.8, 
    5.4, 5.7, 6.2, 5.7, 6.4, 5.9, 5.1, 5.1, 3.3, 1.1, 0.6, 1.8, 1.6, 2.1, 
    1.8, 0.5, 0.6, 1.7, 1, 1.1, 1.5, 2.3, 2.6, 1.3, 1, 1.1, 2, 0.9, 3.4, 2.6, 
    0.5, 1.9, 1.3, 0.4, 1.7, 1.2, 1.6, 1.3, 1.6, 0.8, 1.8, 1.5, 0.9, 1.3, 
    1.1, 1.8, 3.7, 3.9, 3.6, 4.1, 3.9, 3.9, 5.7, 5.7, 2.8, 4, 1.5, 3.2, 1.9, 
    2.4, 1.5, 6.1, 4.3, 2.6, 1.4, 1.9, 1.7, 0.7, 0.7, 0.3, 0.1, 0.6, 0, 3, 
    3.8, 4.6, 2.9, 1.1, 1.3, 1.7, 2.5, 4.7, 3.4, 1.2, 4.6, 5.2, 4.4, 3.3, 
    0.7, 1.1, 0.8, 0.8, 1.3, 1.8, 1.6, 0.1, 0.4, 0.1, 0.6, 1.6, 1.3, 0.8, 
    0.1, 0.1, 0.2, 0, 0, 0.8, 0, 0, 0.6, 0.7, 0.3, 0, 0, 0.7, 0.1, 0.6, 2.3, 
    0.4, 1.1, 0.7, 1.2, 0.3, 0, 0.9, 0.5, 0.5, 0.6, 0.1, 1.2, 1, 0.9, 1.1, 0, 
    0.7, 0, 0.5, 1.1, 0.2, 0.9, 0.3, 0.3, 1.5, 7.1, 3.2, 3.8, 4.2, 3.2, 0.7, 
    2.5, 2.2, 3.9, 4.3, 5.7, 7.4, 4.3, 5.2, 5.6, 4.6, 4.6, 4.8, 6.4, 5.7, 
    4.1, 3.6, 3.8, 5.2, 5.2, 5.2, 4.7, 4.9, 4.7, 4.1, 4.3, 5.4, 5, 4, 2.5, 
    3.2, 3.5, 2.1, 4, 3.5, 1.6, 1.9, 2.9, 1.9, 2.3, 2.9, 3.1, 2.7, 2.7, 2.4, 
    1.6, 1.1, 1.6, 3.3, 2.2, 2.5, 1.3, 0.6, 2.2, 1.3, 1.1, 0.8, 0, 0.6, 1.1, 
    1.8, 3.1, 2.9, 0.8, 0.8, 0.3, 0.5, 1.8, 0.4, 2, 3.9, 0.8, 0.1, 1, 0.8, 
    2.1, 2.4, 3.1, 3.5, 2.3, 2.9, 1.7, 1.3, 0, 0, 0, 0, 0, 0, 0, 0.5, 0.4, 0, 
    0.1, 0.9, 1.1, 4.2, 5.1, 6.1, 4.7, 6.3, 4.3, 5.2, 4.1, 4.6, 3.6, 4.6, 
    3.6, 4.2, 3.8, 3.5, 3.7, 3.7, 3.8, 2.9, 2, 1, 0.7, 1, 0.8, 2.3, 1.5, 1.2, 
    0, 0, 0.3, 0.7, 0.4, 0.2, 0.4, 6, 6.7, 3.3, 3.1, 5.7, 4.7, 3.5, 2.2, 2.4, 
    4.7, 3.3, 3.1, 4.2, 3.9, 2.9, 3.2, 1.9, 0.7, 1.3, 1.4, 1.3, 2, 2.1, 0.3, 
    3, 0.4, 0.3, 1, 0.3, 0, 1.2, 0.9, 0.7, 0.2, 0.1, 0, 0.5, 0.1, 0.1, 0.1, 
    0.1, 0.9, 1.3, 0, 0.8, 1, 0.8, 1.2, 0.1, 1.9, 0, 0.7, 0.6, 0.6, 0.9, 6.4, 
    0.6, 1.2, 1.3, 0.3, 0.5, 4.9, 3.2, 1, 0.5, 1.1, 0, 0.5, 0.9, 2.2, 0.9, 
    1.1, 1.5, 0.1, 0, 0.3, 1, 0.6, 0.3, 0.8, 0, 0.1, 0.5, 0.8, 3, 0.6, 0.6, 
    0.9, 0.8, 1.1, 0, 0.3, 0.1, 0.3, 0.4, 1.1, 1, 2, 3.2, 3, 1.9, 0.5, 0.7, 
    0.1, 0.8, 0.7, 0.8, 0.5, 0.3, 0.5, 0.3, 0.5, 1.6, 3, 1.8, 0.6, 0.7, 1.2, 
    1.4, 0.9, 1.9, 0.7, 0.7, 1.2, 0.3, 0.7, 0.6, 1.4, 0.4, 0.6, 0.9, 1, 0.3, 
    0.8, 2.6, 0.1, 0.1, 0, 0, 0.2, 0.9, 1.3, 0.4, 0.5, 0.2, 0.1, 0.2, 0.2, 
    3.7, 1.9, 2, 2.6, 2.6, 2.1, 0.5, 1.8, 4, 3.7, 0.9, 1.9, 1.4, 1.5, 1.6, 
    0.3, 0.9, 0.4, 0.5, 0.7, 0, 0, 0.2, 0, 0.9, 0.2, 1.4, 0.4, 0.6, 1.9, 1, 
    0.6, 1.1, 0.5, 1.1, 0.1, 0.9, 2.1, 2.2, 2, 2, 2, 2, 1.1, 0.7, 1.1, 0.1, 
    0.4, 0, 0.5, 0.1, 1.2, 0.1, 0.6, 1, 0.6, 0.7, 1.3, 2, 1.6, 0.2, 0.3, 0.2, 
    0.4, 0, 0.7, 0.5, 0.1, 1.1, 1, 2.9, 1.2, 0.5, 0.3, 0.3, 0.8, 0.1, 2, 0.7, 
    0.8, 4.1, 0.8, 0.8, 0.4, 1, 1, 0.8, 0.7, 0.2, 0.4, 0.9, 0.1, 0.5, 0.9, 
    0.7, 0.7, 0, 0.3, 0.9, 0, 1.4, 1, 1.2, 1.3, 2.2, 0.1, 0.1, 0.1, 0.8, 0.6, 
    0.8, 0.4, 0.5, 0.9, 0.2, 1.3, 1.1, 0.8, 1, 0.5, 0.2, 0.5, 0.2, 1.4, 0, 
    0.9, 0.5, 1.7, 0.4, 0.2, 0.3, 0.8, 0.4, 0.9, 0.5, 0.2, 0, 0, 1.1, 0.5, 0, 
    0, 0.2, 0.2, 1, 0.6, 0.2, 0.3, 0.3, 0.9, 0, 0, 2.6, 3.1, 0.2, 0.2, 0.1, 
    0.1, 0.5, 0.4, 0.1, 0.1, 0, 0.5, 0.1, 0.9, 0.7, 1.2, 0.1, 0.9, 0.6, 0.4, 
    0.4, 1.2, 0.9, 0.6, 0.8, 0.7, 0.2, 0.5, 0.1, 0.2, 0.1, 0.3, 0.8, 0.1, 
    0.1, 0.8, 0, 0, 0.1, 0.5, 0, 0, 0, 2.3, 0, 0, 0, 0.1, 0.5, 0.5, 0.9, 0, 
    2.2, 0.3, 0.4, 0.1, 2.7, 0.7, 0.3, 0.7, 1, 1.9, 1.6, 0.6, 4.2, 0.6, 0.7, 
    0.6, 0.7, 0.4, 0.5, 0.3, 0.2, 0.4, 0, 1.4, 1.4, 2.4, 0.9, 1.5, 0.3, 1.3, 
    0.7, 1, 1.3, 0.6, 0.7, 0.6, 2.5, 1.5, 1.7, 1.6, 0.6, 3.6, 1.2, 0.8, 3.1, 
    4.6, 4.6, 5.3, 5.4, 5.4, 5, 4.6, 8.5, 8.1, 8.7, 6.1, 1.4, 4, 5.2, 4.2, 
    4.4, 6.7, 5.8, 10, 9.8, 4.5, 5.9, 5, 6.7, 7.9, 6.2, 6.7, 7, 5.7, 4.9, 
    5.3, 5, 3.9, 5.1, 4.2, 2.6, 4.2, 4.2, 4, 4.9, 3.5, 3.3, 3.3, 3.3, 2.8, 
    2.9, 3, 3.8, 3.8, 1.3, 1.9, 1, 0.4, 0.2, 0, 0.5, 0.8, 2.3, 2.2, 2.2, 0.4, 
    2.8, 1.2, 1.5, 1.5, 1.5, 1.6, 1, 2.7, 1, 0.1, 2, 1.1, 0.7, 0.6, 0.7, 0.3, 
    0.3, 0, 0.6, 0, 0.2, 0.1, 0.1, 0, 0.8, 0.8, 1.6, 0.3, 1, 0.5, 0.4, 0.8, 
    0.6, 0.7, 1.2, 0.9, 0.9, 0.1, 0.1, 0.1, 0.5, 1, 0.5, 0.5, 0.2, 0.3, 0.3, 
    0.1, 0.8, 0.9, 0.9, 0.7, 1.2, 0.6, 0.9, 1.3, 0.7, 0.7, 1, 0.1, 2.1, 0.2, 
    0.8, 0.4, 0.4, 0.6, 0.1, 0.5, 0.8, 0.5, 0.4, 0.4, 0.2, 0.9, 0.7, 1.1, 
    0.3, 0.9, 0.2, 1.2, 0.2, 0.1, 0.4, 0.1, 0.5, 0, 0.1, 0.4, 0.5, 0.6, 0.7, 
    0.5, 2, 1.2, 0.9, 1, 1.7, 2.4, 1.3, 1.1, 0.2, 2.6, 3.1, 0.5, 0.2, 0, 1.6, 
    0, 0, 0.8, 0.9, 1, 0.2, 0.2, 0.3, 0.4, 0.9, 0, 1.1, 0.9, 0.8, 0.2, 0.3, 
    0.6, 1.1, 1.2, 0.9, 0.3, 0.4, 1.5, 0.4, 2.1, 0.7, 1.2, 0.6, 0.9, 0.5, 
    1.1, 0.8, 0, 1, 0, 0.5, 0.1, 0.1, 0.1, 0.8, 0.4, 0, 0, 0.4, 1.1, 0.2, 
    0.4, 0.4, 0.1, 0.9, 1.6, 1.3, 0.1, 0.2, 0, 0, 0.2, 0, 0.3, 0.2, 0, 0, 
    0.2, 0.3, 1.5, 0.1, 2.9, 2.8, 0.1, 0.2, 0.2, 0.1, 0.3, 0.9, 0, 1.3, 1.6, 
    2.8, 0.5, 0.7, 1, 0.7, 0.4, 1.5, 0.5, 1.3, 0.6, 1, 0.7, 1.2, 0.4, 0.4, 
    0.2, 0.6, 0.3, 0.1, 2, 0.3, 0.5, 0.7, 1.1, 0.4, 1.9, 1.3, 0.3, 1.3, 0.8, 
    2.9, 2, 1.3, 0.9, 0.9, 0.5, 0.7, 0.1, 0.3, 4, 0.1, 0.8, 0.4, 0.1, 0.9, 
    0.9, 0.3, 0.7, 1, 1.5, 0.3, 0.9, 0.2, 0.9, 0.9, 0.4, 0.5, 0.1, 0.4, 0.3, 
    0.6, 2, 1.8, 0, 0.2, 0, 0.8, 0.5, 0.1, 0.6, 0.6, 0.2, 0, 0.5, 0, 0.3, 
    0.5, 0, 0.9, 1.6, 1, 0.1, 0.1, 0.4, 0.6, 0.3, 0.2, 0, 0.8, 0, 0, 0.4, 
    1.7, 0.6, 1.4, 2.1, 0.5, 0.4, 2, 0, 1.2, 0.2, 0.8, 0.5, 1, 3.7, 0.4, 0.6, 
    1, 0.6, 1, 3.8, 2.9, 5.5, 5.8, 6.1, 4.4, 2.2, 6.3, 5.1, 4.8, 4, 0.9, 1.4, 
    1.7, 1.3, 0.5, 0.8, 1.8, 0.6, 0.8, 1.1, 0.1, 0.9, 0.6, 0, 0.6, 0.1, 0.2, 
    0.3, 0.3, 0, 0.1, 0.5, 0.2, 0.1, 0, 0, 1, 5.1, 4.7, 2.5, 4.4, 5.1, 4.6, 
    4.6, 4.8, 5.1, 4.6, 5.2, 3.7, 3.6, 6.2, 5, 3.7, 3.4, 1.6, 2.5, 0.5, 0.2, 
    0.2, 0.5, 1.2, 0.6, 0.1, 1.3, 1.1, 0.3, 0.3, 0.5, 1.4, 0.9, 1.9, 4.3, 
    4.2, 2.8, 1.2, 1.6, 0.5, 1.1, 0.3, 1, 0.1, 0.2, 1, 0.3, 1.1, 0.6, 1.1, 
    1.7, 2.2, 1.5, 0.5, 1.3, 0.4, 2.1, 2.2, 0.9, 2.1, 1.3, 1.1, 1.1, 0.1, 1, 
    1, 2.3, 2.1, 0.4, 0, 0.6, 0.8, 1.5, 1.2, 0, 0, 0, 0, 1.1, 2.3, 1, 0.5, 
    7.2, 7.3, 8.5, 7, 6.3, 4.9, 3.6, 4.5, 1.9, 4, 5.8, 6.9, 8.4, 7.5, 9.9, 
    8.9, 9.1, 9.7, 6.3, 8.7, 6.8, 6.4, 5.9, 5.4, 6, 5.1, 3.1, 4.2, 5.4, 4.4, 
    5, 4.5, 3, 2.6, 2.4, 3.3, 2.2, 2.9, 2.9, 3.8, 3.5, 4, 3.1, 3.8, 5.1, 3.6, 
    3.4, 3.8, 4, 3.3, 4, 5.5, 5.9, 7.1, 5.2, 4.7, 5.4, 6, 5.7, 6.1, 6.5, 6.5, 
    5.8, 7.5, 8.6, 9.4, 7.5, 7.2, 6.4, 7.3, 8.5, 7.7, 8.3, 6, 8.2, 8.9, 7.5, 
    8.5, 7.9, 7.2, 7.6, 6.9, 7.6, 6, 6.9, 8.5, 7, 7.7, 7.9, 7.3, 7.9, 7, 7.5, 
    6.6, 7.4, 8.3, 7.2, 9.1, 8.7, 8.8, 9.6, 10.6, 10.2, 10.1, 8.7, 10, 9.8, 
    8.6, 9.8, 9.6, 8, 6.1, 4.7, 3, 1.3, 1.7, 3.1, 1.6, 0.3, 2.5, 2.7, 1, 0.8, 
    0.8, 0.5, 6.2, 6.3, 5.7, 4.8, 5.8, 5.5, 5.7, 5.2, 2.8, 3.6, 2.2, 2.3, 
    2.1, 1.6, 7.1, 6.9, 5.8, 4.6, 7.6, 1.8, 1.4, 4.4, 3.3, 5, 5, 4.8, 3.6, 
    4.5, 3.4, 2.4, 7.7, 9.3, 8.9, 9.8, 7.9, 5.5, 3.7, 6.7, 8, 6.9, 5.6, 2.5, 
    1.4, 1.9, 3.3, 6.2, 5.7, 6.5, 4.9, 1.6, 1.1, 0.5, 2.1, 0.4, 1.5, 1.5, 
    0.3, 1.7, 1.9, 0.7, 0.7, 0.9, 0.5, 0.7, 0.1, 0.1, 2.8, 1, 1.1, 1.2, 0.7, 
    1.2, 0.8, 0.5, 0.6, 0.3, 0.5, 0.2, 0.2, 0.3, 0.1, 0.3, 0.5, 0.6, 0.7, 
    1.1, 0.5, 0.7, 0.2, 1.4, 2.7, 3.6, 3.7, 4.1, 4.3, 4.2, 3.5, 3.6, 3.8, 
    3.8, 2.6, 2.3, 0.2, 1.6, 0.1, 0.5, 0.4, 1.1, 1.3, 1.5, 2.4, 2.1, 1.5, 
    0.3, 1.3, 0.7, 0.6, 0.5, 0, 0.8, 0.1, 0.1, 1, 1.2, 0, 0.9, 1.8, 1.2, 1.9, 
    2, 0.4, 0.6, 0.5, 1.3, 1, 0.3, 0, 0, 4, 2.9, 3.1, 5.4, 5.8, 5.5, 4.4, 
    3.9, 3.9, 4.4, 3.4, 2.9, 4, 5.2, 3.4, 3.1, 4.3, 4.7, 3.3, 3.5, 4, 4.2, 
    5.8, 5.5, 5.4, 4.2, 4.5, 2.8, 3.2, 1.4, 1.2, 0.4, 1.7, 1, 4.4, 1.1, 0.9, 
    0.7, 1.8, 0.2, 1.2, 2.7, 0.9, 0.7, 0.4, 0.8, 0.2, 0.4, 0.3, 0.4, 0.4, 
    0.9, 0.2, 0.2, 0.9, 0.8, 0.4, 0.4, 0.7, 0, 0, 0.1, 0.2, 0, 0.4, 0.2, 0.3, 
    0.1, 0, 0.1, 0.2, 0.6, 0.8, 0, 0.2, 0.3, 1.1, 0.9, 0.9, 2.3, 4.9, 2.9, 
    7.2, 6.3, 5.2, 6.4, 4.9, 4.3, 5.2, 4.3, 5.7, 6.6, 4.7, 4.7, 4, 2.3, 3.8, 
    0.2, 1.1, 1.5, 1.3, 3.8, 0.7, 3.7, 2.8, 0.8, 2.9, 0.1, 0.8, 0.6, 0.7, 
    1.3, 1, 0.4, 1.8, 1.9, 2.8, 1, 3.5, 0.1, 0.2, 0.3, 0.3, 1.3, 0.6, 1, 2, 
    4.9, 5.1, 4.4, 3, 4.3, 6.1, 2.4, 3.3, 1.4, 1.7, 0.6, 3.6, 1.7, 0.5, 1.7, 
    1.8, 3.2, 2.9, 3.1, 4.7, 4, 6.1, 5.3, 3.3, 2.7, 2.2, 1.7, 1.4, 2.2, 2, 
    1.9, 0.9, 0.5, 1.4, 0.2, 0.6, 1, 1.8, 0.9, 0.9, 0.5, 2.5, 2.9, 1.2, 1.1, 
    0.5, 1.8, 0.9, 0.7, 1.1, 1.1, 0.7, 0.1, 0.5, 1.6, 0.8, 1.3, 0.7, 0.8, 
    1.4, 1, 1.4, 0.8, 1.9, 0.2, 1.4, 1, 0.8, 0.6, 1.2, 0.9, 0.3, 0.2, 0.2, 
    0.5, 0.9, 0.5, 0.9, 1.4, 0.2, 1, 1.1, 0.7, 5.2, 1, 1.2, 1, 1.2, 0.9, 0.8, 
    7.8, 0.9, 1, 0.7, 1.9, 2.4, 1.8, 2.2, 1.7, 0.5, 1.3, 0.3, 0.3, 0.9, 5.9, 
    0.1, 2.1, 0.1, 1.3, 1.6, 0.4, 0.9, 1.9, 1.6, 2.1, 1.1, 0.1, 1.5, 0.8, 
    0.7, 1, 1.3, 0.2, 1.3, 0.4, 1.1, 0.4, 1.1, 1.1, 0.8, 4.4, 4.5, 4.8, 6.4, 
    6.4, 7.1, 6, 7.2, 6.4, 6.7, 6.2, 6.9, 7.2, 8.2, 6.9, 7.7, 9.1, 8.3, 6.7, 
    5.9, 7.2, 7.1, 6.1, 5, 5.9, 6.1, 4.6, 5.1, 2.1, 1.7, 0.7, 6.5, 5.2, 4, 
    4.6, 3.3, 4.1, 3.2, 3.5, 2.4, 3.5, 4.8, 6.9, 5.1, 4.5, 3.9, 1.7, 0.7, 
    4.7, 3.1, 3.8, 3.1, 2.7, 3.3, 7.4, 4.4, 4.7, 4.4, 4.5, 3.9, 2.1, 1.9, 
    2.8, 3.1, 3.4, 2.4, 2.8, 4.2, 4.7, 3.8, 4.4, 4.2, 3.2, 4.5, 3.5, 5.4, 
    3.5, 4.1, 3.5, 2.7, 4.9, 4, 4.7, 6.7, 5.5, 6.1, 6.5, 6.1, 6.6, 7.5, 5.7, 
    7.5, 6.5, 8, 8.4, 5.8, 6.5, 5.1, 6.3, 6, 7.5, 7.7, 6.9, 7.3, 6.2, 7, 7.4, 
    6.6, 7, 6.7, 6.3, 4.3, 6.2, 8.5, 9, 7.7, 8.9, 7.5, 6.4, 6.5, 8.1, 7, 7.5, 
    6.8, 3.7, 9.5, 10, 9.6, 6.6, 2.7, 4.2, 4.9, 6.3, 6.2, 6.2, 4.9, 4.5, 5.2, 
    5.2, 3.4, 4.7, 5.1, 3.7, 3.8, 4.7, 5, 4.1, 4.8, 2.7, 5.5, 2.4, 2.4, 3.8, 
    3.4, 2.6, 1.2, 1.1, 0.8, 0.6, 0.7, 0.4, 0.1, 0.5, 0, 0.4, 0.3, 0.5, 1, 
    0.7, 3.1, 3.3, 2.1, 0.9, 0.7, 0.6, 0.7, 3.8, 0.8, 0.8, 0.2, 1.1, 1, 0.2, 
    1.1, 0, 1.2, 3.7, 6.4, 7.8, 7.8, 9.9, 8.1, 3, 5.1, 4.3, 6.7, 5.9, 6, 8.4, 
    5.2, 0.9, 1.2, 1.5, 2.7, 4.9, 5.4, 4.6, 4.5, 0.2, 0.8, 1.2, 3.4, 1.8, 1, 
    1.7, 1.9, 1.3, 1.9, 1.4, 6.1, 2.7, 2.7, 5.7, 6, 4.9, 1.5, 1.7, 1.1, 1.1, 
    0.5, 0.8, 1.5, 1.6, 2.3, 1.1, 0.8, 2.2, 1.2, 1, 1.7, 1.1, 6.5, 1, 1.1, 
    1.1, 1.7, 0.7, 0.5, 0.5, 1.8, 3.6, 2.2, 0.3, 2.2, 3.2, 3.6, 3.3, 0.2, 
    1.8, 3.9, 2.9, 3.3, 3.4, 4.2, 3.8, 2.8, 3.7, 3.4, 3.4, 3.3, 4, 0.2, 0.3, 
    0.5, 0.5, 0.2, 1, 1.2, 1.3, 0.5, 0.9, 0.7, 1.1, 0.7, 0.8, 0, 1.3, 2.1, 
    2.5, 0.6, 3.1, 5.1, 1.4, 0.2, 0.2, 0.7, 1.9, 0.6, 4.2, 4.6, 4.8, 4, 4.7, 
    4.4, 4, 4.4, 1.2, 2, 5.5, 2.9, 4.3, 3.7, 5.4, 5.2, 5.1, 4.5, 4.9, 3.2, 
    2.2, 1, 0.1, 0.2, 1.3, 1.4, 1.6, 2, 4.8, 1.3, 2.4, 2.2, 1.8, 1.4, 2.4, 
    1.9, 5.9, 3.5, 2.9, 1.5, 1.3, 0.7, 2, 1.7, 4.5, 1, 0.9, 0.7, 1.6, 1, 2.4, 
    1.5, 2.3, 3.1, 1.1, 2, 1.8, 0.7, 0.9, 1.6, 1.2, 2.5, 1.3, 0.6, 0.8, 1.3, 
    1.9, 0.7, 0.7, 1.3, 0.6, 1.3, 0.8, 4.9, 4.5, 4.6, 4.9, 4.1, 4.2, 4.4, 
    5.4, 4.4, 4.7, 5, 4.8, 3.6, 1.2, 4.4, 0.8, 4.7, 0.4, 4.2, 4.6, 4.5, 6, 5, 
    5.5, 5.5, 7.3, 5.9, 8.7, 7.4, 8.6, 8.4, 7.6, 7.8, 8.6, 7.7, 6.8, 7.8, 
    8.8, 8.8, 7.9, 8.3, 7.1, 8, 4.7, 9.5, 7.2, 6.7, 8.2, 7.7, 8.8, 8.3, 6.9, 
    8.5, 9.6, 10, 10.1, 8.4, 8.2, 6.8, 7.9, 8.8, 8.8, 10.3, 8.2, 8, 8.6, 7.5, 
    8.7, 7.7, 7.6, 7.1, 7.5, 7.1, 7.3, 6.6, 6.3, 7.8, 8, 7.8, 7.3, 7.2, 7.9, 
    7.1, 8, 7.4, 7.4, 9.7, 10.5, 13.9, 10, 8.8, 5.9, 13.3, 10.7, 10.4, 10.9, 
    5.1, 5.8, 4.7, 6, 4.8, 3.9, 5.6, 3.9, 5.1, 4.7, 2.6, 8.2, 2.9, 3.6, 2.9, 
    4.7, 5, 4.4, 5.3, 5.2, 7.8, 3.7, 4.4, 7.8, 6.1, 4.2, 6.8, 9.6, 9.8, 9.1, 
    9.2, 6.6, 7.9, 9.2, 10.2, 11, 11.3, 12, 13, 11.1, 6.4, 6, 5.4, 6.1, 4.7, 
    4.9, 1.9, 1.8, 1.4, 4.3, 0.8, 3.9, 4.2, 2.7, 0.9, 0.9, 1.3, 0.9, 2, 0.9, 
    1.1, 1.3, 2.6, 2.4, 0.2, 0.9, 1.2, 0.8, 0.2, 1, 0.5, 1.4, 0.8, 0.9, 0.9, 
    1, 0.1, 1.1, 2.2, 0.3, 1.5, 1, 1.2, 5.2, 4, 4.2, 1.8, 1.3, 2.3, 3.9, 4.3, 
    0.9, 2.9, 2, 0.4, 0.8, 1.5, 0.3, 0.6, 0.9, 1.3, 1.3, 1.2, 1.7, 0.5, 1.7, 
    1.3, 1.1, 1.4, 1.7, 4.6, 5.4, 1.7, 2.8, 7.1, 6.5, 7, 7.7, 7.2, 6.7, 5.2, 
    3.4, 2, 1.9, 0.7, 5.2, 1.5, 2, 1.2, 1.2, 0.5, 1.5, 1.3, 0.1, 4.7, 4.2, 
    1.6, 0.1, 1.2, 1.3, 2.6, 1.4, 1.5, 0.7, 1.6, 1.3, 0.9, 10.2, 10.3, 9, 5, 
    9.2, 9, 9, 8.1, 9.8, 7.9, 10.3, 8.9, 8.1, 8.3, 7.6, 9.3, 6.5, 8.5, 5.6, 
    5.8, 5.6, 4.5, 6, 4.4, 4.9, 4.9, 4.4, 2.1, 4.3, 2.8, 2.3, 2.5, 3.3, 1.7, 
    0.8, 1.3, 0.6, 1.9, 0.4, 0.7, 0.6, 0.9, 0.7, 0.5, 0.8, 1, 0.9, 0.6, 2.1, 
    1.5, 0.5, 0.6, 1.2, 2.2, 1.8, 1.2, 0.4, 1.6, 1.3, 2.9, 3.2, 0.6, 0.9, 
    1.3, 0.3, 0.6, 1, 0.7, 0.5, 0.5, 0.9, 0.2, 0.3, 1.3, 1.9, 0.6, 1.6, 1, 
    0.8, 0.9, 0.8, 1.1, 1.1, 0.6, 0.4, 0.4, 0.3, 0.7, 0.4, 0.6, 0.5, 0.2, 
    0.5, 0.4, 0.7, 0.9, 1.5, 0.7, 1.5, 1.1, 1.1, 0.5, 0.7, 1, 0.4, 0.8, 0.9, 
    0.6, 1.5, 0.9, 1, 0.4, 0.3, 0.7, 0.1, 0.1, 0.2, 1.6, 1.2, 3.1, 4.3, 2.7, 
    4.9, 7.3, 5.5, 5.5, 4.3, 4.1, 1.2, 3, 3.2, 7.5, 8.1, 0.3, 1.4, 0.3, 2.6, 
    2.6, 2, 5.5, 7.7, 6.6, 8.2, 8.6, 6.8, 8.1, 7.9, 7, 6.3, 7.1, 5, 3.9, 4.8, 
    3.4, 1.5, 1.2, 0.9, 0.7, 1, 0.3, 1.4, 0.4, 2.2, 1.5, 0.9, 0.8, 0.9, 0.7, 
    1.8, 3.8, 2.2, 1, 0.8, 3, 2.1, 1.8, 1.3, 1.8, 2.5, 1.5, 3.1, 2.8, 1.5, 
    0.8, 2.3, 2.2, 3.6, 1.4, 1.5, 0.8, 1.4, 1.8, 0.9, 1.1, 1.8, 1.4, 0.8, 
    0.9, 1.1, 1, 0.4, 0.6, 0.6, 4.8, 5.3, 0.5, 4.5, 1.2, 1.3, 0.8, 1.1, 1.4, 
    1.4, 0.1, 1.2, 1, 0.6, 1.3, 0.5, 0.4, 0.7, 0.2, 0.4, 0.5, 1, 1, 0.4, 1.1, 
    1.3, 0.8, 0.5, 1.4, 1.2, 1.3, 1.2, 1, 0.3, 1.2, 1, 0.1, 0, 1.6, 1.5, 1.2, 
    1.1, 1.6, 0.9, 6.5, 2, 1.7, 6.7, 3.4, 1.9, 0.6, 0.6, 0.5, 1.9, 1.2, 0.5, 
    2.1, 1.6, 1.1, 0.5, 1.7, 1.3, 1.1, 1.2, 1.1, 0.8, 1.8, 0.8, 1.5, 0.8, 
    0.7, 1, 1.3, 3.6, 1.1, 3.8, 4.8, 3.7, 0.9, 1.4, 0.9, 1, 1.6, 4.2, 6.3, 
    4.7, 9.4, 5.9, 6.2, 8.2, 8.4, 9.4, 5.8, 10.8, 9, 11.2, 11.8, 11.3, 10.3, 
    9.4, 9.7, 10.5, 10.8, 11.3, 11.9, 12.3, 13.7, 14.6, 15, 15.5, 15.7, 15.9, 
    16.1, 16.9, 15.9, 17, 17.8, 19.7, 19.3, 19.2, 19.7, 19.3, 18.3, 17.7, 
    17.3, 19.8, 20, 17.6, 12.1, 3.9, 3.9, 9.4, 9.6, 12.2, 12, 11.7, 10.3, 
    11.5, 8.5, 9.3, 9.6, 10.4, 9.1, 8.3, 11.3, 11.2, 7.9, 6.2, 9, 6, 5.6, 
    6.5, 7.1, 4.7, 4.3, 5.1, 4, 7.3, 4, 5.7, 4.2, 4.3, 2.7, 4, 2.9, 5.3, 4.4, 
    5.2, 2.8, 2.7, 0.5, 1, 1.3, 0.8, 0.2, 1.3, 0.9, 0.7, 0.7, 1.7, 0.5, 1.2, 
    1.5, 0.4, 1.4, 2.1, 0.7, 1, 1.5, 1.1, 0.5, 0.8, 1.2, 1, 2.5, 2, 2.5, 1.4, 
    0.7, 0.7, 0.5, 0.6, 1.1, 0.9, 0.9, 0.6, 1.3, 1.9, 1.2, 1.2, 0.7, 0.4, 
    1.5, 0.9, 0.6, 5.8, 3.3, 4.7, 0.7, 1.4, 2, 5.8, 4.9, 4.8, 5.1, 4.9, 1.1, 
    1.2, 2.3, 2.2, 2.3, 2.2, 2.6, 0.7, 4.2, 4.3, 3.4, 2, 0.9, 1.7, 0.6, 0.4, 
    0.3, 0.5, 0, 0, 0.6, 0.9, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.6, 8.2, 
    3, 4.7, 6.9, 6.1, 5.9, 5.7, 6.8, 6.2, 8, 7.5, 6.5, 5.1, 7, 8.7, 7.9, 8.4, 
    8, 7.5, 6.6, 8.1, 8.8, 10.4, 8.7, 8.2, 9.2, 9.2, 7.9, 8.7, 7.6, 3.8, 4, 
    4.7, 4.8, 3.8, 3.1, 1.9, 3.1, 2.9, 4.2, 3.5, 4.3, 4.3, 3.8, 4.6, 4.6, 4, 
    3.5, 3.2, 6.6, 3.6, 4.1, 3.4, 2.7, 5, 5.4, 4.3, 4.6, 4.8, 4.3, 4.1, 2, 
    1.4, 0.8, 1.2, 2.5, 1, 1.5, 1.2, 1.8, 1.7, 3.1, 3.1, 6.9, 1.7, 3.4, 3.2, 
    0.4, 0.5, 1.2, 0.8, 0.6, 1.8, 0.2, 0.7, 4.3, 4.3, 5.6, 3.7, 3.5, 0.8, 
    1.5, 0.4, 0.6, 2.8, 1.1, 4.6, 3.9, 2.9, 3, 2.1, 1.9, 5.2, 1.3, 1.1, 0.1, 
    0.2, 0.5, 1.4, 0.8, 0.5, 0.6, 1.7, 2.2, 3.8, 0.8, 2.5, 5.3, 5.7, 4.7, 
    1.7, 9.3, 1.8, 1.8, 2, 5.7, 3, 4.1, 3, 4.1, 3.4, 3.4, 1.8, 0.7, 0.6, 1.6, 
    0.7, 2.2, 3, 0.9, 0.2, 1, 0.9, 0.7, 0.5, 1.6, 0.5, 2, 0.4, 0.7, 1.2, 1.2, 
    1.6, 1.3, 1.5, 3.6, 4.1, 5.5, 5.9, 5.2, 1, 5.1, 5, 4.1, 3.4, 4.6, 5.5, 
    5.6, 5.6, 3.7, 4.8, 3.5, 1.2, 0.1, 2.3, 0.7, 0.5, 0.7, 0.4, 0.2, 0.6, 
    1.3, 1.4, 2.6, 1.3, 1.6, 2.2, 3, 0.5, 1, 3.2, 1.7, 1.7, 6.7, 7, 1, 1.4, 
    1.6, 0.5, 2.8, 0.7, 1.8, 1.4, 1.3, 1.4, 1.1, 1.6, 1, 5.1, 6.1, 5.8, 6, 
    10.1, 10.7, 7.4, 6.3, 2.9, 3.3, 0.7, 1, 2.2, 1.2, 3, 1.4, 2.2, 2, 6, 2.9, 
    5.1, 3.9, 0.9, 4, 8, 10.8, 9.8, 7, 5.4, 9, 5.3, 5.4, 3.3, 4.8, 2.8, 2.8, 
    2.5, 2.4, 3, 2.8, 2, 3.1, 2.4, 3.4, 3, 2.9, 2.1, 0.4, 1.3, 1.9, 2.8, 2.3, 
    2.8, 2.4, 2.4, 3.3, 2.8, 2.7, 2.5, 0.8, 2.6, 1.6, 1.8, 1.4, 3.4, 2.5, 
    3.3, 3.5, 3, 2.5, 3.8, 2.8, 2.7, 3.7, 2.4, 2.9, 2.7, 3, 2.8, 1.8, 2.3, 2, 
    1.7, 0.7, 1, 1.6, 2.7, 1.5, 0.4, 1.3, 1.4, 0.6, 1.7, 0.6, 1, 1.9, 0.1, 
    1.1, 0.7, 0.9, 1.2, 1.3, 0.7, 2.8, 0.9, 0.3, 1.2, 0.7, 1, 0.4, 3.3, 3.4, 
    3.8, 2.7, 4.8, 3.5, 2.9, 3.9, 3.8, 4, 2.3, 3, 5.1, 2.9, 4, 3.3, 2.9, 3, 
    3.3, 2.1, 0.8, 0.9, 1, 1, 1.5, 2, 3, 5.1, 2.8, 2, 2, 3.1, 4.1, 5.9, 6.3, 
    7.4, 7.5, 6.9, 6.9, 4.2, 5.4, 5.9, 4.4, 4.6, 4.8, 5, 5.2, 5.4, 4, 3, 1.3, 
    0.8, 1.1, 1.9, 1, 4.4, 4.7, 3.9, 3.6, 2.3, 0.7, 3.3, 3.4, 4.2, 4, 3, 2.5, 
    1.7, 1.9, 1.4, 1, 1, 2.1, 1.3, 0.8, 1, 1.2, 3.6, 3.6, 3, 1, 1.7, 3.7, 
    3.3, 0.7, 1.5, 6, 4.2, 3.8, 4.3, 4.3, 5.1, 5.7, 5.8, 5.6, 5.6, 5.5, 5.9, 
    7.3, 7.5, 7.3, 7.2, 6.4, 6, 6.2, 6.1, 4.1, 5.7, 5, 3.5, 1.6, 0.9, 0.4, 
    0.4, 1.1, 1.7, 2.3, 0.9, 0.6, 0.2, 0.8, 0.2, 0.8, 0, 0.8, 0.2, 0.8, 0.3, 
    0.7, 0.1, 0.2, 0.3, 0.6, 0.1, 0.1, 0.5, 0.1, 0.1, 0.6, 0.2, 0.3, 1.1, 
    0.1, 0.7, 0.7, 0, 0.6, 0.3, 0.5, 0.5, 0, 0.6, 0.5, 0.6, 0.1, 0.6, 0.9, 0, 
    0.1, 0.9, 0.3, 0.7, 0.1, 0.8, 0.3, 0.5, 1, 0.3, 0.8, 1.2, 3.2, 5.4, 4.6, 
    5.3, 3.8, 3.8, 3, 3.5, 2.7, 2.6, 2.7, 4.1, 3.9, 3.2, 3.1, 1.3, 1, 0.4, 
    0.7, 0.8, 0.5, 0, 0, 1, 0.8, 0.9, 0.5, 0.7, 1.1, 1, 2, 0.5, 1, 0.8, 1, 
    0.9, 0.9, 1.3, 0.3, 2, 1, 0.6, 1.2, 1.6, 1, 2.1, 0.4, 1, 5.5, 2.1, 1.5, 
    0.6, 2.5, 1.6, 0.2, 1.4, 1.1, 2.2, 1.9, 2.6, 3.8, 3.4, 4, 1, 1.2, 1.6, 
    1.9, 1.5, 3.7, 1.3, 1.1, 0.6, 4, 1.7, 0.5, 1, 1.6, 1.2, 1.7, 1.6, 0.8, 
    1.9, 0.6, 1, 0.9, 1.7, 1.3, 2.3, 0.6, 0.8, 0.6, 5.1, 4, 5.6, 4.3, 2.1, 
    5.2, 4.8, 2.8, 1.3, 2.3, 1.6, 2.1, 1.2, 1.7, 3.3, 0.6, 1, 2.3, 1.7, 0.9, 
    1.4, 1, 5.7, 2.2, 0.4, 0.9, 0.6, 1.3, 0.7, 5.8, 0.7, 0.5, 2.7, 2.8, 3.1, 
    0.7, 1.2, 0.9, 0.5, 1.6, 1.3, 3.7, 0.3, 0.2, 0.3, 0.1, 0.7, 0.6, 0.9, 
    0.4, 1, 0, 0, 1.1, 0.3, 0.3, 0.6, 0.5, 0.4, 0.5, 0, 0, 0.4, 3, 1.4, 3.9, 
    3.4, 4.1, 3.5, 2.4, 1, 2.6, 0.7, 0.5, 1.5, 0.8, 1.1, 0.8, 0.3, 0.3, 1.1, 
    1.5, 1.5, 2.4, 0.3, 1.1, 0.1, 0.1, 0.5, 0.3, 0.6, 0.5, 0.8, 1.4, 0.5, 
    1.3, 0.7, 0.9, 0.3, 0.8, 0.1, 0.3, 0, 0.8, 0.5, 1, 1, 0.5, 0.4, 0.1, 0.7, 
    0.3, 0.7, 0, 0, 1.1, 2.4, 0.7, 2.1, 2, _, _, 2.5, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2.9, 2.2, 2.5, 1.1, 
    1.3, 2.4, 0.7, 1.8, 1.4, 0.7, 1.3, 1.1, 0.9, 1, 1.1, 2.1, 0.9, 8, 1, 0.8, 
    1.5, 1, 0.7, 0.5, 2, 2.5, 1.9, 0.6, 1.5, 1.6, 1.4, 1.7, 1.6, 1.1, 1.2, 
    0.3, 3.9, 6.6, 3.3, 2.8, 3.6, 3.2, 5.2, 4.5, 4, 6.3, 7.9, 7.2, 9, 9.7, 
    8.2, 9.6, 9.6, 9.5, 9.1, 9.6, 10, 11.1, 6.9, 10.6, 10.8, 9.1, 9.4, 8, 
    8.2, 7, 6.9, 8.2, 6.8, 7.5, 7.2, 5.4, 5.4, 5.8, 5.5, 6, 5.4, 6.9, 4.8, 
    4.3, 4.5, 5.4, 6.4, 5.9, 5.9, 6.1, 5.5, 5, 4.4, 5.8, 5.3, 5.9, 5.7, 5.2, 
    6.4, 6, 5.3, 4.8, 6.3, 3.8, 5.6, 4.8, 4.4, 4.4, 4.5, 6.8, 4, 4.7, 5.8, 
    3.3, 5.5, 4.8, 6.1, 4.2, 3.6, 4.2, 1.2, 5, 4.9, 7, 6.4, 3.9, 1.1, 1.3, 
    0.9, 0.8, 0.2, 0.5, 0.4, 0.3, 0.8, 0.3, 0.5, 0.5, 1.1, 1.5, 0.4, 0.6, 
    1.1, 1.6, 2.2, 5.3, 4.8, 4.3, 5.5, 8, 7, 8.1, 6.9, 7.4, 7.7, 5.5, 7.1, 
    8.4, 5.6, 7.1, 8.3, 7.6, 7.1, 6.7, 6.6, 5.5, 6.9, 8.5, 8.7, 3.9, 2.9, 
    3.8, 4.9, 2.6, 1.9, 3.6, 3.5, 4.3, 1.8, 2.7, 2.9, 1.9, 2.7, 2.3, 4.3, 
    3.3, 1.9, 2.7, 2.3, 2.5, 2.4, 2.6, 5.6, 5.4, 2.3, 5.3, 5.3, 4, 6.6, 4.9, 
    5.7, 6.3, 5.8, 5.5, 5.1, 7, 5.8, 4.8, 4.7, 5.2, 6.7, 8.2, 10.1, 6.3, 5.3, 
    8, 7.5, 7.9, 6.8, 5.4, 2.7, 1.4, 4.9, 7, 3.8, 6.5, 5.6, 9.4, 5, 7.4, 8.6, 
    3.6, 4.3, 8.5, 6, 5.2, 7.9, 6.6, 7.2, 7.7, 6.4, 6.6, 7.5, 3.7, 4.8, 7.4, 
    3.1, 5.3, 3.7, 7.7, 5.1, 6.4, 4.8, 6.6, 3.8, 2.9, 4.7, 6.1, 5, 2.9, 4.4, 
    4.2, 1.2, 4.2, 3.9, 6.4, 4.1, 5.3, 5.3, 4.4, 3.7, 6.2, 4.9, 6.5, 5, 2.8, 
    3.6, 1.5, 3.2, 0.7, 1.1, 1.2, 3.4, 1.5, 0.2, 1.1, 0.6, 2.7, 0.8, 0.7, 
    0.5, 0.9, 0.7, 0.6, 0.6, 0.1, 1.4, 1.4, 0.3, 0.7, 0.5, 1, 0.7, 0.2, 1, 
    0.5, 0.4, 0.9, 1, 2, 2.1, 0.8, 0.7, 1.1, 0.8, 0.2, 0.6, 0.3, 0.9, 0.9, 
    1.1, 1, 1.4, 1.2, 0.8, 1.5, 0.4, 0.7, 0.3, 1.8, 0.3, 0, 1.5, 0.1, 0.7, 
    0.7, 0.5, 1.1, 0.3, 0.9, 1, 0.4, 1.8, 0.9, 0.6, 0.7, 0.5, 0.8, 0.8, 0.4, 
    1.4, 1.1, 2.2, 0.7, 0.7, 0.4, 1.9, 0.8, 1.9, 3.6, 2.8, 0.6, 0.8, 2, 2.7, 
    2.6, 2.5, 3.2, 4.1, 3.9, 3, 1.2, 0.8, 0.3, 1.7, 3.6, 1.9, 0.6, 4.8, 3.4, 
    7.6, 8.1, 8, 7.8, 8.3, 9.9, 10.2, 12.3, 9.2, 8.7, 8.2, 6.6, 7.7, 4.9, 
    3.2, 2.4, 2.4, 1.2, 3.9, 2.9, 2.6, 8.7, 4.4, 4, 6.2, 3.6, 3, 2.4, 2.5, 
    3.7, 2.4, 3, 1.8, 2.2, 1.4, 2.9, 1.5, 1.7, 1, 0.2, 0.5, 2.8, 2, 2.2, 3.1, 
    1.9, 1.6, 2.4, 2.7, 1.8, 2, 1.2, 1, 1.1, 0.8, 0.1, 0.4, 0.1, 0.4, 0.1, 
    0.1, 1, 0.2, 1.2, 0.2, 0.1, 0, 0.1, 0.6, 0, 0.3, 0.8, 0.8, 1, 1.3, 0.5, 
    0.8, 4, 3.5, 3, 4.1, 3.2, 4.4, 3.3, 2.4, 3, 2.9, 0.4, 0.9, 0.5, 0.5, 0.9, 
    0.4, 3.8, 0.7, 1, 1.1, 0.3, 0.6, 0.6, 2.3, 2.6, 0.7, 2.2, 2, 2, 0.7, 1, 
    0.6, 0.1, 0.3, 0.7, 1.8, 0.8, 0.4, 1.4, 1.9, 1.1, 0.9, 0.3, 0.7, 0.3, 0, 
    0.2, 0.8, 1.8, 0.6, 0.6, 1.5, 0.5, 0.7, 1.4, 2, 2.8, 3.3, 3.5, 5.5, 6.6, 
    4.7, 5.5, 4.2, 7.3, 6.2, 4.8, 8.4, 6.6, 7.7, 9.7, 10.4, 8.7, 8.5, 8.3, 6, 
    5.5, 6.1, 4.6, 5.3, 0.7, 0.8, 0.3, 1.3, 1.1, 0.8, 3.3, 1.8, 4.6, 0.7, 
    1.3, 2.6, 2.8, 3.4, 3, 0.9, 1.3, 0.9, 0.1, 0, 0, 0.1, 0.9, 1.2, 0.4, 1.3, 
    0.2, 1.5, 1.9, 0.3, 0.4, 2, 1.6, 0.6, 0.8, 0.5, 0.4, 1.4, 0.5, 1.2, 0.2, 
    0.5, 0.9, 0.2, 0.3, 1, 5.5, 5.9, 4, 3.4, 5.7, 8.1, 6.3, 7.7, 5.8, 6.5, 6, 
    7.3, 6.2, 6.1, 5.3, 3.3, 3.3, 0.6, 0.7, 1.6, 1.3, 1.2, 1.1, 1, 1.4, 0.5, 
    0.8, 0.6, 2.3, 1.5, 1, 0.4, 1, 0.8, 5.4, 2.2, 1.2, 1.3, 0.3, 1, 1.4, 1.4, 
    0.7, 1.3, 1.3, 1.8, 0.2, 0.3, 0.4, 0.6, 0.8, 0.3, 0.5, 0.4, 0.2, 0.4, 
    0.2, 0.6, 0.3, 0.2, 0.3, 1, 0.6, 0.1, 0.5, 1.3, 0.5, 0.4, 0.6, 0.7, 2, 
    1.1, 1.8, 1.3, 0.4, 0.8, 0.3, 0.2, 0.9, 1.1, 0.5, 0.9, 0.9, 0.5, 1.2, 
    0.2, 2.1, 1.8, 0.4, 1.5, 0.7, 1, 0.3, 0.8, 1.9, 0.4, 0.7, 1.3, 1, 1.4, 
    1.9, 5.2, 5.2, 5, 9.5, 6.8, 4.6, 7.5, 4.3, 7.3, 6.5, 5.8, 8.4, 7.2, 5.3, 
    4.2, 5.6, 4.7, 5.1, 6.9, 7.2, 7.3, 4.2, 3.6, 5.9, 6.3, 3.9, 3.5, 1.9, 
    1.4, 1, 1, 1.2, 0.8, 1.6, 0.8, 1.1, 1.1, 1, 0.2, 0.4, 1.5, 2.7, 1.8, 2.2, 
    6.5, 6, 3, 2.3, 2.1, 4.1, 5.8, 6.6, 4.5, 3.1, 3.1, 4.4, 4.6, 2.5, 2.6, 
    4.6, 5.5, 4.6, 4.8, 3.4, 4, 4.7, 4.5, 3.5, 3.7, 5, 4.7, 1.8, 3.7, 2.5, 
    0.9, 1.2, 1.5, 0.6, 1.5, 1.1, 0.1, 0.8, 0.6, 0.2, 1.2, 1, 0.2, 0.1, 0.4, 
    0.7, 0.5, 2.7, 0.5, 1.3, 0.5, 0.8, 1.2, 2.1, 2.2, 1.3, 0.6, 0.5, 0.9, 
    1.4, 1.6, 1, 0.2, 0.7, 0.8, 1.6, 1.5, 1.3, 0.1, 2.7, 1.3, 0.9, 0.8, 0.5, 
    1.5, 1.6, 2.8, 1.1, 1.4, 1.2, 1, 0.4, 1, 0.7, 0.1, 0.7, 1.3, 0.7, 0.8, 
    1.7, 0.5, 0, 1, 0.9, 0.4, 0.9, 0.6, 0.2, 1.1, 0.3, 0.4, 1, 0.7, 1, 0.2, 
    0.8, 0.1, 0.3, 0.9, 0, 0.1, 0.2, 0.5, 0.3, 0.5, 0.4, 1, 0.7, 0.3, 0.1, 
    0.4, 0.2, 0.1, 0.3, 0.3, 0.9, 0.3, 0.6, 0.6, 1.3, 1, 0.2, 0.8, 0.2, 0.1, 
    0.9, 0.3, 0.1, 1.2, 0.3, 0.2, 0.9, 0.2, 0.1, 0.3, 0.4, 0.2, 1, 0.6, 0.4, 
    0, 1.5, 1, 0.4, 0.6, 0.1, 0.7, 0.5, 0.6, 0.7, 1.3, 1.3, 2.4, 0.6, 0.9, 
    0.3, 0.8, 0.1, 1.5, 1.8, 0.8, 0.4, 0.5, 0.4, 0.7, 0.7, 0.5, 0.1, 0.3, 
    0.6, 0.5, 0.7, 3.9, 4.6, 4.4, 4.9, 5.9, 4.5, 2.3, 2.3, 0.6, 2.1, 0.9, 1, 
    0.1, 1.1, 0.5, 0.7, 1.4, 0.4, 7.4, 4, 4, 5.2, 5.2, 6.1, 4.2, 4.4, 3.7, 
    3.6, 4.1, 3.4, 4.6, 6.8, 6.1, 3, 3.9, 3, 1.2, 1.8, 0.2, 1.3, 0.2, 1, 0.4, 
    2.2, 0.9, 1, 3.6, 1.7, 3.4, 0.7, 2, 0.9, 2.5, 0.9, 0.5, 0.7, 0.7, 4.6, 
    4.7, 3.8, 0.8, 0.8, 3, 4.5, 1.9, 1.4, 0.3, 0.1, 0.8, 0.1, 0, 1.2, 0.3, 0, 
    0.3, 0, 0.4, 0, 0.8, 0.8, 0.2, 0.8, 0.2, 0.6, 0.3, 1.2, 1.8, 0.4, 0.7, 
    1.3, 5.3, 4.9, 4.9, 4.3, 3.5, 4.4, 3.3, 3.2, 2.1, 1.3, 0.5, 0.4, 3.1, 
    2.2, 2.7, 3.1, 0.7, 1.4, 0, 0.1, 0, 0.7, 0.5, 0.2, 0.2, 0.1, 0.9, 1.1, 
    0.7, 0.6, 1.7, 0.7, 0.4, 0.1, 0.4, 0.9, 0.2, 0.3, 0.5, 0, 0.3, 1.2, 1, 1, 
    1.8, 0.6, 0.1, 0.3, 0.2, 0.7, 0.1, 1.2, 0.1, 0.4, 0.6, 0.3, 0.3, 0.6, 
    0.1, 0.7, 0.7, 0.7, 0.2, 0.7, 0.5, 1, 0.1, 0.9, 0.7, 0.2, 0.4, 0.4, 1.3, 
    0.3, 1.3, 1.1, 0.2, 0.9, 0.7, 0.4, 0.2, 0.1, 0, 0.7, 0.9, 1.2, 1.3, 1.1, 
    0.5, 0.6, 0.8, 0.7, 1.2, 1.6, 0, 0.5, 0.2, 0.4, 0.6, 1.5, 1, 0.9, 0.3, 
    0.4, 2.3, 0.3, 0.5, 0.8, 0.2, 0.3, 0, 1.1, 0.4, 0.2, 0.3, 0.2, 0.7, 1, 
    0.8, 1.2, 0.3, 1.2, 0.4, 0.7, 1.2, 1, 2, 0.2, 0.9, 0.7, 0.3, 0.3, 1, 0.2, 
    1.1, 0.5, 2.2, 1.9, 1.6, 0.1, 0.9, 2.1, 2, 1, 5.7, 1.6, 2, 1.5, 1.4, 2.6, 
    1.7, 1.6, 4.2, 3.9, 3.2, 3.7, 2.8, 0.1, 0.8, 2.8, 3.1, 4.2, 5.9, 6.2, 
    7.9, 3.7, 7.4, 7.5, 7, 6.7, 5.4, 3.3, 4.1, 8.5, 2.3, 5.3, 3.4, 3, 1.7, 
    0.2, 0.9, 0.8, 1.9, 3.5, 3.1, 5.4, 6.1, 7.3, 9, 8.6, 7.2, 3.7, 7.5, 7.5, 
    5.3, 8, 7.5, 4.3, 9.4, 6.8, 5.9, 4.2, 4.4, 4, 3.7, 2.9, 1.7, 0.4, 1.2, 
    1.2, 0.9, 1, 2, 0.7, 2.3, 2.3, 1.6, 2, 1.8, 2.1, 1.2, 1.2, 2.3, 0.7, 0.5, 
    0.8, 1.5, 2.9, 2.3, 3.4, 7.8, 6.5, 6.5, 3.3, 6.1, 8.7, 8.5, 7.5, 8.1, 
    7.9, 7.2, 2.4, 1.5, 3.8, 1.5, 0.1, 1.2, 1.3, 3.2, 5, 0.5, 5.6, 7.7, 6.3, 
    6.8, 4.9, 5.1, 1.4, 3.5, 2.1, 5.4, 3.6, 1.2, 3.5, 3.2, 1.5, 3.5, 2.5, 
    1.3, 7.1, 2.5, 2.5, 0.8, 1.8, 0.7, 1.6, 1.6, 2.1, 2.1, 2.8, 2.2, 2.2, 
    1.6, 2.8, 3.2, 3.3, 4.9, 4.6, 7.2, 6.9, 2.1, 6.2, 6.5, 2.3, 3.6, 3.6, 4, 
    4.3, 5.5, 3.5, 2.5, 1.7, 2.1, 6.3, 8.6, 2.4, 2.7, 2.5, 4.3, 3.9, 4.2, 
    4.9, 6.2, 2.8, 0.9, 3, 2, 1.3, 1.3, 2.4, 0.7, 0.8, 1.3, 2.4, 1.4, 1.4, 
    1.2, 2.2, 3.1, 1.4, 4.2, 3, 2.2, 3, 4, 1.1, 1, 2.5, 1.2, 1.6, 3.1, 4, 
    0.6, 1.2, 0.7, 2.4, 1.3, 1.1, 2.5, 1.2, 1, 0.8, 0.9, 1.3, 1.6, 0.5, 1, 
    0.8, 0.8, 1, 1.9, 0.2, 2.4, 2.4, 1.9, 2.1, 1.4, 3.1, 1.4, 0.7, 1.9, 2.2, 
    1.5, 0.7, 1.4, 0.7, 1.8, 2.2, 2.7, 1.4, 0.9, 1.4, 1, 0.4, 3.4, 0.8, 0.4, 
    0.5, 0.8, 0.1, 0.5, 0.5, 0.3, 0.3, 0.7, 1.2, 1, 1.5, 1.4, 1.1, 0.3, 0.5, 
    0.9, 0.6, 0.1, 1.3, 1.1, 1.2, 1, 0.9, 1.6, 0.4, 0.6, 1.2, 0.3, 1.9, 0.4, 
    1, 1.6, 0.9, 1.7, 0.7, 2, 0.8, 0.4, 0.3, 2.6, 0.6, 0.4, 0.7, 1.1, 0.3, 
    1.8, 0.4, 0, 0.8, 0.6, 1, 0, 0.8, 0.6, 0.7, 0.2, 0.8, 0.2, 0.8, 0.6, 0.4, 
    1, 0.6, 0.3, 1.1, 0.2, 1.4, 0, 0.6, 0.6, 0.2, 0.2, 0.3, 0.5, 0.3, 0.1, 
    0.1, 0.2, 0.6, 0.9, 0.1, 0.4, 0.6, 0.1, 0.5, 0.9, 0.1, 0.5, 0.3, 1, 1.6, 
    0.7, 0.8, 0.2, 0.7, 0.7, 0.3, 0.9, 0.3, 0.3, 0.4, 1.7, 0.6, 0.7, 1, 0.3, 
    1, 0.8, 1.4, 0.8, 0.9, 2, 1.4, 1.7, 0.7, 1.5, 1, 1.4, 1, 1.8, 1.7, 0.6, 
    1.3, 0.9, 1.4, 0.8, 1.8, 1.1, 5.6, 6.2, 7.9, 7.9, 8.8, 9.2, 8.1, 7, 7.1, 
    7, 4.6, 5.3, 1.7, 7.5, 7.5, 3.9, 3.1, 3.7, 0.8, 0.7, 0.9, 1, 3.6, 4.8, 
    5.4, 3.3, 5.8, 6.7, 5.8, 5.2, 5.4, 6.4, 6.1, 2.9, 1.4, 1.7, 0.9, 1.3, 
    0.9, 5.7, 5, 6, 6.6, 5.4, 6.1, 6, 3.9, 3.9, 4, 4.7, 3.1, 2.2, 2.4, 2.7, 
    0.4, 0.7, 0.2, 0, 0.2, 0.7, 0.8, 1.4, 0.4, 0.5, 0.6, 0.3, 0.8, 0.7, 1.7, 
    0.1, 0.5, 1, 1.4, 0.7, 0.2, 0.4, 0.6, 1, 0.3, 0.5, 0.7, 0.4, 1.9, 3.9, 
    4.4, 2, 2.6, 5.5, 5.3, 6.2, 5.8, 5.6, 5.8, 6.6, 6.8, 8.1, 6.6, 5.1, 5.9, 
    6.2, 5.6, 5.8, 5.6, 6.3, 7, 7.7, 8.5, 6.7, 6.4, 6.4, 6.1, 2.3, 3.8, 1.3, 
    1.3, 2.9, 1.3, 1.5, 2.3, 0.5, 0.1, 0.8, 0.2, 0.2, 1.1, 1, 0.7, 1.3, 0.2, 
    0.7, 0.7, 0.5, 1.5, 0.4, 0.5, 0.1, 0.7, 1.2, 0.2, 0.4, 0.5, 0.8, 0.4, 
    0.6, 0.3, 0.5, 0.7, 1.4, 0.2, 1, 1, 0.5, 0.7, 0.1, 0.2, 0.2, 2, 2.9, 2.3, 
    0.2, 0.3, 0.6, 0, 0.3, 0.3, 0.2, 0.7, 0.4, 0.2, 0.3, 0.1, 0, 0.1, 0.8, 
    2.2, 2.7, 2.6, 3.2, 3.8, 2.2, 1.8, 2.7, 2.5, 0.6, 2.9, 2.9, 1.1, 0.1, 1, 
    2.3, 3.7, 4, 3.6, 3.2, 3, 3.3, 2.6, 2.8, 4.2, 2.7, 2.6, 2.4, 1.2, 2.3, 
    1.8, 2.5, 2.7, 2.5, 1.7, 1.7, 1.5, 1.9, 0.1, 0, 0.9, 0.4, 1.8, 3.1, 3.5, 
    2.8, 2.8, 3, 2.4, 0.9, 0.9, 0.3, 0.9, 1.6, 1.1, 1.9, 1.9, 0.3, 2.2, 1.3, 
    2.3, 0.9, 0.7, 0.1, 0.4, 0.4, 0.2, 0.2, 0.3, 0.2, 0.7, 0.8, 0.9, 0.9, 
    0.4, _, 0.9, 1.6, 0.7, 0.8, 0.2, 0, 1.1, 0.6, 1.2, 0.1, 0.1, 0.1, 1, 0, 
    0, 0, 0.2, 0, 0.5, 0, 0, 0.1, 1.5, 0.8, 0, 0, 0, 0.2, 0.2, 0.2, 1.5, 0, 
    0, 0.8, 0.1, 0.4, 0, 0.2, 0.3, 0.4, 0.1, 0.1, 0, 0, 0.4, 1, 0.5, 0.8, 0, 
    1.2, 0.8, 3.1, 3.1, 0.4, 0.3, 0.2, 0.2, 0.1, 0.1, 0.9, 2.3, 1.3, 0.5, 
    0.1, 0.3, 0, 0.1, 0.5, 1.2, 2, 0.5, 4.6, 2.3, 5.9, 5.4, 5.4, 5.9, 3.5, 
    1.2, 4.1, 2.9, 4, 1, 1.3, 4.6, 4.7, 4.1, 5.4, 3.7, 5.7, 5.3, 3, 5.4, 2, 
    3.4, 5.9, 8.1, 4, 6.5, 2.6, 1.2, 1, 1.2, 6.8, 2.1, 2, 1.7, 1.1, 1.9, 1.9, 
    4.4, 0.5, 3, 5.2, 3.4, 1.8, 4.5, 3.9, 1.6, 1.1, 2.4, 0.8, 4.3, 6.1, 6.5, 
    5.9, 6.7, 3.1, 3.6, 3.6, 1.2, 2.6, 2.2, 1.8, 1.3, 0.9, 1.4, 2.4, 1.3, 
    1.1, 2.4, 0.5, 1, 6, 0.6, 6.5, 6.3, 5.7, 2.7, 1.8, 0.9, 2.3, 1.6, 2, 1.5, 
    5.6, 1.2, 0.9, 0.6, 1.3, 1.8, 1.1, 2.8, 1.2, 1.1, 0.8, 2.1, 2, 1, 0.5, 
    0.4, 0.7, 0.5, 1.2, 0.8, 0.8, 0.2, 0.6, 0.8, 1, 0.8, 1.6, 0.8, 2.6, 2.9, 
    2.3, 3.4, 2.7, 7, 4.7, 3.5, 5.1, 5.1, 4.7, 5, 3.9, 4.3, 7.8, 8.1, 6.4, 2, 
    3, 2.7, 1.2, 2.6, 2.3, 2.1, 3.8, 6.2, 6, 1.9, 6.2, 7.2, 4.6, 3.4, 1, 2.6, 
    1.4, 4.1, 4.2, 4.3, 3.4, 2.9, 1.5, 1.6, 2.2, 1, 0.8, 1.2, 0.8, 0.9, 2.3, 
    0.9, 1, 1.1, 1.3, 0.5, 2, 0.5, 1.6, 1.8, 2, 3.6, 1.1, 1.4, 0.4, 1, 1.6, 
    1.8, 1.2, 1.3, 1.1, 2, 1.2, 3.9, 1.7, 1.9, 2, 2.3, 2.1, 2.6, 2.3, 2.5, 
    4.9, 6.4, 5.9, 6.2, 1.6, 2.1, 6, 7.7, 5.5, 6.2, 5.6, 4, 2.9, 3.5, 1.3, 
    2.6, 2, 1.2, 1.8, 1, 2, 1.7, 2.7, 2.7, 4, 2.5, 2, 2.9, 2.2, 1.3, 0.8, 
    0.7, 0.8, 0.4, 0.6, 1.2, 0.8, 0.5, 0.8, 1.1, 1, 0.1, 0.7, 0.4, 2, 1.7, 
    2.1, 3.8, 2.6, 1.4, 1.4, 1.8, 0.9, 0.6, 0.3, 0.1, 1.3, 0.4, 1, 0.4, 0.4, 
    0.5, 0.8, 0, 0.7, 0.1, 3.1, 0.3, 0.3, 1, 1.2, 0.9, 0.8, 1.3, 1.3, 0.2, 
    1.1, 1.7, 0.5, 0.1, 1.2, 0.4, 0.1, 0.2, 0.3, 0.7, 0.8, 0.5, 0.6, 0.2, 
    0.1, 1.8, 1.9, 1.7, 2, 1.3, 1.3, 1.2, 2.3, 1.1, 0.4, 0.2, 1.6, 1.4, 1.1, 
    1.1, 1.1, 1.1, 0.4, 0.3, 1.6, 0.7, 0.7, 0.4, 1.3, 0.4, 0.3, 0.1, 1, 1.1, 
    0.7, 1.3, 1, 0.2, 0, 1, 1, 0.7, 0.2, 0.9, 0.1, 0, 0.4, 0.5, 0.1, 0.5, 
    0.5, 0.1, 0.5, 0, 0, 1.5, 2, 1.9, 0.6, 0.3, 0.6, 1.3, 0.9, 1, 1, 1.2, 
    0.5, 0.6, 0.8, 6.3, 6.5, 8.6, 6.6, 3.8, 1, 2.1, 1.8, 1.7, 0.6, 0.8, 0.9, 
    1.3, 0.7, 1.6, 0.9, 1, 0.9, 0.5, 1.2, 0.7, 2.1, 0.9, 1.1, 1.2, 0.5, 0.6, 
    0.1, 0.6, 0.4, 0.5, 0.9, 1.2, 1.4, 1.4, 0.9, 1.6, 0.5, 0.5, 0.7, 0, 0, 
    0.4, 0.3, 1, 0, 0, 0, 1.1, 0.4, 0.3, 1, 0.4, 0.7, 0, 2.7, 1.1, 0.3, 1.8, 
    2.2, 1.3, 1.7, 2.1, 1.1, 1.3, 5.1, 2.4, 0.6, 5.7, 5.2, 5.3, 5.8, 6.4, 
    4.4, 1.6, 1.8, 1.5, 0.8, 1.3, 0.2, 1.2, 1.1, 2.7, 1.3, 1, 2.7, 3.4, 4.3, 
    2.6, 0.9, 0.5, 1.3, 0.8, 0.7, 0.5, 0.9, 0.7, 0.8, 0.6, 0.2, 0.5, 0.1, 0, 
    0, 0.1, 0.7, 0.5, 0.8, 2.1, 1, 0.7, 0.9, 0.4, 0, 0.1, 0.6, 0.5, 0.7, 0.5, 
    1.3, 0.4, 0.2, 0.4, 1, 1.5, 0, 0.9, 1.4, 0.6, 0.8, 1.2, 0.9, 0.1, 0.2, 
    2.5, 2.6, 0.1, 0.1, 1.6, 0.3, 0.2, 0.3, 0.6, 1.3, 0, 0.8, 0.6, 0.6, 0.3, 
    0.3, 0.4, 0.2, 0.6, 0.2, 0.4, 0.2, 0.8, 0, 0, 0.6, 0.1, 0.7, 0, 0.6, 0, 
    0.2, 0.3, 0.1, 0, 0.1, 0.2, 0.5, 2.3, 1.2, 0.3, 0.5, 0.3, 0.9, 0.5, 0.2, 
    0.3, 1.9, 2.3, 2.4, 1.4, 1, 0.5, 0.7, 1.6, 0.7, 0.4, 1.6, 0.9, 1.1, 0.3, 
    0.4, 0.3, 0, 0.2, 1.3, 0.3, 1.5, 1.1, 0.4, 0.5, 0.2, 0.4, 0.9, 0.4, 1.5, 
    3.2, 0, 0.2, 0, 0, 0, 0.5, 0.8, 0.4, 0.2, 0.2, 0.9, 0.4, 0.9, 3.4, 1, 
    0.9, 1, 1.1, 0.9, 1.1, 1.7, 2, 0.8, 1.4, 1.4, 0.9, 2.1, 1.6, 1, 0.4, 0.3, 
    0.5, 1.2, 1, 0.9, 0.7, 1, 1.1, 0.9, 0.3, 1.2, 3.5, 0.9, 0.7, 0.8, 0.5, 
    0.4, 0.8, 0.5, 4.4, 4.5, 4.3, 2.7, 3.6, 5, 3.7, 3.6, 3.8, 3.7, 4.9, 4.3, 
    5.3, 4.7, 5.6, 8.1, 9.5, 8.8, 7.7, 6.9, 6.9, 7.1, 5.5, 6.4, 5.6, 3.9, 
    3.3, 4.2, 3.3, 2, 2.4, 1.9, 1.9, 1.3, 1.3, 1.5, 5.1, 0.9, 0.7, 2, 4.3, 
    4.7, 6.1, 5.9, 5, 4.1, 2.9, 3.1, 2.9, 4.6, 4.2, 2.6, 4.4, 4.2, 4.6, 5.3, 
    4.7, 5.4, 3.9, 5.1, 3.4, 4.6, 5.3, 5.2, 4.6, 4.6, 5.1, 4.5, 4.3, 4.6, 
    4.6, 5, 5.1, 4, 4.9, 4.4, 3.5, 3.3, 1.5, 0.8, 2, 1.7, 1.3, 1.1, 2, 4.8, 
    5.1, 3.6, 0.8, 2.4, 2.9, 2.6, 1.5, 2.5, 2.2, 0.8, 1.2, 1.2, 0.2, 0, 0.2, 
    0.2, 0.1, 0.2, 0.6, 1.5, 0.3, 1.4, 2, 1.4, 0.3, 0.8, 0, 0.5, 0.2, 0.8, 
    0.4, 0.4, 0.2, 0.1, 0.7, 2.9, 1.7, 2.3, 1.3, 1, 1.1, 1.2, 2.1, 0.7, 1, 
    1.7, 2.3, 2.3, 2.3, 2.1, 2.4, 1.6, 0.9, 0.6, 1.3, 2.8, 0.3, 0.3, 0.8, 
    0.5, 0.4, 0.3, 0.8, 0.9, 2.1, 2.6, 5.3, 6.6, 5.7, 6.5, 7.4, 8.5, 7.6, 
    8.1, 7.4, 8.2, 7.9, 6.8, 6.8, 9.9, 10, 9.3, 7.7, 9.2, 10.3, 12.6, 11.7, 
    12.4, 9.1, 10.6, 10.3, 5.2, 5.9, 5, 4.9, 4.9, 6, 5.7, 5.9, 5.6, 6.2, 6.5, 
    5.2, 5.5, 6.7, 6.4, 7.1, 7.5, 7.7, 7.6, 7.2, 7.5, 7, 7.7, 7.9, 7.5, 7.1, 
    7.9, 8.4, 8.4, 7.8, 7.9, 7.3, 7.3, 7.1, 7, 5.9, 5.7, 5.9, 5.3, 6.4, 6, 
    6.5, 5.4, 4.7, 4.9, 3.5, 2.5, 2, 3, 4.1, 3.2, 5.7, 3, 3.4, 3.5, 4.9, 4.9, 
    1.2, 2.9, 6.1, 5.1, 4.3, 1.1, 6.2, 3, 4.1, 4.1, 4.2, 3, 4.4, 3.3, 0.7, 
    0.9, 1.7, 1.3, 3.4, 0.8, 1.4, 0.6, 0.7, 0.7, 1.4, 1, 0.7, 1.6, 1.5, 0.8, 
    2.1, 3.3, 2.8, 2.6, 1.9, 3.6, 3.6, 2.7, 4, 3.8, 3.4, 1.9, 4.1, 4, 2.2, 
    2.3, 3.6, 3.3, 2.9, 3.8, 2.4, 1.5, 3.2, 1.2, 0.2, 0.3, 0.2, 0.1, 0.5, 
    0.4, 0, 2.8, 2.6, 0.4, 7, 8.7, 8.8, 7.6, 6.4, 4.6, 3.9, 3.2, 5, 2.3, 1.9, 
    4.5, 5.4, 6, 5.2, 4.4, 4.5, 4.6, 6.5, 1.9, 5.9, 4.7, 6.3, 3.8, 4.2, 5.5, 
    5.3, 6.5, 5.4, 3.5, 3.6, 5.8, 2.3, 4.4, 3.3, 3.7, 3.5, 6.9, 3.9, 4.4, 
    5.7, 6, 6.2, 3.4, 4.5, 4.8, 3.8, 2.9, 1.8, 1.1, 1.7, 1.3, 1.9, 1.6, 2.3, 
    2.2, 2.4, 0.9, 1, 0.5, 1.7, 0.5, 1.5, 1.4, 0.2, 0, 0.1, 0.3, 0.1, 0.5, 
    0.7, 0.5, 0.8, 0.2, 0.8, 0.9, 2.3, 2.8, 1.3, 1.8, 2.2, 2, 1.4, 1.7, 1.3, 
    1.8, 0.8, 0.6, 1.5, 0.1, 0.7, 0.4, 1.4, 1.9, 1.5, 0.7, 1.2, 0.7, 0.9, 
    4.8, 5.7, 4.7, 5.2, 4.7, 5.5, 3.7, 4.2, 4.8, 3.6, 4, 3.6, 3.6, 4.9, 5.3, 
    4.5, 3.5, 3.1, 2.9, 2.8, 2.6, 2.3, 1.7, 1.8, 1.8, 1.3, 1.7, 1.7, 1, 1.8, 
    2.3, 1.6, 1.9, 2.4, 1.7, 1, 0.2, 0, 1.2, 1.1, 0.4, 0.6, 0.7, 1, 0.5, 1, 
    2.3, 1, 1.3, 0.9, 0.9, 1.4, 1.3, 1.3, 0.2, 0.4, 0.8, 0.6, 0, 0.3, 0, 0.2, 
    0.1, 0.4, 0, 0.5, 1.1, 0.2, 0.6, 0.7, 0.6, 0.9, 0.9, 1.1, 1, 0.9, 1.3, 
    2.3, 2.7, 1.5, 2.5, 0.8, 1.1, 1.7, 2.7, 1.1, 1.5, 0.7, 0.7, 1.6, 4, 3.7, 
    3.7, 3.6, 2.9, 2.1, 1, 1.8, 2.2, 2.5, 2.6, 2.6, 2.1, 1.3, 1.1, 2.2, 2, 
    2.7, 2.1, 1.6, 0.8, 2.2, 1.4, 1, 0.4, 2.4, 1.9, 2.3, 1.8, 2, 1.9, 2, 1.6, 
    1.3, 0.9, 0.8, 0.4, 0.7, 0.2, 1.2, 0.1, 0.2, 0.7, 0.1, 0.9, 0.9, 0.6, 
    1.5, 1.4, 2.5, 1.7, 2, 1.7, 1.3, 2.1, 1.6, 5.4, 6.8, 7.8, 6.7, 4.6, 6.5, 
    5.3, 5.4, 7.1, 6.3, 7.7, 5.2, 4.1, 5.3, 6.1, 6, 5.3, 5.7, 7.1, 7.4, 5.3, 
    5.1, 4.9, 5.5, 4.7, 5.2, 5.8, 6.2, 5.2, 5.6, 4.7, 5.2, 3.8, 2.6, 1.1, 
    1.6, 1, 1.9, 0.9, 1.4, 1.6, 0.3, 2.1, 1.3, 1.2, 1.2, 1.4, 1.3, 1.7, 1.7, 
    1.6, 2.6, 2.1, 1.7, 2.5, 1.4, 1.1, 1.1, 0.6, 0.2, 0.6, 1.5, 2, 1.5, 1.9, 
    1.5, 1.2, 2.3, 1.2, 1.4, 1.8, 2, 2, 2.4, 2.7, 2.5, 2.8, 1.5, 2.2, 2, 0.5, 
    0.4, 0.4, 0.2, 0.6, 0.6, 0.6, 0.6, 1.5, 1.6, 1.1, 2.6, 1.7, 1.2, 1.2, 
    0.4, 1, 1.6, 1.7, 1, 0.6, 0.9, 0.8, 0.4, 0.7, 1.3, 0.4, 1.5, 0.9, 1.9, 
    1.2, 1.4, 0.9, 1, 1.1, 1.2, 2, 1.8, 1.2, 1.2, 4.1, 1.9, 3.5, 2.6, 2, 1, 
    1.4, 1.1, 0.9, 1.7, 2.9, 0.9, 1.5, 1.5, 0.2, 1.9, 1.3, 2.5, 1.7, 2.5, 1, 
    2.1, 1.7, 2.1, 1.6, 1.9, 4.4, 5.6, 5.2, 6, 4.9, 5.5, 2.6, 4.7, 2.8, 3.6, 
    3.5, 6, 3.9, 5.6, 3.6, 1.6, 1, 2.5, 8.4, 3.7, 4.2, 2.5, 3.6, 5.5, 2.2, 2, 
    6.9, 5.7, 6.2, 4.5, 3.5, 6.8, 3.5, 5.1, 4.9, 4.1, 4.3, 2.1, 1.8, 5.3, 3, 
    1.3, 3.6, 3.9, 2.2, 2.9, 5, 6.2, 4.6, 5.2, 5.2, 7, 4.2, 5.7, 4.9, 3.2, 
    1.7, 1.1, 0.7, 0.9, 2.5, 2.4, 1.9, 3.8, 5, 4.1, 5.2, 5.2, 5.1, 4.7, 4.4, 
    4.1, 4.2, 3.7, 4.3, 3.9, 4.1, 3.8, 3.1, 3.4, 2.7, 2.5, 0.7, 0.9, 1.1, 
    0.9, 1.4, 2, 2.2, 3.5, 2.4, 5.2, 2.2, 4.5, 4.4, 3.5, 3.5, 2.5, 2.7, 3.2, 
    3.5, 2.1, 1.6, 3.7, 2.2, 4.3, 0.5, 2.2, 0.4, 0.6, 3.3, 1.7, 1.5, 2.1, 2, 
    3.4, 3.2, 2, 3.6, 3.7, 3.4, 1, 1.7, 3.4, 1.3, 3, 1.8, 2.2, 3.2, 0.8, 0.9, 
    0.8, 1.2, 0.3, 3.1, 2.6, 2.4, 5.3, 3.3, 5.4, 4.6, 5.4, 5.2, 1.7, 3.7, 
    2.9, 4, 2.9, 2, 2.1, 0.2, 0.5, 1.7, 0.9, 1.3, 0.2, 2.2, 1.5, 2.2, 0.2, 
    3.2, 1.5, 4.2, 2, 3, 3.6, 4.1, 5.8, 5, 4.5, 4.6, 4.8, 4.3, 4, 3.7, 1.2, 
    1, 2.9, 1.6, 1.8, 2.6, 0.4, 2.3, 1.1, 1.2, 2.4, 4, 2.5, 1.3, 2.4, 4.6, 
    4.3, 4.4, 4.6, 3.5, 1.2, 2.4, 2.6, 4, 4.4, 2.9, 2.7, 2.9, 1.3, 3.1, 4.6, 
    1.6, 5.1, 5.2, 5.5, 6.2, 5.6, 5.2, 4.2, 3.5, 4.6, 4.2, 4.7, 4.7, 5.1, 
    5.8, 5.1, 2.8, 0.7, 2.5, 1.1, 3.3, 1.1, 2.6, 2.9, 4.1, 3.4, 2.4, 2.3, 2, 
    3.1, 1.6, 1.4, 1.5, 2, 2.5, 1.4, 2.2, 3.5, 2.1, 3.2, 0.9, 2.9, 1.1, 2.1, 
    1.4, 0.9, 0.7, 1.1, 2.1, 2.3, 2.7, 2.4, 1.9, 1.6, 2, 2, 2.2, 2.3, 2, 2.5, 
    1.9, 1.6, 1.2, 1.8, 0.9, 1.7, 0.5, 2.8, 0.5, 1, 0.8, 0.9, 1.2, 1.1, 1.8, 
    1.8, 1.4, 0.1, 2, 1.7, 2.2, 2.1, 2.5, 2.2, 2.5, 3.1, 3.5, 3.3, 2.6, 1.8, 
    1.1, 3, 2.7, 2.8, 2.4, 4.9, 1.5, 3.4, 2, 3, 4.6, 2.7, 3.1, 3.3, 1.1, 3.1, 
    4.8, 6.9, 6.1, 5.9, 0.6, 2.6, 2, 2.1, 1.4, 1.1, 0.8, 1, 3.5, 3, 3, 1, 
    3.2, 5, 3.1, 1.4, 1.5, 1.1, 1.2, 0.9, 3.5, 1.3, 0.4, 0.8, 1.3, 5.2, 1.3, 
    1.5, 0.9, 0.2, 1.1, 0.2, 2.6, 2.7, 2.3, 2.9, 2.1, 3, 2.5, 4, 0.7, 1, 1.9, 
    1.2, 0.8, 2.2, 2, 1.9, 1.3, 0.5, 5.6, 0.6, 2.5, 0.9, 1.7, 0.5, 2.1, 3, 
    0.6, 1, 0.8, 0.5, 1.6, 1.6, 2.1, 2.2, 1.7, 0.9, 1.9, 2.1, 2.7, 3.4, 2.4, 
    2.4, 1.8, 1.2, 0, 0.7, 0.7, 0.4, 0.2, 1.6, 2, 1.2, 1.2, 1.7, 1.3, 2.6, 
    4.7, 3.9, 3.7, 4.6, 2.9, 2.5, 2.8, 3.2, 4.1, 3, 3.7, 4.9, 3.4, 4, 2.9, 
    3.2, 3, 2.5, 2.9, 1.9, 3.1, 3.7, 3.4, 2.8, 3.6, 3.6, 4.4, 4.4, 3.7, 4.8, 
    3.4, 4.1, 4.3, 2.9, 2.5, 3.2, 4, 2.5, 4.2, 3.8, 3.6, 4, 3.2, 3.6, 2.1, 
    4.3, 4.6, 3.6, 3.7, 5.2, 4.1, 3.3, 3.3, 2.8, 2.2, 2.8, 3, 2, 1.7, 0.6, 1, 
    2.2, 0.7, 1.4, 1.3, 1.1, 2, 2.2, 2.1, 1.1, 2.8, 2.8, 3.3, 2.8, 3.5, 2.8, 
    3.5, 3.4, 3.8, 3, 4, 3.2, 4.3, 4.2, 3.2, 2, 1.3, 1.9, 2.3, 2.2, 5.2, 3.3, 
    2.1, 5.4, 5.4, 5.2, 4.3, 5.5, 6, 5.2, 6.1, 5.7, 5.2, 5.2, 4.1, 3.7, 5.2, 
    5.2, 3.7, 3.6, 2.9, 3.5, 3.8, 3.6, 3.5, 3.3, 1.8, 2.7, 3.7, 3, 1.7, 3.7, 
    3.2, 3.7, 3.7, 3.1, 4.2, 4, 3.8, 3.7, 4.1, 3.8, 2.3, 2.4, 1.6, 0.8, 0.6, 
    2.1, 1, 1.5, 1.2, 1.7, 2.9, 2.3, 1.9, 0.9, 1.7, 2.9, 3.7, 3.2, 3.5, 2.8, 
    3, 1.5, 1.7, 1.1, 1.7, 0.2, 1.1, 1, 0.1, 1.3, 1.7, 2.4, 1.9, 2.3, 1.5, 
    1.2, 1.2, 1.5, 0.4, 1.7, 2.1, 2.4, 1.7, 1.6, 1.7, 2.3, 1.7, 1.8, 0.7, 
    0.4, 1.6, 2.4, 1.1, 0.7, 1.5, 1.9, 2.5, 1.7, 1, 3.7, 2.5, 2, 3.5, 1.7, 
    2.1, 3, 2.1, 2.7, 1.6, 2.7, 1.6, 1.7, 0, 1.3, 0, 0.5, 0, 0.8, 1, 1.2, 
    0.5, 1.4, 1.8, 1.8, 2.1, 2.1, 1.7, 2.1, 2.2, 2.3, 3.3, 2.3, 1.8, 2.1, 
    1.9, 2.6, 1.4, 2.3, 2.2, 1.2, 1.8, 1.8, 1.2, 2.4, 1.9, 2.1, 3, 2.4, 2.2, 
    2, 1.2, 2.8, 2.9, 2.5, 2.8, 2.2, 1.4, 1.1, 1.4, 1, 2, 2.9, 2.7, 0.7, 1.4, 
    2, 2, 1, 1.5, 1.9, 1.6, 1.1, 1.8, 1.8, 2.4, 2, 1.9, 1.2, 1.4, 1.6, 1.8, 
    1.7, 1.1, 1.7, 1.6, 0.6, 0.6, 0.7, 0.6, 0.9, 0.9, 0.6, 0.7, 1.9, 2.2, 
    2.3, 2.4, 2.1, 2.3, 1.9, 0.3, 2, 1.7, 2.1, 2.8, 2.4, 1.8, 0.8, 0, 0.4, 
    0.1, 0, 0, 0.3, 1.5, 1, 2.2, 2.2, 2.4, 2.9, 3.1, 2.3, 1.3, 2.9, 2.8, 2.9, 
    3.2, 2.9, 2.2, 1.9, 3.4, 1, 1.1, 1.4, 0.4, 0.6, 0, 0.3, 0.2, 1.6, 2.3, 
    2.1, 0.7, 2.2, 3.1, 1.5, 3, 2.1, 3.9, 3.6, 4, 4.5, 6.3, 3.7, 3, 2.1, 1.9, 
    2.1, 1.1, 3.9, 5.6, 1.9, 0.8, 0.8, 1.8, 2.2, 2.3, 1.4, 2.1, 1.5, 0.6, 
    1.5, 2, 2, 1.5, 1.4, 1.3, 1.5, 1.2, 1.1, 1.1, 0.6, 0.1, 0.5, 0.5, 0.7, 
    4.6, 4, 2.4, 2.9, 3.5, 1, 1.4, 2.8, 2.4, 2.7, 2.9, 2.8, 2.5, 3.6, 3.5, 
    1.9, 1.9, 2.2, 1.7, 1.1, 1.4, 1, 0.4, 0.4, 2, 1.6, 1.7, 1.7, 2.2, 2.4, 
    1.7, 1.9, 2.5, 1.9, 3, 2.7, 2.1, 2.7, 2.2, 3.9, 2.2, 3.4, 3.1, 1.7, 2.8, 
    3.9, 3.8, 4.2, 3.5, 3.9, 2.3, 4.5, 4.4, 4.4, 4, 3.9, 5.2, 3.4, 3.6, 3.8, 
    2.4, 3.7, 3.4, 4, 2.6, 3.3, 3.2, 3, 3, 2.4, 3.5, 3.2, 1.8, 1.1, 1.3, 1.8, 
    3.3, 3.1, 2.8, 3.5, 3.6, 2.8, 2.6, 3.1, 3, 3.7, 3.6, 3.1, 3.1, 2.8, 2.7, 
    1, 3.3, 3.2, 2.4, 3.4, 4.4, 3.2, 2.5, 2, 1.7, 2.6, 3.7, 1.3, 2.7, 3.1, 
    2.9, 2.4, 2.7, 4.4, 3.4, 3.2, 2.8, 2, 3.1, 2.3, 1, 1.3, 4.1, 4.1, 4.5, 2, 
    4.2, 3.9, 2.8, 3.2, 3.1, 3.7, 3.4, 3.3, 4.3, 3.9, 3.5, 3.9, 3.9, 3.1, 
    1.6, 3.1, 2.7, 2.1, 2.2, 1.5, 1.4, 2.2, 2.6, 1.8, 2.7, 2.4, 1.4, 3.4, 
    1.4, 1.5, 1.3, 1.2, 1.3, 4.4, 2.8, 4.8, 7, 7.5, 5.2, 4.9, 5.7, 4.9, 7.4, 
    3.4, 5.9, 5.2, 4.8, 5.7, 6.4, 5, 4.7, 4.9, 4.5, 3.6, 5, 5, 5.8, 4, 4.4, 
    3.9, 2.9, 3.4, 1.9, 0.7, 1.4, 0.9, 0.2, 0.5, 0.6, 0.2, 1, 0.3, 0.7, 2.1, 
    1.2, 0.8, 1.3, 1.6, 0.3, 0.7, 1.1, 0.8, 1, 0.1, 1.1, 1.3, 0.2, 0.2, 0.8, 
    1, 0.1, 0.7, 0.2, 0.4, 0.6, 1.4, 1.1, 0.3, 0.9, 0.5, 0.6, 0.5, 1, 1.6, 
    0.5, 1.7, 0.9, 1.3, 1.6, 0.7, 1.1, 0.2, 0.2, 0.2, 0.8, 0.5, 0.3, 0.2, 
    0.9, 0.7, 0.2, 0.8, 1.5, 0.6, 0.3, 0.6, 0.9, 1, 1.2, 1.6, 1.8, 1, 1.3, 
    1.1, 1.4, 0.6, 1.1, 0.2, 1, 1, 0.3, 0.3, 0.8, 0.9, 0.6, 1.1, 0.7, 0.9, 
    0.5, 0.7, 1.3, 1.9, 1.8, 1.5, 2, 2.4, 2, 2.5, 3.2, 1.9, 2.9, 1.9, 2.2, 
    1.6, 1, 0.2, 0.5, 0.4, 0.7, 1.2, 0.9, 0.6, 0.6, 1.4, 0.6, 0.7, 0.3, 1.1, 
    0.7, 1.2, 1.4, 0.9, 0.4, 0.5, 1.8, 1, 1.3, 0.2, 3.1, 4.9, 3.8, 3.5, 2.6, 
    4.7, 3.3, 4.5, 1.5, 3.3, 3.4, 1.4, 4.8, 4.3, 5.4, 2.4, 4, 4.4, 1.4, 5.1, 
    3.2, 8.1, 6.4, 3.8, 3.2, 3.9, 1.6, 4.4, 6.1, 0.8, 2.7, 0.3, 1.4, 3.5, 
    2.6, 1.3, 1.9, 2.1, 1.1, 2.4, 3.3, 1.9, 1.7, 1.7, 0, 0.4, 1.1, 1.4, 0.9, 
    1.3, 3, 2.6, 1.4, 1.6, 1.8, 1, 1.6, 2.5, 1.4, 1.8, 2.3, 1.5, 1.3, 0.7, 
    1.3, 1.4, 1.2, 0.9, 0.6, 3.4, 1.2, 3, 3.5, 2.6, 3.3, 3.6, 3.4, 3.4, 1.9, 
    2.3, 2.9, 4.2, 2.4, 3.8, 4.8, 3.9, 4.2, 3.7, 3.7, 3.4, 4.3, 4.2, 3.3, 
    3.8, 3.8, 3.3, 2.4, 2.2, 1.8, 0.4, 1.3, 1.2, 1.4, 1.3, 2.3, 0.4, 2.6, 
    2.7, 2.9, 3.1, 2.4, 3, 1.7, 2.9, 2.1, 1.9, 2.5, 1.2, 0.2, 1.5, 1.4, 2.3, 
    2.1, 1.9, 1.7, 1.4, 1.4, 2, 2, 2.4, 2.2, 1.8, 1.6, 1.6, 1.6, 1.8, 2.3, 
    0.8, 1, 1.1, 0.1, 1.1, 2.2, 1.3, 1.8, 1.8, 1.1, 2.1, 2.2, 0.3, 1.7, 2.6, 
    3.2, 2.8, 2.4, 3.3, 3.5, 3.2, 2.4, 2.5, 1.9, 1.9, 2.5, 3.6, 1.4, 0.8, 
    2.6, 2.2, 4.9, 3.7, 2.2, 1.2, 3.8, 5, 5, 1, 5.4, 5.3, 2.3, 3.4, 4.3, 2.1, 
    5.3, 6.4, 1.2, 0.1, 3.2, 0.5, 0.8, 0.7, 1.7, 0.5, 2, 0.7, 2.1, 0.4, 0.2, 
    0.3, 1.1, 2.3, 2.3, 2.5, 2.3, 2.5, 2.5, 2.3, 2.8, 3.2, 3, 1.9, 0, 0.9, 
    1.1, 0, 0.7, 0.2, 1.6, 2.1, 2.6, 2, 3.2, 2.7, 3, 2.9, 2.7, 3.4, 3.3, 3.2, 
    3.2, 3.3, 3.9, 3.8, 3.9, 3.1, 1.7, 1.7, 1.8, 1.4, 0.8, 0.1, 1.1, 0.2, 
    0.4, 1.8, 2.1, 3.1, 3.2, 3.9, 3.4, 3.7, 2.9, 4.2, 3.2, 3, 3.2, 2.8, 3.7, 
    3.5, 2.3, 3.2, 3.6, 3.1, 2.5, 2, 2.7, 1.9, 3.1, 0.2, 1.8, 0.4, 0.7, 1.2, 
    3.5, 4.6, 5.8, 3.9, 5.3, 5.6, 3, 2.4, 4, 1.8, 0.5, 1, 0.3, 5.1, 1.1, 3.7, 
    4, 0.2, 1.1, 3.7, 2.5, 4.1, 4.6, 2.8, 2.3, 1.9, 2.7, 2.1, 2, 1.1, 2.8, 
    1.1, 0.6, 3.7, 6.2, 4.2, 5.1, 6.4, 1.5, 4.7, 5.4, 5.5, 4, 3.6, 2.5, 4.5, 
    2.9, 3.8, 3, 3.9, 4.4, 1.5, 3.9, 1.3, 3.2, 5, 1.4, 0.9, 1.4, 1.1, 3.8, 
    3.4, 4.9, 5.7, 2.6, 6.3, 6.4, 6.3, 6, 3.1, 1.1, 0.9, 2.7, 5, 1.7, 3.7, 
    4.1, 1.2, 1.5, 0.4, 3.8, 4.3, 1.3, 3.8, 0.4, 1, 1.3, 0.6, 0.7, 3.8, 0.9, 
    0.7, 2.2, 0.9, 1.2, 1.4, 2.1, 2.5, 2.5, 2.1, 3.1, 3.3, 2.2, 4.6, 3.3, 
    2.9, 3, 3.2, 3.2, 1.9, 2, 2.3, 2.5, 2.5, 1.5, 3.3, 2.5, 3.1, 1.3, 2, 1.5, 
    1.8, 4, 4.4, 3.8, 2.9, 2.9, 3.4, 3.9, 3.6, 3.4, 2.8, 3.3, 2.7, 2.1, 2.5, 
    2.4, 3.1, 3, 1.7, 1.3, 1, 1.6, 3, 0.4, 1, 2.9, 1.6, 3.3, 1.8, 1.9, 1, 3, 
    2.9, 3.2, 2.5, 3.2, 3.2, 2.2, 2.6, 2.7, 1.8, 0.8, 1.1, 0.8, 1.5, 0.6, 2, 
    2, 2.3, 1.6, 1.7, 1.5, 1.6, 2.5, 2.1, 2.3, 1.8, 1.5, 2, 1.4, 1.8, 2.7, 
    2.4, 2.5, 2.4, 1.7, 1.4, 0.5, 0.7, 0.8, 1.1, 1.4, 2, 1.6, 1.8, 1.5, 2.5, 
    3.7, 3.7, 0.2, 2.9, 2.5, 1.8, 1.5, 0.2, 0.6, 1.1, 1.9, 2, 2.1, 2.1, 1.4, 
    0.8, 0.6, 0.3, 0.9, 0.7, 1.6, 1.7, 1.1, 0.7, 0.8, 1.4, 1.1, 0.7, 0.7, 
    1.3, 0.3, 1, 0.1, 0.9, 0.7, 0.6, 0.4, 0.3, 0.2, 0.5, 0.4, 0.9, 1.2, 1, 
    1.1, 1.1, 1.5, 2.1, 5.1, 3.1, 4.1, 4.3, 4.7, 3.2, 5, 4.2, 5.6, 6, 4.1, 
    5.1, 4.3, 3.1, 2, 2.3, 3.7, 4.4, 3.6, 3.9, 2.8, 3.2, 3.2, 2.6, 6.4, 6.2, 
    5.2, 3.9, 3.6, 2.4, 1.6, 0.9, 2.1, 1.3, 1.4, 1, 0.6, 0.6, 0.8, 1, 2.7, 3, 
    7.2, 7.4, 6.8, 5, 7.2, 5.8, 3.3, 4, 4.4, 4.7, 1.3, 6.2, 5.8, 4.6, 3.6, 
    2.9, 2.2, 1.5, 0.8, 1.7, 2.3, 1, 3.7, 3.6, 3.7, 4, 3.9, 2.3, 2, 2, 1.4, 
    1.1, 1.2, 0.8, 0.3, 1.1, 0.1, 0.2, 0.2, 0.5, 1.3, 0.3, 1.1, 2, 1.2, 2.1, 
    2.7, 3.2, 2.8, 2.4, 1, 1.6, 1.5, 1.4, 0.5, 1, 1.3, 1, 0.2, 0.4, 0, 0.5, 
    0, 0, 0, 0, 0.2, 1.2, 2.6, 2.7, 4.1, 3, 2.5, 2.8, 2.2, 1.4, 1.8, 2.5, 
    2.6, 1.4, 2.3, 2.2, 0.4, 1.4, 1, 1.5, 1.4, 1.2, 1, 0.8, 1.9, 4.8, 4.6, 
    2.2, 5, 8.3, 4.7, 6.9, 7.2, 6.4, 7.5, 4.6, 5.6, 4.7, 5.4, 4.5, 4.4, 3.8, 
    3.1, 2.8, 2.5, 2.4, 2.6, 3.4, 2.3, 1.7, 2.5, 2.1, 1.5, 2.7, 2.4, 3, 2.3, 
    3.4, 3.2, 3.6, 3.6, 3.2, 1.9, 1.7, 2.4, 0, 0, 0.8, 0.6, 0, 0, 0.1, 0.4, 
    0.7, 0.8, 0.6, 1.6, 1.7, 1.3, 1.7, 0.8, 2, 1.5, 3, 2.5, 2.2, 1.4, 2.7, 
    1.8, 3.3, 2.5, 1.2, 0.5, 0.5, 0, 0.4, 0, 0.3, 0.7, 1.6, 0.7, 0.1, 0, 1.8, 
    1.4, 1.2, 0.8, 1, 0.4, 3.3, 3.5, 3.6, 3.3, 3.2, 5.8, 5.5, 4.9, 4.8, 5.4, 
    2.2, 2.8, 1.7, 3.5, 4.5, 3, 1, 1.3, 0.9, 0.4, 0.4, 3.8, 2.6, 1, 5, 4.8, 
    4.6, 5.5, 5.5, 4.4, 3.7, 5.5, 4.8, 4.3, 4.5, 3.8, 4.5, 3.4, 4.5, 4.7, 
    3.8, 3.6, 2.8, 0.7, 3, 4.5, 5.3, 4.9, 3.4, 4, 4.3, 2.9, 5.3, 3.8, 4, 2.6, 
    2.1, 2.7, 1.1, 0.5, 1.5, 1.5, 1.2, 1.3, 1, 1.8, 1.3, 0, 0.8, 0.9, 0.3, 
    1.2, 3.6, 3.8, 3.6, 2.7, 4.1, 5, 5.5, 4.3, 4.4, 5.7, 4.5, 3.4, 3.6, 4, 
    4.9, 5.7, 5.6, 3.5, 3.8, 4.7, 5.3, 4.9, 4, 4.2, 3.4, 3.9, 3.9, 4.3, 7.8, 
    4.6, 4.6, 4.8, 4.8, 2.4, 3.4, 4.3, 4.4, 4.9, 4.4, 4.3, 3.9, 5.1, 5.6, 
    5.6, 4.8, 4.5, 4.1, 4.5, 3.6, 2.5, 4.6, 4.2, 1.8, 1.1, 2, 1.2, 4.2, 4.8, 
    5.4, 3.2, 2.3, 2.3, 1.3, 3.9, 4.5, 3.4, 3.1, 4, 1.9, 2.3, 2.2, 2.7, 2.6, 
    2.3, 1.9, 2.5, 2.6, 1.2, 0.8, 0.9, 1, 1.4, 0.1, 1.2, 1.8, 0.3, 1, 1.4, 
    1.3, 1.5, 2, 2.7, 2.4, 2.2, 1.8, 3, 2.3, 1.6, 0, 0.7, 2.2, 1.2, 0.2, 0.1, 
    0.9, 2.5, 3.3, 1, 3.9, 1.8, 6.6, 3.7, 3.1, 3.4, 2.6, 3.7, 6.6, 5.2, 6.4, 
    5.1, 3.7, 0.9, 2.1, 2.2, 2.1, 3.8, 3, 2, 1.7, 2, 1.6, 1, 2.5, 2, 1.4, 
    2.9, 3, 2.6, 2.7, 2, 4.3, 4.3, 2.9, 1.4, 2.2, 0.2, 0.9, 0.2, 0, 0, 0.3, 
    3.7, 0.1, 1.1, 1.2, 1.4, 0.9, 0.1, 0.1, 4.7, 1, 1.7, 1, 1.1, 0.4, 0.3, 
    0.3, 0.2, 0.2, 0.3, 0.3, 0.5, 1, 3.5, 3.3, 1.8, 1.7, 1.1, 5.3, 1.4, 0.4, 
    0.2, 3.1, 4.4, 4.8, 5.1, 3.6, 4.8, 5.3, 4.2, 5.1, 4.5, 4.5, 4.6, 5.2, 7, 
    6.9, 5.1, 5.5, 3.8, 3.3, 3.1, 4.1, 3.1, 4, 3.8, 3.8, 3.3, 4.1, 3.4, 2, 
    3.1, 2.3, 1.8, 2, 2.3, 1.7, 1.3, 0.8, 1, 1.7, 1.6, 1.2, 4, 2.2, 3.9, 2.4, 
    2, 4.6, 4.6, 3.1, 3.9, 3.6, 3.7, 2.6, 3.7, 1.6, 1.8, 2.6, 1.8, 1.1, 0.6, 
    0.6, 0.9, 0.7, 2.8, 0.6, 1.6, 0.7, 1.9, 1.1, 0.1, 1.2, 1.7, 1.1, 0.5, 
    1.4, 0.7, 0.3, 1.3, 0.9, 1.2, 1.6, 1.1, 0.8, 2.2, 3.1, 2.9, 0.1, 0.5, 
    0.2, 2.2, 0.3, 0.5, 0.5, 0.4, 0.6, 0.8, 0.9, 1.6, 2.6, 1.6, 2.2, 1.9, 
    1.2, 0.4, 0.7, 2.7, 2.2, 1.3, 0.9, 0, 0.1, 1.1, 0.3, 0, 0.8, 0, 0.1, 0.3, 
    0.7, 1.1, 1.2, 0.8, 2.8, 4.3, 7.1, 5.9, 5.7, 5.6, 4.2, 4.9, 3.2, 4.4, 
    4.7, 4.3, 4.1, 4.9, 3.3, 2.2, 1.5, 2.4, 1.5, 1.6, 2.2, 1.2, 0.4, 0.7, 
    0.9, 2.2, 1.9, 2.2, 3.2, 3.4, 3.8, 2.6, 2.6, 2.5, 4.4, 1.9, 0.5, 1, 1.4, 
    1.7, 1.8, 0.3, 0.8, 0.4, 1, 0.1, 0.4, 0.8, 1.5, 1.6, 2, 1.8, 1.3, 1, 1.5, 
    0.9, 0.2, 0.3, 0.7, 1, 0.9, 0.5, 0.2, 0.4, 2.3, 0.1, 1.8, 0.3, 0, 0.9, 
    0.8, 1.6, 1.5, 1.6, 1.7, 1.2, 1.9, 1.6, 2.4, 1.5, 2.4, 1.7, 1.4, 0.5, 
    1.7, 1.4, 0.5, 0.6, 1.2, 1.6, 0.6, 0.9, 0, 0.5, 1.7, 1.5, 0.8, 1.4, 1.3, 
    0, 1.6, 1.1, 1.3, 0.6, 0.6, 0.6, 0.5, 0.4, 0.7, 0.6, 0.7, 0.1, 0.6, 0.7, 
    0.2, 1, 0.7, 1, 0.9, 0.1, 1.9, 2.1, 0.9, 0.8, 0.4, 1.3, 1.4, 0.7, 0.8, 
    1.1, 1.3, 1.1, 1, 0.8, 1.1, 0.7, 1.3, 0.3, 0.4, 0, 1.1, 0.9, 1.3, 0.2, 
    0.7, 1.6, 1.9, 1.2, 0.5, 0.5, 0.4, 0.2, 0.6, 0.2, 0, 0.1, 0.4, 0.4, 1, 
    0.6, 0.5, 0.2, 0.3, 0.5, 0.1, 0.7, 0.9, 2, 1.7, 1.4, 1.3, 0.7, 0.2, 0.5, 
    0.4, 2.1, 1.4, 1.8, 1.7, 0, 0.3, 0.5, 0.1, 0.1, 0, 0.1, 0.5, 0.3, 0, 0, 
    1.1, 1.2, 1.2, 1, 1.7, 1.3, 1.3, 0.4, 0.4, 1.8, 1.4, 0.7, 1.3, 0.4, 0.3, 
    0.3, 0.3, 0.4, 0.6, 0.1, 0.1, 1.4, 0.5, 0.1, 0.5, 0.6, 1.6, 2.4, 3, 1.1, 
    0.9, 0, 0.1, 0.2, 0.3, 0.8, 2, 1.3, 0.6, 1.2, 0.7, 0.8, 1.2, 0.7, 0.1, 
    0.2, 0.3, 0, 0.9, 1, 0.4, 0.6, 0.6, 0.2, 0.9, 0.7, 0.1, 0.9, 0.1, 0.2, 0, 
    0.9, 0.6, 0.8, 0.3, 1, 0.7, 0.2, 0.2, 0.3, 0.4, 1.7, 0.1, 0.2, 0, 0.8, 
    1.1, 0.7, 0.9, 1.5, 1.1, 0.9, 0.5, 1, 1, 1, 0.5, 0.9, 1, 1.1, 1, 0.5, 
    0.8, 0.3, 1.4, 1.2, 1.1, 2.4, 1.7, 0.8, 0.8, 1.1, 3.7, 2.4, 1.6, 6.6, 
    4.9, 4.8, 4.9, 5.4, 4.3, 4.9, 5, 3.9, 4, 3.7, 2.6, 3.3, 2.7, 3, 3.4, 2.9, 
    2.2, 1, 2.2, 2.7, 2.7, 4, 0.8, 2.3, 0.7, 0.8, 1, 1.2, 2.2, 0.6, 0.8, 0.7, 
    0, 1.3, 0.8, 1.8, 1.6, 1.8, 1.2, 2.1, 1.2, 1.2, 0.4, 0.6, 1.3, 1, 1.2, 
    2.8, 0.6, 0.9, 2.1, 1.8, 1.4, 0.6, 0.2, 0.7, 2.8, 1.5, 0.6, 0.3, 0.3, 
    0.7, 1.3, 0.1, 1.7, 1.7, 1.3, 1.9, 1.4, 1.1, 3.5, 1, 3.4, 3.8, 3.1, 3.6, 
    3.8, 5.4, 4.7, 4.7, 1, 1.1, 1.1, 0.9, 1.2, 0.9, 1.1, 0.6, 0.9, 0.6, 3.1, 
    2.5, 1.2, 5.1, 1, 0.6, 1.7, 2.6, 7, 12.4, 9.4, 13.9, 13.8, 13.4, 8, 12.6, 
    6.9, 4.4, 2.3, 3.5, 3.5, 3.4, 3.9, 3.7, 3.9, 3.7, 4, 4.3, 2.7, 3.5, 2.5, 
    3.7, 3.1, 2.4, 2.3, 0.3, 0.8, 0.1, 0.3, 0.3, 0.8, 0.3, 1.5, 0.1, 0.8, 0, 
    1, 0.1, 1.2, 1.6, 1.9, 1.4, 1.3, 0.9, 1.1, 0.6, 0.8, 0.1, 0.4, 2.3, 1.9, 
    4.1, 0.5, 1.2, 1.6, 4.5, 1.9, 2.9, 4.5, 7, 6.7, 3.8, 7.7, 6.8, 4.7, 4.9, 
    5.4, 4.4, 3.6, 4.3, 4.2, 4.4, 4, 3.7, 1.9, 1.4, 0.4, 3.9, 0.9, 0.7, 1.2, 
    1.5, 2.1, 1.5, 2.3, 3.5, 3.8, 4.5, 3.8, 3.7, 3, 3.1, 2.6, 4.1, 2.3, 0.9, 
    1.2, 1.9, 1.5, 1.6, 1.1, 1, 0.7, 1, 2.3, 2.1, 0.8, 0.4, 3.1, 1.5, 1, 0.5, 
    0.6, 0.3, 0.8, 0.1, 0, 0.2, 0.8, 0.2, 0, 1.4, 0.1, 1.9, 0.1, 0, 0, 1.1, 
    0.3, 0.6, 0.4, 0, 0, 0.3, 0, 0, 0.5, 0.5, 0.2, 0.8, 0.5, 1.4, 0.4, 0.5, 
    0, 0.8, 0.3, 0.4, 0.8, 0.3, 0, 0.1, 0.5, 0, 0, 0, 0.2, 1.1, 0.4, 0.2, 
    0.4, 0.7, 0, 0.4, 0.2, 0.1, 0.8, 1, 1.1, 0.1, 0.4, 0.7, 1.2, 0.5, 0.5, 
    1.3, 0.6, 0.8, 0.5, 0.8, 0.8, 1.3, 0.6, 1.4, 1.9, 0.5, 1.8, 1.1, 0.8, 
    1.8, 2.2, 1.3, 1.4, 7.1, 1.7, 1.5, 1.3, 1.7, 1.4, 0.9, 1.2, 0.6, 0.1, 
    0.1, 0.2, 0.2, 1.4, 1.5, 0.7, 1, 1.2, 1.5, 1.5, 1.4, 0.4, 1.1, 3.6, 1.6, 
    0.9, 0.5, 0.4, 0.5, 1.4, 1.7, 0.6, 0.8, 1.2, 0.4, 1.8, 0.9, 0.8, 1.2, 
    0.7, 0.5, 0.7, 1.2, 1.4, 0.6, 0.4, 0.4, 0, 1.2, 1.2, 1.1, 3.3, 1.8, 2.6, 
    8.6, 8, 6, 2.6, 2.5, 2.9, 2.6, 3.9, 6.2, 5.2, 4.7, 3.9, 4.2, 6.3, 5, 4.5, 
    3.9, 6.1, 6.2, 5.2, 5.6, 5.3, 4.3, 5, 2.6, 3.9, 2.7, 9.1, 8.1, 9.1, 7.5, 
    9.7, 9.4, 8.6, 7.2, 8.1, 8.6, 8.7, 7.9, 8.8, 7, 7.2, 5.6, 4.3, 8.2, 9.5, 
    9.8, 9.2, 9.9, 10, 7.7, 6.3, 10, 9.2, 4.5, 5.3, 6.8, 9.7, 9.3, 6.4, 4.7, 
    3, 3, 3, 2.5, 3.2, 1.3, 2.4, 2.4, 1.1, 0.6, 0.9, 1.4, 0.8, 0.4, 0.6, 0.5, 
    0.4, 0.5, 0.4, 0.3, 1, 0, 0.1, 1, 1.1, 0.8, 0.5, 1.2, 0.7, 0.7, 0.6, 0.9, 
    1.2, 1.7, 3.5, 4.1, 5.8, 5.5, 4.5, 3.2, 3.5, 2.9, 1.8, 1.4, 1.9, 3.7, 
    2.9, 4.6, 3.7, 4.6, 3.2, 5.2, 4.1, 2.7, 3.2, 1.8, 2.6, 1.6, 0, 0.9, 1, 1, 
    4.1, 2.6, 2.7, 3.1, 1.3, 0.7, 0, 0.3, 0.3, 1.3, 0.9, 0.1, 4.2, 3.5, 0.7, 
    0.5, 1.6, 0.6, 1.6, 2.2, 5.1, 1.2, 1.9, 0.5, 0.9, 1.4, 2.6, 3, 3.6, 2.5, 
    3.5, 3.9, 3.5, 3.7, 2.9, 1.4, 0.9, 0.3, 1.4, 5.6, 1.2, 1.6, 0.2, 1.1, 
    0.4, 1.2, 0.7, 0.1, 0.5, 1.1, 0.8, 1.9, 1.1, 2.7, 0.3, 2.3, 2.3, 1.4, 
    1.5, 1.3, 0.9, 3.8, 4, 1.4, 1.2, 1, 1.5, 6.3, 7, 7.4, 5.1, 8.3, 11, 9.1, 
    10.5, 8.4, 3.4, 3.5, 5.3, 4.1, 3.5, 8.9, 6.4, 5, 3.3, 3.5, 4.8, 5.2, 2.7, 
    3.5, 4.3, 3.5, 2.3, 2.1, 2, 3, 0.8, 1.2, 0.3, 0.2, 0.6, 1.1, 0, 0.2, 0.4, 
    0.1, 0, 1.1, 1, 0.5, 0.3, 0.6, 1, 0.6, 0.5, 1.4, 1.6, 0.7, 1.2, 0.6, 1.5, 
    0.8, 1.5, 3.8, 3.6, 2.7, 1.1, 0.1, 4.4, 3.6, 3.7, 4.4, 4.9, 7.7, 7.6, 
    4.9, 3.8, 4.2, 7, 6.6, 4, 3.6, 3.4, 5.2, 2, 3.6, 3.3, 3.2, 4.5, 3.9, 4.5, 
    4.3, 2.5, 2.2, 2.9, 3.4, 3.1, 2.4, 4, 4.5, 4.1, 2.8, 2.8, 2.6, 3.6, 2.9, 
    2.5, 2.5, 0.8, 1.8, 1.1, 1.1, 1.9, 0.7, 0.6, 0.5, 0, 0.2, 0, 0.3, 0.8, 0, 
    0.1, 0.6, 0.6, 0.3, 0.4, 0.5, 0, 0.4, 1.8, 2.8, 4.3, 3.5, 3.7, 3.4, 3.7, 
    3.7, 1.9, 0.7, 0.5, 0.8, 0, 1.2, 1.6, 1.4, 0.8, 0.4, 0.4, 0.8, 0.1, 0.1, 
    1.6, 1.1, 1.2, 0, 1, 0.8, 1.5, 0.8, 0.7, 0, 0.3, 2.6, 2.7, 1.9, 0.6, 0.7, 
    0.7, 0.6, 1.5, 0.8, 1.1, 2, 2.2, 1, 1.8, 1.3, 2, 0.6, 0.2, 0, 0.6, 0.1, 
    0.4, 5, 4.5, 4.8, 8, 9, 8.8, 7.8, 4.7, 3.3, 4.4, 3.9, 4.9, 4.7, 4.7, 3.4, 
    4.4, 4.8, 5.5, 6.4, 6.2, 6.5, 5.3, 7.9, 6.6, 7, 4.8, 5.7, 7.4, 6.7, 5.7, 
    8.5, 7.8, 5.7, 7.7, 5.8, 7.7, 6.6, 6.3, 5.2, 3.8, 3.8, 3.6, 3.6, 3.6, 
    2.7, 3.1, 2.3, 1.7, 0.7, 0.9, 0.7, 2.7, 1.5, 1.7, 2.5, 3.3, 2.4, 1.5, 
    1.7, 1.6, 0.3, 0.2, 0.9, 0.7, 0.3, 0.1, 0.4, 1, 1.9, 2.1, 0.4, 0.2, 1, 
    1.2, 1.1, 0.6, 0, 1.9, 0.7, 2.1, 1.8, 1.4, 0.8, 2.1, 3.2, 1.9, 0.5, 1.2, 
    0.5, 0.6, 0.8, 0.9, 0.9, 0.2, 1, 1.2, 0.3, 1.3, 0.9, 0.2, 0, 0.4, 0, 0.3, 
    5.4, 3.6, 3.7, 2.6, 2.6, 0.1, 1.2, 0.2, 0.6, 0.1, 0.9, 0.2, 0, 0.2, 1.1, 
    1.2, 0, 0.8, 0.2, 0.4, 1, 0.8, 0.6, 4.6, 0.5, 0.9, 4.4, 1.1, 3.6, 5.1, 
    3.3, 4.3, 4.9, 4.8, 4.9, 5.2, 4.8, 5.2, 2.8, 3.6, 4.3, 5.3, 5.3, 6.2, 
    5.5, 7.6, 5.7, 6.1, 5.6, 8.4, 9.6, 10.3, 11.9, 11.2, 9.8, 9.1, 9.6, 8.8, 
    9.1, 8.8, 6.6, 7.1, 9.1, 7.2, 5.3, 5, 5.5, 4.8, 5, 6.7, 4.9, 4.8, 2.6, 
    3.4, 3.2, 4.8, 6.3, 5.1, 4.4, 4.3, 3.2, 5.3, 4.6, 3.5, 0.4, 1, 0.4, 2.2, 
    0.3, 0.4, 1.5, 0.2, 0.4, 0, 0.2, 0.7, 0, 0.1, 1.4, 1.1, 1.2, 0.3, 0.9, 0, 
    0.1, 0.8, 1.2, 3.7, 5.6, 3.5, 3.3, 4.3, 4.4, 3.7, 3.5, 2.7, 4.7, 4, 4.1, 
    5.5, 5.2, 3, 2.4, 3.1, 3.5, 3.8, 2.9, 1.1, 1, 0.8, 0, 0.8, 0, 0.1, 0.1, 
    0.4, 0.4, 1, 1.6, 0.7, 0.2, 0.1, 0.6, 0.4, 0.7, 1.2, 0.2, 0.9, 0.4, 0.3, 
    0.5, 2.8, 4.2, 4.5, 4.3, 4.6, 2.8, 2.1, 1.4, 0.5, 0.1, 0.4, 0.1, 0.5, 
    0.1, 0.7, 0.4, 0.4, 0.5, 1, 0.6, 0.2, 0.2, 0.3, 0.2, 0.6, 0.7, 0.5, 1.1, 
    0.7, 1.1, 0.4, 0.4, 0.9, 0.8, 1.1, 0.4, 0.8, 4.5, 1.9, 0.4, 1.5, 1.2, 
    1.2, 0.8, 0.9, 3.9, 4.6, 5.3, 5.3, 5.7, 5.4, 3.4, 4.2, 3.3, 4.3, 4.7, 4, 
    5.5, 3.9, 4.4, 4.6, 5, 6.5, 7.3, 8.3, 6.1, 5.8, 6.6, 5.5, 5.6, 4.7, 6.6, 
    7.4, 7.6, 6.7, 9.7, 8.2, 6.4, 6.9, 4.7, 4.3, 7.9, 8.1, 9.4, 8.5, 7.9, 
    5.6, 7, 4.7, 5.8, 3.4, 3.6, 5.6, 6.2, 8.4, 2.8, 1.4, 4.2, 3.2, 3.8, 5.3, 
    3.5, 2.9, 3.2, 1.7, 0.9, 3.1, 1.8, 3.4, 1.1, 2.2, 2, 0.8, 2.7, 5.4, 7.1, 
    5.2, 5.5, 3.9, 4.7, 3.5, 3.2, 3.8, 2.8, 3.7, 3.8, 3.7, 3.1, 2.7, 2, 1.1, 
    0.6, 0.7, 0.9, 3.1, 0.8, 1.5, 2.6, 3, 1.1, 1.6, 1.6, 0.4, 1, 0.7, 1.1, 
    0.1, 0.9, 1, 1.1, 0.4, 0.2, 0, 1.2, 1.4, 0.9, 0.8, 0.7, 0.3, 0.7, 0.6, 
    0.1, 1, 0.6, 0.1, 0.1, 1, 1.1, 0.3, 1, 0.3, 0.2, 0.5, 0.3, 0.9, 0.1, 0.2, 
    0.3, 0.2, 0.2, 0.8, 0.2, 1, 1.3, 1.9, 1.2, 1.2, 1.4, 1.7, 1.7, 1.6, 0.4, 
    0.8, 1.4, 1.3, 0.9, 0.2, 0.7, 0.1, 0.7, 0, 0.5, 1.1, 0, 0.1, 0.3, 0.8, 
    1.8, 0, 0.9, 0.2, 0.2, 0.2, 0.5, 0.4, 0.2, 0, 0.2, 0.1, 0, 0.1, 0.2, 1.7, 
    1.1, 1.1, 1, 0.9, 0, 0.9, 0, 0.1, 0.2, 0.1, 1, 0.7, 0.3, 1, 0.4, 1.2, 
    0.7, 0.4, 0, 0.2, 0.9, 0.4, 0.8, 1.3, 0.9, 1, 0.5, 1.9, 0.5, 0.5, 0.1, 
    0.8, 0.7, 1.4, 0, 4.2, 4.6, 3.1, 3.3, 3, 1.6, 0, 0.1, 0.8, 0.4, 0.7, 0.5, 
    1.7, 2, 2.8, 3.4, 3.9, 2.5, 2.3, 1.8, 1.5, 1.4, 0.6, 0.9, 1, 2, 1.7, 2.4, 
    0.5, 0.8, 0.1, 0.7, 0.8, 0.6, 2.8, 3.1, 3.1, 2.3, 2.5, 2.6, 2.5, 1.9, 
    3.7, 2.9, 5.2, 3.6, 2.1, 3.3, 3.2, 6.2, 5.6, 5.8, 5.5, 5.2, 5.3, 3, 2.7, 
    4.3, 6.6, 6.6, 6.9, 2.9, 2.4, 3.6, 4.7, 5.7, 6.7, 7.1, 5, 3.3, 6.1, 5.6, 
    7.6, 7.2, 9, 10.9, 12.1, 10.2, 10.2, 10.8, 7.7, 6.2, 5.3, 4.9, 6.6, 4.7, 
    4.5, 3.5, 4.3, 3.3, 4.8, 3.9, 1.7, 1.7, 0.8, 0.7, 0.4, 0.5, 1.5, 1.2, 
    0.1, 0.5, 0.3, 0, 0.2, 1.1, 0.5, 0.1, 0.2, 4, 4.4, 5.9, 4.4, 2, 5, 4.5, 
    4.4, 4.7, 5.4, 5.4, 3.3, 4.2, 3, 3.2, 4, 3, 3.5, 3.8, 3.4, 2.5, 2, 2.3, 
    2.3, 2.8, 2.3, 2.5, 0.9, 1.5, 0.1, 1, 0.7, 0.7, 1.1, 0.8, 0.7, 0.2, 0.1, 
    0.7, 0.6, 0.9, 0.9, 1, 0.4, 0.8, 0.6, 0.3, 0.7, 0.4, 0.8, 1.1, 1.5, 1.2, 
    5.4, 0.4, 1, 0.7, 0.9, 0.9, 0.7, 2.4, 1.7, 1.2, 2.1, 1, 0.1, 1.8, 2.5, 
    0.3, 0, 0, 0, 0, 2.7, 0.5, 0.6, 1.1, 1.2, 0.5, 1, 0.8, 2.1, 1.8, 0.9, 
    3.1, 1.3, 1.5, 0.4, 1.2, 1.8, 0.7, 0.3, 0.5, 0.6, 0.3, 1, 0.1, 0.3, 0.8, 
    0.5, 1.4, 0.1, 1.6, 3.3, 0.4, 4.8, 4.6, 0.9, 0.1, 1, 1.6, 2.7, 2.4, 1.5, 
    1.5, 0.7, 0.3, 1.3, 4.9, 5.5, 3.5, 2.8, 2.3, 2.3, 2.2, 7.9, 3.4, 2.3, 
    4.6, 1.4, 1.9, 5.2, 3.9, 6, 8, 8.9, 9.7, 8.2, 6.8, 6.9, 7.5, 7.2, 7.4, 
    7.1, 4.4, 4.6, 4.8, 4.8, 4.7, 4.4, 2.8, 1.7, 0.4, 2, 1.5, 0.9, 2, 1.4, 
    0.5, 0.7, 4.8, 5, 6.4, 6.2, 7.1, 5.6, 4.3, 6.5, 5.1, 7.1, 4.5, 7.1, 6.8, 
    6.6, 5.3, 6.6, 3.9, 4.7, 6.1, 4.5, 3.6, 6, 4.9, 5, 5.6, 6.1, 4.4, 2.5, 
    0.5, 0, 1.8, 1.8, 1.1, 0.2, 0.4, 0.9, 4.3, 4.1, 1.4, 0.9, 1.4, 0.9, 2, 
    1.8, 0.5, 0.7, 0.8, 0.9, 0.6, 0.3, 0.3, 1, 1.5, 0.7, 1.2, 5.3, 4.3, 3.6, 
    3.2, 2, 3.3, 4.4, 5.9, 5.3, 2.2, 1.4, 4.2, 5.7, 6.5, 7.1, 5.7, 6.8, 6.2, 
    7.1, 5.2, 5.2, 3.5, 2.4, 3.8, 6.5, 6.3, 5.6, 4.1, 4.9, 5.4, 3.3, 3.3, 
    4.8, 3.6, 3.7, 2.7, 2.3, 4.5, 4.8, 5.9, 4.8, 4.5, 4.9, 4.1, 4.9, 5.3, 
    6.3, 5.8, 6.7, 3.8, 5.6, 4.3, 6.2, 6.5, 6.3, 4.1, 4.2, 4.6, 4.9, 5, 3.4, 
    4.3, 3.9, 4.5, 4.4, 6.2, 4.3, 4.2, 4.4, 5.9, 5.5, 2.5, 4.2, 4.8, 2.2, 4, 
    4.9, 2.7, 2.3, 1, 1, 0.4, 1.2, 0.8, 1.2, 0.1, 0.5, 0, 0.4, 0.7, 1.7, 1.9, 
    2.3, 2.2, 3.2, 3, 2.1, 0.2, 0.2, 0.5, 0.8, 1, 0.6, 0.9, 2.9, 2.8, 2.5, 
    2.4, 3.3, 3.1, 3.3, 3.3, 3.7, 2, 2.3, 1.7, 2.6, 3.1, 4.4, 2.4, 3.5, 3.1, 
    2.6, 3.1, 4.4, 3.2, 0.7, 2, 2.4, 1.6, 0.8, 0.9, 1, 0.5, 1.2, 2.8, 3.2, 
    3.5, 4.5, 4.1, 3.7, 3.8, 2.2, 1.5, 0, 0.9, 0.7, 0.4, 0.4, 0.4, 0.5, 0.2, 
    0.8, 0.5, 0.8, 0.2, 0.1, 0.9, 0.5, 0.3, 1.1, 0.5, 0, 1, 0.8, 0.6, 1.2, 
    0.9, 0.9, 3.5, 4.3, 5.3, 3.6, 3.4, 4.4, 5.4, 6.4, 6.6, 4, 2, 1, 1.6, 1.5, 
    1, 1.3, 1.7, 1.9, 1.7, 1, 3.3, 2.7, 3.7, 2.5, 2.4, 2.4, 2.5, 2.1, 0.8, 
    1.3, 2, 2.3, 3, 2.9, 1.5, 4.4, 6, 6.8, 6.2, 9, 7.7, 3.9, 5.5, 1.5, 1.4, 
    0.5, 1.8, 1.2, 0.4, 1.9, 0.3, 0.3, 1.5, 0.6, 0.1, 1, 1.2, 1.4, 1.2, 1.5, 
    0.7, 0.2, 0.5, 0.2, 1.2, 1.5, 0.8, 1, 1.5, 0.8, 1.2, 0.6, 1, 0.7, 0.7, 
    0.7, 0.5, 4.3, 3.8, 4, 4, 3.7, 4.8, 4.8, 5.6, 5.8, 5.4, 5.9, 5.6, 7.7, 
    7.6, 8.5, 7.8, 9, 9, 9.5, 10.2, 10.3, 8.4, 8.6, 9.3, 7.8, 7.3, 4.3, 6.7, 
    7.7, 6.6, 6.4, 5.5, 6.9, 7.7, 8.3, 6.9, 4.9, 3.8, 2, 4.3, 3.8, 2.9, 1.4, 
    4, 4.1, 4.2, 3.9, 3.7, 3.1, 3.1, 3.9, 3.2, 4.2, 4, 2.6, 3.4, 4.4, 3.3, 
    3.6, 3.7, 1, 1.9, 4.4, 5.6, 3, 4.8, 1.2, 0.6, 0.6, 0.4, 1.4, 1.4, 1.5, 
    1.4, 1.6, 1.8, 0.8, 1.1, 1.1, 2.3, 1.5, 0.9, 0.7, 1.3, 1.3, 1.4, 0.9, 
    1.2, 1.9, 0.2, 1.3, 0.8, 1, 1.2, 0.7, 1, 1, 1.8, 0.9, 0.7, 1.1, 0.4, 0.2, 
    0.4, 2.2, 2, 3.3, 3.1, 4.4, 4, 4.3, 3.1, 1.5, 2.1, 1.8, 1.5, 2, 0.8, 1.5, 
    1.1, 0.6, 1, 0.8, 2.4, 0.7, 0.4, 0, 0.2, 1.2, 0.6, 2.5, 5, 5.6, 5.5, 4.4, 
    5.8, 6, 7.3, 5.4, 5.1, 4.8, 7.8, 7.8, 7, 6.6, 6.9, 5.5, 4.5, 5.5, 4.6, 
    3.8, 4.3, 1.7, 0.5, 1.7, 1.2, 3, 1.8, 1.7, 0.6, 0.8, 8.2, 8.7, 4.9, 7.8, 
    6, 5.3, 5.6, 5.2, 5, 5.1, 5.3, 1.6, 2.9, 2.7, 1.9, 2, 0.4, 0, 0.6, 0.1, 
    0.7, 0.3, 1.2, 1.8, 2.5, 0.4, 0.4, 1.2, 0.8, 2, 3, 3.4, 0.5, 4.9, 5.1, 
    5.4, 4, 5.6, 3.8, 1.8, 3.5, 4.6, 5.1, 5, 4.9, 5.4, 4.6, 5.5, 4.6, 1.1, 
    1.2, 0.4, 0.5, 2.2, 0.8, 2.1, 1.4, 2, 2.6, 1.3, 2.5, 0.9, 2.7, 3.5, 2.4, 
    3.5, 2.6, 1.3, 1.7, 0.9, 2.6, 1.5, 1.7, 1.7, 1.9, 3.1, 1.1, 0.3, 0.9, 0, 
    1.9, 1.1, 1.1, 1, 0.8, 2, 1.1, 0.8, 1.1, 1, 2.2, 2, 1.1, 0.5, 1.8, 0.7, 
    1.3, 2.4, 1, 1.5, 2.4, 1.4, 1.3, 1.3, 0.9, 1.1, 1.1, 1.2, 0.8, 0.1, 1, 
    0.8, 1.4, 0.7, 1.4, 2.6, 1.7, 1.7, 1.5, 1.2, 2, 0.9, 1.8, 0.7, 1.3, 0.8, 
    1.3, 0.9, 1.6, 1.1, 0.7, 1.1, 0.2, 0.4, 1.5, 1.6, 2.2, 0.2, 1.4, 1.3, 
    1.2, 0.7, 0.2, 2, 2.5, 0.9, 1.3, 0.5, 1.2, 1.4, 1.6, 1.7, 1.8, 0, 0.9, 
    1.5, 0.1, 0.9, 1.4, 1.3, 0.7, 1, 2.2, 1.6, 2, 2.4, 2.3, 1.3, 1.7, 1.1, 
    2.2, 1.3, 1.6, 1.3, 2, 1.7, 1.4, 2.1, 2.2, 1.2, 0.8, 1.1, 2.1, 1.7, 1.7, 
    2.9, 1.6, 2.2, 2.1, 3.2, 1.7, 0.8, 1.3, 1.9, 1.6, 2.1, 2.1, 0.9, 1.5, 
    1.7, 2.5, 2.8, 3.2, 2.4, 1.2, 0.9, 1.5, 0.7, 1.1, 0.4, 0.7, 1.1, 1, 0.9, 
    1, 1.7, 2, 1.1, 1, 0.5, 0.3, 0.8, 0.8, 0.5, 0, 1.3, 1.4, 0.7, 1.1, 1.8, 
    2.3, 0.2, 1.8, 0.8, 0.7, 0.1, 0.8, 0.4, 0.2, 0.3, 0.9, 1.9, 3.1, 0.7, 
    1.1, 0.9, 1.8, 1.6, 1.7, 1, 1, 0.9, 1, 1.6, 0.9, 1.2, 1.5, 2.1, 0.8, 3.1, 
    0.4, 0.9, 0.5, 0, 1, 0.1, 1.5, 1.4, 1, 0.5, 1, 0.8, 1, 1.1, 2.4, 0.3, 
    1.6, 2.1, 1.6, 1.3, 0.7, 0.7, 0.3, 0.9, 0, 0.5, 0.7, 0.5, 0.9, 0.7, 0.5, 
    0.7, 0.5, 1.7, 0.7, 0.2, 0.2, 0.7, 0.4, 0.2, 0.3, 1, 0.9, 2.7, 0.3, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 4.4, 2.5, 2.7, 5.3, 4.3, 5, 4.5, 4.4, 3.3, 4, 
    3.2, 4, 4.2, 3.4, 0.9, 1.5, 2.3, 1.7, 1, 0.6, 3.1, 1.2, 2, 0.5, 2.4, 8.5, 
    4.6, 4.8, 8.3, 8.6, 7.1, 4.8, 2.1, 3.9, 6.9, 6.8, 7.2, 7, 6.9, 5.5, 3.9, 
    3.3, 8.7, 7, 5.4, 5.6, 6.6, 4.7, 4.6, 4.5, 3.4, 7.6, 1.8, 1.3, 1.8, 1, 
    1.4, 1.7, 2.7, 1.7, 0.3, 1.3, 3.3, 7.2, 8.9, 10, 9.1, 6.4, 1.7, 0, 0.2, 
    1.4, 2.5, 3.9, 2.3, 1.4, 1.8, 2.3, 2.5, 2.5, 2.6, 2.6, 1.4, 1.4, 1.2, 
    1.4, 0.4, 1.4, 2.7, 0.6, 1.1, 0.5, 2.5, 3.3, 0.4, 1.6, 2, 2, 1, 0.8, 1, 
    2.7, 5.6, 2.1, 3.3, 5.3, 6, 6, 5.4, 5.6, 6, 4.4, 3.1, 4.1, 3.3, 4.1, 0.4, 
    0.8, 1.2, 1.6, 0.2, 0.7, 1.1, 0.6, 0.5, 0.1, 0.1, 0.5, 0.4, 1.3, 0.1, 
    0.8, 0.5, 0.1, 0.6, 0.4, 0.4, 0.6, 0.7, 1.8, 1.4, 0.9, 0.9, 3, 1.3, 2.5, 
    0.5, 0.8, 1.7, 0.8, 0.7, 0.1, 0.3, 0.4, 0.7, 0.7, 0.4, 0.1, 0.8, 0.4, 
    1.4, 0.6, 0.6, 0.1, 1.6, 1, 0.5, 1.2, 1.5, 1.1, 0.6, 0.7, 2.6, 1.4, 0.1, 
    0.2, 0.2, 1.1, 3.4, 1.5, 1.5, 1.2, 2.4, 0.7, 0.6, 1.8, 0.9, 1, 1.7, 2.3, 
    2.5, 1.9, 2.9, 2.9, 0.6, 1.7, 2, 6.1, 7.1, 7.7, 7.1, 6.3, 4.1, 2.5, 5.2, 
    3, 5.9, 5.5, 5.4, 1.3, 3.5, 7.7, 3.2, 3.1, 3.5, 2.8, 0.7, 2.7, 2.8, 1, 
    0.2, 0.5, 0.6, 0.8, 1, 0.8, 1.7, 1, 1.1, 1.2, 1.2, 1.2, 0.3, 2.1, 1.6, 
    1.7, 1.2, 3.8, 8.4, 9.1, 10.5, 10.4, 12, 11.3, 12.7, 14.1, 16.6, 17.9, 
    16.3, 17.8, 17.1, 18.6, 18.7, 17.8, 15.9, 16.5, 15.5, 16.1, 13.8, 13, 
    13.1, 12.1, 11.6, 11, 9.4, 10, 10.7, 13.1, 12, 12, 11.1, 10, 8.5, 8.8, 9, 
    9.2, 8.8, 8.8, 9.1, 10, 9, 11.5, 12.1, 12.1, 13.3, 11.1, 10.3, 8.5, 10.1, 
    10.8, 9.6, 11, 11, 9.4, 8.5, 9.3, 6.3, 5.5, 5.8, 7.1, 6.8, 4.8, 5.6, 7.4, 
    6.4, 5.7, 4.9, 5.3, 3.2, 5.6, 3.8, 3.1, 5.1, 5.1, 3.4, 3.4, 1.9, 2.6, 
    5.5, 4.3, 4.6, 4.6, 3.8, 2.2, 3.6, 1.1, 4.6, 5.1, 3.3, 3.7, 2.6, 4.7, 
    4.3, 2.8, 1.7, 2.7, 2.7, 4.1, 7.1, 3.9, 2.3, 2.1, 0.6, 0.6, 1.7, 0.8, 
    0.5, 3.5, 1.2, 3.3, 1, 3.1, 1.3, 2.9, 2.1, 1.2, 4.5, 4.9, 2.3, 2, 1.4, 
    1.9, 1.1, 0.5, 1.4, 1.8, 6, 5.4, 5, 4.8, 5.7, 5.6, 5.4, 2.9, 2.4, 2.3, 
    1.7, 1.5, 0.4, 1.5, 1.4, 1.3, 1.4, 0.2, 1, 1.1, 1.3, 1.3, 1.5, 1.4, 2.1, 
    1, 0.4, 0.6, 0.6, 1, 0.7, 0.5, 0.3, 0.4, 1, 0.7, 0.9, 1.6, 2, 0.1, 0.7, 
    0.1, 0.9, 0.7, 1, 0.4, 0.7, 0.9, 1, 1.2, 0.9, 1.8, 0.5, 0.5, 0.1, 1.2, 
    1.3, 0.9, 1.2, 1.3, 1.5, 1.3, 2.9, 1.1, 3.6, 3.7, 3.8, 3.9, 5.2, 7.1, 
    8.6, 2.8, 5, 4.7, 5.6, 2.9, 0.6, 1.5, 1.4, 1.6, 1.3, 0.1, 1.3, 0.1, 0.8, 
    0.7, 1, 0.8, 0.7, 0.9, 1.2, 6.8, 7, 7.1, 7.3, 7.5, 6.4, 5.7, 5.6, 7.2, 
    5.3, 2.7, 3.8, 2.6, 1.9, 4.4, 6.5, 8, 8.1, 8.4, 7, 8.3, 8, 4.6, 4, 5, 
    5.4, 5.6, 5.3, 5.6, 3.2, 3, 2.6, 1.9, 1.5, 1.6, 0.6, 0.8, 1, 1.1, 0.7, 
    0.8, 0.4, 3, 3.3, 2.8, 3.5, 4.3, 5.1, 5.2, 5.9, 4.2, 5.5, 1.4, 3.4, 3.7, 
    1.2, 3.9, 5.8, 5.8, 6, 2, 7.4, 6.8, 7.1, 7.3, 6.8, 7.1, 7.5, 8.2, 8.7, 
    8.2, 7.6, 6, 5.5, 2.4, 2, 1.2, 2.1, 2.4, 2.2, 2.2, 2.9, 3.3, 2.4, 1.8, 
    2.8, 4.3, 2.2, 5.8, 4.2, 4.1, 4.3, 4, 3.9, 3.8, 3.7, 5.6, 5.3, 5.3, 3.4, 
    4, 4.4, 4.3, 5.2, 4.5, 0.9, 0.7, 1.3, 1, 0, 1, 0.3, 0.1, 0.2, 0.5, 0.9, 
    1.2, 0.8, 1, 1.2, 0.2, 0.4, 0.4, 0.7, 0.3, 2, 0.8, 2, 0.6, 0.6, 0.1, 2, 
    4.9, 2.5, 0.9, 1.1, 0, 0.5, 0.6, 0.7, 0.3, 0.4, 0.7, 0.8, 1, 1.1, 0.6, 
    1.4, 1.6, 0.6, 1.9, 3.1, 2.7, 1.3, 0.7, 0.7, 1.3, 1.7, 0.3, 1.4, 1.1, 
    0.7, 1.2, 0.7, 0.9, 0.8, 0.8, 0.9, 0.2, 0.4, 0.5, 1.1, 1, 0.2, 0.4, 1.4, 
    0.8, 0.8, 1.5, 1.8, 1.1, 1.1, 1.7, 2, 1.9, 1.9, 1, 1, 1.7, 1.7, 2.1, 1.2, 
    2.6, 0.8, 1, 1.3, 1, 1.4, 1.1, 0.9, 1.6, 0.2, 0.4, 0.5, 1.1, 0.2, 0.4, 
    0.2, 0.4, 0.6, 0.1, 1, 0.7, 0.3, 0.5, 1.1, 0.9, 0.3, 1, 2.1, 3, 1.1, 1.4, 
    1.2, 1.4, 0.9, 0.3, 1.2, 1.2, 1.5, 0.8, 0.2, 0.4, 1.5, 1.9, 1.8, 0.8, 
    0.4, 2.1, 2.6, 2.6, 2.7, 0.7, 1.1, 6.1, 3.4, 7.6, 4.1, 5.7, 7.1, 4.8, 
    4.5, 4.9, 3.4, 8.6, 9.1, 9.9, 10.3, 11, 11.5, 7.2, 8.1, 7.2, 10.3, 9.7, 
    6.1, 6.1, 5.8, 6.5, 7.3, 6.8, 7.3, 7.1, 6.9, 8.1, 4.2, 3.5, 1.4, 0.2, 
    0.6, 1.7, 0.3, 2.3, 0.5, 1.2, 2.6, 1.5, 0.1, 2, 2.1, 2.3, 6.1, 1, 1.5, 
    4.1, 0.3, 1.2, 0.4, 2.8, 1.5, 3.1, 2.9, 3.4, 1.4, 1.4, 1.3, 1.9, 2.7, 
    1.6, 2.1, 1.3, 1.8, 1, 1, 1.8, 3.6, 3.4, 5.2, 3.8, 4, 3.9, 3.3, 3.7, 2.5, 
    2.9, 2.9, 1.7, 3.8, 1.1, 4, 2.3, 2.3, 5.1, 1.6, 4.7, 4.3, 2.3, 2.5, 4.7, 
    5.7, 5.9, 7.2, 6.5, 6.5, 4.1, 0.6, 2.3, 1.1, 4.4, 5.1, 5.2, 5.1, 4.7, 
    2.7, 4.6, 4.2, 2, 3.4, 3.4, 1.9, 6.7, 2.7, 2.1, 2, 4, 6.3, 6.1, 8.3, 6.4, 
    6.9, 4.1, 2, 1.2, 0.5, 1, 1.2, 1, 3.3, 1.1, 1, 0.2, 1.7, 0.5, 0.5, 0.2, 
    0.7, 0.3, 1, 0.2, 0.6, 0.3, 0.3, 0.6, 0.3, 2, 1, 1.3, 0.7, 0.8, 0.2, 0.2, 
    0.9, 1, 1.4, 0.8, 0.7, 1.2, 0.4, 0.6, 0.6, 0.8, 0.4, 0.6, 0.2, 1.4, 0.8, 
    1.1, 0.6, 0.5, 0, 1.1, 2, 0.3, 0.4, 0.6, 0.4, 0.2, 0.1, 0.7, 0.5, 2.2, 
    1.1, 1.1, 0.3, 0.7, 0.7, 1.1, 1.8, 1.1, 6.9, 7.2, 6.2, 7.7, 4.7, 5.1, 
    6.1, 10.4, 11.1, 11.8, 9.2, 10.9, 11.3, 10, 7.5, 7, 9.1, 9.5, 10, 8.3, 
    8.5, 8.7, 8.3, 8.1, 7.6, 5.9, 6.2, 8.7, 9.7, 10, 10.3, 10.2, 8.2, 6.3, 
    6.1, 6.1, 3.5, 5.6, 1.7, 1.6, 4.9, 1.4, 1.1, 1, 1.3, 2, 1.8, 1.6, 0.7, 
    1.3, 1.3, 1.2, 1.7, 1.4, 1.2, 0.4, 1.7, 1.9, 1.8, 0.9, 1.2, 1.5, 0.4, 
    1.1, 1.6, 2.8, 2.2, 2.1, 6.1, 5, 4.5, 3.5, 3.2, 2.3, 0.7, 1.4, 3, 3.4, 
    2.8, 0.7, 0.7, 1.2, 0.7, 2, 1.6, 2.2, 2, 1.5, 1.1, 0.5, 1.1, 1.9, 0.2, 
    0.3, 0.6, 1.1, 0, 0.5, 1.2, 1.5, 1.4, 0.5, 1.4, 0.4, 0.3, 0.6, 1.5, 0.3, 
    1, 2, 2.1, 1.8, 2.9, 6.5, 6.7, 3.5, 6.2, 3.7, 3.4, 2.9, 1.6, 2.9, 1.4, 
    1.2, 1.7, 2.3, 0.9, 1.2, 1.2, 0.9, 0.8, 3.2, 2.9, 0.4, 1.2, 0.9, 2.1, 
    2.1, 2, 3.3, 5.2, 7.4, 6.3, 6.3, 3.2, 2.2, 2.1, 5.2, 8.2, 7.1, 8.8, 10.6, 
    7.5, 8.8, 8.8, 1.9, 2.3, 2.5, 2.2, 4.1, 4.6, 7.2, 1.1, 1.2, 0.9, 0.8, 
    1.1, 1.9, 1.3, 0.4, 2.3, 1.8, 0.9, 0.6, 0.7, 1.4, 1.3, 0.6, 1.2, 1.8, 
    0.2, 0.8, 1.3, 3.1, 1.2, 1.2, 1.1, 0.2, 2.3, 1.1, 0.4, 1.5, 1.3, 1.1, 
    0.9, 0.8, 1, 1, 0.4, 1, 0.6, 1.2, 1.3, 0.4, 1.7, 2.4, 0.4, 1.2, 1.1, 1.5, 
    1.9, 0.9, 0.6, 1, 0.7, 0.3, 0.8, 0.9, 0.9, 1.2, 0.4, 1.3, 0.5, 0.7, 0.9, 
    1, 1.1, 1.4, 1.3, 0.6, 1, 1.1, 1.3, 1.5, 1, 1.1, 1.3, 0.9, 2.7, 2.5, 2.7, 
    2.8, 2.4, 1, 1.1, 0.4, 0.4, 0.2, 4.7, 3.3, 0.6, 1.4, 0.4, 0.2, 1.1, 0.4, 
    0.3, 0.5, 0.7, 0.8, 0.8, 0.7, 0.2, 1.2, 0.5, 0.7, 1.1, 0.3, 0, 0, 0.4, 
    0.2, 0.8, 1.1, 2, 5.9, 3.8, 4.2, 6, 6, 6.4, 5.5, 5.7, 4.6, 4.7, 2.4, 3.2, 
    5, 4.5, 4.4, 4.5, 4.4, 5, 4.7, 5.2, 5.3, 5.2, 4.6, 1.1, 0.9, 6.4, 4.9, 
    3.4, 3.6, 4.1, 4.2, 4.9, 5, 5.4, 5.1, 4, 5, 7.4, 6.5, 5.3, 6.5, 7.2, 6.9, 
    7.8, 7.2, 7.7, 6.8, 8.3, 6, 6.3, 5.8, 7.2, 6.7, 5.3, 5.5, 4.9, 5.4, 5.5, 
    3.3, 2.1, 1.4, 6.4, 7.1, 6, 3.3, 4.6, 3.8, 4.8, 4.3, 5.5, 5.9, 4.3, 4.1, 
    4, 3.8, 4.1, 4.4, 3.9, 3.2, 4.3, 5.7, 5.6, 4.7, 4.4, 5.2, 4.4, 2.6, 4.8, 
    3.6, 4.2, 4.1, 3.6, 6.1, 5.4, 4.1, 5.3, 4.8, 4, 4.4, 5, 3.5, 3.1, 3.8, 
    3.8, 4.5, 4.2, 4.5, 4.2, 3.5, 2.6, 2.8, 2.1, 3.4, 3.6, 2.4, 1.3, 2.5, 
    3.3, 4.1, 3.5, 4.1, 3.7, 6.7, 5.6, 3.3, 3.6, 3.9, 4.2, 3.6, 3, 3.6, 1.1, 
    4.6, 8.2, 5.9, 9.7, 9.8, 8.9, 7.2, 8, 5.9, 7.5, 6.5, 3, 6.4, 6.6, 7.5, 
    7.5, 6.8, 4.8, 6.9, 3, 5.2, 5.6, 5.3, 4.2, 4.2, 5.9, 5.1, 4.7, 2.3, 5.3, 
    3, 1.6, 1.8, 2.9, 0.7, 1.7, 3.9, 3.9, 4.9, 6.1, 8.1, 8.8, 9.6, 3.2, 2.4, 
    7.2, 4.2, 2.2, 6.4, 6.1, 6, 2.9, 1.9, 7.4, 0.3, 1.1, 0.4, 0.6, 6.3, 6.1, 
    6.4, 7.6, 6.8, 6.8, 8.3, 9.2, 8.7, 9.1, 9, 7.9, 6, 7.6, 5.5, 8.4, 2.3, 
    1.9, 3.5, 2.3, 1.7, 1.5, 0.7, 0.2, 2.1, 2.4, 4.1, 3.7, 1.9, 2.3, 2.5, 
    2.8, 2, 2.9, 2.5, 1.5, 1.9, 2.4, 1.9, 2.4, 0.1, 1.9, 0.7, 1.5, 1, 0.8, 
    0.3, 0.6, 0.8, 0.1, 0.6, 1.1, 3.2, 4, 5.1, 8.5, 8.5, 9.1, 9.3, 10.2, 9.9, 
    9.7, 9.8, 9.9, 8.6, 9.6, 6.8, 6.2, 3.8, 3.3, 4.5, 3.1, 2.9, 1.3, 3.1, 
    2.5, 3.6, 2.2, 1.6, 2.3, 2, 2.2, 2.2, 3.6, 3.5, 2.4, 0.8, 1.6, 1.7, 1, 
    1.1, 0.7, 0.8, 0.8, 2.4, 2.3, 1, 1.1, 1.3, 1.6, 0.6, 0.8, 0.8, 1.8, 1.1, 
    0.5, 0.9, 0.8, 0.4, 1.6, 0.1, 0.6, 0.9, 0.3, 1.6, 1.5, 2, 1.2, 1.4, 1.4, 
    1.3, 1.5, 1.3, 2.3, 1.1, 1.4, 1, 3, 0.9, 1.4, 1.9, 2.2, 2.1, 1.3, 1.7, 
    0.3, 0.5, 0.5, 0, 1, 0.2, 1, 0.3, 0.4, 0.6, 4, 4.3, 5.6, 6.2, 5.7, 6.2, 
    8.5, 12, 11.1, 9.4, 10.3, 3.7, 4.2, 6.9, 8.1, 8.1, 9, 6.4, 9.5, 7.6, 3.6, 
    0.9, 2.3, 2, 2, 1.8, 2, 2.3, 8.8, 10.7, 10.3, 10.8, 9.8, 9.1, 8.4, 8.8, 
    8.6, 6.9, 7.9, 12.7, 12, 11, 10.2, 13.1, 15.3, 15.3, 16.2, 16, 15, 15.8, 
    12.1, 11.9, 11.8, 11.7, 11.5, 8, 6.2, 5.5, 5.6, 7.1, 7.3, 6.4, 9.5, 6.5, 
    7.7, 5.5, 6.4, 4.3, 1.9, 4.1, 0.7, 1.6, 2.5, 1.8, 4, 3.2, 3.7, 3.2, 2.2, 
    3.1, 8.9, 6.7, 6.5, 1.4, 4, 1.6, 1.3, 1.6, 2.3, 2.8, 3.3, 1.8, 3.8, 3, 
    2.4, 2, 2.9, 2.9, 3, 5, 5.8, 6.9, 3.5, 3, 5.7, 4.5, 2.5, 1.6, 2.9, 2.6, 
    3.2, 4.5, 3.8, 3.6, 2.3, 3.3, 1.6, 4.1, 4.6, 6, 6, 9, 10.8, 9.7, 6.8, 
    6.3, 6.1, 4.6, 4.5, 1.6, 3.4, 2.9, 1.4, 1.4, 1, 1.3, 1.9, 1.6, 1.8, 0.9, 
    1.3, 1.4, 2.1, 2.3, 0.7, 0.7, 1.1, 2.3, 1.1, 0.8, 1.2, 0.8, 0.5, 1.2, 
    1.2, 1.1, 1.3, 1.1, 0.2, 1.4, 0.4, 1.3, 1.5, 0.8, 0.5, 0.8, 0.7, 0.8, 
    1.5, 0.4, 0.2, 0.2, 1, 1, 1.9, 1.1, 0.6, 0.5, 0.6, 0.6, 0.7, 0.5, 1.2, 
    0.7, 1.5, 0.6, 0.2, 0.8, 0.2, 0.5, 0.5, 1.5, 0.9, 1.7, 1.3, 1, 2.7, 0.6, 
    0.8, 0.6, 0.6, 0.7, 0.4, 0.6, 0.4, 1.3, 0.4, 0.3, 0.9, 0.1, 1, 0.3, 1, 
    1.5, 0.5, 0.5, 0.1, 0.3, 0.4, 0.4, 0.9, 0.3, 0.7, 0, 0.2, 0.5, 0.1, 0.4, 
    0.4, 1, 0.1, 0.4, 0.2, 0.8, 0.4, 0.7, 1.3, 0.5, 2.6, 1.5, 1, 0.2, 0.1, 
    0.1, 0.2, 0.2, 0, 0.3, 0.4, 1.1, 0.3, 0.1, 0.2, 0.1, 0.2, 0.6, 0.4, 0.7, 
    0.6, 0.4, 0.4, 0.7, 1.2, 0.9, 0.9, 0.2, 0.6, 0.4, 0.9, 0, 0, 0, 0.3, 0.9, 
    0.4, 0.1, 0.3, 0.6, 0.6, 0.2, 0.1, 0.3, 0.2, 1, 0.9, 0.3, 0.7, 0.7, 0.6, 
    0.4, 0, 0.7, 1, 1, 1.1, 0.5, 0.3, 0.2, 0.2, 0.4, 0, 0.3, 1.8, 1.8, 2.4, 
    1, 1.3, 1.5, 3.5, 1.5, 0.6, 1, 0.4, 0, 1.1, 1.2, 0.5, 0.3, 0, 1.1, 1, 
    0.6, 0.6, 0.9, 0.6, 0.5, 0.4, 0.7, 1.2, 1.6, 0.3, 0.3, 0.9, 0, 0.1, 0.9, 
    0.8, 0.3, 0.3, 2.3, 3.4, 3.1, 3, 1.2, 2.1, 5.2, 5.1, 2.5, 2.9, 1.3, 1.9, 
    2.9, 0.8, 1.6, 1.6, 1, 1, 0.8, 1.1, 0.5, 0, 0.9, 0.3, 1, 1.1, 0.9, 0.8, 
    3.5, 2, 1.9, 0.2, 0.4, 1, 0.6, 0.8, 0.7, 0.8, 0.5, 0.6, 0.6, 1.2, 0, 0.1, 
    1.3, 0.1, 0.9, 0.8, 0.6, 0.6, 0.1, 0, 0.1, 0, 1, 0.3, _, _, _, _, _, _, 
    _, _, _, _, _, _, 1.1, 4.8, 3.4, 4.2, 4.7, 3.5, 2.8, 4.6, 6.7, 7.8, 9.6, 
    5, 4.2, 5.6, 1.2, 0.8, 1.4, 2.4, 3.3, 5.1, 4.7, 4.6, 4.4, 4.9, 4.2, 5.1, 
    4.8, 3.8, 4, 4.2, 3.3, 3.5, 1, 0.9, 0.7, 1, 0.3, 1.1, 0.8, 1.3, 1.5, 2.2, 
    0.6, 1, 0.7, 1.3, 0, 1.2, 0, 6.1, 1, 1, 0.8, 0.9, 7.4, 11.6, 7.8, 7, 6.8, 
    3, 1.7, 2.1, 1.9, 1.9, 4.4, 3.7, 5.3, 6.3, 5, 2.6, 4.8, 3.5, 0.6, 4.6, 6, 
    5.4, 3.7, 7, 7.7, 7.5, 7.1, 2.5, 2, 4.7, 1.5, 4.5, 1.8, 1.7, 0.5, 2, 1.8, 
    3.2, 8, 8, 7.5, 1.7, 0.8, 2.1, 2.4, 1.6, 1.6, 0.7, 1.5, 0.3, 1.1, 1.7, 
    1.2, 0.2, 0.8, 0.7, 1.5, 1, 2, 3.4, 2.8, 1.1, 0.5, 0.4, 1.2, 0.1, 1.2, 
    0.4, 0.7, 0.6, 0.6, 0.4, 0.9, 0.6, 0.5, 1, 0.3, 0, 0.4, 0.1, 0.1, 0.2, 0, 
    0.7, 0.5, 0.8, 0.4, 2.6, 0.4, 0.9, 0.8, 0.5, 0.3, 2, 1.1, 1.5, 2.3, 1.9, 
    1.8, 1.2, 0.7, 0.3, 1.3, 1, 0.7, 0.6, 1.4, 0.7, 0.4, 0.1, 0.6, 0.6, 0.7, 
    1.1, 1.7, 0.8, 1.6, 1.3, 1.3, 1.1, 0.8, 3, 1.8, 1.3, 1.8, 2.4, 2.2, 4, 
    2.6, 4.4, 6.3, 6.3, 7, 11, 10.1, 10.9, 11.1, 11.7, 11.8, 11, 10.5, 10.1, 
    10.1, 10.3, 11.4, 12.6, 11.5, 12, 13.1, 11.9, 12.1, 12.2, 12.8, 12.9, 
    11.9, 13.1, 13, 13.3, 11.2, 12.2, 13.1, 10.7, 10.5, 10.1, 10.1, 10.4, 
    8.1, 9.8, 10.2, 9.3, 8.1, 8.9, 5.6, 8, 7.6, 5.5, 6.8, 6.3, 3.7, 2.4, 1.4, 
    4.7, 2, 3, 0.5, 1.3, 0.6, 0.7, 0.8, 1.8, 0.8, 0.6, 2.4, 1, 1.2, 0.4, 0, 
    0.6, 0.6, 0.1, 0.8, 0.5, 0, 0.1, 0, 0, 0.2, 0.1, 0.5, 0.3, 0.3, 0.6, 0.3, 
    0.5, 0.5, 0, 0.9, 0.8, 0.6, 1.1, 0.7, 0.8, 0.2, 0, 0.4, 2.9, 1.2, 1.8, 
    1.4, 1.1, 1.1, 1.7, 0.6, 0.1, 0.5, 0.6, 0.6, 0.3, 0.1, 0.9, 0.2, 1.1, 
    1.3, 1, 0.1, 0.5, 0, 0.1, 0.7, 1.2, 0.2, 0.6, 0.4, 0.8, 0.3, 1, 0.2, 0.4, 
    0.2, 1, 0.5, 0.5, 0.4, 0, 0.4, 0.1, 0, 0.2, 1, 0.3, 0.5, 0.1, 0.5, 1, 
    0.7, 0.1, 0.5, 0.7, 0.4, 0.5, 0.4, 1, 0.4, 0.9, 1.2, 1, 0.5, 0.5, 0.5, 
    0.2, 0.1, 0.1, 0.5, 0.7, 4.1, 1, 1.8, 6.6, 2.6, 1.3, 1.5, 1.5, 0.4, 0.2, 
    0.9, 1.4, 0.7, 0.7, 0.6, 0.2, 1.2, 0.7, 0.7, 0.8, 0.7, 0.6, 3.4, 4.1, 
    6.6, 7.4, 5.9, 4.5, 4.4, 3.3, 3.7, 4.4, 3.9, 3.1, 0.8, 0.8, 0.1, 0.7, 
    0.7, 0.3, 0.3, 0.5, 0.4, 0.6, 0.4, 0, 0.8, 0.7, 1.7, 1.4, 2.1, 1.6, 1, 
    0.7, 0.8, 0.6, 0.6, 0.9, 0.8, 0.8, 0.6, 1.1, 0.4, 0.5, 0.2, 0.3, 0.7, 
    0.3, 0.5, 0.4, 1.8, 4.3, 5.1, 5.6, 4.7, 5.6, 7.6, 7.1, 7.8, 5.9, 6, 6.1, 
    5.9, 7.1, 6, 5.6, 7, 7.4, 10.3, 5.9, 2.9, 5.6, 5.1, 3.1, 2.4, 2.8, 1.7, 
    2, 1.3, 2.2, 2.7, 11.4, 2.6, 5.6, 3, 2.6, 2.6, 1.4, 2.7, 1.2, 1.7, 2, 
    6.6, 10.5, 8, 5, 3.4, 2.8, 2.9, 4.9, 4.2, 6.5, 2.6, 2.6, 2.4, 4.1, 5.1, 
    2.3, 5.3, 7.6, 3.4, 2.4, 2.8, 5.1, 4.8, 10, 10.5, 9.1, 4.1, 3.7, 2.2, 
    2.7, 6.6, 6.2, 2.9, 3.4, 5.1, 2.9, 2, 1.6, 1.4, 1.3, 0.1, 0.6, 0.9, 0.9, 
    1.5, 0.7, 1.7, 2.2, 1.4, 0.8, 2.2, 1.6, 1.5, 1.1, 0.2, 1, 2.2, 0.5, 0.7, 
    2.9, 1.2, 0.5, 1.5, 1.2, 0, 0.3, 0.2, 0.4, 0.9, 0.5, 0.2, 1.1, 0.7, 0.7, 
    1, 1.4, 0.3, 0.1, 0.3, 0.8, 0.9, 0.6, 0.6, 1.6, 3.4, 0.7, 0.4, 0.1, 0, 
    0.1, 0.4, 0.1, 0.4, 0.2, 0.3, 1.1, 0, 0.1, 0.3, 1.5, 0.9, 1.6, 1.5, 1.2, 
    1.5, 0.8, 1.3, 1.3, 1.5, 1.2, 1.9, 0.5, 0.4, 1, 0.9, 0.8, 0.3, 1.3, 1, 1, 
    0.9, 0.3, 1.7, 1.4, 2.7, 2.2, 1.1, 1, 0.7, 1.6, 0.9, 1.1, 0.3, 0.6, 1.1, 
    0.5, 0.2, 0.2, 0.7, 0.1, 0.5, 0.8, 0.4, 0.7, 0, 1.4, 0.7, 0.3, 0.8, 0.6, 
    0.8, 0.8, 0.6, 0.2, 0.4, 0.3, 0.3, 0.8, 0.1, 0.5, 0, 0.6, 0.3, 0.5, 0.1, 
    0.7, 0.8, 0.7, 1.5, 0.9, 2, 0.9, 1.8, 2.7, 1.6, 5.3, 8.2, 5.9, 2.7, 3.4, 
    2.5, 2.6, 1.8, 1.1, 0.5, 1.3, 0.6, 0.9, 0.7, 0.7, 0.8, 0.9, 1.2, 1.1, 
    0.2, 1, 1, 0.8, 1.1, 1.1, 1.4, 0.6, 1.1, 1.1, 0.6, 0.5, 1.3, 0.9, 1.1, 
    1.5, 0.8, 0.8, 0.6, 1, 3.4, 6.6, 6.5, 3.5, 2.6, 4.4, 7, 3.9, 3.9, 3.4, 
    6.1, 4, 5.2, 4.8, 1.8, 1.2, 1.8, 1.3, 1.6, 1.9, 1.6, 1, 0.9, 2, 2.1, 2.3, 
    0.6, 1.6, 2.6, 3.2, 0.8, 2.1, 2.5, 1.5, 1.6, 1.7, 1.4, 1.3, 1.2, 1.1, 
    0.6, 1.1, 1, 1.1, 0.9, 1, 1, 1.1, 1.3, 0.9, 1.5, 0.3, 1.5, 0.3, 0.5, 0.1, 
    1, 0.4, 0.8, 1.2, 0.4, 0.7, 0, 0.7, 0.2, 0.1, 0.7, 0.2, 0.3, 0.5, 0.5, 0, 
    0.2, 0.4, 0.8, 0.3, 0, 0.2, 0.1, 0.2, 0.8, 0.3, 0.7, 0, 1, 1.8, 0.1, 0.2, 
    0.9, 1.1, 0.6, 5.5, 5, 1.4, 0.2, 1.1, 1.1, 0.5, 1.2, 0.6, 1, 3.6, 4.5, 
    4.4, 4.1, 4.8, 4.7, 5.9, 4.7, 5.8, 6.6, 6.8, 6.3, 6.5, 4.6, 5.4, 2.7, 
    4.3, 2.1, 0.4, 2.1, 2.8, 3.7, 3.7, 1.4, 2.5, 3.8, 1.2, 1.1, 1, 1.1, 1.3, 
    0.5, 0.7, 0.8, 1.5, 0.2, 0.2, 0.2, 0.5, 1.4, 1.1, 0.9, 0.7, 0.9, 1.2, 
    0.2, 0.5, 0.7, 0.4, 0, 1.1, 1.1, 0.7, 0.9, 1.1, 0.2, 0.1, 0.4, 0.4, 0.1, 
    0.6, 0.3, 0.5, 0.8, 0.9, 0.5, 0.8, 1.2, 0.4, 2.2, 0.9, 0.6, 0.2, 0.4, 
    0.1, 0.6, 0.9, 0.7, 0.1, 0.2, 0.4, 0.9, 0.1, 0, 0, 0, 0.6, 0.2, 0.5, 0.2, 
    0.7, 0.2, 0.1, 0, 0.9, 0.4, 0.5, 0, 0, 1.4, 0.3, 0.5, 0.3, 0.7, 0.9, 0.6, 
    0.4, 0.7, 0.9, 1.1, 0.3, 1.4, 1.5, 1.5, 1, 1.9, 1.4, 1.9, 2.2, 1.6, 1.8, 
    1.8, 1.1, 1, 0.7, 1.5, 0.8, 0.7, 0.2, 1.4, 1.5, 2.3, 0.5, 1, 0.7, 0.8, 
    0.9, 0.9, 0.8, 1.2, 0.8, 3, 2.6, 2, 1.7, 1.4, 1.9, 2.6, 2.7, 2.1, 2.8, 
    3.8, 1, 1.2, 0.9, 1.7, 1.9, 1.7, 1, 0.6, 1.2, 1.1, 0.4, 0.6, 0.8, 1.6, 1, 
    0.9, 4, 1.3, 3.2, 0.8, 0.3, 0.6, 0.3, 0.2, 0.5, 0.4, 0.1, 0.1, 0.3, 0, 
    0.3, 0.3, 0.9, 0.9, 1, 1, 0.2, 0, 0.1, 1.2, 0.7, 1.2, 1.5, 1, 1, 1.1, 
    0.7, 0.5, 1, 1.2, 3.7, 3.4, 1.3, 0.9, 1.2, 1, 1, 0.7, 1.4, 0.5, 3.1, 2.4, 
    2.1, 1.2, 2.1, 2.1, 2.5, 3, 2.1, 0.5, 0.8, 0.9, 0.8, 1, 0.6, 0.3, 0.1, 
    0.3, 0.2, 1.1, 0.4, 0.7, 0.8, 1, 0.1, 0.7, 2.5, 3.2, 3.5, 3.3, 2.5, 2.7, 
    2.4, 0.5, 1.2, 0.6, 0.5, 0.2, 0.4, 0.8, 1.2, 1.3, 0.7, 0.2, 0.3, 0.5, 
    1.1, 0.6, 0.5, 1.3, 1.3, 1.4, 2.4, 0.5, 1, 1, 1.5, 6.3, 5.4, 6.3, 4.9, 7, 
    6.1, 4.1, 6.6, 6, 5.1, 6, 6.9, 3.8, 4.2, 7.1, 4.2, 6.8, 6, 2.8, 3.6, 4.2, 
    4.3, 5.9, 7.2, 6.5, 4.6, 6.1, 10, 3.8, 1.3, 3.7, 1.9, 2.8, 2.3, 0.8, 1.3, 
    1.3, 1.3, 1.5, 4.2, 4.2, 2.5, 2, 2.1, 1.7, 2, 0.5, 1.9, 1.4, 0.9, 1.3, 
    0.3, 1.1, 2.5, 1.9, 1.4, 1.9, 2, 1.5, 1.5, 6.2, 5.3, 6.3, 2.3, 5.2, 7.5, 
    2.9, 2.2, 2.4, 3.3, 1.8, 4.4, 1.8, 1.7, 3, 0.5, 0.4, 0.7, 2.1, 0.9, 0.9, 
    0.9, 0.9, 0.9, 0.3, 1.2, 1, 1.1, 1.6, 0.2, 1.1, 1.3, 1.6, 1.5, 2.1, 1.2, 
    2.7, 2.1, 0.9, 0.4, 0, 0.2, 0, 0.2, 0.6, 0.5, 0, 0, 0, 0.1, 0.5, 0.3, 
    0.3, 0.3, 0.6, 0.4, 1.1, 0.8, 1, 1.3, 1.5, 1, 0.8, 0, 0.2, 0.2, 0, 0, 
    0.5, 0.5, 0.6, 0.2, 0.3, 0.6, 1, 2.2, 2.8, 3, 2.3, 1.4, 2.4, 1.5, 0.7, 
    1.5, 0.8, 1.4, 0.7, 0.7, 0.9, 1.5, 0.1, 0.8, 4, 4.4, 4.3, 4.3, 3.7, 3.5, 
    1.2, 0.9, 1.5, 0.3, 0.7, 0.4, 0.6, 0.2, 0.8, 0.2, 0.4, 0.8, 0.1, 0.9, 
    0.3, 0.6, 1, 1.2, 1.4, 4.2, 7.7, 4.5, 4.3, 0.3, 4, 4.1, 4.9, 8.8, 4.2, 5, 
    4.5, 5.2, 3.2, 1, 1.4, 0.2, 1.5, 1.7, 5.8, 6.5, 5.9, 7, 6.1, 5, 4.8, 4.2, 
    5.2, 4.4, 5.2, 5.5, 5, 4.2, 5.9, 5.3, 4.9, 1.8, 2.2, 1.7, 1.7, 1.7, 1.5, 
    2.2, 2.4, 2.2, 0, 0.9, 0.2, 0.5, 0.5, 0.8, 4.3, 2.7, 3.1, 3, 2.8, 1.4, 
    1.7, 1.9, 1, 0.6, 2.4, 2.4, 2, 0.8, 2.5, 2.8, 0.6, 1.3, 1.2, 2, 3.3, 2.8, 
    1.3, 1.1, 1.1, 0.4, 1, 1.3, 1.3, 0.5, 1.4, 1.8, 1.3, 1.3, 0.7, 1.8, 0.2, 
    0, 0.4, 0, 1.2, 0.7, 1.1, 0.7, 0.6, 0.7, 0.5, 0.5, 1, 0.9, 0.7, 1, 0.6, 
    1.6, 1, 1, 1.2, 1.4, 1.2, 1.3, 1, 1, 0.8, 0.6, 0.8, 0.6, 0.4, 1, 0.7, 
    0.6, 3.1, 3.1, 2.9, 2.1, 1.3, 2, 1.1, 1.8, 2.1, 2.1, 1.1, 0.3, 1.4, 1.1, 
    1.4, 2.9, 4.1, 1.4, 0.7, 0.6, 0.8, 0.6, 0.4, 0.9, 1.3, 0.2, 0.9, 0.2, 
    1.2, 1.1, 1.1, 1.6, 1.4, 2.2, 4, 2.4, 5.8, 5, 1.7, 8.4, 5.2, 4.5, 1.6, 1, 
    3.1, 3.6, 1.3, 1.5, 1.9, 2, 2.1, 2.3, 3.4, 2.9, 2.9, 3, 2.4, 1.9, 2.6, 
    8.2, 7.9, 4.8, 3.1, 3.3, 1.9, 0.3, 0.4, 0.9, 0.6, 0.8, 2.2, 0.8, 3, 4.5, 
    2.1, 2.9, 3.4, 3.5, 5.5, 8.2, 8.3, 9.9, 7.5, 1.8, 3.5, 2.5, 2.9, 2.8, 
    8.4, 7, 7.3, 1.2, 0.9, 5.5, 1.5, 5.2, 7.4, 1.3, 1.5, 3.6, 3.2, 1.9, 1.5, 
    4.5, 2.5, 1.4, 2.5, 1.6, 1.4, 2.5, 1.3, 2, 2.6, 3, 3.1, 0.5, 1, 0.8, 0.7, 
    1.9, 3.1, 3, 2.6, 2, 1.9, 2.8, 2.7, 2.7, 1.7, 3.7, 3.8, 6.5, 1.7, 3.3, 
    5.4, 1.7, 2.9, 4.3, 0.7, 3.2, 1, 2.1, 0.4, 0.8, 1, 1.1, 1.1, 1.4, 1.6, 
    1.2, 1, 1.7, 1, 1.4, 1.7, 1.8, 1.7, 1.3, 1.1, 1.5, 1.7, 1.2, 1, 1.1, 1.5, 
    1.1, 0.6, 1.4, 2.7, 2.4, 2.4, 1.7, 2, 2.8, 2, 1.7, 1.1, 0.7, 1.7, 1.1, 
    0.8, 1.1, 1, 1.5, 2.3, 0.6, 0.3, 0.5, 0.6, 0.4, 0.1, 0.8, 1, 1, 0.9, 0.4, 
    0.9, 0.9, 1.5, 1.3, 1.1, 2.2, 2, 2.7, 3.5, 3.5, 3.6, 3.5, 3.1, 2.8, 2.9, 
    2.2, 0.7, 0.5, 0.2, 0.5, 0.5, 1, 1.1, 1.4, 1.3, 1.1, 1, 1.2, 1, 1.5, 1.3, 
    1.1, 1.2, 1.2, 0.9, 1.4, 1.4, 2, 1.8, 1.4, 1.7, 1.2, 1, 0.3, 0, 1.8, 0.7, 
    0.6, 0.7, 0.3, 0.9, 2.2, 1.4, 1.2, 0.9, 0.6, 1, 0.6, 0.3, 0.4, 1.6, 0.6, 
    1.6, 0.1, 1.3, 0.9, 0.3, 0.2, 0.4, 0.6, 1, 1.3, 1.3, 2.6, 2.6, 2.7, 1.1, 
    1, 0.8, 0.8, 0.4, 0.9, 1.1, 1.7, 0.3, 2.2, 2, 0.9, 1.9, 1.2, 0.8, 4.3, 
    4.1, 4.3, 4.7, 3.8, 4.6, 4.6, 5.7, 4.6, 5.6, 5.1, 4.4, 3.6, 1.6, 1.2, 
    1.2, 2.5, 1.8, 0.9, 1.3, 1.1, 0.3, 0.3, 0.1, 0.1, 0.3, 0.3, 1.6, 0.7, 
    0.9, 3.2, 2.3, 1.5, 1.5, 1, 1.5, 2.2, 2.6, 0.8, 1.4, 1.4, 1, 1.2, 1.7, 
    0.6, 0.8, 1.2, 1.3, 1, 0.7, 1.5, 0.4, 1.2, 2.6, 4.9, 4.1, 1.3, 2.1, 1.2, 
    1.6, 1.7, 1.6, 1.3, 1.6, 0.7, 0.7, 0.8, 1.6, 1.2, 0.7, 0.9, 1.1, 1.4, 
    1.5, 1.8, 1.9, 1.7, 2.2, 2.4, 2.5, 1.5, 1.4, 1.1, 1.4, 1.1, 1.2, 1, 0.8, 
    1.6, 2.5, 1.6, 1.8, 1.1, 0.4, 0.5, 0.6, 0.6, 0.2, 1.2, 1.8, 2.3, 2.2, 
    1.4, 1.6, 1.7, 1.2, 1.2, 1.2, 1.4, 0.9, 0.9, 0.7, 0.2, 1.1, 0.9, 0.7, 
    0.9, 1.6, 0.8, 0, 0.9, 3.8, 2.6, 1.5, 0.9, 2.8, 0.9, 1.1, 1, 1.4, 1, 1.2, 
    0.6, 1.7, 2.3, 2.4, 2.5, 1.7, 1.4, 0.9, 0.8, 0.4, 0, 0.2, 0.4, 0.5, 0.5, 
    0.3, 0.2, 0.3, 0.4, 0.7, 0.1, 0.9, 0.4, 0, 1.3, 2.1, 1.5, 0.4, 0.2, 1.2, 
    1.7, 1.2, 1.8, 2.6, 1.5, 1.7, 1.8, 1.7, 3.6, 4.7, 3.5, 6.1, 6.1, 5.4, 
    3.5, 7.2, 6.3, 10.3, 3.9, 4.3, 7.3, 1.6, 5.6, 4.7, 3.3, 3, 1.1, 0.8, 0.7, 
    0.4, 1, 1.6, 2, 2.7, 5.3, 2.7, 5.9, 5.3, 5.7, 3.8, 5.7, 3, 3.1, 2.5, 5.2, 
    3.5, 1.4, 1.9, 3.8, 3, 1.6, 1.8, 1.8, 1, 1.6, 1.6, 2.4, 1.9, 0.7, 1.7, 
    1.5, 1.6, 1.9, 2, 1.5, 1.5, 1.8, 1.7, 1.6, 3.5, 2.1, 6, 1.3, 1.2, 0.3, 
    1.6, 2.1, 1.7, 1.5, 1.2, 2.8, 2.6, 2.4, 2.5, 2.8, 1.8, 3.1, 3.3, 1.4, 
    1.8, 1.3, 1.3, 1, 1.5, 0.7, 1.1, 1.6, 1.1, 1.2, 1.6, 1.9, 1.2, 0.9, 1.1, 
    1.3, 1.5, 1.2, 0.8, 1.7, 1.5, 1, 1.3, 4.8, 4.7, 4.2, 4.5, 4.7, 2.8, 0.9, 
    2.2, 1.4, 1.3, 1.5, 2, 0.9, 2.4, 0.4, 1.5, 1.5, 1.7, 1.4, 2.4, 2.3, 2.1, 
    1.4, 1.2, 1.7, 1.5, 1.7, 1.3, 1.2, 1.9, 1.8, 0.4, 2.1, 0.7, 1.5, 1.2, 
    1.2, 1.5, 1.9, 1.5, 1.3, 1.8, 1.3, 1.8, 2.1, 1.6, 3.2, 3.3, 2.4, 3.1, 
    2.4, 2.3, 1.6, 3, 3.5, 3.2, 3.2, 2.1, 1.2, 1.8, 2.6, 1.6, 2.1, 1.8, 1.8, 
    1.5, 4.8, 4.8, 2.4, 2.1, 2.8, 3.3, 3.4, 9, 8.5, 6.1, 3.6, 6, 3, 3.6, 2.3, 
    3.5, 4.9, 6.9, 2.7, 2.7, 2.4, 2.6, 1.5, 2, 4.4, 3.4, 2.5, 2.9, 4.9, 4.3, 
    6.9, 4.8, 7.5, 3.7, 3.3, 4.8, 5.2, 2.5, 3.2, 3.6, 2.7, 5, 5.1, 3.2, 3.5, 
    6, 3.8, 3.6, 2, 3.9, 3.6, 4.7, 1.1, 1, 2.2, 2.1, 4.4, 2.9, 3.2, 4.3, 2.9, 
    3.9, 2.1, 1.8, 1.2, 1.5, 0.6, 0.8, 1.8, 2.1, 2.1, 2.9, 1.5, 1.2, 2.6, 
    2.2, 1.4, 1.6, 1.4, 1.6, 1.9, 1.9, 2, 1.2, 1.3, 1.2, 1, 0, 0, 1, 0.4, 
    0.5, 0.1, 0.5, 0.4, 1.1, 1.9, 1.5, 2.4, 2.5, 1.9, 1.6, 1.7, 1.9, 1.7, 
    2.2, 2.1, 2.4, 1.8, 1.8, 2.2, 1.4, 2.4, 2.1, 1.1, 1.2, 1.4, 0.9, 0.6, 
    0.6, 1.3, 1.8, 1.1, 1.5, 1.1, 1.4, 2.7, 2.1, 2.6, 3.1, 3.1, 2.6, 1.8, 
    2.6, 1.4, 1.7, 1.4, 0.5, 1.1, 1.8, 1.2, 1.6, 1.6, 1.5, 0.2, 1.3, 1.2, 
    1.9, 1.7, 1.7, 1.5, 2, 2.3, 0.7, 1.2, 1, 2.1, 0.2, 0.8, 0.7, 0.7, 0.3, 
    0.1, 0.9, 0.9, 0.6, 1.5, 1, 1.1, 2.2, 1.1, 1.9, 1, 0.8, 1.5, 0.6, 0.5, 
    1.1, 1, 2.2, 1.1, 1.2, 0.1, 0.8, 0.6, 0.1, 0.2, 0.3, 0.8, 0.8, 0.7, 0.5, 
    1.2, 4.6, 2.6, 4, 3.4, 3.8, 1.8, 3.3, 4.1, 3.1, 0.5, 1.6, 1.4, 2.4, 3.2, 
    2.9, 1.3, 0.1, 1.1, 2.9, 1.8, 1.2, 0.2, 0.4, 0.4, 0.7, 1.8, 1.6, 1, 1, 
    1.3, 1.9, 1.4, 2.4, 2.1, 1.7, 1.4, 1.7, 1.7, 1, 1, 1.1, 0.3, 0.5, 0, 0.9, 
    0.1, 0.1, 0.7, 0.6, 1, 2.7, 3.2, 2.6, 1.2, 1.4, 1.2, 1.2, 1.8, 1, 0.9, 
    1.8, 0.6, 1.2, 0.3, 0.8, 0.7, 0.2, 0.2, 0.1, 0.3, 2.4, 1.9, 0.9, 0.8, 
    1.2, 2.4, 1.1, 1.5, 1.4, 1.4, 1.3, 1.7, 1.3, 0.8, 1.1, 1.3, 0.9, 0.4, 
    0.6, 1, 0.2, 1.1, 1, 0.2, 0.8, 0.1, 0.3, 0.8, 0.7, 0.9, 0.4, 1.2, 1.1, 
    0.3, 0, 0.1, 1.7, 0.7, 0.3, 1, 1.2, 0.4, 0.1, 0.1, 0.1, 0.8, 1.3, 0.8, 
    0.9, 1.2, 1.4, 1.4, 1.4, 1.9, 1.4, 1.5, 1.9, 0.8, 1.5, 1.6, 1, 1.2, 1.3, 
    1.3, 0.2, 0.7, 1.2, 0.6, 0, 0.4, 0.7, 0.8, 1, 1.6, 1.7, 2.1, 2.6, 1.8, 
    1.6, 1.9, 1.3, 2.9, 2.7, 1.7, 2.5, 1.7, 0.9, 0.5, 1.3, 3.3, 1.6, 0.8, 
    0.7, 1.3, 0.7, 1.4, 0.7, 3.3, 2, 1, 1.3, 2, 2.1, 2.1, 2, 1.4, 1.8, 2.5, 
    3.2, 1.7, 0.9, 0.8, 0.1, 1, 1, 0.8, 0.3, 0.7, 1, 0.7, 0.7, 0.8, 1.3, 1.3, 
    2.3, 3.3, 2.3, 2.3, 2, 1.8, 2.5, 1.5, 0.8, 0.8, 0.9, 0.5, 0.8, 0.6, 0.2, 
    0.8, 0, 0.7, 0.1, 0.3, 0.6, 0.2, 0.8, 0.8, 1.3, 1.4, 1.2, 1.8, 0.8, 0.9, 
    0.4, 1, 1.3, 1.3, 1.4, 2, 1.4, 1.1, 1.1, 0.8, 0.8, 0.6, 0.6, 1, 0.4, 0.3, 
    0.3, 1, 0, 0.4, 0.8, 0.5, 1, 0.5, 0.9, 1, 1.8, 0.8, 0.4, 1.2, 1, 0.7, 
    0.4, 1, 0.3, 0.6, 0.5, 0.2, 0.6, 0.9, 2.7, 2.3, 2.7, 2, 2, 3.3, 4.2, 1.2, 
    1.3, 2.8, 3.3, 2.4, 0.8, 2.9, 4, 2.5, 3, 1.4, 2.7, 2.4, 1.1, 1.3, 1.4, 
    1.3, 1.5, 1.8, 1.7, 2.1, 2.4, 2.6, 2, 2, 2.3, 1.7, 1.9, 2, 1, 0.8, 1.7, 
    0.1, 0.1, 0.8, 1, 1.2, 1.5, 1.9, 2.7, 1.9, 1.7, 2.5, 2.7, 1.4, 2.2, 2.2, 
    1.6, 2.4, 2.7, 1.1, 1.3, 1.1, 1.4, 2.3, 1.3, 1.5, 2.1, 1, 1.2, 1.1, 0.7, 
    1.3, 1.5, 1.7, 5.6, 2.4, 2, 1.1, 1.7, 3.1, 2.1, 1.1, 1.9, 0.9, 2.3, 1.1, 
    1.8, 1.3, 0.8, 1, 0.4, 1.4, 0.6, 1, 2, 2, 1.1, 1.6, 2.1, 2.3, 2.2, 2.8, 
    2.4, 2.3, 2, 2.3, 2.6, 1.6, 1.9, 1, 1.2, 1.3, 2.5, 2, 4, 4.5, 3.8, 3.4, 
    3.6, 4, 3.3, 3.4, 1.7, 2.1, 3.6, 4.5, 1.3, 0.4, 1.7, 1.2, 2.8, 3.9, 3.3, 
    3.4, 3.8, 2, 2.1, 1.4, 2.5, 1.7, 1.2, 0.5, 0.9, 1.3, 2.6, 4.2, 4.3, 2.6, 
    2.2, 3.8, 4.3, 3, 3.3, 2.6, 2, 1.8, 0.9, 1.3, 1.3, 2.4, 0.8, 4.3, 1.8, 
    1.8, 1.6, 2.1, 2.4, 1, 1.3, 1.5, 1.9, 1.4, 1.8, 1.9, 1.5, 1.3, 3.6, 2.8, 
    1.2, 1.9, 2.4, 2.2, 1.6, 1.6, 1.2, 1.2, 1.5, 0.9, 1.9, 0.5, 1.6, 1.9, 
    2.4, 2.1, 2.8, 3.3, 3.6, 2.4, 2.2, 3.9, 2, 3.3, 1, 2.9, 3.4, 5.2, 3.1, 
    2.9, 3.4, 1.4, 1.5, 3.2, 3, 3.1, 3.5, 3.3, 1.8, 1.3, 2.8, 2.7, 2.8, 4.2, 
    3.9, 3.4, 4.1, 3.4, 2.8, 3.1, 3.2, 4.3, 4, 3.7, 4.4, 3.4, 3.8, 3.8, 4.6, 
    5.1, 4, 2.8, 2.1, 3.7, 3.2, 4.1, 1.7, 3, 4.2, 4.9, 3.7, 3.2, 4, 3.6, 3.2, 
    2.6, 1.5, 2.3, 1.8, 3.3, 1.3, 0.4, 0.5, 1.5, 2.3, 0.9, 2.6, 3, 2.7, 0.9, 
    1.7, 0.7, 1.1, 1.4, 0.9, 1.5, 1.8, 3.2, 2.3, 0.3, 2, 1.4, 4, 4, 4, 3.9, 
    3.4, 3.6, 3.5, 3.6, 3.5, 2.9, 3, 3.8, 3, 2.1, 1.2, 3.3, 2.3, 2.9, 3, 3.5, 
    2.2, 2.2, 2, 1.1, 1.3, 0.9, 1, 0.9, 1.1, 0.8, 1.4, 1.3, 1.6, 1.8, 2.2, 
    2.7, 2.7, 2.9, 3.8, 4.2, 3.4, 3, 3.6, 4, 4, 3.9, 3.5, 3.6, 2.5, 1.6, 1.1, 
    1.1, 1.4, 1.2, 3.3, 2, 3, 1.8, 3.4, 3.9, 2.9, 2, 1.9, 2.9, 2.3, 1.9, 1.9, 
    1.9, 2.9, 2.5, 3, 2.1, 0.7, 1, 1.3, 0.9, 1, 1.1, 1.2, 0.8, 1.2, 1.2, 1.1, 
    1.4, 0.7, 2.6, 1.3, 1.2, 1.4, 3, 3.8, 3.6, 3.9, 4.8, 5, 6.5, 6.9, 5.9, 
    5.7, 5.7, 5.4, 5.1, 3.8, 5.3, 5.1, 4.7, 5.5, 5.7, 6.8, 6.4, 6.2, 5.6, 
    4.9, 5.4, 5.2, 5.9, 5.4, 6.5, 5, 5, 4.4, 4.3, 4.1, 4, 4.4, 4, 4.8, 4, 
    3.1, 1.5, 1.5, 2.3, 2, 2, 1.9, 2.2, 2.2, 1.5, 1.5, 3.4, 3.2, 2.7, 3, 0.5, 
    0, 1, 1, 0.8, 0.4, 0.2, 0.1, 2.5, 0.8, 0.4, 0.8, 4.1, 3.3, 3.3, 4.7, 4, 
    5.8, 5.9, 6.5, 6.7, 4.7, 5.4, 5.5, 5.8, 5.5, 4.2, 3.1, 3.8, 4, 3.5, 3.1, 
    4.3, 4.4, 4.7, 5.7, 5.1, 6.1, 4.1, 5, 4.6, 5, 5.3, 4.4, 2.9, 3, 4.8, 4.8, 
    4.4, 4.1, 2.7, 2.7, 3, 3.1, 3, 2.7, 2.6, 3.3, 2.9, 3.3, 2.9, 2.2, 2.8, 3, 
    3.2, 2.7, 2.9, 2.9, 1.5, 1.9, 1.1, 1.6, 1.1, 1.8, 1.6, 1, 1.4, 1.8, 1.3, 
    0.7, 1, 0.8, 0.4, 1.3, 4, 4.5, 4.6, 3.6, 3.9, 4.8, 4.4, 5, 4.4, 3.3, 4.1, 
    4.1, 4, 3.2, 1.6, 0.5, 1.7, 1.1, 0.7, 1.3, 1.9, 1.2, 0.9, 1.8, 1.9, 2, 
    2.6, 2, 2.2, 2.4, 2.1, 1.9, 1.7, 2.4, 2.1, 1.3, 1.1, 1.3, 1, 1.3, 1.3, 2, 
    0.8, 0.3, 0.8, 1, 1.8, 1.9, 2, 2.4, 2.4, 2.9, 2.8, 2.5, 2.3, 2.4, 2.5, 
    2.1, 2.2, 2.2, 1.9, 2.1, 2.1, 2.3, 2.8, 2.7, 2.2, 3.3, 3.1, 2.5, 2.3, 
    2.7, 2.9, 3.6, 3.7, 4, 4.1, 4.1, 4.3, 3.8, 3.7, 3.4, 3.2, 3, 2.7, 2.2, 
    2.6, 1.8, 1.7, 1.1, 0.7, 1, 1, 0.9, 1.3, 1.8, 2.5, 2.1, 1.6, 1.3, 2.4, 
    2.1, 2.6, 3.2, 3.2, 2.3, 3.4, 2.8, 1.5, 2.6, 1.7, 1.7, 1.2, 2, 1.5, 0.9, 
    1.2, 0.6, 0.8, 0.8, 1.2, 0.2, 0.3, 1, 0.6, 1.5, 1.4, 1.4, 0.9, 0.3, 0.6, 
    0.5, 1.4, 3.9, 4.1, 4.5, 3.9, 2.8, 3.5, 4.1, 4.5, 6.7, 7.5, 6.8, 5.6, 
    6.1, 6, 6.7, 7.5, 6.8, 6.8, 6.7, 8.9, 8.2, 5.5, 5.1, 3.9, 1.5, 2.4, 2.3, 
    2.9, 3, 2.1, 1.7, 3.1, 2.1, 2.4, 2.4, 1.6, 1, 1.8, 1.5, 2.4, 2.2, 2.3, 
    1.2, 1.5, 0.9, 0.3, 1.2, 0.1, 1.2, 0.2, 0.6, 0.6, 0.5, 0.4, 0.4, 1.6, 
    0.7, 2.3, 4.3, 6.2, 8.3, 7.1, 4.8, 4.3, 1.8, 0.4, 1.2, 1.5, 1.6, 2.2, 
    1.8, 2, 1.7, 1, 0.9, 1.3, 0.9, 0.2, 2, 2.7, 5.2, 4.5, 5.1, 2.3, 0.9, 2.5, 
    4, 2.8, 3.4, 1.4, 2.9, 3.7, 3.1, 0.6, 1.2, 2.1, 2, 2.5, 2.6, 0.6, 0.9, 
    0.4, 0.3, 0.7, 0.8, 1.4, 2.2, 1.8, 1.1, 0.9, 1.5, 0.8, 2.2, 0.4, 0.7, 
    0.5, 1, 0.4, 0, 0.3, 0.3, 1.5, 0.2, 0.9, 1, 1.2, 0.8, 1.7, 3.2, 1.1, 0.8, 
    0.9, 2, 2.1, 2.2, 2.3, 1.6, 2, 1.5, 0.7, 1.7, 4.2, 3.2, 4.8, 4.1, 4.6, 
    5.1, 3.7, 2.4, 2.4, 4, 1.7, 3.4, 2.2, 2, 0.8, 0.7, 0.5, 0.2, 1, 1.1, 0.7, 
    0, 0.1, 0.8, 0.7, 0.9, 3.3, 5.2, 5, 4.5, 4.7, 3, 1.6, 2.2, 2, 3.5, 2.1, 
    3.3, 2.9, 2.8, 3.1, 4.4, 4.2, 2, 1.4, 0.8, 1.6, 2.2, 1.7, 1.8, 1.8, 2.1, 
    2.4, 2.6, 1.6, 1.5, 1.3, 1.9, 0.1, 1.4, 2, 2.2, 1.2, 1.7, 1.9, 1.7, 3.2, 
    3.3, 3.2, 3.2, 2.8, 4.9, 7, 7.6, 6.2, 6.9, 7.7, 8.4, 9.2, 5.3, 5, 5.2, 
    5.5, 5, 3.7, 4.1, 4.2, 5.4, 5.5, 2.6, 4.6, 5.4, 3.8, 4.2, 2.3, 2.5, 4.1, 
    3.1, 2, 1.6, 2.6, 1.8, 1.2, 0.8, 1.5, 1.3, 0.8, 1.6, 1.3, 0.7, 2.4, 2.1, 
    2.2, 2.6, 2.7, 3.2, 2, 2, 3, 3.1, 2.8, 3.2, 1.8, 2.1, 2.4, 1.7, 2.1, 0.4, 
    0.3, 1.4, 2.5, 1.7, 1.7, 1.3, 0.7, 1.7, 2, 2.5, 1.2, 0.9, 1.6, 2.1, 2.6, 
    2.7, 2.7, 2.3, 2.9, 3.6, 1.5, 3.2, 2.7, 3.3, 1.6, 2.4, 0.9, 1.7, 1.1, 
    1.5, 1.5, 2.1, 0.7, 1.9, 4, 3.9, 3.5, 5.1, 2.4, 2.3, 2.6, 3.4, 4.1, 3.8, 
    2.9, 2.8, 2.7, 1.8, 0.6, 0.3, 0.3, 3.5, 3.3, 3, 2.7, 2.9, 4.4, 2, 1.8, 
    3.6, 2.9, 1.8, 2.2, 2.7, 2.8, 2, 2.9, 3.7, 4.6, 2.8, 2.4, 3.7, 3.4, 3.2, 
    3.9, 3, 2.5, 1.4, 2.1, 2.8, 2.6, 4.8, 2.1, 6.2, 8, 8, 7.8, 7.3, 8, 8.2, 
    7.1, 4, 1.3, 1.8, 1.4, 2.8, 4.2, 1.6, 1.1, 2.5, 2.7, 5.3, 5.9, 6, 6.4, 
    5.9, 4.6, 3.8, 3.2, 1.7, 1, 1.4, 1.1, 1.1, 2.6, 2, 0.8, 0.8, 1.4, 1.1, 0, 
    0.9, 1.1, 1.9, 1.3, 2, 2.1, 2.3, 2.2, 2.3, 2.3, 2.2, 2.7, 2.7, 2.7, 2.9, 
    2.5, 2.5, 2, 1.2, 0.6, 1.4, 2.2, 1.4, 2, 0.4, 1.9, 2.5, 2.2, 2.9, 2.7, 
    2.5, 2.3, 2.4, 2.8, 3.2, 3.6, 3.5, 3.5, 3.4, 2.7, 3.1, 2.5, 2.6, 1, 0.7, 
    0.4, 2.4, 2, 2.3, 2.4, 2.1, 2.1, 1.4, 2, 2.4, 2.1, 1.5, 2.4, 2.8, 2.3, 
    2.5, 2.1, 2.1, 2.1, 2.1, 2.5, 3.1, 6, 1.2, 1.4, 1.4, 2.2, 2, 1.7, 1.3, 
    1.7, 4.9, 3.5, 3, 1.8, 3.4, 3.5, 3.7, 3.4, 3.1, 4, 4.4, 2.4, 0.7, 1.2, 
    0.8, 0.8, 0.2, 0.1, 0.8, 0.7, 0.4, 1, 2.4, 1.1, 1.2, 1.8, 1.9, 2.4, 3, 4, 
    2.4, 2.9, 2.3, 2.8, 3.6, 3.1, 5.5, 2.3, 3.5, 3.7, 3, 2.8, 1.3, 1.2, 1.6, 
    2.2, 2, 1.6, 1.4, 1.8, 1.8, 2.4, 2.3, 2.1, 2.1, 2.3, 2.7, 2.6, 2.3, 3.5, 
    2.5, 2.3, 2.5, 3.2, 3.4, 4.2, 4.2, 4.3, 4.5, 3, 3, 0.8, 1.6, 1.3, 2.2, 
    1.7, 1.6, 2, 1.3, 1.6, 1.3, 2.4, 2.8, 2.5, 0.7, 1, 0.7, 0.1, 0, 0.2, 0.1, 
    0.2, 0.4, 0.7, 0.5, 0.3, 0.6, 0.6, 1.2, 1.4, 0.9, 0.7, 1.1, 1.1, 0.8, 
    0.7, 1.7, 1.6, 1.8, 1.4, 1.9, 0.6, 1.4, 1.5, 1.4, 0.6, 0.1, 0.9, 2.6, 
    0.7, 2, 1.2, 1.4, 1.3, 2.2, 2.2, 1.7, 2.1, 1.3, 1.4, 2.4, 1, 1.6, 1.5, 
    1.7, 3.9, 3.3, 2.2, 2.7, 3, 2.7, 1.7, 2.3, 2.6, 2.3, 2.7, 2.9, 3.3, 2.6, 
    2.1, 1.9, 1.7, 4.8, 3.4, 1.3, 1.6, 3.5, 3.5, 3.3, 2.4, 2.6, 2.6, 2.8, 
    2.4, 2.3, 3, 2.6, 2, 1.8, 2, 0.8, 2.8, 2.4, 2.5, 2.5, 1.9, 1.5, 1.5, 2.1, 
    1.5, 1.5, 1, 0.5, 1, 0.7, 1.4, 2.2, 0.9, 0.2, 0.9, 0.6, 0.3, 1.6, 1.4, 
    1.7, 1.8, 1.6, 1.8, 1.7, 1.7, 1.5, 0.7, 1.1, 0.4, 0.1, 0, 0.5, 0.3, 0.3, 
    3, 2, 3, 3.6, 4.1, 2.8, 2.1, 3.6, 1.7, 2.7, 3.4, 3.3, 5.3, 3.6, 5.6, 4.6, 
    4.7, 4.5, 4.3, 5.3, 1.9, 0.9, 5.2, 4.5, 5.2, 5.9, 5.3, 4.8, 3.6, 4.9, 
    4.5, 5.1, 4.9, 5.2, 6.2, 6.1, 6.9, 7.8, 6.6, 7.1, 5.5, 5.1, 5.7, 5.1, 
    6.6, 5.3, 5.3, 4.6, 4.6, 6.1, 8.3, 7.4, 8, 8.1, 7.1, 6.8, 8.1, 8.8, 6.1, 
    4.7, 4.1, 4.7, 4.7, 3.8, 4.6, 2.7, 3, 3.1, 1.6, 0.2, 2.4, 1, 0.8, 0.3, 0, 
    0.1, 1.7, 1.5, 0.7, 0.8, 2.1, 1.2, 2.7, 1.6, 4, 2.7, 1.5, 2, 1.6, 1.5, 
    2.6, 4.1, 0.6, 0.3, 0.5, 0.5, 0.5, 1.7, 2.3, 0.8, 0.2, 0.4, 0, 0, 0.1, 1, 
    0.3, 0.9, 0.9, 0.6, 0.9, 1.1, 0.8, 0.1, 1.9, 2.1, 1, 1, 1.4, 0.2, 0.9, 
    2.3, 1.6, 0.1, 0.8, 0.5, 1.1, 0.7, 1.5, 2.8, 1.4, 1, 6.8, 8, 6.1, 7.3, 
    5.8, 4.8, 5.7, 5.1, 3.2, 5.4, 3.6, 3.4, 4.1, 3.1, 4, 2.9, 4.4, 5.7, 4.3, 
    4.5, 6.4, 4.7, 6, 6.5, 6.6, 5.5, 6, 6.2, 6.1, 6.1, 6.1, 6.5, 5.6, 4.6, 
    5.2, 4.3, 3.5, 3.2, 3.1, 2.7, 1.5, 0.5, 1.3, 0.4, 2.5, 2.4, 1.6, 2.1, 
    1.9, 2.5, 2, 2, 2.3, 1.9, 0.9, 1.2, 1.7, 2.9, 3.2, 3.7, 2.1, 3.4, 2.2, 
    0.1, 0.8, 0.5, 0, 0.4, 1.6, 3.7, 4.6, 3.9, 3.9, 3.8, 3.8, 3.8, 2.7, 3.2, 
    3, 2.8, 2.9, 2.1, 2.8, 2.4, 2, 2.1, 2.4, 3, 3.2, 3.2, 1.6, 2.1, 2.1, 2.3, 
    2.9, 3.6, 3.7, 3.1, 3.1, 3.4, 1.1, 1.4, 2.9, 0.5, 0.8, 0.7, 0.7, 0.1, 
    0.6, 0, 0.3, 0.7, 0.1, 0.3, 0.2, 0, 0.9, 2.3, 1.8, 0.8, 2.1, 2.1, 2.2, 
    1.4, 0.9, 1, 1.8, 2.8, 3.4, 3, 3, 3.9, 3.9, 2.4, 2.6, 1.4, 0.5, 2, 1.5, 
    4.2, 4.8, 2, 3.6, 1.7, 0.9, 1.2, 1.3, 2.3, 2.7, 1.3, 0.3, 0.9, 0.7, 0.4, 
    0.4, 0.8, 0.6, 0.4, 0.3, 0.6, 1.1, 0.1, 0.4, 1.7, 0.3, 2.2, 3.1, 4.1, 
    3.4, 3.1, 3.5, 1.8, 1.5, 2, 1.3, 2.9, 3.4, 2.9, 2.1, 2.9, 2.3, 1.7, 1.4, 
    0.5, 0.9, 0.2, 1.4, 1.6, 2, 2.1, 3.1, 2.5, 2.2, 1.5, 1, 2.1, 2.3, 1.6, 
    2.4, 1.4, 0.1, 0.8, 1.2, 2.3, 3.8, 1.2, 1.2, 0.3, 1.9, 0.5, 0.3, 0.7, 
    2.1, 2.8, 1.1, 1.4, 1, 0.3, 1, 4.2, 3.4, 3.3, 3.6, 6.5, 5.8, 4.6, 4.4, 4, 
    3.8, 4.1, 4.4, 3.3, 3.5, 2.8, 4, 4.3, 3.3, 4.4, 3.6, 4.8, 5.5, 6.5, 7.2, 
    6.2, 6, 6.1, 5.1, 4.6, 4.4, 4.2, 1.9, 2.5, 1.8, 2, 1.6, 1.2, 0.7, 0.7, 
    0.7, 0.8, 0.6, 1.3, 1.5, 0.8, 1.4, 1.3, 3.4, 2.5, 3.2, 2.6, 1.1, 0.5, 
    1.2, 0, 0.6, 1.3, 0.5, 0.6, 0.6, 0.6, 0.2, 0.1, 0.2, 0.1, 0, 0.8, 0.2, 
    1.2, 1.1, 2.8, 2, 1.4, 0.2, 0.3, 1.2, 0.4, 0.7, 0.6, 0.5, 0.5, 0.3, 0.2, 
    0.6, 0.7, 0.3, 0.8, 0.1, 2, 1.2, 2.1, 2.1, 1.4, 1.3, 1.2, 1.7, 0.3, 0.9, 
    0.6, 1.4, 1.4, 2.8, 2.8, 1.4, 0.6, 0.6, 1.5, 0.8, 0.7, 1.1, 1, 1.2, 1.9, 
    1.1, 1.1, 2.4, 2.7, 3.8, 2.6, 2.7, 4.4, 2.4, 3.9, 5.7, 6.1, 2.9, 3, 3, 
    4.4, 1.5, 2.9, 3, 2.1, 2.4, 0.8, 1.5, 1, 1.5, 1.1, 2.8, 6.4, 5.7, 4.7, 
    4.5, 4.3, 2.9, 1.3, 1.5, 0.9, 0.8, 0.4, 0.4, 0.4, 0.2, 0.4, 0.4, 0.7, 
    0.7, 0.5, 1.3, 0.7, 0.6, 0.7, 0.8, 0.9, 0.5, 0.1, 0.3, 0, 0, 0.9, 0.9, 
    0.8, 0.8, 1, 0.9, 0.7, 2.2, 0.7, 0.2, 0, 0.5, 1, 0.5, 0.2, 1.8, 0.2, 0, 
    1.1, 0.6, 0.8, 1.1, 1.5, 0.6, 0.7, 1.2, 1, 0.2, 0.8, 0.5, 2.7, 1.2, 3.6, 
    4.4, 4, 1.9, 1.3, 1.2, 1.6, 1.4, 1.8, 3.2, 2.9, 1, 1, 1, 2.1, 3.5, 3.5, 
    8.1, 6.3, 4.4, 3, 5, 7.4, 5.4, 5.6, 3.8, 3.4, 4.6, 4, 4, 4, 4, 3.9, 5.5, 
    5.4, 4.9, 4.8, 5.3, 2.7, 2, 1.9, 1.8, 1.8, 2.2, 0.7, 0.6, 0.2, 1, 0.4, 
    0.4, 0.5, 0.6, 0.9, 0, 0.1, 0.1, 1, 0.5, 0, 0, 0.2, 1.3, 0.2, 1.1, 0.4, 
    0.6, 1.5, 0.3, 0.2, 0, 0.1, 0.8, 0.7, 0.3, 0.6, 0.1, 0.5, 0.4, 0.5, 2, 
    1.9, 0.4, 0.9, 0.9, 1, 1.4, 4.1, 4.1, 4.3, 5.7, 5.7, 5.2, 4.5, 3.9, 3.9, 
    2.1, 1, 2.3, 1.5, 4.6, 1, 2.5, 3.6, 3.8, 3.3, 3.4, 2.9, 3.8, 6.5, 6.1, 
    2.9, 1.2, 0.7, 1.5, 1.4, 0.7, 0.2, 0.8, 0.8, 0.3, 0.1, 0.1, 1, 0, 0.8, 
    0.1, 0, 0.1, 0.6, 0.5, 0.5, 0.2, 0.2, 0.1, 0, 0.5, 1, 0.1, 0, 0.1, 0.2, 
    0.5, 0, 0.1, 1.2, 0.8, 1.5, 0.8, 0.6, 1, 0.2, 0.9, 0.1, 0.8, 1.2, 0.5, 
    2.5, 2, 1.5, 1, 1, 0.7, 0.6, 1.4, 0.7, 0.3, 0.5, 1.3, 0.5, 0.2, 1.1, 0.9, 
    0.1, 0, 1.3, 0.3, 0.9, 1, 1, 1.9, 4.9, 2.7, 3.4, 3.3, 5.8, 4.6, 5.1, 5.3, 
    3.1, 2.7, 4.4, 4.9, 4.9, 5.7, 4.5, 5.4, 5.8, 4.4, 4.4, 5.7, 5.5, 6.2, 
    5.9, 6, 7.2, 7.4, 7, 6.8, 7, 5.8, 7.9, 6.4, 8.5, 7.7, 7, 8.6, 8.4, 9.2, 
    8.6, 8.8, 8.7, 8.5, 9, 9.6, 8.7, 9.6, 9.5, 9.1, 8.7, 8, 7.2, 7.5, 6.9, 
    6.2, 8.5, 7.9, 9.9, 8.6, 7.8, 8.1, 8.8, 6.9, 8, 6.3, 6.4, 8.2, 7.8, 6.9, 
    8.8, 7.9, 7, 5.2, 7.2, 9.1, 8.8, 6.8, 4.2, 3.7, 2.7, 2.7, 5, 5.1, 4.8, 5, 
    4.4, 4.6, 4.5, 5.3, 3.4, 3.6, 4.5, 4.3, 3.4, 3.5, 2.9, 1.8, 1.8, 0.6, 
    1.2, 0.4, 0.6, 0.6, 1.8, 1.1, 1.5, 0.1, 0.4, 0.5, 1.1, 1, 0.4, 0.5, 0.5, 
    0.7, 0.8, 0.3, 1.5, 2.5, 2.2, 1.9, 1.7, 1.1, 0.3, 1.6, 3.7, 2.7, 1.9, 
    0.3, 0.8, 0.7, 0.7, 0.2, 0.2, 0.5, 0.7, 0.9, 1.9, 2.1, 1.9, 1.4, 1.3, 
    1.1, 0.7, 1, 0.9, 0.4, 0.3, 1.4, 0.8, 0.6, 0.8, 0.8, 0, 0.1, 0.3, 0, 0.8, 
    0.3, 0.7, 1.3, 0.6, 0, 0, 1, 0.6, 0.2, 0.3, 0.2, 0.2, 0.1, 1.5, 0.1, 0.1, 
    0.2, 0.8, 0.9, 0.3, 0, 0.2, 0, 1, 1.2, 0.9, 1.1, 1, 0.9, 0.3, 0.5, 0.8, 
    4.1, 3.4, 0.8, 3.7, 3.9, 2.4, 4.9, 6.8, 7.5, 7.2, 8, 7.5, 5.1, 5.9, 5.3, 
    4.2, 5, 6.5, 5.4, 5.4, 4.7, 5.2, 4.1, 0.6, 0.9, 1.8, 0.5, 2.2, 3.8, 5, 5, 
    4.9, 2.8, 0.7, 1, 1.7, 4.1, 2.4, 3.8, 5.3, 1.8, 0.8, 1.5, 0.5, 0.3, 1.1, 
    0.3, 0.3, 2, 0.1, 0.2, 0.2, 1.3, 0.5, 0.4, 0.2, 0, 0.1, 0, 0, 0, 0.7, 
    1.2, 0.2, 0, 0, 0.6, 0.7, 0.1, 0.1, 0.8, 0.4, 0.6, 1.1, 0, 1.1, 0.6, 0.3, 
    0.2, 0, 0, 0.1, 0, 0, 0, 0.5, 0.5, 1, 0, 0, 0.1, 0.6, 1.2, 1.9, 1.2, 0.6, 
    0.3, 1.1, 0.1, 0.3, 0.6, 0.2, 0.5, 0, 0.2, 0.1, 0, 0.5, 0.7, 0.7, 1, 0.3, 
    0.8, 0.8, 0.6, 1.4, 2.2, 3.4, 1.8, 0, 1.2, 6.4, 8, 7.3, 11.5, 11.5, 9.1, 
    8.1, 7.6, 6.3, 4.2, 3.7, 3.5, 4, 2.7, 4, 2.9, 2.7, 0.5, 0.4, 1.4, 0.9, 
    0.6, 0.1, 0.6, 0.6, 1.4, 1.6, 1, 0.3, 0.3, 0.1, 0.5, 1.1, 1.2, 1.3, 0.7, 
    0.8, 1.1, 0.2, 1.2, 1.5, 3.3, 1.5, 0.3, 1.3, 0, 0.8, 0.9, 1.2, 0.8, 3, 
    3.5, 1, 0.9, 0.2, 0.2, 4.4, 5.3, 5.9, 8.4, 8.2, 7.7, 5.2, 5.9, 6.5, 5.8, 
    5.5, 5, 5.7, 6.9, 5.7, 5.1, 3.9, 4.7, 3.4, 4.9, 4.9, 5.4, 5.8, 2.6, 2.2, 
    3.3, 5.4, 3.7, 4.7, 3.7, 4.7, 3.8, 5.2, 4.8, 4, 3.2, 4, 4.6, 4.5, 0.7, 
    0.2, 0.3, 3.3, 2.5, 2.1, 1, 1.3, 0.2, 0.9, 1.1, 0.4, 2.1, 2.6, 3.4, 3.9, 
    5.8, 5.8, 5.7, 4.6, 3.5, 1.8, 4, 1.7, 3.7, 4.4, 3.2, 2.1, 2.1, 4.2, 4.2, 
    5.5, 4.5, 2.2, 0.7, 0.4, 3.7, 3.1, 2.9, 1.3, 2.2, 4.1, 1.6, 2.3, 1, 0.5, 
    1.2, 0, 0.8, 0.6, 1, 0.7, 0.7, 0.1, 0.1, 0.8, 1.5, 0.1, 0.4, 0.3, 0.5, 
    0.3, 0.6, 0.6, 0.1, 0.7, 0.5, 0.8, 0.8, 0, 0, 0.3, 0.4, 0.4, 1.3, 0.7, 1, 
    1.8, 1.4, 1, 0, 0.3, 1.1, 0.3, 0.3, 1.1, 0.5, 1.4, 1.4, 1.8, 0.1, 0.4, 
    0.9, 0.3, 0.3, 0.6, 0.1, 0.4, 0.1, 0.9, 1, 0.3, 0.9, 1.2, 0.1, 0.6, 0.3, 
    1.4, 1.3, 0.9, 0.8, 0.1, 0, 0.3, 0, 0.4, 0.1, 0, 0.3, 0, 0.3, 0.1, 0.3, 
    1, 0.3, 0.2, 0.2, 1.2, 0, 0.4, 0.1, 0.8, 0.6, 0.8, 0.5, 0.8, 0.8, 2, 1, 
    1.4, 0.9, 0.8, 2.6, 0.7, 2.2, 1, 1.3, 0.2, 1, 1, 1, 0.1, 0.7, 0.1, 1.8, 
    0.2, 0.5, 0.1, 0.7, 1.1, 0.5, 0.6, 0.7, 0.4, 1, 0.8, 1.7, 0.4, 1.2, 3.2, 
    1.5, 1, 0.6, 0.7, 2.1, 3.6, 2.7, 2.3, 3.6, 2.7, 2.3, 2.5, 2.1, 1, 0.3, 
    0.2, 0.7, 1.3, 1.6, 3.3, 2.7, 3.4, 3.2, 3.2, 3.6, 4.7, 6.4, 5, 6.4, 4.4, 
    5.3, 5.2, 5.5, 5.2, 3.7, 3, 3, 1.6, 1.8, 0.4, 0.5, 1, 0.7, 1.3, 0.8, 2, 
    2.1, 2.8, 1.1, 2.5, 2.8, 2.8, 2.4, 1.8, 2.4, 0.3, 0.9, 1.8, 0.9, 0.7, 
    0.9, 1.2, 0.6, 0.8, 0.5, 1, 1.3, 1.3, 1.2, 0.5, 1.5, 2, 1.2, 0.6, 0.4, 
    1.2, 1.1, 0.8, 0.1, 0.5, 0.2, 0.7, 0.1, 0.7, 0.8, 1, 1.2, 0.7, 0.4, 0, 
    0.3, 1, 1.3, 0.7, 0.6, 0.7, 0.2, 0, 0, 0, 0.8, 0.5, 0.3, 0.4, 0.5, 0.6, 
    0, 1, 1.5, 0.6, 0, 0, 0, 0, 0, 0, 1.4, 0.6, 0.8, 1.3, 1.6, 4, 2.2, 2.4, 
    0.6, 1.2, 0.7, 0.3, 0.1, 0.2, 0.9, 1, 0.7, 1.1, 0.2, 2.2, 0.3, 0.6, 0.7, 
    1.6, 2.6, 1, 0.4, 1.5, 1.1, 0.6, 0, 0.5, 0, 0.7, 0, 0.9, 0, 0.1, 0.6, 
    0.1, 2.5, 0.4, 0.3, 0.3, 0.8, 0.4, 0.1, 0.2, 0.7, 2, 1.4, 1.4, 0.7, 1.4, 
    0.6, 0, 0, 0.1, 0, 0.4, 0.4, 0.4, 1, 0.6, 1, 1.3, 0.2, 1.2, 1.6, 1.6, 
    0.8, 0.9, 1.6, 1.4, 1, 1.5, 4.3, 1.6, 1.1, 2.3, 1.2, 2, 1, 0.8, 1.5, 1.6, 
    1.5, 3.5, 3.9, 1.3, 0.5, 0.3, 3.5, 4.8, 5, 5.1, 5.2, 3.6, 5.4, 4.7, 4.8, 
    4.6, 4.4, 4.9, 3.8, 3.9, 4.5, 4.2, 0.5, 3.9, 2.9, 3.6, 4.3, 5.7, 5.4, 
    5.2, 4.9, 1.8, 5.1, 5, 5.8, 7.6, 7.3, 8.1, 7, 7.3, 7.6, 8.3, 6.5, 7.4, 
    7.9, 7.6, 7.2, 6.9, 6.5, 6.5, 6.9, 4.9, 6.7, 6.9, 7.2, 6.6, 5.8, 5.7, 
    5.4, 6.3, 6, 6.6, 8.2, 6, 4.8, 5.5, 6.4, 4.8, 4.8, 4.8, 4.3, 4.2, 3.8, 
    5.9, 5.9, 5.2, 5, 6.1, 5.2, 4.3, 6.7, 6.9, 4.6, 6.4, 5.2, 5.1, 5.6, 6.8, 
    5.4, 5, 5.3, 4.7, 4.1, 5.1, 4.7, 4.5, 4, 3, 3.4, 2.9, 5.1, 4.2, 4.3, 2.8, 
    3.4, 1.9, 1.8, 1.1, 1.3, 0.6, 1.6, 0.9, 1, 1, 1.5, 1.9, 2.2, 1.3, 0.1, 
    0.3, 1.4, 2.5, 2.7, 1.7, 3.7, 3.1, 2.4, 2.9, 4.2, 3.6, 3.1, 3.1, 3.4, 
    2.9, 1.6, 1.8, 1.2, 0.8, 1.3, 1.6, 1.7, 1, 1, 1.7, 1.6, 1.4, 0.2, 0.9, 
    1.2, 0.7, 0.3, 1, 0.8, 0.6, 0.5, 1.2, 0.1, 0.3, 0.7, 0.7, 0.4, 0.7, 0.8, 
    0.1, 0.4, 0.9, 0.7, 0.6, 1, 0.4, 1.4, 1.6, 1.2, 0.3, 0.2, 0, 0.2, 1.4, 
    0.5, 0.4, 0.1, 0.2, 0.6, 0.6, 0.5, 0.5, 0.4, 0.2, 0.6, 1.3, 0.9, 0.9, 
    1.1, 0.8, 0, 0, 1, 1.8, 0.8, 1.1, 0.1, 0.8, 0.7, 1, 1, 0.2, 0.4, 0.2, 
    0.6, 0.8, 0, 0.6, 0.5, 0.5, 0.1, 0.4, 0.4, 0.2, 0.6, 0.7, 1.4, 0.9, 1.1, 
    1.1, 1.6, 2.4, 0.5, 0.3, 0.6, 0.5, 0.3, 0.5, 0.1, 1.4, 0.9, 0.2, 2.2, 4, 
    4.6, 3.1, 2.2, 1.4, 1.4, 5.4, 4.9, 6.3, 5.2, 6, 5, 4, 5.1, 3.8, 6.2, 4.9, 
    3.8, 4.2, 2.2, 1.1, 0.2, 1.9, 1.5, 2.2, 1.3, 1.4, 1.3, 0.8, 1.7, 2, 1.7, 
    2.4, 2.4, 1.3, 1.5, 1.1, 1.2, 1, 0.9, 0.1, 0.2, 0.6, 0.8, 1.1, 0.9, 4.9, 
    5, 6.3, 6.1, 5.1, 6.3, 5.8, 5.7, 5.7, 5.5, 4.1, 6.4, 1, 0.8, 0.5, 0.4, 1, 
    1, 0.2, 0.9, 1, 1.2, 2.3, 1.8, 1.4, 1.2, 1, 1.4, 1.4, 0.2, 0.7, 0.4, 2, 
    1.3, 1.2, 0.1, 1.3, 1.2, 2.1, 0.3, 1.3, 0.6, 0.1, 2.7, 2, 0.3, 1.2, 1.2, 
    1.3, 0.6, 3.6, 5.4, 6.8, 6.2, 6.1, 6.3, 5, 5.8, 5.9, 8.2, 8.3, 7.6, 5, 
    3.2, 4.1, 4.4, 3.5, 4.3, 3.3, 2.6, 4.3, 3.9, 2, 3.6, 4.4, 2.6, 1.9, 1.5, 
    3.7, 3.2, 2.3, 2.4, 1.8, 1.6, 3, 3, 2.1, 0.1, 1.9, 3.3, 2.4, 3.5, 3.6, 6, 
    6.1, 4.2, 4.7, 4, 4.5, 3.3, 4, 5.6, 7.2, 7.5, 7.5, 11.7, 5.2, 5.5, 4.4, 
    3.6, 3.2, 3.1, 3.3, 2.6, 2.6, 4.8, 4.5, 3.8, 12.9, 13.1, 13.5, 12.7, 
    11.3, 11.5, 5.5, 6.1, 7.7, 6.1, 6.9, 7.3, 6.7, 5.7, 8.6, 8, 8.7, 4.5, 
    5.6, 5.9, 9, 4.2, 2.9, 1.4, 2.1, 2.7, 2.8, 1.9, 3.1, 1.8, 2.1, 2.6, 1.8, 
    2, 2.8, 2.5, 2.9, 1.8, 1.6, 2.7, 3.1, 1.8, 0.7, 0.8, 1.2, 0.9, 0.9, 1, 1, 
    1, 0.9, 0.2, 0.4, 0.9, 0.1, 0.2, 0.6, 0.7, 0.1, 0.9, 0.8, 0.7, 0, 1.5, 1, 
    0.8, 0.1, 0.3, 0.9, 0.8, 0.5, 1.3, 1.5, 1, 1.4, 0.3, 1, 0.8, 0, 0.4, 0.9, 
    0.5, 3.3, 4.3, 4.5, 4.9, 4.2, 4.7, 6, 5.8, 5.2, 4.2, 3, 1.2, 5.9, 5.3, 
    0.9, 1.3, 2.1, 3.3, 1.3, 4.3, 4, 4.1, 2.6, 5, 2.8, 2.6, 1.9, 4.8, 2.8, 
    3.8, 5.6, 5, 4.8, 2.2, 2.5, 3, 1.3, 2.3, 2.5, 5.7, 5.9, 3.9, 3.5, 3.3, 
    2.1, 2.6, 6.7, 7.4, 3.8, 4.1, 4.6, 3.6, 2.5, 4.6, 9.4, 8.4, 7, 7.6, 7.8, 
    8.5, 7.1, 6.6, 8, 8.6, 6.2, 6.1, 7.1, 6.4, 2.9, 3, 2.2, 1, 1.4, 2.4, 2.6, 
    2.1, 3.2, 6.9, 4.6, 6.4, 6.1, 5.9, 6.3, 2.8, 1.7, 3, 5.1, 1.6, 0.4, 1.3, 
    0.8, 0.1, 0.7, 0.6, 0.9, 0, 1.3, 2.4, 0.9, 0.4, 0.5, 0.5, 0.2, 0.7, 0.6, 
    1.2, 2.5, 1.6, 1.3, 0.6, 2.2, 1.2, 3.1, 1.3, 1.2, 1, 1.6, 0.2, 0.1, 1.1, 
    0.7, 1.4, 0.1, 0.8, 0.1, 1, 0.6, 1.4, 0.9, 1, 2.7, 2.1, 2.3, 0.4, 0.5, 
    1.2, 1.2, 0.9, 1, 3.7, 3.7, 6, 6.8, 6.8, 4.3, 6.2, 6.2, 6.4, 8, 7.5, 9.8, 
    9.8, 9.8, 8.2, 8.8, 8.4, 7.8, 7.7, 8.1, 6.6, 8.3, 9.5, 10.4, 9.7, 9.7, 
    9.4, 10.7, 11.8, 12.4, 10.3, 11, 10.5, 10.4, 11, 10.4, 8.8, 9.9, 9.6, 
    9.5, 8.9, 10.9, 11, 11.2, 9.8, 9, 9.3, 10.8, 11.1, 8, 7.1, 7.6, 4.9, 6.5, 
    9.8, 9.3, 8, 8.2, 8, 7.5, 6.6, 6.5, 7, 7.9, 8.5, 7.8, 8.7, 9.8, 9.2, 9.5, 
    9.6, 11, 10.4, 9.4, 9.4, 6.8, 10, 10.1, 7.3, 7.5, 8.8, 6.5, 8.4, 8.5, 
    10.2, 9, 7.5, 7.1, 8.6, 8, 8.4, 8.2, 8.3, 6.5, 6.4, 6.4, 6.2, 4.9, 5.9, 
    6.4, 6.3, 4.1, 5.2, 6.5, 4.5, 3.1, 2.4, 5.3, 5.7, 3, 5.7, 2.2, 3, 3, 1, 
    0.7, 1.3, 1.3, 1.8, 0.2, 0.8, 0.8, 0.6, 0.4, 0.9, 0, 0.5, 0.1, 1.5, 1, 
    0.7, 1, 1.1, 0.4, 0.4, 0.1, 0.6, 1.3, 0.5, 0.3, 1.1, 0.5, 0.7, 0, 0, 0.2, 
    0.6, 0.8, 0.8, 0.9, 0.6, 0.6, 0.5, 0.4, 0.4, 0, 0.8, 0.8, 0.8, 0.4, 1.4, 
    0.1, 0, 0.5, 0.8, 0.2, 0.4, 0.6, 0.5, 0.4, 1.3, 3.6, 4.4, 2, 2.9, 6.3, 
    4.9, 4.1, 2.6, 4, 4.3, 4.5, 5, 6.2, 4.6, 6.2, 5, 4.3, 3.3, 3.9, 7.1, 8.3, 
    5.3, 5.1, 4, 5.8, 3.8, 5, 6, 6, 4.5, 5, 2.2, 5.9, 5.7, 6.8, 2.5, 3.1, 
    4.9, 4.3, 5.2, 5.2, 5.3, 6.3, 5, 5.2, 6.6, 6, 6.6, 5.7, 7.1, 6.6, 7.5, 
    6.5, 5.3, 7.1, 5.9, 4.7, 4.6, 4.1, 3.2, 5.5, 5, 1.8, 4.7, 4.5, 3.7, 4.3, 
    4.3, 4.3, 3.6, 4.4, 5.3, 5, 5.4, 6.4, 5.6, 4.9, 7.7, 6.6, 8.1, 8.3, 8.1, 
    8.1, 9.4, 7.5, 6.4, 6.5, 6, 4.7, 5, 3.7, 4.7, 5.6, 4.2, 4.6, 3.5, 6.3, 
    5.7, 4.2, 2.2, 4.2, 1.9, 2.3, 4.7, 5, 3.7, 5.1, 5.1, 5.1, 4.1, 4.8, 3.2, 
    4.1, 3.8, 4.1, 4.6, 4.6, 3.7, 4.3, 4.3, 4.7, 3.8, 4.4, 3.8, 3.8, 7.8, 
    8.3, 7.8, 5.6, 4.9, 5, 6.4, 7, 7.3, 6.2, 6, 5.7, 5.6, 6.8, 6.3, 5.4, 4.6, 
    4.2, 3.4, 3.3, 3.9, 3.5, 3.5, 3, 6.5, 5.8, 5.6, 5.6, 5.6, 5.6, 3.6, 3.9, 
    3.6, 4.5, 4.5, 3.9, 4.8, 4, 4.4, 4.3, 3.1, 4.3, 3.9, 4.3, 6, 4.5, 4, 6.9, 
    5.8, 5.8, 7.2, 5.8, 6.3, 6.7, 6.1, 6.8, 6.2, 5.9, 6, 7.8, 6.9, 5.9, 5.3, 
    3.3, 3.7, 5.3, 4.5, 6.9, 7.2, 6.3, 4.8, 4.3, 3.2, 5.6, 6.2, 6, 5.1, 5.7, 
    7.3, 7, 7.2, 8.6, 5.1, 5.9, 6, 5, 7, 6.7, 6.1, 7, 6, 5.9, 8.8, 4.3, 3.8, 
    3.9, 2.9, 2.7, 2.7, 2.7, 2.7, 4.5, 6.3, 4.3, 4.3, 5.8, 4.7, 5, 5.7, 4, 
    1.7, 1.5, 2.2, 1, 1.6, 1, 1.5, 1.3, 2.3, 1.7, 0.5, 0.7, 1.4, 0.8, 0.5, 
    1.2, 1.2, 1.7, 1.1, 2.2, 0.5, 0.3, 0.4, 0.7, 1.2, 0.4, 0.5, 0.8, 0.3, 
    0.9, 0.7, 1.5, 0.9, 1.3, 1.2, 0.5, 0.4, 0.7, 0.5, 1.2, 1.2, 0.3, 0.8, 1, 
    0.6, 1.1, 0.2, 1, 1.1, 1.5, 0.8, 1.1, 0.8, 1, 1.1, 0.2, 0.3, 1.5, 2.8, 
    4.9, 5, 6.2, 6.5, 7.6, 7.1, 6.2, 5.4, 6.4, 3.7, 2.8, 3.4, 3.4, 3.4, 1.2, 
    1.3, 2.1, 1.5, 3.3, 3.3, 3.9, 6, 1.9, 1, 0.8, 1.8, 1.7, 2.6, 1.2, 1.6, 
    1.2, 1.2, 0.8, 2, 1.6, 2.5, 3.4, 3.4, 4.8, 2, 2.4, 0.5, 0.4, 0.5, 2.1, 
    2.3, 1.6, 1.5, 0.9, 0.9, 0.6, 0.7, 0.6, 0.4, 1.5, 1, 0.9, 1.2, 1.4, 0.5, 
    1.1, 0.3, 1.3, 0.8, 1.2, 0.9, 0.2, 1.4, 0.8, 1.4, 1.1, 0.5, 1, 1, 1.2, 1, 
    0.6, 2.6, 4.3, 6, 2.6, 5, 5.4, 2.9, 4.8, 8.7, 9.9, 9.6, 8.3, 8.3, 6.7, 5, 
    4.3, 5, 5.1, 4.5, 3.8, 3.2, 1, 0.5, 1.2, 0.1, 0.5, 1.1, 1.1, 0.7, 0.8, 1, 
    1.5, 1.5, 0.6, 0.2, 1.1, 1.3, 0.8, 1.6, 4.4, 4.4, 6.7, 6.7, 5.9, 5.5, 
    7.3, 8.9, 8.2, 9.1, 6.9, 8.5, 8.7, 4.3, 8.3, 4.1, 8.5, 5.4, 7.3, 5.8, 
    1.8, 2.7, 1.7, 0.7, 4.1, 3.7, 4, 1.3, 1.6, 2.1, 2.3, 5.1, 6.5, 8.5, 7.1, 
    8, 7.3, 7.5, 7.6, 7.4, 8, 7.7, 8.7, 8.2, 7.1, 6.3, 8.7, 7.2, 4.6, 4.1, 
    5.4, 8, 5.5, 5.6, 6.2, 5.9, 4.3, 4.6, 4.8, 6.4, 5, 6.7, 3.7, 3.9, 3.7, 
    2.5, 2.8, 3.6, 2.4, 3.9, 2.4, 2, 0.9, 0.6, 0.7, 1.8, 1.7, 0.4, 0.4, 0.7, 
    2.1, 1.2, 1.6, 1.6, 2.3, 1.7, 2.8, 0.8, 1, 2.6, 2.6, 2.9, 1.4, 0.8, 1.8, 
    1.7, 1.4, 3.1, 2, 4.9, 5.9, 5, 3.4, 3.5, 3.7, 3.9, 4.5, 4.2, 5.4, 5.9, 
    5.8, 6.8, 3.4, 6.9, 6, 3.6, 3.6, 4.4, 7.6, 8.8, 7.4, 5.2, 5.1, 6.4, 5.6, 
    6.9, 6.7, 5.1, 4.4, 5.9, 5.1, 5.4, 7.4, 6.6, 4.9, 5.3, 5.3, 7.6, 7.5, 
    8.5, 9.1, 8.5, 7.7, 6.6, 5.8, 8.6, 10.6, 9.9, 8.9, 6, 5.4, 10.3, 6.4, 
    7.5, 4.4, 5.5, 5.5, 5.9, 6.7, 8, 7.7, 6.6, 7, 8.9, 6.6, 4.3, 2.7, 4.6, 
    5.5, 4.2, 5.4, 5.1, 6.2, 6.8, 7.7, 6.2, 6.3, 5.7, 5, 4.5, 5.5, 4.7, 3.7, 
    2.9, 1, 1.7, 1.2, 1, 1.1, 1.1, 0.6, 1.6, 0.9, 0.2, 1.8, 1.9, 1.2, 0.8, 
    0.9, 0.3, 1.1, 0, 1.6, 0.8, 3.3, 3.3, 3.5, 4, 3.4, 4.6, 6.1, 5, 5.9, 5.8, 
    6.6, 6.6, 8.1, 7.4, 6.7, 5, 2.4, 2.3, 4.3, 4, 6.4, 3.6, 3.3, 3.9, 3.3, 
    2.9, 3.1, 3.6, 2.1, 1, 1.5, 2.4, 4.3, 5.2, 6.6, 7.8, 7.3, 4.2, 5.6, 5.5, 
    5.9, 4.7, 4.7, 5.6, 5.3, 4.9, 6.2, 4.4, 5.5, 5.2, 5.3, 8, 4.8, 3.8, 5.9, 
    4, 2.3, 3.4, 4, 3.4, 1.2, 0.9, 1.2, 0.9, 0.5, 1.3, 1.1, 1.1, 1.9, 0.6, 
    0.9, 1.1, 2.6, 1.6, 1.5, 1, 1.4, 1, 4.2, 4.8, 4.1, 4.1, 2.5, 5.2, 5.2, 
    4.7, 4, 5, 5.6, 3.6, 3.4, 4.8, 5.6, 3.6, 3.5, 3.5, 1.4, 2.8, 3.1, 3.6, 
    4.5, 2, 3.2, 5.5, 1.4, 4, 1.6, 0.7, 1.5, 2.9, 3.2, 2.5, 3.3, 2, 2.1, 1.2, 
    1.1, 2.7, 0.9, 1.8, 1.9, 2, 1.4, 2.2, 2.5, 2.2, 2, 1, 1.4, 1.2, 1.2, 0.1, 
    1, 1.5, 0.4, 2.2, 0.6, 0.3, 0.6, 0.9, 2.5, 2.6, 1.8, 1.5, 1.1, 0.8, 2, 
    1.9, 1.1, 1.6, 2.3, 2.6, 3.1, 0.6, 2.3, 2.1, 1.9, 1.7, 1.7, 1.5, 1.5, 
    1.4, 2.5, 0.8, 1.2, 0.9, 0.9, 0.3, 1.8, 2, 2, 1.5, 0.7, 0.8, 0.3, 0.5, 
    0.6, 0.8, 1.3, 0.8, 1, 1.2, 1.6, 3.2, 2.1, 1.6, 0.9, 1, 0.4, 0.7, 0.3, 
    0.6, 0.9, 0.7, 0.9, 0.5, 0.6, 0.9, 1.8, 1.8, 2.6, 0.7, 0.3, 1.1, 0.7, 
    1.5, 1, 1, 1.2, 1.1, 0.7, 1, 5.1, 2.9, 4.7, 5.7, 8.7, 10.7, 12.3, 11.6, 
    12.2, 12.1, 11.2, 9.8, 9.8, 9.8, 7.2, 5.7, 2.5, 1.4, 0.8, 1, 1.7, 2.6, 
    3.4, 1.2, 2.1, 0.7, 0.9, 0.5, 0.7, 0.2, _, _, _, _, _, _, _, _, _, _, 
    2.6, _, _, _, _, _, 3.8, 3.8, 1.5, 1.4, 0.5, 0.8, 0.5, 1.1, 4.9, 1.2, 1, 
    2.3, 1.6, 1.6, 2, 2.1, 1, 1.1, 1.9, 3.2, 2.5, 2.7, 3.9, 5.6, 3.9, 2.1, 4, 
    3.5, 4.8, 4.5, 3.7, 2.9, 0.7, 0.8, 1, 1.3, 1.9, 0.6, 5.8, 5.8, 5.7, 4.8, 
    1.1, 1.7, 2.2, 2.5, 4.5, 5, 5, 4.8, 4.1, 6.4, 5, 5.9, 2.9, 4, 4.8, 5.8, 
    5.5, 5.7, 5.3, 3.5, 7.7, 7, 6.9, 5.1, 5.1, 5.9, 4.1, 1.6, 1.3, 0.8, 1.3, 
    2, 1, 2.9, 3.3, 2.7, 1.3, 1.7, 2.4, 0.9, 2.2, 1.6, 1.5, 1.8, 3, 2.5, 3.8, 
    2.6, 3.7, 4.1, 1.7, 2.8, 2.6, 5, 5.8, 7, 4.9, 4.6, 4.5, 4.3, 3.6, 3.9, 
    2.2, 2, 1.1, 1.8, 1.9, 0.8, 4.7, 1.2, 4.2, 2.6, 0.9, 2.9, 3.1, 3.1, 4.6, 
    4, 2.6, 6.1, 5.4, 5.5, 3.4, 2, 1.1, 4.1, 2.4, 2.3, 4.5, 1.6, 1.2, 1.8, 
    3.2, 2.2, 1.9, 5, 3, 2.9, 4, 4.6, 5.4, 7.1, 10.2, 11.9, 8.1, 5.5, 3.5, 
    2.6, 2.8, 2.2, 1.5, 2.9, 3.7, 2.2, 3.9, 2.5, 0.4, 3.1, 1.9, 0.6, 0.5, 8, 
    5.8, 10.8, 2.9, 1.7, 3, 4.6, 1.2, 4.5, 5.9, 3.1, 4, 3.2, 3.2, 2.8, 1.3, 
    1.9, 3.6, 1.8, 0.8, 3.2, 2.7, 2.7, 1.9, 2.5, 3.9, 4, 4.2, 4.1, 3.8, 4.5, 
    3.3, 4.7, 4.6, 4, 5.6, 4.9, 3.7, 6, 6, 4.5, 4.6, 5.5, 4.9, 1.4, 4.7, 3.9, 
    1.5, 1.6, 1.3, 3.1, 1.9, 2.1, 1.6, 1.6, 1.8, 1.1, 0.5, 0.7, 1.2, 0.8, 
    0.9, 1.1, 0.8, 1.4, 0.9, 0.4, 0.9, 0.5, 1, 1.2, 0.8, 1.7, 1.9, 2.9, 1.2, 
    1, 2.3, 0.8, 1.8, 1.4, 1.5, 2.5, 0.6, 0.7, 0.7, 1, 0.8, 0.9, 1, 0.7, 1, 
    0.2, 1, 0.3, 0.7, 0.6, 0.6, 0.6, 0.2, 1.1, 0.7, 1.1, 0.6, 0.4, 0.9, 0.9, 
    0.5, 0.3, 0.3, 0.7, 0.1, 0.7, 0.4, 0.1, 0.8, 0.5, 0.6, 0.5, 1, 1, 0.8, 
    0.6, 1.6, 1.2, 0.9, 1.7, 1, 0.3, 1.3, 0.2, 1.3, 1.9, 4.3, 1.9, 0.8, 1.2, 
    0.9, 0.6, 1.3, 1.1, 1, 0.4, 1.1, 1.1, 1.1, 1.4, 1.4, 1.5, 0.4, 0.7, 1.5, 
    0.6, 0.5, 0.6, 0.3, 1.7, 1.7, 1.5, 0.8, 0.5, 0.6, 1.2, 1.4, 0.7, 1, 1, 
    1.6, 1.5, 1.2, 2, 0, 0.9, 1.5, 0.6, 0.7, 1.6, 0.9, 0.2, 1.1, 1.3, 0.9, 
    0.2, 0.9, 0.6, 0.8, 0.8, 0.3, 0.5, 0.6, 2.4, 1.5, 1.2, 0.9, 0.9, 0.2, 
    1.3, 0.5, 0.8, 1.4, 0.4, 0.5, 0.5, 1.9, 5, 5.7, 5.3, 6, 5.9, 3.3, 6, 6.7, 
    5.2, 7.8, 7.3, 7.6, 7.3, 6.2, 6.2, 6.5, 6.9, 6.1, 6.1, 6, 5.7, 2.5, 2.5, 
    0.3, 1.6, 2.1, 1.9, 2.2, 2.2, 1.2, 0.7, 0.4, 0.9, 1, 0.5, 1.4, 0.6, 1.7, 
    1, 0.6, 7.5, 7.7, 4.7, 4.6, 4.6, 7.8, 8, 6.8, 4.2, 6.5, 8.5, 6.5, 6.5, 5, 
    1.7, 2.8, 3.6, 6.1, 5.4, 3, 2.8, 1.6, 1.7, 1.1, 1.7, 0.4, 0.3, 0.3, 1.6, 
    2.3, 0, 1.1, 0.8, 0.6, 1, 1, 0.7, 0.6, 0.3, 0.1, 0, 0.8, 0.7, 0.6, 0.6, 
    1.3, 0.9, 0.6, 0.3, 1, 1.8, 0.4, 0.4, 0.2, 1.1, 2, 2.9, 3.1, 3.2, 3.5, 
    1.4, 1.1, 1.2, 1.7, 0.2, 0.2, 0.6, 0.1, 0.5, 0.4, 0.3, 0.1, 0.1, 1, 0.9, 
    0.5, 0.2, 0.6, 0, 0.8, 0.4, 0.3, 1.4, 0.6, 0.4, 0.1, 0.7, 0, 0, 0, 0, 0, 
    0, 0, 0.4, 0, 2.8, 5.5, 4.7, 3.1, 3, 1.9, 0.3, 0.3, 1.1, 0.9, 0.3, 1.9, 
    0.8, 1.1, 0.9, 0, 2.7, 2.6, 1.2, 0.8, 1.2, 0.5, 0.5, 0.8, 0.9, 1.3, 0.5, 
    0.8, 0.6, 0, 0.8, 1.4, 5.4, 7.9, 5.8, 4.3, 3.4, 2, 0.6, 2.9, 1.1, 1.3, 
    0.7, 1.6, 1.9, 0.5, 0, 0, 0, 0.5, 6.2, 8, 4.1, 6.8, 6.7, 7.9, 10.1, 9.8, 
    7.4, 8, 7.7, 8.3, 12.6, 11.5, 10, 8, 6.8, 7, 9.1, 7.6, 7.8, 6.7, 6.2, 
    4.6, 3.9, 4.3, 4, 2.7, 2.9, 1.1, 0.3, 0.7, 1.4, 0.7, 1, 1.4, 0.4, 0.4, 
    0.2, 0.4, 0.3, 1.1, 0, 0.6, 0.8, 0.4, 0.3, 0.1, 0.4, 0.5, 0.7, 0, 0.1, 
    0.8, 1.8, 1.5, 1.6, 1.7, 1.2, 1.6, 2.2, 2, 2.1, 2, 2.4, 2.3, 1.5, 2.1, 3, 
    4.1, 4.2, 3.5, 4.5, 5.4, 5.5, 5.1, 5.3, 4.3, 3.4, 4.3, 4.2, 3.7, 4.8, 
    5.1, 5.1, 6.9, 5.4, 5.6, 5.6, 6.8, 7.3, 6.6, 7.6, 5.7, 5.2, 5.1, 4.8, 
    5.5, 6.7, 6.1, 6.1, 5.9, 5, 4.8, 4.7, 4.8, 5.2, 4.6, 5.2, 6.3, 5.3, 6.8, 
    6, 5.9, 7.7, 5, 5.7, 6.9, 4.2, 5.4, 6.4, 6.3, 6.1, 8.4, 9.3, 8.2, 6.8, 
    2.3, 2.9, 5.1, 6.7, 3.3, 2.1, 3.3, 2.8, 1.9, 1.7, 3.5, 2.8, 2.7, 3.5, 4, 
    3.6, 4, 3.5, 2.8, 3, 2.7, 3.2, 1.9, 4.1, 3.2, 4, 4.5, 3.7, 4.5, 5.3, 5.6, 
    6, 5.4, 5.4, 5.4, 5, 4.2, 5, 5.2, 5.1, 3, 1.9, 2.5, 3.4, 2.5, 3.3, 6, 
    5.5, 5.7, 4.6, 4.9, 2.2, 1.5, 1.3, 1.4, 1.2, 1.2, 1.3, 1.5, 1.7, 1.8, 
    1.7, 1.7, 1.6, 1.9, 1.8, 1.5, 2, 1.7, 1.9, 2.2, 3.3, 2.5, 1.8, 1.8, 2.4, 
    2.6, 2.9, 2.7, 1.6, 1.4, 2.1, 1.2, 0.5, 0.8, 1.1, 3.3, 1.7, 2.1, 2.5, 
    2.6, 3.9, 2.8, 2.8, 2.9, 3.4, 3.9, 3, 3.4, 2.5, 2, 2, 2.4, 0.8, 0.3, 0.3, 
    0.8, 1.3, 2.7, 3.2, 3.7, 3.1, 3.6, 4.1, 4.3, 4.2, 4, 3.9, 3.8, 4.2, 4.7, 
    3.4, 3.4, 3.4, 3.7, 3.6, 3.4, 3, 1.4, 1.2, 3.7, 2.9, 3.8, 4.4, 4.6, 4.4, 
    4.2, 2.5, 2, 1.7, 1.9, 2.9, 2.2, 2.1, 2.5, 2.9, 2.9, 1.8, 1.8, 2.8, 2.7, 
    2.1, 1.7, 2.5, 2, 1, 1.3, 1.3, 1.9, 2.9, 3.7, 3.2, 3.5, 4.1, 2.9, 1.8, 
    3.3, 3.8, 3.6, 4.1, 5.9, 4.9, 5.7, 7.2, 4.6, 4.2, 4.7, 4.1, 3.1, 5.5, 
    6.1, 6.4, 5.3, 3.9, 3.3, 3.5, 2.9, 1.6, 2.3, 3.3, 2.2, 2.3, 5.3, 4.6, 
    2.4, 3.8, 4.3, 5.3, 4.6, 3.2, 2.5, 1.5, 1, 1.2, 1.1, 0.7, 0.9, 1.5, 2.2, 
    1.2, 1.3, 1.6, 1, 0.9, 1.4, 1.2, 1.4, 1.9, 1.8, 1.4, 1.2, 1.2, 1.5, 1.4, 
    1.5, 0.9, 0.9, 0.8, 1.3, 2.5, 3.3, 4.4, 4.4, 4, 4.5, 4.3, 4.7, 3.7, 2, 
    1.4, 3.3, 5.8, 4.9, 1, 3.4, 1.1, 1, 1.4, 1.5, 1.6, 1.8, 1.4, 1.1, 1, 0.9, 
    2.1, 1.6, 1.3, 1.4, 1.4, 1.3, 1.2, 1, 1, 1.8, 2, 2.4, 0.8, 1.6, 3.3, 3, 
    2, 2.2, 2.7, 3.7, 3.6, 3.7, 5.6, 3.7, 3.6, 3.4, 3.7, 3.1, 2.7, 3.2, 3.9, 
    3.4, 2.1, 2.3, 2.1, 3.1, 1.2, 2.9, 1.9, 1.4, 1.5, 2, 1.7, 1.9, 1.7, 1.6, 
    1.4, 1.2, 1, 2.6, 2.3, 2, 1.9, 1.5, 1.3, 1, 1.3, 2.2, 1.7, 1.3, 1.4, 1.8, 
    2.3, 2, 1.6, 1.2, 1.2, 1.2, 1.8, 4, 3.6, 2.2, 1.9, 1.8, 2.3, 2.5, 2.9, 
    3.2, 3, 2, 1.5, 1.9, 1.8, 1.7, 1.2, 1.7, 1.7, 1.7, 1.4, 2, 2, 1.8, 2, 
    2.6, 3.4, 2.1, 1.4, 1.8, 1.7, 1.4, 1, 0.8, 1.1, 1.8, 2, 1.6, 1.2, 2.3, 
    1.8, 1.5, 1.3, 1.9, 1.9, 1.9, 2.2, 3, 3, 2.8, 3.1, 2.5, 3, 1.9, 2.4, 2.2, 
    1.8, 2, 1, 1.4, 1.9, 0.7, 0.5, 1.9, 1.5, 3.1, 4, 4.6, 5.3, 6.1, 4.6, 5.7, 
    6.2, 6.8, 6.8, 5.5, 4.6, 4.7, 3.8, 9.6, 9.4, 7, 4.2, 9.8, 9, 8.6, 7, 6.4, 
    3.3, 4.4, 9.1, 7.5, 6.9, 9.7, 12.4, 10.9, 16.4, 19.3, 18.1, 18.5, 17, 
    17.1, 15.9, 16.3, 13, 11.5, 9.4, 8.7, 7, 5.9, 5.4, 5.8, 5.7, 4.5, 2.7, 
    5.5, 6.3, 6.8, 7, 6.5, 7, 6, 5.6, 5.3, 7.7, 6.2, 4.2, 2.5, 2.4, 1.9, 2.5, 
    3.9, 3.5, 2.4, 4.7, 6.2, 5.1, 4.9, 5.4, 5.2, 5.3, 5.8, 4.5, 3.1, 3.3, 
    4.6, 4.2, 2.5, 1.1, 4.1, 4.3, 3.3, 2.1, 2, 2.5, 4.1, 2.2, 1.7, 1.4, 1.5, 
    1.9, 2.2, 2.5, 2.3, 2.2, 3.2, 4.7, 4.5, 3.9, 3.8, 8.7, 10.1, 9.2, 8.7, 
    7.8, 7.4, 6.6, 4.9, 3.5, 3.2, 1.4, 1.4, 1, 1.3, 1.5, 1.4, 1.5, 1.6, 1.5, 
    1.7, 2.1, 5.8, 4.4, 4.1, 2.9, 2.4, 3.3, 2.5, 0.6, 2.4, 1.9, 2.4, 3, 2, 
    1.1, 1.6, 3.2, 1.4, 2.7, 2.8, 2.8, 4.2, 3.3, 3.3, 4, 10.9, 6, 4.2, 3.4, 
    5.1, 1.2, 1.3, 4.5, 4.1, 4.8, 7.5, 6.8, 9.3, 7.5, 6.7, 3.3, 2.4, 1.8, 
    2.7, 2.2, 4.9, 13, 11.5, 7.9, 4, 5.4, 5.4, 7.4, 7.7, 5.1, 4.1, 1.5, 7.2, 
    6.4, 10.8, 10.4, 9.1, 7.6, 6.9, 5.3, 4.5, 5.6, 5.1, 4.3, 4.2, 5, 4, 2.2, 
    2.5, 1.9, 1.7, 1.9, 2, 1.1, 1.5, 1.7, 2, 1.7, 1.2, 1.5, 1.5, 1.7, 1.8, 
    1.4, 0.6, 3.6, 5.1, 5, 5.9, 7, 6.7, 6.3, 5.7, 5.9, 6.1, 6.3, 6.6, 5.9, 
    4.3, 3.2, 3, 4.2, 4.9, 4.5, 4.2, 6.2, 6.8, 5.4, 4.2, 5.9, 4.1, 1.4, 1, 
    0.8, 0.5, 0.5, 0.5, 0.2, 0.5, 0.2, 0.3, 0.4, 0.8, 0.7, 1.3, 0.8, 1.1, 
    0.7, 0.5, 0.6, 0.7, 0.7, 0.8, 0.6, 0.8, 0.8, 0.9, 0.7, 0.5, 0.5, 0.5, 
    0.5, 0.6, 0.6, 0.6, 1.1, 1.1, 1.4, 0.8, 0.5, 0.3, 0.3, 0.4, 0.8, 1.5, 
    1.6, 1.6, 1.4, 1.1, 0.7, 0.7, 0.8, 0.8, 0.9, 0.9, 1.1, 1.7, 1.5, 1.4, 
    1.5, 1.5, 1.2, 1.1, 1.1, 1.2, 1.2, 1.3, 1.4, 1.3, 1.2, 1.2, 0.9, 1.3, 
    1.6, 1.4, 1.3, 1.4, 1.3, 1.3, 1.3, 1.4, 1.4, 1.4, 0.9, 1.1, 1, 0.8, 0.8, 
    0.7, 0.8, 1.6, 1.8, 1.8, 1.8, 1.9, 1.7, 1.4, 1.9, 2.2, 2.4, 2.6, 2.8, 
    2.5, 2.3, 2.1, 1.9, 1.7, 1.6, 1.7, 2.1, 2.2, 1.9, 2.2, 2, 1.8, 1.7, 1.4, 
    1.2, 1.4, 0.7, 0.8, 0.7, 1, 1, 0.9, 0.9, 1.1, 1, 1, 0.9, 1, 1.2, 0.7, 
    0.8, 1.2, 1.1, 1.1, 1.1, 1.2, 1.2, 1.3, 1.6, 2.2, 1.7, 1.7, 1.6, 1.2, 
    1.8, 1.5, 1.4, 1.5, 1.6, 1.2, 1.3, 1.3, 1.3, 1.3, 1.5, 1.4, 1.5, 1.2, 
    1.5, 0.9, 0.9, 0.7, 0.9, 0.9, 2.2, 1, 1.9, 1, 1.5, 2.3, 2.9, 5.2, 2.3, 
    1.6, 1.1, 1.2, 1.6, 1.8, 1.6, 2.1, 2, 1.8, 2, 1.8, 1.4, 1.3, 1.2, 1.1, 
    1.3, 1.6, 2.6, 1.7, 1.3, 1.3, 1.1, 1.2, 1.6, 1.6, 2, 1.4, 2, 1.9, 1.6, 
    2.1, 1.9, 1.9, 1.5, 1, 1.7, 1.9, 2.6, 2.4, 2.9, 1.3, 1.3, 2.1, 5.4, 6.7, 
    6.9, 6.2, 6.9, 7.3, 8.6, 8.8, 10.1, 11.3, 11.5, 10.6, 10.5, 10, 9.2, 8.8, 
    8.5, 8.9, 7.6, 6.3, 3.4, 3.9, 4.5, 5.1, 6.4, 6.1, 3.7, 3, 2.7, 2.9, 3.2, 
    2.4, 2.3, 1.1, 1, 1.1, 2.5, 1.7, 0.9, 0.4, 0.5, 0.4, 0.5, 0.7, 1.1, 0.7, 
    1.3, 1.5, 1.5, 1.5, 2, 2.6, 2.2, 2.2, 2.2, 2, 1.3, 1.3, 1.1, 2, 2, 1.5, 
    1.8, 1.5, 0.8, 0.5, 3.3, 4.9, 1.7, 9.9, 12.7, 14, 13.5, 13, 12.6, 12.5, 
    11.1, 9.5, 8.9, 8.3, 6.6, 7.1, 7.6, 8.1, 7.9, 4.6, 9.9, 11.1, 10.4, 11, 
    11.3, 12.1, 11.7, 11.4, 11.5, 11.1, 10.5, 8.4, 8.5, 8.8, 9.3, 7.5, 6.7, 
    6.6, 7.8, 7.2, 7.5, 7.9, 9.9, 11.5, 12.1, 11.6, 11.7, 11.2, 10.8, 8.7, 
    12.3, 12.6, 13.2, 12.9, 12.3, 9.5, 7.8, 6.9, 6.2, 7.8, 9.2, 9, 8.1, 8, 
    7.5, 7.2, 6, 3.9, 0.3, 1.2, 1.7, 2.3, 4.4, 3.8, 4.4, 5.2, 5, 4, 4, 3.8, 
    4, 5.3, 4.4, 3.9, 2.1, 0.7, 1, 0.2, 0.5, 1.1, 0.8, 0.8, 0.6, 0.5, 0.2, 
    0.2, 0.5, 0.6, 0.9, 1.1, 1.7, 0.9, 1.5, 1.5, 1.2, 0.8, 2.7, 0.8, 1.2, 
    1.6, 0.4, 1.6, 1.1, 0.9, 1.3, 1.1, 0.4, 0.3, 1.2, 2.5, 0.6, 0.4, 1.8, 
    3.5, 2.7, 1.9, 2.9, 1.5, 0.7, 0.2, 0.4, 0.2, 0.6, 0.6, 0.7, 3.5, 1.8, 
    0.6, 0.9, 1.5, 1.2, 0.5, 1, 0.9, 1, 1.3, 0.7, 0.6, 1.3, 1.5, 1.3, 2.2, 
    1.5, 1.2, 1.3, 2.8, 3.5, 2.6, 2.3, 1.3, 1.6, 0.9, 0.5, 0.5, 0.7, 0.5, 
    1.6, 0.8, 0.8, 0.7, 0.7, 0.2, 1.3, 1.7, 0.9, 0.3, 1.5, 1.3, 1.2, 1.5, 
    0.5, 0.8, 1.7, 1.5, 1.1, 1.6, 2, 1.5, 0.5, 0.2, 0.2, 0.2, 0.4, 0.5, 0.6, 
    1.3, 0, 1, 0.9, 0.5, 0.3, 0.8, 0.5, 0.7, 1.1, 0.7, 1, 1.1, 0, 0.1, 0.6, 
    0.9, 0.5, 0.4, 1.1, 0.7, 0.3, 1.1, 1.1, 1.3, 0.4, 0.1, 0.9, 0, 0, 0.8, 
    0.2, 0.9, 0.5, 0.6, 0.6, 0.9, 0.5, 0.8, 0.6, 0.1, 0, 1, 0.2, 1.1, 0.2, 
    0.4, 0.1, 0.5, 0.1, 0.6, 0, 0.3, 0.8, 0, 0.4, 0.2, 0.1, 0.4, 0.4, 0.6, 
    0.2, 0.5, 0, 0.4, 0.7, 1.1, 0, 0, 0.6, 0, 0.4, 0.5, 0.1, 0.6, 0.7, 0, 
    0.1, 0.5, 0.7, 0, 0.4, 0.1, 0.1, 0, 0, 0.3, 0.1, 0, 0, 0.1, 0.4, 1.3, 
    0.1, 0.3, 0, 0.4, 0.2, 0.4, 0.1, 0, 0.8, 0.5, 0.5, 0.3, 0.1, 0.1, 1.8, 
    0.2, 1.3, 0.4, 0.2, 0.6, 1, 0.1, 0, 0.1, 0.3, 0.1, 0.5, 0.4, 0.7, 0, 0.8, 
    0.9, 0.9, 0.8, 0.3, 0.5, 0.1, 0.1, 0.2, 0.5, 0.2, 1.5, 0.9, 1, 0.3, 0.1, 
    0.1, 0.2, 0.1, 0.5, 1, 0.9, 0.7, 0.2, 0.1, 0.2, 0.1, 0.7, 0.4, 0, 0.8, 
    0.7, 0, 0.5, 0.1, 0.6, 1, 0.2, 0.5, 0.8, 1.4, 0.3, 0, 0.1, 0, 0.2, 0, 0, 
    0.8, 0.2, 0.5, 0, 1, 0.5, 0, 0.2, 0.3, 1.4, 1.8, 0.1, 0, 1.5, 0.7, 0.4, 
    0.3, 0.1, 0, 0.4, 0.2, 0, 0.1, 0.3, 0.4, 0.5, 0.1, 0.4, 0.3, 1.3, 0.5, 
    0.7, 1.1, 0.3, 0.3, 1.5, 1.4, 1.5, 0.4, 0, 0.3, 0.5, 1.8, 0.1, 1.2, 0.9, 
    0.5, 0.5, 0.5, 0.5, 0.2, 0.3, 0.3, 0.6, 0.2, 0.2, 0.5, 0.5, 0.2, 0.5, 
    0.8, 1.2, 1, 0, 1.1, 0.5, 0.5, 1.1, 0.7, 0.6, 0.6, 0, 0.5, 0.4, 0.3, 0.2, 
    0.1, 0.2, 0.3, 0.8, 0.4, 0.4, 0.3, 1, 0.8, 0.2, 0.7, 1.7, 0, 0.3, 0.5, 
    0.8, 0.5, 0.2, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 6.5, 5.7, 5.9, 7.4, 7.9, 9.7, 
    8.8, 9.7, 9.6, 10.9, 11.1, 10, 10.1, 7.9, 11.8, 11.5, 11.6, 11, 10.9, 
    12.3, 11.1, 11.7, 16.2, 15.8, 14.6, 14.5, 12.4, 11.1, 12.5, 10.7, 8.9, 
    9.1, 9.2, 8.7, 8.4, 7.1, 7, 6.3, 7.5, 7, 6.6, 4.6, 4.7, 3.3, 1.6, 2, 1.9, 
    1.1, 1.4, 0.8, 1.5, 1.1, 1.5, 3.7, 2.1, 3.1, 3, 1, 0.4, 0.2, 1.4, 0.8, 
    0.8, 0.1, 0.3, 0.4, 0.2, 0.4, 1.1, 0.5, 0.6, 0.8, 1.4, 0.5, 0.3, 0.3, 
    0.4, 0.5, 0.5, 0.6, 0.5, 0.8, 1.3, 1.2, 1.3, 1.3, 1.4, 1.2, 1.8, 1.2, 
    1.1, 1, 0.8, 0.7, 1.6, 1.5, 1.7, 0.9, 1.3, 1.7, 1.1, 0.8, 1.6, 1.2, 0.8, 
    0.5, 1.8, 0.8, 0.9, 0.7, 0.7, 0.7, 0.7, 0.7, 0.2, 0.5, 0.5, 0.3, 0.4, 
    0.5, 0.4, 0.8, 0.9, 0, 1.2, 1.3, 1.2, 4.6, 4.9, 3.6, 1.8, 1.3, 3.4, 4.1, 
    3.2, 0.8, 1.8, 3.3, 2.7, 1, 1.2, 6.3, 6.9, 1.6, 3.9, 7.5, 2.5, 2.3, 2, 
    2.6, 2.5, 2.7, 3.4, 1.9, 2.8, 5.3, 4.3, 3.5, 3.6, 3.8, 3.6, 2.1, 1.9, 
    1.3, 1.6, 1.3, 2, 2.9, 3.9, 1.1, 1.5, 2.4, 1.8, 1.1, 1.5, 1.5, 1.5, 2.1, 
    2.7, 1.9, 1.4, 3.5, 2.4, 5.7, 4.1, 2.9, 0.4, 1.6, 0.5, 1.9, 0.5, 0, 1.5, 
    0.6, 0.9, 0.9, 0.6, 1.2, 0.6, 1.3, 2, 0.9, 0.6, 0.1, 1.5, 0.6, 0.5, 0.7, 
    0.8, 0.6, 0.6, 0.6, 1.6, 5.2, 1.4, 1.8, 2.6, 2.9, 2.3, 1.8, 4.5, 3.3, 
    3.3, 1.6, 2.1, 1.7, 1.1, 0.3, 0.5, 2.2, 0.8, 0.7, 1.6, 1.3, 0.4, 0.8, 
    0.6, 1.1, 1.4, 1.6, 0.3, 0.8, 0.2, 0.8, 1.1, 2.9, 1.5, 1.6, 0.3, 0.4, 
    0.5, 0.2, 1.1, 1.1, 0.2, 0, 0.1, 1, 0, 0.4, 0.4, 1, 0.9, 0.6, 0, 0.7, 
    0.1, 0.5, 0.6, 1.5, 2.9, 3.4, 3.6, 3.3, 2.8, 2.4, 1.4, 1.4, 0.8, 0.3, 
    0.3, 0.1, 0.3, 0.6, 0.3, 0.4, 0.4, 0.8, 0.5, 0, 0.4, 0.1, 0.8, 0.8, 0.4, 
    0.6, 0, 0.8, 0.8, 0, 0.3, 1.1, 0.1, 0.1, 0.6, 0.8, 0.3, 0.3, 0.6, 0, 0.3, 
    1, 0.2, 0.8, 0.9, 0.4, 0.3, 1, 0.1, 1.2, 1, 0.3, 1.7, 1.8, 1.6, 1.4, 0.6, 
    0.2, 0.4, 0.1, 0.6, 0.1, 0.6, 0.2, 0.1, 0.6, 0.3, 0.1, 0.7, 0.3, 0, 1, 
    0.9, 1.8, 1.6, 1.4, 1, 1, 1, 1, 0.7, 0.4, 0.2, 0.3, 0.7, 1.5, 1.3, 1, 
    0.8, 1, 1.9, 4.7, 5.7, 5.3, 2.5, 1.7, 2, 1.2, 2.3, 1.5, 0.1, 0.7, 0.9, 
    0.3, 1, 0.3, 0.5, 1.2, 0.4, 0.5, 0.1, 0, 0, 0.1, 0.2, 1.4, 0.8, 0.5, 1.4, 
    0.9, 0.3, 0.6, 0.6, 0.4, 0.2, 1, 0.1, 0.6, 0.3, 0.5, 0.2, 1.1, 1.2, 1.1, 
    0.3, 1.2, 0.1, 1.2, 0.5, 1.2, 0.6, 0.8, 1.2, 0.7, 0.2, 0.7, 1.8, 0, 0.8, 
    0.4, 0.5, 0.5, 0.9, 0.5, 0.4, 0.9, 1.3, 0.9, 1, 1, 0.9, 0.8, 0.7, 0.2, 
    0.4, 0.4, 1, 0.8, 0.5, 0.9, 1.3, 0.5, 0.3, 1.1, 1, 1.5, 0.3, 0.2, 0.5, 
    0.5, 0.1, 0.1, 0.2, 0, 0.1, 0, 1.5, 0.3, 0.5, 0.7, 1.3, 0.1, 0.6, 0.1, 
    0.8, 1, 0, 1.4, 0.3, 0.5, 0.4, 0.1, 0.4, 0, 0.5, 0.7, 0.3, 0.1, 0.5, 0.2, 
    0.3, 0.6, 1.1, 1, 0.4, 0.3, 0.1, 0.4, 0.8, 0.8, 0.5, 0.1, 0.2, 0.5, 1.8, 
    1, 0.8, 0.2, 0.5, 0.6, 0.5, 0.5, 0.5, 0.5, 0.4, 0.4, 0.4, 0.2, 2, 0.1, 1, 
    0.7, 0.3, 0.8, 0.7, 0.2, 0.7, 0, 0.7, 0.1, 0, 1.2, 0.3, 0.1, 0.7, 0.2, 
    1.6, 2, 1.4, 0.6, 0.1, 0.5, 0.3, 0.7, 0.4, 0.9, 0.2, 0.6, 0.1, 1, 0, 0.5, 
    0.9, 0.1, 0.3, 1.4, 0.3, 0, 0.5, 0.6, 1.1, 0.8, 0.3, 0.3, 0.6, 0.9, 0.8, 
    0.6, 1, 0.8, 0.9, 0.8, 0.2, 1.1, 1, 0.3, 6.7, 3.7, 4, 4.2, 3.7, 3.3, 4.1, 
    4.3, 0.8, 1.1, 0.7, 1.1, 1.2, 0.1, 1.1, 0.4, 1.1, 0.2, 0.3, 1.5, 0.1, 
    0.4, 0.9, 1, 0, 1.2, 0.6, 0.1, 0.6, 0.4, 0.1, 1.7, 1.3, 0.3, 1.8, 0.9, 
    0.8, 0.3, 1.7, 0.7, 2.2, 0.8, 3, 3.8, 2.8, 1.3, 1.6, 1, 0.1, 1.3, 0.4, 
    1.3, 1.2, 1.1, 0.5, 0, 0.1, 0.2, 0.2, 0.9, 0.9, 0.6, 0.9, 0.1, 0.9, 1, 
    1.3, 1, 1.1, 1.1, 2.4, 2.3, 2.3, 3.8, 6.3, 5.3, 4, 3.6, 3.8, 3.7, 3.2, 
    3.5, 3.8, 3.4, 3.2, 3.4, 3.5, 5, 2, 1.9, 0.5, 1.7, 0.8, 0.4, 3.1, 0.9, 
    1.6, 0.7, 0.6, 0.6, 0.2, 1.3, 0.9, 0.1, 0.8, 0.5, 0.1, 0, 1.4, 0.2, 0.7, 
    0.8, 0.9, 1.1, 0.1, 0.2, 0.2, 1.4, 0.7, 0, 0.8, 0.2, 0.3, 2.4, 4.8, 4.3, 
    1.6, 0.8, 0.5, 1.8, 0.6, 0.8, 1, 0.5, 0.5, 0.2, 0.9, 0.7, 0.8, 1, 1, 0.5, 
    0.1, 1.4, 0, 2.2, 1.3, 0.7, 1.1, 1, 1.8, 0.1, 0.1, 0.7, 1.2, 0.6, 0.3, 0, 
    0.1, 0.9, 0.9, 0.3, 0.2, 0.2, 0.8, 1.3, 0.1, 0.2, 0.9, 0, 0, 0.2, 0.6, 0, 
    0.1, 0.2, 1.5, 0.1, 2.2, 5.5, 2.3, 2.1, 5.9, 3.7, 1.7, 1.7, 2, 0.2, 4.9, 
    7, 4.8, 1.5, 4.3, 4.5, 5.7, 1.8, 0.8, 0.8, 3, 4, 1.8, 2.5, 3.7, 1, 2.4, 
    2.8, 1.6, 2.1, 1.3, 2.4, 1.9, 0.7, 3, 2.7, 1.3, 1.1, 0.8, 1.7, 0.5, 0.9, 
    0.2, 1.2, 0.8, 0.6, 0.6, 0.9, 0, 1.3, 0.5, 0.2, 1, 0, 0.3, 0.8, 0, 0.4, 
    0.1, 0.6, 0.3, 0.9, 0.4, 0.7, 0, 0.5, 1.3, 0.6, 1.3, 0.1, 0.7, 0.8, 1.1, 
    0.5, 0.3, 0.5, 0.5, 1.3, 0.1, 0, 1.3, 1.1, 0.4, 0.4, 0.4, 0.6, 0.3, 0.6, 
    0.7, 0.8, 0.1, 0, 0, 0.3, 0.1, 0.2, 0.6, 0.2, 0.1, 0.8, 0.4, 0.2, 0.5, 
    0.2, 0.8, 5.4, 5, 3.7, 3.4, 5.4, 4.8, 3.1, 1.6, 3.5, 3.6, 4.1, 4.1, 0.7, 
    3.1, 3.2, 0.2, 0.8, 1.2, 0.8, 0.8, 0.1, 0.2, 0, 0, 0.6, 0.9, 1.6, 1, 0.3, 
    2.5, 0.1, 0.7, 0.3, 0.2, 0, 0.8, 0.5, 0.1, 0.7, 0.2, 0.1, 0.5, 0, 0, 0.1, 
    0.9, 0.7, 0.3, 0.5, 1.8, 2, 5.9, 6.4, 5.5, 5.5, 5.2, 4.6, 3.4, 2.6, 2.3, 
    1.4, 0.6, 0.4, 0.5, 0.7, 1, 0.9, 0.5, 2, 1.7, 2.1, 1.5, 2.2, 2.8, 2.5, 
    0.5, 0, 0.7, 0.5, 0.5, 1.4, 0.3, 0.8, 0.8, 0.3, 0.6, 0, 0.7, 0.2, 0.2, 
    0.2, 0.3, 0.8, 0.4, 0.7, 0.7, 0.6, 0.4, 0.2, 0.7, 0.3, 0, 0.2, 0, 0.2, 
    0.6, 0.6, 0.6, 0, 0.1, 0.4, 0.8, 0.4, 0.3, 0.5, 0.6, 0.1, 0, 0.4, 0.2, 0, 
    1.5, 1.2, 1.5, 0.1, 0.2, 0.2, 0, 0.1, 0.1, 0.2, 0.7, 0, 0.1, 0.1, 0.5, 
    0.8, 0.9, 0.5, 0.1, 0.6, 0.2, 0, 0.2, 0.8, 0.1, 1.1, 0.3, 0.3, 0.3, 0, 
    0.2, 0.5, 0.4, 0.2, 0.2, 0.5, 0.4, 0.3, 0.3, 0, 0.4, 2.4, 1, 0.4, 1.3, 
    2.1, 1.2, 2.5, 1.5, 0.7, 0.2, 0, 0.6, 0.2, 0.9, 0.3, 0.4, 0.4, 0.2, 0.3, 
    0.7, 0.2, 0.6, 0.5, 0.5, 0.8, 0.9, 0.7, 0.7, 0.1, 0.8, 0.1, 0.6, 0.7, 
    0.2, 0.3, 0.3, 0.9, 0.7, 0.5, 1.4, 0.5, 0, 0.2, 0.4, 3, 1.5, 0.8, 0.4, 
    1.4, 0, 0.8, 1.2, 0.8, 0, 0.5, 0.4, 0.1, 0, 0.5, 0, 0.2, 0.4, 0.5, 0.1, 
    0, 0.2, 0, 0.5, 0, 0.4, 0.2, 1.2, 0.8, 0.8, 0, 0.8, 0.6, 1.1, 0, 0.5, 
    0.7, 0, 1.2, 2.1, 0.1, 0.7, 1.3, 0.3, 0.5, 0.1, 0.2, 0.3, 0.6, 0.6, 0.9, 
    1.1, 0.5, 0.7, 0.1, 0.5, 0.3, 0.7, 0.9, 1.2, 0.9, 1.7, 0.3, 1.1, 1.3, 
    0.4, 0.4, 0.5, 1.3, 0.5, 0.4, 0.5, 1, 0.4, 0.5, 1.5, 2.8, 0.7, 2, 1.4, 
    2.2, 0.6, 1.5, 0.4, 1.2, 0.6, 1.8, 2.9, 4.4, 6.7, 4.3, 4.9, 4.6, 4, 4.4, 
    3.9, 2.4, 3, 3.7, 5.9, 3.2, 2.6, 2.7, 1.2, 1.7, 1.8, 4.4, 3, 2.8, 3, 3.4, 
    2, 0.8, 0.7, 1.6, 0.6, 0.6, 0.5, 0.7, 1.7, 0.2, 1.2, 0.3, 1.6, 0.9, 0.2, 
    1, 1.3, 1.8, 2.8, 1.4, 3.1, 1.3, 1.5, 1.4, 1, 8.1, 1.8, 3.2, 2.4, 0.1, 
    2.6, 2.7, 0.8, 0.8, 0.1, 0, 0.5, 1.2, 0.8, 0.5, 6, 5.9, 4.6, 5.3, 4, 1.5, 
    0.6, 1.2, 1.5, 1.5, 1.7, 2, 1, 5.3, 5.2, 4.5, 4.9, 4.7, 4.3, 3.7, 4.3, 
    4.7, 5.3, 3.9, 4.3, 4.1, 2.6, 3.1, 0.6, 0.7, 0.2, 2.6, 2.2, 1.9, 1.2, 
    1.2, 1.8, 2, 1.5, 1, 0.3, 1.2, 1.2, 1.2, 0.9, 0.4, 1.3, 0.7, 0.5, 1.3, 
    1.2, 5.3, 3.2, 4.8, 6.1, 3.5, 5.3, 4.1, 4.5, 4.7, 3.6, 4.9, 2.7, 2.6, 
    1.9, 1.5, 1.6, 1.8, 0.6, 0.3, 2, 1.2, 1, 6.6, 7.4, 7.4, 5.2, 7, 7.3, 6.5, 
    7.6, 7, 7.9, 5.6, 3.4, 3.2, 1, 1.4, 0.9, 1.6, 1.5, 1.9, 2.7, 1.1, 0.8, 
    0.7, 0.3, 1.6, 3, 3.4, 2.9, 2.2, 1.8, 1.9, 3.2, 1.5, 2.7, 0, 0.9, 1.5, 
    0.6, 0.2, 0.3, 0.3, 0.1, 0, 0.7, 1.1, 0.6, 0.5, 0, 0.7, 2.8, 2.5, 3.6, 
    1.1, 0.4, 0.5, 0.6, 1.2, 2.7, 0.1, 0, 0, 0, 0, 2.1, 0.8, 0.6, 0.1, 0.4, 
    4.6, 5.2, 3.8, 3.6, 3.3, 0.9, 0.6, 0, 1.1, 0.8, 1.1, 1, 0.3, 1.4, 1.1, 
    0.1, 0.9, 1, 0.9, 0.5, 1, 0.2, 1.4, 1, 0.6, 2.3, 2.7, 0.4, 0.2, 1.6, 2.9, 
    5, 5.9, 9.6, 4.8, 5.1, 4, 5, 3.9, 3.9, 4.8, 2.5, 1.1, 1, 1.4, 1.5, 1.8, 
    0.4, 2.7, 1.8, 1.5, 1, 1.2, 1.1, 0.6, 1.9, 1.1, 1.4, 1.8, 2, 1.7, 0.1, 
    0.8, 0.2, 0.8, 0.4, 0.1, 0.3, 2.6, 0.1, 0.8, 0.7, 1.5, 0.1, 1.3, 0.4, 
    1.4, 1.4, 1.1, 0.8, 0.7, 0.8, 1.5, 0.7, 0.5, 0.4, 1.9, 1.8, 0.6, 0.2, 
    1.8, 1.9, 1.5, 1.4, 1.3, 2.2, 0.6, 0.7, 0.5, 0.7, 0.1, 0.2, 0.3, 0.8, 
    0.3, 0.3, 1.1, 0.8, 0, 0.4, 2.1, 5.3, 5.4, 4.8, 5.2, 7, 7.5, 8.3, 7.3, 
    9.5, 10.2, 10.9, 8.7, 7.4, 5.5, 6, 7.4, 7.4, 4.9, 4.1, 1.3, 1.7, 3.1, 
    1.2, 2.5, 2.3, 1.5, 1.2, 0.8, 0.5, 0.4, 0.9, 1.6, 3.1, 2.3, 3, 2, 1.9, 
    1.1, 0.7, 0.9, 0.7, 1.1, 1.4, 1.2, 0.6, 3.2, 3, 3.5, 3.7, 3.5, 2.1, 3.5, 
    3.4, 4.3, 4.9, 5.2, 6.1, 5.7, 4.9, 5.1, 3.8, 3.9, 3.2, 2.8, 1.9, 2.2, 
    1.6, 2.1, 3.1, 2.9, 1.6, 0.6, 1.1, 0.7, 0.5, 0.2, 1.1, 1.8, 1.2, 0.7, 
    0.8, 1.1, 0.8, 1.4, 1.9, 1.4, 1.1, 1.2, 1.7, 2.3, 4.2, 4.7, 5.2, 1, 5, 
    5.2, 5, 4.9, 5.6, 2.8, 4.3, 4.4, 4.2, 6.1, 4.3, 4.7, 5.7, 4.6, 3.5, 3.7, 
    3.5, 3.6, 4.5, 4, 3.1, 3.8, 3.4, 3.2, 3.2, 3.2, 3.2, 3, 2.8, 1.7, 1.7, 
    0.5, 0.7, 0.6, 0.9, 0.9, 1.2, 0.8, 0.7, 1.5, 1.5, 1.5, 1.9, 1.4, 2, 2.3, 
    1, 1.3, 1.3, 0.8, 0.8, 1.2, 1.2, 1.2, 0.7, 1.2, 0.9, 0.2, 0.9, 0.6, 4.5, 
    5.8, 5.3, 4.4, 4.6, 3.7, 3.7, 3.1, 3.5, 2, 0.5, 2.4, 0.8, 2.2, 0.1, 2.2, 
    1.6, 0.4, 1.3, 2.1, 2.4, 2.5, 2.9, 1.2, 2, 2.1, 3.1, 0.7, 0.8, 1.6, 1, 
    0.4, 2.4, 0.6, 0.3, 1.4, 1.4, 1.3, 1.4, 1.4, 1, 3.9, 0.8, 0.2, 1.5, 1.1, 
    1.7, 0.8, 1.2, 2.5, 3.3, 2.5, 3.7, 2.1, 3.6, 4.2, 6.6, 6.5, 5.6, 3.4, 
    5.5, 4.8, 4.2, 5, 5.2, 4, 4.8, 4.8, 4.8, 4.6, 4.5, 3.9, 3, 1.3, 1.1, 0.5, 
    3.9, 2.4, 2.6, 3.6, 3.8, 4.9, 3.9, 4.3, 3, 3.4, 2.9, 4.2, 5.2, 2.4, 2, 
    1.6, 1.6, 2.6, 2.9, 5, 4.9, 4.1, 4.2, 4.2, 3.8, 3.9, 2.2, 1.5, 1.3, 1.9, 
    1.6, 1.6, 1, 0.7, 1, 2.8, 2.5, 2.7, 1.3, 0.7, 0.3, 0.6, 1.1, 0.3, 0.5, 
    1.4, 1.3, 1.3, 1.1, 1.3, 1.5, 1.2, 1.1, 1.1, 1.1, 2.7, 2.3, 3.9, 3.7, 
    3.4, 4.2, 5.7, 6.5, 7.4, 6.8, 5.6, 6.2, 5.7, 6.1, 5.5, 6.4, 5.1, 4.4, 
    1.8, 1.4, 2, 0.2, 0.6, 0.7, 0.2, 0.2, 1, 1.9, 1.8, 0.9, 0.6, 0.8, 0.7, 
    0.6, 0.6, 1.2, 1.2, 1.1, 1.6, 3.5, 3.3, 3.5, 2.8, 2.9, 2.9, 1.3, 1.1, 
    1.8, 1.6, 0.9, 0.3, 0.3, 1.1, 0.1, 2.2, 0.3, 0.2, 0.4, 1.7, 1, 1.2, 0.7, 
    0.9, 0.7, 1.8, 3.1, 3.2, 5.2, 3.2, 3.1, 4, 3.9, 3.8, 2.6, 1.4, 1.3, 2.5, 
    2.2, 2.1, 0.9, 1.4, 1.1, 1.9, 1.2, 1.6, 1.2, 1.9, 2.2, 2.5, 1.7, 1.6, 
    1.6, 1.3, 3.1, 3, 3.8, 2.6, 1.8, 1, 1.3, 0.9, 1.7, 1.6, 1.6, 0.9, 0.6, 
    0.9, 1.3, 1.9, 1.2, 1.1, 0.8, 0.8, 0.6, 1.6, 3.9, 4.4, 4.5, 3.9, 3.8, 2, 
    1.9, 3.9, 1, 1.6, 1.9, 1.5, 2.5, 2.7, 1.4, 0.9, 0.8, 1.2, 1.8, 1.4, 1.9, 
    2, 1.9, 1.4, 1.1, 0.9, 1.3, 2, 0.6, 0.6, 0.2, 1.3, 0.7, 0.2, 1.3, 0.8, 
    0.6, 1, 3.2, 0.6, 3.1, 4.6, 4.5, 3, 3.4, 3.8, 4.8, 3.9, 4.4, 4.4, 2.5, 
    2.5, 3.4, 0.2, 3.6, 2.9, 2.7, 2.9, 2.4, 2.2, 1.6, 3.8, 3.9, 2.2, 1.6, 
    1.2, 2, 3, 5, 5.3, 4.3, 4.7, 4.1, 3.7, 2.2, 2.4, 6.6, 6.9, 4.3, 5, 4.3, 
    4.4, 3.9, 4.9, 5.6, 5.7, 4.7, 5.4, 6.4, 6.6, 5.4, 4.1, 1.6, 5.7, 3.1, 
    2.8, 3.7, 2, 5.1, 6.1, 3.3, 5, 5.6, 3.8, 2, 0.7, 6.7, 4.5, 4.8, 5.1, 4.5, 
    5, 5.8, 4.8, 4.1, 6.4, 8.4, 7.2, 7.2, 7.2, 7.7, 7.6, 7, 4.2, 5, 4.9, 2.6, 
    0.4, 1.4, 3, 3.2, 2.7, 1.2, 5.2, 1.3, 3, 0.8, 2, 1.4, 1.5, 1.8, 3, 2.5, 
    1.5, 1.3, 2.6, 2.6, 3.6, 3.9, 4.8, 4.8, 3, 1.6, 1.8, 2.1, 2.5, 2.7, 2.6, 
    2.4, 4.2, 4.2, 3.6, 3.9, 1.5, 1.6, 1.9, 2.8, 2, 2.6, 2.6, 3, 3.1, 3.8, 
    4.6, 4.9, 4, 4.1, 4.3, 4.5, 5.4, 6.4, 5.2, 5.8, 5.3, 5.6, 3.7, 4, 3.1, 
    3.6, 3.5, 4.7, 5.8, 6, 6.5, 5.3, 5.1, 4.7, 3.9, 4.3, 3.4, 2.1, 2.3, 2.7, 
    2.7, 2.1, 3.3, 2.4, 3.6, 4, 2.9, 2, 5.1, 5.2, 4.3, 7.1, 3.4, 7, 5.3, 3.6, 
    4.8, 5.7, 4, 5, 1.9, 4, 4, 2.1, 2.7, 0.8, 1.1, 1.4, 2, 2.6, 4, 2.8, 2, 2, 
    4.4, 3.1, 1.3, 1.5, 2.1, 2.1, 2.6, 1.7, 1.7, 4.1, 4.4, 1.3, 2.7, 0.8, 
    1.1, 1.1, 1.1, 0.9, 0.4, 1.6, 1.9, 1.6, 2.9, 3, 3.1, 4.1, 4.2, 4.2, 4.5, 
    3.7, 2.8, 2.5, 1.9, 1.4, 1.9, 1.5, 4.4, 4, 4.1, 0.6, 2.1, 0.8, 1.9, 2.7, 
    2, 2.3, 3, 3.3, 4.2, 3.6, 3.2, 2.3, 1.9, 3.9, 2.7, 2.3, 2.7, 2.4, 1, 0.8, 
    0.8, 1, 0.5, 0.5, 0.2, 0.3, 0.7, 1.2, 2, 5.7, 5.5, 6.5, 7.7, 6.6, 6.2, 
    6.5, 5.6, 1.3, 4.3, 7.8, 7.1, 9.9, 11.2, 10.3, 11.1, 10.2, 8.4, 7.8, 5.9, 
    1.5, 1.5, 0.5, 1.1, 0.9, 0.7, 1.2, 1.5, 1.5, 1.6, 2.1, 1.4, 6.5, 3.5, 
    2.9, 3.8, 2, 5.4, 7.4, 7.2, 8.2, 7.4, 6.2, 4.4, 2.8, 2.1, 2.1, 5.3, 3.9, 
    2.8, 2.4, 0.9, 6.3, 7.9, 4.7, 6.4, 7.4, 5.1, 3.9, 5.2, 6.3, 5.1, 5.4, 
    4.9, 5.5, 5, 5.8, 6.1, 4.7, 4.7, 5.2, 5.3, 5.8, 4.7, 4.6, 3.6, 4.5, 4.6, 
    3.1, 4.8, 3.7, 2.3, 1.8, 1.2, 1.1, 0, 0, 0.3, 0.4, 0.4, 0.1, 0.4, 2.8, 
    4.4, 5.7, 4.2, 5.7, 6.8, 3.8, 3.6, 6.3, 6.5, 6.8, 7, 8, 6.1, 8.1, 8, 6.5, 
    6.2, 5.3, 1.8, 1.5, 0.7, 0.7, 2.1, 3.5, 1.9, 1.5, 1.4, 1.4, 1.9, 1.8, 
    2.9, 3.7, 1.9, 1.9, 1.3, 1.3, 0.8, 1.1, 0.3, 1.2, 0.5, 1.6, 1, 1.3, 2.5, 
    0.3, 0.2, 1.3, 1.8, 1.9, 1.3, 1.1, 1.3, 2, 1.9, 1.4, 1.6, 1.7, 2.2, 3.7, 
    1.9, 2.6, 2.8, 2.1, 1.8, 1.4, 1.9, 2.6, 2.3, 1.6, 1.6, 1.5, 1.7, 1.7, 
    1.9, 2.2, 1.8, 2.6, 2, 2.8, 1.8, 1.8, 2.8, 1.4, 1.2, 1.5, 1.3, 1, 0, 1.2, 
    0.3, 0, 0.5, 0.9, 1.3, 0.5, 1.7, 1.6, 1.8, 1.2, 2, 1.7, 1.4, 1.9, 1.3, 
    1.1, 0.2, 0.3, 1.5, 1.1, 1.5, 0.9, 1, 0, 0.8, 1.6, 1.8, 2.4, 4.4, 2.9, 
    1.6, 1.6, 1.2, 1, 1.8, 1.9, 1.5, 1.4, 1.4, 1.1, 1.2, 1.6, 2.2, 0.1, 1.5, 
    1.6, 1.4, 1.3, 1.5, 1.9, 0, 0.2, 1.6, 1.9, 1, 0.6, 2.1, 2.5, 0.8, 3.1, 
    2.7, 0.7, 2.7, 2.4, 2.8, 3.3, 3.3, 2.4, 1.7, 2.2, 0.8, 1.1, 2.6, 2.4, 
    1.8, 1.7, 0.5, 1.7, 1.6, 1.9, 1.7, 1.5, 1.4, 2, 2, 2.4, 1.7, 1.4, 0.6, 1, 
    0.3, 0.8, 1, 0.5, 0.9, 0.9, 0.4, 1, 1.5, 1.7, 2.1, 1.3, 1.6, 2.5, 1.5, 
    0.8, 0.6, 1.1, 2, 2, 2.4, 2.3, 2.1, 1.8, 0.6, 1.6, 1.7, 0.7, 1.8, 1.5, 
    0.7, 0.5, 0.9, 0.5, 0.9, 1, 0.7, 0.9, 4.5, 1, 2.5, 1.4, 2.3, 1.2, 1.6, 
    2.8, 1.3, 3.1, 0.7, 2, 1.8, 0.4, 0.6, 1.8, 0.9, 0.3, 0.3, 1.1, 0.2, 0.6, 
    1.3, 2.5, 1.6, 2.1, 2.4, 0.7, 1, 1.2, 4.4, 0.9, 1.9, 3.3, 3, 2.6, 2.8, 
    1.3, 3.8, 2, 0.9, 3.8, 2.9, 4.7, 2.4, 1.2, 3.8, 1.9, 3.6, 2, 2.3, 3.1, 
    2.9, 3.3, 4.1, 4.2, 3, 4.5, 5, 5.2, 5.2, 4.6, 3.7, 2.1, 2.5, 4.4, 2.6, 
    2.3, 0.9, 1.3, 1.7, 2.4, 3.6, 4.8, 5, 4.9, 3.9, 3.1, 2.4, 2.2, 1.4, 1.5, 
    0.1, 0.8, 0.1, 0.9, 1.3, 1.3, 1, 0, 0.8, 0.5, 1.9, 1.2, 1.8, 2.4, 0.2, 
    0.2, 2.2, 2.5, 2.5, 3.2, 1.6, 1.7, 1.9, 2.7, 2.9, 2.4, 2, 3.3, 2, 2.4, 
    1.8, 1.7, 1, 0.3, 0.1, 4.1, 3.7, 4.3, 4.5, 4.3, 5, 4, 2.8, 3.5, 3.3, 3.1, 
    3.3, 2.6, 2.3, 1.9, 2, 1.5, 1.1, 1, 0.4, 1, 1.4, 3.3, 2.2, 2.1, 2.9, 2, 
    2.7, 2.7, 3.2, 3.2, 4.1, 3.8, 4, 3.7, 2.6, 3.3, 1, 0.8, 1.7, 2.2, 2.1, 
    2.6, 1, 2.6, 0.6, 1.4, 2.5, 1.3, 0.4, 2, 1.1, 0.6, 1.6, 1, 0.4, 1.3, 0.8, 
    3.2, 2.4, 1.5, 2, 3.3, 2.7, 3, 3, 3, 2, 1.4, 1.9, 2.8, 3.6, 3.1, 3.1, 
    3.2, 2.7, 2.5, 1.4, 1.6, 1.6, 1.2, 1.8, 1.8, 1.2, 1.7, 1.1, 2, 2, 3.7, 
    3.2, 2.9, 2.7, 1.7, 3, 2, 1.4, 1.1, 1.2, 1.8, 1, 0.5, 1.9, 1.4, 1.2, 4.1, 
    2.4, 3.9, 3.7, 3.6, 3.6, 1.1, 0, 0.7, 1, 1.2, 0.1, 0.7, 2, 1.8, 0.8, 2.1, 
    1.6, 1.4, 2.4, 1, 1.5, 3.9, 4.6, 4.1, 3.2, 3.7, 2.5, 4.5, 4, 3.5, 3.7, 
    4.5, 4.2, 4.7, 3.8, 3.6, 4.7, 3, 6.6, 4.9, 4.7, 4.3, 4.6, 5.7, 4.5, 4.5, 
    4.9, 4.7, 5.5, 4.2, 4.3, 4.7, 3.3, 4.6, 5.7, 3.6, 3.7, 3, 2.9, 2.2, 0.8, 
    0.9, 1.2, 1.2, 0.3, 0.9, 4, 6.8, 5.5, 6.7, 5.8, 6.3, 5.1, 5.3, 5.8, 6, 
    7.5, 7.5, 8.3, 7.4, 6.6, 5.5, 4.6, 4.2, 5.5, 5, 4.4, 3.9, 4.4, 6.3, 5.7, 
    3.2, 5, 4.9, 4, 4.8, 5.1, 4.9, 5, 4, 2.2, 3.8, 4.7, 5.1, 4.3, 3.8, 4.8, 
    3.8, 3.2, 3.4, 2.9, 2.4, 1.3, 1.4, 0.2, 1.1, 1.7, 2.3, 2.2, 1.3, 1.5, 
    5.8, 5.4, 4, 4.9, 4.2, 3.5, 5.1, 4.5, 3.2, 3.7, 4.5, 4.5, 4.6, 4.2, 5.1, 
    3.8, 2.8, 3.7, 3.6, 4.4, 3.9, 4.2, 4.1, 2.1, 4.9, 3.4, 2.9, 4.1, 3.3, 1, 
    2.1, 0.9, 1.1, 1.1, 1.4, 1.9, 1.1, 1.1, 1.2, 0.2, 1, 1.6, 1.4, 1.2, 1, 
    1.8, 2.6, 3.7, 1.9, 3.1, 2, 3.1, 3.8, 2.6, 3.5, 3.1, 2.3, 1.6, 0.5, 1.1, 
    1.5, 1.9, 1.5, 1.5, 1.2, 1.6, 2, 2.4, 3.4, 4.2, 3.8, 3.3, 3.6, 3.4, 3.6, 
    3.4, 3.1, 1.7, 1.2, 0.4, 2.2, 2.5, 0.1, 1, 0.2, 0.3, 0.5, 0.7, 0.3, 1.8, 
    2.6, 2.2, 2.8, 1.1, 2.6, 1.3, 6.5, 5.7, 5.3, 2.1, 1.4, 1.2, 0.9, 1.8, 
    1.3, 1.2, 1.4, 0.5, 1.2, 1.3, 1.3, 1.5, 2.4, 3.1, 3.6, 4.1, 3.4, 4.6, 
    4.9, 3.9, 3.6, 3.3, 3, 2.9, 3.3, 3.5, 3, 3.1, 1.5, 1.5, 1, 1.9, 2.1, 2, 
    0.5, 0.5, 1.7, 1.3, 1.5, 1.7, 2, 1.8, 2.1, 2.3, 1.6, 1.6, 1.5, 1.8, 1.3, 
    1.1, 1.1, 1.6, 1.6, 1.7, 1.3, 0.7, 1.1, 0.6, 0.9, 0.5, 1.2, 2.7, 1.2, 
    0.8, 1.6, 0.5, 1, 0.7, 0.4, 0.9, 1.3, 2.8, 1.1, 1.8, 2.1, 1, 0.8, 3, 4.1, 
    3.9, 5.3, 4.7, 3.5, 2.3, 1.4, 1.4, 0.9, 1, 0.8, 0, 0.1, 0.5, 4.5, 2.4, 
    2.7, 1.7, 1.4, 2.1, 1.6, 0.3, 1.3, 3.9, 4.5, 3.9, 3.4, 3.2, 2.4, 3.5, 
    4.5, 4.3, 4.6, 4.6, 4.6, 6, 5.7, 4.4, 4.3, 4, 4.7, 1.5, 0.6, 1.5, 2.6, 
    1.8, 1.1, 1.9, 1.3, 0.4, 0.6, 1.7, 1.5, 0.7, 1.2, 1, 0.2, 0.6, 1.2, 3.2, 
    3, 1.7, 1.5, 1.9, 2.4, 1.6, 0.6, 0.6, 1.1, 1, 1, 1, 0.8, 1.4, 0.7, 0.7, 
    1.1, 1.8, 0.7, 0.7, 0.9, 1.2, 1.3, 1.2, 0.5, 1, 1.3, 1.3, 2, 1.2, 2.5, 
    3.5, 4, 4.3, 3.1, 2.7, 2.7, 1.3, 3.2, 2.8, 1.9, 0.7, 3.6, 3.2, 2.5, 2.5, 
    2, 1.2, 5.4, 5.7, 5.5, 4.5, 6.3, 7, 4.7, 6.3, 5.2, 4.5, 3.5, 4.3, 3.2, 4, 
    3.3, 3.4, 2.1, 1.2, 1.4, 1, 0.4, 0.6, 0.7, 0.3, 0.9, 0, 0.6, 1, 1.2, 0.9, 
    1.1, 1.7, 2.1, 3.9, 1.2, 1.1, 0, 0.3, 0.6, 0.3, 0.7, 0.1, 4.7, 3.4, 5.9, 
    5.7, 3.6, 4.5, 5.4, 5.1, 5.1, 4.1, 4.6, 4.8, 5.6, 4.2, 3.6, 3.4, 4.7, 
    3.7, 4.2, 4.4, 4.4, 5, 3.7, 4, 4.9, 6.8, 6.4, 5.4, 5.5, 6.1, 5.5, 2.9, 
    4.9, 4.1, 3.8, 4.4, 3.2, 4.1, 1.5, 2.3, 0.5, 0.6, 1.6, 3, 1.7, 0.9, 0.5, 
    0.3, 0.8, 4, 3.2, 2.4, 4.3, 4.7, 3.7, 3.5, 3, 1.4, 2.4, 0.9, 2.1, 4.2, 
    2.6, 0.2, 3.1, 2.6, 1.6, 1.9, 3.3, 2.3, 0.3, 0.6, 2, 2, 0.7, 0.5, 3.5, 
    2.1, 2.1, 3.5, 2, 3.7, 3.4, 4, 3.2, 3.1, 3.4, 0.8, 1.1, 0.6, 1.1, 1.1, 
    0.9, 0.7, 1.4, 2.3, 1.1, 1.4, 1.5, 1.3, 1.4, 1.6, 2.3, 2.4, 2.3, 2.1, 
    2.1, 1.8, 1.2, 0.9, 0.3, 0, 0, 0.4, 0.2, 0.7, 0.5, 0.6, 0.4, 0.5, 0.4, 
    0.7, 0.2, 0.5, 0.5, 0.6, 0.4, 1.2, 0.9, 1.4, 1.2, 0.7, 1.9, 1.6, 1.3, 
    0.6, 1.7, 0, 0, 1.3, 1.5, 0.2, 0.9, 0.2, 0.4, 1.9, 0.8, 0.8, 1.1, 1.2, 
    1.6, 1.6, 1.5, 1.2, 1.3, 0.8, 1.5, 0.1, 0.2, 0.5, 1, 0.9, 0.1, 1.1, 1.1, 
    1.5, 4, 4.1, 5.3, 4, 3.5, 1.4, 3.8, 2.8, 5, 4, 2.5, 3.1, 2.3, 2.4, 2.6, 
    1, 0.3, 1.2, 0.5, 0.5, 0.7, 1, 0.4, 0.7, 1.4, 0.3, 1, 0.6, 1.2, 1.2, 0.8, 
    0.2, 0.7, 0.8, 1.4, 0.2, 1.2, 1.1, 0.7, 0.6, 2, 1, 0.1, 0, 0.2, 0.1, 0, 
    0.6, 0.6, 0, 0.1, 0.6, 0.6, 0.6, 0.7, 0.5, 1.4, 0.6, 0.4, 0.5, 0.7, 1.1, 
    1.9, 1.4, 1.5, 1.8, 0, 1.2, 1.4, 0.5, 1, 1, 0.9, 1.1, 1.4, 1.4, 2.2, 2, 
    1.8, 2.2, 2.2, 2.7, 2.4, 2.1, 2.8, 1, 1.7, 1.9, 1, 0.4, 1, 0.7, 0.9, 0.5, 
    1.7, 1.3, 1.3, 2.8, 2.4, 2.4, 2.2, 2, 2, 0.6, 4.2, 4, 1.2, 1.9, 3.6, 2.5, 
    3.6, 6.8, 2.5, 3.8, 4.2, 2.9, 1.1, 0.7, 3.5, 1.6, 3.9, 5.6, 1, 1.3, 1.5, 
    7.5, 4.8, 2.2, 6.7, 7.7, 7.4, 7, 1.2, 1.6, 5.3, 8.1, 3.1, 1.3, 6, 4.1, 
    3.2, 1.4, 1.1, 4.3, 1.2, 1.7, 2.1, 1.1, 2, 1.1, 3.9, 4, 1.2, 1.2, 0.6, 
    0.4, 0.6, 0.9, 2.1, 1.8, 2.3, 3.3, 2.7, 2.6, 2.7, 1.7, 0.7, 1.3, 2.1, 
    1.9, 2.1, 2, 1.9, 1.5, 2, 2.1, 1.8, 1.4, 0.3, 1.9, 1.9, 1.4, 2.6, 2.6, 
    2.2, 1, 2, 0.9, 0.9, 2.1, 0.5, 0.2, 0.4, 1.6, 1.2, 1.1, 0.8, 1.1, 1.4, 
    0.7, 2.9, 2.5, 1.8, 2.4, 3.1, 2.4, 2.4, 2.5, 0.3, 2.5, 1.6, 1.6, 0.9, 
    0.3, 0.2, 0.6, 1.6, 2.4, 1.6, 2, 2.1, 2.1, 1.9, 2.2, 1.1, 1.3, 2.4, 2.4, 
    1.4, 1, 1, 1.7, 0.9, 3.8, 3.5, 2.8, 0.4, 3, 3.3, 3, 2.9, 2.9, 3.5, 0.7, 
    0.5, 1, 4.1, 2.2, 2.4, 1.5, 1.7, 3.2, 4.3, 4.1, 4.5, 4.5, 4.7, 2.3, 1.1, 
    1.3, 2, 1.6, 2.1, 2, 0.6, 1.3, 0.1, 1.5, 1.3, 1.5, 1.3, 2.3, 2.3, 2.3, 
    1.7, 1.1, 0.5, 0.5, 0.1, 1.2, 0.9, 1.1, 0.9, 0.8, 0.5, 0, 0, 0.2, 0.5, 
    0.4, 0.5, 0.8, 0.9, 1.5, 1.6, 2.2, 1.9, 1.4, 1.9, 1.9, 1.5, 2.3, 2.5, 
    3.2, 3.3, 3.4, 3.6, 2.7, 2.6, 3, 2.8, 1.7, 1.9, 0.9, 0.5, 1.3, 1.6, 1.5, 
    1.9, 1, 3.3, 1.3, 3, 3.9, 2.9, 0.6, 1.6, 1.3, 1.5, 0.2, 1.9, 1.7, 1.8, 
    3.5, 2.4, 1.5, 1.9, 1.6, 0.7, 1, 1.3, 1.7, 1.9, 2.4, 2.5, 2.5, 1.7, 1.8, 
    1.6, 2.2, 1.7, 1.7, 0.6, 0.3, 0, 0, 0.9, 1.9, 3.3, 2.9, 3.8, 3.9, 3.2, 
    3.8, 4, 4.3, 3.5, 0.9, 1.8, 1.8, 0.6, 1, 0.7, 0.7, 0, 0.1, 0.6, 1.7, 1.1, 
    4.4, 4.3, 2.7, 5.1, 6.3, 4.1, 3, 2.1, 3.2, 2.8, 1.1, 0.9, 1.5, 2.5, 5.3, 
    4, 1, 2.7, 1.4, 0.1, 0.5, 0.1, 1.8, 1.5, 1.2, 1, 1.1, 1.4, 0.5, 0, 0.5, 
    0.3, 0.7, 0.7, 0.7, 0.6, 0.5, 0, 1.8, 0.5, 0.5, 0.2, 0.1, 0, 0.1, 0, 0, 
    0.2, 0.2, 1.3, 0, 0, 0.1, 0.3, 0.2, 0, 2.2, 3.8, 2.8, 1.1, 2, 2.4, 3, 
    2.7, 3.8, 2.5, 1.1, 0.2, 0.2, 1.9, 0.2, 0, 0.1, 0.9, 0.1, 0.3, 3, 1.4, 
    2.8, 4.2, 2.9, 2, 2.8, 2.6, 0.9, 3.7, 2.3, 2.1, 3.9, 3.9, 6.3, 3.1, 1.1, 
    0.2, 1.6, 2.2, 0.4, 0.6, 0.2, 0.6, 0.7, 0.1, 0.4, 0, 0, 0.8, 0.9, 1.4, 
    1.2, 1.5, 1.3, 3, 2.1, 1.9, 0.3, 0.5, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.5, 0.5, 0.1, 0, 0.2, 0.2, 0.6, 0.5, 0, 0.1, 1.3, 0.2, 
    3.4, 0.5, 0.4, 0.3, 1.1, 0.4, 0, 0.8, 2.2, 1.6, 3.1, 3.2, 4.2, 4.3, 3.9, 
    4.2, 3.2, 3.7, 3.8, 3.8, 1.2, 4, 4, 2.3, 3.4, 2.6, 0.4, 0, 0, 0, 1.6, 
    2.1, 1.5, 1.6, 3.5, 3.4, 4.8, 4.5, 5.2, 3.3, 3.8, 4.8, 3.2, 1.8, 1, 1.9, 
    2, 0.3, 0.3, 0.3, 1.7, 0.4, 1.3, 0.8, 0.6, 0.1, 0.4, 0.2, 0.6, 0.7, 0.4, 
    0, 0.2, 0.7, 0.3, 0.5, 1.3, 1.3, 0.4, 0.3, 1.1, 0.9, 1.4, 1.2, 0.1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.8, 0.9, 0.4, 0.7, 0.8, 0.2, 0.5, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2, 0.2, 0.4, 0.4, 0.3, 0.6, 1.1, 2.3, 3.4, 2.8, 1.9, 
    0.8, 1.9, 0.7, 1.5, 1.5, 0.3, 0.1, 0, 0, 0, 0.1, 0.3, 0.5, 0.8, 0.9, 1, 
    0.1, 0.7, 0.8, 0.5, 0.6, 0.7, 0.1, 0, 0.2, 0.2, 0, 0.2, 0, 3.2, 2.5, 0.4, 
    0.9, 0.5, 0.1, 0.4, 0, 0.4, 0.2, 0.7, 0.2, 0.8, 1, 0.8, 0.8, 0.4, 1.6, 
    2.3, 9.7, 8.2, 8.8, 7.4, 6.1, 4.7, 6.1, 5.7, 5, 5.3, 5.8, 3.6, 5.1, 4.5, 
    3.7, 4.1, 6.8, 6.4, 2.6, 6.4, 6.6, 6.7, 5.7, 2.9, 4.4, 6.5, 2.8, 2, 3.2, 
    1.1, 0.5, 0.4, 0.3, 0.2, 0.2, 0.2, 0.1, 1.5, 0.2, 0.1, 0.6, 0, 0.6, 0.1, 
    0, 0, 0.3, 0.8, 0.1, 0, 0.4, 0, 0, 0.3, 0, 0, 0, 0, 0.1, 0, 0.1, 0, 1.6, 
    0.5, 0.5, 0.4, 0.5, 0.1, 2, 0.9, 0, 0, 0, 0.1, 0.6, 0, 0, 0, 0.2, 0, 0.3, 
    0, 0, 0.1, 0, 0.4, 0.2, 0.1, 0, 0.2, 4.1, 3, 2.3, 2.7, 1.2, 1.1, 0.1, 1, 
    1.3, 0.1, 0, 0.2, 0.3, 0, 0, 0, 0, 0.1, 0.3, 0, 0, 0, 0, 0, 0.1, 0.3, 
    0.1, 2.9, 0.2, 0.7, 1.2, 1.7, 1.9, 2.8, 1.9, 2.7, 2.3, 2.3, 2.4, 2.3, 
    2.5, 2.5, 3.7, 0.9, 0, 0, 1.2, 1.2, 1.3, 1.5, 1.3, 4.1, 3.8, 1.6, 2.9, 
    2.4, 2.9, 0.5, 0.3, 0.6, 0.1, 0.7, 3.4, 3, 1.6, 1.3, 1, 0.5, 2.9, 2.3, 
    0.3, 2.1, 0.3, 1.2, 2.7, 0.1, 0.3, 1.8, 0.8, 0.1, 1.3, 0.1, 0, 0, 0, 0.3, 
    1.8, 0.7, 0.9, 0.9, 0.1, 0, 0.5, 0.4, 0.1, 1, 2.8, 3, 3.3, 2.7, 2.3, 1.8, 
    1.2, 1.1, 1.5, 2.3, 1.9, 2, 1.7, 1.5, 1, 1, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 
    0.5, 0.3, 0, 0, 0.2, 0.3, 2.6, 2, 0.3, 0, 1.6, 1.2, 0.8, 0.5, 0, 0, 0, 
    1.4, 1.5, 1.3, 0.6, 1.8, 1.8, 2, 2.1, 2.7, 3.6, 2.1, 0.7, 1.6, 0.6, 2.1, 
    0.1, 0, 0.1, 0, 0, 0, 0, 0, 0.7, 0.4, 0, 0.5, 0.6, 0.6, 0.8, 0.4, 0.4, 
    0.6, 0.8, 1.1, 0.1, 1.1, 0.1, 0, 0, 0, 0.2, 1, 1, 0, 0, 0.1, 0, 0.2, 0.7, 
    2.9, 3.4, 4.7, 3.4, 4.4, 3, 2.5, 3.5, 3.4, 3.5, 3.5, 3.7, 3.4, 4.8, 4.2, 
    3.8, 3.3, 3.6, 3.4, 3.7, 1.5, 0, 0.8, 0.5, 2.6, 6.8, 5.8, 6.4, 3.7, 4.9, 
    3.6, 2.1, 4.3, 4.8, 4.1, 3.8, 4.1, 4.2, 3.1, 3.4, 4.2, 3.8, 1.6, 0.9, 
    0.5, 0.4, 0, 0, 0, 0, 0.2, 0.2, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.3, 2.4, 3.5, 4.1, 5.3, 4, 0.2, 0.2, 0.1, 1.3, 1.6, 
    2.4, 1.9, 1.4, 1.2, 1.4, 0.6, 0, 0.4, 0, 0.1, 0, 0, 0.4, 0, 0.1, 0.4, 
    0.1, 0.1, 0, 0, 0.4, 0.5, 0.7, 0.3, 0.5, 0.6, 0, 0, 0.1, 0, 0.1, 0, 0, 
    0.1, 0, 0, 0, 0.1, 0.2, 0, 0.1, 0.3, 0.1, 0.3, 0.2, 1, 0.1, 0.1, 0.3, 0, 
    0, 0, 0.3, 0.3, 0, 0.1, 0.1, 0, 0.6, 0.4, 0, 0.1, 2, 0.1, 0, 3.5, 4.2, 2, 
    2.1, 4.6, 4.5, 5.3, 5.1, 5.1, 5.6, 3.4, 4.2, 2.3, 0.7, 0.2, 0.1, 0, 0, 
    1.2, 0, 0.9, 0, 0, 0.2, 1.1, 0.1, 0.6, 0.8, 0, 0.4, 0.8, 0.6, 0.1, 0, 0, 
    0.1, 0, 0.1, 0, 0.7, 0.5, 0.3, 0.4, 0, 0.1, 0.1, 0, 0.1, 0.6, 0.6, 0.4, 
    0.1, 1.4, 0.1, 2, 1.3, 2.1, 1.4, 0.6, 0.5, 0.8, 0.3, 0, 2.2, 1.1, 1.9, 2, 
    4.2, 4.1, 4.2, 2.5, 2.2, 2.9, 3.4, 3.2, 5.5, 5.4, 6.7, 4, 6.9, 4.7, 3, 
    5.4, 6, 3.9, 4.1, 3.6, 2.3, 3.5, 3.8, 3, 2.3, 3.6, 4.2, 3.8, 3.6, 3, 4.8, 
    3.3, 3.5, 3.4, 3.5, 2.4, 1.8, 1.8, 1.1, 4, 3.1, 0.4, 0.2, 0.6, 1.6, 1.5, 
    0.1, 0, 0.1, 1.6, 1.5, 1.5, 2, 2.4, 1.4, 0.9, 1.6, 0.7, 0.2, 0.6, 2.3, 
    2.4, 2.9, 3.1, 2.8, 1.5, 1.8, 3.4, 3.4, 3.6, 3.7, 6.2, 3.1, 6.8, 3.2, 
    5.6, 3.6, 3.8, 5.1, 5.7, 7.4, 4.7, 4.3, 4.3, 4, 2.6, 3.2, 5.5, 5, 4.3, 
    3.8, 6.6, 6, 2.7, 3.7, 1.2, 5.3, 2.2, 0.3, 0.1, 0.1, 0.6, 0.1, 0.1, 0.1, 
    0.2, 0.2, 0.1, 0.2, 0.5, 0.3, _, _, _, _, _, _, _, _, _, _, _, 5.4, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 11.1, _, _, 
    0, 0.3, 1.1, 0.7, 3.3, 0.8, 1.6, 1.3, 0.2, 0.2, 0, 1.2, 1.1, 1.4, 1.2, 
    1.4, 1.4, 0, 0.2, 0, 0.6, 0.8, 0.6, 0.8, 0.5, 0.1, 0.4, 1.9, 1.6, 1.6, 
    0.7, 0.7, 0.8, 1.4, 0.8, 0.4, 0.6, 1.2, 1.3, 1.9, 1.8, 1.1, 0.6, 1.4, 
    0.6, 0.9, 1, 2.3, 1.4, 1, 2.3, 1.6, 2.2, 2.2, 1, 1.7, 1.2, 0.8, 1, 1, 
    1.7, 1.2, 2, 1.8, 1, 0.7, 2, 1.6, 0.9, 0.7, 0.3, 0, 0, 0, 0, 0, 0, 0, 
    0.1, 0, 0, 0.6, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.4, 0, 0, 0, 
    0.6, 0.6, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0.2, 0, 0, 0.1, 0, 0, 0, 
    0, 0, 0, 0, 0.6, 1.4, 0.8, 0.3, 0.1, 0.3, 1.5, 1.1, 3.9, 3.9, 6.9, 8.1, 
    7.5, 7.4, 4.1, 0.5, 1.9, 1.3, 1.1, 0.3, 0.7, 0, 0, 1, 0.2, 0, 5.9, 7.3, 
    1.1, 2.3, 2.4, 3.2, 5.5, 5.7, 4.9, 5.1, 2.6, 1.7, 3, 1, 1.3, 0.1, 0.1, 
    0.1, 0.3, 0, 1, 0.4, 0, 0.2, 0.3, 0, 0.1, 0, 0.4, 0, 1.2, 0.1, 0, 0.1, 
    0.3, 0.3, 0, 2.3, 0.2, 0, 0, 0.4, 0.6, 0.8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1, 0, 0.9, 1, 0.4, 0.3, 0.5, 0.5, 0.2, 0, 0.4, 0.1, 0, 0.2, 0, 0, 
    0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2, 
    0.5, 1.1, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.1, 0, 0.3, 0, 0, 0, 0.1, 0.1, 0.1, 0, 0.1, 0, 0, 0.1, 0.2, 0.8, 0, 
    0.2, 1.5, 0.7, 0.1, 0.2, 0.5, 0.5, 0.4, 0.3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0.1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2, 0, 0, 0.1, 0, 0, 0, 0, 0.4, 0.4, 0, 0.1, 0.7, 0.3, 0, 0, 0.4, 0, 0, 
    0.2, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0.2, 1, 0.8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3, 1.1, 0.5, 0, 0, 0.2, 0, 0.3, 0, 0, 0, 
    0.1, 0.1, 0.1, 0.3, 0.3, 0.2, 0, 0.4, 3.6, 6, 6.3, 5.8, 8.3, 7.9, 5.9, 
    9.1, 9.2, 8.5, 9.9, 9.4, 7.6, 6.1, 4.8, 6.8, 5.2, 2.2, 1.7, 3.1, 4.8, 
    6.3, 7.2, 7.2, 5.7, 2.3, 0.9, 2.8, 2, 0.4, 0, 0.2, 1, 0.1, 0.2, 0.3, 0.2, 
    0.3, 0.1, 0.1, 0.1, 0.5, 0.1, 0.2, 0.5, 0.3, 1.2, 0.5, 0, 0, 0.6, 0, 0, 
    0, 0, 0.1, 0.1, 0, 0, 0.1, 0, 0.6, 0.1, 0, 0.1, 0, 0, 0.2, 0.1, 0.1, 0, 
    0, 0, 0.1, 0, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    0.4, 0, 0, 0, 0.7, 0.1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 3.7, _, _, _, _, _, _, 
    0.1, 0, 0.1, 0.1, 0.1, 0, 0.1, 0, 0.3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1, 0, 0, 0, 0, 0.1, 0, 0.2, 0, 0, 0, 0, 3.6, 3.2, 4.2, 3.5, 2.5, 1.2, 
    2.3, 3.5, 3.7, 1.9, 5, 6.7, 6, 6.1, 7.2, 7.1, 6.7, 5.5, 7, 8.4, 8.9, 9, 
    8.1, 10.2, 7.4, 7.2, 7.2, 5.8, 6, 5.9, 6.1, 4, 6.1, 6.3, 7.9, 5.9, 8.9, 
    9.6, 10.8, 8.6, 9.2, 10.4, 8.4, 7, 6.7, 6.6, 7.5, 6.1, 6.8, 8.2, 7.3, 
    8.6, 8.2, 7.9, 7.2, 8.5, 7.8, 5.8, 8.5, 8.5, 8.5, 8.8, 9.2, 9.1, 6.6, 
    6.2, 5.5, 6.3, 8.9, 6.5, 4.2, 4.8, 3.6, 2.5, 2.7, 5.5, 4.8, 3.8, 3.3, 
    3.4, 3.7, 3.7, 3.8, 2.5, 2.5, 2.5, 1.7, 1.6, 2.3, 3.4, 2.8, 1.8, 1.5, 
    0.1, 0.4, 3.8, 2.5, 0.6, 4.2, 3.4, 1.9, 0.2, 1.1, 0.3, 0.3, 1.9, 2.3, 
    3.3, 1.5, 1.9, 0.4, 2.3, 2.7, 1.3, 1.1, 0.9, 1.5, 0.4, 0.1, 0.1, 0.1, 
    0.7, 0.7, 0.6, 1, 2.1, 1.1, 1.5, 1.7, 1.5, 0.8, 1, 1.1, 2.3, 1.6, 0.9, 
    1.9, 1.6, 1.3, 0.7, 0.4, 0.8, 0.6, 0.1, 0, 0.1, 0.1, 0, 0, 0.4, 0.7, 0.2, 
    0.2, 0, 0.6, 0.5, 0.9, 1.1, 2.3, 0.7, 0.3, 1.5, 0.5, 0.1, 0.6, 0.3, 0, 
    0.3, 0.1, 0.4, 0.1, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0.3, 0, 0.1, 0.2, 
    0, 0.1, 0.3, 0.4, 0, 0.1, 0, 0.3, 0, 0, 0.2, 0, 0, 0.1, 0.4, 0, 0.5, 0.4, 
    0.4, 0.2, 1.6, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 2.1, 3.3, 3.3, 3, 3.4, 1, 
    3.8, 2.8, 5, 3.4, 2, 2.1, 1.4, 0, 0.5, 0, 0, 0.1, 0.3, 0.2, 0, 0, 0, 0, 
    0, 0, 0.1, 0.5, 0.1, 0.9, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0.1, 0, 0, 0.1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2, 0, 0.4, 0.6, 2, 2.1, 4.8, 3.8, 4.1, 
    4.8, 4.3, 4.2, 3.7, 3.5, 4.7, 3.5, 3.6, 3.1, 2.7, 2.4, 1.8, 1.8, 2.8, 
    1.6, 4.3, 3.6, 3.4, 1.6, 2.6, 2.4, 3.1, 4.3, 5.1, 6.9, 5.5, 4.2, 5.8, 
    3.9, 3.9, 0.2, 0.1, 0, 0.1, 4.4, 2.1, 0.3, 0.1, 0, 4.1, 1.8, 0, 0, 5, 
    4.1, 5.8, 5.6, 4.9, 5.5, 8, 10.1, 7.8, 10.4, 6.8, 6.6, 5.8, 6.5, 4.2, 
    2.7, 2.9, 3.8, 2.5, 3.2, 1.5, 1.8, 2.1, 1.5, 3.5, 2, 1.8, 6.1, 7.8, 8.7, 
    8.1, 8.5, 10.3, 10.1, 8.9, 10.9, 8.5, 10, 10.3, 10.2, 10.2, 9.4, 8.9, 
    7.6, 7.4, 7, 7.4, 5.8, 7.1, 8.3, 9.2, 8.1, 8.9, 8.4, 9.2, 9.3, 8.9, 10, 
    8.5, 9.1, 8.7, 6.8, 7.9, 6.5, 7.3, 5, 7.8, 7.4, 7.3, 8.5, 6.3, 6.3, 4.7, 
    4.2, 3.9, 5.3, 4.1, 2.9, 3.8, 3.5, 2.4, 0.7, 1.1, 1.8, 0.8, 0.1, 0.9, 
    0.2, 0.2, 0.1, 0.1, 0.1, 0.1, 0, 0, 0, 0, 0, 0.2, 0, 0.2, 0.1, 0.1, 0, 0, 
    0.1, 0, 0, 0.1, 0.1, 0, 0, 0, 0.1, 0, 0.9, 0.2, 0, 0.1, 0, 0, 0, 0, 0, 
    0.2, 0, 0.9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0.2, 0.1, 0, 0.1, 0.5, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.7, 0.1, 0, 0, 0.1, 0.3, 0.1, 0.2, 0, 0, 0.3, 
    0.2, 0, 0.1, 0.8, 3.8, 4.2, 4.4, 2.7, 0.2, 0.2, 0, 0, 0, 0, 3.6, 4, 3.6, 
    3.3, 3.2, 3, 4.5, 1.5, 2.7, 5.4, 5.3, 3.3, 1.5, 4.7, 2.2, 1.2, 3.1, 0.2, 
    0.1, 1.2, 0, 0, 0.3, 1.1, 0.6, 0.1, 0.2, 0.9, 1.6, 0.6, 1, 0.8, 0.5, 0.1, 
    0.8, 0.8, 0.5, 0, 0.1, 1, 0.1, 0.6, 0.2, 0.3, 0, 0, 0.1, 0.1, 0, 0, 0.2, 
    0.2, 0.2, 0, 0, 0, 0, 0, 0, 0, 0.5, 0.4, 0, 0.4, 0.1, 0.1, 0.3, 0.4, 0.3, 
    0.1, 0.2, 0.3, 0.6, 1.4, 0.2, 0.1, 0, 0, 0.1, 0, 0.4, 0.3, 0, 0, 0, 0.5, 
    0.1, 0.1, 0.1, 0.2, 0.1, 0.3, 4.4, 3.8, 5.4, 3.9, 7.1, 7.1, 9.3, 8.5, 
    7.8, 8.2, 7.9, 7.7, 7.4, 6, 5.4, 3.2, 0.8, 1, 4.2, 0, 0, 0, 0.1, 0, 0.1, 
    0, 0.6, 0.1, 0.5, 0.4, 0.4, 0, 0, 0, 0, 0, 0.1, 0, 0.1, 0, 0.1, 0.3, 0.2, 
    0.3, 0, 0, 0.1, 0.1, 0.6, 0.5, 0.1, 0, 0, 0, 0.7, 0.3, 0.8, 0, 0, 0.8, 
    1.1, 2, 2.2, 4.7, 4.8, 6.9, 6.1, 5.9, 6.5, 6, 6.1, 2.3, 2, 2.4, 2.5, 3.8, 
    3.6, 4.9, 3.4, 4.6, 1.6, 1.9, 2.3, 1.6, 1.3, 2.9, 8, 5.6, 3.6, 4.1, 6.7, 
    5.1, 4.2, 7.7, 4.2, 5.7, 8.3, 6.8, 5, 3.9, 6.2, 5.3, 4.4, 3.8, 3.3, 1.6, 
    6.5, 3.1, 1.4, 1.9, 2.6, 6.1, 2.1, 2, 0.2, 0.6, 1.7, 1.3, 0.9, 0.8, 0.8, 
    1, 2, 3.5, 0.9, 1.3, 0.8, 0, 1.5, 0.5, 0.7, 0, 0.4, 0.2, 0.2, 0.4, 1, 
    1.1, 1.2, 1, 0, 0.1, 0, 0, 0, 0.1, 0.2, 0.9, 0.2, 0.1, 0.7, 0.1, 0.1, 
    0.1, 0.7, 0.4, 0.1, 0, 0, 0, 0.1, 0.2, 0.2, 0.2, 0.3, 0.1, 0, 0.2, 0.5, 
    0, 0, 0, 0, 0.1, 0.2, 0, 0, 0.2, 0.5, 0.7, 0.5, 2.2, 4.8, 5.1, 4.2, 4.2, 
    6.4, 6.4, 6.4, 5.7, 4.2, 6.6, 5.4, 5.2, 5, 5.8, 3.3, 1.8, 4.6, 4.1, 4.4, 
    4.4, 1.8, 1.2, 1.4, 0.3, 0, 0.2, 0.2, 0.3, 1.7, 0.8, 0, 0.8, 0.1, 0.5, 
    0.1, 1.6, 6.2, 6.3, 4.4, 5.8, 4.5, 0.7, 0.2, 1.6, 2.5, 0.3, 0.7, 0.5, 
    0.9, 0.7, 1.7, 0.1, 0.9, 0, 0, 0, 0.1, 0, 0.1, 0.2, 0.1, 0.1, 0.7, 0.3, 
    0.1, 0, 0, 0.3, 0, 0.4, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5, 0.3, 
    0.1, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0.2, 0.1, 0.1, 
    0, 0.2, 0.6, 4.7, 6.4, 8.5, 8.2, 7.4, 5.4, 1.6, 3.1, 3.4, 3.3, 2.6, 2.7, 
    3.2, 2.1, 1.1, 1.4, 1.4, 0, 0.7, 0.2, 0.8, 0.1, 0, 0.1, 0, 0, 0.1, 0, 
    0.2, 1.6, 5.2, 3.8, 5, 2, 2.9, 12.7, 6.7, 2.3, 0.9, 0.3, 0.1, 0.2, 0.1, 
    0.5, 6.5, 6.7, 6.4, 8.5, 7.6, 3.6, 4.4, 6.4, 6, 3.8, 3.2, 5.2, 4, 4, 4, 
    4.4, 2.3, 3.9, 5.2, 4.2, 5.2, 7.3, 5.1, 5.3, 3.5, 1.9, 1.6, 4.8, 5.5, 
    3.2, 5.4, 1.7, 5, 6.4, 4.9, 6, 7.2, 10.9, 9.3, 8.7, 8.9, 7.9, 5.5, 7.4, 
    8, 7.4, 8.2, 8.1, 6.4, 7.1, 6.9, 6, 6.4, 5.8, 6.3, 6.3, 7.8, 3.7, 4.1, 
    5.8, 8.1, 8, 6.7, 5, 5.7, 6.5, 2.8, 3.2, 4.2, 3.7, 3.9, 2.2, 5.1, 5.5, 
    6.2, 5.3, 4.9, 4.6, 4.7, 4.2, 4.3, 4, 3.4, 3.2, 1.3, 3.3, 5.2, 4, 2.3, 
    1.6, 3.6, 1.8, 5, 5.5, 4.3, 3.9, 4.9, 5.9, 3.3, 2.6, 2.4, 4, 5.2, 2.7, 
    4.3, 2.5, 4.2, 3.5, 3.7, 5.2, 5.2, 4.7, 4.8, 4.4, 7, 6.4, 6.8, 6.8, 6.8, 
    6.8, 6.9, 6.6, 5.6, 4.8, 5.1, 4.8, 4.3, 3.6, 4, 2.3, 1.6, 0.8, 0, 0.4, 
    0.4, 0.1, 0.5, 0.4, 0.6, 0.4, 0.1, 0.6, 5, 4.8, 3.4, 0, 0, 0.2, 0, 0.1, 
    0, 0, 0, 0.1, 0.2, 0.4, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 1.9, 0, 0, 
    0, 0, 0, 0.3, 2.6, 4.4, 6.6, 7.4, 7.4, 7.9, 7.8, 9.2, 7.3, 7.8, 7, 8.1, 
    7.3, 6.6, 4.2, 7.8, 8.5, 7.8, 7.5, 7.1, 6.9, 7.6, 6.9, 7.3, 1.5, 3.6, 
    5.6, 4.8, 5.7, 7.1, 6.1, 7, 4.5, 4.8, 1.3, 1.2, 2.8, 2.1, 2.9, 5.4, 5.6, 
    6, 4.1, 1.6, 5.3, 1.9, 2, 0.4, 2.8, 5.5, 2.9, 0.1, 0.3, 1.2, 0.6, 0, 0.5, 
    0.1, 2.9, 2, 2.9, 6.2, 2.7, 4.5, 5.8, 4.9, 4.7, 4.3, 4.6, 3.3, 0.9, 0, 0, 
    0.1, 0.1, 1.1, 0.4, 0, 0.2, 0, 0.3, 0.6, 2.3, 0.2, 0.2, 0.1, 2.2, 5.3, 
    3.3, 4.3, 5.2, 3.2, 2.2, 0.3, 0.6, 1.8, 0.7, 0.8, 0.3, 0.8, 1.2, 0, 0, 0, 
    0.2, 0.4, 2, 2.3, 1.6, 0.5, 0, 0.1, 0, 0.4, 0.7, 1.9, 3.2, 1.8, 2.3, 2.9, 
    1.9, 2.3, 4.9, 2.4, 4, 4.3, 4.1, 2.5, 2.4, 0.4, 3.5, 3, 2, 0.4, 0.1, 0.1, 
    0.3, 0.6, 0.6, 1, 0.1, 0.1, 0, 0.1, 0.2, 0.2, 0, 0, 0.2, 0.1, 0, 0.1, 0, 
    0, 0.1, 0.1, 1.1, 1.6, 0, 0.1, 0.7, 0.8, 0.1, 0.9, 3.9, 6.5, 5.7, 5.2, 
    4.7, 3.5, 3.6, 4.1, 3.3, 3, 3.9, 2.4, 3.2, 4.7, 4.7, 5, 2.8, 3.1, 1.8, 
    0.6, 0.1, 0.1, 0.8, 0, 0, 1.6, 0.3, 0.3, 0.7, 0, 0, 0, 0, 0.1, 0.2, 0.3, 
    1.4, 0, 0.6, 0.1, 1, 1.5, 1.8, 1, 0.2, 0, 0, 0, 0, 0, 0, 0.2, 0, 0, 0, 
    2.5, 5.2, 5.2, 3.2, 3.6, 3.9, 3.9, 6.1, 7.2, 6.3, 6.2, 3.2, 3.1, 6.1, 
    6.9, 2.7, 4.4, 2.1, 0.7, 0, 0.4, 0.2, 0.2, 0, 0.3, 0.7, 1.9, 2, 1.1, 1.7, 
    2.3, 0, 0, 0.6, 0.2, 3.1, 0, 0.3, 0.1, 0.1, 0.1, 0.9, 1.6, 0, 0.6, 0, 
    0.4, 1, 0.4, 0.6, 0.1, 0.2, 0.4, 1.3, 1.2, 0.4, 1, 0.5, 0.3, 0.1, 0, 0.2, 
    0.4, 0.4, 0.7, 0.3, 0, 0.7, 0.7, 2.2, 0, 0, 0.1, 0.6, 2, 0.1, 0, 0, 0, 0, 
    0.5, 0, 0.4, 0.5, 0.7, 5.9, 10.5, 8.7, 7.4, 7.7, 4.6, 3.7, 3, 3.7, 4.2, 
    4.6, 3.9, 4.5, 3.2, 1.6, 2.7, 3.7, 2.4, 3.1, 3.1, 4.1, 3, 2.5, 2.9, 2.8, 
    2.7, 2.6, 3.4, 1.6, 0.4, 0, 0, 0, 0, 0.3, 0, 1.8, 0.5, 2.3, 2.2, 2.7, 
    1.9, 0.7, 0, 0, 0, 0, 0, 1.4, 3.2, 4.3, 3.2, 4.4, 3.7, 3.2, 4.7, 4.8, 
    3.4, 5.3, 2.6, 3.5, 4, 3.9, 3.8, 3.2, 0.8, 0, 0.2, 0.2, 0.1, 0.1, 0, 0, 
    0.1, 0, 0, 4.8, 5.7, 5.9, 5.7, 6.5, 6.7, 5.6, 6.3, 0.1, 0.4, 7.8, 6.2, 
    9.7, 9.8, 9.3, 10.2, 10.1, 7.9, 10.5, 9.2, 9.5, 9.3, 8.4, 8.9, 8.7, 9.8, 
    7.1, 6.9, 4.1, 4.8, 3.4, 0.3, 5.2, 2.4, 6.7, 4, 2.6, 0, 0.2, 1.9, 0.1, 
    0.9, 0.1, 1.1, 0.6, 0.9, 1.1, 0.9, 0.5, 1.6, 2.2, 2.6, 0.1, 0.7, 0.4, 
    0.6, 0.2, 0.3, 2.5, 0.1, 2.5, 2.1, 2, 0, 0, 0, 2.9, 1.1, 3.4, 6.6, 7.2, 
    6.5, 7.4, 7.5, 7.7, 8.3, 7.4, 7.6, 7.1, 8.5, 7.5, 7.3, 7.3, 8.1, 7.3, 
    7.2, 4.7, 7, 8.2, 9.1, 9.2, 8.4, 8.2, 8.5, 8.2, 7.5, 7.4, 7.4, 7.8, 7.5, 
    8.5, 10, 9.6, 9.8, 8.9, 8.3, 7.6, 8.3, 7.2, 6.8, 7.9, 6.4, 6.5, 5.7, 6, 
    4.8, 4.6, 2.5, 0.4, 0, 1.4, 1.4, 1.6, 1.6, 2.7, 2.9, 1.3, 0.1, 0, 0.4, 
    0.1, 0.2, 0, 0, 0.8, 1, 0.3, 1, 1.8, 1.1, 0.6, 0, 0, 0, 0.4, 0.2, 0.9, 
    4.7, 2.7, 2.1, 1.6, 1, 0.6, 0.5, 1.1, 0.9, 1.2, 0.7, 0.7, 0.5, 0, 0, 0, 
    0, 1.2, 0, 0.5, 1.5, 2.4, 0.7, 0.1, 1, 1.6, 0.4, 2.2, 2.7, 4.7, 3.6, 3.1, 
    2.1, 1.3, 3.4, 3.9, 3.1, 0, 0.9, 0.5, 1, 1.1, 0.2, 0.6, 1.1, 2.4, 4, 4, 
    4, 3.5, 1.7, 2.6, 2.3, 0, 0, 0, 0, 0.5, 0, 0.2, 0.8, 1.8, 0.1, 0.5, 0, 
    1.7, 0.1, 0.9, 1.3, 1.3, 1.4, 0.8, 0.1, 1.3, 1.3, 3.1, 1.1, 0.4, 0.6, 0, 
    0.7, 0.2, 0.2, 0, 0, 0, 0.3, 1, 0.7, 0.7, 0, 0.8, 0.6, 0.2, 0.3, 0.2, 0, 
    0.8, 3.9, 2.2, 1.2, 1.1, 2.2, 1.8, 0.3, 2.8, 1.4, 1.4, 1.4, 2.3, 1.7, 
    1.9, 0.7, 4.4, 4, 3.3, 2.2, 1.1, 0.1, 1, 1.8, 1.6, 0.2, 0.6, 0.2, 0, 0, 
    0.6, 0.9, 2.6, 1.8, 1, 0.7, 0.4, 0, 0, 0, 0, 0, 0, 0.2, 0.1, 0.4, 0, 0.2, 
    0.2, 0.4, 0.1, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 
    0, 0, 0.3, 0, 0, 0, 0, 0, 0, 0.2, 0, 0, _, _, 0.9, 1.4, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 3.5, 5.2, 4.8, 4.8, 5.3, 2.9, 
    4.2, 5.6, 5.6, 5.8, 6, 3.1, 3.1, 3.3, 5.9, 7.5, 9.7, 10.1, 10.5, 11.8, 
    10.5, 11.5, 12.7, 12.2, 12.1, 12.7, 11.6, 11.5, 11, 11.8, 11.4, 9.5, 8.6, 
    8.6, 11.4, 11.5, 11.2, 9.9, 7.6, 5.8, 7.8, 6.5, 7.3, 7.6, 8.1, 7.3, 5.7, 
    10.2, 8.5, 8, 10.1, 10.1, 9, 8.6, 8, 7, 7.9, 7.6, 7.4, 7.7, 6.8, 7.5, 
    7.3, 6.6, 7.1, 5.9, 5.6, 5.1, 5, 1.1, 0.9, 3.1, 2.4, 0.2, 0, 0.2, 0.1, 
    0.7, 0.5, 1.7, 1.1, 0.2, 0.5, 1.6, 1.6, 0.7, 2.6, 3.1, 0.8, 0.2, 0, 1.7, 
    1.2, 3, 2.4, 2.4, 1.1, 1.8, 0, 0.5, 0, 0, 0, 2.3, 0, 0.1, 0, 6.2, 6.9, 
    8.6, 12.3, 11, 10.1, 10.2, 13.8, 11.9, 15.5, 16.1, 12.2, 12.2, 11.2, 
    11.1, 11.5, 12.1, 9.6, 11.3, 9.1, 10.1, 7.8, 8.1, 9, 7.8, 2.9, 3.3, 3.6, 
    2.4, 3, 3.7, 2.5, 2.2, 1.4, 2.4, 5.5, 2.6, 1.6, 4.3, 1, 2.9, 2.1, 0.9, 
    1.6, 1.3, 3.5, 1.6, 1, 0.4, 0.4, 0.3, 2.3, 1.6, 2, 0.7, 0.7, 1.5, 0.5, 
    0.9, 0.4, 0.1, 0.2, 0.3, 0.6, 0.2, 1.3, 0.8, 1, 3.3, 2.7, 0.9, 1, 0.7, 
    1.1, 1.1, 0.7, 2.1, 3.7, 3.2, 4.2, 4.9, 5.6, 3.8, 3.9, 4.5, 3.4, 2.6, 
    1.3, 3.4, 0.3, 2.5, 1, 2.7, 0, 0.1, 0.3, 0.4, 0.6, 2.6, 0.5, 1.1, 0.2, 
    0.9, 1.7, 0, 0.1, 0.5, 0.5, 0.3, 0.2, 0.1, 0.5, 0.1, 0, 0, 0.2, 0.2, 0.2, 
    0.2, 1.5, 0, 0.1, 0.8, 0, 0, 0, 0, 0, 0, 0.2, 0.3, 0.4, 0, 0.4, 0.1, 0.1, 
    0, 0, 0, 0, 0.3, 0.5, 0, 0.5, 0, 0, 0, 0.2, 0.3, 0.1, 0.2, 0, 0, 0, 0.2, 
    0.5, 0.3, 0, 0.1, 0, 0.2, 0, 0, 1.3, 0, 0.1, 1, 2.5, 0.1, 3.2, 0.7, 0.1, 
    0.2, 0, 0.2, 0.6, 0.7, 0.3, 0, 1, 3.2, 2.9, 1, 0.4, 0.1, 0.3, 0, 0.5, 
    0.1, 0.5, 1.4, 3, 3, 0.6, 0.3, 0.2, 0.5, 1.7, 0.3, 1.1, 3.1, 5.5, 5.6, 
    5.9, 5.7, 6.9, 8, 7.4, 6.9, 7.4, 8.1, 7.5, 6.9, 6.6, 8, 6.8, 7.3, 7.8, 
    3.4, 5, 3.5, 1, 1.1, 1.6, 0.7, 0.5, 0.4, 0.6, 0.4, 0, 0.5, 0, 0.1, 0, 
    0.2, 0, 0.1, 0, 0.3, 0, 1.1, 0.5, 0.1, 0.6, 1.5, 0.2, 0.1, 0.3, 0.1, 1, 
    0, 0.6, 0.3, 0, 0, 0.1, 0.1, 0.4, 0, 0, 0.1, 0.4, 0, 0, 0, 0, 0, 0, 0, 
    0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3, 0, 0, 0, 0.2, 0.3, 0.1, 0.3, 
    0, 0.1, 0, 0, 0.2, 0.1, 0, 0.2, 0.3, 0.3, 0.1, 0.4, 0.2, 0, 0.6, 0.6, 
    0.6, 1.2, 0, 0.5, 0, 0.9, 0.3, 0, 0, 0, 0.3, 0, 0, 0, 0, 0, 0.4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.2, 
    0.9, 0, 0.1, 0.3, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 
    0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 
    0.1, 0.3, 0, 0.1, 0, 0.2, 0.1, 0.1, 0.1, 0.1, 0.2, 0, 0, 0.3, 0.1, 0, 
    0.1, 0.3, 0.4, 0.7, 0.6, 0.9, 0.5, 1.5, 0.3, 0.2, 0.2, 0, 0.2, 0, 0.3, 
    0.4, 0.3, 0.2, 0.1, 0.1, 2.5, 1.2, 0.1, 0, 0.9, 2.4, 0, 0.1, 0.5, 0.1, 
    0.5, 0.1, 0.1, 0, 0.4, 0.7, 0.3, 0.9, 0.7, 0.7, 0.2, 4.9, 6.2, 5.5, 5.5, 
    5.5, 5.8, 5.8, 7.7, 7.3, 6.8, 7, 7.9, 7.3, 8, 7.6, 7.5, 7.9, 6.6, 6.7, 
    6.5, 5.7, 5.5, 4.5, 4, 4.2, 4.1, 3.3, 0.3, 0.4, 0.3, 4.4, 4.7, 5.1, 4.5, 
    4.7, 4.8, 4.8, 5.1, 5.7, 5.7, 5.8, 5.2, 5.1, 5.2, 5.5, 5.5, 6.6, 5.7, 
    5.1, 3.8, 1.8, 0, 0.3, 0.8, 0.4, 0.5, 0.2, 1.2, 1, 0.5, 0.6, 1.8, 0.6, 0, 
    0.5, 0.5, 0.1, 0.2, 0, 2.2, 0.1, 3, 3.9, 4.3, 4.1, 4.2, 3.3, 3.4, 3, 3.8, 
    3.9, 3.5, 2.4, 0.3, 0.3, 0.6, 0, 0.1, 1, 0.2, 0.5, 0.2, 0.4, 0.1, 0.1, 0, 
    0.2, 0.1, 0.7, 0.1, 0.3, 0.7, 0, 0, 0.1, 0.5, 0.1, 0.8, 0.5, 1.3, 0.2, 
    0.6, 0, 0.2, 0.5, 1.9, 2.9, 0.2, 1.3, 1.5, 2.4, 2.8, 2.7, 2.3, 1.5, 1.6, 
    0, 0, 0.4, 0.9, 0.8, 0.7, 0.8, 0.1, 0.7, 0.3, 0.7, 0.6, 0.1, 0.1, 0.2, 
    0.9, 0.3, 0, 0, 0.6, 0.5, 0.5, 0.7, 0.2, 0.4, 0, 0, 0, 0.1, 0.4, 0.2, 
    0.6, 1.1, 0.1, 1.1, 0.9, 0.3, 0.9, 0.5, 0.5, 0, 0.1, 0.7, 0.3, 0.2, 0, 
    0.2, 0, 0, 0.9, 0.1, 0.1, 0, 0.1, 0, 0, 0, 0.6, 0, 0, 0, 0.1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1, 0.2, 0.1, 0.1, 0, 0, 0.1, 0.1, 0.1, 0, 0.5, 0.4, 0.5, 
    0.1, 1.2, 0.7, 1.2, 0.7, 0.7, 1.2, 0.2, 3.2, 3.4, 3.5, 3.6, 3.6, 4, 4.5, 
    4.3, 3.2, 4.5, 3.9, 5.2, 4.7, 3.7, 3.9, 3.8, 3.9, 4.2, 4.7, 3.4, 3, 4.1, 
    2.9, 3, 3.2, 3, 3.3, 2.6, 3.1, 3.9, 2.7, 5.1, 3.7, 2.3, 1.2, 0.5, 4.3, 
    1.5, 1.4, 1.4, 4.9, 4.3, 0.7, 1, 1.2, 0.6, 1.2, 1.3, 0.2, 0.4, 0.6, 0.5, 
    0.5, 4.2, 2.2, 0.6, 3.1, 3.3, 0.5, 0, 0.5, 0.4, 0.2, 0, 0.2, 1.3, 0.2, 
    0.1, 0, 0.1, 0.4, 0.3, 0.2, 0.4, 0.1, 0.5, 0.1, 0.2, 3, 0.6, 0.8, 1.5, 
    0.5, 0.2, 1.3, 0.7, 1, 0.2, 0.1, 0.3, 1.4, 0.3, 0.3, 0, 0, 0.5, 0, 0.1, 
    0, 0, 0, 0.4, 0.2, 0.1, 0.2, 0.2, 0.3, 0.8, 0.2, 0.1, 0.4, 1, 2.5, 0.6, 
    2.1, 2, 1.6, 0.2, 1.8, 6.1, 0.3, 4.1, 3.8, 3.6, 1.2, 1.9, 0.1, 5.2, 5.5, 
    1.4, 0.2, 5.3, 5.5, 3.9, 4.9, 4.2, 2.1, 0.9, 1.2, 0.3, 0.3, 0.7, 0.1, 
    0.3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 
    0.6, 0.5, 0, 0.1, 0, 0, 0.1, 0, 0, 0.1, 0.1, 0.2, 0, 0.2, 0.2, 0, 0, 0.2, 
    0, 0, 0.5, 0, 0, 0, 0, 0, 0.3, 0, 0, 0.1, 0, 0.1, 1.5, 0, 0, 0, 0.1, 1.2, 
    0, 0, 0.2, 0.4, 0.7, 0, 0, 0.1, 0, 0.2, 0.1, 4.7, 4.3, 2.3, 0.9, 0.8, 
    0.6, 1.9, 2.9, 5.9, 6.2, 6.8, 5.7, 5.8, 7.8, 7.9, 6.2, 5.6, 2.8, 7.7, 
    0.5, 4.3, 2, 1.7, 3.9, 2.4, 0.2, 2.1, 2.7, 2.5, 3.1, 2.4, 3.6, 2.1, 2.6, 
    2.6, 4.1, 4, 4.8, 5, 4, 3.6, 1.6, 2.1, 1.8, 1.2, 0.8, 1.4, 0.7, 0.3, 0.6, 
    1.6, 2, 0.2, 2.9, 0.4, 1.5, 1.9, 0.6, 1.1, 1.3, 0, 0.3, 0, 1, 0.1, 0, 
    0.3, 1, 0.6, 0.2, 0.7, 0.3, 1.1, 0.3, 0.3, 0, 0.6, 0.2, 0.6, 1, 0.3, 0.2, 
    0, 0, 0.7, 0.2, 0.3, 0.2, 0.1, 0, 0, 0, 0.5, 0.6, 0.1, 0.8, 0.2, 0.3, 
    0.6, 0.5, 0, 0, 0, 0.2, 0.1, 0, 0.1, 0.1, 0, 0, 0.3, 0.1, 0.8, 0.5, 0.2, 
    0.4, 0.5, 0.6, 1.8, 0, 0.1, 0.6, 0, 0.1, 0.4, 0, 0.3, 0.2, 0.3, 0, 0, 
    0.5, 0, 0.8, 0, 0.3, 0.3, 0.2, 0, 0.4, 0, 0, 0, 0, 4.5, 4.8, 6.2, 6, 7.2, 
    7.5, 7, 6.3, 7.4, 7.2, 5.6, 4.7, 9.4, 6.5, 5.3, 5.1, 4, 0.5, 0.5, 0, 1.6, 
    0.2, 0.3, 0.2, 0, 0, 0, 0, 3, 3, 3.5, 0.4, 1.1, 0.6, 1, 2.3, 3.7, 4.5, 
    3.8, 0.1, 0, 0, 0.1, 0.1, 0.3, 0.6, 0.1, 0.3, 0.4, 0.2, 0.4, 0.5, 0.3, 1, 
    0.1, 0, 0.1, 0.1, 3.4, 3.2, 5.2, 6.3, 6.1, 6, 5.8, 5.6, 6.1, 6.5, 10.9, 
    10.6, 10.8, 12.8, 12.2, 11, 3.4, 7, 9.9, 6.2, 8.6, 4.5, 6, 5, 8.5, 3.2, 
    1.2, 1.4, 0.1, 0.4, 0.7, 0.1, 0.2, 0.3, 0, 0.1, 0.7, 0.4, 0.5, 0.4, 0, 0, 
    0, 0.1, 0, 0.1, 0, 0, 0, 1, 0.9, 1.1, 0.9, 0, 0.2, 0.5, 0.8, 0, 0.1, 0, 
    0.2, 1, 0, 0.5, 0.6, 0, 0.1, 0, 0, 0, 0, 0, 0.8, 2.6, 1.6, 0.7, 0.8, 2.9, 
    1.1, 1.7, 0.6, 0.5, 0.5, 0.3, 0.7, 1.7, 2.1, 4.9, 4.2, 3.2, 3.3, 5.4, 
    7.7, 1.9, 8.7, 10.7, 3.2, 2.5, 5.2, 11.2, 9.8, 12.1, 8.6, 6, 5, 2.6, 8.6, 
    2.7, 5.9, 2, 1.2, 3.1, 4.2, 2, 1.7, 0.5, 1.1, 0.5, 1.2, 0.8, 2.7, 1.7, 
    0.6, 0.4, 1.8, 0.3, 1.3, 0.4, 1.2, 0.1, 1.4, 5.5, 2.9, 1.6, 1.7, 1.1, 
    0.1, 0.6, 0, 0, 0.1, 0.3, 2.4, 2.1, 3.5, 3.6, 4.1, 1.3, 1.8, 0.3, 0.4, 
    0.4, 1.2, 1.6, 1.6, 0.9, 0.1, 1.1, 1.6, 3, 1.1, 0.3, 0.2, 0.2, 3, 1.7, 
    2.7, 6.3, 9.7, 5.7, 6.7, 8.5, 6.6, 2.7, 4.3, 4, 4, 9.5, 2, 2.1, 2.8, 1.2, 
    0.8, 2.1, 1.6, 2.6, 2.6, 4.2, 2.4, 0.2, 2.9, 1, 1.1, 3.3, 4.7, 1.8, 2.5, 
    3.9, 1.5, 2.5, 2.3, 0.8, 0.4, 0.7, 1.4, 0.5, 0, 0.1, 0, 0.4, 0.2, 0.4, 
    0.2, 0, 0.3, 0.2, 1.2, 0.5, 1.2, 0.7, 2.8, 2, 1.3, 2.5, 0.2, 1.9, 0.8, 
    1.5, 3.3, 0.7, 3.5, 3.6, 2.1, 2.3, 1.2, 1.3, 1.5, 1.1, 0.5, 1.9, 2.6, 
    2.1, 2.8, 4.7, 2.2, 1.9, 4, 2.5, 4.6, 5.1, 3.3, 3.9, 3.9, 2.8, 0.5, 0.2, 
    0.1, 0.4, 1.6, 2.9, 0.1, 4.5, 6.8, 0.5, 0, 0.8, 0.6, 0, 2.2, 0, 1, 0, 
    1.4, 0.4, 0.4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2, 0, 0, 0.8, 
    0.5, 0.7, 0.5, 0, 0.1, 0.4, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0.2, 
    0.1, 0.2, 0.1, 0, 0.5, 1.2, 0.9, 0.7, 2.3, 0, 0.7, 0.1, 0.4, 1.4, 0.1, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0.2, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.7, 0, 0.4, 0.6, 0.7, 0.2, 0.2, 0.1, 0.1, 0, 0.1, 
    0.1, 0, 0.1, 0, 0, 0, 0, 0, 0.2, 1.1, 0.2, 0, 0.1, 0, 0, 0, 0, 0, 0.1, 0, 
    0, 0, 0, 0, 0, 5.4, 5.3, 4.7, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9.4, 0, 0, 0.1, 0.3, 0, 0, 0, 0, 0.7, 0.9, 0.2, 0.3, 
    0.2, 1.4, 0.2, 0.1, 0.5, 0.1, 0, 0, 0, 0, 0.1, 0, 0.1, 0, 0.3, 0, 0, 0, 
    0.4, 0, 0.5, 0, 0.1, 0, 0, 0, 0.2, 0, 0, 0, 0, 0.8, 0.5, 0, 0.1, 2, 0, 0, 
    0.5, 0.1, 0.1, 0.2, 0, 0.3, 0, 0, 0, 0, 1.2, 0.2, 0.1, 0.7, 0.2, 0.6, 
    0.1, 3, 0.9, 1.6, 2.4, 2, 0.4, 11.3, 10.7, 11.4, 13.2, 13.5, 8.4, 6.1, 
    4.3, 3.7, 5.3, 2, 3.1, 3.1, 3.6, 3.3, 2.5, 2.2, 1.4, 0.2, 1.4, 1.8, 2.4, 
    2.1, 1.7, 0, 0.6, 0, 0.1, 0.5, 3.7, 0.9, 6.1, 7.5, 7.6, 9, 8.6, 9.1, 9.8, 
    8.9, 10.6, 9.3, 2.1, 2.4, 3.4, 2.1, 3.1, 3.1, 3.1, 3.5, 3.5, 2.8, 3.6, 
    3.7, 3.2, 3, 2.8, 2.2, 2.1, 0, 0, 0, 0.1, 0.2, 0, 0.3, 0.1, 0, 0.2, 0.2, 
    0.4, 0.6, 0, 0, 0, 0, 0.4, 0.1, 0.1, 0, 0, 0, 1.1, 0.5, 0.4, 0.9, 0.4, 
    0.4, 2, 0.1, 1.1, 0.4, 0.1, 0.2, 0, 0, 0.2, 0.5, 0.1, 0, 0.1, 0, 0.8, 
    0.2, 0.6, 0.1, 0.1, 0.9, 0.4, 0.3, 0.2, 0.4, 1.5, 1.7, 1.7, 0.5, 1.4, 
    0.4, 3, 6.8, 6.8, 6.7, 6.7, 1.9, 1.2, 1, 0.9, 0, 0.8, 0.5, 0.1, 0.4, 0.6, 
    0.4, 0.5, 3, 2.7, 1.6, 1.8, 1.1, 2.3, 4.6, 5, 3.5, 1.5, 5.4, 0.9, 0.5, 
    0.1, 0.1, 0.2, 0.6, 0.9, 0.2, 0.2, 1.9, 3.3, 1.4, 3.7, 2.2, 6.1, 6.9, 
    3.6, 2.8, 4, 1.4, 3.1, 3, 5.5, 1.3, 3, 0.5, 1.3, 1.7, 1.8, 2.6, 2.5, 0.8, 
    1.4, 0.1, 0.1, 0, 0, 0.4, 0.7, 0.6, 0.6, 0, 0, 1.3, 0.4, 2.8, 3.8, 0.2, 
    0.1, 0.1, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0.1, 0.3, 0.3, 
    0.7, 1, 1.1, 3, 2.9, 2.3, 3.9, 4.1, 0.5, 4.2, 3.5, 2.5, 0.2, 0.3, 0.1, 
    4.7, 4.4, 3.1, 5.3, 6.1, 4.9, 3.6, 6.3, 5.9, 6, 6.8, 7.9, 7.1, 9.3, 8.5, 
    8.9, 7.9, 5.6, 7.2, 4.1, 6, 4.6, 10.1, 2.4, 2.1, 5.3, 3.6, 6.4, 9.2, 9.7, 
    8.3, 4.3, 3.5, 3.4, 4, 3.3, 6.1, 3.8, 4.6, 6.3, 7.5, 7.9, 7.4, 3.5, 3, 
    6.4, 11.4, 10.4, 9.5, 8.2, 8.1, 2.9, 3.6, 4.9, 3.9, 2.6, 5.5, 3, 4.1, 
    4.3, 2.8, 1.7, 1.5, 8.4, 2.3, 2.2, 4.3, 1, 2.1, 0.2, 0.6, 2.3, 4.6, 9, 
    8.2, 1.5, 1.1, 3.1, 2.5, 0.8, 4, 4.7, 1.5, 2.9, 2, 0.9, 1.8, 0.5, 3.2, 
    3.8, 2.2, 4, 5.4, 3.5, 2.4, 1.7, 3.4, 0.7, 3.6, 1, 0.8, 3.4, 0.4, 0.4, 
    0.4, 0.4, 1.8, 0.9, 0.3, 1.4, 4.4, 1, 1.3, 2.1, 7.1, 1.4, 3.1, 0.5, 2.1, 
    1.6, 0.7, 4.3, 0, 0.6, 5.9, 2.8, 4.8, 1.3, 0.7, 1.5, 1.5, 1.3, 3.1, 2.2, 
    0.4, 0.1, 0.2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0.2, 0.3, 
    0, 0.2, 0, 0.3, 0.1, 0, 0.2, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0.2, 0, 0, 0, 0, 
    0.1, 0, 0.2, 0.3, 0.4, 0, 0, 0.1, 1.4, 0.8, 0.8, 2.2, 0.1, 0.8, 0.4, 0, 
    2.3, 0, 0.7, 4.3, 5.9, 5.5, 2.6, 3.6, 3.9, 4.3, 4.5, 6.7, 4.6, 6.5, 4.9, 
    7.4, 6.8, 4.5, 3.4, 4, 2.7, 1.2, 0.1, 0, 0, 1.1, 0.8, 0.1, 0, 0, 0.3, 0, 
    0.1, 0.4, 0.8, 0.6, 0.4, 3.1, 1, 3.8, 2.1, 2.4, 8.1, 2.2, 1.7, 4.6, 5.1, 
    2, 2.3, 1.2, 4.2, 2.7, 3.6, 1.9, 2.9, 1.9, 1, 1.1, 1.9, 2, 0.3, 2.2, 0.1, 
    0.5, 0.1, 0, 0.1, 0.5, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0, 0.2, 0, 0, 0.2, 0, 
    0.4, 0.7, 0.3, 0, 0, 0, 0.2, 0.1, 0, 0, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0, 0, 
    0, 0.1, 0.8, 0.3, 0, 0.2, 0.2, 0, 0, 0, 0, 0.1, 0.1, 0, 0, 0.1, 0, 0, 0, 
    0.1, 0, 0.2, 0, 0, 0.1, 0, 0, 0.3, 0, 0.3, 0, 1.3, 0, 0, 0, 0, 0, 0.3, 
    0.1, 0.1, 0.4, 0.2, 1, 0.1, 0.4, 0.6, 0.2, 0, 1, 1.2, 1.3, 0.6, 1.3, 1.1, 
    0.2, 0.1, 0, 0.1, 0.1, 0.1, 0, 0, 0, 0.1, 0, 0, 0.1, 0, 0, 0.1, 0.1, 0.4, 
    0.1, 0, 0.3, 0.3, 0.3, 0.3, 0.3, 0.1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2, 
    0, 0, 0.3, 0.2, 0.1, 0, 0, 0, 0, 0, 0.2, 0.1, 0, 0.4, 0, 0.1, 0.2, 0.3, 
    0.3, 0, 0.2, 0.4, 0, 0, 0.4, 0.4, 0.2, 0.4, 0.1, 0.1, 0, 0, 0, 0.6, 0.7, 
    1.6, 0, 0.1, 0, 0.5, 4.4, 3.9, 5.1, 4.5, 4.2, 3, 4.6, 3.4, 3.3, 2, 3.3, 
    3.5, 0.1, 0.1, 0, 2.8, 3.2, 2.1, 1.5, 1.4, 0.4, 0.5, 0.6, 0.2, 2.3, 0.3, 
    0, 0, 0, 0, 4.3, 5.8, 5.8, 6.7, 6.3, 4.7, 5.6, 5.4, 4.3, 3.6, 3.3, 4.2, 
    5.2, 4.2, 4.4, 4.5, 5.6, 6.5, 5.1, 5.2, 5, 4.8, 4.6, 4.5, 0.7, 2.9, 2.7, 
    2.5, 1.9, 2.1, 2.3, 5.8, 4.7, 4, 2.6, 0.1, 2.2, 2.4, 3.3, 0.2, 0.4, 1, 
    0.5, 0.1, 0.6, 1, 0.1, 6, 6, 5, 5.6, 4.9, 3.5, 3.9, 2.8, 4.1, 4.8, 2.3, 
    3.6, 2.9, 4.4, 4.4, 5, 5.1, 5.6, 4.4, 1.9, 1.7, 5.1, 6, 8.5, 7, 4.3, 5, 
    6.4, 7.1, 5.2, 4.1, 3.7, 3.7, 2.6, 2.8, 3.5, 3.1, 2.7, 0.8, 0.1, 0, 0, 0, 
    0, 0.2, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.3, 0, 0.5, 
    0.2, 0.7, 0.1, 0.7, 2.6, 1.3, 0.8, 0.9, 1.1, 5.3, 7.5, 8.7, 7.5, 7, 5.5, 
    4.5, 6, 6.8, 5.2, 3.8, 6.1, 2.3, 4, 5.8, 8.2, 5.2, 2.9, 3.2, 5.2, 3.4, 
    2.6, 1.3, 0.9, 1.5, 1, 0.3, 0.2, 0.4, 0.6, 0.1, 0.2, 0.7, 0.3, 0.1, 2, 
    2.5, 0.6, 0.2, 0, 1.7, 0.1, 1.1, 0.7, 0.4, 0, 0.6, 0.8, 0, 0, 0, 0.2, 0, 
    0, 0, 0, 0.3, 0.9, 0.5, 0.1, 0, 0, 0.3, 0.1, 0.8, 0.1, 0.5, 0.3, 0.1, 
    0.1, 0.1, 0, 0, 0, 0, 1, 0.9, 0.2, 0, 0.1, 0.2, 1.1, 0.5, 0.2, 2.1, 2.3, 
    0.3, 0, 1.8, 1.8, 0.4, 0.8, 0.2, 0.3, 0, 0.1, 0, 0.7, 0, 0, 0.1, 3.1, 
    2.2, 0.6, 0.4, 0.2, 0.1, 0, 0, 0, 0, 0, 0, 0.1, _, _, _, _, _, _, _, _, 
    _, _, _, 0, 0, 0, 0, 4.9, 0, 2.1, 0, 0, 0, 0, 0.2, 0, 0.1, 0.9, 1.5, 0.4, 
    0, 0, 0, 0, 0, 0.8, 1.8, 0.1, 0, 0, 0, 0, 0.2, 0.1, 0, 0, 0.2, 0, 0, 0, 
    0, 0, 0, 0.1, 0.9, 0.4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1, 0, 0, 0.1, 
    0.1, 0.1, 0.3, 0, 1.4, 0.3, 0.1, 0.3, 0.3, 0.4, 0, 0.2, 0, 0, 0.2, 0.2, 
    0, 0, 0, 0.2, 3, 2.1, 0.8, 1.5, 2.5, 0.5, 0.2, 1.4, 2.1, 9.1, 11.8, 10.1, 
    7.7, 3.2, 2.8, 1.5, 3.8, 0.1, 2.1, 0.7, 0.3, 1.2, 0.4, 2.6, 6.4, 4.1, 
    1.9, 8.6, 8.5, 6, 6.3, 6.7, 4.6, 4.6, 4.5, 0.2, 0.4, 3.5, 8.1, 5.6, 1.7, 
    1.7, 1.7, 6.9, 1.9, 3, 2.8, 1.8, 2.4, 1.8, 9.4, 9.8, 9.5, 3, 4.4, 3.8, 
    0.8, 3.3, 3.7, 2.9, 2.5, 4.4, 2.7, 3.8, 4.8, 2.5, 3.2, 4.7, 4.7, 2.9, 
    4.1, 5.1, 2.8, 3.3, 1.5, 0.9, 7.6, 2.8, 3.1, 6.8, 5.7, 7.2, 9, 8.5, 6.1, 
    4.8, 8, 7.1, 5.9, 7.3, 8.3, 6.5, 4.2, 5.2, 7.3, 2.5, 6.7, 5.4, 4.6, 3.5, 
    6.4, 6, 3.8, 6.1, 6.5, 4.2, 6.1, 4.3, 4.9, 5.9, 5.1, 7.3, 3.5, 3.6, 3.5, 
    5.9, 5.3, 4.8, 4.2, 2.9, 5.7, 5, 3.7, 2.4, 1.1, 1.7, 0.9, 4.6, 6.9, 5.7, 
    5.8, 2.7, 0.5, 0.8, 0.4, 0.3, 0.7, 0.2, 1.7, 0, 0.3, 0.7, 0.8, 0.9, 1.3, 
    1.1, 1, 0.8, 1.7, 0.8, 0.3, 0.6, 0.9, 2.9, 0.9, 0.5, 1.2, 1.3, 0.2, 0.4, 
    5.7, 5.3, 5.1, 2.6, 3.4, 1.1, 2.4, 3.4, 0.9, 1.2, 2.3, 1.4, 2.7, 1.8, 2, 
    2, 5.5, 0.4, 0.6, 0.8, 1.8, 1.8, 1.8, 0.8, 3.2, 0.7, 1, 1.7, 1.1, 1.2, 2, 
    2.3, 1.9, 2.6, 0.9, 0.8, 0.6, 4.4, 6.4, 7.1, 4.6, 2.6, 3.2, 1.5, 2.1, 
    3.3, 2.1, 0.5, 0.1, 2.9, 4.2, 0.3, 4.7, 3.1, 3.2, 3.3, 3.4, 3.5, 3.6, 
    3.3, 2.2, 2.4, 2.1, 2.9, 2.4, 4.9, 2.4, 1.6, 3, 4.6, 3.9, 4.9, 4.4, 4.5, 
    4.5, 4.7, 5.4, 4.9, 7.7, 4, 4.4, 5.3, 4.7, 4.2, 4.2, 4.2, 5.9, 0.4, 2.8, 
    2.6, 0.3, 2.1, 1.3, 0.5, 0.5, 0.4, 0.4, 0.1, 0.7, 0, 1.1, 1, 1, 1.8, 0.8, 
    0.6, 1.2, 0.5, 1, 0.8, 2, 0.6, 0.7, 1.2, 0.4, 0, 0.1, 0, 0, 0, 0.1, 0, 0, 
    0.6, 0.4, 1.5, 1.7, 2.9, 1.5, 0.5, 0.8, 0.3, 0, 0.1, 0, 0.1, 0.1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.4, 0.5, 0.9, 0.9, 7.1, 5.6, 3.7, 6.3, 4.3, 4, 2.2, 
    5.1, 4.8, 4.5, 7, 6.5, 5.1, 4.6, 4.5, 3.4, 3.8, 3.7, 3.3, 2.5, 2.4, 0, 
    0.5, 5.5, 7.2, 8.2, 4.8, 4.1, 0.1, 3.1, 6.5, 6.4, 7.2, 7.6, 7.6, 6.7, 
    2.4, 1, 1.1, 0.6, 1.2, 1.3, 0.1, 1.7, 1, 0.3, 0.2, 0.7, 0.5, 0, 0.1, 0.3, 
    0, 0.4, 0.3, 0, 0.1, 0.4, 0.3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.3, 
    0.3, 0.2, 0.2, 1.2, 4.9, 5.8, 0.9, 3.9, 4.5, 4.8, 4, 4.4, 3.7, 4, 3.3, 
    3.9, 5.2, 4, 4, 3.7, 2.1, 2.1, 0.5, 1.4, 0.1, 2.9, 0.7, 1.2, 0.8, 0.3, 
    1.5, 5.1, 1.2, 0.8, 0, 1.4, 1.4, 0.9, 0.7, 0.1, 0, 0.2, 0.4, 0.7, 0.4, 
    0.5, 0.4, 0.1, 7.6, 1.1, 0.2, 0.3, 0.2, 0.4, 0.6, 0.3, 0.1, 7.2, 0, 0, 0, 
    6.4, 0, 0.1, 0, 0, 0, 5.4, 0, 0, 0, 0.1, 0.2, 0.1, 0, 0, 0.1, 0.2, 0.1, 
    0.1, 0.4, 0.4, 0, 0, 0, 0.1, 0, 0.1, 0.2, 0, 0.2, 0.5, 0.4, 0.7, 0.1, 
    0.6, 0.6, 0.4, 0.4, 0.6, 0.2, 0.3, 1.3, 0.7, 0.6, 0.5, 0.1, 0, 0, 0, 0.2, 
    0, 0, 0, 0.1, 0, 0.3, 0.2, 0.5, 0.4, 0.1, 1.4, 2.3, 3.1, 4.2, 4.8, 6.1, 
    5.6, 4.5, 5.7, 4.8, 4.5, 3.6, 3.7, 3, 2.8, 2.2, 3, 3.5, 2.1, 0.9, 3, 2, 
    1.1, 3.4, 2.5, 2.1, 1.3, 2.1, 2, 2, 1.4, 1.5, 1.9, 1.7, 3.8, 2.8, 4.8, 
    5.3, 4.8, 1.2, 1.4, 1.5, 1.3, 0.6, 1.2, 0, 0.9, 1.4, 1.7, 0.3, 0.8, 2, 
    1.7, 1.6, 2, 5.1, 1.7, 3.5, 3.5, 1.5, 2.5, 1.6, 1.4, 1, 0.9, 2.5, 3.9, 
    2.6, 3.5, 3.5, 2.1, 2.6, 3.1, 4.6, 5, 1.3, 1.8, 3, 2.6, 4.2, 5.6, 3.5, 
    1.3, 3.4, 1.1, 3.1, 3.7, 3.2, 1.4, 1.3, 2.8, 2.2, 1.3, 3.8, 4.6, 3.2, 
    5.9, 4.9, 5.3, 6.3, 6.3, 5.4, 4.3, 4.1, 1.8, 2.8, 1.7, 1.5, 1.1, 1.9, 
    0.3, 3.3, 0.1, 1.5, 6.4, 4, 3.5, 3.5, 3.6, 1.5, 2.7, 1.9, 3.9, 5.6, 4.4, 
    5.3, 4.7, 1.5, 3.4, 2.3, 3.8, 3.1, 2.9, 2.5, 2.6, 4.4, 3.9, 5.4, 3.1, 
    2.9, 3.6, 4.1, 4.3, 4.3, 3.5, 3.8, 4.3, 3.2, 1.2, 3.3, 1.7, 0.9, 1.1, 
    3.9, 1.9, 1.3, 1.8, 0.7, 1.3, 1.1, 0.1, 1.3, 0.5, 0.4, 1, 2.3, 3.2, 3.1, 
    2.3, 2.3, 1.8, 2.2, 2.1, 2.8, 2.2, 2, 2.3, 0.8, 2.2, 0.9, 0.7, 1, 3.1, 1, 
    1, 0.4, 0.7, 1.6, 0.2, 1, 0.2, 1, 0.9, 0.5, 2.1, 0.9, 1, 1.9, 3.9, 1.1, 
    1.7, 0.7, 0.6, 0.2, 0, 0.3, 0.1, 0.1, 0.4, 0.7, 0.6, 0, 0.1, 1, 0.8, 0.5, 
    0, 0.5, 0.1, 0, 0.1, 0.6, 0.1, 2.2, 2.2, 2.8, 3.8, 4.8, 6.1, 7.5, 5.7, 
    5.8, 4.8, 6.4, 5.2, 5.8, 4.5, 3.3, 5.7, 4.3, 4.5, 1.9, 1.7, 3.9, 4.2, 
    4.6, 3.8, 1, 3.3, 6.4, 5.3, 6.1, 6.9, 7.7, 4.6, 4.5, 7.1, 5.6, 6.1, 5.1, 
    6, 4.5, 3.8, 6.1, 5.5, 4.1, 7.5, 10.5, 5.1, 3.4, 3.6, 5.4, 5.4, 4.6, 3.3, 
    3.2, 1, 4.7, 4.4, 3.1, 3.1, 2.5, 0.9, 4, 4, 4.1, 4.1, 4.6, 5.2, 4.1, 1.6, 
    1.2, 3.9, 5.4, 3.4, 3.1, 1.7, 0.1, 0.7, 0.9, 2.7, 1.9, 0.3, 0, 0, 0.5, 
    0.4, 0.4, 1.6, 3.5, 1.9, 3.3, 1.3, 4.2, 4.1, 2.1, 2.9, 3.2, 2.7, 2.3, 
    1.9, 3.8, 1, 0.3, 0.2, 4.2, 6.3, 3.2, 2.3, 1.8, 1.7, 2, 2.1, 0.6, 0.6, 
    0.6, 2.6, 3.6, 0.8, 0.8, 1, 1.7, 1.7, 1.4, 1, 0.2, 0.8, 1.7, 0.6, 1.1, 
    0.5, 1.1, 1, 0.8, 0.4, 2.7, 2.1, 0.8, 0.4, 0.9, 4.4, 2, 2.1, 1, 1.2, 0.5, 
    0.9, 0.7, 3.7, 3.5, 0.7, 0.3, 1.5, 0.9, 1.1, 0.8, 0.5, 0.5, 0.8, 1, 1.1, 
    1.1, 1.4, 4.9, 4.6, 4, 4.1, 2.3, 1.3, 1.2, 1.6, 1.1, 0.6, 2.4, 2, 1.2, 
    0.5, 3.7, 3.9, 4, 1.5, 3.4, 3.4, 3.1, 3, 4.1, 4, 4.2, 3.6, 3.6, 3.5, 3.5, 
    3.5, 3.5, 4.6, 4.7, 5, 4.7, 4.3, 3.7, 3.1, 4.5, 3.3, 4.1, 3.7, 1.8, 3.1, 
    3.8, 5, 4.9, 5.5, 5.5, 5.4, 4.6, 4.6, 5, 4.5, 4.6, 4.7, 4.3, 4, 4, 3.1, 
    3.4, 3.6, 2.8, 3, 3.9, 3.1, 3.4, 4.6, 3.8, 4.1, 4.2, 3.5, 3.3, 4, 3.6, 
    4.7, 3.3, 2.9, 2.2, 0.6, 1.1, 2.3, 1, 1.2, 0.8, 1.4, 2.7, 3, 2.1, 2.4, 
    2.1, 2.6, 3.7, 5.8, 4.1, 3.8, 4.5, 3, 2.3, 1.4, 4.5, 2, 1.7, 2, 2.4, 2.8, 
    1.9, 2.9, 2.9, 1.1, 1.2, 0.9, 0.7, 0.3, 1, 0.1, 1.8, 2, 2.1, 1, 2.1, 1.5, 
    1.1, 0.9, 3.5, 3.1, 2.6, 2.2, 1.5, 1.2, 0.9, 1.5, 1, 0.2, 0.8, 2.3, 0.2, 
    0, 0, 0, 1, 0.5, 0.3, 0.4, 1.3, 2, 2.2, 2.3, 2.2, 2.5, 2.2, 1.6, 1.9, 2, 
    2, 2.7, 2.9, 3.2, 2.9, 2, 1.6, 1, 1, 0.5, 0.5, 0.6, 3.1, 1, 2.2, 1.8, 
    2.3, 2.1, 2.6, 2.1, 2, 3, 2.5, 2.3, 2.1, 0.8, 2.3, 2.5, 0.6, 0.6, 1, 2.5, 
    1.5, 0.5, 0.2, 1.8, 1.5, 3.2, 3.6, 5.4, 5.5, 5.5, 3.3, 3.1, 3, 2.9, 2.1, 
    0.9, 1.6, 0.9, 1.8, 1.7, 2.1, 1, 0.9, 0.4, 1, 0.7, 1.8, 1.6, 1.4, 1.9, 
    1.5, 1.2, 1, 1.6, 1.6, 1.8, 2, 2.2, 2.5, 1.5, 1.5, 2.5, 0.5, 0.1, 0.2, 
    2.5, 0.9, 0.1, 2.5, 2, 0.9, 1.5, 1.8, 2.4, 2.2, 2.9, 2.6, 0.7, 5.3, 0.9, 
    6.3, 2.3, 2.6, 1.8, 2.5, 1.9, 2.1, 1.1, 1.2, 0.5, 4.4, 0.6, 1.7, 5.3, 
    4.5, 1.1, 1.5, 3.5, 3.6, 0.6, 1.1, 2.9, 3, 6, 2.2, 0.8, 3.7, 1.4, 3.2, 
    2.2, 3.9, 1, 5, 0.7, 1.4, 0.5, 1.1, 0.8, 2.5, 2.7, 1.6, 1.4, 1, 1.3, 0.6, 
    3.8, 2.5, 2, 2.8, 3.6, 2.3, 3.2, 2.2, 2, 1.7, 0.3, 0.6, 1.2, 0.5, 1.1, 
    0.6, 0.7, 0, 1.4, 1.5, 2, 3.1, 1, 6.1, 5.7, 5.6, 6.9, 7.4, 5.9, 2.9, 3.4, 
    5.7, 2.9, 0.6, 0.1, 0, 0, 0.1, 0.6, 0.8, 0.8, 0.3, 0.6, 0.6, 3.2, 4.6, 
    3.8, 1.1, 1.1, 1, 0.3, 1.6, 0.7, 1, 1, 3.2, 1.9, 4.5, 0.3, 1.2, 0.9, 0.6, 
    0.1, 0, 0.2, 0, 0.3, 0.3, 0.8, 2.6, 3.1, 2.6, 2.1, 2.6, 2.1, 2.7, 2.8, 
    3.1, 3.4, 4, 4.2, 4.6, 2.2, 0.2, 0.2, 0, 0.1, 0.4, 1.6, 2.4, 2.2, 1.9, 
    1.6, 1.7, 2.1, 2.4, 2.6, 2.8, 4.6, 4.3, 2, 3.9, 2.9, 3.3, 3.5, 2.2, 1.4, 
    0.9, 0.3, 1.5, 1.7, 1, 1, 1.7, 1.8, 2.2, 1.9, 1.4, 1.9, 1.6, 1.3, 1.5, 
    1.8, 2.5, 2.3, 1.9, 2.3, 1.5, 1.9, 1.7, 1, 1.7, 2, 0.9, 1.3, 1.5, 1.4, 
    1.5, 1, 1.2, 2.3, 2, 2, 2.1, 2, 2.1, 2.1, 2.7, 3.1, 3, 1.8, 2.2, 3.3, 
    2.9, 4, 1, 0.2, 2.1, 0.4, 1, 2.6, 0.8, 1.6, 1.8, 2.4, 1.8, 1.7, 1.9, 1.8, 
    2.5, 2.8, 3.6, 3.9, 3.7, 2.7, 2.3, 0.9, 2.8, 2.5, 1.3, 3, 0.8, 2.5, 1.6, 
    2, 3.3, 4.2, 3.2, 3.3, 2.1, 2.7, 2, 1.2, 2.6, 0.6, 4, 3.3, 4, 3, 4.7, 
    3.7, 4.8, 4.7, 4.6, 3.8, 2.9, 1.5, 2.6, 0.7, 0.2, 1.6, 1.8, 1.8, 1.7, 
    1.1, 1.1, 0.8, 0.6, 1.6, 0.7, 1.2, 1.9, 0.3, 0.8, 0.7, 0.7, 0.9, 0.7, 
    0.6, 0.1, 0.7, 1, 2.2, 1.9, 1.4, 2.5, 1.9, 1.1, 1, 0.6, 1.9, 5.4, 6.4, 6, 
    3.2, 4.7, 4.6, 5.4, 8.5, 7, 6.7, 7.6, 5.8, 2.6, 3.1, 2.7, 3.1, 3.4, 5.1, 
    5.7, 7.4, 3.5, 2.6, 2.4, 2, 2.8, 2.9, 3.8, 3.7, 4.8, 4.1, 2.1, 1.8, 1.7, 
    3.3, 6.8, 3.7, 3.7, 5.6, 8.2, 2.1, 4.1, 5.3, 5.8, 6.8, 1.9, 5.8, 5.6, 
    3.3, 2.9, 3.3, 2.9, 3.9, 2.2, 6.4, 4.8, 3.7, 4.7, 5.2, 1.8, 4.6, 4.8, 
    2.4, 6.2, 1.5, 5.3, 3.9, 3.9, 3.7, 3.2, 3.9, 4.3, 4.6, 3.3, 3.6, 6.4, 
    4.6, 5.7, 6.4, 1.9, 2.3, 7.3, 6.7, 4.3, 5.2, 8.2, 8.9, 6.9, 4.2, 5, 1.7, 
    4.8, 7.8, 2.3, 7.5, 7.2, 6, 6, 6, 3.9, 6.5, 7.3, 4.7, 5.1, 5.9, 5.5, 3.7, 
    6.8, 7.5, 5.6, 4.5, 5.1, 4.1, 2, 2.6, 3.4, 4, 4.9, 3.3, 5, 3.3, 3.4, 3.2, 
    5, 3.5, 2.8, 6, 3.5, 2.5, 3, 3.6, 3.3, 1.5, 0.7, 2.4, 3, 3.4, 3.6, 2.3, 
    1.3, 0.5, 0.8, 0.4, 0.2, 0.2, 0, 0, 0.2, 0.4, 0.6, 2, 0.9, 0.1, 0, 0.1, 
    0.1, 0, 0, 0.1, 0, 0, 0, 0.2, 0.3, 0.5, 0.8, 1.2, 0.6, 1.5, 1.7, 2.1, 
    1.3, 1.8, 1.3, 2.4, 3, 4.6, 4.6, 5.8, 6.6, 6, 4.2, 4.6, 3.2, 3.2, 4.7, 
    5.9, 6.1, 8.3, 6.9, 6.7, 4.2, 3, 0.3, 4.6, 2.3, 4, 3.1, 2.3, 3.2, 3, 2.3, 
    0.1, 2.3, 0.7, 1, 1.1, 0.3, 0.5, 0.6, 0.7, 0.8, 1, 0, 0.1, 0.2, 0.9, 0.2, 
    0.4, 1.6, 1.2, 1.9, 2, 0.2, 0.3, 1.2, 0.8, 0.3, 0.9, 1, 0.9, 0, 0, 0, 
    0.6, 1.1, 0.8, 0.6, 0.8, 1.7, 1.2, 1.2, 1.4, 1.7, 1.5, 1.5, 1.1, 1.2, 
    0.1, 0, 0.1, 0.9, 0, 0.5, 0.6, 0.8, 0.8, 0.2, 2.8, 2, 1.4, 0.1, 0.9, 0.3, 
    0.3, 0.8, 0.9, 0.4, 1.4, 1.2, 2.8, 0.2, 0.4, 0.8, 1.9, 0.5, 0, 0.4, 0.4, 
    0, 0.6, 1.6, 2.3, 0.7, 3, 3.1, 3.5, 3.8, 4.6, 5, 4.2, 4.6, 3.8, 3.4, 5.1, 
    0.7, 1.5, 0, 2.3, 1.3, 0.4, 1.8, 1.6, 2.5, 2.5, 2.8, 2.4, 2.3, 2.7, 2.7, 
    2.8, 2.8, 2.6, 2.5, 2.3, 2.2, 2.2, 2.3, 2.3, 2.3, 2.2, 1, 0.7, 0.8, 1.1, 
    0.4, 1.1, 1.7, 1.6, 1.2, 0.9, 1.2, 1.7, 2, 1.3, 1.5, 1.7, 2.6, 2.3, 2.5, 
    3.1, 3, 3, 2.6, 3.8, 1.3, 1.1, 3.9, 4.9, 3.4, 3.7, 2.6, 1.6, 1.8, 1.9, 3, 
    4, 3.4, 4.2, 4.5, 4.3, 3.9, 4, 2.6, 2.9, 2.8, 3.6, 2.5, 1.9, 2.8, 1.9, 
    2.1, 2.1, 2, 1.8, 2.4, 2.6, 1.7, 3.6, 4.7, 4.7, 3.8, 3.5, 3.2, 3.1, 1.7, 
    0.7, 0.8, 1.9, 1.8, 2.6, 2.5, 1.2, 2.9, 3.5, 3.5, 2.9, 2.5, 0.4, 1.7, 
    1.4, 1, 0.2, 3.9, 4.1, 4.7, 3.9, 4, 4, 4, 4.7, 2.3, 1.9, 3.2, 1.8, 4.3, 
    3.9, 3.2, 2.6, 2.8, 3, 3.4, 3.8, 3.7, 4, 3.8, 3.1, 2.6, 1.8, 1.9, 2, 2.2, 
    2.2, 2.2, 2.3, 2.1, 2.2, 2.1, 2.2, 2.3, 2.7, 2.5, 2.2, 1.9, 1.9, 2, 2.5, 
    2.2, 2, 1.8, 2.6, 2.7, 3.7, 0.9, 2.6, 4.2, 2.7, 5.1, 5.1, 4.4, 4.5, 5.4, 
    4.5, 4.4, 3.9, 3.7, 2.4, 2.5, 2.6, 3.1, 3.9, 2.8, 1.7, 2, 0.9, 1, 1.6, 
    1.7, 1.9, 2.2, 2.1, 4.6, 2.8, 4.7, 2.7, 2, 2.1, 1.8, 1.7, 1.8, 1.2, 1.2, 
    1.2, 0.4, 0, 0, 1.5, 2.6, 3.6, 3.3, 3.2, 3, 3.6, 2.3, 0.9, 1.4, 1.5, 4.2, 
    5, 4.4, 5, 4.3, 4, 2.9, 4.8, 4.1, 5.9, 4.1, 4, 3.8, 3.8, 3.8, 4.5, 3.2, 
    3.4, 3.4, 3.4, 3, 1.1, 1.4, 2.6, 2.7, 3.2, 1.9, 1.3, 0.9, 0.7, 0.3, 0.5, 
    0.5, 0.5, 0.4, 0.2, 0, 0, 0.6, 0.3, 0.7, 0, 1.8, 2.3, 1.6, 2, 2.7, 2.7, 
    1.6, 1.6, 3.3, 1.8, 1.4, 0.5, 0.9, 4, 4, 4.2, 3.4, 3.4, 3.4, 2.4, 2.6, 
    0.8, 0.1, 3, 3.7, 2.3, 2.6, 2.8, 3, 0.8, 4.3, 5.2, 4.6, 3.8, 4, 2, 2.4, 
    2.3, 3.6, 1.5, 1.2, 1.6, 3.1, 2.8, 2.8, 2.7, 2.9, 2.5, 2, 2.9, 3.3, 1.2, 
    1.9, 1.3, 2.7, 4.2, 2.9, 2.5, 1.7, 0.6, 0.5, 0, 0.2, 0.3, 0.3, 0.2, 0, 
    0.4, 1, 0.3, 0.8, 0.9, 0.8, 1.3, 1.1, 0.5, 2.3, 1.3, 0.9, 0.9, 1.4, 1.6, 
    2.2, 1.2, 1.3, 0.6, 1.3, 1, 1.2, 0.7, 0.5, 0.4, 0.5, 1.8, 3, 4.3, 4.6, 
    4.7, 5.8, 1.3, 5.4, 2.8, 2.4, 1.8, 4.4, 5, 3.3, 2.8, 4.5, 2.1, 0.9, 0.5, 
    0.8, 0.9, 1.5, 1.1, 0.6, 0, 0.9, 1.3, 1.2, 1.3, 1.8, 2, 2.5, 3.2, 3.1, 
    3.5, 2.6, 2.3, 2.3, 2.6, 1.8, 1.7, 1.6, 0.5, 0, 0, 0, 0.6, 0.1, 1, 0.1, 
    0.6, 1.7, 1.7, 1.6, 1.7, 1.9, 1.8, 2.1, 2.2, 2.3, 2.3, 2.5, 4.2, 2.4, 3, 
    1.9, 1, 0.6, 0.6, 0.3, 1.6, 1.5, 2.3, 1.5, 0.9, 2, 5.5, 1.8, 4.7, 5.4, 6, 
    4.4, 5.3, 1.8, 1.6, 1.6, 0.4, 2.3, 0.9, 0.5, 0.6, 0.6, 0.5, 0.2, 0.8, 
    1.1, 1.8, 1.7, 0.5, 1.5, 0.9, 1.6, 1.1, 1.7, 1.6, 1.5, 1.6, 1.8, 0.8, 
    0.2, 0.9, 0.6, 0.6, 0.3, 0, 0.3, 1.9, 0.1, 2.2, 2.2, 3.6, 2.8, 2.2, 2.4, 
    2.3, 2.3, 2.7, 2.5, 3, 2.9, 3.3, 2.4, 3.2, 3.6, 2.2, 3, 1.5, 1.2, 0.9, 2, 
    0.4, 0, 1.2, 0.8, 1.3, 1.7, 1.3, 1.5, 1.8, 1, 0.8, 0.9, 1, 0.4, 0.6, 0.8, 
    0.4, 1.6, 1.6, 1.4, 2.4, 0.4, 0.1, 0.3, 0.5, 1.5, 1.8, 0.5, 0.7, 0.7, 
    0.3, 0.9, 1.2, 1.7, 1.9, 0.9, 1.1, 0.2, 0.8, 0.5, 2.3, 3.9, 1.7, 1.9, 
    0.5, 0.6, 0.7, 0.7, 0.5, 0.3, 0, 0.5, 1, 1, 1.9, 2.7, 1.8, 1.3, 1, 1.6, 
    2.1, 2.1, 1.8, 2.5, 1.3, 3.8, 3.3, 1.1, 2.5, 1.4, 1.6, 1.1, 1.6, 0.6, 
    2.8, 2.4, 1.8, 3.5, 2, 2.1, 2.6, 2, 2, 1.6, 2.1, 2.4, 1.8, 2.1, 1.9, 2.1, 
    1.9, 2.6, 0.8, 0.6, 0.9, 0.8, 0.7, 0.5, 0.4, 0.3, 0.6, 1, 0.9, 1.1, 1.5, 
    1.4, 1.4, 2, 2.3, 2.1, 2.8, 3.4, 3.6, 4.2, 3.3, 2.8, 2, 2, 1.9, 1.5, 2, 
    3.5, 2.6, 1.9, 1.4, 1.8, 1.6, 1.5, 1, 0.7, 1.6, 1.1, 1.9, 1.8, 1.3, 1.1, 
    0.7, 0.6, 0.6, 0.3, 1.1, 1.2, 1.1, 1, 0.1, 0.1, 0, 1.6, 1.4, 0.7, 1.4, 
    1.3, 1.7, 2.1, 3, 3, 3.1, 2, 1.1, 1, 2.8, 3, 3.1, 2.1, 2, 1.1, 0.2, 0.3, 
    0.5, 0, 0, 0, 0.1, 0.3, 0.8, 2.2, 3.1, 3.3, 2.9, 2.8, 2.3, 1.7, 2.4, 0.8, 
    0.8, 1, 1.1, 4.7, 6.8, 3.7, 0.7, 3, 5.7, 3.9, 3.7, 5.2, 4, 1.3, 2.4, 4.5, 
    4.7, 2.6, 1.7, 1.9, 2.2, 2.4, 1.5, 1.6, 2.9, 2.6, 2.7, 2.8, 3, 3.2, 2.7, 
    1.1, 0.7, 0.1, 0.4, 1, 0.5, 0.9, 1, 2.5, 2.9, 3, 2.4, 2.8, 2.8, 1.5, 2.4, 
    2, 1.4, 1.4, 1.4, 0.9, 0.4, 0.8, 1.3, 1, 0.9, 0.4, 0.2, 0.1, 0.2, 0.4, 
    0.7, 1.9, 0.6, 0.5, 0.5, 0.5, 0.5, 0.7, 0.9, 0.4, 2.4, 2.5, 1, 3.4, 2.3, 
    1.3, 1.3, 0.3, 0.1, 0.2, 0.1, 3.2, 2.6, 0.8, 1.5, 5.7, 5.4, 5.2, 5.7, 
    5.7, 5.1, 5.7, 4.6, 3.3, 3.9, 6, 3.7, 3.6, 4.9, 1.5, 3.9, 3.9, 1.5, 1.1, 
    2.2, 4, 2.8, 3, 5.7, 5.2, 6.1, 6.3, 5.8, 4.8, 6.6, 6, 6.3, 5, 6.6, 5.4, 
    1.9, 3, 0.9, 5.2, 4.2, 5.1, 4.5, 2.6, 0.6, 5.1, 3.6, 3.4, 1.1, 2.9, 5.3, 
    3.6, 3.7, 6.5, 3.1, 7, 6.9, 6.4, 2.5, 1.5, 1.2, 1.2, 1.7, 4.3, 3.1, 2.2, 
    3.4, 5.7, 4.3, 4.7, 0.9, 3.3, 2.7, 0.9, 4.9, 6, 4.1, 3.6, 3.9, 3.1, 2.3, 
    1.5, 1.7, 0.2, 3.6, 5.1, 3.7, 5.4, 4.6, 6.1, 5.6, 5.6, 5.2, 5.4, 4.9, 
    5.8, 4, 4, 3.2, 3.7, 3.4, 3.2, 4.6, 4.1, 3.6, 4.2, 4, 3.6, 3.3, 1.7, 2.4, 
    0.2, 0.2, 2.8, 0.1, 0.9, 0.4, 0.6, 0.1, 0.9, 0.9, 1.8, 3.1, 1.6, 2.9, 
    0.9, 3, 0.7, 2.3, 0.4, 0.7, 0.9, 0.4, 0.2, 0.8, 2.1, 1.6, 0.2, 0, 0.6, 
    0.1, 3.8, 3, 1.7, 3.9, 3.7, 1.8, 0.7, 1.4, 0.8, 1.1, 2, 1.9, 1.6, 4.6, 
    3.8, 4.7, 3.6, 2.6, 3.9, 2.9, 3.9, 4.6, 4.9, 5.7, 3.7, 4.2, 2.4, 3.1, 
    3.7, 4.5, 4.3, 3.8, 4.8, 4, 4.2, 3.7, 5.3, 4.3, 2.1, 2.8, 2.8, 3.2, 3.5, 
    3.7, 3.9, 3.2, 2.5, 2.8, 0.6, 2.3, 1.5, 1.5, 2.3, 1.7, 1.7, 1.2, 3.1, 
    4.5, 3.1, 0.4, 1.1, 1.7, 2.1, 2.8, 2.3, 1.2, 0.2, 1, 0.2, 0, 0, 0, 0, 
    2.9, 3.2, 0.6, 0.7, 2.8, 2.6, 3.5, 3.5, 3.9, 3.5, 3.5, 2.5, 2.3, 1.8, 
    1.9, 2, 2, 2.1, 1.2, 0.6, 1.1, 0.5, 1, 0.7, 1, 1.3, 1.5, 2, 2.3, 1.8, 
    5.9, 6.6, 7.6, 6.8, 6.8, 6.2, 8.5, 5.1, 3.9, 4.2, 5.4, 6, 8.5, 8, 6.1, 
    6.9, 5.1, 2.7, 1.7, 2.7, 1.8, 3.4, 4.2, 2.2, 2.2, 6.2, 5.6, 4.5, 1.7, 
    1.7, 5.5, 5.8, 4.5, 2.8, 1.1, 0.6, 0.5, 0.5, 0.8, 0.5, 0.1, 0.2, 0.2, 
    0.2, 0.9, 0.2, 0.1, 0.2, 0.5, 0.3, 1.1, 1, 1.1, 1.4, 0.9, 0.5, 0.3, 0, 
    0.1, 0.4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.3, 0.2, 0.9, 0.7, 2.6, 1.9, 
    0.3, 0.6, 0.5, 0.5, 0, 0, 0, 0, 0.2, 0, 0, 0.5, 1.5, 0.5, 0.5, 0, 0.3, 
    1.3, 1.2, 1.1, 0.8, 1.4, 0.8, 2.8, 0.8, 2.9, 2.2, 1.6, 1.3, 0.2, 0, 0.6, 
    0.1, 1, 0.9, 0.8, 0.9, 0, 1, 0.4, 0.6, 0.7, 0.6, 0.8, 0.7, 0.8, 0.1, 0.3, 
    0.9, 0.5, 0, 0.2, 1.4, 0.2, 0, 0, 0.7, 0, 0.1, 0.1, 0.4, 0.6, 0.1, 0.8, 
    1.7, 1.2, 1, 1.6, 2, 2.1, 2.1, 1.2, 1.8, 2.5, 0.1, 0.1, 0.2, 3.8, 3, 4.5, 
    5.5, 1.5, 1, 1.6, 0.1, 0.1, 6.1, 8.2, 6.6, 6.7, 2.4, 6, 8.7, 8.1, 6.7, 
    6.8, 6.2, 6.6, 4.7, 7.8, 8.2, 7, 4.5, 3.4, 3.6, 5.1, 2, 2.1, 2.4, 7, 6.5, 
    3.7, 2, 1.6, 1.5, 2, 0.7, 1.2, 0.8, 0.2, 1.8, 1.6, 0.6, 0.3, 0.1, 0.3, 
    0.7, 0, 0, 0, 0, 1.1, 1.4, 0.6, 0.1, 0.3, 0.7, 0.4, 0.1, 0, 0, 0, 0, 0.2, 
    0.2, 0.1, 0.7, 0.4, 0.5, 0.9, 0.6, 0, 1, 0.4, 0.7, 0.2, 0.8, 0.4, 0.6, 
    0.3, 0.6, 0.4, 0.3, 0.7, 0.2, 0.5, 0.3, 0.2, 0.4, 0.3, 1.3, 0.2, 0.1, 
    0.2, 0.3, 0, 1.2, 3, 3, 3.5, 1.2, 0.6, 0.6, 0.3, 1.5, 0.2, 2.2, 0.1, 0.6, 
    2.5, 3.3, 0.8, 2.2, 1.9, 2.8, 1.7, 0.8, 1.9, 2.5, 1.5, 0.9, 0.5, 0.5, 0, 
    1.5, 0.3, 1.1, 1.2, 0, 0, 1.2, 0.2, 0, 0.9, 0, 0.2, 0, 0.7, 1.2, 0.6, 
    0.2, 0, 1, 1.6, 0.6, 1.3, 1.9, 0.3, 0.5, 1, 1, 1.3, 0.5, 0.3, 2.1, 2.1, 
    3.8, 2.8, 6.6, 6.2, 5.5, 5.9, 4.9, 6.9, 6.1, 1.8, 6.2, 1.9, 4.8, 3.9, 
    4.6, 2.9, 0.8, 1.1, 3.8, 3.4, 4, 4.3, 2 ;

 relative_humidity = 0.95, 0.96, 0.96, 0.95, 0.95, 0.98, 0.99, 1, 0.98, 0.97, 
    0.98, 0.99, 0.98, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.88, 0.88, 
    0.88, 0.86, 0.83, 0.83, 0.83, 0.84, 0.86, 0.84, 0.82, 0.81, 0.86, 0.86, 
    0.85, 0.84, 0.83, 0.83, 0.82, 0.81, 0.82, 0.82, 0.82, 0.82, 0.9, 0.89, 
    0.88, 0.86, 0.85, 0.83, 0.83, 0.84, 0.84, 0.85, 0.83, 0.82, 0.86, 0.86, 
    0.87, 0.9, 0.87, 0.82, 0.83, 0.86, 0.84, 0.86, 0.86, 0.85, 0.9, 0.9, 
    0.92, 0.62, 0.62, 0.63, 0.67, 0.67, 0.62, 0.61, 0.66, 0.62, 0.63, 0.57, 
    0.57, 0.59, 0.6, 0.58, 0.63, 0.58, 0.56, 0.64, 0.6, 0.59, 0.65, 0.69, 
    0.76, 0.87, 0.89, 0.91, 0.89, 0.9, 0.8, 0.75, 0.69, 0.66, 0.65, 0.65, 
    0.64, 0.64, 0.6, 0.62, 0.64, 0.62, 0.6, 0.65, 0.65, 0.61, 0.63, 0.64, 
    0.66, 0.63, 0.66, 0.63, 0.6, 0.59, 0.58, 0.55, 0.54, 0.54, 0.56, 0.56, 
    0.55, 0.61, 0.62, 0.65, 0.65, 0.62, 0.61, 0.69, 0.73, 0.75, 0.73, 0.68, 
    0.67, 0.68, 0.65, 0.65, 0.65, 0.65, 0.59, 0.56, 0.56, 0.56, 0.57, 0.57, 
    0.51, 0.53, 0.53, 0.8, 0.81, 0.82, 0.82, 0.83, 0.85, 0.86, _, _, 0.64, 
    0.55, 0.56, 0.57, 0.57, 0.56, _, 0.56, 0.57, 0.59, 0.58, 0.57, 0.57, 
    0.56, 0.56, 0.58, 0.57, 0.53, 0.6, 0.56, 0.53, 0.55, 0.51, 0.46, 0.51, 
    0.47, 0.54, 0.98, 0.5, 0.55, 0.56, 0.57, 0.56, 0.6, 0.64, 0.81, 0.76, 
    0.57, 0.55, 0.58, 0.57, 0.55, 0.54, 0.6, 0.62, 0.63, 0.64, 0.65, 0.66, 
    0.66, 0.63, 0.8, 0.82, 0.61, 0.59, 0.6, 0.61, 0.61, 0.6, 0.63, 0.63, 
    0.59, 0.6, 0.62, 0.65, 0.62, 0.66, 0.66, 0.63, 0.66, 0.65, 0.62, 0.64, 
    0.65, 0.66, 0.66, 0.67, 0.67, 0.83, 0.72, 0.72, 0.65, 0.68, 0.65, 0.65, 
    0.67, 0.67, 0.64, 0.62, 0.63, 0.61, 0.58, 0.61, 0.64, 0.62, 0.58, 0.58, 
    0.58, 0.51, 0.53, 0.56, 0.54, 0.64, 0.63, 0.61, 0.59, 0.56, 0.55, 0.54, 
    0.52, 0.58, 0.57, 0.54, 0.49, 0.57, 0.56, 0.54, 0.52, 0.51, 0.54, 0.5, 
    0.51, 0.51, 0.5, 0.51, 0.53, 0.53, 0.55, 0.6, 0.55, 0.54, 0.58, 0.58, 
    0.56, 0.56, 0.61, 0.59, 0.59, 0.59, 0.54, 0.51, 0.51, 0.51, 0.51, 0.52, 
    0.53, 0.52, 0.54, 0.57, 0.58, 0.65, 0.68, 0.65, 0.68, 0.55, 0.63, 0.61, 
    0.61, 0.67, 0.64, 0.65, 0.64, 0.69, 0.73, 0.7, 0.65, 0.59, 0.58, 0.61, 
    0.69, 0.61, 0.82, 0.57, 0.55, 0.57, 0.56, 0.56, 0.57, 0.58, 0.64, 0.6, 
    0.6, 0.64, 0.62, 0.6, 0.63, 0.68, 0.68, 0.7, 0.66, 0.71, 0.69, 0.69, 
    0.71, 0.73, 0.73, 0.91, 0.68, 0.69, 0.69, 0.67, 0.67, 0.68, 0.69, 0.68, 
    0.65, 0.67, 0.69, 0.74, 0.73, 0.73, 0.71, 0.73, 0.77, 0.72, 0.81, 0.75, 
    0.99, 0.74, 0.77, 0.76, 0.76, 0.79, 0.78, 0.72, 0.75, 0.79, 0.77, 0.75, 
    0.74, 0.72, 0.72, 0.75, 0.72, 0.68, 0.73, 0.73, 0.73, 0.73, 0.71, 0.72, 
    0.67, 0.69, 0.69, 0.69, 0.7, 0.68, 0.72, 0.78, 0.77, 0.75, 0.78, 0.77, 
    0.74, 0.75, 0.7, 0.74, 0.73, 0.75, 0.8, 0.79, 0.77, 0.8, 0.81, 0.8, 0.81, 
    0.8, 0.8, 0.82, 0.84, 0.83, 0.81, 0.75, 0.73, 0.71, 0.75, 0.72, 0.69, 
    0.7, 0.73, 0.68, 0.71, 0.73, 0.77, 0.75, 0.73, 0.73, 0.77, 0.77, 0.99, 
    0.74, 0.73, 0.75, 0.76, 0.74, 0.74, 0.76, 0.72, 0.81, 0.78, 0.73, 0.77, 
    0.75, 0.81, 0.84, 0.81, 0.85, 0.86, 0.87, 0.88, 0.89, 0.88, 0.86, 0.9, 
    0.9, 0.91, 0.9, 0.92, 0.93, 0.93, 0.92, 0.9, 0.92, 0.91, 0.9, 0.76, 0.74, 
    0.69, 0.71, 0.72, 0.74, 0.68, 0.67, 0.67, 0.64, 0.67, 0.67, 0.69, 0.71, 
    0.69, 0.67, 0.65, 0.67, 0.73, 0.74, 0.77, 0.77, 0.76, 0.81, 0.85, 0.86, 
    0.88, 0.85, 0.84, 0.85, 0.81, 0.83, 0.83, 0.81, 0.82, 0.8, 0.94, 0.74, 
    0.76, 0.7, 0.79, 0.76, 0.73, 0.75, 0.72, 0.72, 0.63, 0.65, 0.7, 0.66, 
    0.74, 0.69, 0.64, 0.73, 0.73, 0.65, 0.66, 0.68, 0.69, 0.84, 0.85, 0.93, 
    0.9, 0.89, 0.92, 0.91, 0.92, 0.92, 0.93, 0.93, 0.96, 0.96, 0.96, 0.96, 
    0.94, 0.86, 0.87, 0.89, 0.87, 0.88, 0.87, 0.88, 0.88, 0.88, 0.91, 0.92, 
    0.87, 0.77, 0.78, 0.8, 0.77, 0.71, 0.71, 0.63, 0.61, 0.68, 0.74, 0.75, 
    0.72, 0.78, 0.78, 0.76, 0.76, 0.72, 0.66, 0.65, 0.73, 0.71, 0.71, 0.71, 
    0.72, 0.72, 0.8, 0.74, 0.78, 0.76, 0.72, 0.72, 0.73, 0.71, 0.77, 0.74, 
    0.69, 0.72, 0.71, 0.7, 0.68, 0.67, 0.69, 0.74, 0.75, 0.74, 0.72, 0.74, 
    0.71, 0.79, 0.74, 0.74, 0.74, 0.74, 0.73, 0.73, 0.73, 0.66, 0.7, 0.75, 
    0.72, 0.69, 0.71, 0.72, 0.66, 0.72, 0.69, 0.69, 0.73, 0.71, 0.68, 0.69, 
    0.71, 0.73, 0.68, 0.72, 0.71, 0.69, 0.72, 0.69, 0.69, 0.71, 0.68, 0.71, 
    0.7, 0.64, 0.66, 0.73, 0.68, 0.66, 0.75, 0.72, 0.72, 0.8, 0.72, 0.72, 
    0.73, 0.71, 0.74, 0.72, 0.76, 0.75, 0.78, 0.75, 0.74, 0.66, 0.66, 0.81, 
    0.81, 0.85, 0.78, 0.8, 0.74, 0.75, 0.75, 0.72, 0.68, 0.7, 0.74, 0.7, 
    0.75, 0.76, 0.8, 0.78, 0.8, 0.83, 0.85, 0.78, 0.84, 0.79, 0.79, 0.82, 
    0.9, 0.9, 0.92, 0.93, 0.76, 0.74, 0.78, 0.73, 0.73, 0.72, 0.6, 0.55, 
    0.51, 0.51, 0.52, 0.5, 0.48, 0.48, 0.46, 0.47, 0.46, 0.48, 0.46, 0.46, 
    0.44, 0.41, 0.47, 0.5, 0.5, 0.5, 0.48, 0.51, 0.53, 0.52, 0.51, 0.5, 0.57, 
    0.54, 0.55, 0.55, 0.6, 0.57, 0.6, 0.59, 0.55, 0.54, 0.54, 0.54, 0.55, 
    0.54, 0.54, 0.59, 0.57, 0.59, 0.72, 0.72, 0.77, 0.82, 0.84, 0.87, 0.89, 
    0.9, 0.91, 0.92, 0.91, 0.91, 0.81, 0.75, 0.65, 0.6, 0.58, 0.62, 0.54, 
    0.54, 0.55, 0.55, 0.47, 0.49, 0.5, 0.5, 0.58, 0.55, 0.84, 0.62, 0.6, 
    0.87, 0.63, 0.59, 0.67, 0.63, 0.7, 0.91, 0.67, 0.65, 0.67, 0.63, 0.64, 
    0.63, 0.63, 0.62, 0.62, 0.6, 0.65, 0.67, 0.74, 0.77, 0.82, 0.87, 0.88, 
    0.9, 0.9, 0.85, 0.84, 0.91, 0.88, 0.94, 0.94, 0.95, 0.95, 0.97, 0.97, 
    0.97, 0.85, 0.8, 0.78, 0.82, 0.83, 0.74, 0.73, 0.72, 0.72, 0.74, 0.71, 
    0.63, 0.8, 0.76, 0.74, 0.72, 0.62, 0.68, 0.63, 0.67, 0.68, 0.76, 0.75, 
    0.65, 0.56, 0.52, 0.51, 0.48, 0.51, 0.57, 0.56, 0.51, 0.52, 0.53, 0.55, 
    0.57, 0.58, 0.58, 0.58, 0.56, 0.58, 0.61, 0.65, 0.64, 0.67, 0.67, 0.62, 
    0.6, 0.68, 0.6, 0.61, 0.62, 0.7, 0.68, 0.66, 0.64, 0.64, 0.62, 0.62, 
    0.67, 0.67, 0.68, 0.66, 0.65, 0.66, 0.67, 0.64, 0.67, 0.59, 0.52, 0.65, 
    0.62, 0.52, 0.45, 0.45, 0.4, 0.34, 0.44, 0.49, 0.45, 0.39, 0.38, 0.42, 
    0.46, 0.54, 0.46, 0.35, 0.41, 0.45, 0.42, 0.5, 0.5, 0.5, 0.49, 0.48, 
    0.55, 0.66, 0.66, 0.63, 0.69, 0.65, 0.58, 0.55, 0.53, 0.53, 0.48, 0.49, 
    0.51, 0.53, 0.51, 0.46, 0.45, 0.47, 0.46, 0.48, 0.51, 0.45, 0.45, 0.44, 
    0.45, 0.4, 0.38, 0.36, 0.4, 0.41, 0.43, 0.45, 0.45, 0.43, 0.49, 0.5, 
    0.49, 0.49, 0.49, 0.47, 0.49, 0.51, 0.54, 0.57, 0.61, 0.69, 0.76, 0.76, 
    0.7, 0.7, 0.65, 0.69, 0.68, 0.66, 0.66, 0.65, 0.65, 0.64, 0.66, 0.64, 
    0.62, 0.6, 0.63, 0.7, 0.72, 0.72, 0.72, 0.72, 0.65, 0.67, 0.66, 0.61, 
    0.62, 0.62, 0.63, 0.59, 0.58, 0.55, 0.53, 0.46, 0.52, 0.47, 0.48, 0.52, 
    0.48, 0.49, 0.46, 0.49, 0.49, 0.58, 0.64, 0.69, 0.83, 0.86, 0.86, 0.85, 
    0.86, 0.85, 0.78, 0.82, 0.81, 0.74, 0.85, 0.89, 0.79, 0.67, 0.58, 0.66, 
    0.57, 0.59, 0.57, 0.61, 0.68, 0.62, 0.6, 0.65, 0.59, 0.55, 0.55, 0.8, 
    0.65, 0.76, 0.86, 0.88, 0.83, 0.79, 0.77, 0.78, 0.74, 0.77, 0.74, 0.74, 
    0.74, 0.74, 0.74, 0.81, 0.84, 0.77, 0.68, 0.71, 0.65, 0.74, 0.74, 0.79, 
    0.78, 0.77, 0.78, 0.8, 0.81, _, _, 0.8, 0.79, 0.81, 0.8, 0.78, 0.81, 
    0.84, 0.89, 0.86, 0.84, 0.83, 0.75, 0.76, 0.78, 0.78, 0.74, 0.75, 0.81, 
    0.77, 0.78, 0.79, 0.76, 0.74, 0.71, 0.68, 0.69, 0.66, 0.68, 0.7, 0.64, 
    0.63, 0.66, 0.68, 0.64, 0.65, 0.64, 0.62, 0.62, 0.66, 0.66, 0.64, 0.62, 
    0.61, 0.63, 0.66, 0.6, 0.65, 0.7, 0.76, 0.74, 0.79, 0.77, 0.67, 0.69, 
    0.66, 0.63, 0.65, 0.66, 0.64, 0.62, 0.66, 0.63, 0.6, 0.59, 0.65, 0.67, 
    0.66, 0.72, 0.71, 0.66, 0.62, 0.7, 0.82, 0.67, 0.75, 0.94, 0.96, 0.96, 
    0.94, 0.92, 0.91, 0.96, 0.97, 0.95, 0.93, 0.74, 0.64, 0.65, 0.64, 0.67, 
    0.65, 0.62, 0.64, 0.64, 0.66, 0.57, 0.59, 0.56, 0.82, 0.62, 0.69, 0.68, 
    0.66, 0.71, 0.67, 0.66, 0.63, 0.66, 0.66, 0.63, 0.67, 0.74, 0.69, 0.66, 
    0.65, 0.64, 0.72, 0.73, 0.74, 0.65, 0.65, 0.65, 0.68, 0.66, 0.72, 0.76, 
    0.77, 0.68, 0.77, 0.78, 0.78, 0.72, 0.7, 0.71, 0.61, 0.62, 0.65, 0.6, 
    0.68, 0.73, 0.9, 0.88, 0.8, 0.76, 0.73, 0.8, 0.76, 0.9, 0.91, 0.9, 0.88, 
    0.86, 0.9, 0.92, 0.95, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.86, 0.85, 0.79, 0.86, 0.8, 0.8, 0.87, 0.76, 0.76, 0.76, 0.82, 0.83, 
    0.76, 0.79, 0.66, 0.69, 0.66, 0.69, 0.72, 0.7, 0.66, 0.68, 0.64, 0.61, 
    0.64, 0.68, 0.67, 0.65, 0.69, 0.63, 0.71, 0.69, 0.69, 0.6, 0.63, 0.63, 
    0.64, 0.65, 0.67, 0.67, 0.64, 0.65, 0.64, 0.68, 0.7, 0.65, 0.65, 0.67, 
    0.66, 0.69, 0.68, 0.68, 0.68, 0.67, 0.66, 0.69, 0.7, 0.72, 0.74, 0.71, 
    0.7, 0.74, 0.7, 0.73, 0.76, 0.76, 0.77, 0.77, 0.77, 0.81, 0.8, 0.79, 
    0.83, 0.83, 0.85, 0.76, 0.76, 0.72, 0.67, 0.71, 0.75, 0.79, 0.88, 0.93, 
    0.83, 0.82, 0.81, 0.86, 0.85, 0.78, 0.76, 0.84, 0.86, 0.85, 0.83, 0.84, 
    0.8, 0.76, 0.65, 0.58, 0.51, 0.62, 0.61, 0.53, 0.58, 0.58, 0.56, 0.55, 
    0.63, 0.63, 0.62, 0.64, 0.69, 0.73, 0.75, 0.7, 0.57, 0.55, 0.58, 0.62, 
    0.57, 0.58, 0.64, 0.69, 0.67, 0.67, 0.66, 0.6, 0.65, 0.61, 0.67, 0.67, 
    0.58, 0.59, 0.55, 0.53, 0.52, 0.5, 0.52, 0.53, 0.51, 0.49, 0.44, 0.45, 
    0.48, 0.48, 0.46, 0.5, 0.45, 0.48, 0.5, 0.5, 0.5, 0.55, 0.55, 0.55, 0.61, 
    0.6, 0.64, 0.62, 0.63, 0.61, 0.63, 0.63, 0.62, 0.61, 0.64, 0.66, 0.63, 
    0.68, 0.69, 0.65, 0.63, 0.66, 0.62, 0.67, 0.65, 0.66, 0.67, 0.67, 0.67, 
    0.65, 0.69, 0.67, 0.64, 0.6, 0.63, 0.65, 0.62, 0.62, 0.63, 0.62, 0.63, 
    0.65, 0.65, 0.59, 0.61, 0.63, 0.58, 0.62, 0.61, 0.61, 0.64, 0.58, 0.62, 
    0.63, 0.59, 0.64, 0.55, 0.59, 0.55, 0.57, 0.61, 0.65, 0.67, 0.61, 0.79, 
    0.88, 0.86, 0.88, 0.87, 0.87, 0.83, 0.73, 0.72, 0.75, 0.82, 0.87, 0.91, 
    0.9, 0.75, 0.7, 0.67, 0.69, 0.65, 0.67, 0.61, 0.58, 0.59, 0.7, 0.7, 0.69, 
    0.6, 0.66, 0.67, 0.69, 0.59, 0.59, 0.6, 0.61, 0.62, 0.62, 0.56, 0.53, 
    0.55, 0.51, 0.62, 0.65, 0.58, 0.55, 0.49, 0.51, 0.5, 0.51, 0.52, 0.52, 
    0.52, 0.48, 0.49, 0.5, 0.55, 0.57, 0.6, 0.59, 0.66, 0.66, 0.63, 0.64, 
    0.6, 0.58, 0.57, 0.57, 0.54, 0.57, 0.59, 0.65, 0.72, 0.74, 0.77, 0.79, 
    0.71, 0.68, 0.71, 0.68, 0.71, 0.73, 0.73, 0.74, 0.74, 0.76, 0.75, 0.75, 
    0.76, 0.78, 0.78, 0.78, 0.73, 0.76, 0.86, 0.86, 0.88, 0.9, 0.89, 0.87, 
    0.89, 0.88, 0.9, 0.92, 0.95, 0.96, 0.96, 0.96, 0.95, 0.92, 0.91, 0.94, 
    0.92, 0.9, 0.76, 0.69, 0.66, 0.69, 0.65, 0.63, 0.77, 0.57, 0.51, 0.5, 
    0.51, 0.51, 0.53, 0.55, 0.6, 0.58, 0.62, 0.65, 0.65, 0.53, 0.51, 0.41, 
    0.38, 0.47, 0.48, 0.51, 0.48, 0.54, 0.5, 0.51, 0.57, 0.55, 0.45, 0.44, 
    0.44, 0.44, 0.47, 0.49, 0.57, 0.49, 0.53, 0.51, 0.52, 0.45, 0.51, 0.51, 
    0.48, 0.57, 0.53, 0.48, 0.42, 0.45, 0.5, 0.45, 0.42, 0.41, 0.51, 0.5, 
    0.47, 0.5, 0.5, 0.51, 0.51, 0.49, 0.49, 0.53, 0.57, 0.46, 0.44, 0.45, 
    0.46, 0.46, 0.47, 0.49, 0.47, 0.45, 0.45, 0.48, 0.55, 0.57, 0.55, 0.54, 
    0.56, 0.56, 0.55, 0.56, 0.57, 0.53, 0.54, 0.53, 0.54, 0.6, 0.54, 0.6, 
    0.53, 0.5, 0.55, 0.56, 0.59, 0.59, 0.6, 0.63, 0.67, 0.63, 0.64, 0.66, 
    0.62, 0.58, 0.63, 0.53, 0.57, 0.61, 0.57, 0.57, 0.59, 0.57, 0.58, 0.59, 
    0.6, 0.6, 0.62, 0.63, 0.61, 0.61, 0.58, 0.57, 0.56, 0.54, 0.56, 0.58, 
    0.55, 0.57, 0.57, 0.58, 0.57, 0.56, 0.6, 0.58, 0.6, 0.6, 0.59, 0.59, 
    0.61, 0.58, 0.58, 0.57, 0.59, 0.61, 0.62, 0.64, 0.63, 0.69, 0.68, 0.64, 
    0.69, 0.69, 0.7, 0.71, 0.72, 0.73, 0.76, 0.73, 0.75, 0.76, 0.71, 0.71, 
    0.71, 0.76, 0.73, 0.78, 0.73, 0.76, 0.73, 0.74, 0.78, 0.74, 0.69, 0.69, 
    0.77, 0.75, 0.71, 0.77, 0.65, 0.78, 0.74, 0.72, 0.74, 0.75, 0.81, 0.76, 
    0.77, 0.78, 0.79, 0.77, 0.77, 0.78, 0.76, 0.78, 0.8, 0.77, 0.8, 0.84, 
    0.85, 0.8, 0.8, 0.8, 0.79, 0.79, 0.78, 0.8, 0.78, 0.78, 0.79, 0.8, 0.79, 
    0.77, 0.76, 0.75, 0.81, 0.78, 0.79, 0.81, 0.78, 0.76, 0.79, 0.8, 0.79, 
    0.78, 0.76, 0.78, 0.79, 0.8, 0.77, 0.74, 0.8, 0.69, 0.69, 0.68, 0.68, 
    0.71, 0.68, 0.62, 0.58, 0.55, 0.6, 0.57, 0.55, 0.53, 0.56, 0.6, 0.55, 
    0.55, 0.53, 0.52, 0.53, 0.51, 0.46, 0.48, 0.52, 0.55, 0.57, 0.53, 0.57, 
    0.62, 0.48, 0.58, 0.46, 0.52, 0.48, 0.48, 0.48, 0.54, 0.47, 0.47, 0.49, 
    0.47, 0.47, 0.45, 0.47, 0.53, 0.45, 0.47, 0.46, 0.44, 0.46, 0.47, 0.44, 
    0.53, 0.58, 0.5, 0.53, 0.54, 0.52, 0.52, 0.51, 0.48, 0.54, 0.52, 0.58, 
    0.46, 0.5, 0.56, 0.49, 0.49, 0.45, 0.51, 0.52, 0.59, 0.56, 0.6, 0.58, 
    0.57, 0.65, 0.65, 0.61, 0.66, 0.65, 0.67, 0.68, 0.68, 0.71, 0.72, 0.7, 
    0.77, 0.72, 0.75, 0.71, 0.67, 0.76, 0.76, 0.71, 0.71, 0.73, 0.77, 0.76, 
    0.73, 0.8, 0.78, 0.81, 0.75, 0.77, 0.76, 0.74, 0.74, 0.74, 0.73, 0.74, 
    0.72, 0.73, 0.71, 0.73, 0.7, 0.74, 0.73, 0.72, 0.68, 0.67, 0.74, 0.7, 
    0.71, 0.73, 0.72, 0.68, 0.64, 0.64, 0.65, 0.72, 0.73, 0.69, 0.61, 0.59, 
    0.65, 0.69, 0.65, 0.63, 0.61, 0.58, 0.57, 0.64, 0.63, 0.6, 0.6, 0.66, 
    0.65, 0.61, 0.67, 0.64, 0.64, 0.69, 0.67, 0.67, 0.64, 0.68, 0.72, 0.68, 
    0.69, 0.77, 0.63, 0.67, 0.7, 0.7, 0.66, 0.77, 0.72, 0.68, 0.7, 0.68, 
    0.71, 0.74, 0.75, 0.7, 0.75, 0.76, 0.72, 0.74, 0.77, 0.71, 0.76, 0.73, 
    0.76, 0.75, 0.77, 0.72, 0.73, 0.73, 0.73, 0.73, 0.74, 0.73, 0.77, 0.75, 
    0.72, 0.7, 0.71, 0.73, 0.78, 0.72, 0.74, 0.77, 0.81, 0.78, 0.74, 0.71, 
    0.77, 0.77, 0.79, 0.76, 0.76, 0.77, 0.89, 0.92, 0.93, 0.92, 0.9, 0.92, 
    0.92, 0.95, 0.93, 0.91, 0.93, 0.91, 0.9, 0.91, 0.89, 0.92, 0.94, 0.92, 
    0.92, 0.92, 0.94, 0.96, 0.94, 0.89, 0.9, 0.9, 0.9, 0.9, 0.94, 0.95, 0.96, 
    0.96, 0.97, 0.98, 0.99, 0.98, 0.99, 0.81, 0.79, 0.74, 0.72, 0.74, 0.74, 
    0.73, 0.75, 0.79, 0.77, 0.77, 0.76, 0.88, 0.83, 0.82, 0.9, 0.95, 0.94, 
    0.86, 0.87, 0.72, 0.69, 0.65, 0.59, 0.64, 0.66, 0.68, 0.73, 0.74, 0.74, 
    0.73, 0.75, 0.71, 0.7, 0.73, 0.73, 0.75, 0.74, 0.76, 0.78, 0.76, 0.79, 
    0.83, 0.86, 0.85, 0.84, 0.84, 0.87, 0.86, 0.8, 0.8, 0.82, 0.83, 0.81, 
    0.8, 0.84, 0.85, 0.8, 0.77, 0.74, 0.74, 0.79, 0.79, 0.81, 0.81, 0.81, 
    0.76, 0.82, 0.79, 0.81, 0.84, 0.78, 0.79, 0.76, 0.74, 0.77, 0.74, 0.75, 
    0.76, 0.82, 0.81, 0.84, 0.83, 0.81, 0.79, 0.83, 0.85, 0.89, 0.88, 0.84, 
    0.9, 0.91, 0.91, 0.89, 0.88, 0.9, 0.91, 0.9, 0.87, 0.87, 0.88, 0.89, 
    0.82, 0.87, 0.88, 0.94, 0.97, 0.96, 0.97, 0.96, 0.96, 0.96, 0.97, 0.97, 
    0.97, 0.95, 0.93, 0.89, 0.82, 0.82, 0.84, 0.88, 0.84, 0.85, 0.82, 0.79, 
    0.77, 0.7, 0.66, 0.64, 0.61, 0.56, 0.51, 0.47, 0.56, 0.57, 0.57, 0.61, 
    0.63, 0.62, 0.63, 0.62, 0.63, 0.62, 0.62, 0.66, 0.66, 0.66, 0.67, 0.65, 
    0.65, 0.66, 0.64, 0.7, 0.75, 0.75, 0.76, 0.73, 0.67, 0.68, 0.63, 0.65, 
    0.62, 0.65, 0.66, 0.73, 0.73, 0.71, 0.72, 0.75, 0.75, 0.71, 0.77, 0.79, 
    0.8, 0.82, 0.83, 0.81, 0.81, 0.84, 0.82, 0.82, 0.84, 0.83, 0.86, 0.83, 
    0.82, 0.79, 0.79, 0.76, 0.73, 0.72, 0.7, 0.67, 0.62, 0.57, 0.55, 0.55, 
    0.54, 0.53, 0.53, 0.53, 0.53, 0.52, 0.54, 0.56, 0.6, 0.59, 0.61, 0.59, 
    0.65, 0.64, 0.65, 0.66, 0.67, 0.64, 0.69, 0.64, 0.7, 0.71, 0.65, 0.67, 
    0.64, 0.63, 0.62, 0.61, 0.6, 0.59, 0.62, 0.62, 0.62, 0.67, 0.68, 0.65, 
    0.65, 0.67, 0.65, 0.63, 0.72, 0.78, 0.72, 0.67, 0.68, 0.69, 0.67, 0.64, 
    0.6, 0.64, 0.57, 0.55, 0.52, 0.52, 0.54, 0.57, 0.53, 0.5, 0.49, 0.51, 
    0.51, 0.38, 0.37, 0.35, 0.35, 0.41, 0.49, 0.43, 0.43, 0.46, 0.51, 0.54, 
    0.56, 0.58, 0.61, 0.56, 0.61, 0.57, 0.56, 0.55, 0.59, 0.56, 0.57, 0.58, 
    0.56, 0.57, 0.6, 0.57, 0.55, 0.58, 0.52, 0.51, 0.5, 0.45, 0.49, 0.47, 
    0.45, 0.45, 0.44, 0.45, 0.57, 0.52, 0.51, 0.49, 0.57, 0.59, 0.59, 0.56, 
    0.52, 0.47, 0.49, 0.51, 0.52, 0.47, 0.43, 0.45, 0.48, 0.47, 0.49, 0.52, 
    0.54, 0.52, 0.53, 0.54, 0.55, 0.56, 0.55, 0.62, 0.58, 0.58, 0.58, 0.59, 
    0.57, 0.6, 0.55, 0.54, 0.51, 0.5, 0.54, 0.52, 0.49, 0.51, 0.47, 0.49, 
    0.54, 0.49, 0.5, 0.52, 0.52, 0.48, 0.55, 0.51, 0.52, 0.52, 0.54, 0.56, 
    0.57, 0.53, 0.51, 0.51, 0.57, 0.5, 0.5, 0.46, 0.46, 0.42, 0.44, 0.44, 
    0.39, 0.5, 0.48, 0.48, 0.5, 0.5, 0.51, 0.46, 0.47, 0.49, 0.51, 0.49, 
    0.51, 0.52, 0.53, 0.54, 0.52, 0.55, 0.5, 0.5, 0.5, 0.48, 0.51, 0.51, 
    0.52, 0.53, 0.52, 0.5, 0.5, 0.51, 0.56, 0.56, 0.59, 0.61, 0.58, 0.57, 
    0.56, 0.55, 0.52, 0.52, 0.49, 0.48, 0.49, 0.43, 0.41, 0.44, 0.41, 0.39, 
    0.37, 0.43, 0.37, 0.35, 0.38, 0.39, 0.41, 0.47, 0.48, 0.53, 0.53, 0.54, 
    0.52, 0.45, 0.47, 0.52, 0.45, 0.42, 0.43, 0.51, 0.49, 0.52, 0.54, 0.49, 
    0.46, 0.44, 0.47, 0.46, 0.49, 0.45, 0.45, 0.51, 0.52, 0.52, 0.53, 0.52, 
    0.44, 0.45, 0.47, 0.5, 0.5, 0.55, 0.47, 0.48, 0.49, 0.49, 0.5, 0.54, 
    0.59, 0.66, 0.63, 0.71, 0.61, 0.6, 0.66, 0.68, 0.7, 0.65, 0.72, 0.79, 
    0.83, 0.81, 0.81, 0.82, 0.82, 0.8, 0.81, 0.83, 0.84, 0.82, 0.83, 0.85, 
    0.84, 0.79, 0.77, 0.82, 0.8, 0.8, 0.8, 0.8, 0.8, 0.83, 0.76, 0.65, 0.66, 
    0.66, 0.58, 0.57, 0.53, 0.59, 0.62, 0.61, 0.63, 0.64, 0.62, 0.62, 0.62, 
    0.6, 0.62, 0.58, 0.59, 0.53, 0.55, 0.61, 0.6, 0.5, 0.47, 0.49, 0.46, 
    0.44, 0.42, 0.41, 0.43, 0.41, 0.48, 0.73, 0.51, 0.53, 0.55, 0.51, 0.55, 
    0.52, 0.55, 0.53, 0.51, 0.48, 0.47, 0.54, 0.55, 0.59, 0.65, 0.73, 0.63, 
    0.59, 0.58, 0.65, 0.51, 0.56, 0.47, 0.44, 0.45, 0.41, 0.47, 0.53, 0.57, 
    0.46, 0.46, 0.52, 0.51, 0.47, 0.46, 0.61, 0.62, 0.58, 0.54, 0.48, 0.44, 
    0.5, 0.45, 0.41, 0.44, 0.4, 0.4, 0.39, 0.39, 0.41, 0.43, 0.42, 0.44, 
    0.49, 0.5, 0.47, 0.47, 0.47, 0.49, 0.52, 0.49, 0.54, 0.55, 0.54, 0.57, 
    0.59, 0.6, 0.67, 0.65, 0.65, 0.66, 0.66, 0.68, 0.7, 0.66, 0.74, 0.75, 
    0.76, 0.77, 0.72, 0.62, 0.6, 0.71, 0.72, 0.72, 0.69, 0.67, 0.67, 0.66, 
    0.67, 0.64, 0.64, 0.64, 0.64, 0.64, 0.65, 0.65, 0.68, 0.66, 0.63, 0.6, 
    0.62, 0.62, 0.59, 0.57, 0.55, 0.63, 0.66, 0.63, 0.63, 0.67, 0.63, 0.66, 
    0.61, 0.63, 0.66, 0.66, 0.69, 0.71, 0.71, 0.68, 0.68, 0.69, 0.63, 0.64, 
    0.63, 0.62, 0.62, 0.63, 0.64, 0.63, 0.63, 0.65, 0.62, 0.54, 0.45, 0.51, 
    0.49, 0.48, 0.43, 0.46, 0.45, 0.51, 0.52, 0.52, 0.53, 0.55, 0.58, 0.59, 
    0.54, 0.55, 0.55, 0.57, 0.63, 0.68, 0.7, 0.73, 0.74, 0.73, 0.73, 0.75, 
    0.71, 0.7, 0.72, 0.63, 0.7, 0.65, 0.66, 0.68, 0.69, 0.7, 0.72, 0.72, 
    0.77, 0.78, 0.81, 0.58, 0.58, 0.62, 0.63, 0.66, 0.59, 0.59, 0.6, 0.61, 
    0.65, 0.58, 0.58, 0.58, 0.59, 0.53, 0.5, 0.48, 0.51, 0.49, 0.51, 0.53, 
    0.55, 0.56, 0.5, 0.49, 0.53, 0.56, 0.59, 0.57, 0.59, 0.6, 0.6, 0.62, 
    0.63, 0.64, 0.67, 0.69, 0.7, 0.71, 0.73, 0.78, 0.82, 0.78, 0.79, 0.77, 
    0.76, 0.78, 0.74, 0.71, 0.71, 0.74, 0.75, 0.75, 0.79, 0.8, 0.81, 0.78, 
    0.73, 0.65, 0.64, 0.59, 0.52, 0.53, 0.5, 0.54, 0.57, 0.63, 0.69, 0.73, 
    0.73, 0.7, 0.71, 0.7, 0.69, 0.68, 0.74, 0.72, 0.71, 0.76, 0.78, 0.75, 
    0.78, 0.73, 0.74, 0.68, 0.68, 0.63, 0.62, 0.62, 0.65, 0.58, 0.56, 0.54, 
    0.55, 0.55, 0.53, 0.62, 0.73, 0.71, 0.68, 0.67, 0.66, 0.64, 0.62, 0.62, 
    0.58, 0.62, 0.6, 0.61, 0.59, 0.58, 0.6, 0.63, 0.63, 0.6, 0.61, 0.64, 
    0.65, 0.62, 0.69, 0.69, 0.69, 0.67, 0.69, 0.7, 0.71, 0.75, 0.68, 0.67, 
    0.69, 0.68, 0.69, 0.65, 0.61, 0.68, 0.65, 0.53, 0.64, 0.64, 0.62, 0.57, 
    0.62, 0.58, 0.54, 0.49, 0.51, 0.56, 0.59, 0.56, 0.6, 0.56, 0.57, 0.6, 
    0.49, 0.53, 0.53, 0.55, 0.59, 0.51, 0.51, 0.53, 0.6, 0.54, 0.7, 0.6, 
    0.57, 0.56, 0.51, 0.56, 0.44, 0.57, 0.51, 0.48, 0.5, 0.5, 0.46, 0.53, 
    0.48, 0.46, 0.48, 0.57, 0.55, 0.54, 0.53, 0.52, 0.56, 0.51, 0.44, 0.54, 
    0.52, 0.51, 0.47, 0.44, 0.44, 0.47, 0.53, 0.5, 0.56, 0.55, 0.59, 0.56, 
    0.53, 0.58, 0.55, 0.58, 0.57, 0.59, 0.58, 0.76, 0.62, 0.67, 0.55, 0.55, 
    0.55, 0.54, 0.49, 0.52, 0.48, 0.52, 0.5, 0.58, 0.61, 0.54, 0.59, 0.53, 
    0.55, 0.6, 0.59, 0.64, 0.62, 0.58, 0.58, 0.59, 0.62, 0.62, 0.57, 0.58, 
    0.54, 0.51, 0.49, 0.55, 0.51, 0.46, 0.57, 0.57, 0.55, 0.54, 0.58, 0.62, 
    0.64, 0.58, 0.61, 0.63, 0.62, 0.62, 0.63, 0.64, 0.65, 0.6, 0.67, 0.63, 
    0.59, 0.59, 0.61, 0.61, 0.48, 0.58, 0.6, 0.67, 0.7, 0.64, 0.74, 0.72, 
    0.71, 0.77, 0.79, 0.78, 0.83, 0.8, 0.84, 0.82, 0.57, 0.6, 0.57, 0.62, 
    0.5, 0.51, 0.48, 0.5, 0.53, 0.5, 0.49, 0.47, 0.55, 0.52, 0.51, 0.53, 
    0.56, 0.53, 0.55, 0.57, 0.61, 0.57, 0.55, 0.54, 0.54, 0.51, 0.53, 0.57, 
    0.55, 0.53, 0.52, 0.53, 0.51, 0.49, 0.53, 0.48, 0.49, 0.52, 0.56, 0.55, 
    0.58, 0.57, 0.6, 0.62, 0.65, 0.65, 0.74, 0.65, 0.65, 0.65, 0.62, 0.58, 
    0.58, 0.58, 0.5, 0.52, 0.5, 0.46, 0.46, 0.49, 0.52, 0.53, 0.57, 0.63, 
    0.61, 0.6, 0.56, 0.57, 0.58, 0.61, 0.62, 0.61, 0.62, 0.63, 0.62, 0.58, 
    0.54, 0.51, 0.52, 0.52, 0.45, 0.49, 0.46, 0.52, 0.5, 0.55, 0.55, 0.58, 
    0.56, 0.57, 0.6, 0.6, 0.6, 0.61, 0.61, 0.61, 0.58, 0.58, 0.57, 0.8, 0.81, 
    0.75, 0.61, 0.53, 0.52, 0.53, 0.48, 0.5, 0.48, 0.5, 0.52, 0.5, 0.52, 
    0.52, 0.54, 0.59, 0.6, 0.61, 0.59, 0.57, 0.59, 0.62, 0.68, 0.72, 0.71, 
    0.8, 0.69, 0.68, 0.67, 0.63, 0.6, 0.57, 0.6, 0.56, 0.54, 0.56, 0.53, 
    0.63, 0.64, 0.63, 0.66, 0.64, 0.66, 0.67, 0.65, 0.61, 0.63, 0.63, 0.61, 
    0.56, 0.57, 0.6, 0.61, 0.64, 0.58, 0.68, 0.64, 0.65, 0.65, 0.66, 0.68, 
    0.69, 0.72, 0.68, 0.59, 0.66, 0.71, 0.76, 0.74, 0.64, 0.63, 0.59, 0.62, 
    0.55, 0.53, 0.54, 0.52, 0.48, 0.5, 0.49, 0.58, 0.58, 0.63, 0.66, 0.73, 
    0.73, 0.74, 0.73, 0.71, 0.66, 0.64, 0.63, 0.64, 0.66, 0.66, 0.62, 0.56, 
    0.57, 0.6, 0.57, 0.58, 0.58, 0.61, 0.64, 0.62, 0.62, 0.68, 0.75, 0.72, 
    0.78, 0.74, 0.73, 0.73, 0.73, 0.75, 0.79, 0.75, 0.74, 0.66, 0.67, 0.65, 
    0.61, 0.53, 0.56, 0.57, 0.5, 0.54, 0.57, 0.63, 0.57, 0.6, 0.64, 0.66, 
    0.64, 0.63, 0.66, 0.68, 0.7, 0.66, 0.64, 0.65, 0.63, 0.6, 0.59, 0.64, 
    0.48, 0.54, 0.5, 0.52, 0.53, 0.51, 0.55, 0.65, 0.65, 0.64, 0.68, 0.65, 
    0.69, 0.73, 0.64, 0.63, 0.78, 0.65, 0.68, 0.74, 0.69, 0.67, 0.59, 0.57, 
    0.5, 0.53, 0.56, 0.48, 0.51, 0.57, 0.56, 0.51, 0.61, 0.59, 0.65, 0.65, 
    0.64, 0.7, 0.68, 0.7, 0.72, 0.71, 0.73, 0.69, 0.69, 0.7, 0.69, 0.69, 
    0.67, 0.62, 0.57, 0.56, 0.59, 0.6, 0.68, 0.58, 0.57, 0.56, 0.52, 0.52, 
    0.56, 0.52, 0.54, 0.52, 0.53, 0.54, 0.54, 0.52, 0.55, 0.48, 0.41, 0.43, 
    0.51, 0.58, 0.58, 0.53, 0.52, 0.52, 0.55, 0.59, 0.57, 0.61, 0.57, 0.53, 
    0.55, 0.55, 0.56, 0.57, 0.58, 0.58, 0.57, 0.58, 0.52, 0.48, 0.49, 0.48, 
    0.45, 0.48, 0.48, 0.46, 0.45, 0.55, 0.5, 0.5, 0.55, 0.6, 0.57, 0.6, 0.59, 
    0.59, 0.52, 0.53, 0.55, 0.5, 0.57, 0.55, 0.54, 0.54, 0.5, 0.48, 0.45, 
    0.42, 0.39, 0.44, 0.42, 0.43, 0.44, 0.46, 0.48, 0.49, 0.6, 0.63, 0.68, 
    0.63, 0.53, 0.48, 0.47, 0.46, 0.46, 0.53, 0.57, 0.58, 0.56, 0.49, 0.48, 
    0.48, 0.46, 0.49, 0.51, 0.5, 0.59, 0.57, 0.59, 0.53, 0.49, 0.5, 0.51, 
    0.49, 0.53, 0.55, 0.56, 0.55, 0.56, 0.57, 0.58, 0.56, 0.51, 0.47, 0.47, 
    0.42, 0.51, 0.52, 0.55, 0.54, 0.54, 0.54, 0.54, 0.56, 0.56, 0.61, 0.61, 
    0.63, 0.61, 0.61, 0.62, 0.64, 0.67, 0.67, 0.65, 0.68, 0.58, 0.61, 0.56, 
    0.54, 0.47, 0.5, 0.55, 0.49, 0.5, 0.51, 0.58, 0.57, 0.61, 0.61, 0.62, 
    0.62, 0.6, 0.51, 0.54, 0.58, 0.58, 0.62, 0.6, 0.6, 0.6, 0.57, 0.53, 0.55, 
    0.53, 0.51, 0.52, 0.51, 0.57, 0.55, 0.58, 0.61, 0.65, 0.69, 0.7, 0.71, 
    0.69, 0.69, 0.73, 0.73, 0.71, 0.73, 0.71, 0.68, 0.57, 0.53, 0.53, 0.49, 
    0.48, 0.57, 0.55, 0.55, 0.6, 0.56, 0.6, 0.63, 0.66, 0.74, 0.74, 0.73, 
    0.73, 0.75, 0.77, 0.72, 0.75, 0.72, 0.7, 0.73, 0.63, 0.61, 0.48, 0.54, 
    0.53, 0.51, 0.55, 0.62, 0.5, 0.59, 0.6, 0.62, 0.67, 0.73, 0.75, 0.74, 
    0.73, 0.73, 0.77, 0.77, 0.76, 0.76, 0.75, 0.68, 0.63, 0.57, 0.58, 0.56, 
    0.62, 0.6, 0.72, 0.7, 0.61, 0.68, 0.65, 0.69, 0.71, 0.67, 0.72, 0.67, 
    0.64, 0.63, 0.64, 0.67, 0.69, 0.65, 0.6, 0.65, 0.56, 0.52, 0.51, 0.51, 
    0.5, 0.47, 0.52, 0.54, 0.51, 0.5, 0.57, 0.53, 0.52, 0.57, 0.62, 0.59, 
    0.57, 0.62, 0.62, 0.57, 0.58, 0.61, 0.55, 0.52, 0.48, 0.45, 0.52, 0.51, 
    0.53, 0.45, 0.5, 0.45, 0.5, 0.43, 0.49, 0.48, 0.5, 0.49, 0.53, 0.49, 
    0.56, 0.57, 0.61, 0.56, 0.56, 0.54, 0.52, 0.5, 0.41, 0.42, 0.41, 0.4, 
    0.4, 0.4, 0.38, 0.44, 0.45, 0.46, 0.49, 0.52, 0.55, 0.56, 0.58, 0.57, 
    0.57, 0.57, 0.59, 0.58, 0.58, 0.58, 0.56, 0.56, 0.49, 0.49, 0.46, 0.45, 
    0.49, 0.49, 0.49, 0.48, 0.55, 0.53, 0.55, 0.57, 0.6, 0.64, 0.67, 0.66, 
    0.64, 0.66, 0.65, 0.68, 0.6, 0.59, 0.53, 0.55, 0.48, 0.45, 0.36, 0.43, 
    0.34, 0.44, 0.49, 0.51, 0.55, 0.57, 0.53, 0.48, 0.48, 0.8, 0.55, 0.57, 
    0.58, 0.57, 0.57, 0.56, 0.57, 0.58, 0.56, 0.49, 0.5, 0.43, 0.46, 0.46, 
    0.41, 0.57, 0.45, 0.61, 0.62, 0.59, 0.64, 0.69, 0.72, 0.69, 0.73, 0.78, 
    0.81, 0.8, 0.83, 0.82, 0.82, 0.82, 0.79, 0.78, 0.64, 0.58, 0.5, 0.55, 
    0.48, 0.58, 0.6, 0.58, 0.66, 0.68, 0.62, 0.57, 0.62, 0.64, 0.61, 0.69, 
    0.65, 0.64, 0.63, 0.64, 0.71, 0.65, 0.65, 0.66, 0.63, 0.61, 0.56, 0.46, 
    0.44, 0.38, 0.34, 0.46, 0.5, 0.48, 0.56, 0.58, 0.73, 0.92, 0.93, 0.9, 
    0.88, 0.86, 0.78, 0.88, 0.91, 0.89, 0.87, 0.87, 0.87, 0.89, 0.85, 0.84, 
    0.79, 0.78, 0.79, 0.81, 0.8, 0.85, 0.85, 0.86, 0.72, 0.85, 0.85, 0.85, 
    0.81, 0.82, 0.8, 0.84, 0.79, 0.71, 0.69, 0.65, 0.69, 0.67, 0.66, 0.66, 
    0.65, 0.68, 0.73, 0.75, 0.79, 0.85, 0.89, 0.91, 0.91, 0.9, 0.9, 0.92, 
    0.92, 0.92, 0.91, 0.93, 0.96, 0.96, 0.93, 0.92, 0.91, 0.86, 0.84, 0.82, 
    0.77, 0.82, 0.78, 0.8, 0.84, 0.82, 0.88, 0.86, 0.84, 0.87, 0.94, 0.94, 
    0.94, 0.94, 0.91, 0.94, 0.89, 0.92, 0.87, 0.87, 0.86, 0.77, 0.73, 0.75, 
    0.7, 0.67, 0.7, 0.81, 0.8, 0.77, 0.79, 0.81, 0.79, 0.77, 0.76, 0.82, 
    0.88, 0.83, 0.82, 0.81, 0.78, 0.79, 0.79, 0.79, 0.78, 0.72, 0.71, 0.68, 
    0.68, 0.66, 0.68, 0.69, 0.68, 0.65, 0.74, 0.71, 0.7, 0.7, 0.72, 0.7, 
    0.68, 0.66, 0.65, 0.66, 0.67, 0.67, 0.66, 0.65, 0.66, 0.65, 0.65, 0.61, 
    0.5, 0.48, 0.49, 0.55, 0.49, 0.58, 0.57, 0.54, 0.6, 0.54, 0.52, 0.57, 
    0.65, 0.6, 0.58, 0.62, 0.63, 0.64, 0.65, 0.62, 0.54, 0.52, 0.52, 0.53, 
    0.64, 0.61, 0.58, 0.61, 0.6, 0.62, 0.63, 0.62, 0.63, 0.69, 0.72, 0.72, 
    0.71, 0.8, 0.83, 0.77, 0.74, 0.77, 0.75, 0.72, 0.62, 0.54, 0.52, 0.53, 
    0.6, 0.46, 0.62, 0.63, 0.55, 0.67, 0.64, 0.7, 0.69, 0.71, 0.72, 0.63, 
    0.62, 0.62, 0.63, 0.65, 0.62, 0.61, 0.63, 0.65, 0.63, 0.58, 0.55, 0.58, 
    0.54, 0.59, 0.52, 0.54, 0.54, 0.62, 0.58, 0.53, 0.59, 0.61, 0.68, 0.68, 
    0.72, 0.78, 0.72, 0.74, 0.75, 0.73, 0.66, 0.68, 0.6, 0.52, 0.59, 0.6, 
    0.48, 0.57, 0.58, 0.46, 0.56, 0.63, 0.62, 0.61, 0.62, 0.67, 0.78, 0.78, 
    0.8, 0.86, 0.85, 0.81, 0.86, 0.81, 0.68, 0.73, 0.58, 0.53, 0.59, 0.47, 
    0.66, 0.66, 0.72, 0.67, 0.71, 0.76, 0.76, 0.75, 0.79, 0.79, 0.82, 0.85, 
    0.87, 0.89, 0.91, 0.93, 0.94, 0.94, 0.92, 0.92, 0.92, 0.89, 0.86, 0.86, 
    0.69, 0.72, 0.64, 0.7, 0.67, 0.61, 0.69, 0.73, 0.78, 0.79, 0.86, 0.87, 
    0.83, 0.84, 0.8, 0.78, 0.76, 0.76, 0.8, 0.85, 0.85, 0.84, 0.78, 0.76, 
    0.74, 0.71, 0.64, 0.65, 0.64, 0.63, 0.65, 0.66, 0.59, 0.6, 0.67, 0.71, 
    0.72, 0.72, 0.73, 0.7, 0.7, 0.72, 0.72, 0.69, 0.64, 0.61, 0.65, 0.65, 
    0.61, 0.64, 0.6, 0.66, 0.63, 0.63, 0.64, 0.68, 0.66, 0.68, 0.75, 0.76, 
    0.74, 0.76, 0.76, 0.71, 0.71, 0.61, 0.63, 0.56, 0.53, 0.62, 0.58, 0.5, 
    0.56, 0.47, 0.59, 0.64, 0.65, 0.61, 0.62, 0.66, 0.7, 0.66, 0.67, 0.68, 
    0.68, 0.71, 0.72, 0.74, 0.69, 0.67, 0.62, 0.66, 0.68, 0.64, 0.57, 0.7, 
    0.73, 0.75, 0.76, 0.79, 0.79, 0.72, 0.85, 0.7, 0.68, 0.71, 0.7, 0.7, 
    0.71, 0.69, 0.69, 0.68, 0.64, 0.62, 0.63, 0.7, 0.63, 0.61, 0.64, 0.68, 
    0.7, 0.75, 0.76, 0.74, 0.77, 0.78, 0.75, 0.79, 0.84, 0.9, 0.9, 0.91, 
    0.91, 0.91, 0.94, 0.95, 0.92, 0.89, 0.88, 0.87, 0.79, 0.77, 0.79, 0.85, 
    0.81, 0.77, 0.81, 0.79, 0.75, 0.73, 0.77, 0.8, 0.78, 0.78, 0.79, 0.81, 
    0.88, 0.89, 0.94, 0.93, 0.92, 0.9, 0.89, 0.88, 0.96, 0.85, 0.8, 0.58, 
    0.61, 0.61, 0.58, 0.68, 0.69, 0.66, 0.66, 0.7, 0.7, 0.71, 0.71, 0.71, 
    0.77, 0.8, 0.79, 0.81, 0.74, 0.68, 0.58, 0.65, 0.59, 0.58, 0.63, 0.61, 
    0.6, 0.62, 0.52, 0.56, 0.6, 0.6, 0.6, 0.63, 0.63, 0.64, 0.71, 0.79, 0.77, 
    0.79, 0.78, 0.78, 0.79, 0.78, 0.71, 0.76, 0.68, 0.67, 0.72, 0.71, 0.64, 
    0.69, 0.66, 0.66, 0.65, 0.68, 0.71, 0.72, 0.71, 0.73, 0.73, 0.74, 0.75, 
    0.76, 0.76, 0.79, 0.81, 0.78, 0.78, 0.77, 0.76, 0.72, 0.72, 0.68, 0.66, 
    0.69, 0.66, 0.65, 0.68, 0.7, 0.74, 0.71, 0.73, 0.73, 0.75, 0.78, 0.77, 
    0.8, 0.76, 0.8, 0.8, 0.78, 0.78, 0.78, 0.76, 0.77, 0.71, 0.71, 0.68, 
    0.71, 0.68, 0.69, 0.68, 0.68, 0.66, 0.69, 0.7, 0.72, 0.67, 0.66, 0.65, 
    0.69, 0.71, 0.72, 0.67, 0.66, 0.65, 0.65, 0.63, 0.68, 0.66, 0.63, 0.59, 
    0.54, 0.55, 0.54, 0.55, 0.5, 0.59, 0.57, 0.61, 0.61, 0.62, 0.63, 0.71, 
    0.73, 0.69, 0.69, 0.67, 0.65, 0.64, 0.63, 0.57, 0.68, 0.62, 0.6, 0.61, 
    0.82, 0.82, 0.75, 0.72, 0.71, 0.65, 0.66, 0.7, 0.67, 0.67, 0.68, 0.7, 
    0.64, 0.66, 0.62, 0.62, 0.67, 0.68, 0.67, 0.7, 0.77, 0.67, 0.7, 0.6, 
    0.62, 0.63, 0.61, 0.61, 0.64, 0.65, 0.71, 0.72, 0.77, 0.75, 0.75, 0.75, 
    0.75, 0.74, 0.75, 0.74, 0.69, 0.74, 0.69, 0.68, 0.63, 0.64, 0.57, 0.62, 
    0.6, 0.6, 0.59, 0.65, 0.66, 0.72, 0.76, 0.73, 0.75, 0.76, 0.78, 0.83, 
    0.85, 0.81, 0.82, 0.87, 0.9, 0.95, 0.94, 0.89, 0.93, 0.92, 0.9, 0.93, 
    0.9, 0.9, 0.89, 0.91, 0.91, 0.92, 0.93, 0.94, 0.94, 0.95, 0.97, 0.96, 
    0.97, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.96, 0.95, 0.93, 0.88, 0.88, 
    0.84, 0.91, 0.85, 0.78, 0.68, 0.63, 0.66, 0.67, 0.66, 0.7, 0.69, 0.71, 
    0.72, 0.69, 0.68, 0.68, 0.67, 0.66, 0.63, 0.65, 0.64, 0.65, 0.62, 0.6, 
    0.6, 0.6, 0.62, 0.63, 0.64, 0.64, 0.67, 0.64, 0.67, 0.66, 0.65, 0.64, 
    0.61, 0.58, 0.6, 0.59, 0.55, 0.67, 0.56, 0.68, 0.84, 0.85, 0.8, 0.78, 
    0.74, 0.8, 0.81, 0.82, 0.83, 0.79, 0.71, 0.77, 0.85, 0.88, 0.91, 0.92, 
    0.92, 0.92, 0.94, 0.92, 0.91, 0.93, 0.92, 0.87, 0.9, 0.87, 0.86, 0.83, 
    0.79, 0.81, 0.82, 0.89, 0.82, 0.86, 0.72, 0.68, 0.64, 0.63, 0.61, 0.59, 
    0.58, 0.58, 0.61, 0.56, 0.55, 0.55, 0.57, 0.56, 0.53, 0.52, 0.53, 0.55, 
    0.55, 0.55, 0.56, 0.57, 0.59, 0.6, 0.57, 0.55, 0.53, 0.53, 0.54, 0.57, 
    0.56, 0.53, 0.62, 0.56, 0.59, 0.6, 0.52, 0.5, 0.49, 0.53, 0.47, 0.47, 
    0.51, 0.54, 0.56, 0.52, 0.57, 0.54, 0.55, 0.57, 0.59, 0.62, 0.65, 0.7, 
    0.7, 0.68, 0.69, 0.75, 0.6, 0.59, 0.6, 0.57, 0.59, 0.56, 0.64, 0.63, 
    0.56, 0.56, 0.62, 0.73, 0.73, 0.77, 0.83, 0.75, 0.8, 0.78, 0.69, 0.63, 
    0.65, 0.66, 0.59, 0.69, 0.64, 0.61, 0.65, 0.63, 0.56, 0.54, 0.51, 0.54, 
    0.58, 0.54, 0.56, 0.51, 0.58, 0.58, 0.65, 0.66, 0.71, 0.76, 0.8, 0.79, 
    0.73, 0.73, 0.81, 0.95, 0.91, 0.78, 0.72, 0.72, 0.72, 0.66, 0.65, 0.66, 
    0.7, 0.66, 0.71, 0.84, 0.78, 0.73, 0.77, 0.79, 0.8, 0.78, 0.81, 0.81, 
    0.9, 0.95, 0.96, 0.95, 0.93, 0.92, 0.92, 0.94, 0.94, 0.9, 0.92, 0.92, 
    0.92, 0.91, 0.86, 0.84, 0.88, 0.9, 0.91, 0.95, 0.96, 0.98, 0.96, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.98, 0.96, 0.97, 
    0.96, 0.95, 0.96, 0.97, 0.97, 0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.94, 0.88, 0.85, 0.85, 0.86, 
    0.83, 0.67, 0.62, 0.68, 0.7, 0.7, 0.67, 0.67, 0.68, 0.7, 0.81, 0.83, 
    0.81, 0.88, 0.86, 0.89, 0.79, 0.72, 0.74, 0.84, 0.78, 0.78, 0.8, 0.71, 
    0.75, 0.8, 0.76, 0.76, 0.75, 0.77, 0.78, 0.75, 0.79, 0.78, 0.84, 0.81, 
    0.8, 0.85, 0.8, 0.88, 0.78, 0.7, 0.77, 0.74, 0.77, 0.73, 0.76, 0.77, 
    0.76, 0.81, 0.82, 0.88, 0.87, 0.9, 0.85, 0.9, 0.85, 0.92, 0.98, 0.99, 
    0.86, 0.87, 0.88, 0.86, 0.82, 0.89, 0.88, 0.85, 0.78, 0.85, 0.85, 0.77, 
    0.81, 0.82, 0.83, 0.83, 0.82, 0.81, 0.78, 0.77, 0.82, 0.81, 0.85, 0.9, 
    0.9, 0.94, 0.96, 0.96, 0.97, 0.98, 0.9, 0.92, 0.93, 0.9, 0.92, 0.93, 
    0.88, 0.89, 0.86, 0.9, 0.9, 0.91, 0.9, 0.86, 0.82, 0.89, 0.84, 0.82, 
    0.86, 0.84, 0.81, 0.81, 0.79, 0.75, 0.77, 0.78, 0.82, 0.81, 0.81, 0.78, 
    0.73, 0.73, 0.73, 0.67, 0.75, 0.71, 0.76, 0.77, 0.76, 0.78, 0.79, 0.76, 
    0.83, 0.86, 0.85, 0.87, 0.92, 0.84, 0.81, 0.76, 0.73, 0.67, 0.58, 0.62, 
    0.58, 0.55, 0.59, 0.57, 0.55, 0.51, 0.52, 0.46, 0.42, 0.5, 0.52, 0.41, 
    0.54, 0.5, 0.48, 0.55, 0.54, 0.51, 0.55, 0.54, 0.56, 0.59, 0.63, 0.6, 
    0.61, 0.64, 0.67, 0.68, 0.69, 0.69, 0.69, 0.68, 0.68, 0.67, 0.73, 0.73, 
    0.75, 0.71, 0.71, 0.74, 0.75, 0.75, 0.76, 0.81, 0.87, 0.87, 0.85, 0.81, 
    0.83, 0.88, 0.87, 0.83, 0.75, 0.66, 0.58, 0.6, 0.58, 0.61, 0.64, 0.62, 
    0.58, 0.58, 0.59, 0.58, 0.59, 0.6, 0.62, 0.56, 0.58, 0.57, 0.6, 0.6, 
    0.57, 0.66, 0.69, 0.7, 0.7, 0.67, 0.64, 0.64, 0.65, 0.69, 0.69, 0.69, 
    0.75, 0.72, 0.7, 0.73, 0.69, 0.66, 0.69, 0.68, 0.63, 0.63, 0.67, 0.71, 
    0.67, 0.76, 0.78, 0.79, 0.76, 0.69, 0.63, 0.64, 0.66, 0.64, 0.67, 0.7, 
    0.75, 0.77, 0.77, 0.77, 0.75, 0.77, 0.72, 0.64, 0.59, 0.65, 0.57, 0.62, 
    0.65, 0.6, 0.58, 0.58, 0.6, 0.63, 0.62, 0.58, 0.54, 0.59, 0.62, 0.54, 
    0.62, 0.64, 0.6, 0.48, 0.48, 0.53, 0.5, 0.5, 0.51, 0.51, 0.47, 0.5, 0.49, 
    0.56, 0.57, 0.6, 0.57, 0.58, 0.6, 0.63, 0.64, 0.7, 0.66, 0.67, 0.68, 
    0.69, 0.68, 0.7, 0.69, 0.67, 0.64, 0.57, 0.55, 0.56, 0.52, 0.5, 0.53, 
    0.54, 0.52, 0.52, 0.54, 0.53, 0.58, 0.58, 0.58, 0.63, 0.66, 0.59, 0.57, 
    0.59, 0.58, 0.63, 0.61, 0.49, 0.51, 0.61, 0.57, 0.52, 0.48, 0.52, 0.58, 
    0.5, 0.59, 0.47, 0.55, 0.54, 0.51, 0.48, 0.53, 0.54, 0.55, 0.55, 0.55, 
    0.54, 0.55, 0.52, 0.45, 0.42, 0.44, 0.42, 0.44, 0.5, 0.58, 0.6, 0.64, 
    0.68, 0.69, 0.72, 0.88, 0.82, 0.86, 0.81, 0.83, 0.85, 0.84, 0.86, 0.88, 
    0.88, 0.9, 0.9, 0.83, 0.88, 0.89, 0.9, 0.87, 0.81, 0.82, 0.76, 0.79, 
    0.75, 0.71, 0.69, 0.71, 0.71, 0.76, 0.76, 0.76, 0.77, 0.81, 0.85, 0.85, 
    0.83, 0.82, 0.86, 0.85, 0.91, 0.89, 0.91, 0.96, 0.96, 0.96, 0.92, 0.97, 
    0.91, 0.96, 0.97, 0.94, 0.88, 0.83, 0.92, 0.87, 0.85, 0.85, 0.86, 0.8, 
    0.82, 0.8, 0.88, 0.87, 0.91, 0.95, 0.97, 0.98, 0.98, 0.97, 0.92, 0.75, 
    0.78, 0.8, 0.76, 0.73, 0.83, 0.76, 0.82, 0.82, 0.81, 0.82, 0.84, 0.87, 
    0.9, 0.91, 0.93, 0.96, 0.98, 0.98, 0.98, 0.82, 0.89, 0.85, 0.87, 0.76, 
    0.71, 0.7, 0.67, 0.64, 0.63, 0.67, 0.69, 0.72, 0.78, 0.79, 0.79, 0.81, 
    0.77, 0.8, 0.82, 0.76, 0.81, 0.77, 0.81, 0.74, 0.79, 0.87, 0.83, 0.81, 
    0.73, 0.71, 0.68, 0.72, 0.73, 0.81, 0.89, 0.92, 0.97, 0.97, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.98, 0.96, 0.98, 0.86, 0.87, 0.89, 0.86, 0.87, 0.77, 
    0.68, 0.73, 0.67, 0.76, 0.73, 0.71, 0.73, 0.66, 0.74, 0.75, 0.73, 0.69, 
    0.72, 0.83, 0.82, 0.88, 0.86, 0.82, 0.78, 0.75, 0.82, 0.87, 0.97, 0.88, 
    0.91, 0.8, 0.73, 0.74, 0.75, 0.78, 0.77, 0.74, 0.71, 0.65, 0.68, 0.71, 
    0.71, 0.73, 0.75, 0.8, 0.82, 0.73, 0.7, 0.76, 0.81, 0.78, 0.76, 0.74, 
    0.73, 0.8, 0.89, 0.85, 0.91, 0.91, 0.91, 0.91, 0.92, 0.92, 0.92, 0.92, 
    0.9, 0.9, 0.9, 0.9, 0.89, 0.91, 0.81, 0.8, 0.79, 0.78, 0.8, 0.81, 0.8, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.83, 0.85, 0.9, 0.88, 0.85, 0.87, 0.8, 0.82, 
    0.86, 0.79, 0.8, 0.83, 0.85, 0.8, 0.8, 0.89, 0.92, 0.95, 0.93, 0.97, 
    0.96, 0.93, 0.94, 0.89, 0.85, 0.84, 0.85, 0.82, 0.82, 0.83, 0.84, 0.85, 
    0.78, 0.82, 0.79, 0.83, 0.84, 0.83, 0.79, 0.79, 0.8, 0.88, 0.89, 0.88, 
    0.87, 0.88, 0.89, 0.94, 0.92, 0.92, 0.9, 0.9, 0.87, 0.89, 0.85, 0.96, 
    0.95, 0.88, 0.9, 0.91, 0.9, 0.89, 0.87, 0.72, 0.65, 0.75, 0.76, 0.75, 
    0.71, 0.76, 0.68, 0.63, 0.72, 0.67, 0.62, 0.67, 0.69, 0.75, 0.75, 0.78, 
    0.69, 0.74, 0.7, 0.77, 0.66, 0.75, 0.75, 0.68, 0.55, 0.52, 0.56, 0.69, 
    0.66, 0.76, 0.78, 0.7, 0.7, 0.83, 0.78, 0.82, 0.84, 0.89, 0.94, 0.92, 
    0.94, 0.94, 0.95, 0.95, 0.92, 0.9, 0.92, 0.96, 0.96, 0.96, 0.98, 0.98, 
    0.97, 0.96, 0.94, 0.94, 0.89, 0.83, 0.86, 0.82, 0.84, 0.86, 0.87, 0.83, 
    0.83, 0.92, 0.92, 0.83, 0.89, 0.89, 0.84, 0.84, 0.86, 0.88, 0.74, 0.83, 
    0.86, 0.86, 0.89, 0.91, 0.91, 0.91, 0.92, 0.98, 0.99, 0.91, 0.93, 0.91, 
    0.9, 0.89, 0.98, 0.99, 0.99, 0.99, 0.97, 0.95, 0.93, 0.91, 0.89, 0.89, 
    0.83, 0.82, 0.79, 0.8, 0.81, 0.91, 0.9, 0.89, 0.91, 0.91, 0.87, 0.91, 
    0.94, 0.94, 0.89, 0.82, 0.83, 0.82, 0.76, 0.75, 0.74, 0.68, 0.68, 0.7, 
    0.77, 0.76, 0.75, 0.76, 0.7, 0.77, 0.72, 0.8, 0.76, 0.74, 0.74, 0.76, 
    0.76, 0.72, 0.74, 0.74, 0.71, 0.67, 0.69, 0.68, 0.76, 0.74, 0.82, 0.81, 
    0.8, 0.83, 0.87, 0.88, 0.96, 0.96, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 
    0.99, 1, 1, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.92, 0.93, 0.89, 0.89, 0.9, 0.82, 0.88, 0.89, 0.86, 
    0.86, 0.9, 0.94, 0.98, 0.99, 0.99, 0.99, 0.96, 0.89, 0.87, 0.88, 0.89, 
    0.8, 0.83, 0.81, 0.84, 0.88, 0.82, 0.89, 0.92, 0.93, 0.93, 0.97, 0.89, 
    0.91, 0.91, 0.71, 0.77, 0.75, 0.72, 0.74, 0.75, 0.79, 0.81, 0.84, 0.87, 
    0.92, 0.75, 0.8, 0.8, 0.79, 0.83, 0.83, 0.85, 0.89, 0.89, 0.9, 0.85, 
    0.85, 0.86, 0.84, 0.76, 0.71, 0.73, 0.71, 0.77, 0.76, 0.77, 0.85, 0.86, 
    0.88, 0.91, 0.93, 0.94, 0.97, 0.97, 0.99, 0.98, 0.97, 0.94, 0.95, 0.94, 
    0.9, 0.92, 0.9, 0.87, 0.85, 0.93, 0.93, 0.92, 0.84, 0.69, 0.67, 0.67, 
    0.66, 0.66, 0.7, 0.7, 0.69, 0.79, 0.8, 0.82, 0.81, 0.81, 0.8, 0.75, 0.76, 
    0.76, 0.8, 0.79, 0.74, 0.76, 0.81, 0.84, 0.81, 0.75, 0.71, 0.66, 0.66, 
    0.66, 0.62, 0.67, 0.63, 0.65, 0.61, 0.61, 0.62, 0.65, 0.63, 0.66, 0.67, 
    0.72, 0.73, 0.75, 0.71, 0.67, 0.72, 0.77, 0.73, 0.7, 0.64, 0.64, 0.66, 
    0.69, 0.74, 0.73, 0.74, 0.75, 0.76, 0.76, 0.78, 0.74, 0.73, 0.72, 0.7, 
    0.69, 0.64, 0.61, 0.63, 0.63, 0.63, 0.62, 0.63, 0.64, 0.63, 0.62, 0.6, 
    0.6, 0.61, 0.64, 0.68, 0.72, 0.74, 0.72, 0.74, 0.72, 0.69, 0.7, 0.76, 
    0.71, 0.69, 0.7, 0.63, 0.57, 0.58, 0.57, 0.56, 0.56, 0.54, 0.52, 0.5, 
    0.52, 0.54, 0.52, 0.54, 0.59, 0.63, 0.67, 0.6, 0.62, 0.58, 0.57, 0.55, 
    0.54, 0.52, 0.5, 0.51, 0.45, 0.5, 0.52, 0.54, 0.54, 0.53, 0.52, 0.53, 
    0.58, 0.58, 0.64, 0.6, 0.64, 0.67, 0.67, 0.74, 0.66, 0.64, 0.62, 0.67, 
    0.66, 0.66, 0.6, 0.64, 0.64, 0.78, 0.78, 0.79, 0.79, 0.79, 0.8, 0.83, 
    0.81, 0.79, 0.7, 0.67, 0.64, 0.64, 0.63, 0.65, 0.64, 0.61, 0.66, 0.65, 
    0.64, 0.62, 0.68, 0.7, 0.69, 0.72, 0.74, 0.76, 0.77, 0.75, 0.73, 0.66, 
    0.71, 0.75, 0.72, 0.73, 0.73, 0.72, 0.71, 0.7, 0.7, 0.64, 0.65, 0.71, 
    0.74, 0.71, 0.8, 0.82, 0.85, 0.83, 0.78, 0.8, 0.8, 0.8, 0.8, 0.84, 0.73, 
    0.72, 0.78, 0.84, 0.86, 0.82, 0.78, 0.79, 0.82, 0.82, 0.71, 0.73, 0.6, 
    0.63, 0.67, 0.73, 0.77, 0.78, 0.73, 0.79, 0.79, 0.8, 0.82, 0.82, 0.8, 
    0.84, 0.87, 0.91, 0.95, 0.91, 0.97, 0.98, 0.98, 0.92, 0.91, 0.92, 0.81, 
    0.72, 0.57, 0.46, 0.42, 0.46, 0.49, 0.51, 0.55, 0.6, 0.64, 0.61, 0.66, 
    0.68, 0.69, 0.71, 0.7, 0.71, 0.69, 0.75, 0.72, 0.7, 0.67, 0.64, 0.63, 
    0.61, 0.68, 0.74, 0.77, 0.74, 0.85, 0.95, 0.96, 0.95, 0.96, 0.96, 0.95, 
    0.95, 0.95, 0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.9, 0.9, 
    0.91, 0.85, 0.87, 0.89, 0.82, 0.82, 0.79, 0.82, 0.76, 0.72, 0.77, 0.83, 
    0.78, 0.86, 0.85, 0.76, 0.82, 0.84, 0.9, 0.87, 0.86, 0.83, 0.82, 0.88, 
    0.79, 0.88, 0.92, 0.8, 0.78, 0.77, 0.81, 0.86, 0.82, 0.79, 0.8, 0.77, 
    0.86, 0.83, 0.85, 0.87, 0.91, 0.87, 0.83, 0.81, 0.85, 0.83, 0.81, 0.79, 
    0.79, 0.83, 0.84, 0.8, 0.83, 0.82, 0.82, 0.83, 0.84, 0.81, 0.86, 0.84, 
    0.85, 0.84, 0.82, 0.8, 0.83, 0.83, 0.85, 0.84, 0.8, 0.8, 0.81, 0.82, 
    0.77, 0.81, 0.78, 0.76, 0.84, 0.82, 0.76, 0.82, 0.84, 0.84, 0.79, 0.84, 
    0.85, 0.83, 0.87, 0.86, 0.88, 0.9, 0.9, 0.9, 0.9, 0.88, 0.82, 0.86, 0.76, 
    0.72, 0.71, 0.71, 0.7, 0.66, 0.66, 0.68, 0.67, 0.67, 0.8, 0.8, 0.77, 
    0.82, 0.78, 0.84, 0.81, 0.79, 0.79, 0.77, 0.78, 0.77, 0.75, 0.75, 0.75, 
    0.75, 0.76, 0.75, 0.77, 0.78, 0.78, 0.76, 0.8, 0.75, 0.73, 0.82, 0.8, 
    0.78, 0.8, 0.81, 0.74, 0.71, 0.65, 0.65, 0.66, 0.7, 0.68, 0.67, 0.65, 
    0.67, 0.65, 0.67, 0.63, 0.68, 0.66, 0.6, 0.71, 0.83, 0.68, 0.66, 0.69, 
    0.72, 0.73, 0.72, 0.72, 0.74, 0.78, 0.77, 0.77, 0.75, 0.74, 0.76, 0.77, 
    0.79, 0.77, 0.75, 0.75, 0.76, 0.76, 0.74, 0.75, 0.77, 0.83, 0.86, 0.94, 
    0.95, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.9, 0.95, 0.93, 0.86, 
    0.88, 0.92, 0.97, 0.96, 0.94, 0.92, 0.88, 0.89, 0.9, 0.84, 0.91, 0.91, 
    0.91, 0.96, 0.98, 0.99, 0.98, 0.98, 0.97, 0.96, 0.92, 0.94, 0.93, 0.92, 
    0.86, 0.87, 0.87, 0.81, 0.78, 0.75, 0.68, 0.69, 0.69, 0.64, 0.6, 0.62, 
    0.66, 0.75, 0.73, 0.74, 0.8, 0.78, 0.8, 0.85, 0.84, 0.85, 0.9, 0.9, 0.89, 
    0.89, 0.83, 0.87, 0.84, 0.84, 0.85, 0.86, 0.88, 0.92, 0.92, 0.9, 0.9, 
    0.87, 0.85, 0.85, 0.79, 0.8, 0.79, 0.77, 0.77, 0.81, 0.84, 0.82, 0.81, 
    0.81, 0.87, 0.88, 0.88, 0.84, 0.77, 0.81, 0.79, 0.8, 0.82, 0.84, 0.85, 
    0.96, 0.98, 0.99, 0.99, 0.99, 1, 0.99, 1, 1, 1, 0.99, 1, 0.99, 0.99, 
    0.96, 0.97, 0.98, 0.99, 0.99, 0.99, 1, 0.99, 1, 1, 0.96, 0.97, 0.94, 0.9, 
    0.89, 0.91, 0.88, 0.81, 0.81, 0.78, 0.78, 0.77, 0.76, 0.72, 0.79, 0.87, 
    0.84, 0.81, 0.75, 0.81, 0.85, 0.85, 0.85, 0.83, 0.84, 0.91, 0.92, 0.89, 
    0.91, 0.88, 0.9, 0.91, 0.93, 0.91, 0.92, 0.94, 0.93, 0.92, 0.91, 0.87, 
    0.88, 0.88, 0.8, 0.81, 0.86, 0.83, 0.82, 0.75, 0.72, 0.7, 0.63, 0.62, 
    0.62, 0.64, 0.69, 0.67, 0.7, 0.75, 0.77, 0.75, 0.72, 0.66, 0.68, 0.66, 
    0.7, 0.64, 0.65, 0.67, 0.69, 0.69, 0.71, 0.72, 0.7, 0.76, 0.76, 0.76, 
    0.75, 0.74, 0.77, 0.8, 0.8, 0.79, 0.78, 0.78, 0.79, 0.77, 0.72, 0.7, 0.7, 
    0.7, 0.73, 0.75, 0.75, 0.69, 0.68, 0.74, 0.76, 0.74, 0.81, 0.82, 0.8, 
    0.8, 0.76, 0.87, 0.88, 0.88, 0.88, 0.87, 0.84, 0.89, 0.88, 0.86, 0.84, 
    0.84, 0.81, 0.9, 0.87, 0.89, 0.97, 0.99, 0.98, 0.99, 1, 1, 0.99, 0.88, 
    0.87, 0.83, 0.79, 0.77, 0.75, 0.77, 0.76, 0.77, 0.74, 0.75, 0.74, 0.76, 
    0.79, 0.74, 0.82, 0.83, 0.84, 0.87, 0.86, 0.87, 0.88, 0.88, 0.81, 0.8, 
    0.82, 0.82, 0.84, 0.83, 0.8, 0.75, 0.75, 0.77, 0.75, 0.75, 0.75, 0.78, 
    0.76, 0.74, 0.74, 0.87, 0.81, 0.84, 0.9, 0.73, 0.6, 0.63, 0.66, 0.68, 
    0.69, 0.68, 0.7, 0.83, 0.84, 0.81, 0.82, 0.76, 0.78, 0.68, 0.63, 0.61, 
    0.67, 0.69, 0.59, 0.61, 0.63, 0.63, 0.64, 0.62, 0.58, 0.61, 0.76, 0.7, 
    0.68, 0.59, 0.57, 0.54, 0.58, 0.57, 0.61, 0.6, 0.66, 0.68, 0.7, 0.72, 
    0.75, 0.7, 0.77, 0.77, 0.77, 0.81, 0.87, 0.83, 0.84, 0.86, 0.86, 0.84, 
    0.83, 0.88, 0.88, 0.87, 0.88, 0.8, 0.76, 0.81, 0.84, 0.82, 0.73, 0.7, 
    0.66, 0.64, 0.69, 0.67, 0.66, 0.7, 0.69, 0.64, 0.62, 0.67, 0.72, 0.7, 
    0.8, 0.83, 0.87, 0.89, 0.93, 0.95, 0.96, 0.95, 0.95, 0.94, 0.92, 0.89, 
    0.77, 0.74, 0.77, 0.75, 0.74, 0.72, 0.74, 0.75, 0.71, 0.81, 0.66, 0.62, 
    0.67, 0.66, 0.62, 0.64, 0.7, 0.76, 0.85, 0.87, 0.92, 0.89, 0.82, 0.89, 
    0.87, 0.93, 0.95, 0.92, 0.88, 0.87, 0.96, 0.92, 0.88, 0.83, 0.8, 0.83, 
    0.81, 0.84, 0.86, 0.87, 0.86, 0.89, 0.98, 0.98, 0.97, 0.96, 0.95, 0.97, 
    0.97, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 1, 1, 
    1, 0.99, 1, 1, 1, 0.99, 1, 1, 1, 1, 1, 0.99, 1, 1, 1, 0.99, 1, 1, 0.99, 
    0.99, 1, 1, 0.99, 0.97, 0.95, 0.98, 0.98, 0.94, 0.93, 0.93, 0.84, 0.81, 
    0.82, 0.74, 0.69, 0.55, 0.73, 0.67, 0.79, 0.76, 0.74, 0.81, 0.78, 0.76, 
    0.75, 0.67, 0.73, 0.68, 0.72, 0.7, 0.7, 0.68, 0.74, 0.72, 0.71, 0.74, 
    0.73, 0.74, 0.69, 0.69, 0.69, 0.69, 0.74, 0.77, 0.78, 0.79, 0.84, 0.92, 
    0.93, 0.9, 0.92, 0.91, 0.9, 0.92, 0.84, 0.88, 0.78, 0.77, 0.74, 0.7, 
    0.63, 0.6, 0.67, 0.71, 0.69, 0.69, 0.72, 0.76, 0.77, 0.77, 0.83, 0.83, 
    0.83, 0.84, 0.86, 0.9, 0.91, 0.9, 0.89, 0.89, 0.88, 0.89, 0.86, 0.87, 
    0.88, 0.98, 0.99, 0.98, 0.99, 0.91, 0.9, 0.9, 0.93, 0.88, 0.9, 0.86, 
    0.86, 0.85, 0.89, 0.92, 0.92, 0.83, 0.9, 0.88, 0.83, 0.77, 0.74, 0.79, 
    0.66, 0.63, 0.63, 0.65, 0.69, 0.73, 0.72, 0.72, 0.76, 0.83, 0.84, 0.82, 
    0.82, 0.82, 0.85, 0.84, 0.84, 0.84, 0.82, 0.79, 0.76, 0.77, 0.78, 0.76, 
    0.78, 0.8, 0.8, 0.81, 0.92, 0.94, 0.94, 0.93, 0.94, 0.95, 0.95, 0.97, 
    0.99, 0.98, 0.97, 0.96, 0.93, 0.91, 0.79, 0.88, 0.94, 0.86, 0.76, 0.7, 
    0.68, 0.72, 0.71, 0.81, 0.85, 0.9, 0.91, 0.89, 0.86, 0.84, 0.86, 0.86, 
    0.86, 0.77, 0.85, 0.85, 0.84, 0.8, 0.73, 0.75, 0.77, 0.78, 0.76, 0.78, 
    0.8, 0.84, 0.78, 0.82, 0.86, 0.86, 0.89, 0.86, 0.9, 0.9, 0.91, 0.91, 
    0.89, 0.91, 0.9, 0.91, 0.89, 0.89, 0.87, 0.81, 0.81, 0.77, 0.75, 0.8, 
    0.84, 0.85, 0.82, 0.83, 0.89, 0.9, 0.92, 0.93, 0.94, 0.91, 0.89, 0.94, 
    0.98, 0.99, 0.97, 0.94, 0.96, 0.97, 0.94, 0.96, 0.94, 0.9, 0.89, 0.93, 
    0.89, 0.78, 0.75, 0.8, 0.77, 0.75, 0.72, 0.72, 0.69, 0.75, 0.71, 0.73, 
    0.77, 0.76, 0.76, 0.74, 0.78, 0.7, 0.7, 0.68, 0.68, 0.72, 0.76, 0.75, 
    0.74, 0.77, 0.76, 0.75, 0.75, 0.77, 0.77, 0.72, 0.74, 0.74, 0.75, 0.74, 
    0.79, 0.77, 0.76, 0.74, 0.78, 0.84, 0.82, 0.7, 0.7, 0.67, 0.77, 0.71, 
    0.72, 0.71, 0.73, 0.72, 0.72, 0.71, 0.71, 0.72, 0.74, 0.77, 0.69, 0.62, 
    0.66, 0.64, 0.66, 0.76, 0.68, 0.63, 0.63, 0.56, 0.66, 0.63, 0.6, 0.62, 
    0.63, 0.63, 0.62, 0.66, 0.58, 0.7, 0.67, 0.67, 0.7, 0.66, 0.63, 0.64, 
    0.67, 0.63, 0.7, 0.72, 0.66, 0.62, 0.6, 0.58, 0.59, 0.56, 0.59, 0.6, 
    0.59, 0.6, 0.66, 0.63, 0.69, 0.69, 0.76, 0.81, 0.78, 0.8, 0.79, 0.76, 
    0.77, 0.71, 0.73, 0.73, 0.72, 0.69, 0.74, 0.73, 0.71, 0.73, 0.75, 0.74, 
    0.71, 0.65, 0.65, 0.66, 0.64, 0.67, 0.71, 0.78, 0.78, 0.87, 0.86, 0.87, 
    0.85, 0.84, 0.83, 0.98, 0.84, 0.84, 0.85, 0.79, 0.78, 0.79, 0.79, 0.78, 
    0.81, 0.83, 0.84, 0.85, 0.87, 0.88, 0.89, 0.9, 0.91, 0.91, 0.92, 0.92, 
    0.94, 0.94, 0.91, 0.89, 0.87, 0.84, 0.85, 0.84, 0.9, 0.86, 0.88, 0.89, 
    0.92, 0.93, 0.88, 0.89, 0.87, 0.87, 0.9, 0.9, 0.95, 0.95, 0.95, 0.88, 
    0.91, 0.91, 0.9, 0.91, 0.88, 0.83, 0.79, 0.71, 0.72, 0.72, 0.7, 0.74, 
    0.7, 0.64, 0.76, 0.7, 0.69, 0.75, 0.76, 0.76, 0.78, 0.77, 0.72, 0.75, 
    0.75, 0.77, 0.82, 0.81, 0.83, 0.86, 0.73, 0.77, 0.77, 0.73, 0.68, 0.63, 
    0.64, 0.65, 0.63, 0.62, 0.63, 0.69, 0.74, 0.77, 0.72, 0.75, 0.68, 0.71, 
    0.72, 0.73, 0.74, 0.67, 0.76, 0.8, 0.85, 0.88, 0.84, 0.82, 0.83, 0.84, 
    0.71, 0.73, 0.86, 0.86, 0.91, 0.84, 0.8, 0.83, 0.84, 0.89, 0.86, 0.8, 
    0.81, 0.82, 0.8, 0.82, 0.78, 0.72, 0.73, 0.72, 0.68, 0.72, 0.71, 0.72, 
    0.68, 0.7, 0.72, 0.71, 0.77, 0.82, 0.85, 0.83, 0.83, 0.79, 0.77, 0.79, 
    0.81, 0.83, 0.82, 0.81, 0.78, 0.77, 0.74, 0.73, 0.72, 0.68, 0.63, 0.63, 
    0.62, 0.6, 0.64, 0.67, 0.69, 0.68, 0.67, 0.73, 0.78, 0.77, 0.84, 0.86, 
    0.96, 0.94, 0.95, 0.95, 0.96, 0.94, 0.92, 0.93, 0.94, 0.93, 0.9, 0.93, 
    0.87, 0.85, 0.82, 0.81, 0.83, 0.84, 0.85, 0.89, 0.88, 0.87, 0.87, 0.87, 
    0.9, 0.91, 0.95, 0.98, 0.99, 0.99, 0.99, 0.98, 0.96, 0.97, 0.95, 0.89, 
    0.9, 0.86, 0.79, 0.68, 0.68, 0.7, 0.69, 0.68, 0.69, 0.68, 0.73, 0.74, 
    0.73, 0.73, 0.74, 0.79, 0.77, 0.78, 0.68, 0.7, 0.57, 0.57, 0.6, 0.65, 
    0.68, 0.69, 0.71, 0.71, 0.71, 0.75, 0.72, 0.77, 0.77, 0.93, 0.97, 0.98, 
    0.95, 0.96, 0.94, 0.88, 0.82, 0.83, 0.78, 0.77, 0.77, 0.74, 0.72, 0.7, 
    0.76, 0.73, 0.76, 0.73, 0.73, 0.81, 0.85, 0.84, 0.8, 0.84, 0.94, 0.85, 
    0.82, 0.91, 0.9, 0.89, 0.88, 0.89, 0.86, 0.78, 0.62, 0.61, 0.64, 0.72, 
    0.71, 0.77, 0.82, 0.84, 0.84, 0.86, 0.88, 0.88, 0.88, 0.85, 0.87, 0.8, 
    0.77, 0.81, 0.86, 0.71, 0.8, 0.77, 0.78, 0.75, 0.7, 0.71, 0.74, 0.68, 
    0.71, 0.7, 0.69, 0.75, 0.73, 0.83, 0.81, 0.78, 0.78, 0.89, 0.91, 0.94, 
    0.94, 0.96, 0.96, 0.94, 0.93, 0.82, 0.8, 0.73, 0.67, 0.72, 0.77, 0.7, 
    0.74, 0.78, 0.75, 0.86, 0.88, 0.87, 0.84, 0.81, 0.79, 0.84, 0.86, 0.89, 
    0.87, 0.84, 0.84, 0.81, 0.88, 0.86, 0.89, 0.87, 0.76, 0.74, 0.71, 0.77, 
    0.72, 0.78, 0.79, 0.8, 0.84, 0.83, 0.85, 0.82, 0.84, 0.81, 0.86, 0.75, 
    0.85, 0.83, 0.83, 0.78, 0.76, 0.74, 0.68, 0.7, 0.73, 0.76, 0.78, 0.79, 
    0.69, 0.65, 0.67, 0.76, 0.85, 0.82, 0.8, 0.72, 0.82, 0.8, 0.7, 0.74, 
    0.86, 0.87, 0.86, 0.85, 0.85, 0.84, 0.87, 0.87, 0.87, 0.87, 0.87, 0.82, 
    0.85, 0.87, 0.83, 0.84, 0.88, 0.91, 0.92, 0.81, 0.83, 0.86, 0.9, 0.9, 1, 
    0.89, 0.95, 0.95, 0.95, 0.9, 0.84, 0.82, 0.81, 0.83, 0.83, 0.85, 0.85, 
    0.8, 0.84, 0.87, 0.91, 0.93, 0.91, 0.93, 0.92, 0.94, 0.89, 0.92, 0.92, 
    0.91, 0.91, 0.95, 0.86, 0.91, 0.86, 0.86, 0.83, 0.81, 0.8, 0.84, 0.77, 
    0.78, 0.83, 0.85, 0.88, 0.92, 0.88, 0.84, 0.91, 0.93, 0.87, 0.9, 0.91, 
    0.93, 0.91, 0.9, 0.95, 0.84, 0.89, 0.85, 0.8, 0.78, 0.8, 0.87, 0.87, 
    0.79, 0.73, 0.81, 0.77, 0.76, 0.74, 0.72, 0.74, 0.72, 0.67, 0.77, 0.78, 
    0.79, 0.82, 0.82, 0.72, 0.86, 0.88, 0.87, 0.75, 0.77, 0.79, 0.76, 0.74, 
    0.71, 0.7, 0.69, 0.68, 0.77, 0.75, 0.74, 0.74, 0.77, 0.76, 0.75, 0.71, 
    0.7, 0.7, 0.65, 0.66, 0.61, 0.67, 0.64, 0.68, 0.61, 0.62, 0.65, 0.56, 
    0.59, 0.6, 0.62, 0.61, 0.61, 0.72, 0.72, 0.71, 0.7, 0.75, 0.77, 0.79, 
    0.74, 0.73, 0.71, 0.7, 0.65, 0.72, 0.73, 0.73, 0.73, 0.69, 0.75, 0.8, 
    0.78, 0.82, 0.79, 0.8, 0.87, 0.82, 0.91, 0.86, 0.86, 0.86, 0.88, 0.9, 
    0.91, 0.9, 0.89, 0.87, 0.86, 0.85, 0.9, 0.91, 0.86, 0.88, 0.86, 0.86, 
    0.87, 0.93, 0.95, 0.95, 0.91, 0.93, 0.96, 0.98, 0.98, 0.89, 0.89, 0.89, 
    0.9, 0.92, 0.92, 0.92, 0.88, 0.88, 0.88, 0.89, 0.89, 0.89, 0.9, 0.94, 
    0.94, 0.96, 0.94, 0.96, 0.98, 0.98, 0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.96, 0.97, 0.96, 0.97, 0.97, 0.97, 0.92, 0.84, 0.78, 0.8, 0.88, 
    0.89, 0.87, 0.85, 0.87, 0.88, 0.83, 0.85, 0.88, 0.85, 0.82, 0.89, 0.83, 
    0.82, 0.8, 0.88, 0.84, 0.76, 0.78, 0.79, 0.79, 0.73, 0.77, 0.79, 0.8, 
    0.79, 0.78, 0.78, 0.77, 0.81, 0.81, 0.81, 0.78, 0.81, 0.82, 0.81, 0.77, 
    0.78, 0.81, 0.85, 0.85, 0.83, 0.78, 0.72, 0.69, 0.67, 0.82, 0.82, 0.82, 
    0.82, 0.84, 0.85, 0.87, 0.9, 0.95, 0.92, 0.92, 0.92, 0.92, 0.94, 0.94, 
    0.95, 0.93, 0.93, 0.94, 0.93, 0.92, 0.93, 0.93, 0.94, 0.79, 0.79, 0.75, 
    0.88, 0.79, 0.81, 0.81, 0.76, 0.87, 0.84, 0.87, 0.9, 0.9, 0.87, 0.85, 
    0.87, 0.85, 0.91, 0.95, 0.92, 0.94, 0.88, 0.81, 0.82, 0.71, 0.66, 0.68, 
    0.71, 0.64, 0.8, 0.81, 0.8, 0.88, 0.88, 0.75, 0.8, 0.81, 0.85, 0.89, 
    0.91, 0.91, 0.93, 0.96, 0.85, 0.82, 0.87, 0.9, 0.9, 0.86, 0.91, 0.92, 
    0.84, 0.83, 0.82, 0.81, 0.81, 0.82, 0.71, 0.78, 0.76, 0.78, 0.76, 0.77, 
    0.82, 0.82, 0.94, 0.81, 0.9, 0.95, 0.96, 0.92, 0.94, 0.97, 0.96, 0.99, 
    0.99, 0.83, 0.76, 0.83, 0.77, 0.72, 0.77, 0.74, 0.73, 0.72, 0.72, 0.71, 
    0.75, 0.74, 0.72, 0.72, 0.69, 0.71, 0.71, 0.71, 0.69, 0.72, 0.76, 0.72, 
    0.73, 0.71, 0.68, 0.72, 0.71, 0.67, 0.57, 0.54, 0.64, 0.59, 0.65, 0.63, 
    0.66, 0.68, 0.64, 0.71, 0.68, 0.71, 0.66, 0.66, 0.68, 0.68, 0.71, 0.76, 
    0.78, 0.77, 0.76, 0.79, 0.76, 0.68, 0.73, 0.57, 0.72, 0.63, 0.71, 0.59, 
    0.65, 0.63, 0.58, 0.59, 0.63, 0.63, 0.64, 0.66, 0.64, 0.69, 0.7, 0.76, 
    0.73, 0.77, 0.79, 0.76, 0.78, 0.83, 0.64, 0.63, 0.55, 0.56, 0.56, 0.56, 
    0.57, 0.57, 0.58, 0.56, 0.56, 0.59, 0.63, 0.64, 0.6, 0.61, 0.65, 0.61, 
    0.63, 0.63, 0.63, 0.61, 0.59, 0.59, 0.63, 0.68, 0.72, 0.67, 0.61, 0.69, 
    0.73, 0.76, 0.72, 0.73, 0.7, 0.71, 0.72, 0.71, 0.66, 0.65, 0.66, 0.68, 
    0.7, 0.73, 0.73, 0.69, 0.7, 0.73, 0.71, 0.72, 0.67, 0.69, 0.68, 0.69, 
    0.69, 0.69, 0.65, 0.66, 0.7, 0.66, 0.7, 0.72, 0.67, 0.67, 0.75, 0.68, 
    0.69, 0.68, 0.67, 0.68, 0.69, 0.67, 0.65, 0.65, 0.68, 0.62, 0.66, 0.68, 
    0.66, 0.69, 0.68, 0.7, 0.68, 0.68, 0.7, 0.76, 0.73, 0.72, 0.72, 0.73, 
    0.73, 0.71, 0.71, 0.67, 0.66, 0.64, 0.63, 0.62, 0.6, 0.67, 0.64, 0.6, 
    0.62, 0.68, 0.73, 0.72, 0.73, 0.72, 0.74, 0.71, 0.71, 0.64, 0.68, 0.73, 
    0.75, 0.74, 0.75, 0.75, 0.75, 0.75, 0.73, 0.73, 0.8, 0.79, 0.77, 0.77, 
    0.72, 0.72, 0.73, 0.72, 0.68, 0.64, 0.67, 0.67, 0.68, 0.56, 0.45, 0.5, 
    0.64, 0.57, 0.51, 0.49, 0.46, 0.45, 0.44, 0.41, 0.47, 0.52, 0.56, 0.57, 
    0.61, 0.58, 0.58, 0.59, 0.56, 0.61, 0.61, 0.59, 0.53, 0.55, 0.53, 0.58, 
    0.58, 0.68, 0.67, 0.68, 0.62, 0.68, 0.73, 0.75, 0.77, 0.8, 0.81, 0.83, 
    0.86, 0.84, 0.82, 0.84, 0.89, 0.9, 0.78, 0.81, 0.8, 0.82, 0.82, 0.83, 
    0.81, 0.81, 0.8, 0.79, 0.8, 0.87, 0.88, 0.89, 0.89, 0.83, 0.8, 0.81, 
    0.77, 0.76, 0.75, 0.78, 0.71, 0.7, 0.66, 0.66, 0.6, 0.61, 0.63, 0.64, 
    0.63, 0.67, 0.6, 0.64, 0.63, 0.6, 0.58, 0.59, 0.53, 0.51, 0.54, 0.52, 
    0.48, 0.5, 0.47, 0.47, 0.46, 0.47, 0.52, 0.57, 0.6, 0.61, 0.59, 0.64, 
    0.63, 0.64, 0.64, 0.57, 0.57, 0.61, 0.6, 0.66, 0.61, 0.54, 0.61, 0.61, 
    0.66, 0.71, 0.68, 0.67, 0.67, 0.7, 0.73, 0.71, 0.76, 0.75, 0.75, 0.77, 
    0.81, 0.84, 0.83, 0.81, 0.72, 0.67, 0.71, 0.71, 0.69, 0.7, 0.72, 0.67, 
    0.68, 0.63, 0.6, 0.56, 0.53, 0.59, 0.63, 0.62, 0.66, 0.57, 0.48, 0.51, 
    0.43, 0.41, 0.43, 0.41, 0.41, 0.42, 0.5, 0.46, 0.45, 0.45, 0.46, 0.43, 
    0.44, 0.44, 0.46, 0.44, 0.46, 0.45, 0.47, 0.47, 0.5, 0.47, 0.53, 0.5, 
    0.56, 0.52, 0.54, 0.53, 0.6, 0.63, 0.66, 0.65, 0.67, 0.64, 0.68, 0.63, 
    0.65, 0.66, 0.68, 0.7, 0.72, 0.73, 0.68, 0.67, 0.7, 0.72, 0.7, 0.71, 0.7, 
    0.7, 0.66, 0.7, 0.71, 0.74, 0.67, 0.65, 0.63, 0.59, 0.58, 0.63, 0.62, 
    0.61, 0.74, 0.75, 0.8, 0.78, 0.75, 0.76, 0.77, 0.78, 0.8, 0.77, 0.79, 
    0.78, 0.79, 0.82, 0.82, 0.82, 0.81, 0.81, 0.81, 0.8, 0.79, 0.79, 0.79, 
    0.78, 0.76, 0.76, 0.77, 0.71, 0.65, 0.62, 0.63, 0.67, 0.59, 0.63, 0.66, 
    0.63, 0.62, 0.62, 0.67, 0.69, 0.69, 0.69, 0.71, 0.68, 0.64, 0.65, 0.66, 
    0.63, 0.63, 0.66, 0.68, 0.67, 0.67, 0.62, 0.65, 0.7, 0.67, 0.68, 0.73, 
    0.72, 0.75, 0.74, 0.77, 0.78, 0.74, 0.75, 0.76, 0.81, 0.79, 0.77, 0.77, 
    0.77, 0.75, 0.77, 0.64, 0.64, 0.62, 0.56, 0.54, 0.56, 0.56, 0.6, 0.64, 
    0.64, 0.67, 0.71, 0.7, 0.7, 0.64, 0.69, 0.62, 0.61, 0.59, 0.55, 0.55, 
    0.6, 0.53, 0.54, 0.56, 0.54, 0.55, 0.57, 0.57, 0.51, 0.54, 0.58, 0.44, 
    0.46, 0.54, 0.58, 0.56, 0.54, 0.56, 0.59, 0.58, 0.61, 0.65, 0.65, 0.65, 
    0.59, 0.57, 0.57, 0.57, 0.53, 0.57, 0.53, 0.57, 0.54, 0.52, 0.51, 0.51, 
    0.87, 0.53, 0.54, 0.57, 0.54, 0.55, 0.52, 0.54, 0.57, 0.56, 0.53, 0.53, 
    0.58, 0.59, 0.61, 0.64, 0.63, 0.65, 0.63, 0.67, 0.69, 0.68, 0.71, 0.66, 
    0.73, 0.74, 0.75, 0.77, 0.79, 0.8, 0.8, 0.81, 0.84, 0.85, 0.8, 0.78, 
    0.76, 0.77, 0.76, 0.76, 0.77, 0.75, 0.76, 0.76, 0.77, 0.87, 0.9, 0.87, 
    0.88, 0.85, 0.89, 0.86, 0.86, 0.84, 0.85, 0.9, 0.92, 0.92, 0.94, 0.94, 
    0.93, 0.93, 0.92, 0.91, 0.92, 0.93, 0.94, 0.91, 0.92, 0.95, 0.95, 0.9, 
    0.88, 0.85, 0.79, 0.79, 0.79, 0.76, 0.71, 0.71, 0.71, 0.66, 0.67, 0.63, 
    0.65, 0.57, 0.52, 0.52, 0.55, 0.54, 0.54, 0.53, 0.57, 0.55, 0.56, 0.56, 
    0.59, 0.54, 0.58, 0.58, 0.59, 0.6, 0.61, 0.58, 0.66, 0.67, 0.7, 0.68, 
    0.68, 0.72, 0.77, 0.86, 0.93, 0.94, 0.89, 0.82, 0.88, 0.91, 0.93, 0.89, 
    0.77, 0.74, 0.69, 0.68, 0.63, 0.62, 0.61, 0.61, 0.66, 0.67, 0.64, 0.67, 
    0.65, 0.68, 0.68, 0.68, 0.74, 0.7, 0.71, 0.73, 0.65, 0.7, 0.68, 0.66, 
    0.71, 0.69, 0.68, 0.7, 0.68, 0.7, 0.72, 0.7, 0.7, 0.74, 0.7, 0.69, 0.7, 
    0.71, 0.66, 0.66, 0.65, 0.65, 0.64, 0.63, 0.64, 0.68, 0.64, 0.64, 0.62, 
    0.65, 0.65, 0.64, 0.62, 0.62, 0.6, 0.63, 0.56, 0.56, 0.56, 0.64, 0.64, 
    0.63, 0.62, 0.59, 0.65, 0.62, 0.57, 0.47, 0.45, 0.48, 0.51, 0.52, 0.57, 
    0.56, 0.51, 0.53, 0.54, 0.57, 0.52, 0.46, 0.48, 0.56, 0.59, 0.63, 0.58, 
    0.58, 0.61, 0.63, 0.62, 0.63, 0.61, 0.62, 0.65, 0.63, 0.63, 0.64, 0.64, 
    0.65, 0.67, 0.7, 0.69, 0.7, 0.74, 0.64, 0.67, 0.58, 0.61, 0.7, 0.71, 
    0.71, 0.75, 0.71, 0.72, 0.72, 0.77, 0.71, 0.62, 0.61, 0.62, 0.65, 0.66, 
    0.64, 0.56, 0.58, 0.67, 0.63, 0.58, 0.65, 0.61, 0.6, 0.6, 0.62, 0.63, 
    0.67, 0.87, 0.87, 0.74, 0.77, 0.76, 0.83, 0.92, 0.94, 0.9, 0.71, 0.64, 
    0.6, 0.6, 0.6, 0.59, 0.9, 0.81, 0.82, 0.84, 0.89, 0.78, 0.84, 0.89, 0.88, 
    0.82, 0.78, 0.77, 0.75, 0.77, 0.74, 0.67, 0.82, 0.71, 0.64, 0.64, 0.78, 
    0.66, 0.7, 0.71, 0.72, 0.71, 0.74, 0.74, 0.73, 0.69, 0.8, 0.78, 0.76, 
    0.78, 0.71, 0.73, 0.8, 0.82, 0.86, 0.86, 0.85, 0.75, 0.76, 0.77, 0.79, 
    0.78, 0.83, 0.91, 0.75, 0.71, 0.72, 0.67, 0.68, 0.65, 0.66, 0.61, 0.55, 
    0.53, 0.56, 0.55, 0.51, 0.55, 0.51, 0.52, 0.54, 0.55, 0.55, 0.55, 0.57, 
    0.63, 0.65, 0.65, 0.66, 0.68, 0.69, 0.69, 0.8, 0.8, 0.82, 0.67, 0.66, 
    0.65, 0.64, 0.63, 0.65, 0.64, 0.67, 0.66, 0.65, 0.65, 0.69, 0.59, 0.66, 
    0.68, 0.67, 0.63, 0.6, 0.65, 0.55, 0.54, 0.63, 0.66, 0.68, 0.68, 0.67, 
    0.61, 0.66, 0.65, 0.68, 0.67, 0.85, 0.95, 0.93, 0.86, 0.89, 0.94, 0.93, 
    0.94, 0.92, 0.9, 0.91, 0.89, 0.87, 0.9, 0.91, 0.89, 0.85, 0.78, 0.72, 
    0.7, 0.65, 0.62, 0.6, 0.6, 0.65, 0.67, 0.6, 0.62, 0.77, 0.84, 0.7, 0.68, 
    0.68, 0.66, 0.69, 0.63, 0.64, 0.58, 0.59, 0.54, 0.54, 0.52, 0.51, 0.54, 
    0.54, 0.56, 0.58, 0.57, 0.66, 0.67, 0.67, 0.67, 0.69, 0.69, 0.7, 0.66, 
    0.66, 0.66, 0.66, 0.67, 0.69, 0.7, 0.84, 0.87, 0.87, 0.84, 0.7, 0.61, 
    0.57, 0.57, 0.49, 0.58, 0.52, 0.57, 0.65, 0.61, 0.64, 0.62, 0.63, 0.64, 
    0.63, 0.63, 0.63, 0.64, 0.66, 0.7, 0.7, 0.61, 0.61, 0.64, 0.64, 0.65, 
    0.64, 0.68, 0.66, 0.68, 0.69, 0.66, 0.73, 0.76, 0.75, 0.73, 0.74, 0.75, 
    0.77, 0.86, 0.9, 0.92, 0.93, 0.89, 0.86, 0.83, 0.84, 0.9, 0.94, 0.86, 
    0.96, 0.9, 0.91, 0.82, 0.73, 0.8, 0.89, 0.97, 0.98, 0.98, 0.95, 0.93, 
    0.9, 0.99, 0.82, 0.76, 0.8, 0.8, 0.78, 0.74, 0.76, 0.81, 0.79, 0.74, 
    0.67, 0.71, 0.64, 0.67, 0.66, 0.6, 0.64, 0.57, 0.52, 0.56, 0.57, 0.54, 
    0.56, 0.59, 0.61, 0.57, 0.57, 0.55, 0.53, 0.56, 0.53, 0.57, 0.6, 0.54, 
    0.52, 0.52, 0.47, 0.53, 0.51, 0.51, 0.55, 0.57, 0.55, 0.57, 0.61, 0.64, 
    0.61, 0.66, 0.64, 0.67, 0.67, 0.66, 0.69, 0.7, 0.69, 0.64, 0.6, 0.59, 
    0.58, 0.63, 0.64, 0.63, 0.59, 0.58, 0.6, 0.54, 0.52, 0.51, 0.5, 0.53, 
    0.59, 0.62, 0.64, 0.63, 0.58, 0.6, 0.62, 0.62, 0.65, 0.62, 0.61, 0.61, 
    0.62, 0.67, 0.64, 0.62, 0.59, 0.54, 0.49, 0.5, 0.51, 0.53, 0.53, 0.56, 
    0.57, 0.56, 0.51, 0.57, 0.59, 0.59, 0.6, 0.57, 0.59, 0.59, 0.59, 0.6, 
    0.63, 0.67, 0.71, 0.74, 0.74, 0.74, 0.76, 0.76, 0.81, 0.75, 0.75, 0.76, 
    0.78, 0.79, 0.75, 0.74, 0.76, 0.79, 0.79, 0.79, 0.74, 0.75, 0.76, 0.75, 
    0.76, 0.77, 0.8, 0.83, 0.9, 0.89, 0.92, 0.88, 0.88, 0.85, 0.85, 0.8, 
    0.84, 0.95, 0.95, 0.98, 1, 1, 0.96, 0.86, 0.86, 0.83, 0.92, 0.77, 0.65, 
    0.63, 0.67, 0.66, 0.73, 0.74, 0.79, 0.8, 0.78, 0.82, 0.9, 0.87, 0.83, 
    0.85, 0.82, 0.77, 0.76, 0.73, 0.7, 0.74, 0.7, 0.66, 0.67, 0.68, 0.68, 
    0.65, 0.69, 0.61, 0.73, 0.8, 0.76, 0.62, 0.56, 0.52, 0.55, 0.52, 0.5, 
    0.43, 0.57, 0.57, 0.58, 0.59, 0.6, 0.49, 0.63, 0.76, 0.73, 0.72, 0.69, 
    0.72, 0.66, 0.58, 0.57, 0.55, 0.64, 0.65, 0.73, 0.62, 0.64, 0.7, 0.71, 
    0.66, 0.6, 0.55, 0.53, 0.63, 0.54, 0.6, 0.61, 0.65, 0.63, 0.6, 0.55, 
    0.55, 0.55, 0.54, 0.57, 0.56, 0.54, 0.58, 0.62, 0.53, 0.51, 0.54, 0.56, 
    0.57, 0.51, 0.52, 0.57, 0.6, 0.59, 0.59, 0.62, 0.6, 0.62, 0.6, 0.62, 
    0.63, 0.61, 0.59, 0.61, 0.63, 0.63, 0.67, 0.63, 0.61, 0.62, 0.64, 0.68, 
    0.69, 0.66, 0.64, 0.64, 0.6, 0.63, 0.66, 0.66, 0.65, 0.6, 0.63, 0.66, 
    0.62, 0.6, 0.62, 0.58, 0.61, 0.62, 0.62, 0.62, 0.62, 0.62, 0.64, 0.61, 
    0.6, 0.59, 0.59, 0.56, 0.59, 0.58, 0.57, 0.59, 0.6, 0.61, 0.62, 0.62, 
    0.6, 0.63, 0.66, 0.66, 0.65, 0.63, 0.6, 0.62, 0.61, 0.61, 0.61, 0.6, 
    0.59, 0.61, 0.59, 0.63, 0.64, 0.6, 0.63, 0.61, 0.6, 0.6, 0.61, 0.61, 
    0.63, 0.59, 0.59, 0.57, 0.55, 0.56, 0.54, 0.54, 0.51, 0.52, 0.54, 0.51, 
    0.52, 0.48, 0.43, 0.41, 0.42, 0.44, 0.45, 0.48, 0.4, 0.4, 0.39, 0.4, 
    0.42, 0.45, 0.46, 0.44, 0.5, 0.57, 0.72, 0.83, 0.67, 0.45, 0.45, 0.47, 
    0.44, 0.44, 0.44, 0.54, 0.5, 0.52, 0.56, 0.59, 0.56, 0.65, 0.58, 0.61, 
    0.57, 0.54, 0.52, 0.52, 0.5, 0.5, 0.46, 0.51, 0.55, 0.57, 0.54, 0.53, 
    0.53, 0.53, 0.52, 0.53, 0.55, 0.6, 0.58, 0.56, 0.53, 0.55, 0.58, 0.55, 
    0.57, 0.55, 0.62, 0.59, 0.6, 0.6, 0.64, 0.59, 0.61, 0.59, 0.56, 0.51, 
    0.56, 0.55, 0.54, 0.54, 0.54, 0.57, 0.63, 0.59, 0.64, 0.59, 0.57, 0.59, 
    0.63, 0.59, 0.59, 0.59, 0.56, 0.56, 0.54, 0.54, 0.57, 0.59, 0.6, 0.62, 
    0.61, 0.62, 0.65, 0.64, 0.63, 0.62, 0.62, 0.6, 0.59, 0.6, 0.6, 0.59, 
    0.58, 0.6, 0.6, 0.57, 0.59, 0.59, 0.59, 0.61, 0.6, 0.63, 0.62, 0.62, 
    0.66, 0.67, 0.65, 0.64, 0.6, 0.59, 0.59, 0.55, 0.56, 0.55, 0.57, 0.59, 
    0.56, 0.54, 0.52, 0.5, 0.52, 0.45, 0.58, 0.55, 0.51, 0.56, 0.71, 0.63, 
    0.66, 0.65, 0.61, 0.55, 0.5, 0.57, 0.6, 0.59, 0.58, 0.63, 0.66, 0.66, 
    0.62, 0.63, 0.62, 0.61, 0.63, 0.7, 0.64, 0.64, 0.58, 0.64, 0.64, 0.62, 
    0.8, 0.57, 0.56, 0.58, 0.61, 0.62, 0.63, 0.64, 0.63, 0.62, 0.62, 0.62, 
    0.62, 0.62, 0.6, 0.64, 0.72, 0.64, 0.62, 0.62, 0.75, 0.73, 0.63, 0.65, 
    0.6, 0.63, 0.53, 0.5, 0.53, 0.56, 0.58, 0.57, 0.58, 0.55, 0.6, 0.6, 0.61, 
    0.6, 0.57, 0.62, 0.68, 0.66, 0.63, 0.66, 0.66, 0.69, 0.67, 0.66, 0.67, 
    0.7, 0.66, 0.69, 0.7, 0.66, 0.62, 0.66, 0.72, 0.74, 0.78, 0.79, 0.79, 
    0.79, 0.8, 0.76, 0.77, 0.76, 0.75, 0.76, 0.75, 0.77, 0.77, 0.8, 0.82, 
    0.81, 0.85, 0.79, 0.71, 0.78, 0.81, 0.76, 0.73, 0.79, 0.74, 0.74, 0.68, 
    0.64, 0.64, 0.64, 0.62, 0.59, 0.7, 0.67, 0.63, 0.67, 0.67, 0.7, 0.64, 
    0.58, 0.56, 0.69, 0.58, 0.61, 0.6, 0.51, 0.44, 0.45, 0.45, 0.45, 0.45, 
    0.47, 0.52, 0.51, 0.48, 0.43, 0.45, 0.5, 0.47, 0.64, 0.51, 0.49, 0.46, 
    0.5, 0.48, 0.45, 0.51, 0.51, 0.5, 0.46, 0.48, 0.45, 0.44, 0.47, 0.51, 
    0.57, 0.52, 0.6, 0.57, 0.57, 0.58, 0.59, 0.61, 0.6, 0.58, 0.62, 0.61, 
    0.6, 0.52, 0.53, 0.58, 0.66, 0.65, 0.67, 0.67, 0.67, 0.67, 0.75, 0.89, 
    0.95, 0.93, 0.91, 0.9, 0.85, 0.8, 0.83, 0.78, 0.76, 0.73, 0.73, 0.72, 
    0.76, 0.74, 0.76, 0.78, 0.86, 0.87, 0.87, 0.86, 0.9, 0.91, 0.98, 0.87, 
    0.79, 0.72, 0.68, 0.68, 0.68, 0.69, 0.77, 0.78, 0.74, 0.68, 0.78, 0.86, 
    0.82, 0.84, 0.83, 0.87, 0.85, 0.85, 0.79, 0.75, 0.8, 0.73, 0.79, 0.81, 
    0.77, 0.79, 0.78, 0.79, 0.77, 0.76, 0.68, 0.73, 0.73, 0.73, 0.75, 0.73, 
    0.73, 0.71, 0.65, 0.71, 0.69, 0.64, 0.69, 0.69, 0.69, 0.71, 0.72, 0.69, 
    0.63, 0.56, 0.64, 0.56, 0.53, 0.64, 0.67, 0.93, 0.78, 0.81, 0.8, 0.75, 
    0.7, 0.89, 0.72, 0.72, 0.82, 0.71, 0.69, 0.68, 0.67, 0.65, 0.69, 0.79, 
    0.67, 0.79, 0.74, 0.72, 0.74, 0.92, 1, 0.92, 0.89, 0.87, 0.87, 0.82, 
    0.85, 0.83, 0.77, 0.78, 0.91, 0.86, 0.77, 0.82, 0.78, 0.75, 0.76, 0.75, 
    0.75, 0.75, 0.75, 0.76, 0.75, 0.7, 0.74, 0.78, 0.77, 0.78, 0.75, 0.65, 
    0.72, 0.65, 0.67, 0.66, 0.75, 0.59, 0.68, 0.67, 0.62, 0.69, 0.7, 0.72, 
    0.79, 0.76, 0.87, 0.97, 0.93, 0.95, 1, 0.99, 1, 0.99, 0.99, 1, 0.99, 
    0.99, 0.99, 1, 1, 1, 1, 0.98, 0.99, 0.98, 0.99, 0.99, 1, 0.99, 0.89, 
    0.89, 0.88, 0.88, 0.87, 0.92, 0.81, 0.83, 0.84, 0.86, 0.79, 0.76, 0.79, 
    0.76, 0.8, 0.8, 0.78, 0.78, 0.77, 0.78, 0.78, 0.76, 0.78, 0.78, 0.77, 
    0.75, 0.68, 0.78, 0.74, 0.77, 0.71, 0.75, 0.77, 0.8, 0.76, 0.68, 0.68, 
    0.72, 0.56, 0.72, 0.64, 0.68, 0.71, 0.72, 0.72, 0.69, 0.61, 0.57, 0.56, 
    0.54, 0.64, 0.57, 0.66, 0.59, 0.61, 0.6, 0.59, 0.54, 0.54, 0.53, 0.55, 
    0.56, 0.59, 0.55, 0.55, 0.59, 0.58, 0.59, 0.52, 0.53, 0.57, 0.55, 0.55, 
    0.58, 0.57, 0.57, 0.56, 0.57, 0.6, 0.61, 0.6, 0.61, 0.57, 0.58, 0.57, 
    0.55, 0.53, 0.51, 0.49, 0.47, 0.47, 0.47, 0.46, 0.48, 0.47, 0.48, 0.46, 
    0.48, 0.46, 0.46, 0.44, 0.44, 0.46, 0.46, 0.47, 0.47, 0.46, 0.49, 0.48, 
    0.48, 0.52, 0.52, 0.54, 0.49, 0.48, 0.48, 0.48, 0.51, 0.53, 0.52, 0.49, 
    0.54, 0.59, 0.58, 0.61, 0.59, 0.57, 0.59, 0.58, 0.59, 0.61, 0.62, 0.67, 
    0.6, 0.59, 0.64, 0.62, 0.62, 0.61, 0.58, 0.59, 0.58, 0.6, 0.59, 0.57, 
    0.58, 0.56, 0.55, 0.54, 0.56, 0.55, 0.53, 0.54, 0.52, 0.52, 0.5, 0.51, 
    0.54, 0.53, 0.56, 0.56, 0.46, 0.46, 0.43, 0.41, 0.4, 0.36, 0.32, 0.45, 
    0.3, 0.3, 0.34, 0.41, 0.47, 0.51, 0.54, 0.53, 0.53, 0.55, 0.57, 0.55, 
    0.54, 0.53, 0.61, 0.63, 0.58, 0.57, 0.53, 0.55, 0.57, 0.58, 0.61, 0.61, 
    0.57, 0.55, 0.55, 0.56, 0.56, 0.56, 0.52, 0.55, 0.59, 0.56, 0.57, 0.59, 
    0.58, 0.57, 0.55, 0.53, 0.53, 0.55, 0.61, 0.57, 0.63, 0.57, 0.62, 0.64, 
    0.62, 0.65, 0.65, 0.62, 0.6, 0.63, 0.59, 0.58, 0.62, 0.6, 0.63, 0.54, 
    0.57, 0.53, 0.57, 0.6, 0.56, 0.56, 0.53, 0.59, 0.58, 0.57, 0.5, 0.6, 
    0.59, 0.56, 0.53, 0.58, 0.51, 0.63, 0.59, 0.82, 0.89, 0.88, 0.85, 0.86, 
    0.83, 0.86, 0.88, 0.88, 0.89, 0.89, 0.89, 0.83, 0.72, 0.68, 0.68, 0.63, 
    0.65, 0.7, 0.68, 0.64, 0.69, 0.73, 0.7, 0.69, 0.71, 0.69, 0.74, 0.76, 
    0.78, 0.88, 0.91, 0.94, 0.93, 0.93, 0.92, 0.95, 0.93, 0.93, 0.97, 0.99, 
    0.99, 0.99, 0.99, 1, 0.91, 0.99, 0.95, 0.99, 0.85, 0.84, 0.82, 0.74, 
    0.72, 0.74, 0.85, 0.83, 0.88, 0.8, 0.83, 0.78, 0.77, 0.81, 0.82, 0.84, 
    0.93, 0.98, 0.94, 0.99, 0.94, 0.99, 0.99, 0.95, 0.99, 0.97, 0.97, 0.88, 
    0.84, 0.85, 0.89, 0.86, 0.83, 0.71, 0.72, 0.82, 0.74, 0.72, 0.71, 0.75, 
    0.68, 0.75, 0.68, 0.72, 0.73, 0.72, 0.69, 0.67, 0.68, 0.67, 0.66, 0.61, 
    0.58, 0.59, 0.58, 0.62, 0.6, 0.57, 0.62, 0.61, 0.59, 0.69, 0.72, 0.67, 
    0.7, 0.69, 0.68, 0.66, 0.64, 0.64, 0.66, 0.69, 0.61, 0.67, 0.66, 0.57, 
    0.53, 0.56, 0.63, 0.63, 0.64, 0.67, 0.58, 0.67, 0.59, 0.62, 0.6, 0.51, 
    0.63, 0.51, 0.59, 0.54, 0.49, 0.48, 0.51, 0.52, 0.54, 0.53, 0.53, 0.56, 
    0.56, 0.54, 0.59, 0.6, 0.58, 0.57, 0.58, 0.57, 0.59, 0.59, 0.65, 0.6, 
    0.61, 0.6, 0.62, 0.66, 0.62, 0.68, 0.67, 0.7, 0.7, 0.73, 0.69, 0.73, 
    0.74, 0.72, 0.69, 0.74, 0.73, 0.71, 0.72, 0.8, 0.69, 0.7, 0.67, 0.67, 
    0.65, 0.66, 0.74, 0.71, 0.7, 0.71, 0.62, 0.55, 0.68, 0.59, 0.6, 0.61, 
    0.61, 0.58, 0.62, 0.6, 0.56, 0.6, 0.61, 0.6, 0.56, 0.56, 0.55, 0.52, 
    0.53, 0.57, 0.51, 0.51, 0.43, 0.67, 0.54, 0.52, 0.51, 0.56, 0.52, 0.53, 
    0.51, 0.56, 0.58, 0.63, 0.57, 0.61, 0.69, 0.64, 0.74, 0.77, 0.81, 0.84, 
    0.9, 0.93, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.99, 0.93, 0.81, 0.82, 
    0.79, 0.8, 0.94, 0.81, 0.87, 0.91, 0.91, 0.95, 0.91, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.84, 0.83, 0.81, 0.84, 0.88, 0.77, 0.85, 0.84, 0.81, 0.79, 
    0.78, 0.84, 0.86, 0.88, 0.9, 0.93, 0.92, 0.93, 0.91, 0.93, 0.93, 0.91, 
    0.87, 0.84, 0.82, 0.8, 0.79, 0.8, 0.81, 0.81, 0.79, 0.77, 0.74, 0.71, 
    0.74, 0.79, 0.83, 0.8, 0.8, 0.85, 0.83, 0.84, 0.81, 0.82, 0.85, 0.82, 
    0.84, 0.83, 0.8, 0.73, 0.72, 0.84, 0.83, 0.75, 0.71, 0.86, 0.79, 0.78, 
    0.79, 0.87, 0.81, 0.85, 0.89, 0.86, 0.89, 0.88, 0.82, 0.84, 0.85, 0.84, 
    0.85, 0.82, 0.83, 0.85, 0.78, 0.64, 0.7, 0.65, 0.66, 0.67, 0.69, 0.71, 
    0.74, 0.71, 0.76, 0.82, 0.83, 0.92, 0.86, 0.79, 0.84, 0.8, 0.85, 0.83, 
    0.76, 0.78, 0.85, 0.81, 0.82, 0.82, 0.78, 0.79, 0.76, 0.85, 0.85, 0.86, 
    0.85, 0.87, 0.85, 0.83, 0.86, 0.9, 0.88, 0.85, 0.96, 0.95, 0.94, 0.9, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 
    0.99, 0.99, 1, 0.72, 0.74, 0.79, 0.79, 0.88, 0.83, 0.75, 0.73, 0.67, 
    0.67, 0.68, 0.66, 0.72, 0.79, 0.82, 0.82, 0.87, 0.96, 0.81, 0.8, 0.84, 
    0.82, 0.84, 0.87, 0.83, 0.8, 0.82, 0.78, 0.76, 0.93, 0.84, 0.83, 0.85, 
    0.9, 0.89, 0.99, 0.88, 0.89, 0.89, 0.89, 0.94, 0.93, 0.9, 0.99, 0.86, 
    0.72, 0.75, 0.78, 0.78, 0.78, 0.86, 0.76, 0.8, 0.79, 0.86, 0.86, 0.83, 
    0.7, 0.67, 0.71, 0.71, 0.71, 0.7, 0.67, 0.63, 0.72, 0.76, 0.77, 0.79, 
    0.8, 0.76, 0.75, 0.84, 0.73, 0.86, 0.86, 0.91, 0.75, 0.78, 0.78, 0.78, 
    0.78, 0.86, 0.8, 0.85, 0.79, 0.83, 0.8, 0.82, 0.83, 0.81, 0.83, 0.81, 
    0.61, 0.78, 0.72, 0.77, 0.74, 0.79, 0.79, 0.85, 0.92, 0.96, 0.99, 0.99, 
    0.99, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.98, 0.9, 0.81, 0.8, 0.75, 
    0.84, 0.83, 0.78, 0.73, 0.78, 0.76, 0.71, 0.7, 0.64, 0.63, 0.61, 0.82, 
    0.71, 0.81, 0.73, 0.68, 0.7, 0.72, 0.74, 0.66, 0.66, 0.69, 0.66, 0.65, 
    0.7, 0.84, 0.75, 0.69, 0.9, 0.86, 0.83, 0.92, 0.99, 1, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.87, 0.97, 0.93, 
    0.9, 0.9, 0.94, 0.95, 0.98, 1, 0.96, 0.99, 0.99, 0.91, 0.88, 0.96, 0.85, 
    0.97, 0.97, 0.96, 0.99, 0.99, 0.96, 0.97, 0.96, 1, 0.99, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 1, 0.99, 
    0.99, 0.99, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.91, 0.96, 0.99, 0.93, 0.99, 
    1, 0.99, 0.97, 0.99, 0.99, 1, 0.99, 0.97, 0.91, 0.85, 0.93, 0.96, 0.83, 
    0.85, 0.82, 0.82, 0.73, 0.74, 0.75, 0.74, 0.72, 0.6, 0.74, 0.63, 0.73, 
    0.63, 0.61, 0.62, 0.66, 0.62, 0.62, 0.73, 0.69, 0.65, 0.74, 0.7, 0.82, 
    0.79, 0.77, 0.8, 0.75, 0.79, 0.75, 0.73, 0.74, 0.75, 0.77, 0.75, 0.77, 
    0.74, 0.74, 0.77, 0.79, 0.81, 0.73, 0.79, 0.8, 0.76, 0.76, 0.74, 0.75, 
    0.79, 0.74, 0.77, 0.71, 0.68, 0.74, 0.71, 0.72, 0.72, 0.69, 0.71, 0.71, 
    0.76, 0.74, 0.66, 0.66, 0.69, 0.66, 0.72, 0.8, 0.81, 0.75, 0.78, 0.72, 
    0.71, 0.75, 0.74, 0.78, 0.81, 0.84, 0.82, 0.86, 0.9, 0.88, 0.84, 0.8, 
    0.76, 0.71, 0.81, 0.76, 0.79, 0.78, 0.85, 0.92, 0.9, 0.86, 0.86, 0.86, 
    0.9, 0.9, 0.9, 0.9, 0.88, 0.93, 0.95, 0.95, 0.9, 0.92, 0.94, 0.98, 0.99, 
    0.99, 1, 0.99, 0.99, 0.97, 0.86, 0.94, 0.87, 0.81, 0.81, 0.78, 0.86, 
    0.94, 0.93, 0.93, 0.92, 0.99, 0.99, 0.99, 0.98, 0.97, 0.99, 0.91, 0.88, 
    0.95, 0.95, 0.99, 0.99, 0.99, 0.99, 0.98, 1, 1, 0.99, 0.99, 0.99, 0.91, 
    0.95, 0.96, 0.95, 0.93, 0.97, 0.99, 1, 0.99, 0.92, 0.9, 1, 1, 0.95, 0.99, 
    1, 0.94, 0.97, 0.99, 0.95, 0.94, 0.91, 0.84, 0.83, 0.76, 0.75, 0.87, 
    0.84, 0.82, 0.82, 0.8, 0.76, 0.71, 0.73, 0.62, 0.7, 0.65, 0.76, 0.7, 
    0.75, 0.66, 0.65, 0.79, 0.76, 0.66, 0.69, 0.73, 0.8, 0.78, 0.77, 0.72, 
    0.71, 0.77, 0.81, 0.84, 0.79, 0.74, 0.74, 0.76, 0.74, 0.78, 0.74, 0.82, 
    0.78, 0.78, 0.82, 0.73, 0.82, 0.85, 0.76, 0.82, 0.78, 0.77, 0.78, 0.83, 
    0.94, 0.82, 0.82, 0.82, 0.88, 0.9, 0.81, 0.89, 0.94, 0.85, 0.94, 0.93, 
    0.89, 0.97, 0.88, 0.94, 0.91, 0.84, 0.87, 0.85, 0.85, 0.96, 0.99, 0.88, 
    0.86, 0.7, 0.79, 0.79, 0.76, 0.69, 0.7, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.95, 0.91, 0.98, 1, 0.96, 0.81, 0.89, 0.84, 0.85, 0.91, 0.84, 0.81, 
    0.77, 0.86, 0.75, 0.8, 0.84, 0.8, 0.76, 0.76, 0.76, 0.82, 0.79, 0.78, 
    0.73, 0.72, 0.7, 0.76, 0.76, 0.72, 0.69, 0.74, 0.77, 0.77, 0.75, 0.73, 
    0.79, 0.77, 0.73, 0.79, 0.88, 0.79, 0.78, 0.73, 0.76, 0.74, 0.69, 0.68, 
    0.74, 0.75, 0.81, 0.78, 0.77, 0.7, 0.67, 0.76, 0.77, 0.66, 0.73, 0.72, 
    0.73, 0.72, 0.7, 0.71, 0.73, 0.76, 0.71, 0.76, 0.7, 0.68, 0.74, 0.77, 
    0.7, 0.65, 0.69, 0.7, 0.82, 0.71, 0.66, 0.65, 0.77, 0.79, 0.8, 0.79, 0.7, 
    0.61, 0.62, 0.65, 0.65, 0.63, 0.65, 0.67, 0.6, 0.62, 0.66, 0.7, 0.73, 
    0.74, 0.82, 0.72, 0.82, 0.84, 0.77, 0.73, 0.82, 0.71, 0.68, 0.65, 0.67, 
    0.65, 0.63, 0.67, 0.74, 0.77, 0.7, 0.72, 0.85, 0.75, 0.84, 0.79, 0.87, 
    0.77, 0.76, 0.78, 0.85, 0.83, 0.82, 0.96, 0.99, 0.99, 0.99, 0.99, 0.95, 
    1, 0.99, 0.91, 0.99, 1, 1, 0.99, 1, 1, 1, 0.99, 0.99, 0.91, 0.88, 0.91, 
    0.95, 0.9, 0.85, 0.82, 0.71, 0.72, 0.69, 0.69, 0.7, 0.68, 0.73, 0.74, 
    0.83, 0.81, 0.77, 0.72, 0.75, 0.8, 0.76, 0.74, 0.73, 0.75, 0.78, 0.81, 
    0.81, 0.76, 0.75, 0.79, 0.76, 0.79, 0.76, 0.78, 0.74, 0.78, 0.81, 0.82, 
    0.82, 0.87, 0.82, 0.86, 0.86, 0.78, 0.78, 0.8, 0.82, 0.74, 0.72, 0.7, 
    0.65, 0.66, 0.68, 0.66, 0.7, 0.67, 0.82, 0.79, 0.79, 0.83, 0.84, 0.81, 
    0.81, 0.79, 0.88, 0.89, 0.88, 0.78, 0.78, 0.84, 0.87, 0.74, 0.7, 0.71, 
    0.69, 0.71, 0.72, 0.73, 0.72, 0.68, 0.58, 0.57, 0.57, 0.56, 0.61, 0.62, 
    0.63, 0.64, 0.6, 0.6, 0.64, 0.63, 0.63, 0.66, 0.65, 0.69, 0.74, 0.56, 
    0.63, 0.69, 0.7, 0.68, 0.62, 0.62, 0.63, 0.63, 0.62, 0.58, 0.55, 0.57, 
    0.7, 0.65, 0.64, 0.65, 0.71, 0.68, 0.7, 0.71, 0.71, 0.71, 0.75, 0.78, 
    0.75, 0.77, 0.72, 0.77, 0.75, 0.71, 0.76, 0.75, 0.7, 0.64, 0.58, 0.58, 
    0.57, 0.59, 0.59, 0.69, 0.66, 0.7, 0.62, 0.6, 0.58, 0.61, 0.62, 0.73, 
    0.75, 0.62, 0.68, 0.67, 0.72, 0.71, 0.68, 0.7, 0.74, 0.75, 0.73, 0.66, 
    0.69, 0.66, 0.68, 0.66, 0.69, 0.72, 0.67, 0.7, 0.72, 0.73, 0.69, 0.67, 
    0.66, 0.67, 0.66, 0.67, 0.72, 0.62, 0.65, 0.66, 0.66, 0.59, 0.75, 0.59, 
    0.55, 0.65, 0.65, 0.68, 0.69, 0.73, 0.71, 0.68, 0.76, 0.75, 0.74, 0.73, 
    0.73, 0.72, 0.71, 0.71, 0.72, 0.69, 0.71, 0.76, 0.82, 0.87, 0.91, 0.85, 
    0.97, 0.99, 0.99, 0.95, 0.9, 0.87, 0.86, 0.82, 0.78, 0.83, 0.82, 0.78, 
    0.74, 0.84, 0.85, 0.82, 0.75, 0.77, 0.78, 0.76, 0.74, 0.73, 0.71, 0.73, 
    0.72, 0.7, 0.72, 0.71, 0.79, 0.76, 0.85, 0.79, 0.85, 0.88, 0.82, 0.82, 
    0.79, 0.77, 0.87, 0.9, 0.89, 0.91, 0.91, 0.84, 0.84, 0.88, 0.93, 0.95, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.96, 0.92, 0.94, 0.92, 0.9, 0.85, 0.79, 
    0.79, 0.65, 0.74, 0.66, 0.63, 0.69, 0.7, 0.73, 0.63, 0.64, 0.67, 0.7, 
    0.67, 0.62, 0.58, 0.62, 0.62, 0.61, 0.6, 0.61, 0.62, 0.62, 0.56, 0.57, 
    0.56, 0.54, 0.53, 0.59, 0.55, 0.55, 0.54, 0.55, 0.52, 0.51, 0.52, 0.52, 
    0.51, 0.51, 0.52, 0.53, 0.58, 0.52, 0.62, 0.54, 0.57, 0.58, 0.58, 0.57, 
    0.54, 0.56, 0.54, 0.58, 0.6, 0.54, 0.57, 0.58, 0.57, 0.57, 0.5, 0.54, 
    0.58, 0.55, 0.58, 0.56, 0.55, 0.57, 0.56, 0.57, 0.57, 0.58, 0.63, 0.55, 
    0.55, 0.51, 0.71, 0.63, 0.65, 0.66, 0.71, 0.71, 0.77, 0.87, 0.82, 0.83, 
    0.89, 0.84, 0.89, 0.88, 0.89, 0.9, 0.81, 0.96, 0.81, 0.83, 0.74, 0.65, 
    0.67, 0.69, 0.71, 0.66, 0.61, 0.6, 0.58, 0.67, 0.71, 0.64, 0.62, 0.73, 
    0.8, 0.77, 0.84, 0.73, 0.7, 0.62, 0.67, 0.63, 0.63, 0.62, 0.61, 0.59, 
    0.7, 0.68, 0.7, 0.78, 0.72, 0.73, 0.74, 0.81, 0.8, 0.8, 0.83, 0.81, 0.8, 
    0.52, 0.53, 0.44, 0.46, 0.44, 0.5, 0.5, 0.46, 0.46, 0.47, 0.5, 0.55, 
    0.55, 0.56, 0.6, 0.56, 0.47, 0.55, 0.57, 0.58, 0.61, 0.6, 0.59, 0.62, 
    0.62, 0.67, 0.66, 0.68, 0.66, 0.64, 0.67, 0.64, 0.64, 0.7, 0.64, 0.7, 
    0.7, 0.7, 0.74, 0.74, 0.71, 0.69, 0.66, 0.69, 0.74, 0.8, 0.88, 0.92, 
    0.94, 0.95, 0.94, 0.9, 0.89, 0.85, 0.81, 0.83, 0.88, 0.92, 0.94, 0.93, 
    0.87, 0.82, 0.92, 0.82, 0.76, 0.71, 0.74, 0.98, 0.99, 0.96, 0.92, 0.89, 
    0.8, 0.82, 0.99, 0.99, 0.99, 1, 0.89, 0.92, 0.87, 0.76, 0.74, 0.73, 0.85, 
    0.87, 0.85, 0.78, 0.68, 0.67, 0.62, 0.62, 0.63, 0.6, 0.64, 0.64, 0.63, 
    0.63, 0.68, 0.68, 0.73, 0.77, 0.7, 0.7, 0.73, 0.77, 0.75, 0.74, 0.68, 
    0.74, 0.74, 0.7, 0.75, 0.73, 0.74, 0.7, 0.76, 0.79, 0.77, 0.75, 0.76, 
    0.86, 0.93, 0.91, 0.81, 0.8, 0.81, 0.92, 0.97, 0.99, 0.99, 0.98, 0.98, 
    0.97, 0.87, 0.84, 0.75, 0.89, 0.8, 0.82, 0.88, 0.71, 0.65, 0.64, 0.74, 
    0.63, 0.72, 0.75, 0.83, 0.78, 0.79, 0.75, 0.7, 0.73, 0.74, 0.77, 0.79, 
    0.75, 0.74, 0.73, 0.69, 0.66, 0.69, 0.74, 0.74, 0.84, 0.96, 0.88, 0.99, 
    0.99, 0.83, 0.69, 0.68, 0.66, 0.7, 0.74, 0.72, 0.69, 0.66, 0.68, 0.66, 
    0.67, 0.69, 0.71, 0.72, 0.79, 0.76, 0.74, 0.68, 0.64, 0.67, 0.69, 0.65, 
    0.73, 0.67, 0.72, 0.7, 0.71, 0.77, 0.69, 0.66, 0.69, 0.73, 0.7, 0.99, 
    0.99, 1, 1, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.91, 0.93, 
    0.93, 0.82, 0.75, 0.8, 0.78, 0.79, 0.77, 0.8, 0.72, 0.71, 0.74, 0.77, 
    0.77, 0.66, 0.74, 0.71, 0.68, 0.75, 0.76, 0.79, 0.74, 0.73, 0.66, 0.62, 
    0.73, 0.81, 0.76, 0.79, 0.82, 0.79, 0.88, 0.88, 0.89, 0.92, 0.91, 0.91, 
    0.92, 0.92, 0.92, 0.97, 0.96, 0.95, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.97, 0.92, 0.91, 0.93, 0.97, 0.94, 0.91, 0.91, 0.91, 0.96, 0.83, 
    0.84, 0.77, 0.75, 0.74, 0.73, 0.68, 0.71, 0.65, 0.57, 0.6, 0.6, 0.56, 
    0.55, 0.54, 0.52, 0.59, 0.62, 0.61, 0.61, 0.62, 0.61, 0.61, 0.71, 0.66, 
    0.63, 0.65, 0.67, 0.74, 0.67, 0.69, 0.65, 0.66, 0.59, 0.65, 0.59, 0.53, 
    0.48, 0.43, 0.42, 0.39, 0.68, 0.54, 0.39, 0.42, 0.44, 0.34, 0.38, 0.38, 
    0.31, 0.38, 0.37, 0.44, 0.39, 0.38, 0.45, 0.47, 0.41, 0.44, 0.47, 0.48, 
    0.44, 0.41, 0.46, 0.56, 0.49, 0.48, 0.57, 0.47, 0.51, 0.46, 0.49, 0.51, 
    0.52, 0.53, 0.53, 0.58, 0.63, 0.63, 0.64, 0.65, 0.66, 0.69, 0.66, 0.66, 
    0.61, 0.6, 0.62, 0.6, 0.65, 0.63, 0.68, 0.68, 0.7, 0.7, 0.68, 0.68, 0.72, 
    0.71, 0.68, 0.69, 0.71, 0.72, 0.69, 0.68, 0.7, 0.72, 0.68, 0.61, 0.63, 
    0.62, 0.55, 0.68, 0.72, 0.6, 0.62, 0.64, 0.68, 0.66, 0.7, 0.59, 0.51, 
    0.53, 0.57, 0.57, 0.57, 0.52, 0.54, 0.61, 0.62, 0.59, 0.66, 0.66, 0.52, 
    0.57, 0.54, 0.51, 0.53, 0.52, 0.55, 0.52, 0.54, 0.57, 0.47, 0.54, 0.56, 
    0.61, 0.67, 0.78, 0.74, 0.64, 0.7, 0.59, 0.53, 0.53, 0.53, 0.6, 0.72, 
    0.62, 0.57, 0.53, 0.53, 0.49, 0.52, 0.49, 0.59, 0.6, 0.52, 0.5, 0.54, 
    0.55, 0.56, 0.52, 0.52, 0.53, 0.62, 0.6, 0.55, 0.55, 0.55, 0.61, 0.53, 
    0.53, 0.49, 0.55, 0.63, 0.62, 0.71, 0.66, 0.63, 0.69, 0.71, 0.65, 0.71, 
    0.77, 0.73, 0.75, 0.71, 0.78, 0.76, 0.78, 0.85, 0.76, 0.76, 0.7, 0.62, 
    0.7, 0.65, 0.63, 0.65, 0.74, 0.77, 0.76, 0.84, 0.85, 0.87, 0.84, 0.88, 
    0.9, 0.95, 0.96, 0.96, 0.96, 0.97, 0.96, 0.94, 0.98, 0.93, 0.77, 0.74, 
    0.75, 0.72, 0.73, 0.63, 0.63, 0.8, 0.83, 0.79, 0.72, 0.73, 0.78, 0.91, 
    0.87, 0.86, 0.8, 0.77, 0.78, 0.77, 0.68, 0.69, 0.71, 0.62, 0.61, 0.6, 
    0.52, 0.54, 0.5, 0.5, 0.61, 0.64, 0.5, 0.6, 0.6, 0.65, 0.62, 0.61, 0.64, 
    0.65, 0.64, 0.62, 0.66, 0.65, 0.62, 0.76, 0.59, 0.52, 0.52, 0.49, 0.47, 
    0.46, 0.44, 0.48, 0.52, 0.54, 0.61, 0.59, 0.64, 0.66, 0.62, 0.61, 0.61, 
    0.59, 0.69, 0.6, 0.61, 0.58, 0.72, 0.65, 0.62, 0.58, 0.54, 0.54, 0.43, 
    0.45, 0.49, 0.51, 0.5, 0.56, 0.64, 0.61, 0.62, 0.61, 0.7, 0.67, 0.62, 
    0.56, 0.56, 0.6, 0.59, 0.61, 0.62, 0.67, 0.77, 0.75, 0.7, 0.76, 0.92, 
    0.91, 0.9, 0.9, 0.75, 0.69, 0.65, 0.64, 0.56, 0.63, 0.61, 0.67, 0.71, 
    0.7, 0.71, 0.72, 0.71, 0.68, 0.71, 0.7, 0.66, 0.65, 0.56, 0.59, 0.63, 
    0.57, 0.48, 0.44, 0.45, 0.45, 0.46, 0.48, 0.54, 0.55, 0.57, 0.56, 0.6, 
    0.65, 0.6, 0.6, 0.64, 0.68, 0.6, 0.62, 0.62, 0.64, 0.7, 0.73, 0.58, 0.66, 
    0.61, 0.74, 0.8, 0.87, 0.96, 0.96, 0.99, 1, 0.89, 1, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.89, 0.84, 0.8, 0.83, 0.79, 0.73, 0.68, 0.66, 0.61, 
    0.62, 0.68, 0.71, 0.69, 0.73, 0.71, 0.61, 0.55, 0.6, 0.54, 0.56, 0.44, 
    0.49, 0.48, 0.47, 0.57, 0.61, 0.58, 0.56, 0.63, 0.6, 0.55, 0.54, 0.57, 
    0.5, 0.55, 0.59, 0.61, 0.56, 0.67, 0.65, 0.6, 0.59, 0.61, 0.56, 0.61, 
    0.62, 0.57, 0.66, 0.61, 0.64, 0.63, 0.59, 0.56, 0.53, 0.55, 0.51, 0.57, 
    0.58, 0.58, 0.59, 0.6, 0.68, 0.68, 0.65, 0.66, 0.64, 0.63, 0.61, 0.69, 
    0.6, 0.62, 0.59, 0.59, 0.61, 0.53, 0.56, 0.53, 0.51, 0.49, 0.48, 0.49, 
    0.56, 0.53, 0.53, 0.53, 0.55, 0.59, 0.59, 0.61, 0.58, 0.6, 0.61, 0.62, 
    0.65, 0.61, 0.63, 0.61, 0.6, 0.6, 0.59, 0.55, 0.55, 0.57, 0.58, 0.59, 
    0.59, 0.58, 0.58, 0.62, 0.66, 0.7, 0.7, 0.66, 0.66, 0.62, 0.66, 0.63, 
    0.65, 0.66, 0.68, 0.65, 0.66, 0.66, 0.56, 0.51, 0.51, 0.49, 0.52, 0.5, 
    0.49, 0.52, 0.55, 0.54, 0.58, 0.58, 0.53, 0.57, 0.62, 0.56, 0.55, 0.53, 
    0.64, 0.56, 0.56, 0.63, 0.59, 0.61, 0.59, 0.48, 0.5, 0.53, 0.41, 0.51, 
    0.52, 0.47, 0.56, 0.55, 0.55, 0.61, 0.62, 0.57, 0.6, 0.64, 0.66, 0.64, 
    0.66, 0.64, 0.66, 0.65, 0.63, 0.63, 0.52, 0.58, 0.47, 0.49, 0.48, 0.45, 
    0.51, 0.53, 0.48, 0.56, 0.51, 0.57, 0.62, 0.61, 0.62, 0.65, 0.57, 0.57, 
    0.62, 0.57, 0.61, 0.56, 0.55, 0.57, 0.48, 0.44, 0.45, 0.49, 0.46, 0.47, 
    0.49, 0.49, 0.52, 0.48, 0.52, 0.58, 0.52, 0.57, 0.61, 0.61, 0.64, 0.64, 
    0.59, 0.51, 0.55, 0.55, 0.5, 0.55, 0.5, 0.47, 0.47, 0.4, 0.49, 0.5, 0.5, 
    0.49, 0.54, 0.53, 0.54, 0.58, 0.54, 0.56, 0.63, 0.57, 0.63, 0.65, 0.65, 
    0.62, 0.62, 0.65, 0.62, 0.58, 0.54, 0.52, 0.48, 0.47, 0.46, 0.46, 0.52, 
    0.54, 0.52, 0.56, 0.65, 0.65, 0.66, 0.62, 0.67, 0.69, 0.65, 0.64, 0.64, 
    0.66, 0.66, 0.7, 0.69, 0.75, 0.76, 0.67, 0.78, 0.68, 0.7, 0.66, 0.75, 
    0.74, 0.83, 0.89, 0.85, 0.89, 0.86, 0.82, 0.88, 0.94, 0.94, 0.96, 0.97, 
    0.98, 0.97, 0.96, 0.93, 0.95, 0.94, 0.89, 0.87, 0.85, 0.9, 0.88, 0.88, 
    0.92, 0.97, 0.98, 0.99, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.95, 0.89, 
    0.91, 0.83, 0.64, 0.63, 0.58, 0.58, 0.57, 0.57, 0.6, 0.55, 0.53, 0.53, 
    0.5, 0.52, 0.52, 0.54, 0.62, 0.59, 0.63, 0.7, 0.76, 0.81, 0.81, 0.8, 
    0.83, 0.84, 0.87, 0.84, 0.82, 0.85, 0.86, 0.85, 0.83, 0.85, 0.67, 0.64, 
    0.63, 0.65, 0.65, 0.6, 0.61, 0.6, 0.59, 0.58, 0.59, 0.59, 0.55, 0.59, 
    0.58, 0.59, 0.56, 0.56, 0.56, 0.52, 0.51, 0.52, 0.51, 0.5, 0.48, 0.53, 
    0.5, 0.51, 0.55, 0.57, 0.65, 0.65, 0.66, 0.66, 0.65, 0.65, 0.63, 0.67, 
    0.66, 0.66, 0.63, 0.62, 0.55, 0.57, 0.56, 0.55, 0.56, 0.46, 0.41, 0.45, 
    0.47, 0.56, 0.54, 0.51, 0.57, 0.65, 0.54, 0.59, 0.62, 0.61, 0.65, 0.66, 
    0.67, 0.66, 0.58, 0.55, 0.52, 0.49, 0.5, 0.46, 0.5, 0.4, 0.48, 0.43, 
    0.46, 0.62, 0.6, 0.62, 0.63, 0.66, 0.63, 0.64, 0.66, 0.68, 0.65, 0.59, 
    0.63, 0.59, 0.6, 0.58, 0.53, 0.52, 0.66, 0.65, 0.53, 0.76, 0.74, 0.78, 
    0.84, 0.88, 0.83, 0.88, 0.94, 0.98, 0.95, 0.95, 0.91, 0.95, 0.92, 0.97, 
    0.85, 0.86, 0.79, 0.73, 0.69, 0.68, 0.68, 0.69, 0.68, 0.69, 0.63, 0.6, 
    0.55, 0.61, 0.6, 0.66, 0.64, 0.61, 0.65, 0.69, 0.69, 0.64, 0.68, 0.73, 
    0.7, 0.68, 0.67, 0.62, 0.59, 0.66, 0.63, 0.61, 0.67, 0.6, 0.61, 0.54, 
    0.57, 0.61, 0.65, 0.6, 0.6, 0.64, 0.62, 0.57, 0.63, 0.61, 0.68, 0.66, 
    0.62, 0.65, 0.65, 0.52, 0.62, 0.52, 0.52, 0.54, 0.56, 0.53, 0.59, 0.53, 
    0.59, 0.52, 0.56, 0.63, 0.64, 0.7, 0.66, 0.73, 0.71, 0.71, 0.68, 0.72, 
    0.69, 0.68, 0.64, 0.58, 0.63, 0.63, 0.62, 0.56, 0.61, 0.59, 0.52, 0.55, 
    0.46, 0.51, 0.51, 0.51, 0.56, 0.61, 0.62, 0.6, 0.64, 0.66, 0.69, 0.68, 
    0.62, 0.69, 0.68, 0.65, 0.56, 0.56, 0.46, 0.55, 0.52, 0.54, 0.6, 0.69, 
    0.76, 0.84, 0.85, 0.82, 0.79, 0.9, 0.9, 0.91, 0.85, 0.9, 0.95, 0.93, 
    0.89, 0.82, 0.84, 0.86, 0.67, 0.63, 0.64, 0.59, 0.55, 0.61, 0.57, 0.56, 
    0.55, 0.52, 0.57, 0.56, 0.6, 0.63, 0.62, 0.61, 0.62, 0.64, 0.6, 0.64, 
    0.62, 0.64, 0.65, 0.6, 0.58, 0.55, 0.58, 0.57, 0.49, 0.53, 0.52, 0.54, 
    0.59, 0.6, 0.59, 0.58, 0.65, 0.68, 0.69, 0.73, 0.68, 0.63, 0.68, 0.7, 
    0.66, 0.71, 0.69, 0.61, 0.58, 0.62, 0.61, 0.62, 0.69, 0.65, 0.69, 0.62, 
    0.57, 0.7, 0.69, 0.74, 0.77, 0.74, 0.75, 0.8, 0.77, 0.76, 0.77, 0.76, 
    0.83, 0.71, 0.7, 0.66, 0.65, 0.58, 0.62, 0.56, 0.51, 0.55, 0.56, 0.55, 
    0.57, 0.55, 0.6, 0.62, 0.68, 0.71, 0.74, 0.74, 0.75, 0.71, 0.64, 0.69, 
    0.62, 0.57, 0.51, 0.59, 0.44, 0.5, 0.46, 0.53, 0.52, 0.48, 0.56, 0.54, 
    0.51, 0.48, 0.5, 0.53, 0.55, 0.57, 0.59, 0.61, 0.58, 0.57, 0.62, 0.56, 
    0.57, 0.51, 0.54, 0.47, 0.49, 0.55, 0.56, 0.53, 0.42, 0.46, 0.44, 0.45, 
    0.75, 0.75, 0.53, 0.58, 0.65, 0.74, 0.73, 0.78, 0.78, 0.78, 0.75, 0.72, 
    0.7, 0.67, 0.62, 0.63, 0.68, 0.64, 0.61, 0.63, 0.58, 0.59, 0.55, 0.55, 
    0.56, 0.59, 0.63, 0.68, 0.6, 0.56, 0.67, 0.72, 0.73, 0.73, 0.71, 0.68, 
    0.6, 0.6, 0.5, 0.48, 0.48, 0.49, 0.52, 0.51, 0.49, 0.39, 0.48, 0.45, 
    0.44, 0.5, 0.58, 0.52, 0.6, 0.63, 0.67, 0.67, 0.7, 0.68, 0.68, 0.67, 
    0.69, 0.7, 0.69, 0.66, 0.63, 0.64, 0.67, 0.65, 0.56, 0.56, 0.59, 0.53, 
    0.53, 0.58, 0.6, 0.66, 0.63, 0.74, 0.75, 0.76, 0.77, 0.76, 0.75, 0.74, 
    0.75, 0.66, 0.64, 0.58, 0.52, 0.55, 0.5, 0.55, 0.52, 0.49, 0.53, 0.5, 
    0.58, 0.59, 0.56, 0.58, 0.59, 0.62, 0.64, 0.64, 0.54, 0.56, 0.6, 0.56, 
    0.53, 0.52, 0.59, 0.58, 0.57, 0.54, 0.54, 0.5, 0.57, 0.6, 0.63, 0.62, 
    0.65, 0.64, 0.61, 0.54, 0.6, 0.61, 0.56, 0.62, 0.61, 0.64, 0.58, 0.62, 
    0.69, 0.79, 0.66, 0.53, 0.53, 0.55, 0.62, 0.58, 0.55, 0.59, 0.54, 0.56, 
    0.59, 0.58, 0.53, 0.59, 0.55, 0.64, 0.68, 0.68, 0.7, 0.74, 0.78, 0.77, 
    0.76, 0.71, 0.69, 0.61, 0.51, 0.56, 0.55, 0.62, 0.61, 0.58, 0.58, 0.64, 
    0.65, 0.64, 0.63, 0.64, 0.67, 0.76, 0.77, 0.81, 0.79, 0.76, 0.76, 0.81, 
    0.78, 0.64, 0.65, 0.58, 0.51, 0.48, 0.51, 0.43, 0.57, 0.47, 0.54, 0.6, 
    0.64, 0.64, 0.6, 0.62, 0.6, 0.75, 0.74, 0.71, 0.75, 0.78, 0.78, 0.68, 
    0.77, 0.74, 0.71, 0.64, 0.65, 0.61, 0.66, 0.61, 0.68, 0.59, 0.68, 0.74, 
    0.71, 0.78, 0.78, 0.75, 0.85, 0.97, 0.99, 0.83, 0.85, 0.93, 0.93, 0.93, 
    0.89, 0.91, 0.92, 0.91, 0.88, 0.93, 0.86, 0.93, 0.91, 0.97, 0.87, 0.87, 
    0.93, 0.95, 0.92, 0.91, 0.86, 0.88, 0.82, 0.85, 0.83, 0.8, 0.8, 0.79, 
    0.78, 0.86, 0.86, 0.88, 0.89, 0.87, 0.89, 0.84, 0.77, 0.83, 0.83, 0.8, 
    0.75, 0.72, 0.77, 0.77, 0.75, 0.7, 0.73, 0.76, 0.78, 0.81, 0.75, 0.83, 
    0.84, 0.84, 0.89, 0.89, 0.79, 0.71, 0.56, 0.5, 0.47, 0.47, 0.55, 0.51, 
    0.52, 0.54, 0.58, 0.6, 0.68, 0.73, 0.72, 0.82, 0.78, 0.88, 0.91, 0.92, 
    0.9, 0.85, 0.82, 0.9, 0.77, 0.81, 0.82, 0.7, 0.65, 0.66, 0.75, 0.65, 
    0.63, 0.63, 0.79, 0.78, 0.71, 0.69, 0.74, 0.69, 0.69, 0.67, 0.68, 0.67, 
    0.62, 0.56, 0.59, 0.62, 0.55, 0.58, 0.5, 0.51, 0.51, 0.6, 0.56, 0.51, 
    0.55, 0.55, 0.61, 0.61, 0.62, 0.61, 0.61, 0.61, 0.63, 0.61, 0.62, 0.63, 
    0.61, 0.61, 0.59, 0.59, 0.6, 0.56, 0.56, 0.56, 0.6, 0.57, 0.55, 0.57, 
    0.56, 0.55, 0.52, 0.51, 0.51, 0.52, 0.6, 0.59, 0.6, 0.69, 0.63, 0.71, 
    0.57, 0.59, 0.58, 0.53, 0.52, 0.54, 0.53, 0.5, 0.51, 0.52, 0.47, 0.38, 
    0.43, 0.48, 0.49, 0.49, 0.54, 0.57, 0.6, 0.63, 0.62, 0.63, 0.6, 0.6, 
    0.53, 0.56, 0.55, 0.52, 0.47, 0.52, 0.51, 0.48, 0.5, 0.5, 0.49, 0.52, 
    0.54, 0.55, 0.54, 0.57, 0.57, 0.6, 0.6, 0.58, 0.72, 0.71, 0.67, 0.65, 
    0.66, 0.64, 0.67, 0.62, 0.57, 0.57, 0.56, 0.5, 0.49, 0.47, 0.5, 0.47, 
    0.52, 0.53, 0.53, 0.52, 0.53, 0.54, 0.57, 0.61, 0.64, 0.66, 0.69, 0.62, 
    0.55, 0.55, 0.52, 0.54, 0.56, 0.53, 0.58, 0.52, 0.55, 0.51, 0.49, 0.5, 
    0.54, 0.6, 0.63, 0.64, 0.62, 0.62, 0.63, 0.62, 0.7, 0.83, 0.81, 0.89, 
    0.92, 0.86, 0.83, 0.87, 0.91, 0.86, 0.88, 0.92, 0.94, 0.91, 0.9, 0.99, 
    0.99, 1, 0.99, 0.99, 1, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.84, 0.73, 0.93, 
    0.84, 0.7, 0.64, 0.62, 0.63, 0.57, 0.56, 0.59, 0.53, 0.55, 0.5, 0.54, 
    0.57, 0.63, 0.68, 0.68, 0.68, 0.68, 0.64, 0.65, 0.63, 0.68, 0.64, 0.64, 
    0.57, 0.58, 0.6, 0.54, 0.55, 0.59, 0.52, 0.62, 0.63, 0.59, 0.56, 0.65, 
    0.59, 0.59, 0.6, 0.67, 0.81, 0.79, 0.87, 0.85, 0.81, 0.74, 0.75, 0.84, 
    0.89, 0.82, 0.76, 0.76, 0.8, 0.79, 0.73, 0.8, 0.99, 0.99, 0.99, 0.99, 
    0.92, 0.93, 1, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.92, 0.92, 
    0.71, 0.72, 0.72, 0.64, 0.67, 0.69, 0.7, 0.71, 0.65, 0.67, 0.69, 0.67, 
    0.61, 0.69, 0.72, 0.74, 0.69, 0.83, 0.68, 0.83, 0.72, 0.51, 0.62, 0.62, 
    0.62, 0.57, 0.53, 0.52, 0.56, 0.53, 0.5, 0.51, 0.57, 0.56, 0.58, 0.58, 
    0.54, 0.57, 0.71, 0.67, 0.68, 0.68, 0.65, 0.68, 0.62, 0.65, 0.54, 0.71, 
    0.62, 0.6, 0.53, 0.53, 0.49, 0.47, 0.5, 0.51, 0.5, 0.55, 0.47, 0.51, 
    0.58, 0.63, 0.63, 0.69, 0.75, 0.73, 0.75, 0.84, 0.9, 0.75, 0.75, 0.67, 
    0.6, 0.63, 0.6, 0.6, 0.57, 0.53, 0.65, 0.69, 0.56, 0.5, 0.6, 0.61, 0.63, 
    0.69, 0.68, 0.61, 0.71, 0.74, 0.78, 0.88, 0.86, 0.91, 0.75, 0.7, 0.74, 
    0.71, 0.66, 0.69, 0.69, 0.6, 0.61, 0.61, 0.57, 0.61, 0.64, 0.68, 0.71, 
    0.67, 0.74, 0.72, 0.75, 0.79, 0.79, 0.94, 0.91, 0.92, 0.8, 0.68, 0.81, 
    0.68, 0.59, 0.64, 0.67, 0.63, 0.65, 0.58, 0.54, 0.63, 0.62, 0.64, 0.56, 
    0.56, 0.62, 0.75, 0.85, 0.82, 0.82, 0.84, 0.85, 0.79, 0.78, 0.67, 0.66, 
    0.62, 0.63, 0.67, 0.63, 0.66, 0.68, 0.67, 0.64, 0.81, 0.82, 0.81, 0.61, 
    0.99, 0.99, 1, 1, 1, 1, 1, 0.99, 1, 0.99, 1, 0.93, 0.97, 0.9, 0.95, 0.95, 
    0.91, 0.88, 0.95, 0.88, 0.95, 0.98, 0.96, 0.99, 0.96, 0.93, 0.93, 0.98, 
    0.99, 1, 1, 1, 1, 1, 0.96, 0.88, 1, 0.88, 0.87, 0.84, 0.82, 0.82, 0.86, 
    0.83, 0.89, 0.91, 0.97, 0.99, 0.95, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    1, 1, 1, 1, 1, 1, 0.87, 0.88, 0.85, 0.79, 0.92, 0.93, 0.99, 0.99, 1, 1, 
    0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 1, 1, 0.91, 1, 1, 0.98, 
    0.99, 1, 1, 1, 0.99, 1, 0.99, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 0.99, 1, 1, 
    0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.89, 0.84, 0.88, 0.79, 0.8, 0.76, 0.83, 
    0.79, 0.82, 0.79, 0.8, 0.79, 0.84, 0.81, 0.82, 0.84, 0.85, 0.88, 0.85, 
    0.87, 0.84, 0.85, 0.82, 0.81, 0.78, 0.76, 0.74, 0.7, 0.72, 0.7, 0.68, 
    0.69, 0.72, 0.7, 0.72, 0.7, 0.68, 0.69, 0.68, 0.77, 0.78, 0.77, 0.84, 
    0.8, 0.72, 0.87, 0.84, 0.72, 0.76, 0.8, 0.82, 0.82, 0.82, 0.93, 0.92, 
    0.83, 0.76, 0.74, 0.76, 0.78, 0.89, 0.84, 0.88, 0.82, 0.81, 0.82, 0.87, 
    0.81, 0.81, 0.72, 0.59, 0.74, 0.64, 0.62, 0.7, 0.74, 0.7, 0.67, 0.62, 
    0.65, 0.63, 0.62, 0.63, 0.68, 0.64, 0.7, 0.71, 0.72, 0.74, 0.94, 0.99, 
    0.88, 0.85, 0.9, 0.8, 0.68, 0.78, 0.75, 0.77, 0.69, 0.68, 0.7, 0.69, 
    0.63, 0.64, 0.66, 0.68, 0.7, 0.71, 0.7, 0.79, 0.86, 0.94, 1, 0.9, 0.86, 
    0.78, 0.75, 0.88, 0.81, 0.89, 0.88, 0.75, 0.93, 0.82, 0.66, 0.63, 0.67, 
    0.72, 0.7, 0.67, 0.68, 0.73, 0.73, 0.74, 0.78, 0.89, 0.89, 0.99, 0.89, 
    0.8, 0.77, 0.85, 0.74, 0.67, 0.72, 0.66, 0.68, 0.62, 0.65, 0.64, 0.89, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.95, 0.99, 0.98, 1, 0.93, 
    0.93, 0.91, 0.96, 0.92, 0.93, 0.88, 0.84, 0.87, 0.85, 0.85, 0.85, 0.79, 
    0.85, 0.94, 0.89, 0.93, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 1, 1, 0.99, 1, 0.99, 1, 0.98, 0.99, 1, 1, 0.9, 0.86, 
    0.92, 0.95, 0.99, 0.9, 0.94, 1, 0.94, 0.89, 0.99, 1, 1, 1, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.97, 1, 0.99, 1, 1, 0.99, 1, 1, 0.99, 0.99, 
    0.99, 1, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 1, 0.83, 0.86, 0.91, 0.96, 
    0.93, 0.93, 0.92, 0.87, 0.89, 0.89, 0.9, 0.97, 1, 0.93, 0.96, 0.97, 0.99, 
    0.92, 0.87, 0.85, 0.77, 0.76, 0.74, 0.88, 0.82, 0.8, 0.75, 0.53, 0.52, 
    0.61, 0.61, 0.56, 0.52, 0.57, 0.61, 0.64, 0.87, 0.95, 0.74, 0.7, 0.73, 
    0.73, 0.8, 0.8, 0.81, 0.81, 0.83, 0.77, 0.77, 0.74, 0.78, 0.77, 0.77, 
    0.76, 0.77, 0.74, 0.64, 0.52, 0.62, 0.46, 0.53, 0.56, 0.54, 0.54, 0.48, 
    0.54, 0.57, 0.56, 0.53, 0.52, 0.56, 0.55, 0.55, 0.64, 0.72, 0.75, 0.79, 
    0.77, 0.76, 0.74, 0.77, 0.72, 0.73, 0.71, 0.68, 0.69, 0.69, 0.67, 0.6, 
    0.64, 0.61, 0.58, 0.55, 0.47, 0.49, 0.53, 0.62, 0.72, 0.86, 0.72, 0.62, 
    0.54, 0.52, 0.48, 0.49, 0.51, 0.52, 0.87, 0.77, 0.74, 0.65, 0.67, 0.7, 
    0.63, 0.66, 0.55, 0.51, 0.57, 0.54, 0.56, 0.63, 0.53, 0.5, 0.51, 0.52, 
    0.54, 0.56, 0.55, 0.57, 0.56, 0.56, 0.58, 0.58, 0.64, 0.6, 0.61, 0.58, 
    0.6, 0.6, 0.59, 0.58, 0.55, 0.57, 0.55, 0.57, 0.53, 0.56, 0.56, 0.59, 
    0.58, 0.61, 0.62, 0.65, 0.98, 1, 1, 1, 1, 0.99, 0.99, 1, 1, 0.73, 0.99, 
    0.99, 1, 0.99, 0.99, 0.87, 0.79, 0.81, 0.83, 0.77, 0.73, 0.72, 0.71, 
    0.72, 0.74, 0.75, 0.71, 0.72, 0.72, 0.69, 0.69, 0.7, 0.69, 0.63, 0.64, 
    0.63, 0.61, 0.61, 0.58, 0.56, 0.53, 0.59, 0.6, 0.57, 0.59, 0.68, 0.62, 
    0.74, 0.67, 0.65, 0.58, 0.58, 0.57, 0.56, 0.6, 0.63, 0.59, 0.66, 0.62, 
    0.65, 0.63, 0.6, 0.6, 0.62, 0.56, 0.58, 0.58, 0.62, 0.57, 0.54, 0.57, 
    0.6, 0.6, 0.61, 0.64, 0.64, 0.65, 0.66, 0.63, 0.63, 0.66, 0.66, 0.65, 
    0.62, 0.6, 0.61, 0.63, 0.63, 0.62, 0.6, 0.56, 0.61, 0.62, 0.64, 0.64, 
    0.66, 0.65, 0.65, 0.66, 0.64, 0.66, 0.7, 0.66, 0.64, 0.65, 0.66, 0.66, 
    0.61, 0.59, 0.58, 0.56, 0.57, 0.59, 0.6, 0.64, 0.71, 0.72, 0.74, 0.72, 
    0.75, 0.76, 0.76, 0.82, 0.92, 0.92, 0.95, 0.96, 0.92, 0.88, 0.8, 0.77, 
    0.75, 0.75, 0.73, 0.78, 0.77, 0.76, 0.74, 0.74, 0.77, 0.86, 0.81, 0.82, 
    0.8, 0.81, 0.95, 0.9, 0.92, 0.92, 0.89, 0.9, 0.93, 0.86, 0.83, 0.76, 
    0.75, 0.78, 0.77, 0.76, 0.78, 0.78, 0.78, 0.74, 0.74, 0.73, 0.68, 0.65, 
    0.67, 0.65, 0.7, 0.71, 0.72, 0.73, 0.75, 0.75, 0.7, 0.64, 0.64, 0.63, 
    0.7, 0.68, 0.72, 0.77, 0.79, 0.73, 0.79, 0.79, 0.98, 0.77, 0.67, 0.63, 
    0.67, 0.68, 0.7, 0.8, 0.92, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 0.99, 
    0.99, 0.98, 0.98, 0.92, 0.99, 0.99, 0.87, 0.75, 0.73, 0.83, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0.97, 0.98, 0.99, 0.98, 0.99, 0.87, 0.94, 0.89, 0.91, 
    0.91, 0.94, 0.93, 0.91, 1, 0.82, 0.84, 1, 1, 1, 1, 1, 0.99, 1, 0.99, 
    0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 1, 0.99, 0.7, 1, 0.99, 0.87, 0.95, 
    1, 1, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 0.99, 0.99, 
    0.99, 0.99, 1, 0.99, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.87, 1, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.85, 0.63, 0.59, 0.56, 0.54, 
    0.64, 0.63, 0.63, 0.64, 0.66, 0.65, 0.68, 0.69, 0.63, 0.6, 0.61, 0.61, 
    0.59, 0.63, 0.6, 0.57, 0.6, 0.62, 0.65, 0.66, 0.64, 0.68, 0.79, 0.92, 
    0.99, 1, 0.95, 0.92, 0.96, 0.85, 0.96, 0.95, 0.96, 0.99, 0.99, 0.97, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.89, 0.99, 0.93, 0.99, 0.98, 1, 0.7, 
    0.77, 0.8, 0.8, 0.81, 0.84, 0.82, 0.83, 0.83, 0.83, 0.99, 0.87, 0.86, 
    0.85, 0.92, 0.91, 0.96, 0.88, 0.82, 0.88, 0.8, 0.78, 0.75, 0.76, 0.83, 
    0.8, 0.76, 0.8, 0.74, 0.77, 0.77, 0.75, 0.77, 0.85, 0.91, 0.89, 0.95, 
    0.98, 0.99, 0.99, 0.99, 1, 1, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 1, 1, 
    0.99, 1, 1, 1, 1, 1, 1, 1, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 1, 1, 0.9, 0.91, 0.94, 0.89, 0.91, 0.95, 0.91, 0.94, 0.9, 0.94, 
    0.96, 0.92, 0.92, 0.93, 0.93, 0.88, 0.86, 0.89, 0.74, 0.65, 0.75, 0.69, 
    0.9, 0.73, 0.83, 0.77, 0.77, 0.87, 0.75, 0.75, 0.84, 0.9, 0.94, 0.95, 
    0.93, 0.96, 0.97, 0.97, 0.95, 0.92, 0.89, 0.85, 0.81, 0.82, 0.79, 0.79, 
    0.86, 0.89, 0.93, 0.96, 1, 0.99, 0.8, 0.95, 0.95, 0.94, 0.92, 0.93, 1, 
    0.99, 1, 1, 1, 0.88, 0.98, 0.94, 0.99, 0.98, 1, 0.96, 0.94, 0.87, 0.97, 
    0.94, 1, 0.95, 0.89, 0.99, 1, 1, 1, 0.99, 1, 1, 0.99, 0.99, 0.98, 0.88, 
    0.85, 0.73, 0.67, 0.66, 0.66, 0.67, 0.75, 0.67, 0.68, 0.68, 0.64, 0.73, 
    0.6, 0.66, 0.68, 1, 0.99, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 
    1, 1, 0.99, 1, 1, 1, 1, 0.99, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 0.99, 1, 0.99, 1, 1, 1, 0.99, 1, 0.99, 0.99, 1, 0.99, 1, 1, 
    0.99, 0.99, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 0.96, 0.99, 0.99, 0.94, 0.99, 
    1, 1, 1, 1, 0.99, 1, 0.99, 0.99, 1, 1, 0.99, 1, 1, 0.99, 1, 0.91, 0.87, 
    0.8, 0.9, 0.86, 0.9, 0.84, 0.82, 0.81, 0.87, 0.67, 0.7, 0.64, 0.65, 0.65, 
    0.65, 0.67, 0.69, 0.72, 0.68, 0.72, 0.7, 0.71, 0.73, 0.75, 0.77, 0.73, 
    0.69, 0.67, 0.68, 0.67, 0.62, 0.59, 0.57, 0.57, 0.59, 0.59, 0.57, 0.58, 
    0.59, 0.56, 0.58, 0.54, 0.55, 0.59, 0.63, 0.63, 0.64, 0.65, 0.63, 0.61, 
    0.6, 0.94, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.96, 0.99, 0.99, 0.95, 1, 
    0.98, 1, 1, 0.99, 0.97, 0.9, 0.86, 0.99, 1, 0.99, 0.86, 0.73, 0.74, 0.75, 
    0.68, 0.73, 0.78, 0.72, 0.7, 0.67, 0.68, 0.71, 0.75, 0.69, 0.72, 0.67, 
    0.67, 0.73, 0.95, 0.96, 0.96, 0.99, 0.99, 0.99, 1, 0.97, 1, 0.92, 1, 
    0.85, 0.77, 0.77, 0.68, 0.59, 0.58, 0.57, 0.62, 0.57, 0.52, 0.54, 0.62, 
    0.61, 0.62, 0.6, 0.58, 0.6, 0.9, 1, 0.99, 0.99, 0.99, 0.99, 0.97, 1, 1, 
    0.99, 0.95, 0.98, 0.93, 1, 0.99, 1, 1, 1, 1, 0.99, 1, 1, 1, 1, 0.97, 
    0.99, 0.99, 1, 1, 0.99, 1, 1, 1, 1, 0.99, 0.99, 0.8, 0.99, 1, 1, 0.99, 
    0.99, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 1, 1, 0.94, 0.99, 1, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 1, 0.99, 0.99, 0.97, 
    0.96, 0.99, 0.99, 1, 1, 0.99, 1, 1, 1, 1, 0.99, 0.8, 0.8, 0.73, 0.75, 
    0.69, 0.76, 0.74, 0.77, 0.83, 0.88, 0.98, 0.99, 0.99, 0.99, 0.99, 1, 1, 
    1, 0.9, 0.94, 0.94, 0.99, 0.97, 0.93, 0.88, 0.84, 0.8, 0.85, 1, 0.92, 
    0.86, 0.99, 0.99, 0.94, 0.95, 1, 0.96, 1, 0.99, 0.97, 0.99, 1, 1, 1, 1, 
    0.99, 0.99, 0.99, 1, 0.95, 1, 0.99, 0.94, 0.89, 0.84, 0.85, 0.85, 0.99, 
    0.97, 1, 0.78, 0.79, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 0.99, 
    0.99, 0.99, 0.99, 1, 1, 1, 1, 0.99, 0.99, 1, 1, 1, 1, 1, 0.99, 1, 1, 1, 
    0.99, 0.99, 1, 1, 0.86, 0.99, 0.98, 0.99, 1, 1, 0.99, 0.99, 0.95, 0.99, 
    0.95, 0.95, 0.92, 0.91, 0.94, 0.96, 0.95, 0.99, 0.99, 0.99, 0.97, 0.96, 
    0.97, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.93, 0.84, 0.84, 0.78, 0.79, 
    0.76, 0.78, 0.83, 0.92, 1, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 1, 0.99, 1, 
    1, 0.99, 0.99, 1, 1, 1, 1, 1, 0.99, 0.99, 1, 0.94, 1, 0.98, 0.86, 0.87, 
    1, 1, 0.99, 0.97, 1, 0.96, 1, 0.81, 1, 0.96, 0.93, 1, 1, 0.97, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 1, 1, 0.97, 1, 0.99, 1, 1, 0.99, 
    1, 1, 1, 0.98, 0.91, 0.87, 0.91, 0.81, 0.8, 1, 1, 1, 1, 1, 1, 0.96, 0.99, 
    0.99, 0.99, 1, 0.97, 0.99, 0.93, 0.97, 0.88, 0.94, 0.77, 0.9, 0.83, 1, 
    0.83, 0.79, 0.83, 0.81, 0.89, 0.9, 0.92, 0.91, 0.92, 0.97, 0.95, 0.91, 
    0.85, 0.84, 0.83, 0.81, 0.66, 0.63, 0.65, 0.59, 0.54, 0.53, 0.53, 0.53, 
    0.52, 0.53, 0.53, 0.53, 0.6, 0.48, 0.57, 0.56, 0.71, 0.67, 0.61, 0.66, 
    0.66, 0.6, 0.6, 0.61, 0.59, 0.57, 0.56, 0.61, 0.63, 0.62, 0.63, 0.6, 0.6, 
    0.62, 0.66, 0.66, 0.62, 0.63, 0.65, 0.68, 0.66, 0.68, 0.77, 0.98, 0.99, 
    0.99, 0.9, 0.82, 0.77, 0.74, 0.68, 0.67, 0.66, 0.7, 0.69, 0.69, 0.67, 
    0.68, 0.7, 0.68, 0.69, 0.7, 0.71, 0.72, 0.96, 1, 0.98, 0.99, 0.97, 0.92, 
    0.91, 0.85, 0.8, 0.77, 0.78, 0.76, 0.75, 0.74, 0.79, 0.66, 0.65, 0.66, 
    0.68, 0.69, 0.72, 0.76, 0.81, 0.87, 0.93, 0.95, 0.96, 0.96, 0.96, 0.96, 
    0.96, 0.94, 0.85, 0.75, 0.67, 0.64, 0.6, 0.57, 0.55, 0.53, 0.5, 0.49, 
    0.5, 0.53, 0.62, 0.66, 0.71, 0.75, 0.81, 0.86, 0.87, 0.89, 0.9, 0.87, 
    0.84, 0.81, 0.65, 0.61, 0.78, 0.83, 0.55, 0.75, 0.71, 0.5, 0.51, 0.54, 
    0.57, 0.61, 0.68, 0.74, 0.77, 0.79, 0.83, 0.87, 0.91, 0.91, 0.92, 0.93, 
    0.93, 0.94, 0.87, 0.78, 0.93, 1, 1, 0.99, 0.99, 0.99, 0.98, 0.95, 0.94, 
    1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.98, 0.99, 0.99, 0.99, 
    0.99, 0.99, 1, 1, 0.99, 1, 0.95, 0.94, 0.93, 0.99, 0.91, 0.89, 0.9, 0.74, 
    0.93, 0.94, 0.95, 0.97, 1, 0.97, 0.98, 0.94, 0.91, 0.8, 0.74, 0.7, 0.69, 
    0.72, 0.73, 0.74, 0.86, 0.86, 0.9, 0.94, 0.97, 0.86, 0.86, 0.9, 0.87, 
    0.99, 0.99, 1, 0.78, 0.8, 1, 0.99, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 1, 1, 1, 0.99, 0.99, 0.99, 0.75, 0.78, 0.79, 0.99, 
    0.99, 0.99, 0.99, 0.94, 0.84, 0.76, 0.73, 0.77, 0.79, 0.75, 0.72, 0.7, 
    0.68, 0.67, 0.65, 0.62, 0.59, 0.59, 0.78, 0.8, 0.98, 0.98, 1, 1, 0.99, 1, 
    0.99, 1, 1, 0.98, 0.87, 0.82, 0.79, 1, 1, 1, 0.99, 0.67, 0.93, 0.94, 
    0.87, 0.98, 0.94, 0.99, 1, 0.88, 0.88, 0.87, 0.86, 0.84, 0.83, 0.77, 
    0.63, 0.67, 0.67, 0.66, 0.63, 0.63, 0.56, 0.65, 0.64, 0.58, 0.6, 0.64, 
    0.66, 0.67, 0.66, 0.65, 0.65, 0.66, 0.67, 0.7, 0.71, 0.7, 0.68, 0.77, 
    0.77, 0.97, 0.74, 0.72, 0.7, 0.73, 0.73, 0.73, 0.71, 0.71, 0.69, 0.75, 
    0.75, 0.8, 0.86, 0.92, 1, 0.92, 0.96, 0.97, 0.97, 0.96, 0.96, 0.93, 0.91, 
    0.88, 0.88, 0.93, 0.92, 0.89, 0.82, 0.94, 0.82, 0.82, 0.9, 0.89, 0.87, 
    0.87, 0.93, 0.94, 0.94, 0.92, 0.92, 0.9, 1, 0.95, 0.99, 1, 0.99, 0.96, 
    0.9, 0.8, 0.75, 0.74, 0.68, 0.68, 0.67, 0.68, 0.67, 1, 0.69, 1, 1, 0.8, 
    1, 0.77, 0.82, 0.9, 0.89, 0.89, 0.91, 0.98, 0.89, 0.83, 0.79, 0.74, 0.66, 
    0.64, 0.68, 0.64, 0.65, 0.72, 0.65, 0.66, 0.67, 0.68, 0.69, 0.71, 0.77, 
    0.81, 0.89, 0.94, 0.96, 0.99, 0.9, 0.89, 0.88, 0.88, 0.83, 0.78, 0.68, 
    0.63, 0.65, 0.7, 0.71, 0.67, 0.69, 0.74, 0.69, 0.68, 0.68, 0.76, 0.85, 
    0.82, 0.87, 0.93, 0.95, 0.87, 0.93, 0.91, 0.88, 0.78, 0.77, 0.73, 0.65, 
    0.66, 0.62, 0.59, 0.58, 0.54, 0.55, 0.56, 0.57, 0.58, 0.6, 0.61, 0.62, 
    0.64, 0.67, 0.68, 0.71, 0.63, 0.67, 0.66, 0.65, 0.76, 0.64, 0.62, 0.59, 
    0.57, 0.56, 0.59, 0.58, 0.57, 0.55, 0.6, 0.69, 0.71, 0.72, 0.76, 0.8, 
    0.84, 0.88, 0.91, 0.91, 0.91, 1, 1, 0.89, 0.83, 0.71, 0.64, 0.67, 0.6, 
    0.59, 0.6, 0.6, 0.59, 0.62, 0.62, 0.64, 0.66, 0.69, 0.72, 0.8, 0.84, 
    0.87, 0.9, 0.91, 0.95, 0.99, 1, 0.84, 0.95, 0.87, 0.79, 0.71, 0.64, 0.58, 
    0.53, 0.51, 0.5, 0.51, 0.5, 0.49, 0.52, 0.51, 0.58, 0.64, 0.72, 0.78, 
    0.81, 0.96, 0.99, 0.99, 1, 0.89, 0.88, 0.86, 0.91, 0.85, 0.74, 0.79, 
    0.71, 0.73, 0.65, 0.7, 0.71, 0.65, 0.68, 0.72, 0.79, 0.83, 0.83, 0.81, 
    0.81, 0.83, 0.85, 0.87, 0.9, 0.92, 0.93, 0.95, 0.93, 0.83, 0.73, 0.64, 
    0.56, 0.57, 0.54, 0.56, 0.73, 0.75, 0.77, 0.78, 0.81, 0.82, 0.95, 0.99, 
    0.99, 0.99, 0.9, 0.86, 0.85, 0.82, 0.79, 0.76, 0.72, 0.69, 0.68, 0.67, 
    0.65, 0.64, 0.64, 0.64, 0.66, 0.7, 0.73, 0.78, 0.82, 0.86, 0.93, 0.97, 
    0.99, 0.98, 0.96, 1, 0.93, 0.96, 0.96, 0.87, 0.76, 0.67, 0.59, 0.53, 
    0.54, 0.54, 0.56, 0.56, 0.6, 0.65, 0.68, 0.64, 0.69, 0.76, 0.83, 0.92, 
    0.99, 1, 0.99, 0.99, 1, 0.84, 0.96, 1, 0.76, 0.71, 0.68, 0.8, 0.76, 0.75, 
    0.8, 0.59, 0.66, 0.65, 0.68, 0.73, 0.84, 0.99, 0.99, 1, 1, 0.99, 1, 0.81, 
    0.8, 0.99, 0.99, 0.98, 0.97, 0.95, 0.91, 0.8, 0.78, 0.76, 0.85, 0.79, 
    0.74, 0.87, 0.78, 0.7, 0.84, 0.86, 0.85, 0.85, 0.93, 0.94, 0.96, 0.99, 
    0.99, 1, 0.99, 0.99, 0.83, 0.84, 0.9, 0.9, 0.9, 0.91, 0.94, 0.9, 0.86, 
    0.87, 0.86, 0.86, 0.94, 0.99, 0.92, 0.98, 0.89, 0.92, 1, 0.98, 1, 1, 1, 
    0.99, 1, 1, 0.99, 1, 1, 1, 0.99, 1, 1, 0.91, 0.83, 0.7, 0.7, 0.81, 0.93, 
    0.87, 0.93, 0.75, 0.8, 0.85, 0.89, 0.86, 0.82, 0.78, 0.79, 0.79, 0.83, 
    0.78, 0.73, 0.69, 0.69, 0.77, 0.7, 0.65, 0.69, 0.64, 0.66, 0.69, 0.72, 
    0.64, 0.61, 0.64, 0.63, 0.68, 0.67, 0.71, 0.68, 0.65, 0.64, 0.58, 0.64, 
    0.63, 0.64, 0.67, 0.99, 0.96, 0.8, 0.82, 0.84, 0.69, 0.67, 0.64, 0.7, 
    0.63, 0.62, 0.66, 0.67, 0.64, 0.65, 0.67, 0.8, 0.69, 0.67, 0.6, 0.57, 
    0.56, 0.58, 0.61, 0.59, 0.61, 0.6, 0.64, 0.63, 0.72, 0.7, 0.68, 0.66, 
    0.7, 0.68, 0.73, 0.73, 0.7, 0.73, 0.8, 0.87, 0.83, 0.67, 0.71, 0.69, 
    0.71, 0.69, 0.68, 0.65, 0.68, 0.66, 0.65, 0.67, 0.72, 0.73, 0.71, 0.76, 
    0.8, 0.99, 1, 0.99, 0.9, 0.81, 0.87, 0.77, 0.79, 0.88, 0.77, 0.67, 0.63, 
    0.64, 0.66, 0.67, 0.66, 0.67, 0.67, 0.64, 0.67, 0.67, 0.67, 0.67, 0.71, 
    0.69, 0.7, 0.7, 0.71, 0.71, 0.67, 0.66, 0.78, 0.83, 0.69, 0.65, 0.68, 
    0.67, 0.63, 0.64, 0.62, 0.64, 0.69, 0.9, 0.73, 0.74, 0.74, 0.75, 0.75, 
    0.76, 0.76, 0.75, 0.87, 0.67, 0.68, 0.67, 0.68, 0.67, 0.66, 0.66, 0.66, 
    0.66, 0.66, 0.65, 0.66, 0.66, 0.65, 0.65, 0.72, 0.68, 0.68, 0.74, 0.74, 
    0.74, 0.77, 0.78, 0.78, 0.82, 0.87, 1, 0.92, 0.91, 0.92, 0.99, 0.99, 
    0.99, 0.99, 0.95, 0.83, 0.88, 0.92, 0.94, 0.9, 0.92, 1, 1, 0.99, 0.99, 
    0.99, 1, 1, 0.99, 0.99, 0.96, 0.95, 0.91, 0.89, 1, 0.99, 0.99, 1, 1, 
    0.99, 0.99, 1, 1, 0.95, 0.97, 0.97, 0.96, 0.84, 0.73, 0.69, 0.64, 0.66, 
    0.65, 0.68, 0.68, 0.71, 0.69, 0.67, 0.66, 0.63, 0.62, 0.62, 0.58, 0.58, 
    0.57, 0.6, 0.56, 0.68, 0.67, 0.71, 0.79, 0.79, 0.84, 0.9, 0.93, 0.92, 
    0.88, 0.91, 0.87, 0.91, 0.9, 0.84, 0.82, 0.79, 0.92, 1, 1, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.84, 1, 1, 1, 0.79, 0.91, 0.73, 
    0.74, 0.7, 0.67, 0.66, 0.65, 0.68, 0.67, 0.66, 0.68, 0.7, 0.71, 0.73, 
    0.79, 0.86, 0.8, 0.84, 0.85, 0.87, 0.88, 0.89, 0.91, 1, 1, 0.99, 0.99, 
    0.99, 1, 0.99, 0.8, 0.68, 0.68, 0.68, 0.68, 0.68, 0.67, 0.72, 0.78, 0.68, 
    0.69, 0.92, 0.92, 0.92, 0.93, 0.92, 0.89, 0.79, 0.81, 0.84, 0.9, 0.86, 
    0.81, 0.68, 0.71, 0.59, 0.58, 0.59, 0.6, 0.61, 0.66, 0.64, 0.71, 0.77, 
    0.77, 0.79, 0.77, 0.72, 0.66, 0.65, 0.68, 0.71, 0.7, 0.73, 0.63, 0.63, 
    0.65, 0.67, 0.63, 0.63, 0.66, 0.72, 0.83, 0.99, 0.99, 0.99, 0.85, 0.88, 
    0.94, 0.99, 1, 1, 0.99, 1, 0.99, 1, 0.99, 0.89, 0.92, 0.89, 0.99, 1, 
    0.99, 1, 1, 1, 0.99, 1, 1, 0.92, 0.89, 0.95, 0.99, 1, 0.99, 0.86, 0.84, 
    0.73, 0.7, 0.74, 0.73, 0.71, 0.73, 0.69, 0.69, 0.62, 0.69, 0.68, 0.66, 
    0.63, 0.68, 0.64, 0.67, 0.65, 0.64, 0.64, 0.65, 0.67, 0.68, 0.69, 0.7, 
    0.71, 0.73, 0.68, 0.7, 0.73, 0.71, 0.69, 0.69, 0.67, 0.62, 0.62, 0.67, 
    0.61, 0.69, 0.65, 0.77, 0.8, 0.81, 0.68, 0.68, 0.79, 0.8, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 1, 1, 0.97, 0.98, 0.99, 0.99, 1, 1, 1, 0.99, 
    0.99, 1, 1, 0.91, 0.96, 0.99, 0.79, 0.99, 1, 0.96, 0.83, 0.78, 0.9, 0.84, 
    0.81, 0.79, 0.76, 0.74, 0.77, 0.71, 0.59, 0.64, 0.76, 0.64, 0.62, 0.7, 
    0.71, 0.71, 0.7, 0.68, 0.67, 0.6, 0.66, 0.7, 0.71, 0.75, 0.81, 0.79, 
    0.72, 0.68, 0.71, 0.68, 0.6, 0.65, 0.56, 0.64, 0.61, 0.63, 0.66, 0.67, 
    0.67, 0.66, 0.66, 0.67, 0.89, 0.92, 0.94, 0.94, 0.79, 0.79, 0.64, 0.7, 
    0.7, 0.67, 0.67, 0.67, 0.64, 0.61, 0.6, 0.6, 0.56, 0.6, 0.56, 0.59, 0.61, 
    0.69, 0.69, 0.7, 0.67, 0.69, 0.77, 0.85, 0.86, 0.87, 0.89, 0.72, 0.73, 1, 
    1, 0.99, 0.73, 0.57, 0.56, 0.56, 0.59, 0.59, 0.58, 0.61, 0.6, 0.58, 0.59, 
    0.56, 0.53, 0.55, 0.54, 0.57, 0.58, 0.6, 0.64, 0.69, 0.66, 0.67, 0.66, 
    0.67, 0.79, 0.79, 0.77, 0.75, 0.74, 0.7, 0.69, 0.68, 0.74, 0.78, 0.79, 
    0.84, 0.87, 0.89, 0.9, 0.92, 0.92, 0.91, 0.88, 0.89, 0.95, 0.9, 0.92, 
    0.92, 0.82, 0.8, 0.79, 0.76, 0.76, 0.77, 0.76, 0.75, 0.73, 0.75, 0.83, 
    0.92, 0.83, 0.89, 0.83, 0.82, 0.99, 1, 1, 0.99, 0.99, 0.93, 0.88, 0.83, 
    0.81, 0.78, 0.77, 0.78, 0.82, 0.81, 0.89, 0.85, 0.85, 0.84, 0.78, 0.75, 
    0.76, 0.77, 0.77, 0.75, 0.74, 0.74, 0.89, 0.73, 0.73, 0.72, 0.75, 0.72, 
    0.71, 0.71, 0.73, 0.75, 0.84, 0.99, 0.86, 0.99, 0.99, 1, 0.91, 0.89, 
    0.89, 0.9, 0.9, 0.91, 0.93, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.97, 0.92, 0.71, 0.69, 0.7, 0.69, 0.68, 0.66, 0.63, 0.57, 0.58, 
    0.64, 0.68, 0.65, 0.66, 0.75, 0.7, 0.72, 0.76, 0.72, 0.66, 0.64, 0.65, 
    0.64, 0.63, 0.65, 0.66, 0.65, 0.62, 0.6, 0.6, 0.61, 0.64, 0.68, 0.72, 
    0.76, 0.75, 0.72, 0.7, 0.69, 0.68, 0.66, 0.6, 0.69, 0.66, 0.69, 0.64, 
    0.6, 0.59, 0.6, 0.62, 0.65, 0.67, 0.8, 0.72, 0.74, 0.75, 0.77, 0.85, 
    0.89, 0.92, 0.94, 0.94, 0.93, 0.99, 0.96, 0.99, 0.99, 0.87, 0.95, 0.99, 
    0.93, 0.77, 0.77, 0.7, 0.63, 0.64, 0.59, 0.55, 0.56, 0.6, 0.68, 0.71, 
    0.8, 0.75, 0.77, 0.81, 0.79, 0.84, 0.93, 0.99, 0.99, 0.96, 0.93, 0.9, 
    0.9, 0.84, 0.8, 0.86, 0.92, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.94, 0.8, 0.71, 0.74, 0.71, 0.68, 0.65, 0.61, 0.58, 0.58, 0.56, 0.63, 
    0.62, 0.61, 0.81, 0.79, 0.75, 0.64, 0.68, 0.65, 0.62, 0.58, 0.52, 0.54, 
    0.57, 0.56, 0.56, 0.57, 0.85, 0.85, 0.84, 0.84, 0.81, 0.7, 0.72, 0.72, 
    0.66, 0.7, 0.74, 0.69, 0.69, 0.63, 0.59, 0.57, 0.62, 0.65, 0.74, 0.81, 
    0.89, 0.96, 0.99, 0.97, 0.93, 0.9, 1, 0.99, 0.99, 1, 1, 0.99, 1, 0.99, 
    0.99, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 1, 1, 0.99, 0.98, 
    0.97, 0.94, 1, 1, 0.99, 0.99, 1, 0.99, 0.89, 0.92, 1, 0.89, 1, 1, 0.79, 
    0.78, 0.82, 0.85, 0.88, 0.89, 0.88, 0.83, 0.79, 0.78, 0.76, 0.73, 0.7, 
    0.69, 0.74, 0.83, 0.91, 0.78, 0.84, 0.81, 0.8, 0.76, 0.92, 1, 0.99, 0.99, 
    0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.98, 1, 0.9, 0.89, 0.87, 0.88, 0.87, 
    0.91, 0.91, 0.91, 0.88, 0.83, 0.97, 0.99, 1, 1, 0.99, 0.79, 0.99, 0.89, 
    0.99, 0.99, 1, 0.99, 0.95, 0.89, 0.83, 0.85, 0.89, 0.88, 0.88, 0.88, 
    0.89, 0.81, 0.8, 0.79, 0.79, 0.82, 0.84, 0.79, 0.77, 0.76, 0.78, 0.79, 
    0.75, 0.71, 0.7, 0.7, 0.72, 0.76, 0.73, 0.73, 0.73, 0.72, 0.71, 0.71, 
    0.7, 0.67, 0.67, 0.72, 0.77, 0.75, 0.78, 0.85, 0.73, 0.68, 0.64, 0.71, 
    0.74, 0.79, 0.8, 0.81, 0.83, 0.84, 0.84, 0.85, 0.81, 0.86, 0.88, 0.87, 
    0.88, 0.81, 0.83, 0.82, 0.84, 0.84, 0.85, 0.87, 0.87, 0.89, 0.91, 0.94, 
    0.97, 0.99, 0.9, 0.87, 0.92, 0.95, 0.89, 0.93, 0.95, 0.81, 0.98, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.92, 0.92, 0.9, 
    0.89, 0.99, 1, 1, 1, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 
    0.99, 0.99, 1, 0.99, 0.99, 0.97, 0.96, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.96, 0.93, 0.87, 0.9, 0.92, 
    0.95, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.97, 0.97, 0.98, 0.99, 
    0.99, 0.99, 0.97, 0.94, 0.87, 0.82, 0.8, 0.8, 0.79, 0.71, 0.75, 0.8, 
    0.85, 0.88, 0.85, 0.88, 0.88, 0.88, 0.88, 0.87, 0.89, 0.81, 0.83, 0.86, 
    0.8, 0.8, 0.83, 0.82, 0.8, 0.79, 0.8, 0.76, 0.73, 0.79, 0.75, 0.75, 0.73, 
    0.72, 0.73, 0.8, 0.77, 0.78, 0.74, 0.76, 0.77, 0.77, 0.79, 0.81, 0.81, 
    0.8, 0.8, 0.82, 0.82, 0.74, 0.65, 0.62, 0.61, 0.59, 0.56, 0.52, 0.54, 
    0.56, 0.59, 0.61, 0.64, 0.63, 0.68, 0.71, 0.7, 0.71, 0.68, 0.7, 0.72, 
    0.72, 0.72, 0.73, 0.75, 0.74, 0.71, 0.72, 0.73, 0.73, 0.84, 0.83, 0.64, 
    0.63, 0.66, 0.63, 0.62, 0.63, 0.64, 0.68, 0.76, 0.85, 0.85, 0.83, 0.96, 
    0.92, 0.71, 0.7, 0.71, 0.65, 0.64, 0.65, 0.7, 0.68, 0.69, 0.71, 0.64, 
    0.63, 0.62, 0.62, 0.65, 0.62, 0.63, 0.64, 0.65, 0.68, 0.67, 0.71, 0.75, 
    0.73, 0.73, 0.72, 0.71, 0.77, 0.71, 0.7, 0.68, 0.67, 0.66, 0.68, 0.66, 
    0.65, 0.63, 0.64, 0.64, 0.85, 0.63, 0.63, 0.62, 0.63, 0.63, 0.66, 0.69, 
    0.69, 0.69, 0.69, 0.9, 0.91, 0.87, 0.83, 0.77, 0.76, 0.77, 0.72, 0.72, 
    0.71, 0.68, 0.69, 0.7, 0.72, 0.86, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.98, 0.96, 0.72, 0.79, 0.8, 0.81, 0.85, 0.82, 0.79, 0.77, 0.89, 
    0.83, 0.83, 0.79, 0.78, 0.78, 0.78, 0.78, 0.87, 0.82, 0.83, 0.8, 0.8, 
    0.86, 0.83, 0.84, 0.87, 0.9, 0.84, 0.86, 0.94, 0.88, 0.8, 0.81, 0.77, 
    0.65, 0.64, 0.73, 0.74, 0.62, 0.54, 0.61, 0.6, 0.59, 0.57, 0.61, 0.68, 
    0.69, 0.94, 0.65, 0.65, 0.66, 0.91, 0.89, 0.7, 0.73, 0.78, 0.79, 0.77, 
    0.84, 0.83, 0.81, 0.81, 0.85, 0.84, 0.88, 0.88, 0.71, 0.69, 0.71, 0.74, 
    0.76, 0.76, 0.73, 0.71, 0.75, 0.75, 0.88, 0.88, 0.88, 0.88, 0.9, 0.9, 
    0.92, 0.78, 0.79, 0.8, 0.86, 0.76, 0.76, 0.87, 0.73, 0.85, 0.82, 0.87, 
    0.91, 0.97, 0.94, 0.88, 0.84, 0.92, 0.9, 0.76, 0.8, 0.79, 0.94, 0.94, 
    0.79, 0.78, 0.74, 0.75, 0.79, 0.76, 0.79, 0.72, 0.76, 0.87, 0.86, 0.84, 
    0.83, 0.92, 0.81, 0.8, 0.79, 0.82, 0.78, 0.76, 0.74, 0.72, 0.7, 0.75, 
    0.76, 0.76, 0.73, 0.73, 0.73, 0.78, 0.7, 0.71, 0.76, 0.81, 0.82, 0.74, 
    0.7, 0.74, 0.77, 0.78, 0.93, 0.91, 0.87, 0.83, 0.78, 0.78, 0.72, 0.77, 
    0.74, 0.76, 0.71, 0.71, 0.68, 0.67, 0.66, 0.66, 0.63, 0.67, 0.65, 0.64, 
    0.65, 0.64, 0.66, 0.68, 0.83, 0.73, 0.74, 0.71, 0.63, 0.63, 0.6, 0.64, 
    0.62, 0.61, 0.6, 0.78, 0.6, 0.6, 0.61, 0.6, 0.6, 0.58, 0.59, 0.61, 0.6, 
    0.6, 0.77, 0.76, 0.73, 0.59, 0.59, 0.58, 0.59, 0.59, 0.61, 0.62, 0.6, 
    0.63, 0.63, 0.68, 0.65, 0.64, 0.66, 0.69, 0.71, 0.67, 0.68, 0.7, 0.68, 
    0.68, 0.66, 0.67, 0.68, 0.69, 0.69, 0.71, 0.71, 0.73, 0.73, 0.71, 0.67, 
    0.66, 0.67, 0.59, 0.63, 0.67, 0.64, 0.65, 0.64, 0.63, 0.61, 0.63, 0.66, 
    0.61, 0.54, 0.58, 0.64, 0.63, 0.58, 0.63, 0.58, 0.6, 0.59, 0.63, 0.61, 
    0.6, 0.6, 0.62, 0.61, 0.68, 0.71, 0.69, 0.69, 0.67, 0.69, 0.72, 0.73, 
    0.71, 0.71, 0.76, 0.75, 0.73, 0.75, 0.72, 0.74, 0.74, 0.75, 0.74, 0.65, 
    0.66, 0.7, 0.73, 0.78, 0.79, 0.78, 0.84, 0.94, 0.99, 0.99, 0.99, 1, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 
    0.94, 0.86, 0.9, 0.92, 0.91, 0.87, 0.87, 0.84, 0.83, 0.89, 0.93, 0.96, 
    0.99, 0.95, 0.93, 0.89, 0.89, 0.88, 0.91, 0.87, 0.88, 0.87, 0.77, 0.79, 
    0.73, 0.72, 0.69, 0.72, 0.67, 0.66, 0.61, 0.62, 0.63, 0.59, 0.59, 0.59, 
    0.55, 0.54, 0.53, 0.52, 0.54, 0.57, 0.56, 0.56, 0.62, 0.58, 0.61, 0.61, 
    0.6, 0.61, 0.66, 0.67, 0.67, 0.66, 0.67, 0.65, 0.64, 0.67, 0.66, 0.67, 
    0.65, 0.66, 0.66, 0.5, 0.62, 0.48, 0.62, 0.62, 0.64, 0.62, 0.6, 0.6, 
    0.63, 0.62, 0.63, 0.66, 0.64, 0.63, 0.64, 0.64, 0.62, 0.63, 0.69, 0.71, 
    0.76, 0.83, 0.91, 0.96, 0.98, 0.93, 0.96, 0.98, 0.99, 0.98, 0.95, 0.86, 
    0.89, 0.85, 0.86, 0.86, 0.85, 0.83, 0.82, 0.77, 0.73, 0.74, 0.68, 0.65, 
    0.65, 0.66, 0.69, 0.64, 0.68, 0.59, 0.6, 0.58, 0.61, 0.61, 0.66, 0.65, 
    0.64, 0.64, 0.66, 0.67, 0.69, 0.69, 0.73, 0.75, 0.77, 0.74, 0.75, 0.74, 
    0.73, 0.74, 0.73, 0.73, 0.73, 0.74, 0.71, 0.69, 0.62, 0.81, 1, 0.99, 
    0.99, 0.99, 0.9, 0.79, 0.94, 0.89, 0.75, 0.89, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.85, 0.75, 0.93, 0.86, 0.75, 0.78, 0.79, 0.73, 0.77, 0.78, 0.75, 
    0.8, 0.79, 0.84, 0.76, 0.73, 0.63, 0.63, 0.65, 0.67, 0.67, 0.65, 0.63, 
    0.66, 0.64, 0.63, 0.66, 0.64, 0.6, 0.61, 0.61, 0.63, 0.63, 0.65, 0.65, 
    0.63, 0.61, 0.59, 0.58, 0.6, 0.57, 0.56, 0.55, 0.58, 0.58, 0.58, 0.59, 
    0.58, 0.62, 0.63, 0.58, 0.63, 0.58, 0.57, 0.6, 0.55, 0.56, 0.6, 0.57, 
    0.57, 0.57, 0.58, 0.55, 0.57, 0.58, 0.59, 0.62, 0.58, 0.6, 0.58, 0.59, 
    0.58, 0.55, 0.55, 0.58, 0.55, 0.55, 0.59, 0.6, 0.59, 0.61, 0.64, 0.66, 
    0.64, 0.62, 0.66, 0.61, 0.57, 0.58, 0.6, 0.64, 0.61, 0.64, 0.68, 0.7, 
    0.71, 0.73, 0.74, 0.73, 0.71, 0.69, 0.69, 0.68, 0.7, 0.65, 0.65, 0.67, 
    0.68, 0.66, 0.7, 0.63, 0.63, 0.64, 0.63, 0.61, 0.62, 0.58, 0.59, 0.6, 
    0.61, 0.6, 0.63, 0.62, 0.64, 0.67, 0.67, 0.66, 0.67, 0.7, 0.7, 0.71, 
    0.71, 0.68, 0.7, 0.71, 0.69, 0.7, 0.71, 0.7, 0.71, 0.71, 0.73, 0.72, 0.7, 
    0.69, 0.73, 0.73, 0.73, 0.72, 0.72, 0.72, 0.72, 0.72, 0.74, 0.73, 0.73, 
    0.75, 0.76, 0.76, 0.78, 0.83, 0.91, 0.88, 0.88, 0.75, 0.78, 0.8, 0.78, 
    0.78, 0.75, 0.76, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.88, 0.99, 1, 1, 0.99, 0.92, 0.86, 0.89, 0.82, 0.81, 0.76, 0.7, 0.67, 
    0.65, 0.65, 0.63, 0.61, 0.6, 0.62, 0.62, 0.63, 0.62, 0.62, 0.6, 0.57, 
    0.59, 0.65, 0.66, 0.68, 0.63, 0.61, 0.63, 0.64, 0.66, 0.65, 0.65, 0.66, 
    0.67, 0.67, 0.65, 0.63, 0.6, 0.65, 0.6, 0.59, 0.58, 0.57, 0.67, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.82, 
    0.76, 0.77, 0.77, 0.81, 0.83, 0.83, 0.82, 0.8, 0.71, 0.71, 0.72, 0.75, 
    0.73, 0.76, 0.78, 0.8, 0.83, 0.77, 0.81, 0.84, 0.87, 0.83, 0.84, 0.84, 
    0.85, 0.87, 0.8, 0.72, 0.69, 0.71, 0.71, 0.72, 0.78, 0.82, 0.87, 0.99, 
    0.82, 0.79, 0.76, 0.67, 0.69, 0.69, 0.64, 0.61, 0.6, 0.64, 0.63, 0.66, 
    0.69, 0.72, 0.73, 0.71, 0.69, 0.7, 0.69, 0.67, 0.67, 0.68, 0.64, 0.65, 
    0.67, 0.63, 0.63, 0.61, 0.57, 0.59, 0.5, 0.48, 0.48, 0.51, 0.74, 0.89, 
    0.93, 0.78, 0.94, 0.99, 0.9, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.98, 0.93, 0.95, 0.93, 0.98, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.92, 0.94, 1, 1, 0.99, 0.99, 0.99, 1, 0.99, 
    0.99, 1, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 1, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 0.96, 0.98, 0.93, 0.99, 
    0.97, 0.99, 0.83, 1, 0.91, 0.93, 1, 0.94, 0.86, 0.75, 0.67, 0.59, 0.63, 
    0.65, 0.7, 0.69, 0.64, 0.67, 0.71, 0.75, 0.76, 0.76, 0.78, 0.76, 0.76, 
    0.75, 0.77, 0.79, 0.79, 0.81, 0.83, 0.9, 1, 1, 0.99, 0.99, 1, 1, 0.99, 
    0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 
    1, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 
    0.88, 0.8, 0.77, 0.75, 0.82, 0.82, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 
    0.99, 0.99, 0.99, 1, 1, 0.99, 0.99, 1, 1, 1, 0.99, 0.99, 0.94, 1, 1, 
    0.99, 0.99, 0.99, 1, 0.99, 0.95, 1, 0.99, 0.84, 0.96, 0.89, 0.83, 0.78, 
    0.73, 0.83, 0.86, 0.88, 0.87, 0.92, 0.94, 0.99, 0.99, 1, 0.99, 0.99, 
    0.99, 0.92, 0.85, 0.97, 0.92, 0.78, 0.72, 0.73, 0.71, 0.64, 0.6, 0.6, 
    0.62, 0.62, 0.61, 0.61, 0.61, 0.6, 0.58, 0.59, 0.63, 0.68, 0.71, 0.68, 
    0.69, 0.69, 0.69, 0.72, 0.72, 0.72, 0.73, 0.75, 0.78, 0.82, 0.82, 0.84, 
    0.81, 0.82, 0.83, 0.95, 0.93, 0.87, 0.92, 0.91, 0.96, 0.94, 0.92, 0.91, 
    0.96, 0.86, 0.97, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.78, 0.75, 0.82, 0.74, 0.74, 0.74, 0.71, 0.72, 0.74, 0.75, 0.72, 
    0.73, 0.72, 0.71, 0.7, 0.73, 0.7, 0.71, 0.69, 0.74, 0.71, 0.73, 0.75, 
    0.73, 0.68, 0.67, 0.69, 0.67, 0.67, 0.66, 0.66, 0.67, 0.64, 0.64, 0.62, 
    0.63, 0.6, 0.6, 0.6, 0.64, 0.64, 0.66, 0.66, 0.64, 0.59, 0.62, 0.58, 
    0.58, 0.54, 0.57, 0.56, 0.53, 0.54, 0.55, 0.53, 0.61, 0.57, 0.61, 0.57, 
    0.56, 0.52, 0.53, 0.56, 0.56, 0.51, 0.52, 0.53, 0.51, 0.51, 0.6, 0.55, 
    0.5, 0.51, 0.57, 0.58, 0.58, 0.59, 0.63, 0.61, 0.64, 0.61, 0.64, 0.61, 
    0.65, 0.62, 0.6, 0.61, 0.57, 0.6, 0.6, 0.6, 0.6, 0.59, 0.59, 0.58, 0.6, 
    0.58, 0.59, 0.6, 0.63, 0.6, 0.56, 0.58, 0.6, 0.58, 0.61, 0.65, 0.63, 
    0.63, 0.62, 0.6, 0.59, 0.63, 0.61, 0.63, 0.62, 0.62, 0.67, 0.6, 0.54, 
    0.5, 0.55, 0.55, 0.52, 0.59, 0.55, 0.6, 0.56, 0.58, 0.57, 0.55, 0.61, 
    0.63, 0.61, 0.56, 0.58, 0.57, 0.57, 0.58, 0.59, 0.61, 0.6, 0.62, 0.7, 
    0.74, 0.58, 0.57, 0.55, 0.55, 0.54, 0.53, 0.52, 0.53, 0.53, 0.5, 0.53, 
    0.52, 0.52, 0.51, 0.51, 0.53, 0.55, 0.52, 0.52, 0.52, 0.51, 0.51, 0.53, 
    0.52, 0.54, 0.56, 0.57, 0.57, 0.57, 0.57, 0.58, 0.59, 0.56, 0.53, 0.52, 
    0.5, 0.51, 0.5, 0.54, 0.55, 0.55, 0.54, 0.55, 0.55, 0.52, 0.54, 0.53, 
    0.56, 0.55, 0.59, 0.63, 0.63, 0.66, 0.7, 0.72, 0.7, 0.73, 0.73, 0.75, 
    0.76, 0.78, 0.82, 0.84, 0.86, 0.94, 0.97, 0.95, 0.89, 0.85, 0.81, 0.75, 
    0.69, 0.79, 0.72, 0.72, 0.69, 0.72, 0.72, 0.74, 0.67, 0.68, 0.65, 0.65, 
    0.58, 0.6, 0.57, 0.54, 0.53, 0.54, 0.53, 0.54, 0.56, 0.66, 0.52, 0.53, 
    0.54, 0.56, 0.58, 0.57, 0.58, 0.6, 0.62, 0.64, 0.68, 0.64, 0.57, 0.57, 
    0.55, 0.59, 0.59, 0.62, 0.62, 0.67, 0.67, 0.7, 0.68, 0.71, 0.74, 0.84, 
    0.74, 0.76, 0.77, 0.79, 0.89, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.77, 
    0.74, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.81, 0.77, 0.68, 0.84, 0.71, 
    0.91, 0.9, 0.85, 0.82, 0.7, 0.74, 0.72, 0.7, 0.67, 0.74, 0.89, 0.95, 
    0.99, 1, 0.9, 0.78, 0.84, 0.86, 0.71, 0.68, 0.65, 0.68, 0.73, 0.69, 0.72, 
    0.71, 0.68, 0.67, 0.67, 0.82, 0.99, 0.99, 0.99, 1, 0.99, 0.99, 1, 0.99, 
    1, 0.99, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.96, 0.92, 0.84, 0.75, 0.76, 0.77, 0.78, 0.76, 0.77, 0.75, 
    0.76, 0.73, 0.73, 0.7, 0.8, 0.81, 0.78, 0.73, 0.72, 0.76, 0.72, 0.74, 
    0.8, 0.67, 0.8, 0.8, 0.82, 0.9, 0.86, 0.89, 0.71, 0.7, 0.7, 0.69, 0.68, 
    0.7, 0.75, 0.67, 0.65, 0.63, 0.63, 0.63, 0.61, 0.59, 0.57, 0.57, 0.58, 
    0.6, 0.63, 0.64, 0.63, 0.63, 0.6, 0.58, 0.64, 0.68, 0.63, 0.69, 0.69, 
    0.69, 0.7, 0.65, 0.59, 0.65, 0.62, 0.63, 0.63, 0.61, 0.61, 0.6, 0.62, 
    0.59, 0.59, 0.66, 0.61, 0.66, 0.67, 0.67, 0.72, 0.66, 0.68, 0.65, 0.64, 
    0.65, 0.65, 0.7, 0.74, 0.78, 0.73, 0.6, 0.59, 0.6, 0.51, 0.48, 0.51, 
    0.55, 0.57, 0.6, 0.57, 0.57, 0.55, 0.61, 0.63, 0.62, 0.68, 0.72, 0.67, 
    0.63, 0.66, 0.62, 0.58, 0.59, 0.58, 0.56, 0.57, 0.6, 0.65, 0.64, 0.63, 
    0.67, 0.66, 0.65, 0.65, 0.64, 0.66, 0.7, 0.69, 0.68, 0.72, 0.74, 0.74, 
    0.75, 0.76, 0.74, 0.77, 0.77, 0.74, 0.73, 0.75, 0.77, 0.71, 0.74, 0.76, 
    0.74, 0.74, 0.72, 0.71, 0.73, 0.71, 0.73, 0.72, 0.7, 0.72, 0.71, 0.69, 
    0.68, 0.66, 0.66, 0.62, 0.62, 0.67, 0.62, 0.63, 0.63, 0.62, 0.64, 0.62, 
    0.67, 0.63, 0.66, 0.68, 0.67, 0.67, 0.7, 0.68, 0.7, 0.73, 0.72, 0.69, 
    0.69, 0.69, 0.71, 0.69, 0.7, 0.69, 0.7, 0.7, 0.69, 0.7, 0.69, 0.69, 0.7, 
    0.71, 0.69, 0.7, 0.71, 0.71, 0.7, 0.69, 0.72, 0.7, 0.68, 0.67, 0.69, 
    0.68, 0.68, 0.7, 0.67, 0.7, 0.65, 0.73, 0.73, 0.72, 0.7, 0.7, 0.71, 0.7, 
    0.73, 0.69, 0.61, 0.67, 0.65, 0.66, 0.67, 0.67, 0.66, 0.69, 0.66, 0.67, 
    0.75, 0.62, 0.57, 0.57, 0.55, 0.53, 0.57, 0.57, 0.56, 0.63, 0.58, 0.56, 
    0.58, 0.6, 0.62, 0.68, 0.68, 0.71, 0.71, 0.69, 0.67, 0.65, 0.68, 0.72, 
    0.73, 0.68, 0.64, 0.64, 0.64, 0.64, 0.64, 0.64, 0.61, 0.62, 0.63, 0.62, 
    0.62, 0.63, 0.66, 0.64, 0.65, 0.65, 0.67, 0.67, 0.69, 0.7, 0.69, 0.69, 
    0.69, 0.7, 0.71, 0.69, 0.67, 0.66, 0.66, 0.66, 0.66, 0.66, 0.65, 0.66, 
    0.65, 0.65, 0.67, 0.68, 0.68, 0.71, 0.74, 0.71, 0.65, 0.64, 0.65, 0.64, 
    0.63, 0.66, 0.63, 0.61, 0.64, 0.66, 0.63, 0.61, 0.55, 0.55, 0.52, 0.55, 
    0.5, 0.55, 0.61, 0.69, 0.62, 0.61, 0.62, 0.58, 0.58, 0.62, 0.63, 0.65, 
    0.64, 0.64, 0.63, 0.64, 0.65, 0.66, 0.59, 0.58, 0.59, 0.6, 0.61, 0.58, 
    0.53, 0.51, 0.58, 0.56, 0.55, 0.55, 0.58, 0.62, 0.65, 0.67, 0.64, 0.65, 
    0.67, 0.62, 0.61, 0.58, 0.68, 0.68, 0.66, 0.64, 0.65, 0.72, 0.77, 0.77, 
    0.7, 0.64, 0.66, 0.59, 0.66, 0.64, 0.62, 0.6, 0.6, 0.55, 0.55, 0.53, 
    0.55, 0.51, 0.49, 0.53, 0.53, 0.56, 0.57, 0.56, 0.55, 0.54, 0.52, 0.52, 
    0.52, 0.53, 0.54, 0.61, 0.64, 0.66, 0.63, 0.64, 0.66, 0.7, 0.84, 0.91, 
    0.93, 0.98, 0.97, 0.96, 0.98, 0.99, 0.96, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.89, 0.92, 0.82, 0.82, 0.83, 0.83, 0.82, 0.85, 0.85, 0.79, 0.83, 
    0.85, 0.78, 0.81, 0.95, 0.89, 0.86, 0.82, 0.81, 0.79, 0.75, 0.82, 0.76, 
    0.73, 0.61, 0.61, 0.7, 0.78, 1, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.97, 0.92, 0.9, 0.88, 0.92, 0.91, 0.92, 0.88, 0.81, 
    0.76, 0.75, 0.66, 0.64, 0.69, 0.73, 0.66, 0.65, 0.66, 0.66, 0.68, 0.68, 
    0.74, 0.85, 0.81, 0.78, 0.76, 0.81, 0.73, 0.73, 0.72, 0.72, 0.72, 0.71, 
    0.75, 0.78, 0.82, 0.89, 0.78, 0.84, 0.76, 0.79, 0.77, 0.77, 0.77, 0.8, 
    0.82, 0.83, 0.79, 0.85, 0.82, 0.81, 0.89, 0.86, 0.89, 0.9, 0.89, 0.86, 
    0.84, 0.87, 0.89, 0.89, 0.88, 0.91, 0.91, 0.91, 0.96, 0.99, 0.98, 0.99, 
    0.99, 0.86, 0.94, 0.82, 0.78, 0.74, 0.71, 0.74, 0.73, 0.65, 0.74, 0.74, 
    0.72, 0.99, 0.99, 1, 0.77, 0.72, 0.76, 0.74, 0.72, 0.71, 0.73, 0.88, 
    0.74, 0.75, 0.72, 0.74, 0.8, 0.89, 1, 1, 0.98, 0.84, 0.99, 0.99, 0.99, 
    0.99, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 1, 
    0.97, 1, 0.93, 0.87, 0.81, 0.77, 0.67, 0.76, 0.7, 0.7, 0.72, 0.7, 0.75, 
    0.77, 0.79, 0.79, 0.75, 0.75, 0.75, 0.74, 0.69, 0.76, 0.79, 0.84, 0.77, 
    0.76, 0.75, 0.76, 0.79, 0.75, 0.75, 0.74, 0.79, 0.74, 0.75, 0.76, 0.76, 
    0.72, 0.71, 0.67, 0.74, 0.71, 0.76, 0.7, 0.72, 0.76, 0.77, 0.83, 0.77, 
    0.78, 0.81, 0.83, 0.81, 0.81, 0.78, 0.8, 0.8, 0.78, 0.79, 0.83, 0.76, 
    0.73, 0.57, 0.59, 0.71, 0.68, 0.68, 0.71, 0.75, 0.75, 0.79, 0.72, 0.65, 
    0.63, 0.62, 0.58, 0.58, 0.59, 0.6, 0.65, 0.66, 0.7, 0.7, 0.71, 0.72, 
    0.73, 0.73, 0.74, 0.76, 0.88, 0.88, 0.82, 0.86, 0.83, 0.81, 0.85, 0.79, 
    0.85, 0.84, 0.83, 0.83, 0.87, 0.79, 0.78, 0.78, 0.8, 0.78, 0.78, 0.8, 
    0.79, 0.78, 0.81, 0.79, 0.76, 0.73, 0.73, 0.66, 0.61, 0.71, 0.62, 0.6, 
    0.66, 0.64, 0.62, 0.61, 0.6, 0.59, 0.6, 0.6, 0.56, 0.64, 0.62, 0.61, 
    0.59, 0.6, 0.61, 0.59, 0.59, 0.58, 0.58, 0.56, 0.52, 0.48, 0.49, 0.47, 
    0.42, 0.43, 0.45, 0.54, 0.5, 0.57, 0.46, 0.49, 0.53, 0.49, 0.49, 0.48, 
    0.54, 0.5, 0.53, 0.59, 0.6, 0.64, 0.65, 0.62, 0.64, 0.64, 0.65, 0.65, 
    0.61, 0.61, 0.62, 0.6, 0.61, 0.6, 0.58, 0.55, 0.47, 0.5, 0.46, 0.47, 
    0.48, 0.5, 0.51, 0.52, 0.59, 0.56, 0.56, 0.55, 0.55, 0.5, 0.5, 0.61, 
    0.55, 0.61, 0.6, 0.63, 0.62, 0.61, 0.66, 0.65, 0.63, 0.68, 0.65, 0.68, 
    0.62, 0.67, 0.7, 0.73, 0.73, 0.74, 0.76, 0.78, 0.8, 0.8, 0.79, 0.8, 0.81, 
    0.81, 0.8, 0.81, 0.79, 0.76, 0.77, 0.75, 0.74, 0.73, 0.69, 0.72, 0.71, 
    0.7, 0.69, 0.68, 0.72, 0.67, 0.69, 0.69, 0.74, 0.73, 0.74, 0.74, 0.81, 
    0.86, 0.9, 0.91, 0.94, 0.95, 0.93, 0.92, 0.74, 0.71, 0.62, 0.65, 0.64, 
    0.58, 0.58, 0.59, 0.63, 0.66, 0.69, 0.68, 0.7, 0.75, 0.83, 0.92, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.92, 0.81, 0.85, 0.83, 0.88, 0.82, 0.82, 0.83, 
    0.82, 0.85, 0.8, 0.78, 0.78, 0.82, 0.81, 0.77, 0.75, 0.83, 0.75, 0.74, 
    0.73, 0.68, 0.69, 0.71, 0.7, 0.7, 0.73, 0.72, 0.76, 0.76, 0.78, 0.81, 
    0.88, 0.87, 0.9, 0.98, 0.8, 0.87, 0.91, 0.89, 0.86, 0.89, 0.84, 0.8, 
    0.83, 0.88, 0.86, 0.87, 0.87, 0.83, 0.85, 0.91, 0.91, 0.98, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.9, 0.94, 0.94, 0.95, 0.87, 
    0.96, 0.99, 0.99, 0.97, 0.99, 0.96, 0.88, 0.85, 0.88, 0.91, 0.93, 0.84, 
    0.86, 0.89, 0.92, 0.99, 0.95, 0.81, 0.9, 0.74, 0.84, 0.84, 0.83, 0.74, 
    0.68, 0.72, 0.78, 0.76, 0.79, 0.81, 0.81, 0.75, 0.8, 0.81, 0.84, 0.77, 
    0.79, 0.79, 0.78, 0.83, 0.8, 0.9, 0.75, 0.82, 0.79, 0.76, 0.74, 0.81, 
    0.79, 0.81, 0.86, 0.93, 0.89, 0.8, 0.79, 0.81, 0.93, 0.78, 0.76, 0.75, 
    0.79, 0.83, 0.78, 0.73, 0.73, 0.79, 0.76, 0.75, 0.73, 0.73, 0.82, 0.95, 
    0.89, 0.85, 0.94, 0.93, 0.94, 0.82, 0.83, 0.77, 0.85, 0.92, 0.81, 0.8, 
    0.74, 0.71, 0.73, 0.74, 0.73, 0.74, 0.74, 0.73, 0.72, 0.71, 0.7, 0.7, 
    0.71, 0.69, 0.71, 0.7, 0.68, 0.65, 0.55, 0.47, 0.54, 0.5, 0.45, 0.41, 
    0.48, 0.45, 0.42, 0.41, 0.42, 0.43, 0.44, 0.45, 0.49, 0.53, 0.5, 0.46, 
    0.49, 0.48, 0.46, 0.47, 0.5, 0.52, 0.49, 0.55, 0.53, 0.52, 0.54, 0.56, 
    0.57, 0.58, 0.58, 0.58, 0.58, 0.61, 0.59, 0.59, 0.6, 0.63, 0.66, 0.63, 
    0.62, 0.63, 0.67, 0.69, 0.72, 0.74, 0.69, 0.68, 0.67, 0.68, 0.68, 0.67, 
    0.65, 0.61, 0.56, 0.61, 0.54, 0.57, 0.5, 0.48, 0.49, 0.55, 0.58, 0.66, 
    0.63, 0.61, 0.6, 0.65, 0.6, 0.64, 0.66, 0.64, 0.66, 0.65, 0.66, 0.65, 
    0.67, 0.68, 0.72, 0.72, 0.71, 0.72, 0.75, 0.74, 0.77, 0.76, 0.76, 0.75, 
    0.69, 0.66, 0.66, 0.68, 0.62, 0.61, 0.66, 0.5, 0.58, 0.59, 0.59, 0.57, 
    0.52, 0.45, 0.47, 0.51, 0.52, 0.49, 0.54, 0.6, 0.52, 0.54, 0.48, 0.51, 
    0.54, 0.56, 0.55, 0.51, 0.47, 0.47, 0.58, 0.49, 0.53, 0.59, 0.54, 0.61, 
    0.62, 0.59, 0.65, 0.64, 0.65, 0.66, 0.63, 0.63, 0.68, 0.72, 0.7, 0.67, 
    0.67, 0.56, 0.52, 0.52, 0.53, 0.48, 0.55, 0.49, 0.49, 0.57, 0.52, 0.5, 
    0.53, 0.54, 0.54, 0.54, 0.55, 0.56, 0.58, 0.51, 0.54, 0.53, 0.47, 0.47, 
    0.53, 0.53, 0.54, 0.54, 0.62, 0.64, 0.62, 0.64, 0.63, 0.64, 0.68, 0.69, 
    0.7, 0.69, 0.74, 0.75, 0.75, 0.74, 0.73, 0.76, 0.79, 0.76, 0.77, 0.8, 
    0.88, 0.96, 0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.8, 0.64, 0.66, 
    0.71, 0.72, 0.78, 0.81, 0.84, 0.9, 0.83, 0.81, 0.78, 0.74, 0.71, 0.67, 
    0.62, 0.68, 0.69, 0.72, 0.74, 0.71, 0.77, 0.79, 0.68, 0.88, 0.83, 0.77, 
    0.76, 0.8, 0.88, 0.83, 0.84, 0.82, 0.82, 0.79, 0.76, 0.77, 0.78, 0.95, 
    0.99, 0.63, 0.66, 0.66, 0.67, 0.99, 0.86, 0.92, 0.94, 0.84, 0.73, 0.65, 
    0.7, 0.69, 0.71, 0.63, 0.64, 0.63, 0.61, 0.56, 0.55, 0.55, 0.55, 0.55, 
    0.62, 0.63, 0.54, 0.54, 0.51, 0.54, 0.49, 0.53, 0.47, 0.53, 0.57, 0.51, 
    0.57, 0.59, 0.69, 0.73, 0.72, 0.7, 0.73, 0.71, 0.66, 0.59, 0.55, 0.52, 
    0.49, 0.48, 0.48, 0.46, 0.46, 0.47, 0.48, 0.51, 0.55, 0.57, 0.54, 0.55, 
    0.6, 0.55, 0.56, 0.56, 0.57, 0.57, 0.56, 0.51, 0.46, 0.5, 0.49, 0.49, 
    0.5, 0.51, 0.52, 0.5, 0.55, 0.55, 0.53, 0.58, 0.61, 0.62, 0.63, 0.66, 
    0.66, 0.65, 0.66, 0.62, 0.64, 0.65, 0.74, 0.66, 0.67, 0.7, 0.66, 0.72, 
    0.71, 0.69, 0.67, 0.66, 0.62, 0.68, 0.62, 0.66, 0.55, 0.63, 0.55, 0.56, 
    0.58, 0.58, 0.56, 0.6, 0.57, 0.6, 0.62, 0.62, 0.62, 0.62, 0.65, 0.64, 
    0.64, 0.61, 0.61, 0.62, 0.62, 0.62, 0.61, 0.64, 0.58, 0.6, 0.6, 0.6, 
    0.57, 0.56, 0.55, 0.57, 0.56, 0.57, 0.56, 0.56, 0.56, 0.53, 0.52, 0.52, 
    0.52, 0.58, 0.59, 0.66, 0.7, 0.73, 0.74, 0.77, 0.79, 0.82, 0.82, 0.82, 
    0.81, 0.79, 0.75, 0.75, 0.7, 0.69, 0.68, 0.65, 0.62, 0.63, 0.64, 0.64, 
    0.62, 0.6, 0.61, 0.63, 0.64, 0.63, 0.68, 0.67, 0.66, 0.66, 0.64, 0.65, 
    0.66, 0.66, 0.64, 0.64, 0.63, 0.66, 0.64, 0.64, 0.64, 0.62, 0.62, 0.62, 
    0.63, 0.62, 0.61, 0.6, 0.6, 0.57, 0.6, 0.62, 0.59, 0.54, 0.52, 0.45, 
    0.53, 0.58, 0.51, 0.48, 0.48, 0.53, 0.51, 0.55, 0.49, 0.54, 0.54, 0.53, 
    0.55, 0.56, 0.6, 0.61, 0.6, 0.58, 0.6, 0.62, 0.64, 0.61, 0.63, 0.64, 
    0.63, 0.62, 0.6, 0.56, 0.59, 0.57, 0.59, 0.57, 0.59, 0.64, 0.69, 0.61, 
    0.79, 0.91, 0.99, 0.96, 1, 0.99, 0.99, 0.99, 0.99, 0.92, 0.99, 1, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 1, 0.99, 0.99, 1, 
    0.79, 0.99, 0.99, 0.95, 0.88, 0.99, 0.99, 0.79, 0.82, 0.67, 0.77, 0.81, 
    0.72, 0.75, 0.77, 0.9, 0.89, 0.86, 0.89, 0.86, 0.86, 0.89, 0.89, 0.89, 
    0.83, 0.83, 0.89, 0.83, 0.97, 0.99, 0.99, 0.81, 0.93, 0.99, 0.96, 0.99, 
    0.99, 0.76, 0.68, 0.63, 0.61, 0.61, 0.59, 0.58, 0.58, 0.58, 0.58, 0.59, 
    0.61, 0.59, 0.59, 0.6, 0.6, 0.6, 0.59, 0.59, 0.62, 0.61, 0.62, 0.61, 0.6, 
    0.6, 0.6, 0.61, 0.59, 0.59, 0.59, 0.58, 0.57, 0.56, 0.55, 0.53, 0.55, 
    0.59, 0.6, 0.63, 0.65, 0.65, 0.64, 0.66, 0.65, 0.66, 0.66, 0.65, 0.66, 
    0.65, 0.63, 0.61, 0.59, 0.59, 0.61, 0.62, 0.64, 0.66, 0.65, 0.68, 0.69, 
    0.69, 0.7, 0.7, 0.69, 0.67, 0.65, 0.67, 0.64, 0.65, 0.64, 0.69, 0.64, 
    0.61, 0.62, 0.62, 0.63, 0.64, 0.67, 0.62, 0.64, 0.63, 0.63, 0.59, 0.61, 
    0.64, 0.62, 0.6, 0.61, 0.6, 0.62, 0.66, 0.6, 0.6, 0.6, 0.61, 0.6, 0.59, 
    0.63, 0.63, 0.65, 0.61, 0.64, 0.61, 0.63, 0.61, 0.64, 0.65, 0.64, 0.63, 
    0.64, 0.67, 0.65, 0.66, 0.64, 0.66, 0.67, 0.66, 0.67, 0.68, 0.66, 0.66, 
    0.67, 0.66, 0.68, 0.68, 0.65, 0.66, 0.69, 0.66, 0.65, 0.61, 0.62, 0.6, 
    0.61, 0.63, 0.61, 0.64, 0.65, 0.57, 0.61, 0.58, 0.59, 0.58, 0.65, 0.71, 
    0.71, 0.69, 0.67, 0.72, 0.73, 0.7, 0.75, 0.69, 0.6, 0.5, 0.42, 0.48, 
    0.42, 0.42, 0.47, 0.35, 0.35, 0.34, 0.35, 0.38, 0.38, 0.38, 0.43, 0.6, 
    0.64, 0.59, 0.64, 0.65, 0.52, 0.53, 0.43, 0.6, 0.63, 0.62, 0.65, 0.65, 
    0.63, 0.59, 0.61, 0.74, 0.87, 0.76, 0.82, 0.88, 0.8, 0.92, 0.99, 0.99, 
    0.99, 0.98, 0.78, 0.71, 0.72, 0.68, 0.65, 0.61, 0.61, 0.58, 0.58, 0.62, 
    0.66, 0.67, 0.67, 0.67, 0.69, 0.69, 0.71, 0.73, 0.74, 0.71, 0.74, 0.75, 
    0.73, 0.7, 0.74, 0.7, 0.58, 0.71, 0.65, 0.58, 0.55, 0.62, 0.65, 0.56, 
    0.59, 0.57, 0.56, 0.57, 0.55, 0.51, 0.55, 0.53, 0.52, 0.56, 0.54, 0.46, 
    0.57, 0.5, 0.58, 0.44, 0.44, 0.54, 0.49, 0.47, 0.51, 0.54, 0.54, 0.51, 
    0.53, 0.6, 0.62, 0.55, 0.54, 0.56, 0.56, 0.56, 0.46, 0.44, 0.52, 0.52, 
    0.52, 0.53, 0.52, 0.51, 0.52, 0.56, 0.57, 0.54, 0.57, 0.58, 0.59, 0.59, 
    0.62, 0.57, 0.6, 0.56, 0.57, 0.66, 0.68, 0.67, 0.63, 0.66, 0.61, 0.66, 
    0.67, 0.68, 0.68, 0.67, 0.66, 0.65, 0.64, 0.58, 0.66, 0.69, 0.66, 0.69, 
    0.73, 0.75, 0.71, 0.64, 0.61, 0.62, 0.58, 0.55, 0.58, 0.6, 0.59, 0.59, 
    0.62, 0.64, 0.71, 0.71, 0.73, 0.96, 0.97, 0.92, 0.99, 0.99, 0.99, 1, 
    0.99, 0.99, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.95, 0.94, 0.93, 
    0.99, 0.94, 0.87, 0.88, 0.89, 0.89, 0.88, 0.88, 0.88, 0.87, 0.88, 0.89, 
    0.88, 0.88, 0.87, 0.86, 0.87, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 0.88, 
    0.9, 0.9, 0.89, 0.89, 0.89, 0.89, 0.9, 0.87, 0.86, 0.88, 0.86, 0.84, 
    0.84, 0.82, 0.85, 0.87, 0.88, 0.89, 0.88, 0.84, 0.87, 0.89, 0.9, 0.9, 
    0.91, 0.9, 0.88, 0.89, 0.87, 0.87, 0.87, 0.88, 0.87, 0.87, 0.88, 0.88, 
    0.9, 0.92, 0.92, 0.92, 0.93, 0.92, 0.92, 0.92, 0.92, 0.91, 0.91, 0.9, 
    0.91, 0.9, 0.89, 0.88, 0.86, 0.86, 0.84, 0.87, 0.9, 0.89, 0.87, 0.87, 
    0.85, 0.86, 0.84, 0.84, 0.84, 0.84, 0.84, 0.83, 0.84, 0.84, 0.84, 0.85, 
    0.87, 0.88, 0.8, 0.8, 0.82, 0.84, 0.87, 0.9, 0.85, 0.82, 0.83, 0.86, 
    0.84, 0.82, 0.89, 0.88, 0.89, 0.88, 0.88, 0.9, 0.89, 0.89, 0.87, 0.87, 
    0.87, 0.86, 0.83, 0.83, 0.83, 0.83, 0.83, 0.82, 0.83, 0.83, 0.84, 0.84, 
    0.85, 0.85, 0.85, 0.85, 0.85, 0.86, 0.85, 0.85, 0.83, 0.81, 0.81, 0.83, 
    0.83, 0.82, 0.84, 0.84, 0.83, 0.78, 0.77, 0.76, 0.77, 0.78, 0.77, 0.74, 
    0.73, 0.77, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 0.76, 
    0.76, 0.77, 0.77, 0.76, 0.76, 0.75, 0.75, 0.75, 0.74, 0.75, 0.75, 0.76, 
    0.76, 0.78, 0.78, 0.78, 0.79, 0.8, 0.83, 0.81, 0.8, 0.8, 0.79, 0.77, 
    0.77, 0.75, 0.72, 0.71, 0.7, 0.68, 0.64, 0.63, 0.64, 0.65, 0.67, 0.68, 
    0.67, 0.66, 0.67, 0.68, 0.68, 0.68, 0.71, 0.75, 0.76, 0.74, 0.77, 0.84, 
    0.85, 0.83, 0.83, 0.82, 0.81, 0.8, 0.8, 0.8, 0.81, 0.83, 0.84, 0.84, 
    0.85, 0.87, 0.88, 0.88, 0.87, 0.86, 0.87, 0.88, 0.87, 0.85, 0.83, 0.83, 
    0.83, 0.8, 0.81, 0.82, 0.82, 0.82, 0.84, 0.85, 0.84, 0.85, 0.87, 0.88, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 0.99, 0.92, 0.84, 0.89, 
    0.91, 0.77, 0.82, 0.79, 0.73, 0.72, 0.68, 0.75, 0.99, 0.99, 0.99, 0.99, 
    0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 0.78, 0.71, 0.68, 0.66, 
    0.79, 0.67, 0.67, 0.67, 0.66, 0.67, 0.66, 0.67, 0.66, 0.67, 0.68, 0.67, 
    0.72, 0.72, 0.73, 0.73, 0.74, 0.76, 0.77, 0.76, 0.76, 0.75, 0.75, 0.76, 
    0.75, 0.76, 0.76, 0.76, 0.76, 0.75, 0.75, 0.75, 0.69, 0.73, 0.77, 0.71, 
    0.71, 0.76, 0.77, 0.76, 0.74, 0.69, 0.8, 0.73, 0.71, 0.72, 0.72, 0.73, 
    0.72, 0.7, 0.68, 0.69, 0.67, 0.67, 0.62, 0.62, 0.63, 0.6, 0.65, 0.63, 
    0.56, 0.56, 0.58, 0.57, 0.52, 0.51, 0.56, 0.6, 0.64, 0.67, 0.68, 0.69, 
    0.55, 0.52, 0.56, 0.58, 0.54, 0.57, 0.55, 0.54, 0.54, 0.53, 0.57, 0.54, 
    0.53, 0.53, 0.52, 0.54, 0.53, 0.52, 0.53, 0.72, 0.57, 0.52, 0.52, 0.54, 
    0.51, 0.56, 0.52, 0.56, 0.61, 0.56, 0.58, 0.63, 0.62, 0.61, 0.65, 0.67, 
    0.67, 0.68, 0.67, 0.72, 0.67, 0.77, 0.77, 0.68, 0.72, 0.73, 0.66, 0.65, 
    0.7, 0.65, 0.63, 0.62, 0.64, 0.62, 0.61, 0.67, 0.62, 0.65, 0.61, 0.67, 
    0.66, 0.69, 0.65, 0.73, 0.58, 0.73, 0.66, 0.67, 0.64, 0.71, 0.78, 0.77, 
    0.72, 0.76, 0.8, 0.78, 0.76, 0.69, 0.67, 0.71, 0.73, 0.7, 0.73, 0.59, 
    0.73, 0.57, 0.6, 0.71, 0.56, 0.57, 0.54, 0.72, 0.6, 0.61, 0.73, 0.55, 
    0.52, 0.73, 0.51, 0.74, 0.47, 0.54, 0.51, 0.53, 0.57, 0.63, 0.62, 0.69, 
    0.69, 0.74, 0.72, 0.74, 0.76, 0.77, 0.72, 0.74, 0.72, 0.74, 0.76, 0.73, 
    0.72, 0.69, 0.65, 0.59, 0.6, 0.58, 0.58, 0.56, 0.63, 0.67, 0.66, 0.74, 
    0.73, 0.73, 0.75, 0.74, 0.71, 0.74, 0.74, 0.78, 0.69, 0.68, 0.63, 0.62, 
    0.67, 0.63, 0.65, 0.69, 0.69, 0.7, 0.71, 0.73, 0.77, 0.79, 0.79, 0.89, 
    0.95, 0.99, 0.99, 0.87, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.99, 
    0.99, 1, 0.99, 0.92, 0.85, 0.95, 0.91, 0.94, 0.94, 0.87, 0.86, 0.87, 
    0.81, 0.93, 0.99, 0.92, 0.99, 0.99, 0.99, 1, 0.88, 0.99, 0.99, 0.91, 
    0.85, 0.84, 0.92, 0.85, 0.93, 0.96, 0.87, 0.95, 0.97, 0.99, 0.99, 0.99, 
    1, 1, 1, 0.99, 0.99, 0.99, 0.99, 0.94, 0.99, 0.99, 1, 0.99, 1, 0.99, 
    0.99, 0.99, 0.99, 0.83, 0.73, 0.73, 0.76, 0.88, 0.77, 0.91, 0.96, 0.86, 
    0.83, 0.87, 0.86, 0.96, 0.93, 0.88, 0.81, 0.75, 0.71, 0.82, 0.83, 0.82, 
    0.8, 0.78, 0.74, 0.7, 0.67, 0.67, 0.71, 0.7, 0.74, 0.71, 0.71, 0.7, 0.7, 
    0.7, 0.7, 0.68, 0.67, 0.69, 0.68, 0.69, 0.7, 0.7, 0.71, 0.57, 0.56, 0.61, 
    0.65, 0.65, 0.64, 0.63, 0.63, 0.66, 0.63, 0.6, 0.58, 0.69, 0.69, 0.69, 
    0.58, 0.59, 0.69, 0.69, 0.69, 0.54, 0.7, 0.56, 0.7, 0.55, 0.61, 0.58, 
    0.74, 0.77, 0.57, 0.6, 0.6, 0.6, 0.57, 0.56, 0.57, 0.57, 0.59, 0.77, 
    0.61, 0.59, 0.58, 0.59, 0.57, 0.57, 0.58, 0.54, 0.54, 0.51, 0.49, 0.46, 
    0.47, 0.48, 0.55, 0.56, 0.6, 0.56, 0.56, 0.57, 0.54, 0.7, 0.58, 0.55, 
    0.52, 0.54, 0.54, 0.56, 0.55, 0.53, 0.55, 0.58, 0.57, 0.57, 0.56, 0.56, 
    0.54, 0.55, 0.55, 0.56, 0.56, 0.46, 0.5, 0.49, 0.51, 0.67, 0.49, 0.51, 
    0.5, 0.51, 0.52, 0.66, 0.67, 0.52, 0.51, 0.5, 0.48, 0.48, 0.51, 0.53, 
    0.54, 0.56, 0.61, 0.63, 0.63, 0.64, 0.64, 0.63, 0.68, 0.61, 0.68, 0.72, 
    0.63, 0.59, 0.58, 0.51, 0.53, 0.56, 0.53, 0.57, 0.62, 0.64, 0.71, 0.74, 
    0.7, 0.79, 0.79, 0.8, 0.92, 0.99, 0.85, 0.88, 0.81, 0.91, 0.89, 0.82, 
    0.91, 0.91, 0.86, 0.93, 0.9, 0.89, 0.83, 0.49, 0.48, 0.44, 0.45, 0.44, 
    0.49, 0.5, 0.48, 0.5, 0.56, 0.56, 0.58, 0.59, 0.58, 0.65, 0.61, 0.56, 
    0.43, 0.48, 0.55, 0.66, 0.78, 0.64, 0.64, 0.65, 0.65, 0.69, 0.6, 0.62, 
    0.6, 0.67, 0.67, 0.7, 0.74, 0.67, 0.7, 0.67, 0.68, 0.69, 0.72, 0.84, 
    0.75, 0.77, 0.87, 0.76, 0.7, 0.79, 0.67, 0.66, 0.66, 0.64, 0.63, 0.64, 
    0.61, 0.59, 0.68, 0.71, 0.71, 0.85, 0.84, 0.72, 0.8, 0.85, 0.72, 0.82, 
    0.8, 0.7, 0.67, 0.7, 0.68, 0.6, 0.6, 0.61, 0.58, 0.63, 0.61, 0.61, 0.65, 
    0.66, 0.74, 0.69, 0.82, 0.86, 0.84, 0.82, 0.83, 0.83, 0.82, 0.77, 0.77, 
    0.82, 0.81, 0.78, 0.75, 0.76, 0.7, 0.7, 0.68, 0.67, 0.63, 0.67, 0.66, 
    0.68, 0.69, 0.72, 0.74, 0.73, 0.75, 0.79, 0.79, 0.81, 0.79, 0.79, 0.74, 
    0.74, 0.77, 0.7, 0.7, 0.69, 0.66, 0.65, 0.62, 0.6, 0.61, 0.57, 0.57, 
    0.57, 0.57, 0.58, 0.58, 0.57, 0.59, 0.64, 0.7, 0.68, 0.72, 0.72, 0.69, 
    0.71, 0.66, 0.7, 0.65, 0.64, 0.67, 0.63, 0.64, 0.63, 0.58, 0.63, 0.75, 
    0.75, 0.79, 0.83, 0.91, 0.91, 0.86, 0.92, 0.89, 0.82, 0.97, 0.93, 0.94, 
    0.75, 0.71, 0.68, 0.7, 0.75, 0.8, 0.89, 0.78, 0.67, 0.68, 0.68, 0.7, 
    0.74, 0.7, 0.7, 0.66, 0.71, 0.92, 0.79, 0.75, 0.69, 0.69, 0.69, 0.73, 
    0.67, 0.63, 0.63, 0.7, 0.72, 0.89, 0.76, 0.71, 0.71, 0.69, 0.77, 0.77, 
    0.76, 0.68, 0.99, 0.78, 0.76, 0.73, 0.8, 0.75, 0.75, 0.76, 0.74, 0.89, 
    0.81, 0.73, 0.8, 0.84, 0.9, 0.87, 0.85, 0.84, 0.74, 0.77, 0.98, 0.8, 
    0.77, 0.8, 0.76, 0.78, 0.64, 0.6, 0.71, 0.71, 0.71, 0.6, 0.61, 0.63, 
    0.74, 0.71, 0.67, 0.75, 0.79, 0.75, 0.79, 1, 0.97, 1, 0.75, 0.99, 0.89, 
    0.88, 0.82, 0.7, 0.58, 0.64, 0.62, 0.61, 0.61, 0.64, 0.63, 0.64, 0.68, 
    0.68, 0.68, 0.68, 0.65, 0.71, 0.78, 0.76, 0.78, 0.82, 0.87, 0.8, 0.77, 
    0.79, 0.79, 0.79, 0.98, 0.88, 0.91, 0.85, 0.91, 0.94, 0.99, 0.99, 0.99, 
    0.99, 0.87, 0.77, 0.75, 0.68, 0.71, 0.72, 0.76, 0.68, 0.77, 0.73, 0.69, 
    0.69, 0.69, 0.6, 0.69, 0.64, 0.62, 0.59, 0.52, 0.53, 0.56, 0.54, 0.56, 
    0.6, 0.67, 0.63, 0.7, 0.72, 0.7, 0.72, 0.67, 0.7, 0.74, 0.75, 0.67, 0.64, 
    0.65, 0.65, 0.68, 0.62, 0.64, 0.53, 0.61, 0.61, 0.64, 0.63, 0.7, 0.72, 
    0.74, 0.75, 0.74, 0.8, 0.81, 0.78, 0.8, 0.78, 0.68, 0.62, 0.67, 0.66, 
    0.68, 0.65, 0.64, 0.63, 0.61, 0.68, 0.69, 0.73, 0.72, 0.69, 0.64, 0.61, 
    0.61, 0.57, 0.59, 0.57, 0.58, 0.57, 0.6, 0.58, 0.58, 0.57, 0.59, 0.58, 
    0.59, 0.58, 0.58, 0.58, 0.56, 0.57, 0.6, 0.61, 0.58, 0.65, 0.61, 0.58, 
    0.53, 0.55, 0.55, 0.62, 0.62, 0.69, 0.7, 0.68, 0.69, 0.71, 0.68, 0.69, 
    0.66, 0.65, 0.69, 0.72, 0.7, 0.69, 0.58, 0.53, 0.59, 0.42, 0.42, 0.46, 
    0.48, 0.54, 0.53, 0.37, 0.43, 0.44, 0.44, 0.45, 0.5, 0.51, 0.5, 0.58, 
    0.57, 0.56, 0.57, 0.58, 0.61, 0.65, 0.66, 0.66, 0.62, 0.63, 0.67, 0.66, 
    0.65, 0.65, 0.56, 0.57, 0.54, 0.53, 0.54, 0.54, 0.61, 0.57, 0.6, 0.54, 
    0.57, 0.6, 0.58, 0.6, 0.5, 0.53, 0.55, 0.54, 0.55, 0.63, 0.6, 0.55, 0.58, 
    0.64, 0.53, 0.61, 0.61, 0.53, 0.52, 0.5, 0.52, 0.54, 0.5, 0.53, 0.54, 
    0.53, 0.6, 0.58, 0.58, 0.59, 0.64, 0.65, 0.62, 0.59, 0.6, 0.57, 0.6, 
    0.62, 0.55, 0.56, 0.62, 0.61, 0.64, 0.67, 0.69, 0.71, 0.67, 0.66, 0.64, 
    0.64, 0.57, 0.64, 0.62, 0.65, 0.63, 0.63, 0.65, 0.68, 0.72, 0.72, 0.74, 
    0.72, 0.7, 0.67, 0.58, 0.55, 0.62, 0.64, 0.57, 0.59, 0.68, 0.68, 0.67, 
    0.68, 0.69, 0.73, 0.76, 0.77, 0.69, 0.68, 0.67, 0.7, 0.66, 0.58, 0.6, 
    0.64, 0.67, 0.64, 0.61, 0.69, 0.61, 0.66, 0.65, 0.75, 0.76, 0.76, 0.7, 
    0.65, 0.64, 0.59, 0.56, 0.54, 0.54, 0.53, 0.5, 0.51, 0.54, 0.57, 0.59, 
    0.57, 0.61, 0.63, 0.62, 0.58, 0.55, 0.54, 0.58, 0.6, 0.56, 0.61, 0.64, 
    0.71, 0.71, 0.74, 0.74, 0.77, 0.77, 0.81, 0.86, 0.88, 0.89, 0.82, 0.82, 
    0.8, 0.77, 0.68, 0.64, 0.71, 0.65, 0.68, 0.68, 0.66, 0.64, 0.69, 0.71, 
    0.67, 0.63, 0.69, 0.7, 0.73, 0.72, 0.71, 0.75, 0.79, 0.74, 0.74, 0.73, 
    0.74, 0.76, 0.63, 0.75, 0.74, 0.68, 0.82, 0.81, 0.86, 0.77, 0.73, 0.65, 
    0.76, 0.68, 0.61, 0.7, 0.78, 0.68, 0.64, 0.63, 0.54, 0.56, 0.53, 0.49, 
    0.44, 0.46, 0.49, 0.5, 0.46, 0.47, 0.55, 0.52, 0.51, 0.58, 0.59, 0.61, 
    0.6, 0.59, 0.56, 0.63, 0.53, 0.49, 0.48, 0.47, 0.47, 0.46, 0.45, 0.51, 
    0.51, 0.51, 0.52, 0.49, 0.52, 0.56, 0.57, 0.63, 0.63, 0.68, 0.69, 0.73, 
    0.77, 0.75, 0.72, 0.69, 0.66, 0.56, 0.58, 0.52, 0.58, 0.58, 0.51, 0.47, 
    0.52, 0.51, 0.49, 0.6, 0.67, 0.59, 0.64, 0.67, 0.68, 0.7, 0.71, 0.67, 
    0.66, 0.68, 0.68, 0.65, 0.65, 0.67, 0.66, 0.65, 0.64, 0.6, 0.63, 0.58, 
    0.56, 0.63, 0.63, 0.67, 0.67, 0.64, 0.65, 0.67, 0.69, 0.66, 0.72, 0.69, 
    0.71, 0.65, 0.65, 0.66, 0.64, 0.67, 0.67, 0.6, 0.69, 0.68, 0.73, 0.71, 
    0.65, 0.68, 0.68, 0.68, 0.65, 0.67, 0.65, 0.7, 0.72, 0.7, 0.69, 0.7, 
    0.66, 0.65, 0.68, 0.6, 0.62, 0.65, 0.62, 0.64, 0.66, 0.65, 0.62, 0.57, 
    0.63, 0.7, 0.71, 0.72, 0.73, 0.73, 0.75, 0.76, 0.78, 0.7, 0.68, 0.64, 
    0.69, 0.68, 0.67, 0.67, 0.66, 0.64, 0.66, 0.67, 0.66, 0.69, 0.72, 0.73, 
    0.81, 0.83, 0.84, 0.85, 0.86, 0.87, 0.88, 0.88, 0.88, 0.87, 0.86, 0.83, 
    0.76, 0.76, 0.73, 0.72, 0.74, 0.76, 0.75, 0.82, 0.85, 0.82, 0.87, 0.88, 
    0.86, 0.86, 0.9, 0.88, 0.85, 0.83, 0.88, 0.87, 0.84, 0.8, 0.7, 0.84, 
    0.84, 0.74, 0.82, 0.89, 0.87, 0.95, 0.99, 1, 1, 1, 0.99, 1, 0.78, 0.89, 
    0.93, 0.88, 0.91, 0.95, 1, 0.99, 0.95, 1, 0.99, 0.94, 0.99, 0.99, 0.89, 
    0.77, 0.74, 0.83, 0.98, 0.97, 0.85, 0.77, 0.78, 0.85, 0.83, 0.74, 0.78, 
    0.69, 0.66, 0.69, 0.68, 0.65, 0.62, 0.63, 0.67, 0.68, 0.7, 0.71, 0.67, 
    0.7, 0.62, 0.71, 0.71, 0.73, 0.74, 0.7, 0.66, 0.64, 0.63, 0.63, 0.64, 
    0.66, 0.66, 0.61, 0.66, 0.64, 0.67, 0.7, 0.71, 0.76, 0.85, 0.9, 0.98, 
    0.99, 0.99, 0.99, 0.99, 0.99, 1, 1, 0.99, 0.89, 0.98, 0.95, 0.86, 0.78, 
    0.74, 0.72, 0.73, 0.71, 0.69, 0.75, 0.79, 0.74, 0.89, 0.9, 0.9, 0.89, 
    0.77, 0.87, 0.86, 0.81, 0.62, 0.67, 0.53, 0.64, 0.59, 0.62, 0.68, 0.56, 
    0.65, 0.62, 0.65, 0.69, 0.67, 0.71, 0.73, 0.74, 0.75, 0.77, 0.84, 0.82, 
    0.83, 0.8, 0.77, 0.73, 0.69, 0.66, 0.65, 0.65, 0.64, 0.67, 0.62, 0.66, 
    0.68, 0.7, 0.64, 0.62, 0.68, 0.73, 0.71, 0.71, 0.7, 0.71, 0.71, 0.69, 
    0.7, 0.73, 0.72, 0.71, 0.67, 0.7, 0.64, 0.67, 0.61, 0.6, 0.6, 0.64, 0.64, 
    0.63, 0.6, 0.59, 0.61, 0.61, 0.6, 0.61, 0.65, 0.65, 0.61, 0.62, 0.59, 
    0.63, 0.62, 0.62, 0.64, 0.64, 0.63, 0.62, 0.63, 0.72, 0.76, 0.79, 0.82, 
    0.74, 0.72, 0.59, 0.66, 0.6, 0.62, 0.65, 0.67, 0.63, 0.64, 0.77, 0.81, 
    0.89, 0.86, 0.8, 0.79, 0.73, 0.7, 0.6, 0.6, 0.59, 0.65, 0.64, 0.63, 0.65, 
    0.71, 0.68, 0.7, 0.64, 0.67, 0.69, 0.72, 0.66, 0.66, 0.62, 0.61, 0.61, 
    0.59, 0.56, 0.53, 0.6, 0.63, 0.61, 0.52, 0.59, 0.61, 0.66, 0.65, 0.78, 
    0.86, 0.86, 0.89, 0.73, 0.69, 0.72, 0.71, 0.65, 0.56, 0.59, 0.58, 0.58, 
    0.57, 0.53, 0.57, 0.57, 0.6, 0.6, 0.62, 0.63, 0.65, 0.76, 0.74, 0.72, 
    0.73, 0.81, 0.8, 0.76, 0.74, 0.76, 0.74, 0.72, 0.69, 0.69, 0.67, 0.7, 
    0.64, 0.58, 0.64, 0.65, 0.64, 0.65, 0.74, 0.76, 0.77, 0.83, 0.77, 0.64, 
    0.79, 0.77, 0.82, 0.83, 0.78, 0.68, 0.69, 0.65, 0.73, 0.78, 0.8, 0.76, 
    0.74, 0.76, 0.73, 0.84, 0.73, 0.77, 0.78, 0.79, 0.79, 0.78, 0.75, 0.68, 
    0.75, 0.74, 0.71, 0.71, 0.75, 0.73, 0.76, 0.78, 0.71, 0.79, 0.72, 0.66, 
    0.68, 0.67, 0.7, 0.72, 0.74, 0.78, 0.73, 0.74, 0.72, 0.78, 0.79, 0.79, 
    0.83, 0.78, 0.82, 0.77, 0.75, 0.73, 0.72, 0.68, 0.65, 0.64, 0.63, 0.66, 
    0.58, 0.61, 0.64, 0.64, 0.65, 0.68, 0.67, 0.69, 0.71, 0.75, 0.76, 0.8, 
    0.81, 0.85, 0.82, 0.73, 0.7, 0.69, 0.66, 0.64, 0.62, 0.59, 0.58, 0.62, 
    0.61, 0.63, 0.63, 0.62, 0.63, 0.65, 0.65, 0.67, 0.69, 0.71, 0.71, 0.71, 
    0.72, 0.67, 0.9, 0.72, 0.71, 0.74, 0.68, 0.72, 0.62, 0.61, 0.61, 0.6, 
    0.58, 0.63, 0.6, 0.6, 0.62, 0.64, 0.67, 0.66, 0.63, 0.63, 0.63, 0.65, 
    0.66, 0.66, 0.63, 0.69, 0.69, 0.66, 0.69, 0.63, 0.65, 0.73, 0.65, 0.64, 
    0.64, 0.63, 0.56, 0.58, 0.56, 0.6, 0.65, 0.67, 0.65, 0.66, 0.74, 0.72, 
    0.64, 0.63, 0.6, 0.61, 0.61, 0.63, 0.65, 0.73, 0.69, 0.68, 0.66, 0.73, 
    0.71, 0.7, 0.7, 0.64, 0.63, 0.67, 0.68, 0.65, 0.59, 0.56, 0.62, 0.59, 
    0.57, 0.6, 0.62, 0.64, 0.59, 0.64, 0.59, 0.57, 0.58, 0.6, 0.56, 0.53, 
    0.58, 0.61, 0.64, 0.63, 0.63, 0.64, 0.6, 0.61, 0.64, 0.65, 0.63, 0.67, 
    0.68, 0.63, 0.63, 0.62, 0.68, 0.6, 0.66, 0.66, 0.68, 0.7, 0.64, 0.68, 
    0.64, 0.64, 0.65, 0.67, 0.67, 0.64, 0.71, 0.82, 0.94, 0.93, 0.91, 0.96, 
    0.99, 0.97, 0.9, 0.96, 0.97, 0.92, 0.88, 0.76, 0.77, 0.71, 0.6, 0.6, 
    0.55, 0.72, 0.7, 0.66, 0.96, 0.79, 0.63, 0.6, 0.62, 0.72, 0.79, 0.78, 
    0.76, 1, 0.83, 0.83, 0.85, 0.81, 0.83, 0.84, 0.86, 0.78, 0.81, 0.75, 
    0.72, 0.75, 0.76, 0.79, 0.86, 0.92, 0.9, 0.89, 0.99, 1, 1, 1, 1, 0.96, 
    0.89, 0.79, 0.74, 0.65, 0.68, 0.65, 0.65, 0.64, 0.62, 0.67, 0.65, 0.6, 
    0.66, 0.67, 0.65, 0.69, 0.68, 0.65, 0.63, 0.63, 0.64, 0.67, 0.68, 0.67, 
    0.66, 0.68, 0.72, 0.71, 0.69, 0.66, 0.65, 0.63, 0.65, 0.61, 0.63, 0.67, 
    0.69, 0.69, 0.7, 0.71, 0.72, 0.69, 0.67, 0.66, 0.7, 0.69, 0.67, 0.71, 
    0.66, 0.62, 0.62, 0.66, 0.68, 0.61, 0.65, 0.63, 0.63, 0.67, 0.68, 0.8, 
    0.73, 0.66, 0.77, 0.89, 0.87, 0.99, 0.99, 0.74, 0.7, 0.68, 0.62, 0.61, 
    0.64, 0.62, 0.62, 0.64, 0.67, 0.68, 0.66, 0.66, 0.67, 0.62, 0.65, 0.65, 
    0.62, 0.66, 0.69, 0.99, 1, 1, 0.65, 0.67, 0.66, 0.69, 0.69, 0.69, 0.64, 
    0.63, 0.58, 0.55, 0.6, 0.64, 0.68, 0.68, 0.69, 0.67, 0.67, 0.66, 0.68, 
    0.71, 0.72, 0.68, 0.71, 0.68, 0.64, 0.66, 0.6, 0.62, 0.62, 0.68, 0.65, 
    0.63, 0.63, 0.62, 0.62, 0.61, 0.61, 0.67, 0.57, 0.65, 0.63, 0.61, 0.64, 
    0.63, 0.64, 0.66, 0.67, 0.68, 0.79, 0.69, 0.64, 0.66, 0.62, 0.63, 0.78, 
    0.69, 0.68, 0.73, 0.75, 0.93, 0.92, 0.69, 0.78, 0.65, 0.65, 0.65, 0.63, 
    0.85, 0.81, 0.75, 0.97, 1, 0.74, 0.74, 1, 0.99, 0.99, 1, 0.83, 0.79, 
    0.76, 0.73, 0.99, 1, 0.74, 0.74, 0.73, 0.7, 0.71, 0.68, 0.72, 0.81, 0.78, 
    0.88, 0.87, 0.9, 0.91, 0.87, 0.89, 0.91, 0.91, 0.91, 0.91, 0.92, 0.91, 
    0.88, 0.87, 0.86, 0.85, 0.84, 0.8, 0.85, 0.86, 0.9, 0.87, 0.84, 0.88, 
    0.9, 0.9, 0.89, 0.85, 0.82, 0.83, 0.81, 0.82, 0.83, 0.84, 0.79, 0.76, 
    0.75, 0.78, 0.75, 0.72, 0.72, 0.72, 0.7, 0.68, 0.66, 0.64, 0.65, 0.64, 
    0.65, 0.66, 0.67, 0.66, 0.64, 0.63, 0.68, 0.72, 0.71, 0.7, 0.69, 0.68, 
    0.65, 0.65, 0.66, 0.69, 0.77, 0.68, 0.7, 0.71, 0.62, 0.66, 0.78, 0.72, 
    0.81, 0.78, 0.78, 0.84, 0.85, 0.86, 0.87, 0.87, 0.83, 0.85, 0.91, 0.88, 
    0.91, 0.82, 0.77, 0.66, 0.63, 0.64, 0.71, 0.66, 0.66, 0.63, 0.63, 0.64, 
    0.62, 0.66, 0.74, 0.78, 0.81, 0.81, 0.79, 0.67, 0.78, 0.78, 0.66, 0.62, 
    0.64, 0.74, 0.73, 0.74, 0.72, 0.74, 0.72, 0.69, 0.61, 0.6, 0.67, 0.63, 
    0.66, 0.74, 0.75, 0.65, 0.63, 0.62, 0.66, 0.66, 0.66, 0.67, 0.63, 0.58, 
    0.54, 0.54, 0.53, 0.51, 0.51, 0.51, 0.5, 0.53, 0.57, 0.53, 0.55, 0.58, 
    0.56, 0.65, 0.57, 0.59, 0.62, 0.64, 0.64, 0.62, 0.62, 0.62, 0.61, 0.64, 
    0.61, 0.59, 0.6, 0.61, 0.75, 0.74, 0.76, 0.83, 0.79, 0.62, 0.75, 0.64, 
    0.61, 0.64, 0.65, 0.65, 0.66, 0.69, 0.72, 0.68, 0.68, 0.7, 0.72, 0.65, 
    0.73, 0.74, 0.8, 0.74, 0.71, 0.7, 0.68, 0.84, 0.76, 0.63, 0.61, 0.64, 
    0.72, 0.69, 0.65, 0.68, 0.68, 0.73, 0.75, 0.75, 0.78, 0.75, 0.73, 0.71, 
    0.69, 0.73, 0.71, 0.74, 0.68, 0.62, 0.69, 0.68, 0.66, 0.62, 0.67, 0.71, 
    0.71, 0.72, 0.71, 0.63, 0.69, 0.69, 0.71, 0.74, 0.76, 0.75, 0.75, 0.73, 
    0.74, 0.77, 0.77, 0.77, 0.79, 0.64, 0.69, 0.63, 0.59, 0.59, 0.59, 0.69, 
    0.65, 0.66, 0.67, 0.65, 0.65, 0.68, 0.66, 0.67, 0.67, 0.67, 0.67, 0.69, 
    0.7, 0.73, 0.78, 0.8, 0.8, 0.81, 0.86, 0.85, 0.85, 0.89, 0.87, 0.89, 
    0.88, 0.81, 0.77, 0.83, 0.8, 0.73, 0.7, 0.71, 0.74, 0.76, 0.73, 0.65, 
    0.67, 0.67, 0.62, 0.58, 0.58, 0.62, 0.59, 0.59, 0.56, 0.61, 0.58, 0.52, 
    0.52, 0.54, 0.49, 0.49, 0.56, 0.54, 0.58, 0.57, 0.61, 0.58, 0.58, 0.59, 
    0.67, 0.69, 0.71, 0.7, 0.64, 0.58, 0.56, 0.57, 0.57, 0.59, 0.59, 0.55, 
    0.6, 0.56, 0.57, 0.6, 0.63, 0.64, 0.7, 0.73, 0.73, 0.73, 0.69, 0.7, 0.72, 
    0.7, 0.67, 0.63, 0.62, 0.63, 0.61, 0.57, 0.57, 0.52, 0.52, 0.6, 0.66, 
    0.56, 0.62, 0.56, 0.6, 0.57, 0.57, 0.59, 0.64, 0.63, 0.68, 0.63, 0.59, 
    0.6, 0.69, 0.67, 0.7, 0.68, 0.68, 0.66, 0.66, 0.63, 0.67, 0.68, 0.72, 
    0.71, 0.7, 0.76, 0.76, 0.79, 0.74, 0.73, 0.7, 0.71, 0.75, 0.74, 0.75, 
    0.72, 0.7, 0.7, 0.71, 0.69, 0.68, 0.68, 0.66, 0.68, 0.7, 0.72, 0.7, 0.69, 
    0.73, 0.77, 0.79, 0.79, 0.77, 0.78, 0.73, 0.66, 0.67, 0.64, 0.63, 0.63, 
    0.62, 0.58, 0.63, 0.62, 0.62, 0.6, 0.6, 0.59, 0.59, 0.59, 0.58, 0.56, 
    0.58, 0.59, 0.58, 0.62, 0.65, 0.66, 0.66, 0.65, 0.63, 0.62, 0.62, 0.63, 
    0.61, 0.65, 0.65, 0.63, 0.62, 0.6, 0.58, 0.54, 0.58, 0.56, 0.57, 0.55, 
    0.53, 0.54, 0.64, 0.65, 0.64, 0.68, 0.69, 0.77, 0.72, 0.75, 0.8, 0.78, 
    0.78, 0.75, 0.74, 0.72, 0.69, 0.7, 0.62, 0.67, 0.64, 0.66, 0.58, 0.6, 
    0.61, 0.58, 0.62, 0.67, 0.64, 0.68, 0.7, 0.73, 0.72, 0.61, 0.69, 0.7, 
    0.66, 0.7, 0.69, 0.68, 0.65, 0.65, 0.64, 0.55, 0.57, 0.55, 0.56, 0.5, 
    0.56, 0.52, 0.55, 0.52, 0.54, 0.57, 0.6, 0.56, 0.61, 0.53, 0.58, 0.58, 
    0.55, 0.66, 0.59, 0.64, 0.62, 0.6, 0.57, 0.57, 0.58, 0.58, 0.56, 0.56, 
    0.55, 0.5, 0.57, 0.56, 0.5, 0.52, 0.46, 0.49, 0.5, 0.52, 0.56, 0.55, 
    0.55, 0.59, 0.56, 0.6, 0.66, 0.64, 0.67, 0.66, 0.69, 0.69, 0.64, 0.61, 
    0.61, 0.6, 0.58, 0.57, 0.59, 0.57, 0.55, 0.57, 0.59, 0.59, 0.62, 0.56, 
    0.49, 0.47, 0.45, 0.47, 0.47, 0.4, 0.41, 0.4, 0.39, 0.41, 0.44, 0.46, 
    0.47, 0.48, 0.5, 0.53, 0.53, 0.56, 0.6, 0.63, 0.62, 0.63, 0.63, 0.62, 
    0.62, 0.62, 0.61, 0.61, 0.65, 0.68, 0.68, 0.64, 0.64, 0.65, 0.59, 0.54, 
    0.59, 0.62, 0.63, 0.69, 0.73, 0.8, 0.79, 0.75, 0.74, 0.81, 0.9, 0.95, 
    0.92, 0.92, 0.93, 0.89, 0.87, 0.88, 0.86, 0.86, 0.87, 0.88, 0.89, 0.95, 
    0.96, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.96, 0.96, 0.94, 0.92, 0.88, 0.82, 0.9, 0.9, 0.92, 0.95, 
    0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.99, 0.99, 0.98, 0.98, 
    0.98, 0.98, 0.96, 0.95, 0.93, 0.93, 0.91, 0.87, 0.86, 0.86, 0.88, 0.89, 
    0.88, 0.9, 0.9, 0.84, 0.82, 0.8, 0.79, 0.78, 0.77, 0.78, 0.76, 0.73, 
    0.68, 0.66, 0.62, 0.59, 0.57, 0.58, 0.59, 0.58, 0.56, 0.55, 0.56, 0.56, 
    0.59, 0.6, 0.66, 0.72, 0.73, 0.74, 0.74, 0.74, 0.75, 0.72, 0.73, 0.73, 
    0.7, 0.7, 0.69, 0.64, 0.6, 0.6, 0.64, 0.7, 0.52, 0.6, 0.66, 0.65, 0.68, 
    0.69, 0.6, 0.62, 0.69, 0.7, 0.66, 0.76, 0.77, 0.7, 0.63, 0.63, 0.67, 
    0.57, 0.54, 0.61, 0.65, 0.73, 0.75, 0.69, 0.66, 0.63, 0.63, 0.61, 0.66, 
    0.72, 0.75, 0.8, 0.73, 0.71, 0.69, 0.66, 0.68, 0.66, 0.67, 0.69, 0.66, 
    0.6, 0.6, 0.58, 0.61, 0.52, 0.6, 0.61, 0.62, 0.62, 0.63, 0.65, 0.67, 
    0.68, 0.67, 0.66, 0.65, 0.68, 0.7, 0.73, 0.7, 0.68, 0.61, 0.65, 0.64, 
    0.56, 0.51, 0.52, 0.54, 0.58, 0.63, 0.59, 0.62, 0.64, 0.65, 0.63, 0.64, 
    0.62, 0.6, 0.59, 0.61, 0.59, 0.61, 0.64, 0.65, 0.71, 0.74, 0.66, 0.63, 
    0.63, 0.64, 0.68, 0.64, 0.67, 0.65, 0.66, 0.59, 0.58, 0.61, 0.61, 0.61, 
    0.61, 0.61, 0.56, 0.67, 0.59, 0.68, 0.75, 0.69, 0.76, 0.7, 0.73, 0.62, 
    0.61, 0.55, 0.61, 0.59, 0.63, 0.64, 0.6, 0.56, 0.58, 0.6, 0.61, 0.59, 
    0.6, 0.66, 0.73, 0.71, 0.7, 0.76, 0.73, 0.69, 0.82, 0.78, 0.73, 0.66, 
    0.69, 0.56, 0.56, 0.56, 0.55, 0.53, 0.53, 0.53, 0.52, 0.54, 0.54, 0.55, 
    0.57, 0.55, 0.58, 0.57, 0.62, 0.65, 0.68, 0.68, 0.69, 0.68, 0.67, 0.69, 
    0.7, 0.69, 0.68, 0.73, 0.68, 0.69, 0.7, 0.7, 0.7, 0.7, 0.68, 0.58, 0.71, 
    0.68, 0.62, 0.63, 0.6, 0.54, 0.58, 0.56, 0.56, 0.53, 0.52, 0.53, 0.55, 
    0.58, 0.57, 0.64, 0.67, 0.67, 0.63, 0.59, 0.61, 0.61, 0.63, 0.64, 0.62, 
    0.64, 0.64, 0.64, 0.64, 0.65, 0.67, 0.66, 0.69, 0.68, 0.68, 0.73, 0.73, 
    0.71, 0.71, 0.7, 0.7, 0.73, 0.76, 0.76, 0.78, 0.8, 0.77, 0.78, 0.8, 0.77, 
    0.83, 0.87, 0.82, 0.86, 0.91, 0.9, 0.91, 0.88, 0.87, 0.87, 0.91, 0.88, 
    0.89, 0.88, 0.83, 0.84, 0.85, 0.72, 0.67, 0.83, 0.67, 0.68, 0.68, 0.71, 
    0.76, 0.73, 0.71, 0.73, 0.82, 0.76, 0.75, 0.71, 0.79, 0.79, 0.74, 0.68, 
    0.68, 0.79, 0.74, 0.76, 0.75, 0.75, 0.79, 0.7, 0.73, 0.76, 0.75, 0.84, 
    0.79, 0.75, 0.69, 0.75, 0.74, 0.72, 0.73, 0.7, 0.68, 0.7, 0.66, 0.67, 
    0.65, 0.64, 0.63, 0.62, 0.66, 0.56, 0.57, 0.61, 0.61, 0.62, 0.64, 0.66, 
    0.69, 0.66, 0.67, 0.72, 0.72, 0.74, 0.68, 0.72, 0.74, 0.72, 0.7, 0.69, 
    0.66, 0.63, 0.65, 0.63, 0.65, 0.67, 0.69, 0.71, 0.69, 0.74, 0.73, 0.71, 
    0.75, 0.72, 0.75, 0.72, 0.75, 0.75, 0.75, 0.73, 0.75, 0.73, 0.7, 0.66, 
    0.69, 0.7, 0.65, 0.69, 0.68, 0.66, 0.62, 0.73, 0.78, 0.79, 0.73, 0.74, 
    0.77, 0.82, 0.78, 0.81, 0.81, 0.78, 0.83, 0.84, 0.87, 0.79, 0.65, 0.64, 
    0.68, 0.58, 0.49, 0.64, 0.56, 0.48, 0.36, 0.37, 0.35, 0.34, 0.34, 0.36, 
    0.44, 0.51, 0.45, 0.51, 0.44, 0.52, 0.56, 0.5, 0.5, 0.46, 0.38, 0.37, 
    0.36, 0.38, 0.36, 0.3, 0.33, 0.33, 0.33, 0.33, 0.34, 0.43, 0.34, 0.37, 
    0.4, 0.36, 0.45, 0.41, 0.43, 0.45, 0.45, 0.44, 0.48, 0.43, 0.5, 0.51, 
    0.4, 0.41, 0.41, 0.44, 0.43, 0.41, 0.39, 0.37, 0.41, 0.42, 0.4, 0.45, 
    0.47, 0.51, 0.54, 0.56, 0.53, 0.54, 0.57, 0.58, 0.61, 0.61, 0.51, 0.44, 
    0.48, 0.42, 0.49, 0.41, 0.46, 0.43, 0.43, 0.46, 0.4, 0.44, 0.47, 0.39, 
    0.46, 0.46, 0.46, 0.5, 0.47, 0.59, 0.57, 0.63, 0.7, 0.59, 0.58, 0.6, 0.6, 
    0.54, 0.42, 0.65, 0.64, 0.59, 0.58, 0.61, 0.67, 0.84, 0.89, 0.87, 0.87, 
    0.88, 0.88, 0.85, 0.87, 0.88, 0.87, 0.86, 0.87, 0.84, 0.86, 0.85, 0.87, 
    0.88, 0.84, 0.82, 0.8, 0.79, 0.78, 0.8, 0.79, 0.78, 0.77, 0.77, 0.75, 
    0.75, 0.82, 0.84, 0.88, 0.87, 0.89, 0.86, 0.9, 0.91, 0.9, 0.84, 0.84, 
    0.87, 0.86, 0.81, 0.66, 0.71, 0.52, 0.51, 0.48, 0.49, 0.6, 0.73, 0.73, 
    0.72, 0.72, 0.74, 0.79, 0.8, 0.82, 0.81, 0.84, 0.82, 0.81, 0.81, 0.83, 
    0.85, 0.91, 0.9, 0.91, 0.91, 0.92, 0.93, 0.93, 0.92, 0.89, 0.85, 0.89, 
    0.88, 0.89, 0.91, 0.94, 0.95, 0.95, 0.95, 0.94, 0.92, 0.91, 0.9, 0.88, 
    0.92, 0.91, 0.86, 0.85, 0.85, 0.83, 0.89, 0.85, 0.84, 0.9, 0.89, 0.9, 
    0.91, 0.9, 0.89, 0.88, 0.87, 0.9, 0.91, 0.9, 0.89, 0.86, 0.85, 0.84, 
    0.82, 0.81, 0.81, 0.81, 0.82, 0.83, 0.85, 0.84, 0.83, 0.79, 0.75, 0.71, 
    0.69, 0.69, 0.7, 0.72, 0.72, 0.71, 0.74, 0.73, 0.73, 0.7, 0.72, 0.69, 
    0.67, 0.7, 0.73, 0.7, 0.66, 0.64, 0.64, 0.66, 0.76, 0.78, 0.72, 0.79, 
    0.78, 0.82, 0.84, 0.88, 0.9, 0.86, 0.86, 0.86, 0.85, 0.85, 0.84, 0.86, 
    0.82, 0.85, 0.84, 0.81, 0.83, 0.85, 0.85, 0.84, 0.86, 0.85, 0.84, 0.82, 
    0.85, 0.84, 0.86, 0.82, 0.85, 0.84, 0.81, 0.81, 0.73, 0.66, 0.68, 0.69, 
    0.67, 0.68, 0.67, 0.74, 0.72, 0.81, 0.85, 0.83, 0.82, 0.81, 0.82, 0.85, 
    0.87, 0.87, 0.87, 0.89, 0.87, 0.87, 0.87, 0.86, 0.89, 0.8, 0.75, 0.79, 
    0.77, 0.81, 0.78, 0.8, 0.69, 0.67, 0.66, 0.64, 0.64, 0.63, 0.64, 0.63, 
    0.65, 0.66, 0.66, 0.68, 0.68, 0.68, 0.68, 0.69, 0.67, 0.66, 0.64, 0.6, 
    0.61, 0.57, 0.55, 0.56, 0.56, 0.56, 0.57, 0.58, 0.62, 0.63, 0.68, 0.71, 
    0.73, 0.75, 0.8, 0.8, 0.81, 0.83, 0.76, 0.74, 0.68, 0.61, 0.58, 0.73, 
    0.86, 0.86, 0.86, 0.84, 0.86, 0.82, 0.84, 0.86, 0.86, 0.88, 0.88, 0.88, 
    0.91, 0.93, 0.94, 0.96, 0.92, 0.91, 0.9, 0.91, 0.89, 0.87, 0.82, 0.84, 
    0.85, 0.85, 0.84, 0.85, 0.84, 0.83, 0.83, 0.82, 0.85, 0.88, 0.89, 0.93, 
    0.92, 0.92, 0.92, 0.94, 0.94, 0.92, 0.9, 0.9, 0.87, 0.86, 0.87, 0.86, 
    0.86, 0.87, 0.86, 0.91, 0.88, 0.85, 0.86, 0.8, 0.78, 0.82, 0.84, 0.87, 
    0.84, 0.81, 0.86, 0.89, 0.91, 0.9, 0.89, 0.86, 0.85, 0.87, 0.87, 0.84, 
    0.86, 0.79, 0.83, 0.82, 0.85, 0.87, 0.84, 0.89, 0.92, 0.92, 0.94, 0.96, 
    0.93, 0.87, 0.74, 0.77, 0.76, 0.81, 0.89, 0.89, 0.83, 0.79, 0.84, 0.77, 
    0.77, 0.77, 0.73, 0.78, 0.81, 0.78, 0.79, 0.86, 0.88, 0.8, 0.8, 0.82, 
    0.78, 0.83, 0.84, 0.78, 0.75, 0.82, 0.8, 0.78, 0.79, 0.75, 0.75, 0.75, 
    0.78, 0.76, 0.77, 0.76, 0.73, 0.72, 0.74, 0.77, 0.79, 0.82, 0.81, 0.82, 
    0.84, 0.81, 0.8, 0.81, 0.79, 0.83, 0.76, 0.74, 0.71, 0.75, 0.74, 0.74, 
    0.72, 0.69, 0.67, 0.62, 0.68, 0.7, 0.71, 0.66, 0.67, 0.69, 0.75, 0.77, 
    0.75, 0.72, 0.71, 0.72, 0.72, 0.72, 0.75, 0.77, 0.78, 0.72, 0.71, 0.67, 
    0.68, 0.66, 0.67, 0.64, 0.72, 0.66, 0.7, 0.72, 0.67, 0.68, 0.7, 0.72, 
    0.72, 0.74, 0.76, 0.76, 0.76, 0.76, 0.75, 0.74, 0.73, 0.72, 0.64, 0.62, 
    0.53, 0.53, 0.55, 0.58, 0.62, 0.65, 0.66, 0.63, 0.64, 0.63, 0.64, 0.75, 
    0.75, 0.76, 0.75, 0.82, 0.79, 0.77, 0.74, 0.74, 0.74, 0.76, 0.75, 0.73, 
    0.77, 0.77, 0.73, 0.76, 0.8, 0.83, 0.84, 0.86, 0.89, 0.86, 0.87, 0.93, 
    0.96, 0.97, 0.97, 0.97, 0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.97, 0.97, 0.98, 0.98, 0.97, 0.98, 0.96, 0.89, 0.83, 0.83, 
    0.83, 0.86, 0.91, 0.92, 0.93, 0.96, 0.96, 0.97, 0.97, 0.96, 0.94, 0.9, 
    0.89, 0.88, 0.89, 0.84, 0.85, 0.86, 0.86, 0.82, 0.87, 0.88, 0.8, 0.79, 
    0.81, 0.85, 0.83, 0.84, 0.85, 0.81, 0.82, 0.82, 0.77, 0.73, 0.71, 0.74, 
    0.75, 0.68, 0.71, 0.73, 0.78, 0.82, 0.86, 0.85, 0.85, 0.84, 0.81, 0.85, 
    0.87, 0.91, 0.81, 0.73, 0.76, 0.75, 0.75, 0.74, 0.73, 0.72, 0.71, 0.7, 
    0.68, 0.72, 0.72, 0.72, 0.78, 0.8, 0.8, 0.72, 0.76, 0.77, 0.76, 0.75, 
    0.82, 0.82, 0.84, 0.84, 0.89, 0.88, 0.89, 1, 0.85, 0.69, 0.7, 0.66, 0.69, 
    0.67, 0.67, 0.65, 0.64, 0.63, 0.61, 0.6, 0.6, 0.62, 0.64, 0.65, 0.64, 
    0.66, 0.67, 0.75, 0.74, 0.78, 0.73, 0.76, 0.95, 0.95, 0.96, 0.95, 0.95, 
    0.95, 0.93, 0.86, 0.76, 0.7, 0.63, 0.66, 0.62, 0.61, 0.62, 0.65, 0.57, 
    0.59, 0.58, 0.6, 0.62, 0.63, 0.61, 0.6, 0.61, 0.63, 0.61, 0.62, 0.64, 
    0.6, 0.6, 0.59, 0.61, 0.6, 0.6, 0.62, 0.65, 0.69, 0.7, 0.77, 0.72, 0.73, 
    0.7, 0.64, 0.66, 0.75, 0.7, 0.65, 0.65, 0.72, 0.6, 0.62, 0.72, 0.75, 
    0.74, 0.76, 0.72, 0.66, 0.62, 0.6, 0.62, 0.63, 0.64, 0.61, 0.63, 0.64, 
    0.6, 0.62, 0.6, 0.59, 0.59, 0.58, 0.58, 0.59, 0.6, 0.61, 0.51, 0.59, 
    0.59, 0.58, 0.56, 0.55, 0.54, 0.56, 0.61, 0.61, 0.55, 0.56, 0.57, 0.57, 
    0.53, 0.55, 0.6, 0.62, 0.62, 0.55, 0.53, 0.52, 0.55, 0.58, 0.6, 0.61, 
    0.62, 0.61, 0.66, 0.63, 0.65, 0.62, 0.61, 0.62, 0.6, 0.6, 0.6, 0.6, 0.66, 
    0.64, 0.62, 0.62, 0.65, 0.61, 0.58, 0.63, 0.62, 0.59, 0.56, 0.57, 0.56, 
    0.6, 0.6, 0.58, 0.58, 0.61, 0.64, 0.62, 0.6, 0.55, 0.55, 0.62, 0.61, 
    0.62, 0.62, 0.64, 0.63, 0.65, 0.68, 0.73, 0.72, 0.69, 0.66, 0.62, 0.62, 
    0.62, 0.61, 0.56, 0.6, 0.59, 0.59, 0.61, 0.62, 0.64, 0.62, 0.6, 0.62, 
    0.64, 0.67, 0.63, 0.67, 0.7, 0.71, 0.69, 0.69, 0.69, 0.66, 0.66, 0.67, 
    0.74, 0.74, 0.75, 0.76, 0.77, 0.79, 0.82, 0.84, 0.85, 0.86, 0.88, 0.89, 
    0.86, 0.85, 0.87, 0.88, 0.87, 0.89, 0.87, 0.84, 0.81, 0.81, 0.8, 0.79, 
    0.78, 0.76, 0.76, 0.77, 0.72, 0.81, 0.83, 0.82, 0.8, 0.82, 0.78, 0.79, 
    0.79, 0.79, 0.78, 0.82, 0.83, 0.81, 0.77, 0.74, 0.69, 0.75, 0.82, 0.8, 
    0.75, 0.73, 0.83, 0.82, 0.8, 0.76, 0.75, 0.73, 0.65, 0.66, 0.74, 0.76, 
    0.76, 0.75, 0.73, 0.74, 0.69, 0.7, 0.71, 0.7, 0.69, 0.68, 0.67, 0.67, 
    0.66, 0.67, 0.65, 0.66, 0.66, 0.7, 0.7, 0.74, 0.68, 0.65, 0.6, 0.55, 
    0.53, 0.54, 0.56, 0.54, 0.54, 0.57, 0.51, 0.52, 0.52, 0.52, 0.5, 0.49, 
    0.5, 0.49, 0.53, 0.57, 0.57, 0.58, 0.66, 0.68, 0.69, 0.66, 0.72, 0.72, 
    0.74, 0.69, 0.74, 0.65, 0.66, 0.67, 0.66, 0.64, 0.67, 0.75, 0.83, 0.85, 
    0.86, 0.87, 0.88, 0.89, 0.8, 0.79, 0.74, 0.68, 0.65, 0.69, 0.64, 0.69, 
    0.76, 0.92, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 0.96, 0.96, 0.95, 0.95, 
    0.96, 0.98, 0.9, 0.88, 0.87, 0.87, 0.87, 0.88, 0.88, 0.83, 0.82, 0.8, 
    0.81, 0.8, 0.75, 0.74, 0.75, 0.74, 0.76, 0.74, 0.72, 0.71, 0.71, 0.79, 
    0.91, 0.95, 0.95, 0.95, 0.95, 0.95, 0.96, 0.97, 0.97, 0.98, 0.97, 0.98, 
    0.92, 0.91, 0.9, 0.88, 0.88, 0.87, 0.86, 0.87, 0.88, 0.89, 0.9, 0.88, 
    0.81, 0.83, 0.81, 0.81, 0.8, 0.79, 0.8, 0.83, 0.86, 0.92, 0.94, 0.93, 
    0.9, 0.89, 0.93, 0.94, 0.93, 0.95, 0.93, 0.93, 0.94, 0.96, 0.96, 0.95, 
    0.95, 0.96, 0.95, 0.97, 0.97, 0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.97, 
    0.98, 0.9, 0.89, 0.89, 0.85, 0.84, 0.78, 0.75, 0.73, 0.74, 0.73, 0.66, 
    0.68, 0.71, 0.7, 0.71, 0.76, 0.72, 0.72, 0.76, 0.81, 0.81, 0.81, 0.84, 
    0.8, 0.87, 0.87, 0.89, 0.87, 0.83, 0.79, 0.82, 0.8, 0.83, 0.81, 0.79, 
    0.8, 0.82, 0.83, 0.83, 0.83, 0.84, 0.83, 0.82, 0.87, 0.85, 0.82, 0.85, 
    0.79, 0.8, 0.77, 0.81, 0.76, 0.82, 0.83, 0.84, 0.85, 0.86, 0.85, 0.78, 
    0.73, 0.69, 0.71, 0.8, 0.79, 0.78, 0.81, 0.82, 0.8, 0.81, 0.81, 0.83, 
    0.85, 0.86, 0.88, 0.88, 0.89, 0.9, 0.91, 0.92, 0.94, 0.94, 0.95, 0.96, 
    0.96, 0.97, 0.96, 0.93, 0.94, 0.92, 0.87, 0.88, 0.88, 0.87, 0.8, 0.78, 
    0.8, 0.77, 0.71, 0.79, 0.79, 0.77, 0.73, 0.73, 0.67, 0.66, 0.7, 0.68, 
    0.7, 0.73, 0.74, 0.69, 0.71, 0.78, 0.8, 0.83, 0.82, 0.84, 0.83, 0.83, 
    0.86, 0.87, 0.86, 0.87, 0.88, 0.88, 0.86, 0.87, 0.83, 0.84, 0.89, 0.88, 
    0.85, 0.91, 0.94, 0.93, 0.83, 0.75, 0.76, 0.76, 0.74, 0.75, 0.75, 0.71, 
    0.69, 0.68, 0.77, 0.68, 0.77, 0.71, 0.77, 0.76, 0.74, 0.76, 0.88, 0.91, 
    0.91, 0.94, 0.95, 0.94, 0.94, 0.95, 0.96, 0.97, 0.97, 0.97, 0.98, 0.97, 
    0.97, 0.96, 0.95, 0.96, 0.96, 0.95, 0.95, 0.93, 0.94, 0.94, 0.93, 0.93, 
    0.93, 0.94, 0.96, 0.93, 0.9, 0.92, 0.9, 0.9, 0.91, 0.91, 0.92, 0.93, 
    0.89, 0.9, 0.91, 0.91, 0.92, 0.9, 0.89, 0.9, 0.86, 0.87, 0.9, 0.91, 0.91, 
    0.88, 0.9, 0.9, 0.85, 0.79, 0.78, 0.79, 0.77, 0.79, 0.75, 0.75, 0.75, 
    0.75, 0.77, 0.76, 0.79, 0.79, 0.79, 0.79, 0.81, 0.84, 0.79, 0.77, 0.77, 
    0.81, 0.83, 0.81, 0.85, 0.89, 0.86, 0.86, 0.9, 0.88, 0.9, 0.88, 0.9, 
    0.87, 0.89, 0.91, 0.91, 0.9, 0.89, 0.88, 0.87, 0.86, 0.88, 0.87, 0.87, 
    0.86, 0.84, 0.8, 0.85, 0.82, 0.84, 0.86, 0.9, 0.91, 0.88, 0.87, 0.87, 
    0.85, 0.88, 0.83, 0.83, 0.84, 0.8, 0.8, 0.79, 0.77, 0.76, 0.76, 0.77, 
    0.79, 0.79, 0.82, 0.84, 0.88, 0.85, 0.85, 0.85, 0.88, 0.85, 0.88, 0.87, 
    0.89, 0.89, 0.92, 0.91, 0.93, 0.95, 0.96, 0.96, 0.96, 0.95, 0.94, 0.95, 
    0.95, 0.95, 0.95, 0.94, 0.94, 0.94, 0.94, 0.95, 0.96, 0.97, 0.97, 0.97, 
    0.96, 0.95, 0.94, 0.91, 0.89, 0.93, 0.95, 0.93, 0.93, 0.94, 0.91, 0.89, 
    0.9, 0.92, 0.89, 0.91, 0.92, 0.9, 0.94, 0.96, 0.97, 0.96, 0.94, 0.94, 
    0.88, 0.93, 0.95, 0.7, 0.82, 0.75, 0.86, 0.81, 0.84, 0.85, 0.79, 0.65, 
    0.69, 0.75, 0.64, 0.63, 0.73, 0.74, 0.71, 0.69, 0.71, 0.69, 0.65, 0.7, 
    0.65, 0.65, 0.78, 0.75, 0.65, 0.61, 0.58, 0.56, 0.53, 0.49, 0.58, 0.61, 
    0.62, 0.6, 0.61, 0.61, 0.61, 0.61, 0.61, 0.58, 0.56, 0.59, 0.53, 0.53, 
    0.52, 0.55, 0.56, 0.54, 0.51, 0.52, 0.49, 0.47, 0.53, 0.52, 0.54, 0.55, 
    0.56, 0.57, 0.57, 0.61, 0.6, 0.6, 0.63, 0.7, 0.68, 0.61, 0.6, 0.56, 0.63, 
    0.67, 0.6, 0.66, 0.63, 0.64, 0.62, 0.6, 0.61, 0.64, 0.64, 0.62, 0.59, 
    0.66, 0.67, 0.65, 0.66, 0.68, 0.69, 0.7, 0.69, 0.72, 0.72, 0.71, 0.71, 
    0.69, 0.71, 0.65, 0.7, 0.73, 0.71, 0.68, 0.66, 0.64, 0.61, 0.51, 0.53, 
    0.58, 0.56, 0.6, 0.6, 0.57, 0.6, 0.53, 0.6, 0.54, 0.64, 0.58, 0.55, 0.6, 
    0.58, 0.5, 0.51, 0.48, 0.54, 0.54, 0.47, 0.48, 0.52, 0.64, 0.61, 0.58, 
    0.63, 0.65, 0.67, 0.64, 0.64, 0.68, 0.67, 0.65, 0.66, 0.66, 0.66, 0.68, 
    0.64, 0.69, 0.67, 0.71, 0.63, 0.69, 0.67, 0.65, 0.68, 0.64, 0.69, 0.69, 
    0.71, 0.75, 0.75, 0.73, 0.75, 0.74, 0.76, 0.75, 0.75, 0.76, 0.75, 0.78, 
    0.77, 0.77, 0.76, 0.78, 0.79, 0.8, 0.8, 0.77, 0.81, 0.91, 0.93, 0.95, 
    0.95, 0.95, 0.92, 0.89, 0.88, 0.86, 0.88, 0.85, 0.85, 0.83, 0.87, 0.87, 
    0.92, 0.91, 0.93, 0.94, 0.92, 0.92, 0.91, 0.91, 0.91, 0.9, 0.91, 0.93, 
    0.94, 0.91, 0.93, 0.92, 0.91, 0.89, 0.94, 0.93, 0.94, 0.94, 0.94, 0.92, 
    0.94, 0.94, 0.94, 0.91, 0.91, 0.91, 0.9, 0.9, 0.89, 0.9, 0.92, 0.85, 
    0.85, 0.84, 0.85, 0.87, 0.87, 0.9, 0.83, 0.86, 0.86, 0.88, 0.85, 0.88, 
    0.9, 0.77, 0.81, 0.82, 0.8, 0.76, 0.76, 0.84, 0.89, 0.87, 0.87, 0.73, 
    0.81, 0.82, 0.77, 0.85, 0.85, 0.84, 0.86, 0.85, 0.87, 0.88, 0.87, 0.85, 
    0.86, 0.89, 0.92, 0.94, 0.92, 0.91, 0.92, 0.92, 0.92, 0.95, 0.95, 0.94, 
    0.93, 0.93, 0.95, 0.92, 0.9, 0.95, 0.93, 0.94, 0.91, 0.85, 0.78, 0.91, 
    0.88, 0.88, 0.92, 0.9, 0.89, 0.93, 0.9, 0.87, 0.82, 0.85, 0.81, 0.78, 
    0.84, 0.77, 0.72, 0.72, 0.77, 0.81, 0.82, 0.77, 0.82, 0.83, 0.85, 0.85, 
    0.87, 0.86, 0.92, 0.91, 0.92, 0.94, 0.95, 0.96, 0.96, 0.96, 0.95, 0.96, 
    0.96, 0.92, 0.93, 0.95, 0.96, 0.97, 0.97, 0.97, 0.97, 0.97, 0.93, 0.89, 
    0.92, 0.92, 0.92, 0.89, 0.94, 0.95, 0.96, 0.97, 0.95, 0.96, 0.95, 0.86, 
    0.83, 0.83, 0.81, 0.87, 0.84, 0.78, 0.84, 0.85, 0.83, 0.86, 0.88, 0.87, 
    0.86, 0.86, 0.88, 0.79, 0.74, 0.71, 0.67, 0.65, 0.67, 0.64, 0.66, 0.71, 
    0.95, 0.95, 0.92, 0.88, 0.81, 0.84, 0.89, 0.87, 0.77, 0.81, 0.77, 0.77, 
    0.82, 0.79, 0.88, 0.84, 0.84, 0.84, 0.84, 0.83, 0.86, 0.85, 0.91, 0.95, 
    0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.91, 0.78, 0.82, 0.87, 0.87, 
    0.86, 0.93, 0.93, 0.9, 0.9, 0.92, 0.84, 0.83, 0.82, 0.78, 0.8, 0.79, 
    0.78, 0.75, 0.73, 0.76, 0.76, 0.77, 0.75, 0.76, 0.74, 0.73, 0.73, 0.72, 
    0.78, 0.79, 0.82, 0.78, 0.79, 0.7, 0.67, 0.67, 0.68, 0.7, 0.73, 0.71, 
    0.72, 0.7, 0.68, 0.71, 0.72, 0.74, 0.75, 0.74, 0.75, 0.73, 0.77, 0.7, 
    0.78, 0.77, 0.76, 0.77, 0.8, 0.83, 0.87, 0.92, 0.93, 0.93, 0.94, 0.93, 
    0.95, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.97, 0.96, 0.95, 0.97, 0.96, 
    0.97, 0.97, 0.91, 0.87, 0.93, 0.92, 0.85, 0.79, 0.78, 0.76, 0.72, 0.72, 
    0.82, 0.82, 0.79, 0.75, 0.67, 0.74, 0.71, 0.66, 0.64, 0.66, 0.71, 0.66, 
    0.66, 0.65, 0.62, 0.59, 0.54, 0.55, 0.55, 0.56, 0.54, 0.59, 0.61, 0.62, 
    0.63, 0.6, 0.63, 0.62, 0.57, 0.56, 0.56, 0.55, 0.56, 0.55, 0.57, 0.54, 
    0.54, 0.54, 0.6, 0.62, 0.58, 0.58, 0.59, 0.63, 0.57, 0.58, 0.63, 0.61, 
    0.59, 0.53, 0.54, 0.53, 0.56, 0.56, 0.54, 0.53, 0.54, 0.58, 0.61, 0.63, 
    0.61, 0.59, 0.6, 0.62, 0.65, 0.63, 0.65, 0.6, 0.65, 0.61, 0.65, 0.65, 
    0.62, 0.62, 0.64, 0.64, 0.65, 0.63, 0.6, 0.63, 0.6, 0.61, 0.64, 0.61, 
    0.6, 0.6, 0.61, 0.63, 0.63, 0.62, 0.63, 0.57, 0.61, 0.6, 0.67, 0.63, 0.6, 
    0.6, 0.6, 0.59, 0.64, 0.78, 0.65, 0.62, 0.61, 0.6, 0.55, 0.53, 0.6, 0.57, 
    0.54, 0.63, 0.68, 0.72, 0.75, 0.73, 0.68, 0.64, 0.6, 0.55, 0.56, 0.56, 
    0.58, 0.57, 0.63, 0.55, 0.6, 0.63, 0.57, 0.55, 0.57, 0.61, 0.57, 0.58, 
    0.57, 0.56, 0.61, 0.6, 0.62, 0.63, 0.62, 0.66, 0.62, 0.66, 0.66, 0.64, 
    0.63, 0.57, 0.49, 0.48, 0.51, 0.5, 0.49, 0.59, 0.56, 0.57, 0.56, 0.53, 
    0.54, 0.53, 0.55, 0.58, 0.55, 0.49, 0.5, 0.51, 0.52, 0.55, 0.58, 0.59, 
    0.63, 0.6, 0.6, 0.62, 0.6, 0.67, 0.63, 0.61, 0.65, 0.67, 0.67, 0.7, 0.69, 
    0.7, 0.72, 0.73, 0.73, 0.71, 0.7, 0.7, 0.69, 0.74, 0.71, 0.68, 0.68, 
    0.67, 0.67, 0.63, 0.62, 0.67, 0.64, 0.6, 0.6, 0.64, 0.63, 0.64, 0.62, 
    0.64, 0.59, 0.57, 0.52, 0.55, 0.55, 0.53, 0.52, 0.54, 0.59, 0.57, 0.58, 
    0.57, 0.57, 0.58, 0.59, 0.64, 0.68, 0.71, 0.72, 0.78, 0.8, 0.8, 0.74, 
    0.75, 0.75, 0.75, 0.72, 0.72, 0.75, 0.84, 0.83, 0.88, 0.89, 0.91, 0.89, 
    0.88, 0.88, 0.92, 0.92, 0.93, 0.93, 0.94, 0.94, 0.94, 0.94, 0.94, 0.95, 
    0.95, 0.96, 0.95, 0.88, 0.84, 0.84, 0.85, 0.83, 0.83, 0.84, 0.86, 0.86, 
    0.89, 0.83, 0.87, 0.86, 0.83, 0.86, 0.88, 0.92, 0.9, 0.87, 0.88, 0.91, 
    0.91, 0.88, 0.88, 0.88, 0.89, 0.88, 0.83, 0.81, 0.85, 0.85, 0.89, 0.87, 
    0.86, 0.9, 0.93, 0.94, 0.9, 0.94, 0.97, 0.97, 0.89, 0.85, 0.9, 0.89, 
    0.82, 0.83, 0.84, 0.87, 0.87, 0.89, 0.94, 0.94, 0.93, 0.9, 0.9, 0.91, 
    0.85, 0.88, 0.89, 0.91, 0.9, 0.89, 0.82, 0.9, 0.87, 0.89, 0.85, 0.87, 
    0.81, 0.84, 0.83, 0.89, 0.88, 0.86, 0.89, 0.9, 0.75, 0.71, 0.72, 0.68, 
    0.69, 0.67, 0.67, 0.69, 0.69, 0.7, 0.7, 0.69, 0.66, 0.68, 0.68, 0.69, 
    0.71, 0.7, 0.69, 0.72, 0.71, 0.71, 0.71, 0.7, 0.69, 0.69, 0.68, 0.72, 
    0.7, 0.68, 0.75, 0.75, 0.84, 0.81, 0.75, 0.75, 0.68, 0.6, 0.64, 0.73, 
    0.77, 0.8, 0.8, 0.79, 0.73, 0.7, 0.78, 0.83, 0.81, 0.63, 0.59, 0.58, 
    0.59, 0.55, 0.58, 0.62, 0.6, 0.66, 0.77, 0.77, 0.78, 0.8, 0.82, 0.72, 
    0.65, 0.66, 0.6, 0.59, 0.58, 0.59, 0.52, 0.5, 0.48, 0.5, 0.51, 0.55, 
    0.56, 0.55, 0.6, 0.61, 0.61, 0.62, 0.6, 0.61, 0.65, 0.66, 0.66, 0.67, 
    0.7, 0.74, 0.71, 0.73, 0.75, 0.77, 0.79, 0.78, 0.75, 0.81, 0.78, 0.77, 
    0.79, 0.78, 0.81, 0.77, 0.86, 0.79, 0.78, 0.77, 0.76, 0.77, 0.78, 0.79, 
    0.79, 0.79, 0.82, 0.82, 0.83, 0.82, 0.81, 0.81, 0.8, 0.78, 0.79, 0.76, 
    0.77, 0.74, 0.75, 0.71, 0.71, 0.75, 0.74, 0.72, 0.68, 0.65, 0.7, 0.7, 
    0.65, 0.66, 0.68, 0.68, 0.69, 0.72, 0.72, 0.81, 0.87, 0.88, 0.85, 0.85, 
    0.85, 0.88, 0.87, 0.91, 0.87, 0.89, 0.92, 0.81, 0.91, 0.91, 0.82, 0.77, 
    0.71, 0.74, 0.74, 0.72, 0.8, 0.82, 0.82, 0.83, 0.83, 0.8, 0.79, 0.81, 
    0.76, 0.77, 0.85, 0.78, 0.7, 0.74, 0.72, 0.66, 0.65, 0.65, 0.67, 0.68, 
    0.68, 0.68, 0.73, 0.69, 0.71, 0.69, 0.69, 0.67, 0.68, 0.64, 0.64, 0.66, 
    0.64, 0.67, 0.65, 0.67, 0.68, 0.68, 0.67, 0.68, 0.66, 0.64, 0.66, 0.68, 
    0.71, 0.72, 0.71, 0.71, 0.72, 0.67, 0.71, 0.71, 0.72, 0.71, 0.71, 0.73, 
    0.73, 0.69, 0.62, 0.61, 0.65, 0.86, 0.85, 0.67, 0.66, 0.63, 0.6, 0.61, 
    0.64, 0.62, 0.59, 0.6, 0.57, 0.61, 0.64, 0.63, 0.7, 0.65, 0.66, 0.68, 
    0.7, 0.66, 0.69, 0.63, 0.64, 0.66, 0.67, 0.65, 0.62, 0.57, 0.73, 0.71, 
    0.63, 0.74, 0.75, 0.76, 0.78, 0.62, 0.65, 0.67, 0.71, 0.58, 0.72, 0.73, 
    0.69, 0.66, 0.7, 0.73, 0.7, 0.65, 0.62, 0.6, 0.61, 0.65, 0.66, 0.59, 
    0.59, 0.75, 0.66, 0.63, 0.62, 0.69, 0.59, 0.62, 0.56, 0.58, 0.52, 0.6, 
    0.68, 0.76, 0.58, 0.56, 0.54, 0.53, 0.5, 0.54, 0.6, 0.61, 0.6, 0.62, 
    0.65, 0.64, 0.61, 0.6, 0.6, 0.62, 0.61, 0.61, 0.65, 0.72, 0.61, 0.57, 
    0.57, 0.59, 0.59, 0.59, 0.67, 0.59, 0.64, 0.63, 0.66, 0.62, 0.7, 0.83, 
    0.93, 0.74, 0.65, 0.6, 0.6, 0.59, 0.56, 0.65, 0.68, 0.66, 0.64, 0.69, 
    0.67, 0.7, 0.74, 0.76, 0.75, 0.78, 0.74, 0.76, 0.76, 0.77, 0.77, 0.78, 
    0.8, 0.8, 0.78, 0.78, 0.79, 0.81, 0.8, 0.79, 0.78, 0.76, 0.69, 0.69, 
    0.64, 0.66, 0.68, 0.64, 0.6, 0.6, 0.61, 0.56, 0.59, 0.58, 0.62, 0.63, 
    0.61, 0.6, 0.6, 0.64, 0.64, 0.66, 0.64, 0.62, 0.65, 0.65, 0.69, 0.65, 
    0.64, 0.63, 0.64, 0.64, 0.64, 0.64, 0.65, 0.64, 0.64, 0.64, 0.64, 0.64, 
    0.66, 0.63, 0.65, 0.68, 0.68, 0.67, 0.69, 0.67, 0.68, 0.69, 0.68, 0.66, 
    0.64, 0.68, 0.7, 0.67, 0.7, 0.72, 0.67, 0.65, 0.67, 0.69, 0.68, 0.72, 
    0.79, 0.78, 0.77, 0.71, 0.69, 0.69, 0.69, 0.7, 0.66, 0.62, 0.6, 0.57, 
    0.54, 0.59, 0.58, 0.58, 0.58, 0.56, 0.57, 0.57, 0.59, 0.59, 0.59, 0.58, 
    0.58, 0.61, 0.64, 0.66, 0.69, 0.7, 0.72, 0.7, 0.71, 0.71, 0.75, 0.71, 
    0.73, 0.7, 0.72, 0.71, 0.75, 0.76, 0.78, 0.75, 0.77, 0.76, 0.74, 0.72, 
    0.72, 0.76, 0.83, 0.9, 0.9, 0.78, 0.64, 0.64, 0.6, 0.55, 0.52, 0.58, 
    0.53, 0.55, 0.52, 0.63, 0.63, 0.57, 0.64, 0.58, 0.61, 0.67, 0.68, 0.64, 
    0.61, 0.57, 0.57, 0.65, 0.7, 0.57, 0.57, 0.55, 0.57, 0.61, 0.65, 0.64, 
    0.61, 0.62, 0.61, 0.63, 0.64, 0.64, 0.63, 0.65, 0.64, 0.64, 0.68, 0.63, 
    0.65, 0.67, 0.69, 0.67, 0.64, 0.6, 0.58, 0.59, 0.61, 0.61, 0.61, 0.62, 
    0.59, 0.62, 0.64, 0.66, 0.66, 0.69, 0.64, 0.66, 0.65, 0.64, 0.64, 0.66, 
    0.64, 0.65, 0.65, 0.68, 0.65, 0.66, 0.61, 0.61, 0.61, 0.61, 0.61, 0.63, 
    0.61, 0.61, 0.6, 0.64, 0.65, 0.64, 0.64, 0.65, 0.66, 0.66, 0.68, 0.69, 
    0.63, 0.6, 0.59, 0.61, 0.61, 0.64, 0.67, 0.7, 0.7, 0.71, 0.64, 0.62, 
    0.65, 0.6, 0.62, 0.61, 0.53, 0.51, 0.52, 0.56, 0.55, 0.56, 0.73, 0.6, 
    0.54, 0.52, 0.54, 0.57, 0.58, 0.63, 0.63, 0.63, 0.74, 0.73, 0.62, 0.56, 
    0.55, 0.53, 0.58, 0.48, 0.55, 0.51, 0.57, 0.54, 0.52, 0.53, 0.53, 0.51, 
    0.5, 0.53, 0.54, 0.54, 0.52, 0.53, 0.57, 0.58, 0.57, 0.58, 0.54, 0.59, 
    0.58, 0.57, 0.58, 0.54, 0.56, 0.5, 0.54, 0.53, 0.54, 0.64, 0.55, 0.56, 
    0.54, 0.47, 0.5, 0.53, 0.44, 0.47, 0.49, 0.47, 0.47, 0.5, 0.47, 0.44, 
    0.44, 0.43, 0.44, 0.46, 0.45, 0.44, 0.44, 0.43, 0.45, 0.46, 0.44, 0.44, 
    0.45, 0.49, 0.5, 0.49, 0.53, 0.53, 0.53, 0.54, 0.59, 0.66, 0.68, 0.62, 
    0.66, 0.61, 0.57, 0.6, 0.55, 0.59, 0.55, 0.58, 0.51, 0.5, 0.51, 0.54, 
    0.55, 0.64, 0.67, 0.67, 0.73, 0.72, 0.67, 0.65, 0.83, 0.65, 0.62, 0.6, 
    0.74, 0.86, 0.87, 0.88, 0.91, 0.91, 0.93, 0.94, 0.9, 0.87, 0.83, 0.8, 
    0.8, 0.86, 0.92, 0.92, 0.91, 0.86, 0.82, 0.76, 0.79, 0.77, 0.77, 0.82, 
    0.86, 0.88, 0.87, 0.84, 0.75, 0.69, 0.66, 0.67, 0.67, 0.79, 0.58, 0.59, 
    0.58, 0.6, 0.62, 0.65, 0.69, 0.71, 0.73, 0.74, 0.75, 0.72, 0.73, 0.76, 
    0.76, 0.76, 0.75, 0.7, 0.7, 0.71, 0.71, 0.72, 0.72, 0.74, 0.74, 0.72, 
    0.69, 0.66, 0.64, 0.63, 0.63, 0.65, 0.64, 0.62, 0.62, 0.68, 0.72, 0.71, 
    0.7, 0.68, 0.74, 0.85, 0.84, 0.82, 0.81, 0.78, 0.78, 0.81, 0.83, 0.8, 
    0.92, 0.8, 0.73, 0.66, 0.66, 0.67, 0.77, 0.78, 0.84, 0.69, 0.69, 0.67, 
    0.66, 0.64, 0.65, 0.64, 0.63, 0.59, 0.56, 0.57, 0.59, 0.55, 0.53, 0.51, 
    0.54, 0.49, 0.48, 0.48, 0.48, 0.5, 0.47, 0.46, 0.47, 0.46, 0.46, 0.48, 
    0.49, 0.5, 0.5, 0.5, 0.48, 0.49, 0.53, 0.6, 0.63, 0.64, 0.63, 0.7, 0.68, 
    0.68, 0.68, 0.7, 0.64, 0.66, 0.63, 0.62, 0.66, 0.59, 0.53, 0.52, 0.62, 
    0.57, 0.6, 0.63, 0.65, 0.61, 0.64, 0.57, 0.56, 0.56, 0.57, 0.59, 0.62, 
    0.64, 0.61, 0.63, 0.64, 0.66, 0.66, 0.65, 0.71, 0.69, 0.68, 0.69, 0.67, 
    0.68, 0.71, 0.7, 0.69, 0.71, 0.68, 0.62, 0.65, 0.69, 0.61, 0.6, 0.59, 
    0.65, 0.63, 0.67, 0.67, 0.68, 0.71, 0.66, 0.65, 0.62, 0.65, 0.65, 0.62, 
    0.65, 0.68, 0.71, 0.69, 0.72, 0.73, 0.72, 0.73, 0.75, 0.77, 0.81, 0.83, 
    0.85, 0.86, 0.85, 0.86, 0.91, 0.88, 0.89, 0.77, 0.68, 0.64, 0.64, 0.66, 
    0.61, 0.57, 0.59, 0.56, 0.54, 0.52, 0.48, 0.48, 0.51, 0.55, 0.63, 0.58, 
    0.51, 0.54, 0.52, 0.53, 0.58, 0.57, 0.58, 0.59, 0.57, 0.58, 0.61, 0.58, 
    0.59, 0.58, 0.58, 0.58, 0.6, 0.65, 0.63, 0.66, 0.61, 0.63, 0.61, 0.64, 
    0.62, 0.59, 0.58, 0.59, 0.61, 0.61, 0.58, 0.62, 0.59, 0.56, 0.58, 0.59, 
    0.59, 0.56, 0.58, 0.6, 0.6, 0.59, 0.61, 0.6, 0.57, 0.59, 0.6, 0.61, 0.6, 
    0.62, 0.61, 0.6, 0.59, 0.62, 0.6, 0.59, 0.6, 0.56, 0.56, 0.59, 0.59, 0.6, 
    0.62, 0.65, 0.63, 0.69, 0.66, 0.62, 0.58, 0.55, 0.54, 0.53, 0.53, 0.48, 
    0.5, 0.48, 0.55, 0.58, 0.63, 0.74, 0.75, 0.73, 0.67, 0.73, 0.77, 0.82, 
    0.81, 0.84, 0.81, 0.84, 0.77, 0.64, 0.64, 0.62, 0.57, 0.55, 0.52, 0.52, 
    0.49, 0.57, 0.61, 0.69, 0.71, 0.73, 0.83, 0.85, 0.75, 0.64, 0.64, 0.64, 
    0.63, 0.61, 0.6, 0.59, 0.56, 0.51, 0.49, 0.53, 0.53, 0.55, 0.46, 0.54, 
    0.55, 0.51, 0.53, 0.53, 0.54, 0.56, 0.59, 0.58, 0.56, 0.61, 0.6, 0.59, 
    0.56, 0.55, 0.56, 0.58, 0.6, 0.61, 0.61, 0.6, 0.59, 0.59, 0.6, 0.61, 
    0.63, 0.64, 0.67, 0.63, 0.63, 0.64, 0.61, 0.69, 0.65, 0.64, 0.7, 0.65, 
    0.7, 0.57, 0.65, 0.64, 0.65, 0.64, 0.73, 0.8, 0.82, 0.76, 0.7, 0.67, 
    0.69, 0.78, 0.79, 0.81, 0.72, 0.82, 0.86, 0.89, 0.87, 0.9, 0.92, 0.94, 
    0.94, 0.93, 0.92, 0.91, 0.92, 0.92, 0.92, 0.92, 0.92, 0.9, 0.9, 0.91, 
    0.82, 0.9, 0.73, 0.71, 0.75, 0.77, 0.71, 0.67, 0.75, 0.74, 0.72, 0.7, 
    0.68, 0.79, 0.82, 0.72, 0.65, 0.69, 0.66, 0.64, 0.63, 0.67, 0.67, 0.62, 
    0.63, 0.73, 0.64, 0.73, 0.64, 0.62, 0.72, 0.62, 0.65, 0.66, 0.64, 0.6, 
    0.56, 0.58, 0.61, 0.56, 0.54, 0.54, 0.56, 0.68, 0.68, 0.67, 0.71, 0.72, 
    0.72, 0.67, 0.73, 0.68, 0.72, 0.72, 0.76, 0.75, 0.75, 0.72, 0.65, 0.71, 
    0.63, 0.66, 0.65, 0.67, 0.63, 0.61, 0.6, 0.53, 0.51, 0.57, 0.56, 0.64, 
    0.64, 0.64, 0.66, 0.67, 0.61, 0.63, 0.61, 0.62, 0.64, 0.62, 0.64, 0.7, 
    0.71, 0.66, 0.68, 0.66, 0.62, 0.61, 0.69, 0.79, 0.84, 0.75, 0.7, 0.78, 
    0.82, 0.84, 0.84, 0.89, 0.89, 0.89, 0.9, 0.92, 0.92, 0.91, 0.94, 0.84, 
    0.81, 0.75, 0.8, 0.86, 0.88, 0.9, 0.92, 0.93, 0.93, 0.92, 0.9, 0.88, 0.9, 
    0.89, 0.91, 0.93, 0.92, 0.92, 0.92, 0.93, 0.93, 0.93, 0.94, 0.92, 0.81, 
    0.75, 0.78, 0.78, 0.77, 0.78, 0.75, 0.74, 0.67, 0.67, 0.69, 0.64, 0.59, 
    0.58, 0.53, 0.5, 0.48, 0.48, 0.49, 0.47, 0.46, 0.47, 0.46, 0.49, 0.5, 
    0.49, 0.49, 0.51, 0.55, 0.57, 0.55, 0.53, 0.54, 0.57, 0.48, 0.48, 0.43, 
    0.41, 0.42, 0.37, 0.41, 0.42, 0.42, 0.46, 0.51, 0.51, 0.54, 0.54, 0.54, 
    0.53, 0.5, 0.47, 0.43, 0.48, 0.48, 0.46, 0.47, 0.48, 0.45, 0.43, 0.44, 
    0.42, 0.46, 0.44, 0.47, 0.55, 0.5, 0.48, 0.54, 0.56, 0.65, 0.75, 0.77, 
    0.85, 0.86, 0.87, 0.87, 0.85, 0.84, 0.87, 0.82, 0.86, 0.8, 0.82, 0.82, 
    0.8, 0.73, 0.75, 0.76, 0.74, 0.72, 0.75, 0.84, 0.86, 0.9, 0.88, 0.87, 
    0.82, 0.86, 0.83, 0.77, 0.79, 0.81, 0.84, 0.86, 0.8, 0.89, 0.91, 0.93, 
    0.9, 0.92, 0.93, 0.87, 0.93, 0.88, 0.86, 0.95, 0.9, 0.68, 0.64, 0.59, 
    0.6, 0.58, 0.56, 0.57, 0.56, 0.68, 0.67, 0.71, 0.71, 0.78, 0.84, 0.81, 
    0.86, 0.91, 0.95, 0.96, 0.97, 0.94, 0.91, 0.89, 0.88, 0.92, 0.95, 0.93, 
    0.91, 0.77, 0.94, 0.87, 0.7, 0.7, 0.64, 0.67, 0.64, 0.71, 0.75, 0.79, 
    0.82, 0.8, 0.8, 0.76, 0.86, 0.82, 0.82, 0.76, 0.79, 0.81, 0.82, 0.75, 
    0.68, 0.73, 0.65, 0.74, 0.72, 0.74, 0.75, 0.76, 0.78, 0.72, 0.72, 0.77, 
    0.69, 0.74, 0.8, 0.82, 0.88, 0.85, 0.84, 0.85, 0.85, 0.89, 0.85, 0.85, 
    0.88, 0.83, 0.77, 0.83, 0.86, 0.89, 0.88, 0.85, 0.82, 0.87, 0.87, 0.77, 
    0.82, 0.91, 0.94, 0.95, 0.88, 0.88, 0.87, 0.87, 0.78, 0.81, 0.76, 0.72, 
    0.78, 0.89, 0.93, 0.88, 0.84, 0.78, 0.73, 0.74, 0.77, 0.72, 0.64, 0.71, 
    0.77, 0.71, 0.76, 0.79, 0.76, 0.76, 0.67, 0.62, 0.68, 0.69, 0.71, 0.72, 
    0.71, 0.69, 0.68, 0.71, 0.69, 0.68, 0.69, 0.7, 0.68, 0.7, 0.71, 0.71, 
    0.73, 0.8, 0.8, 0.77, 0.74, 0.7, 0.7, 0.74, 0.72, 0.7, 0.69, 0.63, 0.69, 
    0.67, 0.64, 0.65, 0.68, 0.7, 0.69, 0.72, 0.7, 0.71, 0.75, 0.75, 0.78, 
    0.8, 0.8, 0.79, 0.78, 0.81, 0.79, 0.78, 0.83, 0.84, 0.86, 0.79, 0.77, 
    0.77, 0.77, 0.79, 0.78, 0.78, 0.78, 0.77, 0.78, 0.76, 0.77, 0.77, 0.75, 
    0.77, 0.75, 0.74, 0.77, 0.78, 0.76, 0.76, 0.71, 0.7, 0.71, 0.71, 0.69, 
    0.66, 0.62, 0.59, 0.63, 0.57, 0.52, 0.5, 0.53, 0.54, 0.52, 0.46, 0.42, 
    0.43, 0.52, 0.48, 0.47, 0.48, 0.45, 0.48, 0.43, 0.45, 0.46, 0.48, 0.45, 
    0.45, 0.57, 0.6, 0.6, 0.58, 0.54, 0.52, 0.52, 0.55, 0.59, 0.62, 0.61, 
    0.59, 0.57, 0.58, 0.58, 0.59, 0.57, 0.55, 0.56, 0.53, 0.56, 0.62, 0.58, 
    0.58, 0.78, 0.78, 0.59, 0.59, 0.58, 0.6, 0.64, 0.63, 0.64, 0.64, 0.62, 
    0.6, 0.63, 0.57, 0.56, 0.54, 0.63, 0.58, 0.57, 0.55, 0.58, 0.58, 0.58, 
    0.68, 0.63, 0.62, 0.67, 0.65, 0.68, 0.66, 0.65, 0.64, 0.66, 0.57, 0.58, 
    0.56, 0.58, 0.62, 0.58, 0.56, 0.61, 0.61, 0.58, 0.6, 0.6, 0.66, 0.63, 
    0.63, 0.64, 0.62, 0.62, 0.62, 0.62, 0.6, 0.62, 0.64, 0.65, 0.63, 0.61, 
    0.63, 0.62, 0.58, 0.55, 0.54, 0.54, 0.53, 0.58, 0.59, 0.61, 0.65, 0.59, 
    0.61, 0.63, 0.62, 0.65, 0.65, 0.64, 0.63, 0.61, 0.68, 0.65, 0.67, 0.67, 
    0.68, 0.72, 0.68, 0.7, 0.7, 0.7, 0.68, 0.7, 0.7, 0.72, 0.68, 0.69, 0.67, 
    0.75, 0.68, 0.72, 0.68, 0.68, 0.73, 0.73, 0.77, 0.76, 0.74, 0.8, 0.77, 
    0.78, 0.79, 0.77, 0.78, 0.78, 0.78, 0.77, 0.81, 0.78, 0.78, 0.8, 0.79, 
    0.72, 0.74, 0.71, 0.79, 0.82, 0.82, 0.76, 0.67, 0.69, 0.66, 0.71, 0.76, 
    0.72, 0.66, 0.69, 0.72, 0.65, 0.64, 0.64, 0.67, 0.68, 0.66, 0.65, 0.68, 
    0.67, 0.7, 0.72, 0.75, 0.73, 0.71, 0.68, 0.65, 0.67, 0.68, 0.72, 0.73, 
    0.72, 0.67, 0.67, 0.67, 0.76, 0.78, 0.77, 0.72, 0.73, 0.62, 0.68, 0.81, 
    0.88, 0.86, 0.82, 0.83, 0.7, 0.7, 0.69, 0.68, 0.67, 0.68, 0.61, 0.64, 
    0.73, 0.65, 0.61, 0.65, 0.6, 0.67, 0.69, 0.73, 0.74, 0.71, 0.66, 0.63, 
    0.61, 0.69, 0.63, 0.71, 0.7, 0.71, 0.63, 0.59, 0.65, 0.7, 0.63, 0.66, 
    0.62, 0.62, 0.62, 0.63, 0.65, 0.64, 0.68, 0.76, 0.88, 0.79, 0.72, 0.78, 
    0.73, 0.71, 0.66, 0.68, 0.7, 0.72, 0.64, 0.61, 0.58, 0.67, 0.66, 0.76, 
    0.71, 0.67, 0.64, 0.6, 0.69, 0.63, 0.63, 0.6, 0.74, 0.72, 0.71, 0.64, 
    0.58, 0.63, 0.62, 0.61, 0.61, 0.63, 0.64, 0.65, 0.64, 0.62, 0.6, 0.64, 
    0.65, 0.67, 0.68, 0.72, 0.71, 0.68, 0.7, 0.72, 0.73, 0.68, 0.72, 0.67, 
    0.7, 0.72, 0.68, 0.64, 0.72, 0.73, 0.66, 0.69, 0.68, 0.73, 0.86, 0.9, 
    0.92, 0.91, 0.89, 0.87, 0.71, 0.77, 0.71, 0.69, 0.67, 0.67, 0.68, 0.74, 
    0.73, 0.75, 0.69, 0.72, 0.75, 0.76, 0.77, 0.73, 0.72, 0.74, 0.74, 0.7, 
    0.66, 0.67, 0.75, 0.82, 0.87, 0.89, 0.88, 0.86, 0.84, 0.82, 0.81, 0.83, 
    0.88, 0.9, 0.93, 0.91, 0.92, 0.92, 0.95, 0.96, 0.96, 0.96, 0.96, 0.95, 
    0.95, 0.94, 0.95, 0.91, 0.93, 0.91, 0.89, 0.88, 0.86, 0.92, 0.93, 0.95, 
    0.93, 0.95, 0.95, 0.96, 0.96, 0.95, 0.96, 0.96, 0.96, 0.97, 0.96, 0.97, 
    0.97, 0.97, 0.95, 0.96, 0.97, 0.97, 0.95, 0.93, 0.9, 0.9, 0.93, 0.91, 
    0.89, 0.88, 0.85, 0.82, 0.81, 0.82, 0.79, 0.76, 0.75, 0.81, 0.83, 0.72, 
    0.78, 0.71, 0.65, 0.69, 0.68, 0.69, 0.71, 0.79, 0.7, 0.72, 0.78, 0.85, 
    0.85, 0.79, 0.79, 0.73, 0.72, 0.72, 0.72, 0.73, 0.71, 0.73, 0.7, 0.7, 
    0.69, 0.7, 0.68, 0.64, 0.67, 0.63, 0.63, 0.63, 0.6, 0.66, 0.62, 0.68, 
    0.63, 0.68, 0.73, 0.7, 0.66, 0.67, 0.69, 0.71, 0.74, 0.73, 0.72, 0.71, 
    0.71, 0.72, 0.67, 0.68, 0.69, 0.67, 0.65, 0.61, 0.61, 0.61, 0.61, 0.63, 
    0.58, 0.63, 0.6, 0.58, 0.57, 0.6, 0.53, 0.55, 0.55, 0.52, 0.51, 0.49, 
    0.51, 0.48, 0.49, 0.52, 0.53, 0.5, 0.53, 0.51, 0.5, 0.5, 0.49, 0.47, 0.5, 
    0.51, 0.5, 0.46, 0.51, 0.49, 0.5, 0.52, 0.47, 0.48, 0.5, 0.48, 0.45, 0.5, 
    0.51, 0.47, 0.46, 0.44, 0.45, 0.46, 0.44, 0.45, 0.43, 0.44, 0.46, 0.48, 
    0.5, 0.52, 0.54, 0.54, 0.54, 0.6, 0.64, 0.64, 0.68, 0.73, 0.68, 0.65, 
    0.66, 0.65, 0.65, 0.63, 0.6, 0.55, 0.6, 0.64, 0.84, 0.87, 0.79, 0.69, 
    0.6, 0.59, 0.77, 0.59, 0.64, 0.67, 0.67, 0.65, 0.63, 0.68, 0.64, 0.62, 
    0.62, 0.61, 0.6, 0.59, 0.54, 0.54, 0.54, 0.57, 0.54, 0.51, 0.52, 0.51, 
    0.5, 0.5, 0.5, 0.49, 0.55, 0.57, 0.59, 0.62, 0.64, 0.6, 0.57, 0.55, 0.56, 
    0.62, 0.56, 0.49, 0.51, 0.51, 0.5, 0.54, 0.56, 0.53, 0.48, 0.5, 0.49, 
    0.54, 0.53, 0.55, 0.55, 0.49, 0.5, 0.5, 0.5, 0.5, 0.5, 0.49, 0.5, 0.5, 
    0.52, 0.53, 0.55, 0.57, 0.52, 0.55, 0.51, 0.52, 0.52, 0.53, 0.52, 0.51, 
    0.47, 0.48, 0.52, 0.45, 0.51, 0.52, 0.55, 0.51, 0.5, 0.5, 0.49, 0.51, 
    0.52, 0.53, 0.5, 0.55, 0.49, 0.5, 0.51, 0.52, 0.53, 0.56, 0.55, 0.55, 
    0.54, 0.57, 0.54, 0.51, 0.49, 0.52, 0.45, 0.43, 0.43, 0.43, 0.43, 0.44, 
    0.47, 0.46, 0.47, 0.48, 0.47, 0.46, 0.47, 0.47, 0.46, 0.47, 0.49, 0.48, 
    0.5, 0.49, 0.49, 0.5, 0.53, 0.55, 0.52, 0.54, 0.5, 0.49, 0.51, 0.61, 0.6, 
    0.58, 0.63, 0.58, 0.62, 0.64, 0.59, 0.64, 0.63, 0.62, 0.63, 0.68, 0.69, 
    0.69, 0.71, 0.75, 0.75, 0.71, 0.7, 0.73, 0.78, 0.8, 0.8, 0.78, 0.81, 0.8, 
    0.78, 0.79, 0.77, 0.76, 0.75, 0.73, 0.71, 0.67, 0.64, 0.7, 0.67, 0.65, 
    0.7, 0.63, 0.62, 0.62, 0.63, 0.6, 0.63, 0.6, 0.6, 0.61, 0.63, 0.6, 0.62, 
    0.65, 0.62, 0.59, 0.61, 0.62, 0.56, 0.59, 0.59, 0.59, 0.6, 0.58, 0.6, 
    0.52, 0.57, 0.54, 0.53, 0.61, 0.56, 0.58, 0.56, 0.51, 0.55, 0.57, 0.6, 
    0.63, 0.61, 0.61, 0.59, 0.55, 0.51, 0.53, 0.59, 0.62, 0.57, 0.54, 0.56, 
    0.57, 0.59, 0.58, 0.55, 0.54, 0.62, 0.57, 0.57, 0.47, 0.43, 0.43, 0.5, 
    0.43, 0.43, 0.43, 0.69, 0.44, 0.45, 0.46, 0.46, 0.46, 0.59, 0.55, 0.54, 
    0.49, 0.49, 0.55, 0.64, 0.6, 0.59, 0.51, 0.5, 0.5, 0.5, 0.48, 0.49, 0.5, 
    0.46, 0.47, 0.51, 0.51, 0.49, 0.51, 0.51, 0.5, 0.5, 0.49, 0.52, 0.54, 
    0.55, 0.56, 0.59, 0.59, 0.61, 0.65, 0.58, 0.62, 0.61, 0.61, 0.62, 0.65, 
    0.63, 0.64, 0.65, 0.64, 0.67, 0.66, 0.65, 0.72, 0.72, 0.72, 0.75, 0.74, 
    0.71, 0.73, 0.74, 0.73, 0.73, 0.76, 0.77, 0.75, 0.75, 0.71, 0.74, 0.77, 
    0.72, 0.7, 0.88, 0.68, 0.68, 0.72, 0.65, 0.65, 0.65, 0.63, 0.61, 0.6, 
    0.58, 0.62, 0.63, 0.64, 0.68, 0.66, 0.68, 0.67, 0.7, 0.69, 0.7, 0.72, 
    0.76, 0.78, 0.83, 0.72, 0.66, 0.59, 0.59, 0.61, 0.59, 0.59, 0.57, 0.65, 
    0.68, 0.64, 0.66, 0.66, 0.64, 0.64, 0.62, 0.63, 0.6, 0.61, 0.63, 0.61, 
    0.62, 0.57, 0.56, 0.56, 0.64, 0.67, 0.68, 0.74, 0.72, 0.66, 0.68, 0.72, 
    0.69, 0.57, 0.56, 0.69, 0.63, 0.64, 0.67, 0.71, 0.67, 0.71, 0.7, 0.7, 
    0.68, 0.68, 0.62, 0.61, 0.61, 0.59, 0.64, 0.63, 0.72, 0.71, 0.73, 0.68, 
    0.67, 0.69, 0.79, 0.81, 0.78, 0.72, 0.66, 0.68, 0.61, 0.67, 0.64, 0.62, 
    0.71, 0.81, 0.89, 0.87, 0.86, 0.85, 0.81, 0.86, 0.82, 0.83, 0.85, 0.93, 
    0.94, 0.88, 0.89, 0.86, 0.88, 0.91, 0.91, 0.94, 0.95, 0.89, 0.84, 0.85, 
    0.84, 0.77, 0.81, 0.8, 0.8, 0.81, 0.79, 0.74, 0.72, 0.69, 0.68, 0.73, 
    0.71, 0.71, 0.7, 0.68, 0.61, 0.71, 0.71, 0.72, 0.57, 0.65, 0.61, 0.7, 
    0.68, 0.67, 0.67, 0.64, 0.61, 0.67, 0.69, 0.76, 0.85, 0.88, 0.87, 0.84, 
    0.82, 0.8, 0.82, 0.83, 0.76, 0.77, 0.77, 0.78, 0.79, 0.81, 0.8, 0.69, 
    0.9, 0.93, 0.92, 0.91, 0.79, 0.74, 0.73, 0.73, 0.72, 0.73, 0.75, 0.74, 
    0.77, 0.65, 0.79, 0.76, 0.77, 0.72, 0.77, 0.71, 0.79, 0.74, 0.68, 0.7, 
    0.7, 0.67, 0.69, 0.73, 0.7, 0.7, 0.67, 0.71, 0.71, 0.68, 0.82, 0.89, 
    0.86, 0.85, 0.89, 0.87, 0.85, 0.81, 0.85, 0.87, 0.88, 0.91, 0.92, 0.91, 
    0.92, 0.93, 0.94, 0.93, 0.93, 0.92, 0.9, 0.88, 0.84, 0.81, 0.79, 0.72, 
    0.79, 0.75, 0.66, 0.62, 0.61, 0.6, 0.58, 0.6, 0.62, 0.57, 0.58, 0.58, 
    0.58, 0.57, 0.56, 0.58, 0.6, 0.59, 0.58, 0.56, 0.56, 0.58, 0.59, 0.6, 
    0.65, 0.65, 0.62, 0.64, 0.68, 0.68, 0.63, 0.61, 0.64, 0.7, 0.69, 0.68, 
    0.69, 0.73, 0.66, 0.67, 0.68, 0.66, 0.65, 0.71, 0.67, 0.64, 0.69, 0.64, 
    0.68, 0.64, 0.66, 0.59, 0.66, 0.66, 0.71, 0.71, 0.64, 0.55, 0.56, 0.56, 
    0.57, 0.62, 0.62, 0.63, 0.65, 0.62, 0.6, 0.63, 0.61, 0.55, 0.57, 0.61, 
    0.64, 0.62, 0.57, 0.59, 0.57, 0.57, 0.57, 0.63, 0.62, 0.6, 0.62, 0.64, 
    0.62, 0.67, 0.63, 0.66, 0.67, 0.63, 0.65, 0.66, 0.68, 0.71, 0.69, 0.7, 
    0.66, 0.71, 0.71, 0.7, 0.68, 0.73, 0.71, 0.73, 0.76, 0.77, 0.77, 0.71, 
    0.75, 0.63, 0.64, 0.69, 0.68, 0.66, 0.66, 0.7, 0.63, 0.71, 0.61, 0.69, 
    0.7, 0.68, 0.67, 0.66, 0.69, 0.67, 0.64, 0.7, 0.69, 0.7, 0.7, 0.73, 0.73, 
    0.75, 0.69, 0.72, 0.75, 0.71, 0.73, 0.76, 0.73, 0.73, 0.72, 0.71, 0.72, 
    0.73, 0.72, 0.73, 0.73, 0.75, 0.75, 0.72, 0.73, 0.74, 0.83, 0.84, 0.86, 
    0.86, 0.87, 0.82, 0.85, 0.85, 0.86, 0.86, 0.89, 0.85, 0.82, 0.75, 0.79, 
    0.79, 0.72, 0.77, 0.73, 0.73, 0.75, 0.71, 0.79, 0.77, 0.73, 0.72, 0.75, 
    0.74, 0.75, 0.76, 0.76, 0.73, 0.76, 0.72, 0.73, 0.72, 0.72, 0.7, 0.7, 
    0.72, 0.73, 0.75, 0.73, 0.7, 0.73, 0.74, 0.74, 0.75, 0.76, 0.7, 0.71, 
    0.69, 0.67, 0.67, 0.69, 0.64, 0.66, 0.71, 0.77, 0.88, 0.9, 0.89, 0.85, 
    0.84, 0.84, 0.85, 0.79, 0.83, 0.87, 0.81, 0.83, 0.79, 0.76, 0.76, 0.71, 
    0.66, 0.66, 0.58, 0.57, 0.56, 0.58, 0.57, 0.76, 0.74, 0.83, 0.93, 0.87, 
    0.88, 0.85, 0.89, 0.92, 0.88, 0.92, 0.95, 0.94, 0.83, 0.78, 0.7, 0.71, 
    0.69, 0.69, 0.78, 0.88, 0.82, 0.73, 0.68, 0.65, 0.69, 0.74, 0.71, 0.68, 
    0.66, 0.68, 0.77, 0.88, 0.87, 0.85, 0.81, 0.75, 0.71, 0.7, 0.72, 0.7, 
    0.65, 0.71, 0.75, 0.73, 0.82, 0.83, 0.81, 0.8, 0.81, 0.8, 0.7, 0.63, 
    0.63, 0.65, 0.7, 0.71, 0.71, 0.76, 0.78, 0.84, 0.85, 0.86, 0.88, 0.94, 
    0.95, 0.96, 0.95, 0.95, 0.96, 0.95, 0.95, 0.94, 0.94, 0.89, 0.93, 0.95, 
    0.9, 0.89, 0.83, 0.84, 0.88, 0.92, 0.92, 0.93, 0.87, 0.77, 0.77, 0.76, 
    0.75, 0.73, 0.72, 0.72, 0.73, 0.71, 0.74, 0.75, 0.72, 0.73, 0.74, 0.75, 
    0.76, 0.77, 0.79, 0.84, 0.87, 0.85, 0.83, 0.86, 0.86, 0.88, 0.88, 0.86, 
    0.89, 0.86, 0.85, 0.85, 0.86, 0.89, 0.88, 0.87, 0.84, 0.82, 0.82, 0.78, 
    0.79, 0.83, 0.79, 0.78, 0.78, 0.78, 0.78, 0.73, 0.75, 0.72, 0.68, 0.71, 
    0.64, 0.66, 0.71, 0.67, 0.75, 0.76, 0.75, 0.76, 0.68, 0.71, 0.7, 0.71, 
    0.72, 0.68, 0.68, 0.65, 0.67, 0.69, 0.73, 0.74, 0.74, 0.74, 0.73, 0.82, 
    0.69, 0.72, 0.71, 0.69, 0.68, 0.73, 0.71, 0.71, 0.66, 0.68, 0.75, 0.7, 
    0.71, 0.73, 0.69, 0.72, 0.75, 0.7, 0.79, 0.8, 0.8, 0.87, 0.81, 0.81, 
    0.77, 0.82, 0.78, 0.78, 0.8, 0.81, 0.78, 0.79, 0.79, 0.81, 0.81, 0.8, 
    0.8, 0.82, 0.83, 0.84, 0.85, 0.85, 0.82, 0.8, 0.79, 0.78, 0.79, 0.77, 
    0.76, 0.77, 0.78, 0.78, 0.81, 0.81, 0.87, 0.88, 0.88, 0.9, 0.9, 0.84, 
    0.79, 0.89, 0.86, 0.93, 0.91, 0.82, 0.78, 0.81, 0.77, 0.71, 0.84, 0.93, 
    0.95, 0.93, 0.92, 0.91, 0.77, 0.71, 0.75, 0.77, 0.69, 0.66, 0.71, 0.74, 
    0.68, 0.6, 0.67, 0.64, 0.73, 0.67, 0.6, 0.64, 0.65, 0.75, 0.78, 0.84, 
    0.82, 0.76, 0.82, 0.76, 0.8, 0.76, 0.79, 0.85, 0.8, 0.81, 0.85, 0.85, 
    0.79, 0.85, 0.79, 0.74, 0.77, 0.75, 0.75, 0.8, 0.75, 0.8, 0.81, 0.75, 
    0.63, 0.65, 0.68, 0.64, 0.61, 0.54, 0.59, 0.58, 0.56, 0.58, 0.6, 0.62, 
    0.65, 0.66, 0.66, 0.7, 0.72, 0.77, 0.84, 0.85, 0.88, 0.91, 0.92, 0.92, 
    0.94, 0.94, 0.93, 0.94, 0.93, 0.94, 0.93, 0.7, 0.66, 0.61, 0.6, 0.64, 
    0.68, 0.67, 0.74, 0.68, 0.69, 0.64, 0.66, 0.65, 0.63, 0.63, 0.68, 0.58, 
    0.61, 0.66, 0.67, 0.7, 0.64, 0.64, 0.64, 0.69, 0.71, 0.64, 0.59, 0.5, 
    0.46, 0.45, 0.44, 0.46, 0.51, 0.58, 0.59, 0.47, 0.45, 0.53, 0.49, 0.45, 
    0.45, 0.44, 0.44, 0.46, 0.49, 0.47, 0.53, 0.54, 0.51, 0.5, 0.47, 0.46, 
    0.45, 0.48, 0.57, 0.52, 0.5, 0.48, 0.49, 0.5, 0.59, 0.56, 0.53, 0.51, 
    0.51, 0.5, 0.49, 0.51, 0.5, 0.55, 0.54, 0.57, 0.57, 0.6, 0.57, 0.61, 
    0.61, 0.49, 0.49, 0.55, 0.51, 0.51, 0.51, 0.51, 0.51, 0.51, 0.54, 0.59, 
    0.61, 0.68, 0.61, 0.61, 0.63, 0.61, 0.65, 0.6, 0.64, 0.62, 0.61, 0.68, 
    0.59, 0.59, 0.58, 0.59, 0.61, 0.63, 0.59, 0.64, 0.65, 0.62, 0.62, 0.62, 
    0.62, 0.66, 0.7, 0.67, 0.66, 0.68, 0.67, 0.68, 0.64, 0.63, 0.61, 0.59, 
    0.56, 0.59, 0.59, 0.64, 0.57, 0.66, 0.62, 0.65, 0.65, 0.67, 0.65, 0.66, 
    0.66, 0.65, 0.68, 0.65, 0.66, 0.67, 0.68, 0.64, 0.67, 0.67, 0.66, 0.64, 
    0.59, 0.59, 0.59, 0.57, 0.58, 0.62, 0.63, 0.65, 0.64, 0.63, 0.62, 0.66, 
    0.66, 0.69, 0.69, 0.67, 0.67, 0.69, 0.69, 0.64, 0.66, 0.61, 0.61, 0.57, 
    0.57, 0.54, 0.59, 0.56, 0.61, 0.63, 0.6, 0.67, 0.64, 0.62, 0.66, 0.68, 
    0.69, 0.66, 0.69, 0.66, 0.68, 0.67, 0.64, 0.68, 0.66, 0.57, 0.6, 0.58, 
    0.59, 0.53, 0.57, 0.6, 0.57, 0.57, 0.56, 0.62, 0.63, 0.63, 0.69, 0.71, 
    0.71, 0.72, 0.74, 0.79, 0.79, 0.78, 0.77, 0.77, 0.72, 0.67, 0.62, 0.63, 
    0.6, 0.57, 0.57, 0.61, 0.54, 0.6, 0.63, 0.69, 0.7, 0.7, 0.7, 0.68, 0.7, 
    0.72, 0.71, 0.69, 0.66, 0.62, 0.65, 0.62, 0.68, 0.59, 0.55, 0.55, 0.54, 
    0.49, 0.55, 0.51, 0.56, 0.59, 0.57, 0.6, 0.62, 0.63, 0.61, 0.6, 0.59, 
    0.62, 0.71, 0.65, 0.68, 0.65, 0.69, 0.7, 0.63, 0.6, 0.58, 0.56, 0.55, 
    0.57, 0.55, 0.57, 0.6, 0.56, 0.6, 0.6, 0.62, 0.64, 0.63, 0.65, 0.65, 
    0.67, 0.76, 0.8, 0.89, 0.81, 0.76, 0.62, 0.59, 0.62, 0.61, 0.62, 0.61, 
    0.57, 0.53, 0.49, 0.57, 0.54, 0.57, 0.54, 0.56, 0.57, 0.56, 0.59, 0.58, 
    0.63, 0.63, 0.65, 0.7, 0.61, 0.6, 0.69, 0.69, 0.68, 0.69, 0.63, 0.64, 
    0.7, 0.66, 0.65, 0.69, 0.73, 0.89, 0.92, 0.94, 0.94, 0.8, 0.85, 0.84, 
    0.77, 0.77, 0.69, 0.7, 0.73, 0.65, 0.59, 0.66, 0.67, 0.66, 0.66, 0.67, 
    0.6, 0.68, 0.63, 0.57, 0.61, 0.63, 0.65, 0.69, 0.56, 0.63, 0.65, 0.62, 
    0.66, 0.6, 0.61, 0.59, 0.64, 0.61, 0.55, 0.55, 0.53, 0.6, 0.59, 0.56, 
    0.51, 0.55, 0.56, 0.55, 0.52, 0.51, 0.52, 0.52, 0.5, 0.5, 0.53, 0.55, 
    0.58, 0.58, 0.6, 0.56, 0.53, 0.57, 0.57, 0.54, 0.56, 0.53, 0.51, 0.5, 
    0.49, 0.49, 0.55, 0.55, 0.55, 0.57, 0.56, 0.54, 0.57, 0.54, 0.52, 0.61, 
    0.64, 0.64, 0.62, 0.66, 0.65, 0.67, 0.7, 0.61, 0.57, 0.56, 0.58, 0.58, 
    0.57, 0.54, 0.51, 0.59, 0.59, 0.57, 0.61, 0.66, 0.71, 0.65, 0.62, 0.62, 
    0.69, 0.72, 0.72, 0.69, 0.73, 0.76, 0.74, 0.76, 0.76, 0.8, 0.78, 0.81, 
    0.8, 0.79, 0.83, 0.84, 0.83, 0.84, 0.84, 0.84, 0.85, 0.86, 0.87, 0.89, 
    0.89, 0.89, 0.89, 0.89, 0.87, 0.9, 0.88, 0.88, 0.85, 0.85, 0.79, 0.84, 
    0.73, 0.75, 0.75, 0.78, 0.82, 0.77, 0.75, 0.75, 0.77, 0.79, 0.76, 0.76, 
    0.81, 0.84, 0.82, 0.76, 0.77, 0.78, 0.75, 0.76, 0.79, 0.77, 0.74, 0.62, 
    0.62, 0.64, 0.63, 0.63, 0.65, 0.66, 0.65, 0.68, 0.68, 0.68, 0.68, 0.69, 
    0.71, 0.69, 0.71, 0.73, 0.76, 0.75, 0.72, 0.73, 0.72, 0.69, 0.7, 0.68, 
    0.66, 0.67, 0.7, 0.7, 0.75, 0.77, 0.74, 0.74, 0.73, 0.71, 0.69, 0.71, 
    0.71, 0.72, 0.72, 0.77, 0.81, 0.79, 0.76, 0.69, 0.64, 0.62, 0.63, 0.65, 
    0.65, 0.65, 0.63, 0.64, 0.68, 0.7, 0.68, 0.71, 0.74, 0.75, 0.78, 0.8, 
    0.78, 0.77, 0.82, 0.76, 0.77, 0.75, 0.81, 0.78, 0.79, 0.75, 0.8, 0.77, 
    0.79, 0.8, 0.8, 0.8, 0.74, 0.76, 0.8, 0.84, 0.86, 0.87, 0.87, 0.87, 0.9, 
    0.86, 0.85, 0.88, 0.88, 0.87, 0.85, 0.82, 0.81, 0.77, 0.78, 0.73, 0.78, 
    0.73, 0.74, 0.7, 0.75, 0.74, 0.78, 0.8, 0.82, 0.83, 0.83, 0.84, 0.78, 
    0.8, 0.79, 0.76, 0.78, 0.81, 0.75, 0.8, 0.85, 0.77, 0.82, 0.81, 0.85, 
    0.82, 0.82, 0.78, 0.76, 0.65, 0.64, 0.64, 0.64, 0.63, 0.63, 0.61, 0.63, 
    0.61, 0.63, 0.63, 0.6, 0.59, 0.59, 0.59, 0.57, 0.57, 0.59, 0.56, 0.58, 
    0.55, 0.57, 0.59, 0.6, 0.54, 0.55, 0.55, 0.58, 0.64, 0.66, 0.6, 0.61, 
    0.67, 0.6, 0.66, 0.66, 0.55, 0.58, 0.52, 0.51, 0.56, 0.53, 0.52, 0.57, 
    0.56, 0.51, 0.56, 0.52, 0.52, 0.55, 0.56, 0.56, 0.57, 0.59, 0.59, 0.58, 
    0.6, 0.59, 0.62, 0.62, 0.61, 0.57, 0.6, 0.6, 0.58, 0.59, 0.62, 0.64, 
    0.63, 0.6, 0.57, 0.55, 0.55, 0.55, 0.54, 0.59, 0.61, 0.59, 0.6, 0.62, 
    0.61, 0.62, 0.62, 0.63, 0.66, 0.62, 0.63, 0.59, 0.59, 0.62, 0.57, 0.56, 
    0.6, 0.62, 0.62, 0.6, 0.61, 0.62, 0.64, 0.69, 0.69, 0.68, 0.72, 0.69, 
    0.71, 0.66, 0.71, 0.64, 0.6, 0.66, 0.61, 0.58, 0.59, 0.5, 0.51, 0.51, 
    0.53, 0.55, 0.55, 0.51, 0.52, 0.5, 0.52, 0.55, 0.57, 0.57, 0.55, 0.58, 
    0.58, 0.6, 0.61, 0.6, 0.6, 0.58, 0.54, 0.57, 0.56, 0.53, 0.52, 0.56, 
    0.58, 0.52, 0.53, 0.55, 0.56, 0.58, 0.56, 0.6, 0.59, 0.61, 0.61, 0.64, 
    0.65, 0.67, 0.68, 0.7, 0.69, 0.64, 0.61, 0.61, 0.59, 0.57, 0.55, 0.57, 
    0.6, 0.59, 0.59, 0.62, 0.61, 0.63, 0.63, 0.67, 0.68, 0.68, 0.68, 0.7, 
    0.7, 0.67, 0.7, 0.65, 0.67, 0.62, 0.59, 0.58, 0.6, 0.59, 0.57, 0.53, 
    0.51, 0.55, 0.54, 0.58, 0.58, 0.58, 0.59, 0.6, 0.61, 0.61, 0.6, 0.59, 
    0.59, 0.61, 0.58, 0.63, 0.63, 0.63, 0.6, 0.63, 0.61, 0.56, 0.58, 0.58, 
    0.58, 0.63, 0.6, 0.57, 0.62, 0.6, 0.63, 0.64, 0.68, 0.66, 0.67, 0.67, 
    0.69, 0.71, 0.73, 0.67, 0.7, 0.67, 0.64, 0.53, 0.59, 0.51, 0.61, 0.62, 
    0.62, 0.62, 0.62, 0.62, 0.6, 0.64, 0.66, 0.67, 0.67, 0.68, 0.69, 0.7, 
    0.69, 0.68, 0.75, 0.7, 0.65, 0.63, 0.62, 0.56, 0.56, 0.56, 0.54, 0.56, 
    0.59, 0.59, 0.57, 0.57, 0.6, 0.57, 0.58, 0.63, 0.67, 0.66, 0.68, 0.74, 
    0.69, 0.76, 0.71, 0.68, 0.64, 0.64, 0.6, 0.51, 0.54, 0.61, 0.62, 0.62, 
    0.62, 0.64, 0.61, 0.58, 0.6, 0.56, 0.58, 0.63, 0.66, 0.69, 0.71, 0.65, 
    0.76, 0.76, 0.78, 0.72, 0.65, 0.7, 0.73, 0.72, 0.82, 0.76, 0.73, 0.68, 
    0.71, 0.68, 0.66, 0.68, 0.73, 0.73, 0.72, 0.77, 0.75, 0.82, 0.86, 0.9, 
    0.91, 0.92, 0.92, 0.88, 0.88, 0.85, 0.72, 0.74, 0.75, 0.64, 0.6, 0.57, 
    0.51, 0.62, 0.67, 0.6, 0.64, 0.68, 0.67, 0.69, 0.73, 0.76, 0.75, 0.74, 
    0.73, 0.7, 0.69, 0.67, 0.68, 0.67, 0.64, 0.66, 0.6, 0.59, 0.57, 0.57, 
    0.56, 0.58, 0.58, 0.6, 0.62, 0.65, 0.66, 0.68, 0.68, 0.72, 0.69, 0.7, 
    0.72, 0.7, 0.69, 0.73, 0.68, 0.67, 0.61, 0.6, 0.63, 0.61, 0.6, 0.59, 
    0.56, 0.62, 0.58, 0.57, 0.69, 0.63, 0.64, 0.67, 0.7, 0.72, 0.73, 0.75, 
    0.75, 0.73, 0.75, 0.77, 0.75, 0.73, 0.67, 0.54, 0.59, 0.58, 0.53, 0.57, 
    0.57, 0.62, 0.56, 0.57, 0.57, 0.56, 0.54, 0.56, 0.59, 0.51, 0.53, 0.59, 
    0.49, 0.59, 0.54, 0.54, 0.56, 0.55, 0.56, 0.56, 0.5, 0.55, 0.61, 0.58, 
    0.6, 0.59, 0.65, 0.58, 0.61, 0.57, 0.58, 0.63, 0.71, 0.72, 0.69, 0.71, 
    0.65, 0.65, 0.69, 0.78, 0.63, 0.72, 0.59, 0.53, 0.49, 0.56, 0.61, 0.61, 
    0.61, 0.63, 0.68, 0.65, 0.65, 0.61, 0.61, 0.67, 0.73, 0.7, 0.68, 0.75, 
    0.72, 0.67, 0.67, 0.72, 0.64, 0.67, 0.58, 0.58, 0.57, 0.62, 0.58, 0.59, 
    0.6, 0.56, 0.62, 0.6, 0.58, 0.66, 0.64, 0.65, 0.7, 0.71, 0.79, 0.78, 
    0.79, 0.8, 0.82, 0.7, 0.65, 0.68, 0.61, 0.63, 0.52, 0.52, 0.59, 0.66, 
    0.57, 0.64, 0.59, 0.54, 0.63, 0.62, 0.73, 0.71, 0.77, 0.84, 0.81, 0.81, 
    0.82, 0.82, 0.83, 0.79, 0.79, 0.9, 0.9, 0.9, 0.89, 0.9, 0.9, 0.92, 0.9, 
    0.92, 0.93, 0.91, 0.9, 0.88, 0.9, 0.89, 0.9, 0.88, 0.84, 0.83, 0.92, 
    0.94, 0.95, 0.93, 0.93, 0.92, 0.85, 0.78, 0.69, 0.65, 0.76, 0.69, 0.73, 
    0.76, 0.76, 0.84, 0.85, 0.85, 0.84, 0.85, 0.86, 0.86, 0.87, 0.88, 0.87, 
    0.87, 0.87, 0.87, 0.88, 0.84, 0.82, 0.81, 0.8, 0.81, 0.82, 0.81, 0.79, 
    0.8, 0.82, 0.84, 0.78, 0.79, 0.79, 0.79, 0.8, 0.8, 0.79, 0.79, 0.8, 0.78, 
    0.83, 0.8, 0.8, 0.8, 0.79, 0.77, 0.77, 0.75, 0.75, 0.72, 0.76, 0.74, 
    0.75, 0.74, 0.72, 0.74, 0.77, 0.77, 0.76, 0.69, 0.67, 0.65, 0.62, 0.61, 
    0.63, 0.61, 0.61, 0.61, 0.61, 0.63, 0.62, 0.59, 0.62, 0.57, 0.61, 0.63, 
    0.6, 0.62, 0.65, 0.61, 0.65, 0.62, 0.62, 0.65, 0.67, 0.67, 0.64, 0.63, 
    0.63, 0.76, 0.73, 0.71, 0.65, 0.64, 0.63, 0.63, 0.63, 0.63, 0.65, 0.68, 
    0.7, 0.71, 0.67, 0.67, 0.67, 0.67, 0.7, 0.69, 0.66, 0.67, 0.69, 0.68, 
    0.67, 0.66, 0.69, 0.67, 0.67, 0.65, 0.69, 0.66, 0.67, 0.69, 0.72, 0.68, 
    0.66, 0.7, 0.68, 0.66, 0.69, 0.68, 0.66, 0.7, 0.65, 0.68, 0.62, 0.62, 
    0.64, 0.69, 0.73, 0.68, 0.7, 0.67, 0.68, 0.63, 0.67, 0.68, 0.71, 0.67, 
    0.63, 0.64, 0.63, 0.64, 0.71, 0.67, 0.76, 0.72, 0.75, 0.78, 0.79, 0.81, 
    0.83, 0.86, 0.85, 0.87, 0.86, 0.81, 0.88, 0.85, 0.82, 0.83, 0.88, 0.87, 
    0.88, 0.87, 0.89, 0.88, 0.88, 0.89, 0.92, 0.92, 0.75, 0.77, 0.73, 0.71, 
    0.76, 0.8, 0.77, 0.71, 0.65, 0.65, 0.66, 0.67, 0.72, 0.73, 0.64, 0.72, 
    0.8, 0.7, 0.67, 0.7, 0.67, 0.71, 0.71, 0.73, 0.71, 0.74, 0.77, 0.82, 
    0.87, 0.78, 0.7, 0.72, 0.71, 0.7, 0.67, 0.66, 0.68, 0.64, 0.62, 0.64, 
    0.66, 0.66, 0.67, 0.68, 0.66, 0.64, 0.64, 0.65, 0.61, 0.62, 0.58, 0.57, 
    0.55, 0.56, 0.57, 0.57, 0.55, 0.59, 0.58, 0.6, 0.61, 0.63, 0.66, 0.68, 
    0.7, 0.69, 0.68, 0.66, 0.68, 0.66, 0.66, 0.68, 0.66, 0.66, 0.67, 0.7, 
    0.71, 0.71, 0.68, 0.68, 0.7, 0.71, 0.7, 0.71, 0.71, 0.71, 0.68, 0.7, 
    0.67, 0.67, 0.68, 0.7, 0.7, 0.69, 0.69, 0.71, 0.7, 0.72, 0.74, 0.68, 
    0.64, 0.6, 0.56, 0.54, 0.58, 0.56, 0.54, 0.53, 0.54, 0.57, 0.56, 0.6, 
    0.65, 0.85, 0.72, 0.61, 0.62, 0.59, 0.58, 0.6, 0.59, 0.59, 0.58, 0.6, 
    0.62, 0.62, 0.67, 0.73, 0.75, 0.75, 0.79, 0.87, 0.86, 0.88, 0.91, 0.91, 
    0.92, 0.86, 0.86, 0.85, 0.84, 0.85, 0.83, 0.67, 0.67, 0.68, 0.65, 0.67, 
    0.65, 0.64, 0.63, 0.64, 0.64, 0.65, 0.66, 0.66, 0.65, 0.77, 0.63, 0.61, 
    0.6, 0.64, 0.56, 0.63, 0.63, 0.55, 0.57, 0.68, 0.68, 0.72, 0.74, 0.73, 
    0.7, 0.72, 0.71, 0.68, 0.59, 0.61, 0.6, 0.59, 0.6, 0.6, 0.61, 0.56, 0.53, 
    0.52, 0.47, 0.49, 0.44, 0.43, 0.39, 0.44, 0.52, 0.47, 0.51, 0.46, 0.44, 
    0.52, 0.51, 0.51, 0.52, 0.51, 0.52, 0.53, 0.55, 0.61, 0.59, 0.67, 0.65, 
    0.63, 0.63, 0.63, 0.62, 0.65, 0.64, 0.65, 0.64, 0.65, 0.64, 0.64, 0.62, 
    0.62, 0.63, 0.63, 0.61, 0.61, 0.62, 0.61, 0.67, 0.72, 0.82, 0.86, 0.89, 
    0.89, 0.87, 0.83, 0.78, 0.84, 0.83, 0.77, 0.78, 0.79, 0.84, 0.86, 0.88, 
    0.86, 0.88, 0.87, 0.86, 0.84, 0.79, 0.72, 0.71, 0.6, 0.64, 0.58, 0.61, 
    0.63, 0.68, 0.69, 0.64, 0.58, 0.64, 0.7, 0.66, 0.67, 0.73, 0.73, 0.72, 
    0.7, 0.73, 0.72, 0.75, 0.76, 0.84, 0.82, 0.64, 0.71, 0.72, 0.64, 0.7, 
    0.68, 0.68, 0.74, 0.71, 0.74, 0.76, 0.77, 0.77, 0.75, 0.77, 0.75, 0.74, 
    0.72, 0.69, 0.66, 0.65, 0.6, 0.79, 0.73, 0.76, 0.66, 0.7, 0.68, 0.58, 
    0.61, 0.62, 0.6, 0.63, 0.62, 0.63, 0.67, 0.7, 0.74, 0.64, 0.61, 0.68, 
    0.67, 0.68, 0.69, 0.72, 0.77, 0.78, 0.86, 0.85, 0.87, 0.85, 0.83, 0.8, 
    0.8, 0.81, 0.8, 0.82, 0.86, 0.88, 0.88, 0.86, 0.88, 0.88, 0.87, 0.79, 
    0.8, 0.78, 0.82, 0.84, 0.8, 0.73, 0.72, 0.72, 0.69, 0.66, 0.68, 0.68, 
    0.69, 0.72, 0.72, 0.69, 0.7, 0.73, 0.74, 0.76, 0.76, 0.74, 0.74, 0.75, 
    0.74, 0.74, 0.76, 0.72, 0.71, 0.71, 0.69, 0.71, 0.67, 0.77, 0.88, 0.84, 
    0.86, 0.87, 0.87, 0.87, 0.83, 0.77, 0.76, 0.74, 0.77, 0.71, 0.68, 0.7, 
    0.69, 0.67, 0.66, 0.68, 0.68, 0.68, 0.67, 0.7, 0.71, 0.75, 0.79, 0.79, 
    0.77, 0.81, 0.81, 0.78, 0.78, 0.79, 0.78, 0.81, 0.84, 0.78, 0.81, 0.82, 
    0.76, 0.72, 0.69, 0.71, 0.73, 0.69, 0.66, 0.64, 0.7, 0.74, 0.72, 0.69, 
    0.72, 0.67, 0.86, 0.75, 0.77, 0.7, 0.68, 0.74, 0.69, 0.74, 0.82, 0.8, 
    0.74, 0.74, 0.76, 0.75, 0.73, 0.68, 0.66, 0.69, 0.69, 0.67, 0.65, 0.67, 
    0.67, 0.69, 0.69, 0.68, 0.74, 0.73, 0.73, 0.77, 0.79, 0.82, 0.81, 0.87, 
    0.82, 0.86, 0.79, 0.83, 0.82, 0.77, 0.75, 0.8, 0.74, 0.7, 0.66, 0.64, 
    0.63, 0.63, 0.63, 0.67, 0.66, 0.76, 0.73, 0.78, 0.78, 0.74, 0.72, 0.72, 
    0.7, 0.7, 0.74, 0.74, 0.7, 0.7, 0.72, 0.74, 0.73, 0.71, 0.7, 0.78, 0.78, 
    0.8, 0.75, 0.78, 0.8, 0.8, 0.75, 0.76, 0.8, 0.8, 0.8, 0.84, 0.78, 0.84, 
    0.77, 0.78, 0.77, 0.78, 0.76, 0.8, 0.75, 0.79, 0.85, 0.84, 0.86, 0.86, 
    0.87, 0.86, 0.84, 0.86, 0.9, 0.92, 0.94, 0.94, 0.94, 0.93, 0.94, 0.91, 
    0.89, 0.89, 0.87, 0.85, 0.85, 0.75, 0.7, 0.69, 0.65, 0.69, 0.65, 0.68, 
    0.68, 0.71, 0.72, 0.73, 0.82, 0.78, 0.77, 0.82, 0.9, 0.86, 0.9, 0.88, 
    0.88, 0.86, 0.87, 0.83, 0.83, 0.8, 0.79, 0.75, 0.75, 0.72, 0.72, 0.7, 
    0.66, 0.63, 0.61, 0.61, 0.54, 0.56, 0.54, 0.59, 0.55, 0.53, 0.57, 0.48, 
    0.57, 0.53, 0.51, 0.56, 0.58, 0.57, 0.57, 0.57, 0.61, 0.56, 0.61, 0.57, 
    0.57, 0.61, 0.61, 0.59, 0.64, 0.64, 0.65, 0.61, 0.61, 0.6, 0.57, 0.53, 
    0.55, 0.54, 0.52, 0.53, 0.54, 0.57, 0.55, 0.51, 0.54, 0.54, 0.53, 0.5, 
    0.57, 0.54, 0.58, 0.57, 0.61, 0.6, 0.62, 0.65, 0.65, 0.65, 0.66, 0.63, 
    0.67, 0.67, 0.66, 0.68, 0.66, 0.65, 0.63, 0.63, 0.63, 0.61, 0.62, 0.62, 
    0.63, 0.62, 0.63, 0.63, 0.63, 0.64, 0.64, 0.63, 0.65, 0.66, 0.69, 0.71, 
    0.71, 0.7, 0.69, 0.68, 0.63, 0.59, 0.57, 0.57, 0.55, 0.53, 0.53, 0.54, 
    0.55, 0.53, 0.51, 0.51, 0.48, 0.51, 0.55, 0.56, 0.6, 0.62, 0.59, 0.65, 
    0.64, 0.65, 0.67, 0.64, 0.74, 0.75, 0.7, 0.74, 0.73, 0.71, 0.69, 0.65, 
    0.68, 0.67, 0.72, 0.66, 0.69, 0.69, 0.72, 0.82, 0.84, 0.88, 0.8, 0.68, 
    0.65, 0.64, 0.59, 0.55, 0.52, 0.55, 0.52, 0.49, 0.48, 0.47, 0.53, 0.53, 
    0.56, 0.6, 0.61, 0.59, 0.59, 0.62, 0.62, 0.63, 0.65, 0.65, 0.65, 0.65, 
    0.63, 0.61, 0.62, 0.63, 0.61, 0.64, 0.6, 0.59, 0.6, 0.57, 0.59, 0.59, 
    0.58, 0.61, 0.59, 0.6, 0.66, 0.64, 0.7, 0.76, 0.7, 0.75, 0.74, 0.73, 
    0.71, 0.78, 0.76, 0.86, 0.77, 0.7, 0.65, 0.64, 0.66, 0.71, 0.7, 0.71, 
    0.75, 0.73, 0.73, 0.7, 0.68, 0.66, 0.7, 0.71, 0.68, 0.64, 0.62, 0.49, 
    0.59, 0.51, 0.54, 0.58, 0.54, 0.52, 0.53, 0.52, 0.52, 0.55, 0.57, 0.57, 
    0.6, 0.58, 0.6, 0.57, 0.59, 0.59, 0.58, 0.64, 0.6, 0.61, 0.67, 0.62, 
    0.61, 0.62, 0.61, 0.56, 0.62, 0.6, 0.59, 0.61, 0.62, 0.62, 0.66, 0.69, 
    0.66, 0.73, 0.74, 0.67, 0.79, 0.72, 0.71, 0.69, 0.7, 0.7, 0.72, 0.71, 
    0.68, 0.72, 0.72, 0.65, 0.65, 0.65, 0.65, 0.69, 0.57, 0.58, 0.62, 0.66, 
    0.72, 0.59, 0.59, 0.56, 0.6, 0.66, 0.67, 0.67, 0.73, 0.76, 0.68, 0.66, 
    0.69, 0.66, 0.65, 0.66, 0.62, 0.62, 0.56, 0.56, 0.55, 0.52, 0.58, 0.55, 
    0.52, 0.4, 0.52, 0.55, 0.59, 0.62, 0.61, 0.61, 0.51, 0.55, 0.51, 0.55, 
    0.52, 0.67, 0.65, 0.55, 0.42, 0.58, 0.54, 0.53, 0.54, 0.58, 0.58, 0.58, 
    0.62, 0.61, 0.63, 0.65, 0.66, 0.7, 0.71, 0.7, 0.74, 0.7, 0.71, 0.68, 
    0.68, 0.64, 0.6, 0.66, 0.73, 0.72, 0.77, 0.68, 0.68, 0.73, 0.73, 0.72, 
    0.74, 0.74, 0.75, 0.71, 0.68, 0.69, 0.68, 0.7, 0.67, 0.76, 0.75, 0.72, 
    0.76, 0.7, 0.76, 0.73, 0.74, 0.8, 0.72, 0.77, 0.77, 0.75, 0.74, 0.76, 
    0.75, 0.73, 0.76, 0.81, 0.85, 0.86, 0.82, 0.83, 0.78, 0.8, 0.83, 0.8, 
    0.82, 0.78, 0.68, 0.72, 0.78, 0.78, 0.74, 0.75, 0.75, 0.76, 0.83, 0.82, 
    0.82, 0.77, 0.72, 0.77, 0.86, 0.87, 0.91, 0.89, 0.91, 0.88, 0.86, 0.84, 
    0.81, 0.81, 0.81, 0.68, 0.64, 0.62, 0.6, 0.6, 0.62, 0.59, 0.63, 0.65, 
    0.63, 0.64, 0.63, 0.66, 0.65, 0.65, 0.67, 0.64, 0.66, 0.66, 0.71, 0.68, 
    0.67, 0.79, 0.74, 0.72, 0.74, 0.72, 0.74, 0.71, 0.7, 0.7, 0.73, 0.76, 
    0.73, 0.75, 0.76, 0.77, 0.78, 0.79, 0.8, 0.8, 0.83, 0.84, 0.82, 0.79, 
    0.78, 0.84, 0.79, 0.76, 0.76, 0.75, 0.73, 0.71, 0.71, 0.71, 0.71, 0.72, 
    0.75, 0.76, 0.76, 0.82, 0.85, 0.85, 0.87, 0.9, 0.92, 0.91, 0.91, 0.87, 
    0.85, 0.86, 0.85, 0.84, 0.8, 0.76, 0.8, 0.65, 0.65, 0.63, 0.67, 0.72, 
    0.71, 0.76, 0.74, 0.76, 0.77, 0.73, 0.76, 0.71, 0.72, 0.76, 0.79, 0.81, 
    0.81, 0.83, 0.82, 0.81, 0.82, 0.8, 0.79, 0.8, 0.79, 0.84, 0.77, 0.78, 
    0.83, 0.84, 0.84, 0.83, 0.8, 0.78, 0.81, 0.87, 0.82, 0.81, 0.77, 0.8, 
    0.77, 0.78, 0.7, 0.71, 0.72, 0.77, 0.78, 0.78, 0.77, 0.77, 0.77, 0.77, 
    0.78, 0.8, 0.83, 0.83, 0.83, 0.82, 0.91, 0.88, 0.9, 0.82, 0.73, 0.81, 
    0.82, 0.75, 0.72, 0.8, 0.78, 0.81, 0.77, 0.8, 0.84, 0.84, 0.85, 0.85, 
    0.8, 0.81, 0.78, 0.78, 0.79, 0.71, 0.74, 0.78, 0.78, 0.78, 0.76, 0.75, 
    0.74, 0.74, 0.82, 0.8, 0.8, 0.78, 0.77, 0.73, 0.77, 0.74, 0.75, 0.78, 
    0.79, 0.81, 0.79, 0.77, 0.77, 0.85, 0.85, 0.85, 0.93, 0.94, 0.95, 0.95, 
    0.95, 0.93, 0.91, 0.9, 0.86, 0.92, 0.92, 0.83, 0.87, 0.87, 0.88, 0.91, 
    0.9, 0.91, 0.88, 0.91, 0.9, 0.9, 0.91, 0.91, 0.89, 0.89, 0.77, 0.78, 
    0.79, 0.77, 0.73, 0.79, 0.78, 0.76, 0.72, 0.71, 0.69, 0.63, 0.62, 0.69, 
    0.73, 0.72, 0.72, 0.69, 0.68, 0.73, 0.69, 0.7, 0.7, 0.72, 0.73, 0.76, 
    0.77, 0.79, 0.86, 0.85, 0.86, 0.87, 0.77, 0.74, 0.63, 0.66, 0.75, 0.74, 
    0.75, 0.72, 0.66, 0.75, 0.78, 0.67, 0.67, 0.66, 0.66, 0.68, 0.85, 0.86, 
    0.83, 0.82, 0.82, 0.82, 0.83, 0.83, 0.8, 0.76, 0.76, 0.76, 0.77, 0.84, 
    0.84, 0.85, 0.88, 0.88, 0.89, 0.87, 0.86, 0.87, 0.83, 0.82, 0.82, 0.79, 
    0.79, 0.79, 0.77, 0.75, 0.76, 0.8, 0.77, 0.77, 0.75, 0.7, 0.68, 0.66, 
    0.63, 0.64, 0.61, 0.62, 0.68, 0.69, 0.75, 0.8, 0.76, 0.75, 0.67, 0.67, 
    0.66, 0.65, 0.61, 0.5, 0.48, 0.47, 0.43, 0.43, 0.39, 0.38, 0.35, 0.39, 
    0.39, 0.44, 0.54, 0.58, 0.64, 0.68, 0.71, 0.73, 0.74, 0.77, 0.65, 0.63, 
    0.69, 0.68, 0.61, 0.59, 0.55, 0.54, 0.57, 0.56, 0.6, 0.58, 0.6, 0.6, 
    0.59, 0.62, 0.62, 0.67, 0.76, 0.72, 0.76, 0.82, 0.75, 0.73, 0.87, 0.86, 
    0.8, 0.74, 0.72, 0.8, 0.83, 0.76, 0.78, 0.79, 0.72, 0.69, 0.7, 0.74, 
    0.71, 0.67, 0.68, 0.67, 0.71, 0.78, 0.88, 0.85, 0.8, 0.79, 0.75, 0.74, 
    0.73, 0.72, 0.71, 0.72, 0.69, 0.71, 0.74, 0.7, 0.73, 0.7, 0.68, 0.7, 
    0.73, 0.69, 0.64, 0.68, 0.71, 0.69, 0.7, 0.73, 0.75, 0.76, 0.67, 0.66, 
    0.65, 0.62, 0.71, 0.72, 0.74, 0.73, 0.69, 0.67, 0.74, 0.63, 0.59, 0.49, 
    0.49, 0.48, 0.5, 0.48, 0.53, 0.56, 0.55, 0.51, 0.59, 0.55, 0.58, 0.56, 
    0.52, 0.49, 0.47, 0.45, 0.48, 0.5, 0.55, 0.51, 0.57, 0.59, 0.57, 0.54, 
    0.47, 0.58, 0.55, 0.6, 0.6, 0.61, 0.58, 0.55, 0.54, 0.51, 0.49, 0.54, 
    0.61, 0.65, 0.46, 0.46, 0.49, 0.53, 0.53, 0.48, 0.54, 0.53, 0.48, 0.43, 
    0.51, 0.45, 0.52, 0.51, 0.54, 0.49, 0.61, 0.57, 0.56, 0.57, 0.51, 0.54, 
    0.51, 0.55, 0.45, 0.47, 0.46, 0.54, 0.48, 0.42, 0.44, 0.42, 0.44, 0.5, 
    0.45, 0.45, 0.44, 0.48, 0.5, 0.52, 0.57, 0.64, 0.58, 0.44, 0.53, 0.44, 
    0.48, 0.46, 0.42, 0.38, 0.48, 0.55, 0.42, 0.46, 0.51, 0.45, 0.49, 0.49, 
    0.51, 0.54, 0.53, 0.56, 0.64, 0.59, 0.58, 0.59, 0.7, 0.75, 0.82, 0.81, 
    0.79, 0.79, 0.74, 0.72, 0.71, 0.64, 0.66, 0.68, 0.67, 0.67, 0.69, 0.71, 
    0.68, 0.69, 0.71, 0.73, 0.75, 0.72, 0.72, 0.77, 0.73, 0.72, 0.73, 0.72, 
    0.69, 0.74, 0.7, 0.68, 0.7, 0.68, 0.66, 0.71, 0.74, 0.69, 0.77, 0.77, 
    0.78, 0.81, 0.76, 0.81, 0.82, 0.74, 0.88, 0.87, 0.87, 0.91, 0.92, 0.92, 
    0.93, 0.94, 0.94, 0.93, 0.93, 0.95, 0.95, 0.9, 0.91, 0.91, 0.9, 0.89, 
    0.89, 0.87, 0.86, 0.9, 0.91, 0.91, 0.91, 0.92, 0.91, 0.9, 0.89, 0.81, 
    0.87, 0.83, 0.82, 0.79, 0.76, 0.74, 0.72, 0.69, 0.65, 0.64, 0.61, 0.63, 
    0.67, 0.75, 0.8, 0.82, 0.82, 0.83, 0.81, 0.83, 0.82, 0.84, 0.85, 0.81, 
    0.87, 0.86, 0.83, 0.8, 0.77, 0.81, 0.8, 0.83, 0.83, 0.81, 0.82, 0.82, 
    0.85, 0.83, 0.91, 0.93, 0.9, 0.88, 0.87, 0.85, 0.85, 0.85, 0.86, 0.86, 
    0.82, 0.85, 0.83, 0.86, 0.85, 0.83, 0.83, 0.86, 0.88, 0.93, 0.93, 0.93, 
    0.92, 0.91, 0.9, 0.91, 0.92, 0.92, 0.94, 0.92, 0.92, 0.94, 0.94, 0.95, 
    0.96, 0.95, 0.94, 0.91, 0.89, 0.88, 0.88, 0.85, 0.87, 0.85, 0.85, 0.85, 
    0.82, 0.86, 0.78, 0.76, 0.75, 0.78, 0.8, 0.79, 0.75, 0.77, 0.75, 0.75, 
    0.76, 0.74, 0.79, 0.76, 0.77, 0.78, 0.77, 0.75, 0.73, 0.73, 0.73, 0.67, 
    0.67, 0.66, 0.65, 0.66, 0.62, 0.62, 0.64, 0.66, 0.64, 0.71, 0.72, 0.65, 
    0.62, 0.65, 0.67, 0.68, 0.72, 0.75, 0.72, 0.85, 0.72, 0.76, 0.74, 0.72, 
    0.69, 0.71, 0.77, 0.71, 0.73, 0.72, 0.82, 0.83, 0.8, 0.77, 0.77, 0.79, 
    0.81, 0.84, 0.81, 0.81, 0.77, 0.82, 0.87, 0.93, 0.95, 0.94, 0.93, 0.93, 
    0.92, 0.89, 0.89, 0.89, 0.89, 0.87, 0.87, 0.82, 0.81, 0.85, 0.88, 0.83, 
    0.76, 0.78, 0.7, 0.68, 0.67, 0.69, 0.71, 0.69, 0.74, 0.78, 0.77, 0.78, 
    0.75, 0.76, 0.76, 0.77, 0.77, 0.79, 0.82, 0.83, 0.85, 0.86, 0.87, 0.9, 
    0.93, 0.88, 0.87, 0.86, 0.83, 0.8, 0.83, 0.72, 0.73, 0.71, 0.71, 0.7, 
    0.7, 0.71, 0.8, 0.8, 0.81, 0.73, 0.76, 0.82, 0.86, 0.92, 0.91, 0.85, 
    0.87, 0.85, 0.75, 0.8, 0.76, 0.76, 0.75, 0.75, 0.74, 0.74, 0.75, 0.82, 
    0.85, 0.83, 0.77, 0.79, 0.84, 0.83, 0.81, 0.9, 0.89, 0.93, 0.92, 0.92, 
    0.93, 0.92, 0.89, 0.85, 0.83, 0.86, 0.84, 0.78, 0.83, 0.8, 0.81, 0.81, 
    0.82, 0.81, 0.78, 0.8, 0.89, 0.77, 0.74, 0.71, 0.7, 0.78, 0.63, 0.69, 
    0.65, 0.58, 0.6, 0.66, 0.62, 0.65, 0.63, 0.63, 0.65, 0.63, 0.61, 0.66, 
    0.7, 0.66, 0.68, 0.7, 0.7, 0.68, 0.7, 0.72, 0.73, 0.68, 0.73, 0.73, 0.73, 
    0.74, 0.7, 0.69, 0.75, 0.68, 0.7, 0.71, 0.72, 0.74, 0.74, 0.73, 0.69, 
    0.71, 0.71, 0.72, 0.73, 0.77, 0.76, 0.79, 0.79, 0.84, 0.91, 0.84, 0.81, 
    0.8, 0.75, 0.75, 0.75, 0.71, 0.75, 0.74, 0.74, 0.7, 0.71, 0.71, 0.71, 
    0.7, 0.62, 0.67, 0.71, 0.74, 0.78, 0.78, 0.8, 0.79, 0.77, 0.8, 0.71, 
    0.64, 0.64, 0.65, 0.64, 0.64, 0.65, 0.64, 0.66, 0.63, 0.64, 0.63, 0.65, 
    0.69, 0.73, 0.78, 0.78, 0.83, 0.82, 0.82, 0.81, 0.85, 0.87, 0.89, 0.85, 
    0.85, 0.85, 0.83, 0.8, 0.77, 0.78, 0.75, 0.73, 0.74, 0.76, 0.77, 0.75, 
    0.75, 0.7, 0.71, 0.68, 0.69, 0.7, 0.69, 0.71, 0.68, 0.7, 0.68, 0.69, 
    0.68, 0.69, 0.67, 0.61, 0.59, 0.59, 0.64, 0.62, 0.61, 0.62, 0.68, 0.68, 
    0.67, 0.68, 0.67, 0.64, 0.68, 0.71, 0.68, 0.7, 0.69, 0.67, 0.67, 0.66, 
    0.66, 0.65, 0.63, 0.6, 0.62, 0.64, 0.69, 0.66, 0.72, 0.71, 0.73, 0.75, 
    0.72, 0.71, 0.71, 0.7, 0.75, 0.77, 0.77, 0.77, 0.69, 0.71, 0.7, 0.68, 
    0.69, 0.68, 0.68, 0.69, 0.72, 0.74, 0.69, 0.72, 0.7, 0.71, 0.72, 0.72, 
    0.71, 0.75, 0.78, 0.79, 0.81, 0.79, 0.8, 0.79, 0.79, 0.79, 0.76, 0.74, 
    0.67, 0.71, 0.72, 0.65, 0.61, 0.61, 0.64, 0.62, 0.67, 0.68, 0.57, 0.52, 
    0.55, 0.57, 0.7, 0.79, 0.77, 0.72, 0.71, 0.74, 0.8, 0.81, 0.73, 0.79, 
    0.71, 0.7, 0.69, 0.67, 0.65, 0.66, 0.75, 0.79, 0.62, 0.59, 0.6, 0.63, 
    0.67, 0.69, 0.69, 0.71, 0.7, 0.72, 0.73, 0.73, 0.72, 0.74, 0.75, 0.71, 
    0.72, 0.69, 0.67, 0.73, 0.66, 0.64, 0.69, 0.64, 0.68, 0.65, 0.63, 0.62, 
    0.66, 0.68, 0.7, 0.7, 0.75, 0.76, 0.75, 0.76, 0.75, 0.74, 0.75, 0.72, 
    0.72, 0.73, 0.72, 0.73, 0.75, 0.76, 0.75, 0.74, 0.74, 0.75, 0.74, 0.74, 
    0.72, 0.71, 0.67, 0.7, 0.73, 0.69, 0.7, 0.7, 0.7, 0.71, 0.68, 0.7, 0.71, 
    0.66, 0.67, 0.65, 0.63, 0.66, 0.64, 0.65, 0.66, 0.74, 0.74, 0.76, 0.76, 
    0.81, 0.8, 0.84, 0.81, 0.88, 0.89, 0.87, 0.82, 0.84, 1, 0.85, 0.85, 0.84, 
    0.84, 0.86, 0.89, 0.9, 0.9, 0.88, 0.85, 0.85, 0.86, 0.87, 0.87, 0.87, 
    0.88, 0.9, 0.91, 0.92, 0.95, 0.94, 1, 1, 0.96, 0.95, 0.91, 0.77, 0.78, 
    0.77, 0.76, 0.74, 0.74, 0.73, 0.74, 0.72, 0.69, 0.66, 0.69, 0.66, 0.67, 
    0.62, 0.67, 0.7, 0.69, 0.71, 0.7, 0.67, 0.69, 0.66, 0.67, 0.66, 0.61, 
    0.62, 0.58, 0.62, 0.62, 0.6, 0.61, 0.6, 0.6, 0.61, 0.63, 0.61, 0.64, 
    0.66, 0.7, 0.73, 0.73, 0.72, 0.7, 0.9, 0.71, 0.65, 0.63, 0.61, 0.63, 0.6, 
    0.61, 0.63, 0.63, 0.61, 0.58, 0.59, 0.56, 0.58, 0.58, 0.59, 0.6, 0.62, 
    0.62, 0.63, 0.63, 0.86, 0.9, 0.68, 0.66, 0.63, 0.63, 0.61, 0.63, 0.65, 
    0.67, 0.66, 0.65, 0.63, 0.58, 0.63, 0.65, 0.7, 0.72, 0.71, 0.71, 0.73, 
    0.75, 0.75, 0.74, 0.74, 0.77, 0.73, 0.77, 0.76, 0.76, 0.78, 0.87, 0.9, 
    0.93, 0.85, 0.85, 0.85, 0.87, 0.87, 0.82, 0.81, 0.89, 0.87, 0.86, 0.91, 
    0.92, 0.93, 0.93, 0.91, 0.91, 0.91, 0.88, 0.83, 0.65, 0.7, 0.65, 0.66, 
    0.66, 0.66, 0.7, 0.64, 0.69, 0.68, 0.62, 0.64, 0.7, 0.74, 0.78, 0.74, 
    0.77, 0.79, 0.82, 0.84, 0.85, 0.9, 0.79, 0.77, 0.78, 0.79, 0.69, 0.77, 
    0.79, 0.72, 0.71, 0.73, 0.74, 0.76, 0.78, 0.85, 0.84, 0.79, 0.77, 1, 
    0.79, 1, 0.75, 0.73, 0.71, 0.67, 0.67, 0.68, 0.63, 0.61, 0.62, 0.6, 0.62, 
    0.64, 0.62, 0.65, 0.64, 0.7, 0.74, 0.74, 0.72, 0.78, 0.81, 0.79, 0.82, 
    0.82, 0.91, 0.93, 0.94, 0.95, 0.93, 0.94, 0.93, 0.92, 0.87, 0.87, 0.84, 
    0.81, 0.81, 0.81, 0.81, 0.83, 0.81, 0.84, 0.82, 0.84, 0.81, 0.85, 0.84, 
    0.86, 0.89, 0.91, 0.9, 0.9, 0.89, 0.86, 0.83, 0.79, 0.75, 0.86, 0.84, 
    0.89, 0.88, 0.9, 0.94, 0.96, 0.96, 0.92, 1, 0.9, 0.89, 0.88, 0.86, 0.85, 
    0.84, 0.84, 0.84, 0.75, 0.77, 0.78, 0.83, 0.85, 0.81, 0.8, 0.83, 0.87, 
    0.92, 0.94, 0.94, 0.94, 0.94, 0.86, 1, 0.86, 0.83, 0.81, 0.86, 0.86, 
    0.88, 0.86, 0.85, 0.86, 0.89, 0.9, 0.88, 0.9, 0.89, 0.85, 0.84, 0.85, 
    0.88, 0.86, 0.86, 0.86, 0.81, 0.82, 0.82, 0.86, 0.85, 0.81, 0.82, 0.81, 
    0.82, 0.83, 0.8, 0.86, 0.89, 0.91, 0.93, 0.91, 0.89, 0.89, 0.88, 0.88, 
    0.89, 0.89, 0.9, 0.9, 0.91, 0.88, 0.89, 0.8, 0.91, 0.9, 0.81, 0.83, 0.77, 
    0.8, 0.78, 0.79, 0.78, 0.78, 0.79, 0.8, 0.79, 0.78, 0.78, 0.71, 0.68, 
    0.68, 0.66, 0.63, 0.58, 0.55, 0.61, 0.62, 0.65, 0.67, 0.65, 0.66, 0.66, 
    0.67, 0.69, 0.7, 0.69, 0.7, 0.73, 0.72, 0.71, 0.81, 0.75, 0.73, 0.73, 
    0.7, 0.63, 0.57, 0.59, 0.63, 0.62, 0.66, 0.67, 0.67, 0.67, 0.64, 0.7, 
    0.65, 0.69, 0.48, 0.48, 0.42, 0.48, 0.52, 0.51, 0.49, 0.48, 0.46, 0.46, 
    0.46, 0.46, 0.43, 0.44, 0.47, 0.49, 0.5, 0.59, 0.62, 0.59, 0.61, 0.71, 
    0.66, 0.68, 0.68, 0.64, 0.6, 0.57, 0.62, 0.62, 0.59, 0.58, 0.65, 0.62, 
    0.64, 0.64, 0.62, 0.67, 0.72, 0.76, 0.78, 0.9, 0.95, 0.94, 0.95, 0.95, 
    0.96, 0.87, 0.84, 0.82, 0.69, 0.65, 0.59, 0.59, 0.59, 0.6, 0.56, 0.57, 
    0.65, 0.61, 0.65, 0.64, 0.58, 0.57, 0.61, 0.65, 0.61, 0.66, 0.66, 0.68, 
    0.62, 0.68, 0.62, 0.64, 0.6, 0.59, 0.61, 0.6, 0.6, 0.54, 0.52, 0.58, 
    0.63, 0.6, 0.55, 0.54, 0.53, 0.59, 0.64, 0.68, 0.68, 0.68, 0.71, 0.74, 
    0.77, 0.73, 0.78, 0.72, 0.72, 0.68, 0.7, 0.65, 0.62, 0.66, 0.67, 0.68, 
    0.69, 0.68, 0.72, 0.71, 0.73, 0.76, 0.79, 0.81, 0.82, 0.68, 0.53, 0.61, 
    0.66, 0.71, 0.72, 0.68, 0.73, 0.67, 0.75, 0.7, 0.64, 0.61, 0.61, 0.6, 
    0.6, 0.58, 0.59, 0.61, 0.62, 0.62, 0.71, 0.73, 0.72, 0.66, 0.64, 0.68, 
    0.68, 0.67, 0.7, 0.77, 0.7, 0.67, 0.61, 0.59, 0.71, 0.59, 0.59, 0.64, 
    0.64, 0.64, 0.71, 0.79, 0.78, 0.74, 0.73, 0.76, 0.72, 0.71, 0.7, 0.67, 
    0.64, 0.66, 0.67, 0.62, 0.65, 0.63, 0.62, 0.61, 0.61, 0.61, 0.61, 0.62, 
    0.61, 0.61, 0.62, 0.63, 0.63, 0.67, 0.68, 0.72, 0.7, 0.72, 0.75, 0.83, 
    0.82, 0.83, 0.81, 0.84, 0.76, 0.72, 0.81, 0.78, 0.75, 0.72, 0.7, 0.66, 
    0.67, 0.64, 0.62, 0.64, 0.59, 0.59, 0.64, 0.65, 0.66, 0.67, 0.72, 0.75, 
    0.78, 0.78, 0.76, 0.74, 0.7, 0.6, 0.59, 0.58, 0.57, 0.55, 0.56, 0.55, 
    0.55, 0.56, 0.57, 0.6, 0.66, 0.64, 0.68, 0.73, 0.78, 0.83, 0.87, 0.87, 
    0.88, 0.86, 0.88, 0.79, 0.78, 0.74, 0.69, 0.65, 0.56, 0.54, 0.56, 0.57, 
    0.55, 0.54, 0.59, 0.59, 0.63, 0.63, 0.67, 0.67, 0.66, 0.66, 0.69, 0.69, 
    0.71, 0.64, 0.65, 0.62, 0.59, 0.56, 0.55, 0.55, 0.52, 0.59, 0.56, 0.53, 
    0.55, 0.55, 0.53, 0.54, 0.55, 0.54, 0.55, 0.57, 0.64, 0.61, 0.64, 0.67, 
    0.7, 0.72, 0.72, 0.73, 0.75, 0.73, 0.7, 0.67, 0.71, 0.71, 0.73, 0.75, 
    0.7, 0.76, 0.75, 0.77, 0.82, 0.83, 0.85, 0.8, 0.76, 0.79, 0.87, 0.79, 
    0.82, 0.87, 0.86, 0.85, 0.75, 0.79, 0.75, 0.76, 0.77, 0.76, 0.77, 0.77, 
    0.77, 0.8, 0.85, 0.83, 0.79, 0.83, 0.85, 0.86, 0.83, 0.85, 0.85, 0.87, 
    0.85, 0.87, 0.89, 0.89, 0.87, 0.86, 0.83, 0.79, 0.73, 0.77, 0.78, 0.73, 
    0.74, 0.77, 0.77, 0.77, 0.76, 0.8, 0.83, 0.8, 0.83, 0.81, 0.79, 0.81, 
    0.85, 0.83, 0.85, 0.81, 0.78, 0.8, 0.79, 0.78, 0.81, 0.8, 0.8, 0.81, 0.8, 
    0.81, 0.85, 0.85, 0.83, 0.87, 0.89, 0.9, 0.87, 0.89, 0.88, 0.89, 0.91, 
    0.9, 0.88, 0.89, 0.88, 0.88, 0.84, 0.82, 0.82, 0.83, 0.81, 0.79, 0.78, 
    0.81, 0.83, 0.84, 0.86, 0.89, 0.89, 0.9, 0.88, 0.86, 0.81, 0.86, 0.85, 
    0.84, 0.83, 0.83, 0.83, 0.73, 0.69, 0.7, 0.73, 0.7, 0.75, 0.73, 0.73, 
    0.74, 0.79, 0.73, 0.78, 0.79, 0.82, 0.82, 0.81, 0.85, 0.81, 0.85, 0.87, 
    0.82, 0.84, 0.84, 0.78, 0.79, 0.77, 0.72, 0.77, 0.75, 0.78, 0.78, 0.77, 
    0.74, 0.78, 0.78, 0.79, 0.83, 0.77, 0.75, 0.86, 0.82, 0.82, 0.82, 0.75, 
    0.75, 0.67, 0.7, 0.66, 0.66, 0.7, 0.65, 0.69, 0.67, 0.6, 0.68, 0.76, 
    0.77, 0.78, 0.72, 0.69, 0.72, 0.73, 0.65, 0.67, 0.69, 0.71, 0.64, 0.63, 
    0.73, 0.67, 0.69, 0.62, 0.68, 0.64, 0.69, 0.66, 0.7, 0.72, 0.71, 0.68, 
    0.74, 0.76, 0.71, 0.8, 0.73, 0.79, 0.79, 0.76, 0.85, 0.84, 0.73, 0.76, 
    0.79, 0.81, 0.82, 0.82, 0.8, 0.78, 0.82, 0.79, 0.81, 0.81, 0.78, 0.8, 
    0.88, 0.88, 0.88, 0.92, 0.86, 0.83, 0.73, 0.8, 0.84, 0.81, 0.82, 0.83, 
    0.8, 0.85, 0.85, 0.84, 0.84, 0.83, 0.8, 0.77, 0.84, 0.87, 0.93, 0.93, 
    0.84, 0.87, 0.86, 0.88, 0.9, 0.83, 0.81, 0.76, 0.76, 0.77, 0.79, 0.78, 
    0.73, 0.76, 0.72, 0.73, 0.71, 0.72, 0.71, 0.69, 0.74, 0.68, 0.77, 0.71, 
    0.74, 0.7, 0.73, 0.73, 0.76, 0.74, 0.71, 0.68, 0.72, 0.8, 0.79, 0.81, 
    0.87, 0.85, 0.81, 0.87, 0.87, 0.79, 0.86, 0.85, 0.8, 0.78, 0.77, 0.7, 
    0.72, 0.74, 0.77, 0.82, 0.86, 0.9, 0.91, 0.9, 0.89, 0.87, 0.86, 0.88, 
    0.91, 0.93, 0.94, 0.92, 0.89, 0.85, 0.81, 0.79, 0.88, 0.88, 0.89, 0.89, 
    0.88, 0.77, 0.79, 0.72, 0.76, 0.77, 0.74, 0.78, 0.78, 0.82, 0.83, 0.86, 
    0.87, 0.92, 0.9, 0.91, 0.91, 0.89, 0.93, 0.94, 0.86, 0.72, 0.74, 0.82, 
    0.68, 0.69, 0.73, 0.8, 0.87, 0.8, 0.77, 0.76, 0.78, 0.81, 0.78, 0.73, 
    0.75, 0.75, 0.76, 0.8, 0.8, 0.79, 0.81, 0.8, 0.77, 0.77, 0.84, 0.82, 
    0.81, 0.79, 0.81, 0.8, 0.8, 0.79, 0.77, 0.78, 0.83, 0.83, 0.86, 0.84, 
    0.86, 0.86, 0.82, 0.82, 0.82, 0.81, 0.8, 0.85, 0.83, 0.85, 0.86, 0.87, 
    0.91, 0.92, 0.94, 0.95, 0.95, 0.95, 0.95, 0.94, 0.92, 0.91, 0.9, 0.92, 
    0.86, 0.8, 0.76, 0.84, 0.86, 0.77, 0.76, 0.78, 0.8, 0.74, 0.78, 0.85, 
    0.84, 0.82, 0.83, 0.8, 0.84, 0.83, 0.81, 0.85, 0.87, 0.82, 0.85, 0.87, 
    0.89, 0.89, 0.91, 0.92, 0.85, 0.9, 0.92, 0.79, 0.74, 0.72, 0.71, 0.69, 
    0.72, 0.75, 0.73, 0.74, 0.73, 0.73, 0.73, 0.71, 0.71, 0.72, 0.75, 0.77, 
    0.81, 0.82, 0.78, 0.79, 0.77, 0.75, 0.69, 0.64, 0.77, 0.83, 0.85, 0.84, 
    0.91, 0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.97, 0.98, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 1, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.99, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.98, 0.99, 0.99, 0.99, 0.99, 0.98, 0.99, 0.98, 0.98, 0.99, 0.98, 
    0.98, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 0.98, 0.98, 0.98, 0.94, 0.94, 
    0.95, 0.91, 0.83, 0.75, 0.73, 0.76, 0.77, 0.74, 0.77, 0.82, 0.87, 0.91, 
    0.9, 0.91, 0.94, 0.9, 0.93, 0.95, 0.96, 0.96, 0.97, 0.97, 0.97, 0.96, 
    0.96, 0.95, 0.95, 0.9, 0.93, 0.95, 0.97, 0.98, 0.98, 0.97, 0.98, 0.98, 
    0.98, 0.96, 0.96, 0.96, 0.94, 0.92, 0.9, 0.89, 0.91, 0.92, 0.86, 0.91, 
    0.91, 0.92, 0.92, 0.9, 0.82, 0.87, 0.9, 0.89, 0.88, 0.9, 0.88, 0.8, 0.72, 
    0.71, 0.66, 0.66, 0.62, 0.64, 0.61, 0.62, 0.61, 0.62, 0.6, 0.56, 0.56, 
    0.55, 0.52, 0.52, 0.51, 0.52, 0.53, 0.51, 0.52, 0.53, 0.54, 0.53, 0.53, 
    0.56, 0.59, 0.58, 0.59, 0.55, 0.57, 0.58, 0.59, 0.6, 0.66, 0.65, 0.62, 
    0.63, 0.64, 0.64, 0.64, 0.63, 0.62, 0.63, 0.65, 0.67, 0.65, 0.64, 0.68, 
    0.65, 0.66, 0.68, 0.7, 0.67, 0.63, 0.62, 0.64, 0.63, 0.66, 0.7, 0.68, 
    0.66, 0.68, 0.7, 0.72, 0.72, 0.71, 0.69, 0.76, 0.77, 0.77, 0.78, 0.76, 
    0.76, 0.8, 0.85, 0.84, 0.86, 0.84, 0.83, 0.87, 0.89, 0.85, 0.86, 0.87, 
    0.91, 0.92, 0.91, 0.9, 0.9, 0.87, 0.85, 0.82, 0.81, 0.8, 0.78, 0.73, 0.7, 
    0.65, 0.64, 0.58, 0.56, 0.57, 0.6, 0.65, 0.64, 0.64, 0.87, 0.8, 0.66, 
    0.75, 0.7, 0.62, 0.6, 0.62, 0.63, 0.64, 0.65, 0.63, 0.66, 0.69, 0.73, 
    0.71, 0.72, 0.74, 0.76, 0.75, 0.82, 0.89, 0.91, 0.89, 0.9, 0.94, 0.96, 
    0.97, 0.97, 0.93, 0.91, 0.91, 0.96, 0.96, 0.96, 0.94, 0.97, 0.96, 0.94, 
    0.94, 0.87, 0.93, 0.95, 0.96, 0.96, 0.87, 0.85, 0.86, 0.86, 0.87, 0.87, 
    0.84, 0.81, 0.84, 0.89, 0.9, 0.87, 0.89, 0.88, 0.86, 0.8, 0.78, 0.79, 
    0.78, 0.82, 0.85, 0.88, 0.86, 0.72, 0.59, 0.67, 0.76, 0.78, 0.78, 0.86, 
    0.91, 0.94, 0.96, 0.96, 0.98, 0.97, 0.96, 0.96, 0.97, 0.97, 0.89, 0.86, 
    0.84, 0.81, 0.83, 0.8, 0.82, 0.82, 0.8, 0.76, 0.76, 0.72, 0.75, 0.72, 
    0.74, 0.74, 0.64, 0.67, 0.7, 0.67, 0.69, 0.7, 0.7, 0.71, 0.71, 0.73, 
    0.76, 0.72, 0.74, 0.79, 0.79, 0.71, 0.77, 0.8, 0.76, 0.74, 0.78, 0.8, 
    0.81, 0.83, 0.87, 0.82, 0.87, 0.83, 0.82, 0.81, 0.83, 0.81, 0.85, 0.81, 
    0.83, 0.8, 0.79, 0.88, 0.95, 0.96, 0.86, 0.85, 0.87, 0.91, 0.94, 0.87, 
    0.85, 0.87, 0.9, 0.88, 0.85, 0.86, 0.86, 0.88, 0.88, 0.82, 0.86, 0.91, 
    0.86, 0.87, 0.84, 0.85, 0.88, 0.87, 0.86, 0.89, 0.85, 0.84, 0.84, 0.82, 
    0.83, 0.85, 0.83, 0.84, 0.85, 0.89, 0.9, 0.89, 0.91, 0.89, 0.88, 0.9, 
    0.88, 0.85, 0.83, 0.93, 0.94, 0.95, 0.93, 0.88, 0.85, 0.92, 0.93, 0.92, 
    0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.97, 0.97, 0.97, 
    0.97, 0.92, 0.87, 0.86, 0.85, 0.86, 0.83, 0.82, 0.81, 0.78, 0.77, 0.85, 
    0.81, 0.86, 0.82, 0.82, 0.83, 0.82, 0.83, 0.81, 0.81, 0.86, 0.85, 0.82, 
    0.8, 0.85, 0.87, 0.9, 0.92, 0.89, 0.9, 0.89, 0.91, 0.93, 0.81, 0.81, 
    0.83, 0.83, 0.83, 0.81, 0.88, 0.93, 0.92, 0.92, 0.9, 0.89, 0.9, 0.89, 
    0.92, 0.92, 0.92, 0.91, 0.94, 0.95, 0.96, 0.96, 0.93, 0.87, 0.86, 0.82, 
    0.81, 0.79, 0.8, 0.89, 0.84, 0.8, 0.79, 0.84, 0.84, 0.84, 0.85, 0.83, 
    0.82, 0.79, 0.75, 0.72, 0.66, 0.68, 0.76, 0.75, 0.59, 0.55, 0.63, 0.65, 
    0.63, 0.65, 0.63, 0.63, 0.68, 0.66, 0.62, 0.57, 0.56, 0.56, 0.56, 0.58, 
    0.57, 0.61, 0.59, 0.62, 0.64, 0.65, 0.64, 0.6, 0.64, 0.63, 0.67, 0.66, 
    0.66, 0.68, 0.69, 0.73, 0.79, 0.81, 0.87, 0.94, 0.94, 0.94, 0.92, 0.92, 
    0.92, 0.93, 0.94, 0.91, 0.89, 0.95, 0.95, 0.95, 0.96, 0.96, 0.91, 0.88, 
    0.92, 0.9, 0.89, 0.81, 0.79, 0.8, 0.81, 0.81, 0.84, 0.8, 0.84, 0.86, 
    0.87, 0.85, 0.89, 0.87, 0.86, 0.88, 0.86, 0.88, 0.86, 0.9, 0.94, 0.92, 
    0.95, 0.96, 0.97, 0.97, 0.98, 0.94, 0.89, 0.87, 0.86, 0.89, 0.88, 0.9, 
    0.9, 0.91, 0.94, 0.95, 0.95, 0.95, 0.95, 0.96, 0.95, 0.96, 0.97, 0.97, 
    0.97, 0.97, 0.96, 0.99, 0.97, 0.95, 0.96, 0.96, 0.91, 0.87, 0.91, 0.9, 
    0.87, 0.9, 0.91, 0.91, 0.92, 0.9, 0.89, 0.88, 0.91, 0.92, 0.9, 0.85, 
    0.84, 0.82, 0.82, 0.78, 0.79, 0.74, 0.71, 0.73, 0.76, 0.77, 0.79, 0.83, 
    0.83, 0.83, 0.84, 0.83, 0.86, 0.83, 0.77, 0.76, 0.77, 0.79, 0.78, 0.76, 
    0.79, 0.77, 0.78, 0.8, 0.83, 0.88, 0.86, 0.86, 0.87, 0.88, 0.86, 0.85, 
    0.77, 0.82, 0.82, 0.81, 0.81, 0.81, 0.87, 0.86, 0.9, 0.9, 0.9, 0.93, 0.9, 
    0.91, 0.92, 0.95, 0.93, 0.94, 0.94, 0.96, 0.96, 0.96, 0.96, 0.95, 0.94, 
    0.95, 0.97, 0.94, 0.85, 0.87, 0.87, 0.88, 0.89, 0.87, 0.87, 0.83, 0.83, 
    0.79, 0.8, 0.81, 0.81, 0.76, 0.71, 0.76, 0.78, 0.78, 0.76, 0.86, 0.86, 
    0.92, 0.92, 0.94, 0.94, 0.94, 0.95, 0.95, 0.94, 0.89, 0.87, 0.84, 0.84, 
    0.89, 0.88, 0.78, 0.89, 0.89, 0.88, 0.92, 0.85, 0.79, 0.78, 0.69, 0.68, 
    0.71, 0.7, 0.64, 0.64, 0.65, 0.73, 0.72, 0.75, 0.72, 0.77, 0.84, 0.83, 
    0.84, 0.86, 0.87, 0.89, 0.89, 0.9, 0.88, 0.84, 0.86, 0.85, 0.89, 0.89, 
    0.93, 0.93, 0.94, 0.89, 0.9, 0.94, 0.92, 0.92, 0.76, 0.78, 0.8, 0.68, 
    0.73, 0.81, 0.81, 0.89, 0.86, 0.83, 0.74, 0.63, 1, 0.67, 0.67, 0.7, 0.72, 
    0.71, 0.67, 0.69, 0.71, 0.73, 0.71, 0.7, 0.71, 0.69, 0.75, 0.72, 0.72, 
    0.68, 0.72, 0.73, 0.71, 0.76, 0.75, 0.73, 0.77, 0.75, 0.68, 0.66, 0.72, 
    0.69, 0.64, 0.64, 0.62, 0.65, 0.58, 0.61, 0.59, 0.61, 0.54, 0.55, 0.56, 
    0.51, 0.51, 0.56, 0.58, 0.57, 0.56, 0.52, 0.57, 0.57, 0.52, 0.52, 0.55, 
    0.55, 0.58, 0.54, 0.61, 0.59, 0.56, 0.59, 0.56, 0.54, 0.53, 0.56, 0.64, 
    0.69, 0.68, 0.68, 0.66, 0.65, 0.63, 0.6, 0.59, 0.64, 0.62, 0.63, 0.66, 
    0.68, 0.66, 0.68, 0.66, 0.66, 0.62, 0.63, 0.63, 0.75, 0.71, 0.69, 0.71, 
    0.72, 0.73, 0.83, 0.8, 0.81, 0.79, 0.8, 0.81, 0.85, 0.81, 0.81, 0.82, 
    0.85, 0.85, 0.9, 0.92, 0.92, 0.91, 0.91, 0.88, 0.85, 0.78, 0.83, 0.82, 
    0.81, 0.79, 0.78, 0.8, 0.78, 0.79, 0.81, 0.77, 0.76, 0.77, 0.8, 0.8, 
    0.81, 0.77, 0.77, 0.81, 0.8, 0.81, 0.82, 0.81, 0.76, 0.83, 0.8, 0.74, 
    0.79, 0.84, 0.86, 0.87, 0.88, 0.89, 0.87, 0.84, 0.83, 0.86, 0.82, 0.85, 
    0.85, 0.86, 0.87, 0.85, 0.83, 0.84, 0.85, 0.86, 0.85, 0.87, 0.81, 0.84, 
    0.87, 0.88, 0.86, 0.86, 0.86, 0.86, 0.85, 0.85, 0.83, 0.84, 0.82, 0.84, 
    0.84, 0.85, 0.82, 0.76, 0.82, 0.85, 0.85, 0.86, 0.84, 0.77, 0.75, 0.83, 
    0.84, 0.88, 0.82, 0.84, 0.86, 0.85, 0.85, 0.85, 0.86, 0.84, 0.87, 0.83, 
    0.81, 0.8, 0.81, 0.82, 0.78, 0.81, 0.81, 0.84, 0.85, 0.88, 0.88, 0.95, 
    0.94, 0.96, 0.96, 0.83, 0.74, 0.75, 0.76, 0.75, 0.79, 0.87, 0.87, 0.86, 
    0.86, 0.87, 0.88, 0.86, 0.83, 0.77, 0.72, 0.7, 0.71, 0.68, 0.71, 0.71, 
    0.72, 0.79, 0.75, 0.75, 0.73, 0.74, 0.8, 0.83, 0.87, 0.88, 0.88, 0.92, 
    0.91, 0.73, 0.75, 0.75, 0.8, 0.8, 0.78, 0.8, 0.83, 0.82, 0.74, 0.74, 
    0.81, 0.82, 0.87, 0.86, 0.78, 0.78, 0.76, 0.78, 0.77, 0.77, 0.81, 0.81, 
    0.8, 0.77, 0.77, 0.78, 0.85, 0.86, 0.84, 0.83, 0.84, 0.85, 0.8, 0.83, 
    0.85, 0.79, 0.76, 0.77, 0.76, 0.75, 0.76, 0.78, 0.75, 0.75, 0.79, 0.72, 
    0.68, 0.71, 0.73, 0.72, 0.72, 0.74, 0.66, 0.69, 0.7, 0.7, 0.72, 0.7, 
    0.71, 0.7, 0.74, 0.77, 0.85, 0.9, 0.91, 0.93, 0.96, 0.96, 0.96, 0.97, 
    0.97, 0.97, 0.97, 0.95, 0.91, 0.87, 0.85, 0.85, 0.84, 0.81, 0.83, 0.83, 
    0.82, 0.8, 0.77, 0.75, 0.71, 0.65, 0.7, 0.67, 0.73, 0.69, 0.68, 0.69, 
    0.67, 0.62, 0.63, 0.69, 0.63, 0.7, 0.67, 0.75, 0.75, 0.76, 0.74, 0.72, 
    0.76, 0.79, 0.81, 0.81, 0.83, 0.82, 0.71, 0.79, 0.68, 0.74, 0.69, 0.77, 
    0.71, 0.75, 0.71, 0.73, 0.76, 0.74, 0.68, 0.7, 0.73, 0.74, 0.7, 0.64, 
    0.76, 0.75, 0.73, 0.7, 0.72, 0.69, 0.7, 0.72, 0.74, 0.9, 0.93, 0.93, 
    0.92, 0.94, 0.95, 0.93, 0.85, 0.81, 0.76, 0.79, 0.76, 0.78, 0.76, 0.77, 
    0.77, 0.75, 0.75, 0.75, 0.76, 0.77, 0.77, 0.79, 0.76, 0.75, 0.79, 0.76, 
    0.78, 0.85, 0.79, 0.79, 0.78, 0.78, 0.81, 0.84, 0.79, 0.83, 0.89, 0.92, 
    0.93, 0.88, 0.86, 0.9, 0.85, 0.84, 0.89, 0.9, 0.89, 0.86, 0.83, 0.83, 
    0.82, 0.71, 0.65, 0.7, 0.65, 0.67, 0.69, 0.67, 0.7, 0.7, 0.78, 0.72, 
    0.67, 0.58, 0.66, 0.74, 0.76, 0.8, 0.79, 0.74, 0.69, 0.75, 0.66, 0.69, 
    0.68, 0.73, 0.71, 0.71, 0.78, 0.75, 0.83, 0.75, 0.72, 0.8, 0.81, 0.82, 
    0.84, 0.86, 0.84, 0.87, 0.87, 0.91, 0.91, 0.88, 0.65, 0.6, 0.62, 0.65, 
    0.63, 0.64, 0.64, 0.67, 0.61, 0.65, 0.64, 0.64, 0.65, 0.67, 0.69, 0.71, 
    0.72, 0.77, 0.76, 0.8, 0.85, 0.77, 0.75, 0.85, 0.81, 0.83, 0.77, 0.76, 
    0.78, 0.77, 0.8, 0.81, 0.79, 0.76, 0.76, 0.73, 0.68, 0.68, 0.68, 0.67, 
    0.66, 0.69, 0.71, 0.66, 0.72, 0.77, 0.71, 0.76, 0.77, 0.81, 0.79, 0.78, 
    0.75, 0.72, 0.7, 0.62, 0.6, 0.59, 0.61, 0.65, 0.66, 0.64, 0.59, 0.59, 
    0.64, 0.64, 0.58, 0.64, 0.66, 0.63, 0.61, 0.58, 0.54, 0.61, 0.6, 0.59, 
    0.59, 0.56, 0.56, 0.67, 0.64, 0.66, 0.67, 0.63, 0.6, 0.55, 0.54, 0.54, 
    0.53, 0.53, 0.57, 0.58, 0.57, 0.57, 0.56, 0.56, 0.57, 0.57, 0.57, 0.58, 
    0.57, 0.56, 0.6, 0.62, 0.53, 0.53, 0.51, 0.52, 0.54, 0.53, 0.59, 0.67, 
    0.61, 0.64, 0.58, 0.59, 0.53, 0.52, 0.65, 0.67, 0.59, 0.55, 0.53, 0.51, 
    0.61, 0.6, 0.57, 0.63, 0.6, 0.63, 0.61, 0.62, 0.6, 0.61, 0.7, 0.68, 0.69, 
    0.68, 0.72, 0.71, 0.7, 0.7, 0.66, 0.69, 0.7, 0.63, 0.64, 0.64, 0.63, 
    0.65, 0.64, 0.63, 0.65, 0.67, 0.68, 0.66, 0.69, 0.69, 0.67, 0.61, 0.58, 
    0.59, 0.6, 0.58, 0.57, 0.54, 0.57, 0.56, 0.59, 0.59, 0.59, 0.56, 0.57, 
    0.57, 0.58, 0.59, 0.57, 0.58, 0.56, 0.57, 0.55, 0.59, 0.61, 0.61, 0.59, 
    0.6, 0.61, 0.65, 0.64, 0.69, 0.67, 0.62, 0.63, 0.65, 0.66, 0.66, 0.65, 
    0.68, 0.71, 0.81, 0.88, 0.87, 0.86, 0.87, 0.85, 0.84, 0.87, 0.88, 0.9, 
    0.88, 0.89, 0.89, 0.92, 0.91, 0.91, 0.91, 0.88, 0.91, 0.9, 0.87, 0.85, 
    0.87, 0.85, 0.83, 0.66, 0.6, 0.55, 0.51, 0.48, 0.5, 0.6, 0.62, 0.61, 
    0.47, 0.46, 0.46, 0.53, 0.46, 0.5, 0.47, 0.48, 0.5, 0.47, 0.46, 0.47, 
    0.46, 0.48, 0.44, 0.5, 0.5, 0.52, 0.58, 0.75, 0.83, 0.64, 0.5, 0.52, 
    0.52, 0.53, 0.5, 0.5, 0.44, 0.45, 0.44, 0.47, 0.48, 0.54, 0.55, 0.59, 
    0.64, 0.59, 0.64, 0.64, 0.68, 0.67, 0.68, 0.64, 0.62, 0.68, 0.65, 0.65, 
    0.65, 0.65, 0.68, 0.63, 0.66, 0.61, 0.63, 0.61, 0.62, 0.62, 0.61, 0.66, 
    0.69, 0.65, 0.65, 0.67, 0.7, 0.67, 0.68, 0.67, 0.64, 0.61, 0.62, 0.64, 
    0.62, 0.51, 0.6, 0.6, 0.61, 0.63, 0.61, 0.63, 0.68, 0.62, 0.64, 0.65, 
    0.67, 0.66, 0.7, 0.68, 0.59, 0.63, 0.6, 0.58, 0.55, 0.52, 0.47, 0.44, 
    0.46, 0.52, 0.58, 0.6, 0.58, 0.58, 0.59, 0.58, 0.49, 0.47, 0.45, 0.39, 
    0.36, 0.35, 0.44, 0.45, 0.48, 0.49, 0.5, 0.5, 0.49, 0.5, 0.47, 0.46, 
    0.49, 0.47, 0.46, 0.48, 0.45, 0.46, 0.46, 0.47, 0.53, 0.51, 0.44, 0.43, 
    0.44, 0.41, 0.5, 0.55, 0.59, 0.6, 0.56, 0.59, 0.55, 0.55, 0.54, 0.54, 
    0.57, 0.57, 0.6, 0.59, 0.58, 0.65, 0.68, 0.67, 0.72, 0.72, 0.72, 0.72, 
    0.72, 0.75, 0.82, 0.82, 0.84, 0.84, 0.85, 0.83, 0.84, 0.88, 0.88, 0.9, 
    0.9, 0.91, 0.91, 0.92, 0.83, 0.85, 0.81, 0.79, 0.81, 0.89, 0.78, 0.8, 
    0.74, 0.66, 0.69, 0.66, 0.74, 0.78, 0.75, 0.81, 0.82, 0.8, 0.8, 0.78, 
    0.78, 0.76, 0.79, 0.74, 0.72, 0.75, 0.66, 0.63, 0.71, 0.72, 0.77, 0.78, 
    0.76, 0.73, 0.7, 0.58, 0.63, 0.58, 0.52, 0.54, 0.59, 0.61, 0.59, 0.55, 
    0.54, 0.55, 0.59, 0.6, 0.49, 0.54, 0.61, 0.58, 0.6, 0.57, 0.6, 0.58, 
    0.61, 0.68, 0.72, 0.62, 0.64, 0.59, 0.59, 0.52, 0.6, 0.6, 0.56, 0.49, 
    0.41, 0.38, 0.49, 0.54, 0.53, 0.54, 0.57, 0.59, 0.62, 0.58, 0.58, 0.55, 
    0.55, 0.52, 0.49, 0.5, 0.4, 0.4, 0.4, 0.4, 0.41, 0.45, 0.46, 0.47, 0.45, 
    0.43, 0.43, 0.46, 0.46, 0.48, 0.47, 0.45, 0.45, 0.42, 0.39, 0.42, 0.38, 
    0.41, 0.49, 0.53, 0.53, 0.53, 0.52, 0.52, 0.55, 0.57, 0.57, 0.56, 0.56, 
    0.56, 0.56, 0.58, 0.53, 0.53, 0.56, 0.55, 0.56, 0.54, 0.57, 0.57, 0.61, 
    0.59, 0.62, 0.65, 0.6, 0.57, 0.63, 0.62, 0.64, 0.67, 0.63, 0.72, 0.75, 
    0.71, 0.69, 0.63, 0.58, 0.59, 0.64, 0.65, 0.73, 0.66, 0.56, 0.6, 0.6, 
    0.55, 0.55, 0.54, 0.53, 0.55, 0.54, 0.54, 0.5, 0.52, 0.55, 0.58, 0.6, 
    0.59, 0.62, 0.6, 0.66, 0.65, 0.62, 0.66, 0.66, 0.66, 0.65, 0.68, 0.66, 
    0.66, 0.65, 0.6, 0.6, 0.59, 0.57, 0.58, 0.63, 0.62, 0.62, 0.6, 0.64, 
    0.63, 0.64, 0.62, 0.64, 0.63, 0.63, 0.62, 0.65, 0.66, 0.64, 0.67, 0.67, 
    0.63, 0.71, 0.72, 0.72, 0.74, 0.73, 0.73, 0.73, 0.73, 0.75, 0.65, 0.64, 
    0.7, 0.61, 0.62, 0.64, 0.69, 0.69, 0.67, 0.73, 0.68, 0.7, 0.7, 0.67, 
    0.71, 0.72, 0.74, 0.71, 0.72, 0.72, 0.74, 0.73, 0.71, 0.71, 0.71, 0.68, 
    0.74, 0.7, 0.72, 0.67, 0.66, 0.66, 0.65, 0.67, 0.65, 0.65, 0.64, 0.66, 
    0.64, 0.65, 0.66, 0.63, 0.66, 0.69, 0.67, 0.69, 0.67, 0.68, 0.67, 0.66, 
    0.64, 0.63, 0.61, 0.66, 0.66, 0.63, 0.68, 0.69, 0.67, 0.66, 0.67, 0.68, 
    0.65, 0.63, 0.67, 0.68, 0.7, 0.67, 0.67, 0.66, 0.69, 0.77, 0.88, 0.92, 
    0.91, 0.85, 0.89, 0.87, 0.92, 0.93, 0.93, 0.93, 0.96, 0.95, 0.96, 0.96, 
    0.97, 0.84, 0.77, 0.87, 0.83, 0.84, 0.89, 0.88, 0.84, 0.79, 0.79, 0.81, 
    0.93, 0.95, 0.95, 0.94, 0.94, 0.94, 0.93, 0.91, 0.87, 0.79, 0.84, 0.88, 
    0.79, 0.89, 0.93, 0.89, 0.88, 0.88, 0.86, 0.9, 0.9, 0.92, 0.88, 0.9, 
    0.93, 0.87, 0.88, 0.91, 0.91, 0.92, 0.85, 0.88, 0.9, 0.91, 0.89, 0.87, 
    0.89, 0.89, 0.9, 0.93, 0.95, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.94, 
    0.91, 0.87, 0.88, 0.91, 0.94, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 0.96, 
    0.97, 0.97, 0.84, 0.79, 0.79, 0.77, 0.83, 0.79, 0.8, 0.8, 0.79, 0.83, 
    0.76, 0.76, 0.78, 0.76, 0.76, 0.73, 0.7, 0.66, 0.69, 0.7, 0.74, 0.75, 
    0.72, 0.73, 0.7, 0.89, 0.84, 0.81, 0.83, 0.88, 0.92, 0.91, 0.78, 0.92, 
    0.9, 0.88, 0.76, 0.66, 0.65, 0.66, 0.68, 0.75, 0.81, 0.79, 0.73, 0.75, 
    0.77, 0.74, 0.68, 0.76, 0.75, 0.72, 0.68, 0.66, 0.74, 0.88, 0.9, 0.91, 
    0.94, 0.9, 0.81, 0.88, 0.84, 0.62, 0.7, 0.69, 0.72, 0.75, 0.86, 0.81, 
    0.92, 0.95, 0.96, 0.95, 0.78, 0.71, 0.66, 0.75, 0.7, 0.81, 0.82, 0.82, 
    0.86, 0.77, 0.91, 0.95, 0.95, 0.9, 0.9, 0.88, 0.77, 0.82, 0.8, 0.76, 
    0.88, 0.87, 0.71, 0.66, 0.65, 0.67, 0.7, 0.73, 0.64, 0.68, 0.68, 0.62, 
    0.7, 0.65, 0.66, 0.62, 0.66, 0.67, 0.68, 0.7, 0.64, 0.64, 0.64, 0.67, 
    0.67, 0.67, 0.67, 0.7, 0.72, 0.66, 0.64, 0.69, 0.7, 0.76, 0.77, 0.83, 
    0.84, 0.86, 0.88, 0.88, 0.9, 0.88, 0.89, 0.82, 0.78, 0.74, 0.71, 0.72, 
    0.76, 0.78, 0.65, 0.66, 0.66, 0.75, 0.76, 0.78, 0.79, 0.8, 0.8, 0.8, 
    0.79, 0.79, 0.82, 0.83, 0.79, 0.79, 0.8, 0.76, 0.73, 0.74, 0.75, 0.73, 
    0.76, 0.79, 0.75, 0.75, 0.79, 0.81, 0.79, 0.77, 0.88, 0.9, 0.91, 0.87, 
    0.83, 0.86, 0.81, 0.8, 0.81, 0.79, 0.79, 0.84, 0.78, 0.77, 0.77, 0.71, 
    0.7, 0.65, 0.7, 0.59, 0.59, 0.62, 0.78, 0.81, 0.77, 0.72, 0.71, 0.64, 
    0.59, 0.56, 0.54, 0.54, 0.5, 0.53, 0.51, 0.59, 0.54, 0.5, 0.6, 0.56, 
    0.53, 0.57, 0.55, 0.62, 0.62, 0.65, 0.8, 0.85, 0.9, 0.9, 0.91, 0.91, 
    0.87, 0.84, 0.81, 0.77, 0.73, 0.78, 0.81, 0.85, 0.8, 0.87, 0.76, 0.76, 
    0.74, 0.71, 0.68, 0.79, 0.8, 0.76, 0.74, 0.8, 0.84, 0.86, 0.87, 0.82, 
    0.89, 0.92, 0.92, 0.91, 0.86, 0.9, 0.91, 0.91, 0.89, 0.84, 0.82, 0.77, 
    0.75, 0.75, 0.68, 0.63, 0.64, 0.63, 0.64, 0.63, 0.61, 0.62, 0.6, 0.57, 
    0.62, 0.59, 0.56, 0.57, 0.6, 0.63, 0.63, 0.6, 0.64, 0.63, 0.65, 0.62, 
    0.62, 0.6, 0.61, 0.61, 0.7, 0.66, 0.63, 0.76, 0.65, 0.56, 0.44, 0.46, 
    0.47, 0.5, 0.5, 0.49, 0.53, 0.58, 0.52, 0.54, 0.54, 0.49, 0.49, 0.49, 
    0.5, 0.47, 0.47, 0.44, 0.47, 0.47, 0.46, 0.47, 0.44, 0.48, 0.51, 0.5, 
    0.49, 0.51, 0.49, 0.51, 0.5, 0.42, 0.49, 0.46, 0.48, 0.46, 0.44, 0.44, 
    0.45, 0.43, 0.43, 0.44, 0.47, 0.44, 0.45, 0.46, 0.49, 0.54, 0.56, 0.52, 
    0.56, 0.58, 0.53, 0.59, 0.57, 0.61, 0.6, 0.64, 0.59, 0.64, 0.56, 0.59, 
    0.63, 0.63, 0.62, 0.62, 0.64, 0.64, 0.67, 0.67, 0.67, 0.56, 0.57, 0.56, 
    0.64, 0.58, 0.57, 0.58, 0.54, 0.53, 0.52, 0.54, 0.61, 0.63, 0.6, 0.57, 
    0.61, 0.65, 0.68, 0.61, 0.63, 0.64, 0.65, 0.66, 0.67, 0.68, 0.69, 0.68, 
    0.65, 0.72, 0.74, 0.7, 0.73, 0.75, 0.72, 0.7, 0.69, 0.72, 0.65, 0.74, 
    0.69, 0.72, 0.69, 0.64, 0.81, 0.9, 0.9, 0.92, 0.91, 0.9, 0.89, 0.88, 
    0.71, 0.81, 0.73, 0.74, 0.74, 0.73, 0.78, 0.76, 0.71, 0.76, 0.78, 0.81, 
    0.71, 0.66, 0.64, 0.68, 0.75, 0.92, 0.81, 0.79, 0.72, 0.68, 0.64, 0.62, 
    0.64, 0.63, 0.62, 0.62, 0.6, 0.58, 0.68, 0.63, 0.66, 0.69, 0.71, 0.67, 
    0.67, 0.62, 0.61, 0.64, 0.62, 0.58, 0.58, 0.57, 0.56, 0.55, 0.54, 0.53, 
    0.48, 0.49, 0.51, 0.56, 0.64, 0.64, 0.6, 0.63, 0.63, 0.56, 0.57, 0.59, 
    0.6, 0.58, 0.58, 0.53, 0.56, 0.56, 0.58, 0.54, 0.5, 0.5, 0.51, 0.53, 
    0.54, 0.5, 0.55, 0.57, 0.59, 0.55, 0.58, 0.55, 0.52, 0.52, 0.52, 0.51, 
    0.5, 0.48, 0.51, 0.48, 0.46, 0.45, 0.46, 0.42, 0.41, 0.39, 0.41, 0.4, 
    0.41, 0.39, 0.4, 0.4, 0.39, 0.42, 0.45, 0.5, 0.55, 0.55, 0.53, 0.52, 
    0.52, 0.5, 0.52, 0.51, 0.47, 0.45, 0.5, 0.53, 0.55, 0.57, 0.56, 0.57, 
    0.55, 0.54, 0.58, 0.53, 0.53, 0.48, 0.41, 0.43, 0.48, 0.49, 0.48, 0.5, 
    0.49, 0.48, 0.48, 0.48, 0.5, 0.53, 0.54, 0.53, 0.52, 0.51, 0.49, 0.51, 
    0.5, 0.51, 0.56, 0.52, 0.56, 0.61, 0.54, 0.59, 0.59, 0.6, 0.61, 0.62, 
    0.66, 0.69, 0.79, 0.8, 0.76, 0.74, 0.73, 0.73, 0.71, 0.63, 0.61, 0.62, 
    0.62, 0.63, 0.63, 0.64, 0.64, 0.7, 0.63, 0.65, 0.7, 0.68, 0.62, 0.6, 
    0.61, 0.64, 0.61, 0.59, 0.61, 0.63, 0.58, 0.59, 0.6, 0.6, 0.64, 0.65, 
    0.64, 0.59, 0.61, 0.64, 0.62, 0.63, 0.57, 0.65, 0.66, 0.68, 0.76, 0.77, 
    0.84, 0.81, 0.75, 0.71, 0.7, 0.72, 0.69, 0.7, 0.7, 0.7, 0.63, 0.67, 0.66, 
    0.65, 0.62, 0.63, 0.62, 0.63, 0.64, 0.65, 0.67, 0.69, 0.68, 0.66, 0.64, 
    0.62, 0.64, 0.64, 0.62, 0.63, 0.65, 0.6, 0.62, 0.62, 0.67, 0.69, 0.64, 
    0.68, 0.6, 0.63, 0.67, 0.65, 0.71, 0.68, 0.72, 0.7, 0.7, 0.72, 0.73, 
    0.75, 0.69, 0.74, 0.75, 0.74, 0.68, 0.67, 0.68, 0.61, 0.68, 0.74, 0.72, 
    0.77, 0.82, 0.85, 0.88, 0.88, 0.88, 0.88, 0.89, 0.82, 0.71, 0.76, 0.73, 
    0.8, 0.78, 0.68, 0.68, 0.71, 0.82, 0.86, 0.87, 0.82, 0.7, 0.69, 0.65, 
    0.58, 0.58, 0.65, 0.7, 0.7, 0.69, 0.72, 0.7, 0.72, 0.72, 0.78, 0.8, 0.76, 
    0.82, 0.82, 0.74, 0.66, 0.69, 0.67, 0.74, 0.72, 0.51, 0.55, 0.61, 0.6, 
    0.4, 0.36, 0.39, 0.43, 0.48, 0.6, 0.73, 0.56, 0.5, 0.58, 0.59, 0.71, 
    0.75, 0.82, 0.74, 0.65, 0.59, 0.53, 0.54, 0.57, 0.53, 0.59, 0.58, 0.56, 
    0.6, 0.63, 0.66, 0.66, 0.76, 0.74, 0.78, 0.77, 0.7, 0.67, 0.68, 0.64, 
    0.63, 0.63, 0.56, 0.56, 0.53, 0.51, 0.39, 0.38, 0.43, 0.42, 0.43, 0.45, 
    0.49, 0.49, 0.49, 0.49, 0.45, 0.48, 0.52, 0.49, 0.48, 0.54, 0.46, 0.48, 
    0.46, 0.46, 0.47, 0.45, 0.46, 0.51, 0.48, 0.48, 0.5, 0.51, 0.55, 0.55, 
    0.64, 0.63, 0.54, 0.53, 0.52, 0.56, 0.59, 0.76, 0.47, 0.51, 0.52, 0.58, 
    0.61, 0.51, 0.48, 0.48, 0.54, 0.47, 0.44, 0.53, 0.52, 0.52, 0.55, 0.56, 
    0.58, 0.59, 0.64, 0.64, 0.66, 0.68, 0.63, 0.62, 0.62, 0.63, 0.67, 0.58, 
    0.6, 0.62, 0.64, 0.58, 0.6, 0.58, 0.59, 0.61, 0.62, 0.65, 0.65, 0.64, 
    0.63, 0.6, 0.63, 0.64, 0.66, 0.69, 0.66, 0.72, 0.69, 0.67, 0.65, 0.61, 
    0.63, 0.55, 0.53, 0.58, 0.57, 0.55, 0.52, 0.58, 0.54, 0.53, 0.63, 0.58, 
    0.65, 0.68, 0.69, 0.72, 0.73, 0.79, 0.84, 0.85, 0.88, 0.91, 0.92, 0.93, 
    0.94, 0.95, 0.95, 0.94, 0.95, 0.96, 0.95, 0.88, 0.74, 0.66, 0.65, 0.6, 
    0.58, 0.56, 0.55, 0.59, 0.58, 0.59, 0.54, 0.59, 0.59, 0.57, 0.57, 0.57, 
    0.58, 0.59, 0.56, 0.58, 0.55, 0.54, 0.53, 0.49, 0.48, 0.45, 0.45, 0.44, 
    0.47, 0.49, 0.51, 0.49, 0.51, 0.53, 0.52, 0.45, 0.49, 0.54, 0.52, 0.55, 
    0.56, 0.51, 0.53, 0.56, 0.56, 0.59, 0.56, 0.57, 0.58, 0.57, 0.61, 0.59, 
    0.64, 0.54, 0.52, 0.58, 0.61, 0.61, 0.6, 0.62, 0.66, 0.63, 0.6, 0.63, 
    0.62, 0.62, 0.59, 0.55, 0.52, 0.54, 0.54, 0.56, 0.52, 0.55, 0.53, 0.58, 
    0.55, 0.53, 0.54, 0.53, 0.52, 0.54, 0.54, 0.62, 0.59, 0.57, 0.56, 0.57, 
    0.59, 0.6, 0.57, 0.64, 0.54, 0.61, 0.54, 0.52, 0.56, 0.57, 0.57, 0.55, 
    0.52, 0.5, 0.57, 0.51, 0.56, 0.54, 0.55, 0.55, 0.57, 0.56, 0.58, 0.6, 
    0.58, 0.53, 0.53, 0.54, 0.52, 0.55, 0.54, 0.53, 0.55, 0.56, 0.55, 0.58, 
    0.59, 0.61, 0.6, 0.57, 0.56, 0.59, 0.56, 0.56, 0.52, 0.49, 0.57, 0.53, 
    0.46, 0.54, 0.51, 0.5, 0.53, 0.55, 0.66, 0.6, 0.55, 0.55, 0.51, 0.51, 
    0.55, 0.56, 0.52, 0.46, 0.5, 0.49, 0.44, 0.48, 0.48, 0.55, 0.55, 0.52, 
    0.46, 0.5, 0.55, 0.59, 0.54, 0.49, 0.5, 0.51, 0.55, 0.48, 0.52, 0.53, 
    0.54, 0.55, 0.54, 0.62, 0.61, 0.57, 0.6, 0.6, 0.53, 0.54, 0.53, 0.51, 
    0.47, 0.57, 0.57, 0.56, 0.58, 0.49, 0.44, 0.42, 0.4, 0.34, 0.31, 0.45, 
    0.5, 0.57, 0.59, 0.63, 0.66, 0.64, 0.62, 0.57, 0.59, 0.6, 0.59, 0.65, 
    0.66, 0.61, 0.59, 0.6, 0.59, 0.62, 0.61, 0.62, 0.63, 0.66, 0.69, 0.72, 
    0.71, 0.69, 0.69, 0.7, 0.68, 0.69, 0.67, 0.71, 0.79, 0.85, 0.82, 0.84, 
    0.91, 0.9, 0.91, 0.93, 0.95, 0.95, 0.95, 0.95, 0.94, 0.93, 0.9, 0.89, 
    0.9, 0.94, 0.93, 0.95, 0.96, 0.82, 0.78, 0.81, 0.8, 0.79, 0.8, 0.79, 0.8, 
    0.81, 0.81, 0.84, 0.86, 0.89, 0.88, 0.88, 0.85, 0.84, 0.85, 0.84, 0.85, 
    0.91, 0.92, 0.94, 0.93, 0.94, 0.94, 0.95, 0.9, 0.88, 0.91, 0.84, 0.87, 
    0.83, 0.84, 0.85, 0.85, 0.8, 0.84, 0.76, 0.76, 0.79, 0.8, 0.79, 0.79, 
    0.79, 0.8, 0.8, 0.85, 0.84, 0.83, 0.9, 0.91, 0.83, 0.81, 0.84, 0.82, 
    0.78, 0.78, 0.83, 0.86, 0.79, 0.85, 0.85, 0.85, 0.78, 0.8, 0.85, 0.75, 
    0.74, 0.77, 0.76, 0.78, 0.79, 0.8, 0.77, 0.8, 0.78, 0.82, 0.82, 0.81, 
    0.84, 0.78, 0.73, 0.7, 0.73, 0.72, 0.72, 0.75, 0.77, 0.75, 0.75, 0.73, 
    0.78, 0.78, 0.77, 0.8, 0.82, 0.83, 0.81, 0.81, 0.82, 0.78, 0.83, 0.82, 
    0.81, 0.79, 0.84, 0.84, 0.84, 0.86, 0.86, 0.87, 0.85, 0.88, 0.84, 0.83, 
    0.78, 0.82, 0.83, 0.81, 0.85, 0.8, 0.81, 0.77, 0.86, 0.79, 0.81, 0.78, 
    0.8, 0.82, 0.82, 0.79, 0.74, 0.66, 0.64, 0.71, 0.68, 0.72, 0.72, 0.66, 
    0.83, 0.79, 0.78, 0.72, 0.67, 0.68, 0.77, 0.85, 0.83, 0.68, 0.64, 0.71, 
    0.62, 0.77, 0.71, 0.68, 0.76, 0.81, 0.82, 0.8, 0.78, 0.82, 0.76, 0.77, 
    0.79, 0.73, 0.73, 0.72, 0.7, 0.67, 0.7, 0.73, 0.73, 0.72, 0.71, 0.73, 
    0.73, 0.78, 0.89, 0.85, 0.9, 0.84, 0.86, 0.81, 0.82, 0.8, 0.8, 0.83, 
    0.85, 0.74, 0.77, 0.92, 0.9, 0.9, 0.89, 0.62, 0.57, 0.62, 0.6, 0.59, 
    0.52, 0.56, 0.6, 0.65, 0.68, 0.58, 0.57, 0.59, 0.61, 0.59, 0.51, 0.56, 
    0.59, 0.6, 0.58, 0.63, 0.62, 0.67, 0.66, 0.65, 0.64, 0.63, 0.64, 0.61, 
    0.57, 0.57, 0.56, 0.57, 0.51, 0.5, 0.47, 0.5, 0.47, 0.59, 0.49, 0.59, 
    0.54, 0.47, 0.54, 0.51, 0.53, 0.46, 0.43, 0.5, 0.48, 0.47, 0.51, 0.52, 
    0.49, 0.48, 0.53, 0.57, 0.55, 0.65, 0.78, 0.8, 0.79, 0.79, 0.77, 0.78, 
    0.83, 0.84, 0.83, 0.83, 0.85, 0.85, 0.84, 0.84, 0.81, 0.66, 0.68, 0.71, 
    0.74, 0.76, 0.74, 0.72, 0.7, 0.7, 0.65, 0.63, 0.58, 0.57, 0.58, 0.52, 
    0.5, 0.56, 0.52, 0.56, 0.53, 0.5, 0.51, 0.53, 0.53, 0.51, 0.57, 0.57, 
    0.6, 0.57, 0.57, 0.56, 0.56, 0.58, 0.6, 0.59, 0.6, 0.57, 0.62, 0.61, 
    0.58, 0.59, 0.59, 0.6, 0.62, 0.63, 0.61, 0.61, 0.59, 0.58, 0.59, 0.59, 
    0.54, 0.59, 0.61, 0.57, 0.59, 0.6, 0.62, 0.62, 0.64, 0.62, 0.63, 0.62, 
    0.62, 0.62, 0.63, 0.61, 0.61, 0.62, 0.61, 0.62, 0.62, 0.64, 0.65, 0.65, 
    0.65, 0.65, 0.64, 0.65, 0.65, 0.66, 0.66, 0.59, 0.62, 0.64, 0.67, 0.72, 
    0.77, 0.81, 0.83, 0.83, 0.84, 0.85, 0.77, 0.79, 0.8, 0.76, 0.73, 0.76, 
    0.82, 0.77, 0.74, 0.7, 0.73, 0.61, 0.57, 0.6, 0.62, 0.65, 0.67, 0.6, 
    0.64, 0.59, 0.66, 0.8, 0.8, 0.74, 0.79, 0.71, 0.71, 0.7, 0.67, 0.68, 
    0.68, 0.76, 0.87, 0.88, 0.85, 0.81, 0.81, 0.74, 0.82, 0.85, 0.82, 0.85, 
    0.81, 0.85, 0.88, 0.92, 0.91, 0.84, 0.85, 0.81, 0.73, 0.68, 0.64, 0.59, 
    0.49, 0.42, 0.54, 0.59, 0.52, 0.57, 0.48, 0.52, 0.55, 0.49, 0.49, 0.48, 
    0.46, 0.49, 0.47, 0.55, 0.69, 0.59, 0.59, 0.52, 0.47, 0.43, 0.43, 0.52, 
    0.52, 0.45, 0.48, 0.47, 0.49, 0.54, 0.54, 0.6, 0.61, 0.54, 0.57, 0.58, 
    0.53, 0.53, 0.57, 0.57, 0.55, 0.56, 0.55, 0.54, 0.54, 0.55, 0.51, 0.52, 
    0.54, 0.58, 0.58, 0.6, 0.63, 0.66, 0.65, 0.65, 0.66, 0.7, 0.66, 0.57, 
    0.53, 0.55, 0.52, 0.51, 0.46, 0.47, 0.45, 0.53, 0.57, 0.58, 0.55, 0.56, 
    0.53, 0.48, 0.46, 0.53, 0.53, 0.56, 0.58, 0.61, 0.6, 0.63, 0.64, 0.64, 
    0.63, 0.67, 0.64, 0.63, 0.68, 0.67, 0.69, 0.67, 0.67, 0.67, 0.66, 0.64, 
    0.69, 0.68, 0.66, 0.64, 0.67, 0.65, 0.66, 0.68, 0.68, 0.67, 0.68, 0.64, 
    0.58, 0.61, 0.59, 0.6, 0.58, 0.67, 0.61, 0.71, 0.67, 0.64, 0.67, 0.67, 
    0.66, 0.65, 0.68, 0.69, 0.69, 0.68, 0.65, 0.6, 0.68, 0.66, 0.69, 0.74, 
    0.7, 0.68, 0.73, 0.76, 0.74, 0.73, 0.73, 0.79, 0.68, 0.69, 0.63, 0.66, 
    0.64, 0.62, 0.64, 0.63, 0.59, 0.62, 0.63, 0.63, 0.53, 0.61, 0.62, 0.6, 
    0.57, 0.68, 0.65, 0.61, 0.69, 0.62, 0.63, 0.66, 0.69, 0.68, 0.63, 0.64, 
    0.68, 0.71, 0.7, 0.65, 0.7, 0.68, 0.64, 0.66, 0.66, 0.69, 0.67, 0.64, 
    0.69, 0.69, 0.66, 0.7, 0.62, 0.7, 0.67, 0.62, 0.61, 0.63, 0.68, 0.72, 
    0.73, 0.68, 0.68, 0.7, 0.71, 0.67, 0.69, 0.66, 0.68, 0.64, 0.65, 0.61, 
    0.63, 0.55, 0.61, 0.63, 0.69, 0.63, 0.57, 0.58, 0.55, 0.61, 0.55, 0.57, 
    0.57, 0.58, 0.63, 0.59, 0.66, 0.65, 0.64, 0.65, 0.59, 0.59, 0.62, 0.61, 
    0.62, 0.69, 0.68, 0.67, 0.66, 0.66, 0.66, 0.6, 0.64, 0.64, 0.69, 0.63, 
    0.67, 0.66, 0.66, 0.67, 0.72, 0.68, 0.72, 0.72, 0.71, 0.71, 0.72, 0.7, 
    0.78, 0.79, 0.78, 0.76, 0.78, 0.8, 0.8, 0.84, 0.83, 0.82, 0.84, 0.87, 
    0.86, 0.89, 0.94, 0.94, 0.94, 0.95, 0.94, 0.94, 0.94, 0.95, 0.94, 0.94, 
    0.94, 0.94, 0.95, 0.94, 0.95, 0.95, 0.94, 0.94, 0.94, 0.83, 0.71, 0.71, 
    0.69, 0.66, 0.64, 0.64, 0.6, 0.57, 0.55, 0.54, 0.54, 0.52, 0.55, 0.57, 
    0.57, 0.56, 0.58, 0.6, 0.59, 0.64, 0.64, 0.66, 0.69, 0.71, 0.73, 0.75, 
    0.77, 0.77, 0.75, 0.81, 0.82, 0.81, 0.79, 0.8, 0.81, 0.78, 0.83, 0.86, 
    0.85, 0.85, 0.86, 0.87, 0.86, 0.86, 0.88, 0.87, 0.87, 0.87, 0.87, 0.88, 
    0.86, 0.89, 0.88, 0.9, 0.92, 0.91, 0.92, 0.92, 0.91, 0.91, 0.89, 0.91, 
    0.91, 0.91, 0.91, 0.93, 0.84, 0.81, 0.81, 0.77, 0.78, 0.71, 0.66, 0.65, 
    0.66, 0.67, 0.66, 0.66, 0.64, 0.64, 0.63, 0.64, 0.67, 0.64, 0.6, 0.6, 
    0.6, 0.59, 0.59, 0.59, 0.59, 0.59, 0.58, 0.58, 0.59, 0.58, 0.58, 0.58, 
    0.59, 0.6, 0.62, 0.63, 0.66, 0.66, 0.67, 0.66, 0.65, 0.67, 0.72, 0.76, 
    0.8, 0.77, 0.82, 0.85, 0.87, 0.88, 0.71, 0.76, 0.71, 0.67, 0.64, 0.65, 
    0.7, 0.66, 0.6, 0.62, 0.54, 0.55, 0.59, 0.6, 0.56, 0.47, 0.5, 0.56, 0.57, 
    0.63, 0.57, 0.62, 0.6, 0.57, 0.53, 0.49, 0.51, 0.47, 0.61, 0.63, 0.65, 
    0.64, 0.58, 0.53, 0.48, 0.52, 0.54, 0.58, 0.63, 0.69, 0.65, 0.69, 0.64, 
    0.59, 0.54, 0.5, 0.51, 0.54, 0.53, 0.57, 0.54, 0.54, 0.54, 0.56, 0.56, 
    0.6, 0.6, 0.58, 0.6, 0.59, 0.66, 0.58, 0.67, 0.71, 0.7, 0.7, 0.7, 0.72, 
    0.78, 0.82, 0.83, 0.86, 0.87, 0.88, 0.88, 0.87, 0.87, 0.85, 0.88, 0.87, 
    0.9, 0.89, 0.89, 0.9, 0.88, 0.88, 0.88, 0.87, 0.87, 0.87, 0.85, 0.87, 
    0.86, 0.88, 0.86, 0.92, 0.93, 0.95, 0.84, 0.87, 0.89, 0.8, 0.89, 0.89, 
    0.83, 0.85, 0.82, 0.9, 0.93, 0.93, 0.88, 0.89, 0.88, 0.94, 0.95, 0.92, 
    0.88, 0.86, 0.82, 0.79, 0.71, 0.69, 0.73, 0.73, 0.72, 0.66, 0.67, 0.67, 
    0.69, 0.71, 0.66, 0.66, 0.69, 0.66, 0.71, 0.7, 0.69, 0.68, 0.67, 0.71, 
    0.7, 0.74, 0.68, 0.68, 0.64, 0.66, 0.63, 0.61, 0.65, 0.64, 0.67, 0.67, 
    0.64, 0.64, 0.69, 0.64, 0.6, 0.62, 0.62, 0.6, 0.66, 0.62, 0.64, 0.56, 
    0.59, 0.66, 0.6, 0.58, 0.57, 0.58, 0.6, 0.55, 0.6, 0.53, 0.57, 0.53, 
    0.54, 0.53, 0.58, 0.6, 0.58, 0.58, 0.59, 0.57, 0.56, 0.59, 0.52, 0.55, 
    0.56, 0.57, 0.55, 0.59, 0.58, 0.57, 0.57, 0.54, 0.54, 0.59, 0.56, 0.65, 
    0.63, 0.65, 0.64, 0.7, 0.68, 0.66, 0.67, 0.64, 0.66, 0.64, 0.7, 0.67, 
    0.64, 0.66, 0.69, 0.68, 0.64, 0.64, 0.64, 0.64, 0.57, 0.68, 0.69, 0.71, 
    0.77, 0.79, 0.77, 0.77, 0.78, 0.83, 0.71, 0.76, 0.76, 0.76, 0.74, 0.75, 
    0.76, 0.78, 0.78, 0.78, 0.79, 0.77, 0.73, 0.65, 0.65, 0.59, 0.61, 0.65, 
    0.68, 0.69, 0.68, 0.7, 0.71, 0.67, 0.69, 0.64, 0.66, 0.66, 0.71, 0.69, 
    0.7, 0.7, 0.65, 0.65, 0.62, 0.63, 0.59, 0.55, 0.52, 0.55, 0.53, 0.56, 
    0.6, 0.67, 0.61, 0.65, 0.68, 0.68, 0.63, 0.67, 0.65, 0.59, 0.67, 0.61, 
    0.69, 0.64, 0.56, 0.61, 0.66, 0.62, 0.63, 0.63, 0.58, 0.58, 0.6, 0.64, 
    0.66, 0.68, 0.67, 0.62, 0.69, 0.65, 0.69, 0.7, 0.72, 0.77, 0.83, 0.86, 
    0.85, 0.84, 0.84, 0.84, 0.83, 0.84, 0.86, 0.84, 0.86, 0.84, 0.84, 0.86, 
    0.84, 0.71, 0.64, 0.66, 0.61, 0.58, 0.57, 0.56, 0.57, 0.58, 0.57, 0.59, 
    0.61, 0.63, 0.64, 0.64, 0.61, 0.61, 0.64, 0.67, 0.66, 0.68, 0.63, 0.63, 
    0.63, 0.65, 0.61, 0.59, 0.58, 0.56, 0.58, 0.56, 0.57, 0.59, 0.57, 0.54, 
    0.59, 0.56, 0.59, 0.58, 0.5, 0.52, 0.52, 0.51, 0.47, 0.51, 0.51, 0.53, 
    0.51, 0.52, 0.63, 0.64, 0.58, 0.55, 0.58, 0.66, 0.56, 0.55, 0.54, 0.56, 
    0.58, 0.53, 0.56, 0.53, 0.5, 0.51, 0.54, 0.59, 0.54, 0.51, 0.55, 0.53, 
    0.55, 0.55, 0.54, 0.56, 0.59, 0.56, 0.56, 0.58, 0.64, 0.6, 0.6, 0.54, 
    0.53, 0.53, 0.53, 0.53, 0.54, 0.53, 0.52, 0.51, 0.57, 0.6, 0.59, 0.53, 
    0.53, 0.5, 0.51, 0.53, 0.55, 0.55, 0.55, 0.53, 0.5, 0.53, 0.57, 0.52, 
    0.49, 0.51, 0.5, 0.54, 0.51, 0.58, 0.54, 0.51, 0.55, 0.51, 0.56, 0.51, 
    0.57, 0.48, 0.47, 0.48, 0.49, 0.5, 0.54, 0.54, 0.57, 0.57, 0.62, 0.65, 
    0.65, 0.64, 0.62, 0.58, 0.58, 0.58, 0.58, 0.6, 0.55, 0.6, 0.57, 0.57, 
    0.51, 0.49, 0.47, 0.53, 0.54, 0.56, 0.55, 0.57, 0.58, 0.58, 0.57, 0.56, 
    0.57, 0.59, 0.56, 0.57, 0.62, 0.61, 0.63, 0.6, 0.57, 0.53, 0.5, 0.52, 
    0.56, 0.62, 0.58, 0.6, 0.57, 0.61, 0.57, 0.53, 0.57, 0.6, 0.6, 0.63, 0.6, 
    0.6, 0.61, 0.6, 0.62, 0.55, 0.53, 0.47, 0.49, 0.48, 0.54, 0.54, 0.58, 
    0.55, 0.55, 0.58, 0.59, 0.59, 0.6, 0.59, 0.59, 0.58, 0.6, 0.57, 0.59, 
    0.59, 0.61, 0.63, 0.62, 0.59, 0.56, 0.55, 0.52, 0.53, 0.56, 0.59, 0.56, 
    0.55, 0.57, 0.6, 0.64, 0.61, 0.63, 0.6, 0.62, 0.63, 0.69, 0.64, 0.62, 
    0.63, 0.67, 0.67, 0.65, 0.56, 0.61, 0.54, 0.61, 0.53, 0.5, 0.6, 0.59, 
    0.63, 0.58, 0.65, 0.66, 0.66, 0.7, 0.79, 0.84, 0.86, 0.86, 0.87, 0.85, 
    0.87, 0.85, 0.86, 0.8, 0.73, 0.69, 0.63, 0.57, 0.55, 0.54, 0.51, 0.49, 
    0.51, 0.48, 0.49, 0.57, 0.51, 0.52, 0.53, 0.52, 0.55, 0.58, 0.61, 0.6, 
    0.59, 0.58, 0.57, 0.56, 0.55, 0.54, 0.53, 0.52, 0.49, 0.52, 0.56, 0.57, 
    0.53, 0.53, 0.54, 0.55, 0.58, 0.59, 0.57, 0.57, 0.58, 0.6, 0.66, 0.73, 
    0.77, 0.77, 0.74, 0.66, 0.45, 0.43, 0.43, 0.35, 0.37, 0.35, 0.35, 0.37, 
    0.33, 0.46, 0.38, 0.31, 0.25, 0.24, 0.35, 0.38, 0.47, 0.54, 0.53, 0.54, 
    0.57, 0.59, 0.55, 0.52, 0.5, 0.5, 0.47, 0.5, 0.5, 0.52, 0.51, 0.53, 0.58, 
    0.55, 0.54, 0.6, 0.59, 0.61, 0.61, 0.59, 0.68, 0.65, 0.68, 0.69, 0.7, 
    0.67, 0.63, 0.59, 0.56, 0.56, 0.55, 0.52, 0.55, 0.57, 0.58, 0.53, 0.58, 
    0.58, 0.59, 0.67, 0.63, 0.66, 0.65, 0.67, 0.62, 0.68, 0.65, 0.65, 0.71, 
    0.72, 0.69, 0.61, 0.56, 0.66, 0.6, 0.62, 0.67, 0.77, 0.79, 0.86, 0.8, 
    0.74, 0.82, 0.82, 0.83, 0.81, 0.87, 0.92, 0.9, 0.86, 0.89, 0.8, 0.81, 
    0.84, 0.87, 0.9, 0.91, 0.88, 0.85, 0.68, 0.65, 0.59, 0.6, 0.58, 0.58, 
    0.59, 0.6, 0.64, 0.58, 0.61, 0.65, 0.65, 0.67, 0.66, 0.7, 0.66, 0.62, 
    0.6, 0.61, 0.59, 0.55, 0.53, 0.54, 0.55, 0.55, 0.51, 0.54, 0.54, 0.54, 
    0.58, 0.56, 0.6, 0.62, 0.62, 0.63, 0.67, 0.66, 0.59, 0.72, 0.69, 0.66, 
    0.68, 0.71, 0.57, 0.55, 0.56, 0.53, 0.52, 0.51, 0.48, 0.51, 0.55, 0.57, 
    0.56, 0.63, 0.64, 0.72, 0.64, 0.68, 0.73, 0.72, 0.77, 0.68, 0.73, 0.6, 
    0.5, 0.5, 0.5, 0.53, 0.49, 0.51, 0.48, 0.49, 0.45, 0.48, 0.5, 0.5, 0.54, 
    0.61, 0.61, 0.66, 0.68, 0.7, 0.69, 0.7, 0.69, 0.7, 0.77, 0.68, 0.68, 
    0.68, 0.66, 0.62, 0.58, 0.53, 0.59, 0.55, 0.63, 0.54, 0.54, 0.67, 0.67, 
    0.71, 0.74, 0.75, 0.78, 0.74, 0.74, 0.77, 0.84, 0.87, 0.88, 0.85, 0.8, 
    0.76, 0.69, 0.66, 0.59, 0.54, 0.51, 0.48, 0.46, 0.45, 0.46, 0.47, 0.49, 
    0.5, 0.5, 0.56, 0.6, 0.59, 0.63, 0.64, 0.69, 0.64, 0.64, 0.62, 0.6, 0.59, 
    0.57, 0.55, 0.53, 0.55, 0.54, 0.53, 0.54, 0.52, 0.54, 0.51, 0.53, 0.54, 
    0.56, 0.61, 0.61, 0.6, 0.56, 0.6, 0.59, 0.62, 0.62, 0.61, 0.6, 0.62, 
    0.64, 0.63, 0.6, 0.6, 0.55, 0.52, 0.57, 0.51, 0.59, 0.54, 0.54, 0.59, 
    0.62, 0.66, 0.69, 0.73, 0.73, 0.72, 0.68, 0.71, 0.67, 0.67, 0.66, 0.65, 
    0.62, 0.64, 0.58, 0.57, 0.54, 0.59, 0.57, 0.59, 0.53, 0.53, 0.57, 0.68, 
    0.68, 0.72, 0.74, 0.7, 0.58, 0.58, 0.58, 0.59, 0.6, 0.61, 0.61, 0.59, 
    0.62, 0.54, 0.53, 0.47, 0.47, 0.51, 0.61, 0.59, 0.58, 0.62, 0.57, 0.58, 
    0.65, 0.61, 0.68, 0.72, 0.69, 0.75, 0.7, 0.72, 0.7, 0.72, 0.64, 0.62, 
    0.56, 0.58, 0.6, 0.63, 0.57, 0.57, 0.6, 0.6, 0.57, 0.57, 0.58, 0.58, 0.6, 
    0.63, 0.65, 0.68, 0.7, 0.64, 0.64, 0.65, 0.62, 0.6, 0.63, 0.69, 0.7, 
    0.59, 0.55, 0.51, 0.5, 0.52, 0.55, 0.53, 0.48, 0.46, 0.5, 0.48, 0.49, 
    0.54, 0.52, 0.52, 0.44, 0.47, 0.51, 0.51, 0.5, 0.47, 0.46, 0.45, 0.47, 
    0.48, 0.49, 0.46, 0.46, 0.45, 0.48, 0.47, 0.49, 0.52, 0.54, 0.53, 0.53, 
    0.53, 0.54, 0.52, 0.56, 0.53, 0.54, 0.56, 0.59, 0.62, 0.65, 0.64, 0.61, 
    0.57, 0.54, 0.58, 0.54, 0.54, 0.6, 0.55, 0.58, 0.57, 0.62, 0.59, 0.61, 
    0.66, 0.69, 0.69, 0.71, 0.71, 0.72, 0.69, 0.69, 0.69, 0.64, 0.6, 0.59, 
    0.55, 0.53, 0.61, 0.59, 0.57, 0.53, 0.55, 0.54, 0.53, 0.57, 0.56, 0.6, 
    0.62, 0.67, 0.67, 0.69, 0.7, 0.7, 0.68, 0.67, 0.69, 0.71, 0.72, 0.65, 
    0.6, 0.57, 0.6, 0.49, 0.57, 0.58, 0.59, 0.6, 0.61, 0.63, 0.66, 0.65, 
    0.71, 0.74, 0.75, 0.77, 0.76, 0.77, 0.78, 0.78, 0.78, 0.71, 0.69, 0.64, 
    0.59, 0.54, 0.54, 0.56, 0.59, 0.55, 0.61, 0.63, 0.63, 0.68, 0.67, 0.69, 
    0.68, 0.74, 0.74, 0.79, 0.74, 0.75, 0.78, 0.79, 0.79, 0.67, 0.71, 0.65, 
    0.64, 0.67, 0.68, 0.68, 0.7, 0.65, 0.66, 0.68, 0.64, 0.68, 0.68, 0.72, 
    0.76, 0.8, 0.84, 0.88, 0.88, 0.88, 0.74, 0.68, 0.7, 0.71, 0.79, 0.78, 
    0.65, 0.67, 0.67, 0.69, 0.74, 0.75, 0.81, 0.79, 0.78, 0.82, 0.83, 0.85, 
    0.86, 0.83, 0.85, 0.83, 0.87, 0.88, 0.84, 0.76, 0.7, 0.72, 0.74, 0.81, 
    0.8, 0.77, 0.71, 0.71, 0.7, 0.69, 0.75, 0.8, 0.74, 0.68, 0.83, 0.87, 
    0.88, 0.87, 0.87, 0.86, 0.83, 0.87, 0.85, 0.82, 0.76, 0.81, 0.77, 0.79, 
    0.79, 0.79, 0.8, 0.75, 0.74, 0.77, 0.72, 0.67, 0.57, 0.66, 0.68, 0.69, 
    0.7, 0.71, 0.72, 0.74, 0.76, 0.82, 0.79, 0.76, 0.77, 0.78, 0.72, 0.71, 
    0.67, 0.65, 0.6, 0.6, 0.62, 0.66, 0.63, 0.63, 0.68, 0.68, 0.67, 0.73, 
    0.69, 0.72, 0.71, 0.72, 0.76, 0.75, 0.77, 0.79, 0.8, 0.82, 0.81, 0.78, 
    0.77, 0.72, 0.71, 0.69, 0.73, 0.74, 0.74, 0.74, 0.74, 0.77, 0.77, 0.84, 
    0.84, 0.84, 0.84, 0.82, 0.81, 0.82, 0.78, 0.77, 0.75, 0.73, 0.73, 0.72, 
    0.7, 0.66, 0.64, 0.62, 0.61, 0.62, 0.62, 0.64, 0.65, 0.66, 0.66, 0.7, 
    0.69, 0.73, 0.76, 0.77, 0.77, 0.74, 0.78, 0.78, 0.73, 0.69, 0.68, 0.66, 
    0.69, 0.69, 0.75, 0.84, 0.91, 0.91, 0.91, 0.91, 0.92, 0.89, 0.83, 0.86, 
    0.89, 0.87, 0.89, 0.88, 0.91, 0.94, 0.94, 0.94, 0.95, 0.94, 0.91, 0.79, 
    0.79, 0.8, 0.78, 0.8, 0.78, 0.77, 0.75, 0.69, 0.69, 0.69, 0.67, 0.68, 
    0.66, 0.65, 0.65, 0.65, 0.65, 0.61, 0.6, 0.6, 0.58, 0.58, 0.56, 0.54, 
    0.52, 0.48, 0.52, 0.49, 0.52, 0.51, 0.51, 0.61, 0.59, 0.49, 0.56, 0.57, 
    0.55, 0.6, 0.62, 0.62, 0.63, 0.65, 0.64, 0.7, 0.67, 0.64, 0.64, 0.6, 
    0.57, 0.58, 0.59, 0.64, 0.51, 0.56, 0.48, 0.48, 0.5, 0.5, 0.55, 0.51, 
    0.54, 0.57, 0.55, 0.53, 0.57, 0.56, 0.55, 0.54, 0.59, 0.55, 0.54, 0.55, 
    0.51, 0.52, 0.5, 0.54, 0.51, 0.52, 0.52, 0.51, 0.52, 0.54, 0.54, 0.57, 
    0.58, 0.59, 0.61, 0.59, 0.62, 0.62, 0.62, 0.62, 0.62, 0.61, 0.59, 0.57, 
    0.55, 0.56, 0.54, 0.54, 0.55, 0.57, 0.59, 0.6, 0.58, 0.6, 0.61, 0.58, 
    0.64, 0.65, 0.63, 0.64, 0.65, 0.64, 0.64, 0.64, 0.63, 0.61, 0.61, 0.57, 
    0.56, 0.57, 0.54, 0.56, 0.55, 0.57, 0.55, 0.58, 0.59, 0.56, 0.54, 0.58, 
    0.59, 0.6, 0.6, 0.59, 0.6, 0.59, 0.58, 0.6, 0.57, 0.56, 0.56, 0.56, 0.6, 
    0.59, 0.58, 0.58, 0.59, 0.53, 0.58, 0.6, 0.59, 0.62, 0.62, 0.64, 0.68, 
    0.7, 0.71, 0.71, 0.68, 0.73, 0.72, 0.7, 0.69, 0.68, 0.66, 0.64, 0.61, 
    0.61, 0.64, 0.62, 0.61, 0.6, 0.59, 0.61, 0.62, 0.64, 0.65, 0.66, 0.65, 
    0.68, 0.69, 0.7, 0.73, 0.73, 0.76, 0.72, 0.7, 0.69, 0.72, 0.68, 0.68, 
    0.65, 0.64, 0.65, 0.65, 0.68, 0.67, 0.68, 0.68, 0.69, 0.69, 0.7, 0.69, 
    0.71, 0.72, 0.72, 0.73, 0.74, 0.74, 0.81, 0.73, 0.73, 0.69, 0.68, 0.66, 
    0.59, 0.64, 0.68, 0.67, 0.66, 0.63, 0.66, 0.64, 0.56, 0.61, 0.64, 0.66, 
    0.65, 0.73, 0.74, 0.7, 0.75, 0.74, 0.72, 0.67, 0.69, 0.66, 0.62, 0.58, 
    0.58, 0.63, 0.59, 0.58, 0.57, 0.6, 0.58, 0.55, 0.6, 0.56, 0.62, 0.56, 
    0.58, 0.66, 0.86, 0.85, 0.91, 0.93, 0.9, 0.78, 0.71, 0.69, 0.6, 0.66, 
    0.63, 0.62, 0.68, 0.68, 0.65, 0.59, 0.61, 0.62, 0.61, 0.61, 0.66, 0.66, 
    0.68, 0.7, 0.73, 0.75, 0.77, 0.78, 0.81, 0.71, 0.7, 0.69, 0.64, 0.6, 
    0.63, 0.6, 0.51, 0.53, 0.5, 0.45, 0.47, 0.48, 0.45, 0.48, 0.5, 0.52, 
    0.57, 0.68, 0.67, 0.67, 0.67, 0.67, 0.67, 0.67, 0.66, 0.63, 0.61, 0.56, 
    0.63, 0.61, 0.55, 0.59, 0.55, 0.54, 0.58, 0.6, 0.58, 0.62, 0.63, 0.64, 
    0.63, 0.68, 0.66, 0.66, 0.67, 0.68, 0.68, 0.68, 0.68, 0.68, 0.69, 0.65, 
    0.68, 0.63, 0.64, 0.63, 0.61, 0.55, 0.58, 0.64, 0.69, 0.68, 0.66, 0.64, 
    0.67, 0.67, 0.66, 0.7, 0.72, 0.72, 0.72, 0.73, 0.78, 0.76, 0.71, 0.7, 
    0.68, 0.64, 0.63, 0.62, 0.65, 0.67, 0.68, 0.66, 0.64, 0.69, 0.72, 0.76, 
    0.74, 0.77, 0.78, 0.79, 0.77, 0.76, 0.77, 0.76, 0.74, 0.71, 0.71, 0.7, 
    0.63, 0.66, 0.62, 0.66, 0.64, 0.62, 0.62, 0.6, 0.62, 0.71, 0.77, 0.83, 
    0.88, 0.85, 0.87, 0.88, 0.88, 0.87, 0.9, 0.89, 0.89, 0.87, 0.86, 0.88, 
    0.82, 0.83, 0.76, 0.81, 0.78, 0.78, 0.62, 0.75, 0.84, 0.92, 0.92, 0.93, 
    0.84, 0.72, 0.68, 0.73, 0.71, 0.66, 0.65, 0.62, 0.58, 0.56, 0.54, 0.61, 
    0.59, 0.58, 0.57, 0.63, 0.62, 0.66, 0.55, 0.59, 0.6, 0.52, 0.58, 0.56, 
    0.58, 0.56, 0.59, 0.62, 0.63, 0.61, 0.6, 0.58, 0.62, 0.64, 0.64, 0.59, 
    0.65, 0.64, 0.64, 0.56, 0.57, 0.55, 0.53, 0.49, 0.54, 0.54, 0.5, 0.54, 
    0.54, 0.55, 0.6, 0.61, 0.62, 0.64, 0.63, 0.62, 0.62, 0.61, 0.54, 0.56, 
    0.58, 0.57, 0.57, 0.58, 0.57, 0.57, 0.58, 0.58, 0.57, 0.59, 0.58, 0.66, 
    0.63, 0.64, 0.65, 0.65, 0.64, 0.64, 0.61, 0.59, 0.6, 0.62, 0.6, 0.58, 
    0.6, 0.59, 0.6, 0.6, 0.57, 0.59, 0.58, 0.58, 0.6, 0.64, 0.63, 0.64, 0.66, 
    0.68, 0.66, 0.67, 0.7, 0.71, 0.73, 0.7, 0.67, 0.64, 0.63, 0.61, 0.62, 
    0.67, 0.67, 0.68, 0.65, 0.67, 0.74, 0.7, 0.71, 0.72, 0.71, 0.72, 0.66, 
    0.64, 0.63, 0.6, 0.62, 0.61, 0.63, 0.62, 0.61, 0.63, 0.61, 0.56, 0.56, 
    0.58, 0.54, 0.55, 0.57, 0.53, 0.54, 0.58, 0.56, 0.6, 0.55, 0.56, 0.65, 
    0.61, 0.63, 0.7, 0.74, 0.76, 0.77, 0.71, 0.63, 0.55, 0.55, 0.54, 0.54, 
    0.53, 0.49, 0.51, 0.51, 0.59, 0.54, 0.48, 0.51, 0.57, 0.56, 0.57, 0.57, 
    0.61, 0.61, 0.65, 0.64, 0.59, 0.6, 0.58, 0.55, 0.53, 0.56, 0.58, 0.61, 
    0.57, 0.56, 0.57, 0.58, 0.58, 0.56, 0.62, 0.63, 0.63, 0.56, 0.66, 0.74, 
    0.56, 0.56, 0.6, 0.55, 0.54, 0.52, 0.55, 0.55, 0.53, 0.58, 0.58, 0.56, 
    0.55, 0.51, 0.46, 0.35, 0.33, 0.24, 0.32, 0.36, 0.37, 0.4, 0.41, 0.42, 
    0.33, 0.3, 0.29, 0.27, 0.29, 0.3, 0.27, 0.34, 0.38, 0.38, 0.36, 0.36, 
    0.36, 0.35, 0.36, 0.4, 0.36, 0.46, 0.3, 0.42, 0.46, 0.42, 0.34, 0.41, 
    0.44, 0.48, 0.71, 0.63, 0.69, 0.67, 0.62, 0.6, 0.63, 0.64, 0.66, 0.72, 
    0.66, 0.62, 0.68, 0.62, 0.66, 0.69, 0.73, 0.76, 0.73, 0.68, 0.68, 0.67, 
    0.76, 0.82, 0.83, 0.85, 0.85, 0.86, 0.74, 0.74, 0.79, 0.78, 0.81, 0.83, 
    0.78, 0.83, 0.81, 0.82, 0.81, 0.82, 0.84, 0.83, 0.82, 0.83, 0.86, 0.87, 
    0.85, 0.76, 0.74, 0.76, 0.74, 0.78, 0.81, 0.8, 0.77, 0.79, 0.85, 0.86, 
    0.86, 0.85, 0.82, 0.84, 0.81, 0.78, 0.84, 0.86, 0.88, 0.86, 0.85, 0.85, 
    0.87, 0.84, 0.8, 0.85, 0.8, 0.8, 0.77, 0.76, 0.75, 0.74, 0.77, 0.76, 
    0.75, 0.75, 0.77, 0.74, 0.73, 0.71, 0.75, 0.77, 0.72, 0.76, 0.74, 0.75, 
    0.8, 0.81, 0.83, 0.86, 0.84, 0.82, 0.82, 0.84, 0.86, 0.86, 0.89, 0.84, 
    0.86, 0.82, 0.8, 0.79, 0.73, 0.66, 0.66, 0.66, 0.75, 0.71, 0.66, 0.67, 
    0.71, 0.7, 0.7, 0.76, 0.78, 0.59, 0.45, 0.43, 0.43, 0.37, 0.37, 0.42, 
    0.41, 0.51, 0.62, 0.67, 0.59, 0.63, 0.65, 0.71, 0.77, 0.73, 0.74, 0.77, 
    0.77, 0.87, 0.88, 0.86, 0.78, 0.82, 0.83, 0.83, 0.8, 0.77, 0.78, 0.75, 
    0.74, 0.72, 0.71, 0.76, 0.81, 0.81, 0.9, 0.92, 0.93, 0.94, 0.95, 0.93, 
    0.94, 0.92, 0.93, 0.93, 0.92, 0.92, 0.93, 0.94, 0.91, 0.89, 0.88, 0.87, 
    0.85, 0.82, 0.81, 0.77, 0.76, 0.79, 0.72, 0.74, 0.73, 0.72, 0.7, 0.73, 
    0.86, 0.85, 0.88, 0.87, 0.91, 0.82, 0.76, 0.78, 0.87, 0.88, 0.84, 0.79, 
    0.84, 0.83, 0.81, 0.83, 0.75, 0.86, 0.83, 0.88, 0.86, 0.87, 0.89, 0.89, 
    0.89, 0.92, 0.91, 0.9, 0.91, 0.92, 0.9, 0.92, 0.93, 0.93, 0.92, 0.9, 0.9, 
    0.87, 0.87, 0.87, 0.87, 0.9, 0.82, 0.88, 0.8, 0.89, 0.9, 0.87, 0.89, 
    0.88, 0.93, 0.92, 0.94, 0.93, 0.91, 0.91, 0.86, 0.82, 0.82, 0.83, 0.83, 
    0.83, 0.82, 0.8, 0.78, 0.75, 0.77, 0.74, 0.75, 0.83, 0.83, 0.85, 0.88, 
    0.92, 0.92, 0.93, 0.94, 0.95, 0.86, 0.84, 0.85, 0.88, 0.93, 0.94, 0.96, 
    0.94, 0.88, 0.91, 0.9, 0.85, 0.77, 0.83, 0.84, 0.83, 0.83, 0.82, 0.81, 
    0.81, 0.8, 0.81, 0.77, 0.79, 0.78, 0.76, 0.73, 0.69, 0.7, 0.71, 0.73, 
    0.73, 0.75, 0.8, 0.86, 0.87, 0.87, 0.87, 0.87, 0.86, 0.88, 0.88, 0.9, 
    0.93, 0.95, 0.96, 0.94, 0.95, 0.96, 0.97, 0.92, 0.87, 0.77, 0.75, 0.7, 
    0.7, 0.68, 0.66, 0.65, 0.65, 0.65, 0.66, 0.66, 0.69, 0.74, 0.76, 0.76, 
    0.76, 0.8, 0.81, 0.82, 0.81, 0.83, 0.77, 0.78, 0.74, 0.74, 0.69, 0.68, 
    0.69, 0.68, 0.71, 0.74, 0.76, 0.77, 0.81, 0.79, 0.79, 0.82, 0.8, 0.85, 
    0.84, 0.84, 0.88, 0.89, 0.91, 0.89, 0.88, 0.89, 0.82, 0.79, 0.78, 0.77, 
    0.77, 0.76, 0.72, 0.7, 0.7, 0.7, 0.7, 0.71, 0.71, 0.69, 0.71, 0.72, 0.73, 
    0.74, 0.72, 0.77, 0.78, 0.8, 0.76, 0.72, 0.72, 0.63, 0.58, 0.58, 0.59, 
    0.63, 0.76, 0.82, 0.79, 0.67, 0.66, 0.69, 0.74, 0.71, 0.76, 0.81, 0.76, 
    0.79, 0.79, 0.8, 0.82, 0.79, 1, 0.77, 0.75, 0.8, 0.78, 0.76, 0.78, 0.7, 
    0.68, 0.68, 0.66, 0.68, 0.62, 0.65, 0.67, 0.69, 0.7, 0.67, 0.75, 0.77, 
    0.78, 1, 0.71, 0.77, 0.74, 0.73, 0.63, 0.67, 0.71, 0.69, 0.72, 0.57, 
    0.56, 0.58, 0.66, 0.71, 0.69, 0.7, 0.77, 0.75, 0.81, 0.75, 0.72, 0.72, 
    0.73, 0.74, 0.75, 0.72, 0.72, 0.71, 0.68, 0.71, 0.69, 0.67, 0.66, 0.64, 
    0.59, 0.59, 0.62, 0.65, 0.66, 0.61, 0.6, 0.59, 0.57, 0.57, 0.6, 0.6, 0.6, 
    0.59, 0.61, 0.64, 0.66, 0.65, 0.63, 0.63, 0.64, 0.69, 0.73, 0.59, 0.6, 
    0.58, 0.55, 0.56, 0.55, 0.54, 0.56, 0.54, 0.56, 0.69, 0.58, 0.65, 0.67, 
    0.69, 0.68, 0.69, 0.68, 0.68, 0.68, 0.69, 0.68, 0.73, 0.77, 0.66, 0.67, 
    0.66, 0.69, 0.76, 0.74, 0.73, 0.74, 0.76, 0.74, 0.76, 0.75, 0.78, 0.76, 
    0.76, 0.76, 0.76, 0.75, 0.73, 0.72, 0.71, 0.67, 0.67, 0.67, 0.65, 0.65, 
    0.6, 0.63, 0.66, 0.61, 0.71, 0.71, 0.73, 0.75, 0.7, 0.73, 0.75, 0.7, 
    0.69, 0.75, 0.71, 0.68, 0.69, 0.68, 0.65, 0.62, 0.6, 0.56, 0.59, 0.59, 
    0.59, 0.56, 0.57, 0.6, 0.61, 0.68, 0.67, 0.63, 0.63, 0.63, 0.65, 0.7, 
    0.78, 0.75, 0.7, 0.61, 0.65, 0.78, 0.79, 0.72, 0.69, 0.67, 0.67, 0.78, 
    0.65, 0.75, 0.72, 0.84, 0.88, 0.84, 0.8, 0.8, 0.78, 0.76, 0.74, 0.71, 
    0.72, 0.71, 0.69, 0.68, 0.74, 0.64, 0.67, 0.65, 0.73, 0.75, 0.67, 0.62, 
    0.64, 0.65, 0.67, 0.68, 0.7, 0.69, 0.71, 0.77, 0.75, 0.76, 0.75, 0.79, 
    0.76, 0.8, 0.81, 0.84, 0.82, 0.86, 0.84, 0.83, 0.77, 0.66, 0.65, 0.63, 
    0.62, 0.61, 0.63, 0.69, 0.76, 0.78, 0.82, 0.82, 0.83, 0.79, 0.8, 0.85, 
    0.87, 0.86, 0.88, 0.83, 0.69, 0.65, 0.64, 0.61, 0.61, 0.58, 0.57, 0.6, 
    0.65, 0.62, 0.58, 0.64, 0.64, 0.68, 0.7, 0.7, 0.68, 0.72, 0.73, 0.76, 
    0.78, 0.81, 0.79, 0.8, 0.82, 0.82, 0.81, 0.8, 0.82, 0.73, 0.68, 0.7, 
    0.72, 0.81, 0.72, 0.73, 0.7, 0.75, 0.76, 0.77, 0.76, 0.77, 0.77, 0.77, 
    0.78, 0.77, 0.77, 0.74, 0.76, 0.75, 0.75, 0.76, 0.74, 0.69, 0.72, 0.68, 
    0.67, 0.69, 0.7, 0.73, 0.65, 0.69, 0.69, 0.67, 0.65, 0.65, 0.67, 0.64, 
    0.61, 0.6, 0.59, 0.57, 0.59, 0.58, 0.58, 0.62, 0.58, 0.55, 0.53, 0.53, 
    0.49, 0.49, 0.48, 0.49, 0.49, 0.5, 0.52, 0.48, 0.48, 0.54, 0.6, 0.64, 
    0.64, 0.64, 0.64, 0.64, 0.63, 0.64, 0.7, 0.66, 0.61, 0.67, 0.63, 0.54, 
    0.55, 0.55, 0.58, 0.56, 0.52, 0.52, 0.52, 0.52, 0.53, 0.57, 0.59, 0.6, 
    0.61, 0.61, 0.56, 0.6, 0.58, 0.54, 0.54, 0.54, 0.57, 0.57, 0.56, 0.54, 
    0.5, 0.49, 0.5, 0.48, 0.49, 0.5, 0.51, 0.53, 0.51, 0.53, 0.53, 0.52, 
    0.55, 0.58, 0.61, 0.6, 0.58, 0.62, 0.59, 0.59, 0.58, 0.59, 0.6, 0.59, 
    0.62, 0.59, 0.62, 0.68, 0.71, 0.71, 0.73, 0.75, 0.75, 0.74, 0.77, 0.78, 
    0.79, 0.79, 0.79, 0.8, 0.79, 0.77, 0.73, 0.63, 0.63, 0.61, 0.61, 0.6, 
    0.59, 0.57, 0.62, 0.64, 0.66, 0.71, 0.67, 0.72, 0.71, 0.72, 0.71, 0.73, 
    0.7, 0.71, 0.68, 0.75, 0.7, 0.65, 0.65, 0.67, 0.68, 0.64, 0.67, 0.7, 
    0.66, 0.65, 0.69, 0.74, 0.77, 0.77, 0.77, 0.78, 0.77, 0.77, 0.81, 0.74, 
    0.78, 0.77, 0.77, 0.78, 0.8, 0.78, 0.79, 0.75, 0.73, 0.77, 0.79, 0.75, 
    0.74, 0.75, 0.75, 0.71, 0.73, 0.74, 0.74, 0.78, 0.78, 0.77, 0.78, 0.78, 
    0.79, 0.78, 0.83, 0.81, 0.79, 0.76, 0.71, 0.67, 0.68, 0.69, 0.7, 0.72, 
    0.69, 0.67, 0.68, 0.71, 0.74, 0.72, 0.72, 0.74, 0.72, 0.73, 0.74, 0.75, 
    0.76, 0.78, 0.77, 0.76, 0.75, 0.79, 0.73, 0.77, 0.73, 0.72, 0.71, 0.7, 
    0.67, 0.63, 0.66, 0.63, 0.67, 0.64, 0.65, 0.66, 0.68, 0.69, 0.7, 0.7, 
    0.67, 0.69, 0.68, 0.66, 0.71, 0.69, 0.66, 0.67, 0.68, 0.64, 0.65, 0.64, 
    0.61, 0.6, 0.58, 0.57, 0.64, 0.75, 0.77, 0.78, 0.82, 0.86, 0.84, 0.74, 
    0.73, 0.82, 0.8, 0.76, 0.78, 0.72, 0.72, 0.72, 0.72, 0.75, 0.69, 0.69, 
    0.71, 0.74, 0.72, 0.71, 0.7, 0.73, 0.73, 0.79, 0.79, 0.77, 0.82, 0.75, 
    0.79, 0.84, 0.76, 0.79, 0.78, 0.78, 0.72, 0.67, 0.7, 0.7, 0.69, 0.64, 
    0.6, 0.71, 0.76, 0.77, 0.69, 0.75, 0.81, 0.75, 0.75, 0.78, 0.81, 0.77, 
    0.77, 0.82, 0.84, 0.86, 0.87, 0.88, 0.9, 0.92, 0.92, 0.92, 0.92, 0.91, 
    0.89, 0.85, 0.86, 0.86, 0.85, 0.85, 0.82, 0.85, 0.75, 0.76, 0.76, 0.79, 
    0.8, 0.81, 0.79, 0.78, 0.78, 0.74, 0.74, 0.73, 0.76, 0.77, 0.81, 0.84, 
    0.82, 0.8, 0.79, 0.81, 0.77, 0.76, 0.73, 0.72, 0.76, 0.8, 0.81, 0.79, 
    0.8, 0.79, 0.77, 0.83, 0.84, 0.82, 0.89, 0.83, 0.85, 0.86, 0.83, 0.84, 
    0.87, 0.84, 0.85, 0.83, 0.82, 0.83, 0.8, 0.79, 0.79, 0.77, 0.79, 0.76, 
    0.74, 0.76, 0.65, 0.63, 0.58, 0.53, 0.58, 0.58, 0.66, 0.75, 0.75, 0.77, 
    0.73, 0.71, 0.82, 0.8, 0.8, 0.81, 0.79, 0.8, 0.78, 0.78, 0.8, 0.79, 0.81, 
    0.84, 0.75, 0.72, 0.71, 0.72, 0.74, 0.71, 0.64, 0.64, 0.6, 0.68, 0.7, 
    0.69, 0.66, 0.69, 0.66, 0.69, 0.63, 0.65, 0.67, 0.68, 0.68, 0.69, 0.69, 
    0.82, 0.73, 0.74, 0.76, 0.78, 0.74, 0.79, 0.75, 0.75, 0.78, 0.78, 0.86, 
    0.85, 0.89, 0.86, 0.89, 0.9, 0.93, 0.95, 0.94, 0.92, 0.93, 0.93, 0.9, 
    0.87, 0.93, 0.94, 0.95, 0.96, 0.96, 0.95, 0.94, 0.92, 0.92, 0.95, 0.97, 
    0.97, 0.96, 0.96, 0.93, 0.85, 0.84, 0.84, 0.85, 0.86, 0.85, 0.84, 0.81, 
    0.82, 0.89, 0.87, 0.9, 0.89, 0.88, 0.84, 0.84, 0.82, 0.85, 0.84, 0.85, 
    0.82, 0.82, 0.85, 0.93, 0.95, 0.91, 0.89, 0.88, 0.86, 0.82, 0.85, 0.86, 
    0.83, 0.87, 0.9, 0.91, 0.85, 0.81, 0.82, 0.8, 0.78, 0.8, 0.79, 0.81, 0.8, 
    0.81, 0.78, 0.84, 0.82, 0.87, 0.89, 0.87, 0.85, 0.82, 0.8, 0.82, 0.82, 
    0.83, 0.79, 0.84, 0.84, 0.86, 0.85, 0.84, 0.84, 0.82, 0.83, 0.85, 0.85, 
    0.85, 0.83, 0.8, 0.76, 0.75, 0.77, 0.77, 0.77, 0.82, 0.8, 0.83, 0.8, 
    0.74, 0.75, 0.75, 0.76, 0.77, 0.75, 0.73, 0.72, 0.68, 0.81, 0.82, 0.69, 
    0.75, 0.66, 0.72, 0.81, 1, 0.81, 0.82, 0.85, 0.83, 0.84, 0.85, 0.83, 
    0.82, 0.79, 0.76, 0.78, 0.77, 0.79, 0.79, 0.75, 0.78, 0.77, 0.73, 0.74, 
    0.76, 0.76, 0.79, 0.79, 0.83, 0.84, 1, 0.82, 0.85, 0.82, 0.82, 0.82, 
    0.84, 0.86, 0.86, 0.87, 0.86, 0.86, 0.85, 0.8, 0.83, 0.82, 0.81, 0.81, 
    0.78, 0.8, 0.77, 0.77, 0.8, 0.82, 0.89, 0.8, 0.84, 0.84, 0.84, 0.84, 
    0.81, 0.89, 0.91, 0.89, 0.87, 0.85, 0.77, 0.71, 0.69, 0.67, 0.74, 0.77, 
    0.78, 0.71, 0.71, 0.67, 0.66, 0.65, 0.66, 0.68, 0.73, 0.68, 0.74, 0.76, 
    0.82, 0.76, 0.72, 0.7, 0.73, 0.68, 0.75, 0.85, 0.63, 0.61, 0.76, 0.76, 
    0.68, 0.67, 0.7, 0.72, 0.74, 1, 1, 0.9, 0.74, 0.75, 0.73, 0.72, 0.7, 0.7, 
    0.69, 0.66, 0.69, 0.7, 0.65, 0.64, 0.67, 0.65, 0.65, 0.62, 0.6, 0.61, 
    0.59, 0.62, 0.66, 0.66, 0.58, 0.61, 0.66, 0.68, 0.67, 0.69, 0.67, 0.62, 
    0.64, 0.63, 0.64, 0.64, 0.63, 0.63, 0.62, 0.63, 0.61, 0.61, 0.59, 0.58, 
    0.61, 0.61, 0.63, 0.64, 0.65, 0.65, 0.68, 0.7, 0.7, 0.7, 0.66, 0.67, 
    0.67, 0.69, 0.71, 0.7, 0.75, 0.76, 0.76, 0.75, 0.76, 0.74, 0.66, 0.68, 
    0.71, 0.73, 0.78, 0.77, 0.66, 0.67, 0.66, 0.66, 0.62, 0.62, 0.66, 0.67, 
    0.78, 0.75, 0.72, 0.77, 0.77, 0.72, 0.72, 0.72, 0.76, 0.84, 0.84, 0.8, 
    0.84, 0.79, 0.82, 0.88, 0.86, 0.91, 0.96, 0.94, 0.89, 0.88, 0.89, 0.9, 
    0.9, 0.91, 0.89, 0.88, 0.88, 0.86, 0.84, 0.89, 0.86, 0.81, 0.78, 0.79, 
    0.79, 0.78, 0.77, 0.76, 0.76, 0.79, 0.77, 0.77, 0.77, 0.72, 0.69, 0.64, 
    0.65, 0.6, 0.6, 0.61, 0.61, 0.68, 0.68, 0.67, 0.52, 0.7, 0.68, 0.54, 
    0.54, 0.56, 0.57, 0.59, 0.63, 0.65, 0.72, 0.72, 0.76, 0.75, 0.75, 0.74, 
    0.74, 0.78, 0.78, 0.76, 0.79, 0.77, 0.76, 0.77, 0.72, 0.73, 0.72, 0.66, 
    0.68, 0.76, 0.81, 0.71, 0.76, 0.82, 0.82, 0.81, 0.86, 0.93, 0.9, 0.91, 
    0.84, 0.8, 0.78, 0.78, 0.75, 0.76, 0.75, 0.75, 0.73, 0.74, 0.76, 0.76, 
    0.76, 0.83, 0.82, 0.8, 0.76, 0.74, 0.75, 0.77, 0.77, 0.76, 0.75, 0.69, 
    0.71, 0.72, 0.71, 0.68, 0.71, 0.71, 0.73, 0.72, 0.71, 0.72, 0.7, 0.71, 
    0.73, 0.7, 0.66, 0.69, 0.68, 0.67, 0.7, 0.77, 0.75, 0.75, 0.77, 0.8, 
    0.73, 0.7, 0.69, 0.68, 0.79, 0.74, 0.76, 0.75, 0.79, 0.76, 0.82, 0.77, 
    0.82, 0.84, 0.81, 0.79, 0.82, 0.86, 0.97, 0.97, 1, 1, 1, 1, 0.93, 0.89, 
    0.86, 0.93, 0.94, 0.98, 1, 1, 0.91, 0.84, 0.84, 0.77, 0.85, 0.8, 0.78, 
    0.75, 0.74, 0.74, 0.73, 0.74, 0.73, 0.71, 0.72, 0.72, 0.7, 0.71, 0.69, 
    0.67, 0.62, 0.63, 0.64, 0.63, 0.6, 0.6, 0.66, 0.63, 0.59, 0.61, 0.63, 
    0.64, 0.65, 0.68, 0.68, 0.69, 0.7, 0.7, 0.71, 0.72, 0.71, 0.71, 0.71, 
    0.69, 0.66, 0.73, 0.72, 0.73, 0.72, 0.72, 0.72, 0.71, 0.71, 0.69, 0.7, 
    0.7, 0.76, 0.73, 0.77, 0.72, 0.7, 0.77, 0.76, 0.76, 0.78, 0.75, 0.76, 
    0.81, 0.8, 0.94, 0.96, 0.99, 0.95, 0.94, 0.97, 1, 0.92, 0.95, 0.96, 0.96, 
    1, 0.97, 0.9, 0.74, 0.73, 0.73, 0.68, 0.69, 0.65, 0.65, 0.65, 0.65, 0.65, 
    0.65, 0.64, 0.66, 0.64, 0.68, 0.63, 0.62, 0.6, 0.59, 0.59, 0.59, 0.64, 
    0.65, 0.66, 0.67, 0.67, 0.65, 0.63, 0.56, 0.64, 0.63, 0.58, 0.61, 0.66, 
    0.64, 0.61, 0.65, 0.64, 0.55, 0.68, 0.67, 0.66, 0.64, 0.66, 0.61, 0.65, 
    0.66, 0.68, 0.69, 0.66, 0.72, 0.68, 0.65, 0.65, 0.66, 0.71, 0.69, 0.65, 
    0.63, 0.62, 0.64, 0.62, 0.62, 0.66, 0.67, 0.63, 0.64, 0.67, 0.68, 0.68, 
    0.62, 0.74, 0.71, 0.75, 0.76, 0.76, 0.77, 0.79, 0.74, 0.72, 0.73, 0.68, 
    0.76, 0.73, 0.84, 0.73, 0.74, 0.73, 0.74, 0.76, 0.76, 0.77, 0.75, 0.77, 
    0.76, 0.77, 0.78, 0.8, 0.82, 0.82, 0.82, 0.96, 1, 0.97, 0.96, 1, 0.89, 
    0.94, 1, 0.99, 0.97, 0.95, 0.85, 0.82, 0.79, 0.8, 0.8, 0.82, 0.82, 0.87, 
    0.77, 0.84, 0.85, 0.82, 0.78, 0.86, 0.97, 1, 1, 0.93, 0.86, 0.79, 0.71, 
    0.59, 0.58, 0.61, 0.58, 0.58, 0.63, 0.63, 0.62, 0.6, 0.63, 0.65, 0.66, 
    0.66, 0.64, 0.63, 0.6, 0.57, 0.56, 0.53, 0.53, 0.52, 0.51, 0.53, 0.54, 
    0.54, 0.53, 0.55, 0.56, 0.55, 0.57, 0.58, 0.6, 0.61, 0.61, 0.62, 0.63, 
    0.64, 0.62, 0.63, 0.6, 0.65, 0.67, 0.67, 0.72, 0.68, 0.64, 0.62, 0.66, 
    0.6, 0.61, 0.61, 0.6, 0.58, 0.6, 0.62, 0.64, 0.65, 0.66, 0.66, 0.71, 0.7, 
    0.72, 0.76, 0.78, 0.75, 0.74, 0.72, 0.73, 0.74, 0.76, 0.73, 0.76, 0.74, 
    0.66, 0.59, 0.6, 0.55, 0.56, 0.53, 0.53, 0.55, 0.59, 0.6, 0.6, 0.59, 0.6, 
    0.61, 0.61, 0.6, 0.57, 0.61, 0.59, 0.59, 0.65, 0.68, 0.66, 0.65, 0.66, 
    0.67, 0.64, 0.64, 0.65, 0.64, 0.68, 0.7, 0.74, 0.76, 0.81, 0.82, 0.85, 
    0.84, 0.83, 0.78, 0.76, 0.76, 0.7, 0.75, 0.74, 0.74, 0.72, 0.68, 0.69, 
    0.7, 0.64, 0.67, 0.58, 0.45, 0.46, 0.46, 0.49, 0.44, 0.47, 0.48, 0.53, 
    0.61, 0.66, 0.63, 0.64, 0.69, 0.71, 0.68, 0.71, 0.68, 0.67, 0.65, 0.67, 
    0.67, 0.63, 0.62, 0.62, 0.66, 0.7, 0.72, 0.76, 0.76, 0.77, 0.79, 0.8, 
    0.79, 0.8, 0.81, 0.79, 0.79, 0.75, 0.73, 0.73, 0.78, 0.76, 0.75, 0.74, 
    0.68, 0.68, 0.71, 0.79, 0.78, 0.76, 0.79, 0.77, 0.75, 0.7, 0.72, 0.7, 
    0.74, 0.73, 0.87, 0.97, 0.95, 0.92, 0.95, 0.85, 0.83, 0.82, 0.76, 0.73, 
    0.82, 0.98, 0.95, 0.88, 0.82, 0.9, 0.95, 0.94, 0.93, 0.87, 0.91, 0.87, 
    0.93, 0.92, 0.92, 0.94, 1, 1, 0.85, 0.99, 0.95, 1, 0.99, 0.93, 0.78, 
    0.81, 0.77, 0.82, 0.82, 0.74, 0.72, 0.77, 0.78, 0.79, 0.79, 0.78, 0.73, 
    0.76, 0.69, 0.68, 0.64, 0.63, 0.63, 0.64, 0.61, 0.59, 0.6, 0.55, 0.56, 
    0.56, 0.6, 0.57, 0.59, 0.61, 0.61, 0.69, 0.69, 0.7, 0.7, 0.72, 0.74, 
    0.75, 0.75, 0.74, 0.75, 0.79, 0.95, 0.9, 0.74, 0.72, 0.8, 0.8, 0.77, 
    0.83, 0.8, 0.76, 0.78, 0.8, 0.84, 0.87, 0.82, 0.77, 0.79, 0.73, 0.75, 
    0.78, 0.79, 0.79, 0.75, 0.71, 0.69, 0.66, 0.68, 0.67, 0.68, 0.69, 0.71, 
    0.73, 0.79, 0.84, 0.85, 0.86, 0.89, 1, 0.89, 1, 1, 1, 1, 1, 1, 1, 0.94, 
    0.99, 0.92, 1, 0.96, 0.92, 0.88, 0.82, 0.87, 0.85, 0.85, 0.75, 0.68, 
    0.68, 0.66, 0.75, 0.73, 0.85, 0.84, 0.91, 0.89, 0.87, 0.82, 0.84, 0.76, 
    0.78, 0.78, 0.78, 0.73, 0.69, 0.73, 0.69, 0.68, 0.67, 0.66, 0.65, 0.66, 
    0.65, 0.64, 0.64, 0.64, 0.66, 0.64, 0.64, 0.63, 0.58, 0.61, 0.59, 0.6, 
    0.57, 0.56, 0.6, 0.64, 0.62, 0.6, 0.61, 0.6, 0.58, 0.6, 0.61, 0.67, 0.67, 
    0.7, 0.75, 0.77, 0.78, 0.77, 0.79, 0.75, 0.75, 0.72, 0.67, 0.65, 0.67, 
    0.7, 0.7, 0.71, 0.68, 0.69, 0.71, 0.71, 0.71, 0.71, 0.75, 0.77, 0.78, 
    0.8, 0.79, 0.81, 0.81, 0.83, 0.84, 0.83, 0.82, 0.79, 0.79, 0.79, 0.82, 
    0.8, 0.84, 0.8, 0.8, 0.93, 0.95, 0.96, 0.87, 0.83, 0.86, 0.79, 0.75, 
    0.75, 0.73, 0.76, 0.77, 0.76, 0.76, 0.74, 0.78, 0.93, 0.9, 0.84, 0.85, 
    0.87, 0.93, 0.91, 0.86, 0.8, 0.81, 0.79, 0.89, 1, 0.85, 0.79, 0.77, 0.78, 
    0.74, 0.73, 0.75, 0.74, 0.76, 0.75, 0.75, 0.74, 0.75, 0.71, 0.71, 0.72, 
    0.69, 0.71, 0.69, 0.69, 0.7, 0.72, 0.67, 0.67, 0.7, 0.74, 0.78, 0.8, 
    0.85, 0.89, 0.88, 0.92, 0.82, 0.85, 0.87, 0.82, 0.81, 0.82, 0.82, 0.81, 
    0.83, 0.81, 0.81, 0.79, 0.75, 0.75, 0.83, 0.87, 0.83, 0.96, 0.89, 0.96, 
    0.94, 0.98, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.91, 0.9, 0.9, 0.79, 0.73, 
    0.67, 0.67, 0.7, 0.63, 0.63, 0.58, 0.63, 0.63, 0.59, 0.58, 0.67, 0.7, 
    0.71, 0.63, 0.69, 0.68, 0.67, 0.73, 0.74, 0.74, 0.7, 0.66, 0.69, 0.69, 
    0.71, 0.65, 0.68, 0.68, 0.69, 0.69, 0.72, 0.75, 0.76, 0.8, 0.84, 0.9, 
    0.87, 0.9, 0.96, 0.96, 0.96, 0.93, 0.9, 0.81, 0.89, 0.88, 0.85, 0.83, 
    0.84, 0.86, 0.89, 0.96, 0.94, 0.88, 0.88, 0.89, 0.93, 1, 0.97, 1, 0.98, 
    1, 1, 1, 1, 0.99, 0.98, 1, 1, 1, 1, 0.95, 1, 0.92, 0.92, 0.95, 0.98, 1, 
    1, 1, 0.96, 0.95, 0.92, 0.87, 0.81, 0.77, 0.83, 0.77, 0.76, 0.76, 0.71, 
    0.69, 0.66, 0.62, 0.62, 0.61, 0.6, 0.64, 0.65, 0.68, 0.69, 0.68, 0.7, 
    0.65, 0.69, 0.64, 0.64, 0.66, 0.65, 0.67, 0.66, 0.65, 0.62, 0.65, 0.65, 
    0.66, 0.62, 0.61, 0.61, 0.59, 0.62, 0.64, 0.65, 0.64, 0.7, 0.7, 0.62, 
    0.64, 0.65, 0.63, 0.63, 0.65, 0.66, 0.65, 0.64, 0.65, 0.63, 0.62, 0.61, 
    0.61, 0.62, 0.62, 0.62, 0.63, 0.67, 0.61, 0.62, 0.64, 0.63, 0.61, 0.64, 
    0.64, 0.6, 0.61, 0.63, 0.61, 0.63, 0.63, 0.63, 0.63, 0.65, 0.61, 0.59, 
    0.59, 0.62, 0.63, 0.64, 0.64, 0.64, 0.66, 0.68, 0.71, 0.73, 0.7, 0.63, 
    0.66, 0.72, 0.74, 0.67, 0.63, 0.65, 0.66, 0.62, 0.63, 0.59, 0.58, 0.62, 
    0.63, 0.56, 0.62, 0.68, 0.62, 0.62, 0.64, 0.66, 0.75, 0.79, 0.79, 0.69, 
    0.71, 0.71, 0.71, 0.74, 0.72, 0.69, 0.71, 0.73, 0.74, 0.73, 0.75, 0.76, 
    0.64, 0.7, 0.68, 0.65, 0.63, 0.65, 0.69, 0.73, 0.75, 0.77, 0.8, 0.81, 
    0.85, 0.83, 0.83, 0.85, 0.85, 0.81, 0.83, 0.8, 0.77, 0.77, 0.76, 0.76, 
    0.76, 0.82, 0.8, 0.78, 0.77, 0.78, 0.93, 1, 1, 1, 0.99, 1, 1, 1, 1, 0.99, 
    0.97, 1, 0.98, 0.93, 0.95, 0.95, 0.92, 0.88, 0.88, 0.84, 0.79, 0.77, 
    0.85, 0.81, 0.83, 0.89, 0.92, 0.95, 0.93, 0.92, 0.89, 0.9, 0.95, 0.93, 
    0.94, 0.96, 0.93, 0.96, 0.93, 0.9, 0.92, 0.9, 0.83, 0.81, 0.82, 0.97, 1, 
    0.99, 0.89, 0.79, 0.79, 0.81, 0.81, 0.86, 0.95, 0.89, 0.91, 0.9, 0.91, 
    0.89, 0.92, 0.93, 0.95, 0.87, 0.89, 0.87, 0.82, 0.93, 0.91, 0.77, 0.72, 
    0.7, 0.71, 0.64, 0.64, 0.65, 0.66, 0.65, 0.59, 0.6, 0.65, 0.65, 0.66, 
    0.65, 0.64, 0.7, 0.68, 0.7, 0.73, 0.66, 0.68, 0.69, 0.7, 0.7, 0.7, 0.7, 
    0.74, 0.71, 0.71, 0.75, 0.8, 0.81, 0.8, 0.79, 0.84, 0.88, 0.9, 0.91, 
    0.89, 0.91, 0.87, 0.85, 0.81, 0.81, 0.81, 0.83, 0.81, 0.85, 0.85, 0.85, 
    0.87, 0.85, 0.88, 0.89, 0.93, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0.99, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.94, 0.94, 
    0.98, 0.94, 1, 1, 0.8, 0.79, 0.74, 0.77, 0.78, 0.74, 0.74, 0.71, 0.72, 
    0.74, 0.75, 0.73, 0.71, 0.71, 0.75, 0.76, 0.78, 0.8, 0.82, 0.88, 0.95, 
    0.96, 0.97, 0.97, 0.87, 0.9, 0.94, 0.94, 1, 1, 1, 1, 1, 1, 0.99, 0.89, 
    0.92, 0.86, 0.91, 0.89, 0.88, 0.97, 0.99, 1, 1, 1, 1, 1, 1, 1, 0.95, 
    0.95, 1, 1, 1, 1, 0.86, 0.89, 0.86, 0.84, 0.86, 0.82, 0.89, 0.83, 0.73, 
    0.75, 0.77, 0.77, 0.74, 0.73, 0.73, 0.74, 0.77, 0.81, 0.8, 0.85, 0.85, 
    0.85, 0.85, 0.86, 0.86, 0.85, 0.86, 0.88, 0.88, 0.85, 0.82, 0.84, 0.84, 
    0.83, 0.86, 0.84, 0.84, 0.83, 0.81, 0.8, 0.86, 0.84, 0.78, 0.82, 0.87, 
    0.93, 0.93, 0.96, 1, 1, 1, 1, 0.88, 0.85, 0.87, 0.86, 0.94, 0.91, 0.86, 
    0.87, 0.88, 1, 1, 0.93, 0.91, 0.94, 0.94, 0.95, 0.96, 0.94, 0.96, 0.92, 
    0.94, 1, 1, 0.93, 0.92, 0.93, 0.9, 0.84, 0.87, 0.89, 0.98, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.98, 1, 1, 1, 0.9, 1, 1, 1, 1, 0.99, 0.94, 0.98, 0.97, 0.94, 
    0.96, 0.87, 0.9, 0.98, 0.9, 0.88, 0.92, 0.8, 0.88, 0.89, 0.85, 0.84, 
    0.89, 0.9, 0.93, 0.95, 0.92, 0.87, 0.89, 0.81, 0.87, 0.89, 0.95, 0.99, 1, 
    1, 0.96, 0.96, 0.94, 0.95, 0.88, 0.86, 0.79, 0.78, 0.73, 0.75, 0.75, 
    0.76, 0.74, 0.76, 0.71, 0.7, 0.71, 0.72, 0.72, 0.7, 0.72, 0.72, 0.7, 
    0.74, 0.75, 0.74, 0.73, 0.63, 0.63, 0.61, 0.6, 0.6, 0.58, 0.59, 0.61, 
    0.61, 0.61, 0.66, 0.66, 0.63, 0.64, 0.65, 0.65, 0.64, 0.66, 0.69, 0.64, 
    0.64, 0.71, 0.73, 0.71, 0.74, 0.7, 0.69, 0.65, 0.62, 0.59, 0.69, 0.65, 
    0.65, 0.64, 0.69, 0.68, 0.68, 0.7, 0.73, 0.71, 0.75, 0.77, 0.8, 0.8, 
    0.75, 0.76, 0.77, 0.74, 0.75, 0.8, 0.76, 0.79, 0.76, 0.72, 0.73, 0.74, 
    0.7, 0.74, 0.69, 0.75, 0.79, 0.76, 0.73, 0.68, 0.71, 0.74, 0.77, 0.78, 
    0.73, 0.73, 0.74, 0.74, 0.79, 0.81, 0.9, 0.94, 0.94, 0.94, 0.91, 0.93, 
    0.94, 0.94, 0.94, 0.97, 0.98, 0.99, 1, 1, 1, 0.99, 1, 1, 1, 1, 1, 1, 
    0.95, 1, 1, 1, 1, 1, 0.98, 0.84, 0.88, 0.82, 0.89, 0.95, 0.96, 1, 1, 1, 
    1, 1, 1, 0.98, 0.9, 0.89, 0.91, 0.95, 0.96, 0.86, 0.84, 0.9, 0.9, 0.95, 
    1, 0.98, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.99, 0.93, 1, 0.98, 1, 
    1, 1, 1, 0.98, 0.93, 0.98, 0.98, 1, 0.98, 0.98, 0.98, 1, 1, 0.98, 0.98, 
    0.98, 0.96, 0.9, 0.94, 0.82, 0.79, 0.76, 0.77, 0.72, 0.78, 0.79, 0.77, 
    0.72, 0.69, 0.69, 0.7, 0.72, 0.75, 0.69, 0.79, 0.7, 0.7, 0.65, 0.67, 
    0.67, 0.67, 0.72, 0.73, 0.74, 0.69, 0.69, 0.7, 0.71, 0.71, 0.71, 0.72, 
    0.71, 0.68, 0.66, 0.67, 0.67, 0.65, 0.67, 0.67, 0.69, 0.69, 0.66, 0.67, 
    0.67, 0.68, 0.68, 0.68, 0.69, 0.7, 0.74, 0.7, 0.7, 0.72, 0.7, 0.73, 0.76, 
    0.76, 0.77, 0.71, 0.74, 0.71, 0.73, 0.74, 0.73, 0.73, 0.75, 0.73, 0.71, 
    0.72, 0.69, 0.74, 0.72, 0.73, 0.74, 0.74, 0.73, 0.72, 0.68, 0.72, 0.71, 
    0.69, 0.7, 0.68, 0.71, 0.69, 0.67, 0.72, 0.71, 0.72, 0.7, 0.71, 0.71, 
    0.75, 0.7, 0.76, 0.71, 0.75, 0.73, 0.71, 0.73, 0.7, 0.72, 0.66, 0.64, 
    0.71, 0.63, 0.6, 0.62, 0.66, 0.66, 0.65, 0.63, 0.61, 0.68, 0.59, 0.55, 
    0.61, 0.63, 0.66, 0.67, 0.66, 0.62, 0.72, 0.76, 0.86, 0.87, 0.83, 0.82, 
    0.78, 0.74, 0.75, 0.74, 0.74, 0.69, 0.69, 0.76, 0.76, 0.74, 0.8, 0.7, 
    0.65, 0.67, 0.64, 0.64, 0.58, 0.55, 0.61, 0.6, 0.64, 0.63, 0.61, 0.61, 
    0.61, 0.62, 0.67, 0.65, 0.71, 0.73, 0.72, 0.66, 0.68, 0.72, 0.79, 0.73, 
    0.76, 0.74, 0.79, 0.77, 0.79, 0.79, 0.79, 0.79, 0.79, 0.77, 0.77, 0.76, 
    0.78, 0.81, 0.79, 0.8, 0.81, 0.83, 0.87, 0.9, 0.92, 0.9, 0.87, 0.89, 
    0.87, 0.86, 0.96, 0.97, 0.96, 0.93, 0.91, 0.88, 0.86, 0.88, 0.87, 0.86, 
    0.81, 0.82, 0.85, 0.82, 0.85, 0.81, 0.86, 0.78, 0.78, 0.72, 0.67, 0.76, 
    0.77, 0.78, 0.78, 0.81, 0.88, 0.95, 0.97, 0.99, 1, 0.94, 0.94, 0.98, 
    0.97, 1, 0.97, 1, 1, 1, 1, 1, 1, 0.98, 0.98, 0.95, 0.95, 0.86, 0.84, 
    0.85, 0.89, 0.85, 0.85, 0.94, 0.96, 0.97, 1, 1, 1, 0.93, 1, 1, 1, 1, 
    0.98, 0.85, 0.81, 0.85, 0.86, 0.97, 1, 0.91, 0.93, 0.93, 0.92, 0.89, 
    0.92, 0.95, 0.93, 0.79, 0.79, 0.84, 0.88, 0.89, 0.83, 0.79, 0.83, 0.92, 
    0.89, 0.76, 0.74, 0.72, 0.72, 0.74, 0.76, 0.74, 0.7, 0.72, 0.71, 0.71, 
    0.68, 0.69, 0.71, 0.75, 0.8, 0.84, 0.79, 0.82, 0.87, 0.89, 0.86, 0.69, 
    0.68, 0.67, 0.66, 0.67, 0.69, 0.69, 0.66, 0.7, 0.66, 0.65, 0.66, 0.66, 
    0.67, 0.67, 0.7, 0.67, 0.69, 0.71, 0.69, 0.68, 0.67, 0.7, 0.67, 0.68, 
    0.7, 0.68, 0.68, 0.7, 0.72, 0.72, 0.7, 0.73, 0.71, 0.72, 0.7, 0.74, 0.74, 
    0.73, 0.73, 0.73, 0.69, 0.71, 0.75, 0.87, 0.94, 0.98, 0.98, 0.94, 0.94, 
    0.66, 0.66, 0.64, 0.6, 0.6, 0.57, 0.56, 0.53, 0.53, 0.57, 0.57, 0.57, 
    0.56, 0.51, 0.52, 0.52, 0.52, 0.5, 0.47, 0.47, 0.49, 0.5, 0.48, 0.48, 
    0.5, 0.49, 0.49, 0.49, 0.47, 0.5, 0.52, 0.53, 0.55, 0.6, 0.71, 0.74, 
    0.77, 0.89, 0.91, 0.57, 0.5, 0.51, 0.53, 0.55, 0.52, 0.52, 0.55, 0.62, 
    0.64, 0.62, 0.57, 0.54, 0.55, 0.57, 0.51, 0.53, 0.56, 0.56, 0.54, 0.53, 
    0.55, 0.53, 0.48, 0.48, 0.47, 0.42, 0.42, 0.43, 0.45, 0.47, 0.5, 0.49, 
    0.52, 0.46, 0.48, 0.51, 0.49, 0.49, 0.49, 0.49, 0.48, 0.5, 0.48, 0.46, 
    0.46, 0.48, 0.5, 0.53, 0.54, 0.52, 0.57, 0.51, 0.5, 0.49, 0.55, 0.53, 
    0.5, 0.52, 0.54, 0.55, 0.54, 0.55, 0.54, 0.54, 0.62, 0.53, 0.54, 0.6, 
    0.62, 0.65, 0.66, 0.7, 0.67, 0.67, 0.66, 0.65, 0.62, 0.6, 0.66, 0.67, 
    0.64, 0.67, 0.67, 0.7, 0.72, 0.71, 0.74, 0.77, 0.7, 0.75, 0.74, 0.73, 
    0.71, 0.69, 0.7, 0.71, 0.69, 0.73, 0.76, 0.74, 0.72, 0.74, 0.75, 0.72, 
    0.72, 0.7, 0.71, 0.61, 0.63, 0.62, 0.61, 0.57, 0.55, 0.56, 0.56, 0.56, 
    0.55, 0.52, 0.53, 0.52, 0.53, 0.54, 0.52, 0.59, 0.63, 0.61, 0.61, 0.54, 
    0.59, 0.58, 0.58, 0.62, 0.59, 0.59, 0.56, 0.58, 0.58, 0.56, 0.55, 0.53, 
    0.54, 0.54, 0.58, 0.6, 0.6, 0.62, 0.6, 0.61, 0.56, 0.5, 0.46, 0.48, 0.5, 
    0.52, 0.53, 0.52, 0.58, 0.6, 0.58, 0.59, 0.59, 0.61, 0.6, 0.56, 0.62, 
    0.61, 0.54, 0.54, 0.56, 0.56, 0.55, 0.59, 0.52, 0.53, 0.49, 0.49, 0.47, 
    0.46, 0.46, 0.58, 0.6, 0.56, 0.54, 0.5, 0.49, 0.47, 0.45, 0.51, 0.48, 
    0.51, 0.53, 0.55, 0.56, 0.55, 0.57, 0.56, 0.56, 0.59, 0.6, 0.62, 0.64, 
    0.66, 0.67, 0.7, 0.69, 0.7, 0.7, 0.66, 0.68, 0.7, 0.72, 0.74, 0.73, 0.73, 
    0.73, 0.74, 0.7, 0.72, 0.73, 0.75, 0.76, 0.76, 0.7, 0.7, 0.69, 0.67, 
    0.69, 0.76, 0.78, 0.77, 0.78, 0.77, 0.77, 0.77, 0.78, 0.77, 0.78, 0.77, 
    0.79, 0.76, 0.72, 0.69, 0.69, 0.67, 0.67, 0.69, 0.67, 0.69, 0.67, 0.57, 
    0.54, 0.6, 0.58, 0.57, 0.6, 0.61, 0.61, 0.59, 0.66, 0.68, 0.57, 0.63, 
    0.62, 0.59, 0.61, 0.56, 0.6, 0.62, 0.63, 0.6, 0.63, 0.71, 0.69, 0.76, 
    0.75, 0.68, 0.62, 0.68, 0.61, 0.62, 0.59, 0.63, 0.54, 0.53, 0.59, 0.53, 
    0.52, 0.53, 0.54, 0.54, 0.55, 0.54, 0.55, 0.58, 0.56, 0.52, 0.5, 0.53, 
    0.52, 0.57, 0.58, 0.56, 0.58, 0.65, 0.63, 0.65, 0.63, 0.62, 0.57, 0.51, 
    0.57, 0.66, 0.67, 0.73, 0.63, 0.57, 0.56, 0.56, 0.58, 0.54, 0.5, 0.49, 
    0.49, 0.48, 0.49, 0.47, 0.52, 0.5, 0.49, 0.52, 0.56, 0.58, 0.59, 0.54, 
    0.55, 0.55, 0.53, 0.55, 0.54, 0.53, 0.54, 0.53, 0.49, 0.5, 0.5, 0.5, 
    0.49, 0.49, 0.49, 0.5, 0.49, 0.46, 0.45, 0.46, 0.46, 0.45, 0.46, 0.5, 
    0.51, 0.53, 0.63, 0.56, 0.56, 0.59, 0.63, 0.68, 0.68, 0.66, 0.67, 0.66, 
    0.67, 0.73, 0.71, 0.76, 0.74, 0.73, 0.76, 0.79, 0.79, 0.76, 0.75, 0.75, 
    0.74, 0.79, 0.79, 0.8, 0.97, 0.94, 0.95, 0.84, 0.78, 0.81, 0.8, 0.83, 
    0.88, 0.88, 0.85, 0.82, 0.87, 0.83, 0.9, 0.8, 0.79, 0.83, 0.8, 0.77, 
    0.79, 0.81, 0.81, 0.74, 0.74, 0.76, 0.7, 0.71, 0.73, 0.73, 0.75, 0.75, 
    0.79, 0.77, 0.64, 0.66, 0.64, 0.63, 0.65, 0.6, 0.6, 0.6, 0.64, 0.66, 
    0.65, 0.67, 0.64, 0.63, 0.61, 0.6, 0.57, 0.54, 0.57, 0.6, 0.6, 0.6, 0.62, 
    0.62, 0.65, 0.6, 0.63, 0.64, 0.61, 0.58, 0.59, 0.59, 0.57, 0.59, 0.54, 
    0.51, 0.5, 0.51, 0.52, 0.55, 0.57, 0.57, 0.54, 0.58, 0.54, 0.54, 0.55, 
    0.56, 0.55, 0.52, 0.53, 0.54, 0.55, 0.56, 0.51, 0.53, 0.47, 0.49, 0.47, 
    0.46, 0.51, 0.52, 0.53, 0.5, 0.5, 0.48, 0.48, 0.46, 0.53, 0.52, 0.52, 
    0.51, 0.53, 0.55, 0.56, 0.57, 0.47, 0.58, 0.6, 0.55, 0.49, 0.53, 0.6, 
    0.58, 0.56, 0.59, 0.55, 0.54, 0.52, 0.49, 0.51, 0.52, 0.47, 0.47, 0.48, 
    0.5, 0.53, 0.51, 0.46, 0.45, 0.48, 0.45, 0.49, 0.46, 0.44, 0.46, 0.45, 
    0.47, 0.49, 0.48, 0.48, 0.49, 0.49, 0.47, 0.46, 0.4, 0.41, 0.43, 0.43, 
    0.43, 0.45, 0.43, 0.45, 0.48, 0.46, 0.57, 0.51, 0.44, 0.51, 0.51, 0.51, 
    0.53, 0.56, 0.62, 0.56, 0.58, 0.6, 0.58, 0.57, 0.56, 0.53, 0.53, 0.51, 
    0.51, 0.48, 0.48, 0.49, 0.52, 0.5, 0.55, 0.51, 0.49, 0.49, 0.44, 0.39, 
    0.44, 0.47, 0.44, 0.52, 0.48, 0.48, 0.49, 0.5, 0.51, 0.53, 0.48, 0.5, 
    0.46, 0.5, 0.46, 0.48, 0.5, 0.51, 0.6, 0.54, 0.58, 0.62, 0.63, 0.54, 
    0.54, 0.54, 0.51, 0.52, 0.53, 0.53, 0.52, 0.53, 0.56, 0.53, 0.49, 0.6, 
    0.54, 0.49, 0.52, 0.58, 0.54, 0.57, 0.54, 0.56, 0.6, 0.58, 0.58, 0.59, 
    0.57, 0.59, 0.63, 0.67, 0.53, 0.56, 0.55, 0.56, 0.54, 0.56, 0.55, 0.56, 
    0.52, 0.53, 0.56, 0.51, 0.5, 0.51, 0.51, 0.5, 0.5, 0.48, 0.5, 0.53, 0.58, 
    0.56, 0.54, 0.57, 0.6, 0.6, 0.59, 0.59, 0.66, 0.64, 0.64, 0.64, 0.65, 
    0.67, 0.67, 0.65, 0.65, 0.65, 0.68, 0.67, 0.65, 0.63, 0.7, 0.64, 0.65, 
    0.66, 0.64, 0.63, 0.68, 0.66, 0.65, 0.65, 0.64, 0.67, 0.64, 0.69, 0.67, 
    0.7, 0.69, 0.7, 0.68, 0.68, 0.66, 0.7, 0.7, 0.66, 0.7, 0.7, 0.69, 0.68, 
    0.69, 0.7, 0.7, 0.7, 0.71, 0.72, 0.72, 0.72, 0.73, 0.71, 0.72, 0.73, 
    0.74, 0.74, 0.73, 0.77, 0.65, 0.7, 0.63, 0.53, 0.51, 0.48, 0.47, 0.48, 
    0.45, 0.44, 0.45, 0.44, 0.46, 0.47, 0.45, 0.45, 0.42, 0.43, 0.47, 0.41, 
    0.42, 0.39, 0.43, 0.49, 0.54, 0.58, 0.58, 0.67, 0.61, 0.66, 0.69, 0.73, 
    0.78, 0.77, 0.67, 0.58, 0.57, 0.46, 0.44, 0.44, 0.43, 0.45, 0.56, 0.58, 
    0.57, 0.53, 0.52, 0.5, 0.51, 0.61, 0.56, 0.6, 0.66, 0.67, 0.66, 0.67, 
    0.67, 0.66, 0.66, 0.68, 0.69, 0.68, 0.67, 0.68, 0.7, 0.7, 0.7, 0.67, 
    0.68, 0.68, 0.65, 0.61, 0.59, 0.57, 0.68, 0.84, 0.83, 0.83, 0.93, 0.92, 
    0.76, 0.69, 0.72, 0.79, 0.78, 0.7, 0.8, 0.73, 0.85, 0.72, 0.67, 0.59, 
    0.59, 0.6, 0.67, 0.67, 0.61, 1, 1, 0.98, 0.98, 0.98, 0.95, 0.96, 0.95, 
    0.92, 0.84, 0.86, 0.77, 0.79, 0.74, 0.79, 0.78, 0.76, 0.75, 0.7, 0.71, 
    0.66, 0.68, 0.64, 0.71, 0.72, 0.69, 0.67, 0.69, 0.69, 0.67, 0.57, 0.61, 
    0.63, 0.57, 0.62, 0.6, 0.65, 0.61, 0.59, 0.59, 0.62, 0.65, 0.66, 0.69, 
    0.74, 0.88, 0.89, 0.86, 0.82, 0.77, 0.67, 0.64, 0.59, 0.61, 0.6, 0.59, 
    0.61, 0.58, 0.6, 0.57, 0.65, 0.67, 0.66, 0.63, 0.61, 0.56, 0.6, 0.63, 
    0.55, 0.52, 0.53, 0.52, 0.5, 0.5, 0.5, 0.49, 0.46, 0.45, 0.46, 0.45, 
    0.48, 0.47, 0.49, 0.5, 0.53, 0.53, 0.53, 0.54, 0.51, 0.53, 0.58, 0.6, 
    0.63, 0.67, 0.67, 0.61, 0.58, 0.64, 0.62, 0.64, 0.65, 0.66, 0.66, 0.61, 
    0.57, 0.6, 0.54, 0.61, 0.63, 0.7, 0.52, 0.47, 0.5, 0.57, 0.57, 0.53, 
    0.55, 0.52, 0.54, 0.52, 0.51, 0.52, 0.49, 0.49, 0.48, 0.48, 0.49, 0.49, 
    0.51, 0.51, 0.53, 0.54, 0.51, 0.54, 0.49, 0.48, 0.44, 0.46, 0.6, 0.56, 
    0.56, 0.56, 0.53, 0.54, 0.53, 0.55, 0.51, 0.45, 0.49, 0.5, 0.51, 0.48, 
    0.55, 0.56, 0.44, 0.43, 0.45, 0.5, 0.5, 0.54, 0.57, 0.56, 0.52, 0.5, 
    0.49, 0.55, 0.56, 0.53, 0.49, 0.48, 0.49, 0.49, 0.49, 0.5, 0.5, 0.5, 0.5, 
    0.5, 0.56, 0.61, 0.59, 0.64, 0.6, 0.55, 0.59, 0.59, 0.5, 0.51, 0.55, 
    0.56, 0.6, 0.59, 0.61, 0.7, 0.69, 0.59, 0.57, 0.57, 0.57, 0.56, 0.57, 
    0.52, 0.5, 0.5, 0.58, 0.56, 0.56, 0.65, 0.79, 0.8, 0.79, 0.74, 0.76, 
    0.78, 0.77, 0.77, 0.97, 1, 0.96, 0.88, 0.86, 0.82, 0.75, 0.76, 0.62, 
    0.61, 0.59, 0.58, 0.55, 0.54, 0.57, 0.54, 0.58, 0.58, 0.55, 0.6, 0.6, 
    0.62, 0.63, 0.6, 0.52, 0.49, 0.44, 0.54, 0.58, 0.49, 0.47, 0.5, 0.5, 
    0.54, 0.66, 0.56, 0.59, 0.6, 0.64, 0.64, 0.6, 0.61, 0.65, 0.7, 0.68, 0.7, 
    0.65, 0.58, 0.59, 0.59, 0.55, 0.56, 0.56, 0.57, 0.6, 0.58, 0.56, 0.62, 
    0.62, 0.54, 0.58, 0.52, 0.53, 0.51, 0.5, 0.51, 0.51, 0.5, 0.59, 0.67, 
    0.64, 0.65, 0.67, 0.62, 0.62, 0.6, 0.62, 0.67, 0.68, 0.62, 0.55, 0.58, 
    0.62, 0.64, 0.63, 0.65, 0.54, 0.55, 0.56, 0.5, 0.52, 0.51, 0.56, 0.52, 
    0.56, 0.52, 0.47, 0.43, 0.47, 0.45, 0.47, 0.48, 0.46, 0.49, 0.5, 0.5, 
    0.55, 0.53, 0.5, 0.51, 0.54, 0.52, 0.5, 0.51, 0.51, 0.55, 0.55, 0.51, 
    0.58, 0.58, 0.58, 0.58, 0.63, 0.62, 0.64, 0.67, 0.66, 0.64, 0.61, 0.59, 
    0.6, 0.62, 0.67, 0.73, 0.75, 0.75, 0.77, 0.77, 0.75, 0.72, 0.68, 0.67, 
    0.7, 0.7, 0.71, 0.73, 0.74, 0.73, 0.77, 0.75, 0.73, 0.69, 0.71, 0.69, 
    0.72, 0.66, 0.63, 0.63, 0.64, 0.61, 0.64, 0.65, 0.68, 0.69, 0.72, 0.78, 
    0.82, 0.77, 0.75, 0.65, 0.65, 0.76, 0.77, 0.69, 0.76, 0.83, 0.75, 0.72, 
    0.76, 0.79, 0.81, 0.85, 0.87, 0.94, 0.89, 0.85, 0.81, 0.76, 0.71, 0.67, 
    0.67, 0.68, 0.7, 0.7, 0.64, 0.67, 0.71, 0.75, 0.77, 0.75, 0.78, 0.71, 
    0.78, 0.78, 0.76, 0.73, 0.74, 0.77, 0.78, 0.77, 0.76, 0.76, 0.81, 0.76, 
    0.76, 0.76, 0.71, 0.69, 0.72, 0.69, 0.67, 0.61, 0.65, 0.66, 0.65, 0.66, 
    0.91, 1, 1, 1, 1, 1, 0.99, 1, 1, 0.91, 0.93, 0.93, 0.94, 0.86, 0.84, 
    0.76, 0.75, 0.77, 0.76, 0.72, 0.82, 0.74, 0.84, 0.99, 1, 1, 1, 1, 1, 
    0.92, 0.92, 0.78, 0.84, 0.81, 0.84, 0.88, 0.94, 0.9, 0.86, 0.88, 0.91, 
    0.91, 0.87, 0.89, 0.84, 0.92, 0.97, 0.98, 0.67, 0.72, 0.95, 0.99, 0.91, 
    0.77, 0.64, 0.74, 0.77, 0.7, 0.72, 0.7, 0.73, 0.64, 0.58, 0.62, 0.61, 
    0.59, 0.57, 0.57, 0.56, 0.58, 0.6, 0.6, 0.63, 0.71, 0.69, 0.66, 0.66, 
    0.66, 0.57, 0.57, 0.64, 0.65, 0.64, 0.64, 0.64, 0.62, 0.63, 0.62, 0.61, 
    0.58, 0.58, 0.56, 0.54, 0.53, 0.55, 0.6, 0.57, 0.58, 0.55, 0.59, 0.55, 
    0.55, 0.57, 0.57, 0.55, 0.62, 0.55, 0.51, 0.54, 0.49, 0.56, 0.56, 0.58, 
    0.56, 0.61, 0.62, 0.59, 0.51, 0.51, 0.53, 0.59, 0.54, 0.57, 0.61, 0.54, 
    0.52, 0.54, 0.53, 0.54, 0.51, 0.52, 0.49, 0.47, 0.5, 0.49, 0.5, 0.51, 
    0.53, 0.6, 0.58, 0.55, 0.54, 0.57, 0.55, 0.55, 0.61, 0.64, 0.69, 0.58, 
    0.65, 0.53, 0.57, 0.52, 0.53, 0.49, 0.48, 0.49, 0.47, 0.44, 0.44, 0.46, 
    0.42, 0.44, 0.45, 0.49, 0.55, 0.55, 0.54, 0.52, 0.56, 0.55, 0.57, 0.62, 
    0.6, 0.61, 0.53, 0.53, 0.48, 0.48, 0.49, 0.46, 0.48, 0.44, 0.41, 0.41, 
    0.42, 0.4, 0.4, 0.42, 0.45, 0.51, 0.47, 0.58, 0.51, 0.62, 0.56, 0.58, 
    0.64, 0.63, 0.71, 0.68, 0.82, 0.78, 0.68, 0.69, 0.8, 0.63, 0.61, 0.6, 
    0.58, 0.59, 0.58, 0.58, 0.56, 0.58, 0.57, 0.48, 0.48, 0.46, 0.45, 0.43, 
    0.38, 0.36, 0.35, 0.3, 0.32, 0.42, 0.42, 0.39, 0.42, 0.46, 0.49, 0.51, 
    0.5, 0.48, 0.46, 0.44, 0.44, 0.45, 0.46, 0.49, 0.47, 0.44, 0.46, 0.45, 
    0.45, 0.47, 0.51, 0.46, 0.44, 0.45, 0.47, 0.51, 0.55, 0.57, 0.57, 0.61, 
    0.59, 0.6, 0.58, 0.6, 0.6, 0.6, 0.54, 0.58, 0.52, 0.48, 0.53, 0.46, 0.52, 
    0.49, 0.54, 0.52, 0.55, 0.52, 0.54, 0.55, 0.51, 0.52, 0.54, 0.54, 0.52, 
    0.54, 0.54, 0.58, 0.51, 0.6, 0.57, 0.61, 0.62, 0.58, 0.6, 0.61, 0.63, 
    0.59, 0.65, 0.63, 0.62, 0.67, 0.67, 0.66, 0.67, 0.68, 0.72, 0.64, 0.72, 
    0.76, 0.74, 0.68, 0.68, 0.72, 0.67, 0.74, 0.75, 0.7, 0.69, 0.67, 0.69, 
    0.71, 0.71, 0.75, 0.74, 0.76, 0.77, 0.78, 0.8, 0.8, 0.85, 0.8, 0.74, 
    0.75, 0.71, 0.63, 0.61, 0.59, 0.51, 0.51, 0.53, 0.6, 0.56, 0.61, 0.59, 
    0.58, 0.61, 0.63, 0.65, 0.62, 0.61, 0.59, 0.59, 0.6, 0.61, 0.64, 0.63, 
    0.64, 0.61, 0.66, 0.64, 0.67, 0.63, 0.62, 0.66, 0.64, 0.67, 0.64, 0.62, 
    0.6, 0.62, 0.58, 0.57, 0.57, 0.56, 0.57, 0.56, 0.58, 0.63, 0.55, 0.57, 
    0.6, 0.55, 0.54, 0.55, 0.53, 0.5, 0.56, 0.51, 0.51, 0.56, 0.51, 0.52, 
    0.55, 0.56, 0.47, 0.6, 0.61, 0.62, 0.58, 0.51, 0.54, 0.48, 0.54, 0.54, 
    0.58, 0.55, 0.59, 0.63, 0.5, 0.47, 0.41, 0.36, 0.35, 0.42, 0.44, 0.41, 
    0.42, 0.36, 0.33, 0.42, 0.5, 0.5, 0.5, 0.55, 0.54, 0.5, 0.5, 0.53, 0.56, 
    0.59, 0.52, 0.48, 0.57, 0.55, 0.54, 0.6, 0.61, 0.65, 0.67, 0.66, 0.67, 
    0.65, 0.7, 0.67, 0.64, 0.64, 0.58, 0.53, 0.48, 0.41, 0.43, 0.47, 0.46, 
    0.44, 0.45, 0.51, 0.5, 0.54, 0.54, 0.54, 0.52, 0.51, 0.5, 0.59, 0.54, 
    0.55, 0.57, 0.56, 0.57, 0.59, 0.6, 0.63, 0.64, 0.69, 0.71, 0.7, 0.73, 
    0.67, 0.71, 0.74, 0.75, 0.75, 0.72, 0.76, 0.78, 0.77, 0.86, 0.9, 0.92, 
    0.92, 0.91, 0.94, 0.95, 0.95, 0.98, 0.87, 0.86, 0.92, 0.85, 0.83, 0.78, 
    0.78, 0.76, 0.68, 0.7, 0.65, 0.65, 0.64, 0.63, 0.69, 0.7, 0.74, 0.73, 
    0.71, 0.69, 0.73, 0.7, 0.72, 0.75, 0.73, 0.72, 0.73, 0.73, 0.73, 0.78, 
    0.76, 0.87, 0.93, 0.93, 0.96, 0.95, 0.98, 0.99, 0.99, 0.98, 1, 1, 0.99, 
    1, 0.93, 0.94, 0.98, 0.96, 0.91, 0.98, 0.87, 0.73, 0.73, 0.72, 0.74, 
    0.71, 0.78, 0.79, 0.78, 0.79, 0.82, 0.92, 0.91, 0.87, 0.87, 0.86, 0.85, 
    0.97, 0.98, 1, 1, 0.99, 1, 0.95, 0.98, 0.97, 0.93, 0.96, 1, 1, 1, 1, 
    0.81, 0.76, 0.78, 0.82, 0.83, 0.82, 0.83, 0.91, 0.99, 1, 1, 1, 1, 1, 
    0.95, 1, 1, 1, 0.87, 0.78, 0.78, 0.78, 0.84, 0.79, 0.77, 0.75, 0.79, 
    0.77, 0.75, 0.76, 0.76, 0.8, 0.81, 0.8, 0.81, 0.76, 0.74, 0.68, 0.7, 
    0.72, 0.73, 0.75, 0.7, 0.75, 0.73, 0.73, 0.73, 0.75, 0.78, 0.83, 0.87, 
    0.89, 0.9, 0.9, 0.94, 0.97, 0.98, 0.96, 0.96, 0.93, 0.88, 0.93, 0.92, 
    0.95, 0.96, 0.98, 0.98, 0.93, 0.97, 0.98, 0.9, 0.94, 0.94, 0.95, 0.95, 
    0.94, 0.97, 0.97, 0.97, 0.91, 0.92, 0.93, 0.92, 0.9, 0.9, 0.88, 0.85, 
    0.84, 0.81, 0.85, 0.83, 0.81, 0.81, 0.83, 0.83, 0.83, 0.79, 0.78, 0.78, 
    0.83, 0.81, 0.81, 0.84, 0.82, 0.79, 0.84, 0.8, 0.84, 0.84, 0.83, 0.81, 
    0.82, 0.79, 0.8, 0.84, 0.82, 0.81, 0.83, 0.8, 0.78, 0.79, 0.78, 0.79, 
    0.78, 0.79, 0.79, 0.79, 0.8, 0.8, 0.82, 0.81, 0.79, 0.79, 0.78, 0.77, 
    0.78, 0.79, 0.8, 0.78, 0.77, 0.72, 0.74, 0.79, 0.8, 0.78, 0.81, 0.81, 
    0.77, 0.81, 0.87, 0.92, 0.88, 0.91, 0.9, 0.94, 0.91, 0.91, 0.86, 0.85, 
    0.85, 0.87, 0.84, 0.83, 0.83, 0.84, 0.87, 0.89, 0.88, 0.87, 0.87, 0.81, 
    0.83, 0.82, 0.86, 0.86, 0.86, 0.85, 0.83, 0.83, 0.79, 0.77, 0.77, 0.77, 
    0.78, 0.75, 0.75, 0.77, 0.74, 0.82, 0.83, 0.79, 0.73, 0.74, 0.74, 0.75, 
    0.75, 0.79, 0.87, 0.91, 0.95, 0.96, 0.97, 0.97, 0.96, 0.98, 1, 0.98, 
    0.95, 0.95, 1, 0.94, 0.95, 0.91, 0.86, 0.82, 0.84, 0.74, 0.77, 0.87, 
    0.92, 0.8, 0.8, 0.83, 0.81, 0.87, 0.92, 0.86, 0.91, 0.92, 0.97, 0.95, 
    0.9, 0.89, 0.87, 0.86, 0.87, 0.89, 0.87, 0.89, 0.94, 0.92, 0.87, 0.86, 
    0.87, 0.88, 0.94, 0.89, 0.9, 0.95, 0.97, 0.93, 0.93, 0.95, 0.91, 0.9, 
    0.91, 0.89, 0.92, 0.91, 0.9, 0.91, 0.9, 0.89, 0.9, 0.88, 0.83, 0.87, 
    0.89, 0.9, 0.89, 0.88, 0.87, 0.88, 0.89, 0.92, 0.9, 0.92, 0.88, 0.85, 
    0.83, 0.83, 0.85, 0.85, 0.82, 0.8, 0.87, 0.81, 0.83, 0.84, 0.85, 0.83, 
    0.85, 0.93, 0.95, 0.89, 0.85, 0.85, 0.9, 0.88, 0.87, 0.92, 0.83, 0.79, 
    0.87, 0.75, 0.73, 0.73, 0.75, 0.74, 0.76, 0.85, 0.77, 0.77, 0.74, 0.72, 
    0.71, 0.72, 0.71, 0.72, 0.72, 0.71, 0.69, 0.66, 0.64, 0.6, 0.59, 0.59, 
    0.59, 0.69, 0.7, 0.71, 0.71, 0.82, 0.89, 0.8, 0.85, 0.88, 0.8, 0.73, 
    0.71, 0.73, 0.71, 0.68, 0.68, 0.7, 0.72, 0.83, 0.83, 0.79, 0.74, 0.76, 
    0.78, 0.69, 0.68, 0.7, 0.7, 0.71, 0.71, 0.72, 0.72, 0.72, 0.71, 0.65, 
    0.69, 0.9, 0.92, 0.96, 0.93, 0.96, 0.93, 0.95, 0.94, 0.95, 0.94, 0.91, 
    0.91, 0.88, 0.86, 0.81, 0.79, 0.78, 0.78, 0.8, 0.82, 0.87, 0.73, 0.69, 
    0.68, 0.88, 0.82, 0.83, 0.95, 0.87, 0.88, 0.89, 0.89, 0.93, 0.94, 0.94, 
    0.95, 0.81, 0.88, 0.91, 0.91, 0.89, 0.87, 0.86, 0.86, 0.87, 0.9, 0.93, 
    0.95, 0.91, 0.94, 0.85, 0.84, 0.86, 0.84, 0.85, 0.86, 0.85, 0.84, 0.82, 
    0.84, 0.81, 0.81, 0.8, 0.78, 0.78, 0.78, 0.78, 0.77, 0.77, 0.76, 0.75, 
    0.72, 0.87, 0.81, 0.84, 0.9, 0.87, 0.86, 0.85, 0.84, 0.84, 0.85, 0.85, 
    0.9, 0.79, 0.79, 0.81, 0.82, 0.84, 0.83, 0.83, 0.83, 0.8, 0.84, 0.85, 
    0.88, 0.8, 0.77, 0.79, 0.83, 0.88, 0.89, 0.88, 0.8, 0.78, 0.73, 0.76, 
    0.78, 0.81, 0.84, 0.84, 0.85, 0.74, 0.72, 0.72, 0.81, 0.89, 0.87, 0.94, 
    0.88, 0.75, 0.77, 0.78, 0.79, 0.77, 0.79, 0.81, 0.82, 0.86, 0.92, 0.7, 
    0.74, 0.86, 1, 0.9, 0.94, 0.95, 0.95, 0.93, 0.94, 0.95, 0.96, 1, 1, 0.96, 
    0.97, 0.95, 0.99, 1, 1, 0.94, 0.93, 0.91, 0.92, 0.96, 0.95, 0.93, 0.95, 
    0.95, 0.94, 0.96, 0.96, 0.96, 0.91, 0.88, 0.99, 0.94, 0.95, 0.99, 0.92, 
    0.91, 0.91, 0.9, 0.91, 0.93, 0.93, 0.96, 0.89, 0.9, 0.91, 0.91, 0.92, 
    0.93, 0.94, 0.88, 0.9, 0.92, 0.91, 0.9, 0.87, 0.9, 0.84, 0.9, 0.92, 0.86, 
    0.92, 0.94, 0.94, 0.9, 0.91, 0.91, 0.91, 0.87, 0.86, 0.87, 0.86, 0.86, 
    0.85, 0.89, 0.88, 0.89, 0.89, 0.88, 0.86, 0.86, 0.89, 0.85, 0.85, 0.89, 
    0.9, 0.9, 0.9, 0.9, 0.89, 0.88, 0.86, 0.86, 0.88, 0.82, 0.82, 0.84, 0.84, 
    0.84, 0.8, 0.79, 0.81, 0.84, 0.88, 0.85, 0.9, 0.85, 0.84, 0.82, 0.81, 
    0.81, 0.79, 0.74, 0.63, 0.54, 0.54, 0.51, 0.52, 0.76, 0.58, 0.69, 0.76, 
    0.8, 0.81, 0.81, 0.81, 0.87, 0.86, 0.9, 0.94, 0.94, 0.99, 1, 1, 1, 0.96, 
    0.85, 0.83, 0.81, 0.79, 0.79, 0.85, 0.85, 0.83, 0.83, 0.83, 0.83, 0.83, 
    0.87, 0.86, 0.93, 0.99, 0.99, 1, 1, 1, 1, 1, 1, 1, 0.96, 0.82, 0.72, 
    0.69, 0.76, 0.81, 0.75, 0.84, 0.92, 0.96, 0.96, 1, 0.89, 0.91, 0.91, 
    0.89, 0.85, 0.9, 0.87, 0.88, 0.86, 0.84, 0.84, 0.84, 0.88, 0.9, 0.93, 
    0.96, 0.97, 0.96, 0.93, 0.97, 0.96, 0.91, 0.87, 0.85, 0.85, 0.82, 0.84, 
    0.81, 0.82, 0.8, 0.81, 0.83, 0.95, 0.92, 0.89, 0.83, 0.81, 0.87, 0.86, 
    0.9, 0.91, 0.89, 0.94, 0.91, 0.95, 0.95, 0.93, 0.92, 0.91, 0.92, 0.92, 
    0.91, 0.91, 0.91, 0.87, 0.9, 0.93, 0.91, 0.89, 0.85, 0.85, 0.87, 0.88, 
    0.94, 1, 0.97, 0.93, 0.94, 0.93, 0.91, 0.9, 0.93, 0.84, 0.78, 0.79, 0.85, 
    0.73, 0.66, 0.53, 0.61, 0.65, 0.68, 0.71, 0.73, 0.73, 0.71, 0.71, 0.71, 
    0.71, 0.72, 0.66, 0.63, 0.61, 0.61, 0.62, 0.65, 0.65, 0.64, 0.65, 0.66, 
    0.66, 0.64, 0.6, 0.61, 0.73, 0.85, 0.85, 0.76, 0.82, 0.86, 0.86, 0.95, 
    0.96, 0.92, 0.91, 0.86, 0.89, 0.95, 0.96, 0.88, 0.91, 0.97, 0.97, 0.97, 
    0.97, 0.97, 0.94, 0.93, 0.93, 0.94, 0.95, 1, 0.99, 1, 1, 1, 1, 0.98, 1, 
    1, 1, 0.69, 0.68, 0.74, 0.66, 0.7, 0.68, 0.98, 0.97, 0.96, 0.79, 0.8, 
    0.81, 0.87, 0.88, 0.82, 0.77, 0.85, 0.91, 0.84, 0.81, 0.82, 0.88, 0.86, 
    0.86, 0.88, 0.93, 0.96, 0.99, 0.99, 0.95, 0.89, 0.86, 0.86, 0.68, 0.67, 
    0.68, 0.68, 0.65, 0.66, 0.69, 0.73, 0.74, 0.72, 0.72, 0.73, 0.73, 0.79, 
    0.74, 0.73, 0.77, 0.84, 0.86, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0.92, 0.96, 0.96, 0.95, 0.96, 0.97, 0.98, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.98, 0.98, 0.96, 0.96, 0.94, 
    0.93, 0.92, 0.93, 0.98, 0.94, 0.97, 1, 1, 1, 0.98, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.91, 0.95, 1, 1, 
    1, 1, 1, 0.96, 0.98, 1, 0.99, 0.83, 0.72, 0.75, 0.83, 0.83, 0.81, 0.92, 
    0.78, 0.84, 0.96, 0.95, 0.94, 0.9, 0.96, 1, 1, 1, 1, 0.98, 0.88, 0.96, 
    0.94, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.96, 0.84, 0.79, 0.79, 0.79, 
    0.79, 0.81, 0.81, 0.81, 0.8, 0.8, 0.82, 0.82, 0.84, 0.84, 0.84, 0.85, 
    0.86, 0.85, 0.86, 0.92, 0.91, 0.9, 0.9, 0.88, 0.87, 0.88, 0.87, 0.88, 
    0.88, 0.87, 0.86, 0.9, 0.91, 0.89, 0.88, 0.78, 0.65, 0.69, 0.7, 0.69, 
    0.71, 0.73, 0.73, 0.73, 0.74, 0.91, 0.98, 0.91, 0.95, 1, 0.97, 0.96, 
    0.99, 0.99, 1, 0.9, 0.92, 0.94, 0.99, 1, 1, 0.99, 1, 0.97, 0.95, 1, 0.88, 
    0.93, 0.9, 0.91, 0.93, 0.97, 0.96, 0.93, 0.91, 0.91, 0.91, 0.91, 0.91, 
    0.94, 0.95, 0.95, 0.97, 0.97, 0.95, 0.94, 0.94, 0.91, 0.92, 0.91, 0.92, 
    0.94, 0.93, 0.93, 0.94, 0.95, 0.94, 0.94, 0.94, 0.95, 0.96, 0.95, 0.95, 
    0.95, 0.95, 0.96, 0.95, 0.95, 0.95, 0.93, 0.93, 0.94, 0.95, 0.93, 0.91, 
    0.83, 0.8, 0.81, 0.76, 0.75, 0.72, 0.71, 0.75, 0.81, 0.69, 0.73, 0.72, 
    0.72, 0.7, 0.67, 0.69, 0.63, 0.62, 0.59, 0.39, 0.39, 0.43, 0.43, 0.52, 
    0.54, 0.53, 0.53, 0.53, 0.53, 0.54, 0.55, 0.56, 0.58, 0.54, 0.61, 0.61, 
    0.56, 0.62, 0.63, 0.62, 0.58, 0.62, 0.63, 0.65, 0.65, 0.61, 0.65, 0.64, 
    0.64, 0.61, 0.62, 0.64, 0.59, 0.61, 0.63, 0.6, 0.66, 0.51, 0.54, 0.59, 
    0.61, 0.53, 0.61, 0.58, 0.64, 0.63, 0.79, 0.77, 0.6, 0.64, 0.58, 0.57, 
    0.63, 0.57, 0.54, 0.46, 0.52, 0.54, 0.61, 0.61, 0.6, 0.59, 0.62, 0.63, 
    0.66, 0.56, 0.57, 0.57, 0.53, 0.51, 0.55, 0.6, 0.59, 0.55, 0.56, 0.62, 
    0.62, 0.64, 0.65, 0.65, 0.68, 0.81, 0.76, 0.7, 0.7, 0.65, 0.56, 0.59, 
    0.58, 0.62, 0.61, 0.54, 0.54, 0.59, 0.59, 0.57, 0.59, 0.59, 0.58, 0.61, 
    0.63, 0.66, 0.59, 0.58, 0.57, 0.57, 0.56, 0.54, 0.57, 0.6, 0.62, 0.59, 
    0.58, 0.57, 0.59, 0.54, 0.54, 0.53, 0.61, 0.61, 0.6, 0.65, 0.65, 0.65, 
    0.61, 0.6, 0.62, 0.62, 0.6, 0.63, 0.61, 0.58, 0.61, 0.63, 0.6, 0.59, 
    0.59, 0.57, 0.6, 0.63, 0.59, 0.61, 0.64, 0.65, 0.63, 0.64, 0.6, 0.71, 
    0.71, 0.68, 0.59, 0.68, 0.58, 0.59, 0.72, 0.65, 0.63, 0.7, 0.65, 0.63, 
    0.67, 0.62, 0.64, 0.61, 0.58, 0.57, 0.66, 0.7, 0.63, 0.74, 0.7, 0.66, 
    0.66, 0.69, 0.65, 0.65, 0.72, 0.68, 0.63, 0.72, 0.66, 0.7, 0.7, 0.67, 
    0.73, 0.69, 0.69, 0.69, 0.58, 0.64, 0.71, 0.72, 0.63, 0.73, 0.69, 0.7, 
    0.69, 0.69, 0.73, 0.72, 0.7, 0.65, 0.65, 0.73, 0.73, 0.68, 0.73, 0.71, 
    0.71, 0.73, 0.72, 0.63, 0.66, 0.58, 0.71, 0.71, 0.69, 0.68, 0.71, 0.68, 
    0.69, 0.73, 0.67, 0.68, 0.69, 0.64, 0.67, 0.7, 0.66, 0.63, 0.63, 0.64, 
    0.67, 0.62, 0.51, 0.52, 0.54, 0.59, 0.61, 0.61, 0.56, 0.52, 0.54, 0.54, 
    0.48, 0.46, 0.49, 0.53, 0.55, 0.53, 0.5, 0.44, 0.44, 0.59, 0.46, 0.54, 
    0.51, 0.5, 0.46, 0.49, 0.42, 0.51, 0.53, 0.48, 0.64, 0.49, 0.56, 0.6, 
    0.58, 0.63, 0.61, 0.61, 0.66, 0.56, 0.65, 0.64, 0.56, 0.66, 0.65, 0.66, 
    0.67, 0.58, 0.59, 0.57, 0.51, 0.5, 0.58, 0.64, 0.63, 0.6, 0.55, 0.63, 
    0.54, 0.56, 0.56, 0.52, 0.51, 0.53, 0.57, 0.6, 0.54, 0.53, 0.6, 0.48, 
    0.58, 0.54, 0.51, 0.55, 0.49, 0.56, 0.58, 0.59, 0.52, 0.69, 0.7, 0.6, 
    0.54, 0.59, 0.6, 0.59, 0.94, 0.57, 0.57, 0.6, 0.62, 0.56, 0.54, 0.63, 
    0.71, 0.56, 0.59, 0.62, 0.7, 0.68, 0.62, 0.68, 0.77, 0.8, 0.83, 0.81, 
    0.83, 0.85, 0.85, 0.85, 0.85, 0.8, 0.83, 0.86, 0.87, 0.86, 0.83, 0.84, 
    0.84, 0.83, 0.83, 0.83, 0.82, 0.8, 0.78, 0.78, 0.82, 0.75, 0.83, 0.72, 
    0.83, 0.82, 0.81, 0.86, 0.86, 0.87, 0.88, 0.88, 0.89, 0.88, 0.88, 0.9, 
    0.88, 0.86, 0.86, 0.84, 0.8, 0.83, 0.86, 0.86, 0.86, 0.87, 0.88, 0.93, 
    0.95, 0.91, 0.93, 0.93, 0.95, 0.96, 0.97, 0.96, 0.95, 0.98, 0.7, 0.72, 
    0.74, 0.8, 0.74, 0.7, 0.68, 0.68, 0.69, 0.71, 0.72, 0.7, 0.7, 0.68, 0.76, 
    0.72, 0.72, 0.67, 0.64, 0.69, 0.68, 0.66, 0.81, 0.87, 0.82, 0.86, 0.81, 
    0.73, 0.67, 0.64, 0.65, 0.6, 0.6, 0.56, 0.64, 0.52, 0.52, 0.52, 0.52, 
    0.54, 0.55, 0.55, 0.53, 0.5, 0.51, 0.56, 0.58, 0.59, 0.58, 0.61, 0.59, 
    0.58, 0.52, 0.51, 0.53, 0.52, 0.51, 0.53, 0.6, 0.57, 0.54, 0.56, 0.61, 
    0.63, 0.63, 0.6, 0.65, 0.52, 0.66, 0.6, 0.6, 0.59, 0.65, 0.61, 0.53, 
    0.58, 0.56, 0.59, 0.61, 0.55, 0.55, 0.54, 0.54, 0.55, 0.54, 0.53, 0.56, 
    0.57, 0.61, 0.57, 0.59, 0.59, 0.6, 0.59, 0.56, 0.55, 0.56, 0.58, 0.56, 
    0.54, 0.57, 0.59, 0.57, 0.52, 0.5, 0.51, 0.55, 0.61, 0.54, 0.6, 0.6, 
    0.58, 0.56, 0.64, 0.64, 0.62, 0.82, 0.66, 0.58, 0.64, 0.64, 0.6, 0.68, 
    0.65, 0.66, 0.67, 0.65, 0.54, 0.49, 0.48, 0.46, 0.5, 0.44, 0.43, 0.45, 
    0.49, 0.49, 0.47, 0.5, 0.54, 0.53, 0.5, 0.47, 0.54, 0.56, 0.49, 0.46, 
    0.52, 0.55, 0.52, 0.45, 0.44, 0.44, 0.41, 0.4, 0.42, 0.44, 0.42, 0.42, 
    0.42, 0.45, 0.39, 0.56, 0.49, 0.49, 0.61, 0.56, 0.5, 0.52, 0.42, 0.45, 
    0.43, 0.49, 0.53, 0.49, 0.51, 0.52, 0.46, 0.48, 0.48, 0.44, 0.43, 0.42, 
    0.43, 0.39, 0.38, 0.42, 0.39, 0.47, 0.52, 0.59, 0.58, 0.61, 0.62, 0.62, 
    0.62, 0.58, 0.58, 0.53, 0.47, 0.39, 0.46, 0.5, 0.54, 0.57, 0.6, 0.55, 
    0.6, 0.63, 0.65, 0.63, 0.61, 0.63, 0.53, 0.65, 0.65, 0.58, 0.59, 0.57, 
    0.61, 0.55, 0.5, 0.44, 0.46, 0.57, 0.53, 0.55, 0.56, 0.55, 0.55, 0.6, 
    0.61, 0.58, 0.57, 0.55, 0.58, 0.57, 0.57, 0.56, 0.6, 0.59, 0.59, 0.57, 
    0.58, 0.58, 0.57, 0.61, 0.62, 0.54, 0.62, 0.65, 0.67, 0.68, 0.67, 0.66, 
    0.72, 0.74, 0.73, 0.69, 0.69, 0.69, 0.7, 0.69, 0.67, 0.74, 0.69, 0.76, 
    0.75, 0.73, 0.71, 0.56, 0.57, 0.56, 0.55, 0.47, 0.56, 0.51, 0.49, 0.57, 
    0.61, 0.63, 0.63, 0.61, 0.58, 0.63, 0.62, 0.61, 0.63, 0.64, 0.72, 0.58, 
    0.63, 0.61, 0.62, 0.55, 0.54, 0.52, 0.56, 0.54, 0.57, 0.59, 0.6, 0.72, 
    0.64, 0.65, 0.65, 0.65, 0.64, 0.65, 0.67, 0.64, 0.64, 0.62, 0.59, 0.61, 
    0.6, 0.56, 0.55, 0.53, 0.57, 0.58, 0.53, 0.56, 0.55, 0.56, 0.58, 0.64, 
    0.63, 0.66, 0.65, 0.7, 0.7, 0.66, 0.7, 0.65, 0.7, 0.64, 0.59, 0.55, 0.53, 
    0.48, 0.48, 0.49, 0.51, 0.52, 0.52, 0.51, 0.5, 0.52, 0.51, 0.54, 0.6, 
    0.61, 0.58, 0.62, 0.56, 0.58, 0.59, 0.59, 0.59, 0.58, 0.52, 0.54, 0.53, 
    0.48, 0.51, 0.52, 0.53, 0.54, 0.54, 0.51, 0.5, 0.58, 0.59, 0.66, 0.65, 
    0.65, 0.64, 0.67, 0.6, 0.6, 0.68, 0.65, 0.62, 0.63, 0.57, 0.54, 0.63, 
    0.57, 0.55, 0.54, 0.59, 0.56, 0.61, 0.56, 0.65, 0.6, 0.68, 0.67, 0.72, 
    0.61, 0.67, 0.61, 0.69, 0.65, 0.66, 0.65, 0.66, 0.64, 0.64, 0.63, 0.63, 
    0.59, 0.6, 0.62, 0.62, 0.59, 0.56, 0.65, 0.6, 0.61, 0.62, 0.58, 0.59, 
    0.62, 0.6, 0.54, 0.54, 0.56, 0.59, 0.6, 0.58, 0.56, 0.54, 0.55, 0.51, 
    0.56, 0.47, 0.51, 0.49, 0.56, 0.61, 0.57, 0.59, 0.63, 0.65, 0.65, 0.62, 
    0.63, 0.58, 0.64, 0.63, 0.66, 0.6, 0.65, 0.67, 0.6, 0.66, 0.57, 0.52, 
    0.56, 0.54, 0.53, 0.48, 0.53, 0.58, 0.53, 0.55, 0.51, 0.63, 0.61, 0.64, 
    0.61, 0.65, 0.67, 0.64, 0.68, 0.66, 0.68, 0.7, 0.67, 0.68, 0.61, 0.62, 
    0.61, 0.57, 0.53, 0.63, 0.58, 0.6, 0.59, 0.52, 0.54, 0.56, 0.58, 0.6, 
    0.6, 0.64, 0.61, 0.63, 0.63, 0.62, 0.62, 0.63, 0.62, 0.65, 0.63, 0.55, 
    0.57, 0.52, 0.59, 0.57, 0.61, 0.59, 0.63, 0.61, 0.65, 0.62, 0.63, 0.65, 
    0.71, 0.69, 0.6, 0.65, 0.63, 0.63, 0.67, 0.65, 0.64, 0.63, 0.63, 0.61, 
    0.72, 0.71, 0.62, 0.62, 0.6, 0.61, 0.6, 0.59, 0.73, 0.74, 0.73, 0.8, 
    0.78, 0.79, 0.79, 0.76, 0.76, 0.75, 0.77, 0.83, 0.83, 0.81, 0.82, 0.72, 
    0.73, 0.69, 0.69, 0.54, 0.58, 0.63, 0.62, 0.76, 0.84, 0.84, 0.6, 0.63, 
    0.54, 0.57, 0.58, 0.61, 0.6, 0.58, 0.61, 0.63, 0.68, 0.65, 0.6, 0.56, 
    0.6, 0.57, 0.6, 0.54, 0.52, 0.6, 0.49, 0.58, 0.59, 0.6, 0.58, 0.68, 0.62, 
    0.65, 0.57, 0.63, 0.64, 0.64, 0.7, 0.71, 0.71, 0.7, 0.74, 0.76, 0.76, 
    0.8, 0.83, 0.81, 0.8, 0.85, 0.86, 0.84, 0.87, 0.88, 0.88, 0.9, 0.83, 
    0.84, 0.78, 0.77, 0.79, 0.8, 0.85, 0.85, 0.87, 0.88, 0.86, 0.83, 0.84, 
    0.83, 0.81, 0.81, 0.82, 0.84, 0.87, 0.9, 0.93, 0.95, 0.95, 0.92, 0.86, 
    0.83, 0.81, 0.78, 0.76, 0.74, 0.7, 0.67, 0.71, 0.68, 0.66, 0.64, 0.62, 
    0.59, 0.58, 0.58, 0.54, 0.6, 0.59, 0.55, 0.54, 0.56, 0.59, 0.65, 0.61, 
    0.64, 0.63, 0.69, 0.67, 0.74, 0.73, 0.78, 0.7, 0.69, 0.65, 0.64, 0.6, 
    0.61, 0.59, 0.72, 0.63, 0.62, 0.68, 0.74, 0.77, 0.76, 0.78, 0.8, 0.84, 
    0.66, 0.66, 0.63, 0.71, 0.72, 0.7, 0.74, 0.74, 0.68, 0.64, 0.63, 0.62, 
    0.61, 0.52, 0.68, 0.7, 0.64, 0.67, 0.73, 0.74, 0.72, 0.77, 0.87, 0.91, 
    0.92, 0.92, 0.92, 0.9, 0.91, 0.9, 0.91, 0.89, 0.85, 0.86, 0.76, 0.77, 
    0.81, 0.78, 0.77, 0.77, 0.74, 0.83, 0.82, 0.88, 0.86, 0.91, 0.93, 0.96, 
    0.97, 0.99, 0.99, 0.99, 0.97, 0.98, 0.88, 0.76, 0.69, 0.67, 0.65, 0.6, 
    0.58, 0.54, 0.5, 0.51, 0.44, 0.48, 0.53, 0.49, 0.53, 0.54, 0.53, 0.54, 
    0.57, 0.6, 0.59, 0.56, 0.54, 0.56, 0.6, 0.6, 0.59, 0.52, 0.52, 0.51, 
    0.52, 0.53, 0.56, 0.55, 0.53, 0.6, 0.58, 0.56, 0.6, 0.61, 0.67, 0.67, 
    0.69, 0.67, 0.71, 0.71, 0.68, 0.65, 0.67, 0.62, 0.64, 0.57, 0.53, 0.51, 
    0.52, 0.56, 0.58, 0.49, 0.58, 0.54, 0.59, 0.56, 0.58, 0.65, 0.68, 0.71, 
    0.68, 0.67, 0.75, 0.75, 0.74, 0.74, 0.65, 0.63, 0.68, 0.59, 0.61, 0.51, 
    0.58, 0.6, 0.48, 0.62, 0.61, 0.62, 0.61, 0.62, 0.65, 0.8, 0.9, 0.93, 
    0.85, 0.87, 0.88, 0.9, 0.9, 0.89, 0.9, 0.87, 0.84, 0.81, 0.83, 0.83, 0.8, 
    0.8, 0.83, 0.84, 0.74, 0.73, 0.67, 0.62, 0.61, 0.61, 0.63, 0.69, 0.7, 
    0.69, 0.63, 0.6, 0.7, 0.65, 0.62, 0.72, 0.7, 0.69, 0.68, 0.66, 0.61, 
    0.58, 0.48, 0.51, 0.55, 0.5, 0.59, 0.58, 0.57, 0.59, 0.58, 0.65, 0.67, 
    0.7, 0.67, 0.66, 0.72, 0.69, 0.67, 0.67, 0.58, 0.65, 0.53, 0.52, 0.48, 
    0.51, 0.56, 0.55, 0.56, 0.62, 0.56, 0.6, 0.58, 0.58, 0.53, 0.48, 0.49, 
    0.48, 0.48, 0.5, 0.56, 0.62, 0.56, 0.55, 0.57, 0.54, 0.51, 0.52, 0.5, 
    0.52, 0.54, 0.53, 0.56, 0.56, 0.55, 0.48, 0.46, 0.57, 0.62, 0.63, 0.58, 
    0.61, 0.65, 0.68, 0.66, 0.7, 0.62, 0.6, 0.61, 0.56, 0.5, 0.54, 0.49, 
    0.51, 0.6, 0.56, 0.5, 0.5, 0.54, 0.55, 0.58, 0.59, 0.63, 0.7, 0.7, 0.7, 
    0.71, 0.73, 0.66, 0.75, 0.68, 0.65, 0.71, 0.61, 0.54, 0.52, 0.51, 0.52, 
    0.53, 0.54, 0.5, 0.62, 0.62, 0.62, 0.6, 0.62, 0.91, 0.75, 0.79, 0.77, 
    0.8, 0.79, 0.82, 0.81, 0.76, 0.7, 0.74, 0.64, 0.66, 0.58, 0.49, 0.62, 
    0.55, 0.55, 0.62, 0.52, 0.61, 0.64, 0.72, 0.7, 0.68, 0.73, 0.72, 0.7, 
    0.74, 0.72, 0.72, 0.68, 0.71, 0.69, 0.68, 0.62, 0.69, 0.66, 0.61, 0.69, 
    0.75, 0.75, 0.82, 0.8, 0.78, 0.79, 0.82, 0.86, 0.87, 0.89, 0.83, 0.83, 
    0.78, 0.84, 0.79, 0.81, 0.86, 0.85, 0.79, 0.75, 0.72, 0.73, 0.61, 0.6, 
    0.48, 0.6, 0.51, 0.65, 0.63, 0.64, 0.65, 0.74, 0.73, 0.72, 0.71, 0.68, 
    0.71, 0.75, 0.7, 0.68, 0.65, 0.71, 0.69, 0.63, 0.66, 0.62, 0.68, 0.69, 
    0.71, 0.69, 0.76, 0.74, 0.8, 0.79, 0.83, 0.76, 0.85, 0.93, 0.97, 0.95, 
    0.91, 0.91, 0.93, 0.93, 0.86, 0.84, 0.8, 0.79, 0.75, 0.76, 0.73, 0.74, 
    0.68, 0.69, 0.7, 0.63, 0.7, 0.71, 0.78, 0.79, 0.8, 0.84, 0.84, 0.81, 
    0.91, 0.83, 0.87, 0.81, 0.79, 0.85, 0.83, 0.83, 0.72, 0.79, 0.73, 0.78, 
    0.79, 0.76, 0.72, 0.8, 0.8, 0.79, 0.73, 0.74, 0.74, 0.83, 0.95, 0.89, 
    0.95, 0.88, 0.8, 0.81, 0.68, 0.63, 0.66, 0.61, 0.65, 0.58, 0.61, 0.58, 
    0.58, 0.57, 0.56, 0.57, 0.6, 0.62, 0.59, 0.56, 0.53, 0.5, 0.52, 0.56, 
    0.65, 0.67, 0.7, 0.69, 0.7, 0.65, 0.7, 0.67, 0.66, 0.7, 0.65, 0.66, 0.61, 
    0.73, 0.72, 0.7, 0.68, 0.68, 0.71, 0.81, 0.82, 0.85, 0.84, 0.83, 0.78, 
    0.85, 0.82, 0.94, 0.7, 0.72, 0.69, 0.66, 0.66, 0.67, 0.63, 0.66, 0.66, 
    0.65, 0.7, 0.63, 0.68, 0.68, 0.71, 0.74, 0.83, 0.77, 0.71, 0.69, 0.73, 
    0.75, 0.73, 0.75, 0.69, 0.65, 0.73, 0.78, 0.64, 0.61, 0.56, 0.62, 0.64, 
    0.73, 0.67, 0.71, 0.94, 0.96, 0.95, 0.94, 0.97, 1, 1, 0.97, 0.71, 0.71, 
    0.69, 0.73, 0.71, 0.71, 0.66, 0.65, 0.74, 0.75, 0.67, 0.66, 0.69, 0.67, 
    0.64, 0.68, 0.67, 0.67, 0.83, 0.87, 0.85, 0.78, 0.72, 0.7, 0.75, 0.79, 
    0.82, 0.83, 0.88, 0.92, 0.85, 0.71, 0.68, 0.84, 0.92, 0.9, 0.94, 0.88, 
    0.67, 0.69, 0.76, 0.75, 0.71, 0.77, 0.8, 0.82, 0.86, 0.83, 0.78, 0.78, 
    0.73, 0.71, 0.76, 0.75, 0.8, 0.79, 0.76, 0.8, 0.72, 0.72, 0.62, 0.61, 
    0.6, 0.72, 0.75, 0.81, 0.81, 0.69, 0.75, 0.7, 0.67, 0.7, 0.61, 0.63, 
    0.67, 0.69, 0.75, 0.82, 0.78, 0.74, 0.8, 0.77, 0.67, 0.7, 0.7, 0.64, 
    0.61, 0.66, 0.61, 0.71, 0.84, 0.9, 0.92, 0.87, 0.93, 0.94, 0.88, 0.84, 
    0.85, 0.83, 0.8, 0.76, 0.7, 0.74, 0.72, 0.69, 0.67, 0.66, 0.66, 0.67, 
    0.76, 0.83, 0.91, 0.97, 0.98, 1, 0.99, 1, 1, 1, 1, 1, 1, 0.98, 0.97, 
    0.91, 0.91, 0.82, 0.74, 0.71, 0.75, 0.75, 0.76, 0.76, 0.77, 0.76, 0.78, 
    0.77, 0.77, 0.77, 0.77, 0.8, 0.92, 0.91, 0.92, 0.83, 0.81, 0.81, 0.87, 
    0.87, 0.86, 0.77, 0.81, 0.79, 0.88, 0.93, 0.95, 0.97, 0.74, 0.73, 0.67, 
    0.69, 0.68, 0.62, 0.62, 0.65, 0.65, 0.68, 0.66, 0.59, 0.62, 0.66, 0.67, 
    0.69, 0.68, 0.69, 0.63, 0.62, 0.71, 0.68, 0.74, 0.73, 0.65, 0.63, 0.68, 
    0.64, 0.66, 0.68, 0.7, 0.74, 0.72, 0.77, 0.76, 0.82, 0.76, 0.79, 0.74, 
    0.75, 0.76, 0.78, 0.75, 0.72, 0.76, 0.7, 0.76, 0.74, 0.7, 0.71, 0.7, 
    0.71, 0.73, 0.74, 0.77, 0.8, 0.77, 0.79, 0.81, 0.82, 0.81, 0.76, 0.82, 
    0.76, 0.82, 0.85, 0.82, 0.78, 0.84, 0.88, 0.87, 0.85, 0.89, 0.92, 0.9, 
    0.92, 0.95, 0.94, 0.96, 0.98, 0.76, 0.69, 0.68, 0.68, 0.68, 0.64, 0.65, 
    0.66, 0.64, 0.63, 0.65, 0.66, 0.66, 0.66, 0.73, 0.73, 0.7, 0.67, 0.64, 
    0.74, 0.73, 0.67, 0.69, 0.65, 0.66, 0.69, 0.67, 0.66, 0.68, 0.65, 0.63, 
    0.66, 0.66, 0.72, 0.66, 0.71, 0.72, 0.72, 0.72, 0.72, 0.68, 0.64, 0.63, 
    0.69, 0.73, 0.66, 0.65, 0.66, 0.68, 0.66, 0.66, 0.66, 0.67, 0.62, 0.64, 
    0.65, 0.69, 0.71, 0.71, 0.68, 0.64, 0.65, 0.63, 0.63, 0.67, 0.65, 0.63, 
    0.66, 0.76, 0.82, 0.82, 0.77, 0.79, 0.79, 0.8, 0.76, 0.86, 0.77, 0.78, 
    0.8, 0.87, 0.82, 0.92, 0.87, 0.86, 0.77, 0.86, 0.75, 0.8, 0.79, 0.69, 
    0.66, 0.58, 0.64, 0.59, 0.69, 0.64, 0.59, 0.64, 0.57, 0.61, 0.6, 0.63, 
    0.57, 0.54, 0.56, 0.57, 0.59, 0.58, 0.58, 0.63, 0.64, 0.62, 0.64, 0.66, 
    0.64, 0.66, 0.7, 0.69, 0.68, 0.68, 0.67, 0.71, 0.68, 0.72, 0.68, 0.66, 
    0.68, 0.71, 0.68, 0.68, 0.69, 0.67, 0.66, 0.71, 0.72, 0.72, 0.72, 0.74, 
    0.74, 0.76, 0.69, 0.71, 0.76, 0.75, 0.74, 0.74, 0.78, 0.76, 0.76, 0.77, 
    0.75, 0.73, 0.78, 0.79, 0.79, 0.63, 0.53, 0.58, 0.54, 0.58, 0.68, 0.71, 
    0.74, 0.75, 0.82, 0.99, 1, 1, 0.94, 0.85, 0.78, 0.8, 0.88, 0.93, 0.85, 
    0.86, 0.92, 0.92, 0.83, 0.79, 0.74, 0.74, 0.74, 0.79, 0.76, 0.73, 0.77, 
    0.89, 0.94, 0.96, 0.98, 0.99, 0.99, 0.98, 0.97, 0.91, 0.85, 0.94, 0.91, 
    0.78, 0.74, 0.71, 0.71, 0.73, 0.71, 0.68, 0.7, 0.67, 0.65, 0.62, 0.66, 
    0.64, 0.64, 0.61, 0.6, 0.61, 0.64, 0.65, 0.66, 0.61, 0.61, 0.61, 0.61, 
    0.61, 0.61, 0.62, 0.61, 0.56, 0.56, 0.51, 0.49, 0.49, 0.54, 0.52, 0.49, 
    0.51, 0.5, 0.54, 0.53, 0.57, 0.57, 0.63, 0.6, 0.63, 0.67, 0.71, 0.73, 
    0.76, 0.78, 0.64, 0.64, 0.66, 0.61, 0.67, 0.63, 0.63, 0.62, 0.64, 0.72, 
    0.64, 0.66, 0.66, 0.69, 0.68, 0.7, 0.66, 0.71, 0.76, 0.74, 0.88, 0.82, 
    0.83, 0.83, 0.78, 0.8, 0.79, 0.73, 0.71, 0.76, 0.75, 0.77, 0.79, 0.78, 
    0.81, 0.8, 0.68, 0.71, 0.66, 0.69, 0.69, 0.61, 0.71, 0.68, 0.7, 0.73, 
    0.73, 0.72, 0.69, 0.68, 0.66, 0.68, 0.68, 0.65, 0.58, 0.59, 0.58, 0.58, 
    0.57, 0.58, 0.59, 0.62, 0.62, 0.7, 0.74, 0.76, 0.84, 0.81, 0.83, 0.83, 
    0.85, 0.91, 0.85, 0.85, 0.9, 0.91, 0.9, 0.89, 0.8, 0.69, 0.71, 0.8, 0.73, 
    0.76, 0.75, 0.76, 0.9, 0.88, 0.92, 0.92, 0.95, 0.93, 0.9, 0.9, 0.73, 
    0.69, 0.66, 0.62, 0.67, 0.73, 0.79, 0.76, 0.79, 0.8, 0.76, 0.77, 0.73, 
    0.71, 0.65, 0.69, 0.72, 0.79, 0.8, 0.82, 0.86, 0.82, 0.85, 0.78, 0.84, 
    0.79, 0.76, 0.77, 0.76, 0.76, 0.74, 0.78, 0.71, 0.72, 0.67, 0.7, 0.71, 
    0.71, 0.72, 0.73, 0.75, 0.82, 0.77, 0.79, 0.82, 0.84, 0.8, 0.84, 0.87, 
    0.84, 0.9, 0.88, 0.87, 0.84, 0.84, 0.79, 0.75, 0.85, 0.77, 0.78, 0.72, 
    0.75, 0.82, 0.77, 0.75, 0.72, 0.74, 0.75, 0.77, 0.8, 0.75, 0.76, 0.79, 
    0.8, 0.83, 0.79, 0.77, 0.73, 0.7, 0.7, 0.69, 0.68, 0.66, 0.68, 0.69, 
    0.71, 0.68, 0.7, 0.75, 0.73, 0.74, 0.78, 0.74, 0.77, 0.76, 0.71, 0.67, 
    0.63, 0.64, 0.63, 0.6, 0.65, 0.66, 0.65, 0.63, 0.64, 0.64, 0.57, 0.56, 
    0.63, 0.61, 0.68, 0.71, 0.73, 0.73, 0.74, 0.74, 0.74, 0.71, 0.71, 0.67, 
    0.64, 0.64, 0.6, 0.59, 0.6, 0.57, 0.54, 0.54, 0.57, 0.58, 0.61, 0.57, 
    0.61, 0.55, 0.58, 0.56, 0.56, 0.55, 0.55, 0.56, 0.56, 0.56, 0.55, 0.52, 
    0.54, 0.54, 0.54, 0.54, 0.52, 0.56, 0.56, 0.56, 0.56, 0.56, 0.6, 0.61, 
    0.59, 0.59, 0.6, 0.58, 0.6, 0.59, 0.61, 0.62, 0.58, 0.6, 0.56, 0.58, 
    0.59, 0.6, 0.53, 0.6, 0.6, 0.61, 0.59, 0.57, 0.59, 0.56, 0.56, 0.51, 
    0.54, 0.54, 0.52, 0.54, 0.54, 0.55, 0.54, 0.59, 0.56, 0.6, 0.6, 0.56, 
    0.56, 0.55, 0.52, 0.5, 0.51, 0.57, 0.6, 0.56, 0.58, 0.53, 0.56, 0.56, 
    0.54, 0.58, 0.62, 0.64, 0.63, 0.63, 0.66, 0.69, 0.7, 0.7, 0.7, 0.69, 
    0.67, 0.66, 0.65, 0.62, 0.62, 0.61, 0.61, 0.63, 0.64, 0.65, 0.62, 0.64, 
    0.65, 0.63, 0.64, 0.65, 0.66, 0.66, 0.64, 0.62, 0.63, 0.66, 0.65, 0.64, 
    0.64, 0.58, 0.63, 0.67, 0.64, 0.62, 0.65, 0.64, 0.75, 0.67, 0.64, 0.63, 
    0.65, 0.64, 0.64, 0.6, 0.6, 0.62, 0.63, 0.62, 0.59, 0.55, 0.52, 0.52, 
    0.56, 0.55, 0.54, 0.61, 0.57, 0.55, 0.57, 0.56, 0.55, 0.56, 0.54, 0.56, 
    0.6, 0.52, 0.57, 0.58, 0.58, 0.56, 0.57, 0.63, 0.79, 0.8, 0.76, 0.68, 
    0.68, 0.74, 0.72, 0.64, 0.54, 0.59, 0.6, 0.55, 0.54, 0.52, 0.52, 0.53, 
    0.54, 0.54, 0.59, 0.62, 0.61, 0.66, 0.73, 0.73, 0.75, 0.76, 0.76, 0.75, 
    0.76, 0.74, 0.68, 0.72, 0.74, 0.76, 0.8, 0.83, 0.9, 0.96, 0.98, 0.94, 
    0.97, 0.96, 0.97, 0.95, 0.8, 0.8, 0.8, 0.79, 0.81, 0.88, 0.89, 0.77, 
    0.76, 0.78, 0.7, 0.65, 0.62, 0.58, 0.6, 0.61, 0.61, 0.6, 0.54, 0.58, 
    0.63, 0.59, 0.69, 0.62, 0.66, 0.65, 0.67, 0.74, 0.67, 0.66, 0.62, 0.6, 
    0.56, 0.5, 0.51, 0.51, 0.56, 0.58, 0.55, 0.51, 0.57, 0.67, 0.62, 0.53, 
    0.54, 0.59, 0.65, 0.66, 0.62, 0.6, 0.65, 0.69, 0.72, 0.74, 0.73, 0.81, 
    0.79, 0.73, 0.71, 0.71, 0.68, 0.68, 0.71, 0.7, 0.7, 0.69, 0.64, 0.66, 
    0.68, 0.68, 0.75, 0.69, 0.71, 0.68, 0.72, 0.72, 0.74, 0.73, 0.71, 0.75, 
    0.77, 0.79, 0.78, 0.77, 0.94, 1, 0.9, 0.8, 0.81, 0.75, 0.74, 0.79, 0.8, 
    0.77, 0.78, 0.8, 0.78, 0.73, 0.73, 0.73, 0.71, 0.69, 0.71, 0.71, 0.68, 
    0.64, 0.59, 0.58, 0.59, 0.57, 0.58, 0.54, 0.53, 0.69, 0.62, 0.55, 0.65, 
    0.61, 0.62, 0.67, 0.71, 0.66, 0.61, 0.62, 0.51, 0.53, 0.42, 0.51, 0.62, 
    0.6, 0.71, 0.74, 0.68, 0.63, 0.62, 0.61, 0.63, 0.6, 0.58, 0.61, 0.6, 
    0.65, 0.66, 0.68, 0.7, 0.68, 0.73, 0.7, 0.78, 0.75, 0.78, 0.74, 0.71, 
    0.75, 0.75, 0.81, 0.78, 0.85, 0.89, 0.9, 0.88, 0.87, 0.83, 0.75, 0.82, 
    0.82, 0.8, 0.85, 0.82, 0.78, 0.79, 0.8, 0.8, 0.79, 0.77, 0.72, 0.71, 0.7, 
    0.69, 0.76, 0.68, 0.68, 0.78, 0.75, 0.76, 0.75, 0.79, 0.64, 0.65, 0.65, 
    0.66, 0.75, 0.7, 0.82, 0.8, 0.92, 0.95, 0.95, 0.9, 0.88, 0.8, 0.8, 0.81, 
    0.77, 0.81, 0.81, 0.92, 0.83, 0.9, 0.96, 0.85, 0.73, 0.75, 0.82, 0.7, 
    0.75, 0.88, 0.73, 0.86, 0.95, 0.81, 0.75, 0.77, 0.83, 0.82, 0.8, 0.76, 
    0.8, 0.84, 0.83, 0.77, 0.75, 0.82, 0.77, 0.72, 0.68, 0.69, 0.6, 0.55, 
    0.69, 0.66, 0.73, 0.62, 0.45, 0.47, 0.36, 0.62, 0.68, 0.71, 0.72, 0.78, 
    0.8, 0.82, 0.84, 0.84, 0.89, 0.87, 0.83, 0.83, 0.83, 0.8, 0.84, 0.8, 0.8, 
    0.82, 0.82, 0.82, 1, 1, 1, 1, 1, 1, 0.98, 1, 1, 0.97, 0.95, 0.85, 0.9, 
    0.94, 0.88, 0.95, 0.93, 0.79, 0.93, 0.99, 1, 0.94, 1, 1, 1, 1, 1, 1, 1, 
    0.97, 0.94, 0.9, 0.82, 0.86, 0.82, 0.78, 0.75, 0.79, 0.84, 0.77, 0.75, 
    0.7, 0.72, 0.71, 0.72, 0.73, 0.77, 0.76, 0.8, 0.98, 0.93, 0.83, 0.74, 
    0.68, 0.76, 0.77, 0.74, 0.73, 0.72, 0.77, 0.86, 0.82, 0.78, 0.79, 0.75, 
    0.73, 0.7, 0.69, 0.68, 0.67, 0.71, 0.71, 0.69, 0.7, 0.71, 0.72, 0.71, 
    0.69, 0.73, 0.7, 0.72, 0.78, 0.8, 0.76, 0.72, 0.75, 0.74, 0.74, 0.72, 
    0.7, 0.7, 0.74, 0.78, 0.77, 0.77, 0.72, 0.72, 0.72, 0.66, 0.69, 0.7, 
    0.73, 0.7, 0.68, 0.66, 0.62, 0.63, 0.62, 0.67, 0.64, 0.64, 0.64, 0.63, 
    0.61, 0.61, 0.62, 0.64, 0.64, 0.65, 0.66, 0.65, 0.67, 0.63, 0.65, 0.66, 
    0.63, 0.61, 0.62, 0.73, 0.76, 0.69, 0.73, 0.78, 0.68, 0.69, 0.71, 0.73, 
    0.79, 0.82, 0.92, 0.92, 0.8, 0.83, 0.83, 0.82, 0.87, 0.82, 0.83, 0.86, 
    0.82, 0.78, 0.75, 0.81, 0.86, 0.81, 0.79, 0.74, 0.81, 0.82, 0.81, 0.83, 
    0.88, 0.85, 0.93, 0.93, 0.92, 0.91, 0.92, 0.91, 0.91, 0.9, 0.89, 0.85, 
    0.85, 0.76, 0.76, 0.78, 0.76, 0.82, 0.84, 0.83, 0.8, 0.81, 0.82, 0.84, 
    0.88, 1, 0.98, 0.89, 0.93, 0.93, 0.93, 0.95, 0.98, 0.89, 0.83, 0.8, 0.79, 
    0.71, 0.7, 0.65, 0.64, 0.63, 0.65, 0.67, 0.66, 0.71, 0.69, 0.62, 0.61, 
    0.59, 0.56, 0.61, 0.66, 0.64, 0.62, 0.57, 0.62, 0.71, 0.84, 0.81, 0.76, 
    0.81, 0.79, 0.79, 0.79, 0.8, 0.82, 0.82, 0.83, 0.79, 0.78, 0.77, 0.76, 
    0.79, 0.84, 0.85, 0.75, 0.82, 0.79, 0.78, 0.8, 0.82, 0.91, 0.79, 0.85, 
    0.84, 0.85, 0.96, 0.99, 1, 1, 1, 0.94, 0.83, 0.87, 0.84, 0.72, 0.74, 
    0.79, 0.74, 0.72, 0.69, 0.69, 0.82, 0.82, 0.89, 0.91, 0.9, 0.79, 0.81, 
    0.86, 0.68, 0.69, 0.76, 0.73, 0.69, 0.65, 0.64, 0.64, 0.6, 0.55, 0.65, 
    0.61, 0.63, 0.6, 0.61, 0.63, 0.58, 0.57, 0.53, 0.52, 0.66, 0.71, 0.67, 
    0.63, 0.72, 0.71, 0.7, 0.66, 0.62, 0.75, 0.72, 0.75, 0.76, 0.78, 0.73, 
    0.76, 0.77, 0.8, 0.82, 0.67, 0.7, 0.68, 0.68, 0.67, 0.68, 0.67, 0.69, 
    0.67, 0.66, 0.61, 0.72, 0.69, 0.68, 0.79, 0.73, 0.81, 0.82, 0.89, 0.82, 
    0.94, 0.89, 0.88, 0.9, 0.9, 0.8, 0.85, 0.77, 0.77, 0.79, 0.78, 0.77, 
    0.73, 0.73, 0.75, 0.91, 0.93, 0.83, 0.79, 0.78, 0.77, 0.81, 0.85, 0.98, 
    0.82, 0.89, 0.94, 0.85, 1, 1, 1, 1, 1, 1, 1, 0.92, 0.84, 0.84, 0.82, 
    0.84, 0.81, 0.79, 0.74, 0.81, 0.8, 0.78, 0.8, 0.8, 0.8, 0.88, 0.86, 0.81, 
    0.84, 0.82, 0.79, 0.8, 0.8, 0.83, 0.81, 0.74, 0.77, 0.79, 0.74, 0.77, 
    0.87, 0.79, 0.75, 0.77, 0.77, 0.75, 0.75, 0.77, 0.76, 0.81, 0.87, 0.79, 
    0.87, 0.9, 0.89, 0.83, 0.9, 0.82, 0.89, 0.87, 0.85, 0.81, 0.89, 0.9, 
    0.96, 0.87, 0.78, 0.79, 0.82, 0.81, 0.79, 0.78, 0.75, 0.75, 0.75, 0.77, 
    0.76, 0.84, 0.83, 0.82, 0.81, 0.79, 0.71, 0.67, 0.71, 0.72, 0.73, 0.71, 
    0.66, 0.67, 0.78, 0.78, 0.8, 0.84, 0.71, 0.76, 0.78, 0.77, 0.79, 0.78, 
    0.81, 0.84, 0.8, 0.79, 0.82, 0.76, 0.81, 0.8, 0.76, 0.78, 0.78, 0.82, 
    0.73, 0.75, 0.75, 0.81, 0.79, 0.94, 0.86, 0.74, 0.69, 0.69, 0.78, 0.77, 
    0.76, 0.82, 0.81, 0.86, 0.8, 0.77, 0.62, 0.59, 0.56, 0.55, 0.59, 0.56, 
    0.57, 0.56, 0.61, 0.61, 0.61, 0.66, 0.7, 0.64, 0.65, 0.69, 0.77, 0.91, 
    0.96, 0.98, 0.97, 0.91, 0.89, 0.84, 0.8, 0.72, 0.72, 0.69, 0.67, 0.67, 
    0.64, 0.64, 0.65, 0.58, 0.62, 0.61, 0.64, 0.65, 0.65, 0.66, 0.69, 0.69, 
    0.75, 0.77, 0.77, 0.78, 0.77, 0.8, 0.82, 0.77, 0.79, 0.75, 0.73, 0.76, 
    0.76, 0.76, 0.72, 0.67, 0.68, 0.74, 0.79, 0.82, 0.86, 0.82, 0.79, 0.79, 
    0.8, 0.8, 0.78, 0.75, 0.73, 0.71, 0.72, 0.71, 1, 0.65, 0.64, 0.66, 0.68, 
    0.67, 0.67, 1, 0.7, 0.72, 0.66, 0.69, 0.73, 0.83, 0.82, 0.83, 0.88, 0.91, 
    0.86, 0.86, 0.88, 0.89, 0.84, 0.8, 0.84, 0.82, 0.72, 0.72, 0.79, 0.75, 
    0.71, 0.66, 0.8, 0.76, 0.93, 0.82, 0.91, 0.85, 0.91, 0.85, 0.86, 0.89, 
    0.85, 0.81, 0.78, 0.8, 0.76, 0.94, 0.95, 0.79, 0.89, 0.85, 0.84, 0.85, 
    0.86, 0.95, 0.81, 1, 0.98, 1, 0.99, 1, 1, 1, 0.78, 0.77, 0.79, 0.84, 
    0.87, 0.91, 0.88, 0.82, 0.88, 0.98, 0.87, 0.78, 0.77, 0.77, 0.77, 0.78, 
    0.82, 0.78, 0.8, 0.81, 0.82, 0.82, 0.84, 0.85, 0.81, 0.78, 0.75, 0.78, 
    0.78, 0.79, 0.79, 0.79, 0.79, 0.8, 0.64, 0.65, 0.72, 0.73, 0.73, 0.71, 
    0.64, 0.7, 0.66, 0.74, 0.74, 0.73, 0.76, 0.75, 0.79, 0.76, 0.76, 0.84, 
    0.79, 0.81, 0.85, 0.81, 0.81, 0.8, 0.79, 0.77, 0.77, 0.77, 0.79, 0.79, 
    0.82, 0.75, 0.66, 0.67, 0.66, 0.68, 0.72, 0.69, 0.69, 0.67, 0.7, 0.68, 
    0.73, 0.74, 0.79, 0.81, 0.78, 0.78, 0.85, 0.86, 0.81, 0.75, 0.73, 0.78, 
    0.73, 0.75, 0.79, 0.76, 0.73, 0.72, 0.73, 0.78, 0.87, 0.78, 0.75, 0.73, 
    0.7, 0.67, 0.72, 0.85, 0.67, 0.67, 0.73, 0.69, 0.75, 0.73, 0.78, 0.79, 
    0.79, 0.77, 0.75, 0.75, 0.91, 0.83, 0.77, 0.85, 0.97, 0.98, 1, 1, 1, 1, 
    0.84, 0.85, 0.75, 0.71, 0.76, 0.81, 0.74, 0.71, 0.68, 0.75, 0.74, 0.75, 
    0.8, 0.8, 0.79, 0.81, 0.79, 0.88, 0.79, 0.75, 0.74, 0.8, 0.84, 0.81, 
    0.81, 0.73, 0.68, 0.66, 0.66, 0.67, 0.7, 0.61, 0.67, 0.69, 0.72, 0.72, 
    0.79, 0.85, 0.86, 0.9, 0.96, 1, 1, 1, 1, 1, 1, 1, 1, 0.96, 0.95, 0.95, 
    0.9, 0.93, 0.85, 0.91, 0.89, 0.9, 0.94, 0.93, 0.91, 0.91, 0.92, 0.93, 
    0.86, 0.91, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.98, 1, 0.9, 0.96, 0.91, 
    0.94, 0.97, 0.97, 0.94, 0.9, 0.87, 0.83, 0.85, 0.8, 0.82, 0.77, 0.89, 
    0.86, 0.83, 0.77, 0.82, 0.77, 0.59, 0.65, 0.63, 0.69, 0.68, 0.74, 0.67, 
    0.65, 0.66, 0.64, 0.69, 0.7, 0.76, 0.74, 0.78, 0.77, 0.77, 0.77, 0.75, 
    0.75, 0.8, 0.78, 0.75, 0.71, 0.69, 0.65, 0.68, 0.57, 0.58, 0.67, 0.69, 
    0.68, 0.69, 0.84, 0.69, 0.8, 0.85, 0.87, 0.86, 0.81, 0.78, 1, 1, 0.98, 
    0.94, 0.91, 0.86, 0.86, 0.87, 0.78, 0.83, 0.78, 0.73, 0.71, 0.68, 0.7, 
    0.62, 0.63, 0.74, 0.73, 0.72, 0.74, 0.7, 0.73, 0.73, 0.72, 0.71, 0.66, 
    0.66, 0.69, 0.68, 0.67, 0.66, 0.67, 0.7, 0.67, 0.66, 0.74, 0.8, 0.81, 
    0.84, 0.92, 1, 0.99, 1, 0.77, 0.95, 0.98, 0.93, 0.92, 0.98, 1, 0.91, 
    0.82, 0.81, 0.81, 0.81, 0.85, 0.83, 0.88, 0.86, 0.91, 0.89, 0.88, 0.84, 
    0.86, 0.8, 0.86, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.95, 0.9, 0.93, 0.82, 
    0.8, 0.8, 0.79, 0.74, 0.74, 0.79, 0.9, 0.8, 0.8, 0.85, 0.82, 0.85, 0.88, 
    0.86, 0.87, 0.79, 0.77, 0.75, 0.75, 0.74, 0.72, 0.68, 0.67, 0.61, 0.57, 
    0.51, 0.56, 0.59, 0.56, 0.62, 0.63, 0.64, 0.73, 0.76, 0.8, 0.82, 0.88, 
    0.92, 0.84, 0.79, 0.73, 0.69, 0.6, 0.61, 0.62, 0.59, 0.6, 0.6, 0.64, 
    0.69, 0.66, 0.64, 0.64, 0.65, 0.62, 0.61, 0.53, 0.5, 0.57, 0.49, 0.54, 
    0.55, 0.51, 0.55, 0.62, 0.68, 0.64, 0.68, 0.64, 0.71, 0.63, 0.63, 0.65, 
    0.72, 0.75, 0.72, 0.75, 0.74, 0.73, 0.75, 0.71, 0.69, 0.7, 0.74, 0.73, 
    0.71, 0.72, 0.72, 0.74, 0.71, 0.68, 0.7, 0.71, 0.7, 0.72, 0.73, 0.72, 
    0.71, 0.71, 0.71, 0.69, 0.7, 0.79, 0.92, 0.94, 0.96, 0.96, 0.96, 0.95, 
    0.89, 0.94, 0.98, 1, 1, 1, 1, 1, 0.91, 0.89, 0.88, 0.83, 0.84, 0.83, 
    0.81, 0.8, 0.8, 0.71, 0.73, 0.72, 0.75, 0.71, 0.72, 0.75, 0.86, 0.9, 1, 
    1, 0.99, 0.98, 1, 0.86, 0.88, 0.86, 0.84, 0.91, 0.86, 0.81, 0.81, 0.86, 
    0.83, 0.81, 0.8, 0.8, 0.79, 0.75, 0.79, 0.81, 0.83, 0.83, 0.74, 0.77, 
    0.77, 0.79, 0.79, 0.8, 0.79, 0.76, 0.78, 0.75, 0.77, 0.81, 0.76, 0.78, 
    0.77, 0.74, 0.75, 0.75, 0.71, 0.71, 0.71, 0.73, 0.72, 0.73, 0.74, 0.75, 
    0.75, 0.78, 0.77, 0.74, 0.72, 0.7, 0.68, 0.67, 0.65, 0.63, 0.63, 0.67, 
    0.68, 0.7, 0.7, 0.72, 0.72, 0.74, 0.74, 0.76, 0.75, 0.76, 0.79, 0.79, 
    0.78, 0.74, 0.72, 0.7, 0.72, 0.69, 0.69, 0.69, 0.69, 0.7, 0.69, 0.68, 
    0.69, 0.71, 0.74, 0.76, 0.78, 0.81, 0.88, 0.9, 0.9, 0.88, 0.94, 0.92, 
    0.88, 0.86, 0.87, 0.88, 0.88, 0.89, 0.95, 0.94, 0.93, 0.93, 0.98, 0.94, 
    0.94, 0.96, 0.95, 0.92, 0.91, 0.9, 0.88, 0.87, 0.86, 0.83, 0.82, 0.84, 
    0.79, 0.78, 0.85, 0.86, 0.89, 0.91, 0.88, 0.78, 0.72, 0.8, 0.81, 0.74, 
    0.67, 0.66, 0.68, 0.68, 0.68, 0.69, 0.71, 0.76, 0.82, 0.79, 0.73, 0.68, 
    0.74, 0.72, 0.76, 0.75, 0.72, 0.74, 0.76, 0.74, 0.75, 0.79, 0.83, 0.82, 
    0.79, 0.84, 0.82, 0.88, 0.95, 0.93, 0.93, 0.7, 0.64, 0.61, 0.61, 0.64, 
    0.64, 0.61, 0.63, 0.61, 0.63, 0.63, 0.61, 0.64, 0.63, 0.65, 0.74, 0.73, 
    0.7, 0.72, 0.76, 0.82, 0.73, 0.7, 0.71, 0.63, 0.6, 0.57, 0.58, 0.59, 0.6, 
    0.6, 0.66, 0.85, 0.95, 0.92, 0.95, 0.85, 0.77, 0.77, 0.77, 0.84, 0.89, 
    0.91, 0.94, 0.93, 0.99, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.96, 0.9, 0.89, 0.92, 
    0.79, 0.74, 0.8, 0.86, 0.89, 0.92, 0.87, 0.84, 0.85, 0.85, 0.86, 0.79, 
    0.81, 0.83, 0.85, 0.86, 0.84, 0.83, 0.82, 0.77, 0.76, 0.74, 0.73, 0.66, 
    0.65, 0.62, 0.67, 0.64, 0.63, 0.67, 0.69, 0.69, 0.68, 0.7, 0.78, 0.84, 
    0.86, 0.71, 0.76, 0.85, 0.73, 0.71, 0.68, 0.66, 0.65, 0.6, 0.67, 0.57, 
    0.56, 0.59, 0.6, 0.61, 0.61, 0.65, 0.7, 0.64, 0.69, 0.68, 0.68, 0.69, 
    0.67, 0.7, 0.7, 0.7, 0.64, 0.69, 0.74, 0.74, 0.66, 0.64, 0.62, 0.66, 
    0.68, 0.63, 0.62, 0.69, 0.67, 0.66, 0.64, 0.63, 0.66, 0.66, 0.65, 0.72, 
    0.76, 0.78, 0.73, 0.71, 0.75, 0.7, 0.76, 0.78, 0.77, 0.73, 0.74, 0.67, 
    0.62, 0.6, 0.63, 0.57, 0.49, 0.46, 0.49, 0.5, 0.62, 0.58, 0.57, 0.51, 
    0.55, 0.63, 0.62, 0.65, 0.71, 0.7, 0.65, 0.72, 0.67, 0.62, 0.61, 0.57, 
    0.56, 0.59, 0.58, 0.6, 0.59, 0.58, 0.61, 0.61, 0.62, 0.62, 0.69, 0.68, 
    0.66, 0.67, 0.77, 0.67, 0.71, 0.7, 0.63, 0.6, 0.6, 0.65, 0.57, 0.63, 
    0.67, 0.64, 0.64, 0.64, 0.63, 0.64, 0.62, 0.61, 0.58, 0.58, 0.57, 0.56, 
    0.56, 0.67, 0.67, 0.64, 0.69, 0.57, 0.57, 0.61, 0.57, 0.56, 0.57, 0.55, 
    0.56, 0.56, 0.57, 0.61, 0.55, 0.57, 0.61, 0.63, 0.67, 0.72, 0.8, 0.86, 
    0.82, 0.88, 0.86, 0.88, 0.85, 0.85, 0.84, 0.77, 0.8, 0.69, 0.6, 0.58, 
    0.62, 0.66, 0.65, 0.63, 0.62, 0.63, 0.67, 0.64, 0.67, 0.72, 0.75, 0.76, 
    0.78, 0.8, 0.79, 0.8, 0.82, 0.78, 0.78, 0.71, 0.78, 0.77, 0.76, 0.79, 
    0.73, 0.67, 0.52, 0.53, 0.54, 0.54, 0.65, 0.63, 0.68, 0.69, 0.72, 0.74, 
    0.76, 0.79, 0.83, 0.84, 0.82, 0.77, 0.85, 0.82, 0.8, 0.84, 0.84, 0.87, 
    0.87, 0.9, 0.91, 0.88, 0.86, 0.85, 0.82, 0.84, 0.86, 0.86, 0.76, 0.72, 
    0.71, 0.74, 0.73, 0.75, 0.76, 0.78, 0.79, 0.76, 0.85, 0.8, 0.88, 0.86, 
    0.84, 0.78, 0.73, 0.76, 0.73, 0.67, 0.75, 0.79, 0.77, 0.79, 0.78, 0.79, 
    0.77, 0.77, 0.74, 0.74, 0.74, 0.76, 0.74, 0.75, 0.72, 0.64, 0.61, 0.52, 
    0.52, 0.55, 0.52, 0.54, 0.56, 0.59, 0.62, 0.69, 0.67, 0.71, 0.67, 0.7, 
    0.71, 0.69, 0.73, 0.82, 0.92, 0.93, 0.93, 0.92, 0.92, 0.9, 0.88, 0.89, 
    0.89, 0.91, 0.92, 0.96, 0.95, 0.93, 0.93, 0.95, 0.95, 0.93, 0.91, 0.91, 
    0.92, 0.88, 0.81, 0.78, 0.77, 0.81, 0.72, 0.76, 0.78, 0.78, 0.81, 0.86, 
    0.85, 0.9, 0.83, 0.9, 0.9, 0.91, 0.91, 0.93, 0.87, 0.92, 0.94, 0.91, 
    0.93, 0.94, 0.94, 0.88, 0.84, 0.88, 0.88, 0.88, 0.87, 0.81, 0.73, 0.73, 
    0.65, 0.58, 0.6, 0.59, 0.58, 0.6, 0.69, 0.71, 0.7, 0.74, 0.79, 0.77, 
    0.78, 0.83, 0.81, 0.85, 0.85, 0.81, 0.84, 0.87, 0.82, 0.83, 0.8, 0.75, 
    0.73, 0.81, 0.79, 0.91, 0.92, 0.8, 0.69, 0.78, 0.8, 0.78, 0.77, 0.79, 
    0.76, 0.74, 0.79, 0.78, 0.78, 0.84, 0.79, 0.74, 0.74, 0.76, 0.88, 0.81, 
    0.77, 0.74, 0.78, 0.77, 0.76, 0.76, 0.82, 0.8, 0.79, 0.84, 0.85, 0.85, 
    0.89, 0.87, 0.73, 0.72, 0.73, 0.74, 0.75, 0.73, 0.75, 0.73, 0.7, 0.75, 
    0.71, 0.78, 0.74, 0.69, 0.73, 0.69, 0.66, 0.67, 0.72, 0.73, 0.75, 0.76, 
    0.72, 0.71, 0.71, 0.73, 0.71, 0.68, 0.72, 0.75, 0.74, 0.81, 0.92, 0.86, 
    0.82, 0.85, 0.82, 0.78, 0.79, 0.8, 0.82, 0.81, 0.81, 0.78, 0.8, 0.8, 
    0.75, 0.77, 0.76, 0.8, 0.83, 0.82, 0.84, 0.84, 0.8, 0.8, 0.82, 0.84, 
    0.89, 0.88, 0.91, 0.94, 0.95, 0.9, 0.79, 0.83, 0.88, 0.94, 0.84, 0.85, 
    0.83, 0.85, 0.92, 0.91, 0.92, 0.84, 0.83, 0.83, 0.83, 0.75, 0.71, 0.73, 
    0.77, 0.72, 0.74, 0.75, 0.8, 0.81, 0.83, 0.85, 0.85, 0.87, 0.9, 0.92, 
    0.92, 0.93, 0.93, 0.94, 0.89, 0.94, 0.94, 0.82, 0.9, 0.87, 0.85, 0.86, 
    0.84, 0.83, 0.88, 0.86, 0.87, 0.86, 0.82, 0.82, 0.83, 0.85, 0.9, 0.9, 
    0.87, 0.88, 0.86, 0.87, 0.88, 0.82, 0.74, 0.74, 0.71, 0.67, 0.69, 0.68, 
    0.67, 0.66, 0.68, 0.68, 0.67, 0.7, 0.69, 0.69, 0.73, 0.69, 0.63, 0.62, 
    0.64, 0.67, 0.64, 0.62, 0.66, 0.54, 0.5, 0.48, 0.51, 0.42, 0.53, 0.51, 
    0.57, 0.45, 0.52, 0.51, 0.55, 0.52, 0.59, 0.56, 0.56, 0.55, 0.61, 0.62, 
    0.6, 0.6, 0.55, 0.65, 0.68, 0.69, 0.65, 0.64, 0.65, 0.62, 0.65, 0.67, 
    0.71, 0.71, 0.71, 0.72, 0.7, 0.71, 0.71, 0.73, 0.75, 0.79, 0.77, 0.79, 
    0.82, 0.82, 0.79, 0.81, 0.76, 0.73, 0.69, 0.67, 0.66, 0.65, 0.6, 0.6, 
    0.62, 0.64, 0.6, 0.59, 0.59, 0.59, 0.62, 0.61, 0.63, 0.64, 0.7, 0.7, 
    0.75, 0.78, 0.82, 0.8, 0.87, 0.89, 0.87, 0.88, 0.94, 0.96, 0.94, 0.93, 
    0.86, 0.89, 0.85, 0.78, 0.76, 0.74, 0.76, 0.83, 0.81, 0.81, 0.79, 0.82, 
    0.82, 0.82, 0.8, 0.83, 0.8, 0.75, 0.74, 0.74, 0.72, 0.68, 0.67, 0.65, 
    0.63, 0.67, 0.65, 0.67, 0.69, 0.82, 0.69, 0.79, 0.82, 0.79, 0.81, 0.84, 
    0.79, 0.8, 0.82, 0.8, 0.8, 0.76, 0.74, 0.75, 0.72, 0.66, 0.64, 0.58, 
    0.59, 0.64, 0.63, 0.65, 0.82, 0.67, 0.66, 0.64, 0.64, 0.64, 0.63, 0.71, 
    0.7, 0.78, 0.75, 0.72, 0.73, 0.7, 0.73, 0.69, 0.69, 0.72, 0.7, 0.68, 
    0.63, 0.64, 0.66, 0.68, 0.71, 0.71, 0.75, 0.78, 0.77, 0.82, 0.8, 0.85, 
    0.79, 0.8, 0.8, 0.76, 0.75, 0.72, 0.72, 0.73, 0.68, 0.67, 0.68, 0.65, 
    0.64, 0.63, 0.65, 0.6, 0.61, 0.62, 0.61, 0.6, 0.74, 0.69, 0.73, 0.76, 
    0.65, 0.63, 0.65, 0.64, 0.61, 0.65, 0.61, 0.55, 0.57, 0.54, 0.55, 0.6, 
    0.61, 0.61, 0.63, 0.63, 0.65, 0.65, 0.6, 0.59, 0.6, 0.56, 0.58, 0.58, 
    0.55, 0.53, 0.52, 0.52, 0.5, 0.47, 0.48, 0.51, 0.53, 0.55, 0.53, 0.51, 
    0.51, 0.49, 0.51, 0.53, 0.55, 0.54, 0.57, 0.54, 0.52, 0.5, 0.61, 0.68, 
    0.61, 0.62, 0.65, 0.63, 0.57, 0.58, 0.55, 0.5, 0.51, 0.5, 0.52, 0.52, 
    0.53, 0.53, 0.55, 0.52, 0.55, 0.55, 0.58, 0.59, 0.52, 0.57, 0.57, 0.52, 
    0.51, 0.54, 0.62, 0.57, 0.53, 0.53, 0.51, 0.54, 0.55, 0.53, 0.54, 0.53, 
    0.54, 0.52, 0.54, 0.54, 0.53, 0.49, 0.5, 0.53, 0.52, 0.53, 0.52, 0.62, 
    0.57, 0.59, 0.58, 0.6, 0.6, 0.6, 0.61, 0.65, 0.69, 0.7, 0.75, 0.75, 0.73, 
    0.72, 0.73, 0.71, 0.77, 0.77, 0.85, 0.87, 0.87, 0.87, 0.89, 0.88, 0.9, 
    0.91, 0.92, 0.92, 0.9, 0.93, 0.94, 0.94, 0.96, 0.96, 0.97, 0.97, 0.96, 
    0.89, 0.85, 0.89, 0.92, 0.94, 0.93, 0.95, 0.94, 0.93, 0.95, 0.94, 0.93, 
    0.89, 0.89, 0.85, 0.84, 0.83, 0.74, 0.73, 0.72, 0.68, 0.61, 0.6, 0.66, 
    0.61, 0.62, 0.6, 0.62, 0.63, 0.65, 0.67, 0.66, 0.65, 0.62, 0.63, 0.62, 
    0.61, 0.61, 0.61, 0.62, 0.66, 0.64, 0.65, 0.65, 0.61, 0.64, 0.65, 0.67, 
    0.65, 0.68, 0.67, 0.71, 0.69, 0.67, 0.64, 0.63, 0.64, 0.7, 0.71, 0.7, 
    0.69, 0.68, 0.72, 0.73, 0.69, 0.72, 0.74, 0.75, 0.69, 0.68, 0.65, 0.66, 
    0.68, 0.66, 0.66, 0.66, 0.69, 0.65, 0.69, 0.71, 0.72, 0.66, 0.65, 0.73, 
    0.75, 0.75, 0.77, 0.76, 0.69, 0.7, 0.74, 0.72, 0.74, 0.68, 0.68, 0.68, 
    0.72, 0.73, 0.76, 0.72, 0.71, 0.71, 0.71, 0.7, 0.74, 0.73, 0.75, 0.68, 
    0.7, 0.72, 0.74, 0.72, 0.69, 0.69, 0.69, 0.68, 0.66, 0.67, 0.69, 0.66, 
    0.71, 0.66, 0.69, 0.71, 0.7, 0.7, 0.72, 0.72, 0.74, 0.75, 0.75, 0.79, 
    0.71, 0.71, 0.7, 0.69, 0.71, 0.73, 0.75, 0.68, 0.71, 0.64, 0.63, 0.55, 
    0.52, 0.51, 0.5, 0.55, 0.55, 0.53, 0.54, 0.52, 0.51, 0.54, 0.54, 0.54, 
    0.55, 0.58, 0.54, 0.59, 0.6, 0.61, 0.6, 0.66, 0.67, 0.67, 0.71, 0.72, 
    0.7, 0.54, 0.54, 0.57, 0.57, 0.55, 0.54, 0.58, 0.61, 0.62, 0.64, 0.63, 
    0.64, 0.63, 0.62, 0.69, 0.72, 0.73, 0.8, 0.8, 0.78, 0.75, 0.76, 0.75, 
    0.72, 0.67, 0.76, 0.71, 0.7, 0.66, 0.68, 0.62, 0.74, 0.74, 0.68, 0.69, 
    0.7, 0.68, 0.7, 0.75, 0.9, 0.91, 0.69, 0.61, 0.68, 0.72, 0.7, 0.65, 0.73, 
    0.72, 0.75, 0.77, 0.77, 0.76, 0.79, 0.79, 0.76, 0.73, 0.74, 0.74, 0.75, 
    0.77, 0.76, 0.75, 0.77, 0.78, 0.84, 0.87, 0.9, 0.9, 0.9, 0.88, 0.88, 
    0.89, 0.9, 0.91, 0.88, 0.88, 0.85, 0.88, 0.91, 0.9, 0.9, 0.91, 0.92, 
    0.91, 0.83, 0.88, 0.86, 0.83, 0.85, 0.85, 0.82, 0.76, 0.78, 0.81, 0.77, 
    0.77, 0.79, 0.81, 0.81, 0.8, 0.79, 0.81, 0.81, 0.87, 0.89, 0.92, 0.92, 
    0.91, 0.83, 0.92, 0.85, 0.85, 0.82, 0.89, 0.81, 0.78, 0.81, 0.79, 0.81, 
    0.8, 0.79, 0.83, 0.85, 0.84, 0.84, 0.84, 0.81, 0.8, 0.83, 0.78, 0.8, 
    0.82, 0.83, 0.86, 0.78, 0.77, 0.83, 0.78, 0.79, 0.76, 0.73, 0.72, 0.75, 
    0.75, 0.77, 0.8, 0.82, 0.77, 0.79, 0.82, 0.77, 0.78, 0.82, 0.81, 0.79, 
    0.82, 0.78, 0.84, 0.8, 0.78, 0.79, 0.76, 0.78, 0.78, 0.77, 0.75, 0.76, 
    0.78, 0.8, 0.77, 0.78, 0.76, 0.78, 0.82, 0.81, 0.81, 0.81, 0.79, 0.83, 
    0.73, 0.66, 0.71, 0.75, 0.69, 0.67, 0.67, 0.67, 0.69, 0.6, 0.59, 0.64, 
    0.68, 0.64, 0.68, 0.64, 0.65, 0.65, 0.66, 0.63, 0.66, 0.63, 0.68, 0.68, 
    0.69, 0.63, 0.68, 0.68, 0.83, 0.78, 0.76, 0.78, 0.79, 0.75, 0.78, 0.75, 
    0.77, 0.77, 0.78, 0.74, 0.78, 0.79, 0.79, 0.79, 0.78, 0.8, 0.79, 0.78, 
    0.76, 0.75, 0.85, 0.89, 0.93, 0.94, 0.94, 0.95, 0.96, 0.95, 0.95, 0.97, 
    0.96, 0.95, 0.96, 0.98, 0.98, 0.98, 0.95, 0.9, 0.86, 0.85, 0.86, 0.84, 
    0.8, 0.89, 0.92, 0.86, 0.84, 0.85, 0.87, 0.83, 0.76, 0.78, 0.74, 0.6, 
    0.53, 0.5, 0.51, 0.51, 0.57, 0.61, 0.69, 0.72, 0.7, 0.63, 0.7, 0.7, 0.68, 
    0.67, 0.68, 0.65, 0.67, 0.69, 0.68, 0.62, 0.68, 0.65, 0.67, 0.71, 0.78, 
    0.79, 0.85, 0.8, 0.77, 0.84, 0.9, 0.9, 0.9, 0.88, 0.83, 0.88, 0.86, 0.89, 
    0.8, 0.89, 0.79, 0.77, 0.78, 0.78, 0.78, 0.81, 0.81, 0.99, 0.86, 0.88, 
    0.89, 0.89, 0.91, 0.91, 0.88, 0.88, 0.87, 0.88, 0.85, 0.77, 0.86, 0.81, 
    0.84, 0.78, 0.71, 0.79, 0.77, 0.8, 0.82, 0.8, 0.77, 0.75, 0.77, 0.88, 
    0.85, 0.88, 0.89, 0.92, 0.93, 0.94, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 
    0.98, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.99, 0.98, 0.95, 0.95, 0.94, 
    0.89, 0.84, 0.89, 0.94, 0.9, 0.9, 0.87, 0.88, 0.83, 0.85, 0.83, 0.85, 
    0.84, 0.83, 0.84, 0.84, 0.81, 0.83, 0.81, 0.78, 0.84, 0.81, 0.83, 0.84, 
    0.83, 0.84, 0.8, 0.85, 0.81, 0.82, 0.81, 0.86, 0.83, 0.8, 0.8, 0.8, 0.85, 
    0.87, 0.86, 0.83, 0.86, 0.84, 0.81, 0.84, 0.86, 0.84, 0.85, 0.89, 0.84, 
    0.88, 0.86, 0.88, 0.87, 0.89, 0.84, 0.88, 0.87, 0.86, 0.91, 0.88, 0.86, 
    0.84, 0.87, 0.87, 0.84, 0.78, 0.78, 0.74, 0.71, 0.66, 0.69, 0.71, 0.75, 
    0.77, 0.69, 0.64, 0.67, 0.69, 0.67, 0.66, 0.69, 0.72, 0.75, 0.74, 0.73, 
    0.68, 0.71, 0.68, 0.72, 0.72, 0.72, 0.7, 0.69, 0.7, 0.69, 0.67, 0.69, 
    0.65, 0.66, 0.67, 0.65, 0.69, 0.67, 0.64, 0.59, 0.62, 0.65, 0.71, 0.66, 
    0.64, 0.71, 0.64, 0.7, 0.71, 0.69, 0.71, 0.69, 0.67, 0.66, 0.65, 0.62, 
    0.64, 0.65, 0.65, 0.64, 0.62, 0.61, 0.58, 0.64, 0.67, 0.68, 0.68, 0.68, 
    0.67, 0.67, 0.67, 0.67, 0.67, 0.68, 0.67, 0.66, 0.55, 0.59, 0.55, 0.65, 
    0.58, 0.58, 0.53, 0.57, 0.54, 0.56, 0.58, 0.57, 0.51, 0.52, 0.52, 0.58, 
    0.56, 0.55, 0.61, 0.58, 0.55, 0.52, 0.52, 0.54, 0.57, 0.55, 0.55, 0.53, 
    0.53, 0.49, 0.46, 0.5, 0.48, 0.47, 0.48, 0.48, 0.46, 0.46, 0.48, 0.47, 
    0.46, 0.46, 0.48, 0.49, 0.49, 0.49, 0.48, 0.52, 0.55, 0.57, 0.51, 0.57, 
    0.57, 0.66, 0.47, 0.49, 0.47, 0.48, 0.48, 0.5, 0.55, 0.49, 0.5, 0.5, 
    0.49, 0.53, 0.48, 0.49, 0.48, 0.48, 0.48, 0.49, 0.49, 0.47, 0.49, 0.5, 
    0.48, 0.56, 0.55, 0.57, 0.56, 0.6, 0.5, 0.52, 0.54, 0.55, 0.6, 0.64, 
    0.62, 0.59, 0.6, 0.6, 0.57, 0.61, 0.62, 0.6, 0.64, 0.65, 0.67, 0.68, 
    0.68, 0.67, 0.66, 0.67, 0.71, 0.73, 0.74, 0.74, 0.74, 0.76, 0.74, 0.75, 
    0.71, 0.7, 0.68, 0.7, 0.71, 0.7, 0.72, 0.72, 0.7, 0.67, 0.63, 0.62, 0.58, 
    0.62, 0.67, 0.66, 0.66, 0.81, 0.91, 0.93, 0.92, 0.88, 0.86, 0.88, 1, 
    0.89, 0.82, 0.85, 0.82, 0.87, 0.92, 0.94, 0.96, 0.97, 0.96, 0.97, 0.98, 
    0.85, 0.74, 0.71, 0.71, 0.72, 0.72, 0.69, 0.64, 0.68, 0.72, 0.7, 0.68, 
    0.67, 0.74, 0.72, 0.74, 0.77, 0.74, 0.75, 0.72, 0.76, 0.73, 0.74, 0.73, 
    0.67, 0.7, 0.61, 0.67, 0.69, 0.77, 0.89, 0.87, 0.88, 0.9, 0.91, 0.92, 
    0.93, 0.94, 0.95, 0.95, 0.94, 0.95, 0.93, 0.93, 0.92, 0.93, 0.95, 0.95, 
    0.96, 0.96, 0.97, 0.98, 0.98, 0.98, 0.98, 0.98, 0.97, 0.95, 0.91, 0.87, 
    0.82, 0.82, 0.84, 0.86, 0.85, 0.88, 0.91, 0.93, 0.94, 0.95, 0.96, 0.96, 
    0.96, 0.96, 0.96, 0.91, 0.9, 0.88, 0.83, 0.77, 0.74, 0.71, 0.71, 0.69, 
    0.67, 0.65, 0.67, 0.69, 0.67, 0.67, 0.67, 0.65, 0.62, 0.63, 0.6, 0.6, 
    0.58, 0.61, 0.63, 0.61, 0.61, 0.6, 0.6, 0.61, 0.6, 0.61, 0.6, 0.62, 0.63, 
    0.65, 0.61, 0.62, 0.64, 0.63, 0.64, 0.64, 0.63, 0.7, 0.67, 0.67, 0.63, 
    0.66, 0.71, 0.65, 0.64, 0.64, 0.67, 0.7, 0.66, 0.62, 0.64, 0.59, 0.62, 
    0.62, 0.65, 0.66, 0.65, 0.59, 0.61, 0.63, 0.6, 0.59, 0.6, 0.57, 0.57, 
    0.56, 0.56, 0.55, 0.62, 0.55, 0.6, 0.6, 0.54, 0.56, 0.53, 0.6, 0.57, 
    0.58, 0.58, 0.58, 0.56, 0.57, 0.57, 0.57, 0.6, 0.53, 0.6, 0.61, 0.59, 
    0.6, 0.62, 0.62, 0.64, 0.65, 0.6, 0.6, 0.58, 0.6, 0.63, 0.6, 0.66, 0.59, 
    0.68, 0.68, 0.67, 0.61, 0.66, 0.68, 0.65, 0.65, 0.67, 0.59, 0.69, 0.63, 
    0.66, 0.6, 0.64, 0.62, 0.63, 0.63, 0.6, 0.61, 0.61, 0.59, 0.59, 0.58, 
    0.59, 0.59, 0.76, 0.84, 0.77, 0.72, 0.7, 0.83, 0.88, 0.85, 0.85, 0.82, 
    0.85, 0.83, 0.82, 0.77, 0.73, 0.72, 0.71, 0.72, 0.72, 0.75, 0.76, 0.78, 
    0.76, 0.79, 0.77, 0.8, 0.78, 0.77, 0.73, 0.74, 0.74, 0.77, 0.74, 0.71, 
    0.73, 0.72, 0.74, 0.74, 0.75, 0.75, 0.75, 0.74, 0.78, 0.88, 0.86, 0.82, 
    0.81, 0.77, 0.78, 0.81, 0.79, 0.8, 0.83, 0.81, 0.83, 0.82, 0.77, 0.79, 
    0.76, 0.8, 0.79, 0.8, 0.8, 0.83, 0.85, 0.86, 0.85, 0.8, 0.79, 0.8, 0.87, 
    0.84, 0.8, 0.85, 0.89, 0.92, 0.95, 0.93, 0.95, 0.97, 0.97, 0.97, 0.96, 
    0.98, 0.97, 0.98, 0.96, 0.89, 0.9, 0.83, 0.83, 0.83, 0.86, 0.9, 0.91, 
    0.93, 0.94, 0.83, 0.8, 0.8, 0.77, 0.72, 0.8, 0.68, 0.64, 0.7, 0.68, 0.68, 
    0.61, 0.67, 0.62, 0.62, 0.62, 0.58, 0.54, 0.52, 0.55, 0.61, 0.58, 0.6, 
    0.54, 0.55, 0.55, 0.56, 0.52, 0.56, 0.55, 0.53, 0.55, 0.57, 0.57, 0.61, 
    0.59, 0.63, 0.67, 0.63, 0.63, 0.62, 0.67, 0.68, 0.69, 0.71, 0.73, 0.74, 
    0.74, 0.73, 0.68, 0.66, 0.67, 0.66, 0.65, 0.67, 0.66, 0.67, 0.66, 0.65, 
    0.66, 0.68, 0.69, 0.7, 0.72, 0.67, 0.68, 0.67, 0.69, 0.65, 0.67, 0.71, 
    0.73, 0.77, 0.81, 0.83, 0.85, 0.88, 0.89, 0.9, 0.91, 0.92, 0.89, 0.92, 
    0.91, 0.91, 0.88, 0.87, 0.85, 0.81, 0.74, 0.79, 0.72, 0.69, 0.66, 0.66, 
    0.64, 0.66, 0.67, 0.66, 0.65, 0.67, 0.66, 0.65, 0.64, 0.64, 0.63, 0.61, 
    0.61, 0.59, 0.6, 0.64, 0.64, 0.65, 0.64, 0.67, 0.69, 0.68, 0.69, 0.7, 
    0.71, 0.72, 0.72, 0.74, 0.72, 0.72, 0.73, 0.68, 0.63, 0.63, 0.62, 0.65, 
    0.66, 0.63, 0.66, 0.66, 0.66, 0.68, 0.69, 0.71, 0.74, 0.75, 0.75, 0.75, 
    0.76, 0.76, 0.78, 0.8, 0.79, 0.77, 0.78, 0.78, 0.8, 0.8, 0.72, 0.74, 
    0.84, 0.85, 0.78, 0.82, 0.85, 0.8, 0.86, 0.87, 0.85, 0.86, 0.95, 0.95, 
    0.92, 0.88, 0.85, 0.87, 0.88, 0.87, 0.9, 0.86, 0.86, 0.84, 0.91, 0.82, 
    0.91, 0.87, 0.88, 0.87, 0.86, 0.88, 0.77, 0.83, 0.76, 0.76, 0.77, 0.75, 
    0.76, 0.81, 0.8, 0.78, 0.76, 0.62, 0.56, 0.64, 0.52, 0.55, 0.59, 0.48, 
    0.54, 0.51, 0.55, 0.57, 0.55, 0.49, 0.52, 0.53, 0.47, 0.59, 0.54, 0.5, 
    0.55, 0.54, 0.53, 0.55, 0.54, 0.56, 0.56, 0.51, 0.47, 0.5, 0.52, 0.55, 
    0.57, 0.62, 0.71, 0.75, 0.8, 0.76, 0.77, 0.81, 0.84, 0.82, 0.79, 0.71, 
    0.69, 0.72, 0.7, 0.69, 0.7, 0.68, 0.66, 0.69, 0.66, 0.68, 0.68, 0.66, 
    0.68, 0.64, 0.62, 0.61, 0.61, 0.56, 0.65, 0.64, 0.66, 0.54, 0.48, 0.47, 
    0.5, 0.59, 0.6, 0.75, 0.82, 0.82, 0.82, 0.78, 0.81, 0.83, 0.72, 0.69, 
    0.69, 0.65, 0.64, 0.66, 0.63, 0.62, 0.58, 0.56, 0.61, 0.58, 0.58, 0.57, 
    0.55, 0.57, 0.51, 0.55, 0.55, 0.58, 0.61, 0.58, 0.58, 0.59, 0.56, 0.62, 
    0.67, 0.63, 0.68, 0.74, 0.63, 0.67, 0.62, 0.7, 0.61, 0.59, 0.55, 0.53, 
    0.58, 0.57, 0.59, 0.59, 0.61, 0.63, 0.56, 0.58, 0.59, 0.61, 0.59, 0.54, 
    0.56, 0.57, 0.59, 0.62, 0.63, 0.65, 0.66, 0.66, 0.71, 0.73, 0.66, 0.63, 
    0.63, 0.58, 0.62, 0.6, 0.65, 0.62, 0.61, 0.65, 0.63, 0.67, 0.66, 0.68, 
    0.67, 0.67, 0.69, 0.71, 0.65, 0.64, 0.7, 0.64, 0.65, 0.66, 0.66, 0.66, 
    0.66, 0.66, 0.63, 0.69, 0.64, 0.64, 0.67, 0.63, 0.63, 0.64, 0.59, 0.59, 
    0.64, 0.57, 0.58, 0.62, 0.61, 0.63, 0.62, 0.69, 0.73, 0.65, 0.66, 0.64, 
    0.78, 0.72, 0.68, 0.88, 0.9, 0.91, 0.92, 0.92, 0.91, 0.9, 0.88, 0.84, 
    0.83, 0.81, 0.85, 0.75, 0.76, 0.72, 0.76, 0.79, 0.77, 0.71, 0.73, 0.65, 
    0.57, 0.56, 0.56, 0.5, 0.37, 0.63, 0.66, 0.74, 0.73, 0.64, 0.59, 0.67, 
    0.8, 0.88, 0.8, 0.72, 0.72, 0.67, 0.69, 0.75, 0.68, 0.62, 0.66, 0.63, 
    0.6, 0.53, 0.52, 0.49, 0.5, 0.55, 0.52, 0.51, 0.51, 0.49, 0.45, 0.5, 
    0.48, 0.53, 0.52, 0.54, 0.57, 0.56, 0.56, 0.58, 0.61, 0.61, 0.59, 0.59, 
    0.58, 0.62, 0.63, 0.8, 0.77, 0.73, 0.79, 0.73, 0.58, 0.55, 0.6, 0.65, 
    0.59, 0.64, 0.61, 0.56, 0.55, 0.68, 0.55, 0.58, 0.57, 0.53, 0.55, 0.53, 
    0.52, 0.52, 0.51, 0.52, 0.55, 0.57, 0.54, 0.54, 0.54, 0.52, 0.56, 0.48, 
    0.48, 0.5, 0.49, 0.49, 0.48, 0.5, 0.48, 0.5, 0.49, 0.49, 0.5, 0.48, 0.5, 
    0.51, 0.49, 0.49, 0.51, 0.5, 0.46, 0.47, 0.5, 0.48, 0.47, 0.49, 0.54, 
    0.56, 0.57, 0.6, 0.6, 0.62, 0.62, 0.63, 0.56, 0.55, 0.52, 0.54, 0.59, 
    0.58, 0.53, 0.55, 0.58, 0.58, 0.57, 0.54, 0.55, 0.56, 0.56, 0.57, 0.57, 
    0.6, 0.57, 0.57, 0.58, 0.58, 0.58, 0.58, 0.6, 0.57, 0.55, 0.54, 0.59, 
    0.63, 0.58, 0.6, 0.67, 0.68, 0.68, 0.72, 0.66, 0.72, 0.88, 0.91, 0.85, 
    0.82, 0.73, 0.67, 0.67, 0.67, 0.7, 0.75, 0.69, 0.71, 0.71, 0.74, 0.76, 
    0.81, 0.81, 0.74, 0.75, 0.81, 0.8, 0.91, 0.94, 0.95, 0.94, 0.97, 0.97, 
    0.97, 0.97, 0.98, 0.98, 0.98, 0.97, 0.92, 0.92, 0.89, 0.83, 0.74, 0.72, 
    0.71, 0.74, 0.73, 0.72, 0.71, 0.69, 0.67, 0.66, 0.65, 0.63, 0.63, 0.64, 
    0.6, 0.57, 0.59, 0.57, 0.56, 0.58, 0.61, 0.63, 0.61, 0.63, 0.61, 0.64, 
    0.64, 0.57, 0.61, 0.62, 0.59, 0.63, 0.63, 0.7, 0.62, 0.62, 0.62, 0.61, 
    0.58, 0.61, 0.6, 0.62, 0.59, 0.62, 0.63, 0.66, 0.68, 0.66, 0.64, 0.62, 
    0.64, 0.62, 0.65, 0.5, 0.55, 0.64, 0.77, 0.81, 0.8, 0.54, 0.5, 0.49, 
    0.49, 0.53, 0.51, 0.56, 0.58, 0.6, 0.59, 0.61, 0.56, 0.65, 0.64, 0.62, 
    0.62, 0.68, 0.69, 0.71, 0.71, 0.64, 0.61, 0.62, 0.54, 0.55, 0.61, 0.6, 
    0.61, 0.6, 0.56, 0.51, 0.59, 0.56, 0.52, 0.52, 0.54, 0.53, 0.53, 0.54, 
    0.51, 0.53, 0.53, 0.7, 0.71, 0.81, 0.76, 0.6, 0.57, 0.54, 0.59, 0.57, 
    0.5, 0.53, 0.57, 0.61, 0.68, 0.72, 0.73, 0.7, 0.68, 0.72, 0.75, 0.7, 
    0.64, 0.67, 0.75, 0.68, 0.69, 0.56, 0.58, 0.64, 0.7, 0.65, 0.56, 0.66, 
    0.69, 0.64, 0.57, 0.55, 0.62, 0.59, 0.63, 0.65, 0.63, 0.62, 0.62, 0.67, 
    0.67, 0.68, 0.68, 0.73, 0.71, 0.74, 0.73, 0.75, 0.72, 0.78, 0.89, 0.87, 
    0.91, 0.93, 0.95, 0.96, 0.96, 0.97, 0.95, 0.91, 0.79, 0.75, 0.76, 0.75, 
    0.8, 0.83, 0.78, 0.82, 0.86, 0.78, 0.84, 0.77, 0.75, 0.7, 0.69, 0.7, 
    0.74, 0.73, 0.73, 0.68, 0.76, 0.78, 0.74, 0.81, 0.82, 0.79, 0.76, 0.75, 
    0.82, 0.77, 0.81, 0.8, 0.79, 0.76, 0.77, 0.79, 0.69, 0.75, 0.76, 0.81, 
    0.85, 0.87, 0.93, 0.95, 0.95, 0.95, 0.96, 0.96, 0.96, 0.97, 0.97, 0.96, 
    0.97, 0.97, 0.87, 0.87, 0.89, 0.9, 0.84, 0.82, 0.79, 0.77, 0.76, 0.84, 
    0.84, 0.66, 0.56, 0.59, 0.63, 0.6, 0.56, 0.52, 0.54, 0.58, 0.55, 0.57, 
    0.54, 0.47, 0.48, 0.48, 0.46, 0.5, 0.57, 0.62, 0.65, 0.7, 0.64, 0.64, 
    0.58, 0.49, 0.55, 0.52, 0.49, 0.53, 0.53, 0.52, 0.51, 0.57, 0.55, 0.58, 
    0.62, 0.57, 0.64, 0.57, 0.58, 0.64, 0.57, 0.61, 0.6, 0.6, 0.64, 0.62, 
    0.64, 0.63, 0.65, 0.64, 0.65, 0.66, 0.7, 0.74, 0.78, 0.78, 0.78, 0.83, 
    0.88, 0.88, 0.89, 0.88, 0.86, 0.86, 0.88, 0.88, 0.91, 0.93, 0.91, 0.92, 
    0.96, 0.96, 0.87, 0.77, 0.78, 0.77, 0.76, 0.8, 0.85, 0.86, 0.8, 0.81, 
    0.79, 0.77, 0.82, 0.85, 0.83, 0.82, 0.76, 0.8, 0.79, 0.76, 0.74, 0.73, 
    0.75, 0.72, 0.75, 0.75, 0.76, 0.77, 0.77, 0.73, 0.76, 0.77, 0.78, 0.78, 
    0.84, 0.89, 0.89, 0.8, 0.81, 0.81, 0.78, 0.81, 0.76, 0.78, 0.86, 0.89, 
    0.93, 0.9, 0.91, 0.87, 0.82, 0.84, 0.87, 0.87, 0.87, 0.82, 0.82, 0.83, 
    0.8, 0.85, 0.82, 0.85, 0.84, 0.82, 0.82, 0.85, 0.87, 0.9, 0.9, 0.92, 
    0.93, 0.91, 0.92, 0.89, 0.82, 0.85, 0.77, 0.56, 0.63, 0.76, 0.82, 0.79, 
    0.68, 0.61, 0.73, 0.84, 0.74, 0.74, 0.75, 0.73, 0.76, 0.77, 0.78, 0.74, 
    0.63, 0.6, 0.62, 0.65, 0.54, 0.51, 0.51, 0.51, 0.51, 0.49, 0.52, 0.51, 
    0.49, 0.49, 0.54, 0.54, 0.47, 0.49, 0.47, 0.54, 0.56, 0.56, 0.58, 0.6, 
    0.56, 0.59, 0.6, 0.61, 0.62, 0.6, 0.63, 0.61, 0.63, 0.64, 0.62, 0.58, 
    0.55, 0.56, 0.54, 0.53, 0.52, 0.56, 0.55, 0.76, 0.81, 0.83, 0.84, 0.84, 
    0.84, 0.67, 0.68, 0.65, 0.64, 0.68, 0.66, 0.65, 0.64, 0.66, 0.65, 0.59, 
    0.61, 0.61, 0.65, 0.64, 0.6, 0.58, 0.63, 0.67, 0.67, 0.64, 0.67, 0.7, 
    0.7, 0.7, 0.67, 0.66, 0.65, 0.63, 0.6, 0.6, 0.58, 0.58, 0.58, 0.59, 0.63, 
    0.6, 0.55, 0.52, 0.52, 0.51, 0.51, 0.52, 0.52, 0.5, 0.5, 0.47, 0.47, 
    0.47, 0.48, 0.48, 0.48, 0.54, 0.52, 0.55, 0.56, 0.57, 0.57, 0.56, 0.56, 
    0.54, 0.51, 0.53, 0.53, 0.52, 0.52, 0.52, 0.53, 0.55, 0.56, 0.55, 0.55, 
    0.56, 0.75, 0.76, 0.79, 0.77, 0.66, 0.62, 0.56, 0.61, 0.41, 0.39, 0.35, 
    0.4, 0.39, 0.41, 0.42, 0.45, 0.49, 0.61, 0.72, 0.75, 0.72, 0.68, 0.63, 
    0.61, 0.62, 0.66, 0.72, 0.75, 0.74, 0.49, 0.59, 0.7, 0.62, 0.58, 0.55, 
    0.54, 0.5, 0.56, 0.57, 0.52, 0.49, 0.5, 0.59, 0.52, 0.55, 0.56, 0.51, 
    0.57, 0.58, 0.56, 0.62, 0.59, 0.53, 0.49, 0.5, 0.5, 0.49, 0.48, 0.47, 
    0.51, 0.5, 0.53, 0.56, 0.54, 0.63, 0.59, 0.62, 0.58, 0.55, 0.5, 0.51, 
    0.56, 0.52, 0.48, 0.47, 0.47, 0.47, 0.47, 0.44, 0.52, 0.56, 0.53, 0.55, 
    0.56, 0.6, 0.6, 0.65, 0.6, 0.6, 0.56, 0.57, 0.55, 0.61, 0.66, 0.63, 0.61, 
    0.53, 0.53, 0.52, 0.54, 0.53, 0.48, 0.51, 0.54, 0.51, 0.52, 0.46, 0.53, 
    0.54, 0.58, 0.52, 0.51, 0.49, 0.5, 0.5, 0.5, 0.5, 0.5, 0.53, 0.5, 0.5, 
    0.51, 0.53, 0.49, 0.5, 0.47, 0.49, 0.52, 0.53, 0.53, 0.6, 0.56, 0.59, 
    0.59, 0.63, 0.58, 0.62, 0.6, 0.61, 0.6, 0.54, 0.57, 0.55, 0.59, 0.67, 
    0.7, 0.67, 0.69, 0.66, 0.78, 0.86, 0.86, 0.86, 0.83, 0.8, 0.76, 0.72, 
    0.72, 0.74, 0.7, 0.68, 0.69, 0.67, 0.72, 0.73, 0.73, 0.72, 0.71, 0.65, 
    0.72, 0.73, 0.67, 0.71, 0.73, 0.77, 0.75, 0.77, 0.76, 0.76, 0.81, 0.78, 
    0.75, 0.88, 0.94, 0.95, 0.94, 0.94, 0.94, 0.95, 0.95, 0.95, 0.96, 0.97, 
    0.96, 0.96, 0.96, 0.94, 0.95, 0.92, 0.95, 0.92, 0.94, 0.91, 0.92, 0.84, 
    0.83, 0.82, 0.8, 0.75, 0.67, 0.64, 0.65, 0.65, 0.71, 0.67, 0.71, 0.66, 
    0.68, 0.68, 0.7, 0.72, 0.68, 0.64, 0.63, 0.68, 0.65, 0.65, 0.68, 0.69, 
    0.67, 0.65, 0.67, 0.67, 0.66, 0.65, 0.64, 0.64, 0.64, 0.64, 0.59, 0.61, 
    0.61, 0.6, 0.56, 0.58, 0.58, 0.57, 0.56, 0.55, 0.58, 0.53, 0.52, 0.51, 
    0.54, 0.54, 0.49, 0.53, 0.6, 0.62, 0.65, 0.67, 0.63, 0.65, 0.63, 0.58, 
    0.59, 0.58, 0.56, 0.55, 0.57, 0.57, 0.6, 0.62, 0.62, 0.63, 0.64, 0.6, 
    0.63, 0.62, 0.59, 0.61, 0.61, 0.63, 0.71, 0.67, 0.69, 0.74, 0.75, 0.78, 
    0.85, 0.89, 0.88, 0.87, 0.89, 0.9, 0.86, 0.85, 0.8, 0.67, 0.72, 0.67, 
    0.64, 0.63, 0.6, 0.61, 0.65, 0.67, 0.68, 0.7, 0.7, 0.73, 0.76, 0.73, 
    0.75, 0.72, 0.75, 0.62, 0.68, 0.7, 0.74, 0.65, 0.68, 0.66, 0.67, 0.59, 
    0.64, 0.67, 0.74, 0.68, 0.74, 0.67, 0.67, 0.64, 0.59, 0.59, 0.57, 0.52, 
    0.5, 0.45, 0.46, 0.46, 0.43, 0.44, 0.43, 0.41, 0.45, 0.42, 0.42, 0.41, 
    0.42, 0.42, 0.42, 0.41, 0.41, 0.41, 0.42, 0.4, 0.39, 0.4, 0.4, 0.45, 
    0.39, 0.39, 0.42, 0.45, 0.48, 0.5, 0.41, 0.41, 0.38, 0.41, 0.47, 0.46, 
    0.5, 0.47, 0.5, 0.52, 0.5, 0.52, 0.51, 0.5, 0.46, 0.4, 0.38, 0.39, 0.41, 
    0.45, 0.45, 0.49, 0.46, 0.47, 0.46, 0.5, 0.47, 0.49, 0.48, 0.46, 0.49, 
    0.46, 0.46, 0.43, 0.42, 0.43, 0.47, 0.51, 0.5, 0.5, 0.48, 0.45, 0.58, 
    0.57, 0.55, 0.58, 0.55, 0.56, 0.55, 0.56, 0.54, 0.57, 0.56, 0.56, 0.59, 
    0.57, 0.61, 0.6, 0.59, 0.65, 0.59, 0.62, 0.61, 0.63, 0.64, 0.75, 0.61, 
    0.62, 0.69, 0.65, 0.63, 0.68, 0.67, 0.68, 0.63, 0.66, 0.65, 0.61, 0.65, 
    0.65, 0.63, 0.64, 0.65, 0.67, 0.63, 0.68, 0.65, 0.64, 0.66, 0.64, 0.62, 
    0.64, 0.66, 0.64, 0.67, 0.67, 0.67, 0.62, 0.57, 0.67, 0.66, 0.64, 0.79, 
    0.84, 0.84, 0.83, 0.81, 0.8, 0.76, 0.79, 0.74, 0.69, 0.67, 0.58, 0.58, 
    0.6, 0.55, 0.58, 0.52, 0.54, 0.56, 0.64, 0.65, 0.63, 0.65, 0.66, 0.66, 
    0.63, 0.59, 0.54, 0.55, 0.55, 0.56, 0.59, 0.65, 0.65, 0.58, 0.59, 0.6, 
    0.49, 0.45, 0.44, 0.54, 0.52, 0.53, 0.48, 0.44, 0.45, 0.44, 0.43, 0.44, 
    0.45, 0.44, 0.46, 0.47, 0.47, 0.5, 0.5, 0.5, 0.49, 0.53, 0.5, 0.52, 0.55, 
    0.53, 0.52, 0.5, 0.53, 0.51, 0.52, 0.57, 0.59, 0.59, 0.59, 0.6, 0.6, 
    0.58, 0.62, 0.61, 0.58, 0.65, 0.64, 0.6, 0.6, 0.6, 0.6, 0.62, 0.58, 0.61, 
    0.61, 0.61, 0.62, 0.61, 0.62, 0.6, 0.62, 0.61, 0.6, 0.59, 0.62, 0.61, 
    0.62, 0.63, 0.66, 0.66, 0.63, 0.67, 0.69, 0.69, 0.68, 0.72, 0.68, 0.68, 
    0.68, 0.66, 0.67, 0.67, 0.64, 0.65, 0.68, 0.67, 0.7, 0.67, 0.67, 0.66, 
    0.67, 0.66, 0.66, 0.65, 0.59, 0.57, 0.64, 0.57, 0.53, 0.57, 0.51, 0.58, 
    0.5, 0.45, 0.49, 0.52, 0.49, 0.5, 0.53, 0.57, 0.62, 0.58, 0.62, 0.68, 
    0.67, 0.59, 0.7, 0.58, 0.68, 0.6, 0.58, 0.61, 0.64, 0.64, 0.61, 0.63, 
    0.58, 0.55, 0.54, 0.54, 0.54, 0.59, 0.58, 0.59, 0.59, 0.57, 0.55, 0.6, 
    0.59, 0.6, 0.6, 0.68, 0.6, 0.65, 0.69, 0.68, 0.69, 0.64, 0.71, 0.62, 
    0.69, 0.65, 0.64, 0.7, 0.7, 0.68, 0.66, 0.73, 0.73, 0.75, 0.73, 0.7, 
    0.74, 0.73, 0.71, 0.72, 0.77, 0.73, 0.75, 0.75, 0.74, 0.74, 0.74, 0.76, 
    0.74, 0.78, 0.77, 0.76, 0.78, 0.81, 0.79, 0.82, 0.81, 0.8, 0.8, 0.78, 
    0.69, 0.7, 0.75, 0.83, 0.88, 0.84, 0.8, 0.83, 0.83, 0.8, 0.8, 0.74, 0.82, 
    0.77, 0.74, 0.81, 0.73, 0.74, 0.7, 0.64, 0.76, 0.65, 0.71, 0.73, 0.7, 
    0.73, 0.71, 0.68, 0.73, 0.75, 0.74, 0.72, 0.73, 0.7, 0.72, 0.7, 0.63, 
    0.7, 0.74, 0.71, 0.7, 0.72, 0.75, 0.74, 0.72, 0.75, 0.7, 0.71, 0.62, 
    0.68, 0.64, 0.64, 0.59, 0.58, 0.6, 0.63, 0.62, 0.66, 0.72, 0.65, 0.65, 
    0.7, 0.68, 0.69, 0.68, 0.63, 0.61, 0.62, 0.64, 0.62, 0.69, 0.66, 0.6, 
    0.56, 0.6, 0.62, 0.63, 0.61, 0.59, 0.55, 0.58, 0.61, 0.66, 0.67, 0.61, 
    0.61, 0.62, 0.64, 0.65, 0.69, 0.73, 0.72, 0.74, 0.73, 0.68, 0.69, 0.69, 
    0.67, 0.64, 0.64, 0.58, 0.6, 0.64, 0.67, 0.73, 0.68, 0.63, 0.64, 0.65, 
    0.65, 0.67, 0.67, 0.65, 0.68, 0.79, 0.76, 0.69, 0.7, 0.73, 0.72, 0.74, 
    0.74, 0.77, 0.71, 0.67, 0.67, 0.7, 0.67, 0.66, 0.65, 0.66, 0.69, 0.75, 
    0.72, 0.67, 0.64, 0.67, 0.64, 0.69, 0.67, 0.69, 0.67, 0.69, 0.75, 0.66, 
    0.7, 0.68, 0.66, 0.6, 0.61, 0.62, 0.61, 0.6, 0.6, 0.62, 0.63, 0.67, 0.65, 
    0.67, 0.73, 0.75, 0.75, 0.69, 0.69, 0.7, 0.69, 0.71, 0.72, 0.71, 0.68, 
    0.7, 0.68, 0.73, 0.69, 0.7, 0.72, 0.73, 0.65, 0.64, 0.65, 0.59, 0.59, 
    0.57, 0.57, 0.58, 0.58, 0.55, 0.6, 0.63, 0.61, 0.62, 0.64, 0.66, 0.63, 
    0.61, 0.62, 0.63, 0.67, 0.65, 0.64, 0.62, 0.66, 0.64, 0.64, 0.63, 0.65, 
    0.65, 0.63, 0.64, 0.62, 0.64, 0.63, 0.63, 0.65, 0.66, 0.65, 0.68, 0.74, 
    0.72, 0.72, 0.71, 0.69, 0.66, 0.67, 0.66, 0.69, 0.62, 0.65, 0.67, 0.69, 
    0.67, 0.72, 0.68, 0.66, 0.65, 0.69, 0.65, 0.7, 0.71, 0.66, 0.68, 0.68, 
    0.71, 0.71, 0.7, 0.74, 0.72, 0.72, 0.72, 0.72, 0.73, 0.78, 0.75, 0.8, 
    0.76, 0.77, 0.75, 0.76, 0.76, 0.77, 0.74, 0.75, 0.77, 0.71, 0.79, 0.73, 
    0.75, 0.76, 0.75, 0.72, 0.72, 0.66, 0.71, 0.68, 0.67, 0.64, 0.73, 0.64, 
    0.66, 0.68, 0.72, 0.68, 0.67, 0.66, 0.64, 0.62, 0.63, 0.62, 0.67, 0.63, 
    0.63, 0.68, 0.56, 0.56, 0.54, 0.58, 0.57, 0.55, 0.56, 0.55, 0.53, 0.52, 
    0.5, 0.51, 0.52, 0.49, 0.5, 0.51, 0.52, 0.5, 0.52, 0.5, 0.51, 0.5, 0.46, 
    0.47, 0.48, 0.48, 0.47, 0.45, 0.48, 0.47, 0.51, 0.47, 0.48, 0.5, 0.46, 
    0.58, 0.5, 0.51, 0.57, 0.45, 0.45, 0.43, 0.45, 0.47, 0.48, 0.54, 0.48, 
    0.54, 0.54, 0.54, 0.51, 0.52, 0.49, 0.45, 0.44, 0.46, 0.47, 0.48, 0.55, 
    0.57, 0.56, 0.56, 0.55, 0.57, 0.57, 0.51, 0.56, 0.59, 0.57, 0.55, 0.55, 
    0.54, 0.54, 0.55, 0.58, 0.54, 0.54, 0.52, 0.46, 0.48, 0.51, 0.52, 0.54, 
    0.55, 0.58, 0.56, 0.59, 0.6, 0.59, 0.6, 0.58, 0.6, 0.63, 0.61, 0.65, 
    0.61, 0.55, 0.54, 0.5, 0.48, 0.47, 0.52, 0.5, 0.55, 0.54, 0.55, 0.58, 
    0.64, 0.62, 0.61, 0.6, 0.61, 0.64, 0.7, 0.69, 0.73, 0.77, 0.77, 0.68, 
    0.63, 0.68, 0.63, 0.63, 0.62, 0.62, 0.6, 0.63, 0.62, 0.63, 0.62, 0.64, 
    0.63, 0.63, 0.61, 0.63, 0.63, 0.65, 0.64, 0.67, 0.67, 0.72, 0.71, 0.7, 
    0.68, 0.74, 0.71, 0.71, 0.72, 0.73, 0.73, 0.76, 0.73, 0.74, 0.7, 0.71, 
    0.66, 0.69, 0.62, 0.64, 0.67, 0.62, 0.62, 0.59, 0.56, 0.62, 0.59, 0.63, 
    0.59, 0.63, 0.7, 0.68, 0.64, 0.68, 0.66, 0.68, 0.68, 0.71, 0.66, 0.73, 
    0.68, 0.7, 0.69, 0.74, 0.66, 0.66, 0.72, 0.66, 0.69, 0.73, 0.62, 0.7, 
    0.66, 0.68, 0.69, 0.66, 0.68, 0.69, 0.68, 0.61, 0.61, 0.62, 0.66, 0.64, 
    0.62, 0.65, 0.59, 0.67, 0.63, 0.61, 0.69, 0.7, 0.6, 0.64, 0.6, 0.63, 
    0.57, 0.56, 0.59, 0.59, 0.59, 0.6, 0.61, 0.58, 0.55, 0.54, 0.54, 0.53, 
    0.51, 0.53, 0.52, 0.48, 0.47, 0.43, 0.45, 0.43, 0.45, 0.44, 0.43, 0.33, 
    0.4, 0.4, 0.47, 0.47, 0.48, 0.49, 0.48, 0.51, 0.51, 0.51, 0.55, 0.56, 
    0.55, 0.53, 0.52, 0.52, 0.48, 0.47, 0.5, 0.49, 0.48, 0.47, 0.48, 0.48, 
    0.49, 0.45, 0.48, 0.48, 0.52, 0.47, 0.48, 0.46, 0.46, 0.45, 0.52, 0.51, 
    0.53, 0.52, 0.56, 0.55, 0.57, 0.57, 0.55, 0.56, 0.54, 0.52, 0.53, 0.53, 
    0.52, 0.52, 0.52, 0.57, 0.57, 0.62, 0.62, 0.61, 0.6, 0.62, 0.6, 0.61, 
    0.58, 0.58, 0.6, 0.61, 0.56, 0.57, 0.61, 0.61, 0.6, 0.58, 0.57, 0.55, 
    0.59, 0.59, 0.56, 0.63, 0.61, 0.62, 0.64, 0.64, 0.62, 0.59, 0.59, 0.6, 
    0.63, 0.61, 0.61, 0.6, 0.6, 0.61, 0.6, 0.63, 0.64, 0.66, 0.72, 0.73, 
    0.73, 0.76, 0.8, 0.77, 0.77, 0.81, 0.78, 0.78, 0.74, 0.68, 0.68, 0.71, 
    0.72, 0.71, 0.71, 0.74, 0.72, 0.73, 0.77, 0.8, 0.84, 0.86, 0.87, 0.89, 
    0.87, 0.76, 0.89, 0.87, 0.84, 0.86, 0.82, 0.84, 0.85, 0.82, 0.87, 0.8, 
    0.79, 0.79, 0.89, 0.89, 0.84, 0.86, 0.9, 0.95, 0.95, 0.96, 0.97, 0.98, 
    0.98, 0.97, 0.96, 0.97, 0.76, 0.73, 0.73, 0.78, 0.76, 0.73, 0.69, 0.67, 
    0.64, 0.62, 0.62, 0.69, 0.72, 0.67, 0.75, 0.76, 0.77, 0.78, 0.83, 0.78, 
    0.73, 0.79, 0.74, 0.79, 0.75, 0.76, 0.77, 0.76, 0.76, 0.76, 0.62, 0.58, 
    0.59, 0.59, 0.6, 0.58, 0.57, 0.57, 0.62, 0.67, 0.73, 0.67, 0.63, 0.61, 
    0.59, 0.54, 0.43, 0.44, 0.44, 0.42, 0.44, 0.43, 0.47, 0.46, 0.49, 0.46, 
    0.49, 0.54, 0.57, 0.54, 0.57, 0.55, 0.57, 0.6, 0.63, 0.59, 0.56, 0.55, 
    0.55, 0.56, 0.58, 0.63, 0.59, 0.62, 0.59, 0.59, 0.66, 0.61, 0.59, 0.6, 
    0.55, 0.63, 0.6, 0.6, 0.55, 0.58, 0.54, 0.62, 0.61, 0.61, 0.63, 0.69, 
    0.68, 0.74, 0.77, 0.76, 0.79, 0.81, 0.81, 0.81, 0.8, 0.76, 0.75, 0.68, 
    0.71, 0.71, 0.65, 0.59, 0.6, 0.61, 0.58, 0.59, 0.6, 0.62, 0.62, 0.57, 
    0.56, 0.55, 0.56, 0.51, 0.49, 0.5, 0.54, 0.48, 0.48, 0.49, 0.42, 0.43, 
    0.44, 0.5, 0.46, 0.46, 0.48, 0.47, 0.46, 0.45, 0.52, 0.5, 0.52, 0.53, 
    0.55, 0.54, 0.5, 0.5, 0.52, 0.55, 0.56, 0.58, 0.61, 0.58, 0.59, 0.6, 
    0.63, 0.62, 0.58, 0.61, 0.6, 0.58, 0.58, 0.58, 0.54, 0.61, 0.62, 0.61, 
    0.64, 0.63, 0.66, 0.69, 0.69, 0.66, 0.67, 0.67, 0.6, 0.59, 0.55, 0.55, 
    0.58, 0.57, 0.53, 0.57, 0.55, 0.56, 0.62, 0.6, 0.57, 0.62, 0.61, 0.69, 
    0.66, 0.63, 0.62, 0.63, 0.62, 0.65, 0.54, 0.53, 0.52, 0.55, 0.49, 0.54, 
    0.5, 0.53, 0.45, 0.47, 0.47, 0.44, 0.45, 0.47, 0.44, 0.47, 0.5, 0.5, 
    0.51, 0.51, 0.52, 0.52, 0.52, 0.47, 0.52, 0.52, 0.49, 0.55, 0.52, 0.51, 
    0.5, 0.56, 0.55, 0.49, 0.49, 0.5, 0.49, 0.54, 0.57, 0.57, 0.57, 0.58, 
    0.65, 0.62, 0.64, 0.61, 0.62, 0.61, 0.59, 0.6, 0.62, 0.61, 0.59, 0.55, 
    0.57, 0.58, 0.55, 0.54, 0.53, 0.56, 0.57, 0.6, 0.6, 0.56, 0.56, 0.55, 
    0.48, 0.51, 0.53, 0.55, 0.57, 0.56, 0.58, 0.55, 0.53, 0.53, 0.53, 0.59, 
    0.62, 0.56, 0.56, 0.54, 0.47, 0.51, 0.45, 0.42, 0.44, 0.46, 0.39, 0.39, 
    0.45, 0.48, 0.43, 0.41, 0.38, 0.38, 0.44, 0.37, 0.41, 0.44, 0.49, 0.46, 
    0.48, 0.52, 0.4, 0.48, 0.44, 0.48, 0.49, 0.48, 0.49, 0.46, 0.45, 0.44, 
    0.44, 0.46, 0.43, 0.43, 0.45, 0.45, 0.48, 0.5, 0.49, 0.48, 0.52, 0.49, 
    0.52, 0.51, 0.49, 0.56, 0.59, 0.6, 0.58, 0.6, 0.58, 0.65, 0.58, 0.54, 
    0.52, 0.54, 0.59, 0.55, 0.52, 0.54, 0.55, 0.54, 0.53, 0.54, 0.48, 0.59, 
    0.54, 0.49, 0.62, 0.56, 0.58, 0.6, 0.53, 0.62, 0.61, 0.54, 0.61, 0.54, 
    0.49, 0.64, 0.61, 0.69, 0.77, 0.73, 0.78, 0.79, 0.75, 0.72, 0.73, 0.74, 
    0.67, 0.77, 0.69, 0.66, 0.63, 0.69, 0.72, 0.75, 0.74, 0.69, 0.68, 0.69, 
    0.71, 0.73, 0.72, 0.7, 0.67, 0.71, 0.67, 0.72, 0.63, 0.66, 0.64, 0.69, 
    0.62, 0.66, 0.61, 0.55, 0.59, 0.6, 0.63, 0.59, 0.55, 0.6, 0.58, 0.57, 
    0.58, 0.59, 0.51, 0.58, 0.59, 0.61, 0.53, 0.6, 0.6, 0.58, 0.57, 0.7, 
    0.57, 0.64, 0.55, 0.63, 0.57, 0.62, 0.64, 0.65, 0.65, 0.61, 0.6, 0.61, 
    0.73, 0.78, 0.77, 0.76, 0.77, 0.79, 0.79, 0.75, 0.8, 0.77, 0.73, 0.74, 
    0.73, 0.72, 0.72, 0.7, 0.67, 0.69, 0.67, 0.66, 0.7, 0.73, 0.7, 0.67, 
    0.73, 0.7, 0.67, 0.7, 0.61, 0.74, 0.73, 0.72, 0.67, 0.71, 0.69, 0.68, 
    0.68, 0.62, 0.62, 0.58, 0.54, 0.61, 0.64, 0.64, 0.65, 0.65, 0.65, 0.65, 
    0.65, 0.67, 0.63, 0.7, 0.62, 0.69, 0.66, 0.66, 0.66, 0.62, 0.63, 0.62, 
    0.75, 0.76, 0.77, 0.78, 0.78, 0.77, 0.78, 0.79, 0.72, 0.69, 0.64, 0.62, 
    0.6, 0.59, 0.58, 0.58, 0.6, 0.59, 0.59, 0.59, 0.6, 0.6, 0.63, 0.63, 0.58, 
    0.53, 0.52, 0.53, 0.48, 0.5, 0.56, 0.56, 0.58, 0.63, 0.52, 0.62, 0.56, 
    0.67, 0.57, 0.6, 0.65, 0.59, 0.59, 0.54, 0.65, 0.61, 0.57, 0.5, 0.55, 
    0.49, 0.47, 0.55, 0.57, 0.52, 0.59, 0.63, 0.64, 0.61, 0.58, 0.55, 0.64, 
    0.7, 0.61, 0.57, 0.66, 0.68, 0.84, 0.82, 0.81, 0.75, 0.85, 0.82, 0.77, 
    0.76, 0.6, 0.61, 0.66, 0.67, 0.83, 0.93, 0.89, 0.84, 0.79, 0.84, 0.8, 
    0.8, 0.79, 0.66, 0.66, 0.69, 0.69, 0.68, 0.69, 0.65, 0.6, 0.59, 0.57, 
    0.57, 0.58, 0.58, 0.6, 0.59, 0.62, 0.63, 0.67, 0.67, 0.69, 0.71, 0.71, 
    0.69, 0.69, 0.64, 0.67, 0.7, 0.7, 0.81, 0.76, 0.7, 0.78, 0.69, 0.67, 
    0.64, 0.67, 0.63, 0.7, 0.69, 0.65, 0.77, 0.88, 0.84, 0.8, 0.78, 0.75, 
    0.73, 0.74, 0.71, 0.71, 0.69, 0.75, 0.75, 0.76, 0.83, 0.77, 0.77, 0.81, 
    0.72, 0.69, 0.71, 0.75, 0.78, 0.76, 0.74, 0.76, 0.75, 0.73, 0.73, 0.78, 
    0.79, 0.86, 0.85, 0.87, 0.81, 0.83, 0.77, 0.78, 0.66, 0.73, 0.64, 0.68, 
    0.65, 0.68, 0.67, 0.77, 0.84, 0.83, 0.75, 0.72, 0.68, 0.71, 0.79, 0.81, 
    0.75, 0.7, 0.78, 0.79, 0.82, 0.81, 0.79, 0.77, 0.77, 0.79, 0.77, 0.77, 
    0.77, 0.75, 0.74, 0.66, 0.54, 0.57, 0.58, 0.57, 0.58, 0.56, 0.64, 0.65, 
    0.71, 0.75, 0.83, 0.76, 0.74, 0.73, 0.67, 0.65, 0.67, 0.57, 0.65, 0.58, 
    0.59, 0.56, 0.51, 0.53, 0.55, 0.56, 0.58, 0.61, 0.61, 0.62, 0.64, 0.64, 
    0.64, 0.68, 0.68, 0.69, 0.74, 0.83, 0.86, 0.78, 0.62, 0.58, 0.58, 0.56, 
    0.53, 0.52, 0.54, 0.5, 0.51, 0.53, 0.58, 0.53, 0.54, 0.57, 0.57, 0.55, 
    0.56, 0.58, 0.59, 0.6, 0.6, 0.64, 0.67, 0.71, 0.69, 0.65, 0.65, 0.66, 
    0.67, 0.61, 0.61, 0.6, 0.64, 0.61, 0.67, 0.69, 0.7, 0.72, 0.77, 0.76, 
    0.8, 0.82, 0.84, 0.84, 0.86, 0.91, 0.86, 0.79, 0.77, 0.74, 0.7, 0.68, 
    0.67, 0.64, 0.63, 0.58, 0.53, 0.48, 0.48, 0.5, 0.5, 0.54, 0.59, 0.59, 
    0.61, 0.62, 0.66, 0.66, 0.64, 0.62, 0.6, 0.59, 0.6, 0.6, 0.63, 0.65, 
    0.62, 0.57, 0.57, 0.55, 0.55, 0.57, 0.58, 0.57, 0.65, 0.6, 0.57, 0.63, 
    0.55, 0.54, 0.55, 0.51, 0.51, 0.49, 0.58, 0.63, 0.6, 0.56, 0.57, 0.58, 
    0.58, 0.56, 0.53, 0.54, 0.53, 0.53, 0.5, 0.52, 0.56, 0.58, 0.53, 0.57, 
    0.57, 0.57, 0.59, 0.61, 0.6, 0.63, 0.63, 0.58, 0.54, 0.49, 0.5, 0.48, 
    0.47, 0.47, 0.45, 0.51, 0.61, 0.58, 0.54, 0.47, 0.47, 0.43, 0.39, 0.44, 
    0.46, 0.54, 0.59, 0.59, 0.57, 0.54, 0.55, 0.48, 0.54, 0.57, 0.55, 0.49, 
    0.52, 0.51, 0.51, 0.47, 0.46, 0.47, 0.48, 0.48, 0.46, 0.47, 0.48, 0.52, 
    0.5, 0.52, 0.52, 0.53, 0.56, 0.57, 0.58, 0.57, 0.59, 0.59, 0.59, 0.57, 
    0.58, 0.56, 0.54, 0.59, 0.6, 0.56, 0.54, 0.54, 0.57, 0.57, 0.58, 0.54, 
    0.55, 0.58, 0.6, 0.55, 0.56, 0.63, 0.58, 0.66, 0.63, 0.63, 0.62, 0.62, 
    0.59, 0.58, 0.56, 0.56, 0.56, 0.56, 0.56, 0.54, 0.6, 0.62, 0.67, 0.66, 
    0.65, 0.66, 0.68, 0.68, 0.69, 0.7, 0.69, 0.69, 0.66, 0.69, 0.67, 0.67, 
    0.62, 0.64, 0.6, 0.62, 0.65, 0.59, 0.62, 0.64, 0.65, 0.69, 0.7, 0.72, 
    0.74, 0.73, 0.75, 0.76, 0.72, 0.72, 0.74, 0.72, 0.78, 0.75, 0.68, 0.67, 
    0.69, 0.68, 0.66, 0.7, 0.64, 0.66, 0.7, 0.71, 0.73, 0.75, 0.8, 0.87, 
    0.89, 0.9, 0.94, 0.94, 0.93, 0.9, 0.84, 0.8, 0.78, 0.86, 0.81, 0.76, 
    0.69, 0.7, 0.61, 0.63, 0.6, 0.57, 0.59, 0.55, 0.54, 0.65, 0.7, 0.7, 0.68, 
    0.7, 0.71, 0.77, 0.73, 0.74, 0.66, 0.71, 0.73, 0.73, 0.69, 0.65, 0.61, 
    0.56, 0.55, 0.57, 0.7, 0.64, 0.69, 0.63, 0.54, 0.51, 0.54, 0.51, 0.63, 
    0.56, 0.53, 0.56, 0.55, 0.52, 0.53, 0.58, 0.59, 0.58, 0.58, 0.6, 0.59, 
    0.6, 0.59, 0.58, 0.6, 0.53, 0.56, 0.56, 0.62, 0.66, 0.68, 0.73, 0.75, 
    0.74, 0.7, 0.7, 0.76, 0.72, 0.77, 0.68, 0.68, 0.69, 0.62, 0.64, 0.54, 
    0.59, 0.62, 0.6, 0.58, 0.55, 0.54, 0.57, 0.63, 0.64, 0.65, 0.68, 0.69, 
    0.73, 0.69, 0.71, 0.8, 0.81, 0.84, 0.82, 0.84, 0.84, 0.83, 0.82, 0.77, 
    0.83, 0.79, 0.83, 0.82, 0.81, 0.83, 0.83, 0.86, 0.85, 0.83, 0.85, 0.88, 
    0.88, 0.86, 0.87, 0.87, 0.86, 0.89, 0.9, 0.9, 0.91, 0.9, 0.9, 0.9, 0.88, 
    0.9, 0.88, 0.9, 0.86, 0.83, 0.82, 0.87, 0.92, 0.88, 0.78, 0.75, 0.73, 
    0.74, 0.71, 0.7, 0.71, 0.72, 0.71, 0.71, 0.69, 0.7, 0.75, 0.62, 0.61, 
    0.61, 0.55, 0.55, 0.57, 0.65, 0.71, 0.7, 0.68, 0.72, 0.74, 0.74, 0.75, 
    0.79, 0.79, 0.81, 0.79, 0.81, 0.81, 0.79, 0.79, 0.79, 0.8, 0.81, 0.8, 
    0.76, 0.75, 0.82, 0.79, 0.81, 0.84, 0.83, 0.85, 0.89, 0.91, 0.92, 0.93, 
    0.92, 0.94, 0.93, 0.95, 0.94, 0.93, 0.92, 0.87, 0.88, 0.88, 0.81, 0.84, 
    0.85, 0.8, 0.83, 0.87, 0.83, 0.83, 0.78, 0.71, 0.8, 0.88, 0.86, 0.83, 
    0.82, 0.79, 0.81, 0.79, 0.84, 0.81, 0.8, 0.79, 0.77, 0.81, 0.88, 0.91, 
    0.9, 0.89, 0.87, 0.82, 0.85, 0.85, 0.75, 0.73, 0.74, 0.72, 0.74, 0.73, 
    0.74, 0.74, 0.69, 0.67, 0.69, 0.69, 0.72, 0.68, 0.67, 0.68, 0.71, 0.71, 
    0.74, 0.74, 0.76, 0.79, 0.84, 0.88, 0.86, 0.85, 0.9, 0.92, 0.93, 0.96, 
    0.84, 0.81, 0.78, 0.82, 0.84, 0.91, 0.86, 0.84, 0.8, 0.79, 0.8, 0.83, 
    0.83, 0.82, 0.82, 0.83, 0.87, 0.84, 0.86, 0.84, 0.85, 0.88, 0.89, 0.88, 
    0.9, 0.88, 0.93, 0.94, 0.92, 0.85, 0.8, 0.84, 0.8, 0.79, 0.77, 0.79, 
    0.74, 0.77, 0.82, 0.89, 0.89, 0.84, 0.91, 0.92, 0.96, 0.97, 0.98, 1, 
    0.89, 0.86, 0.87, 0.89, 0.9, 0.89, 0.87, 0.88, 0.85, 0.86, 0.9, 0.88, 
    0.88, 0.87, 0.88, 0.88, 0.88, 0.89, 0.89, 0.93, 0.9, 0.83, 0.85, 0.76, 
    0.77, 0.89, 0.81, 0.78, 0.85, 0.87, 0.89, 0.88, 0.89, 0.9, 0.86, 0.82, 
    0.84, 0.87, 0.85, 0.87, 0.92, 0.92, 0.94, 0.95, 0.96, 0.97, 0.98, 0.96, 
    0.97, 0.97, 0.93, 0.84, 0.75, 0.72, 0.71, 0.68, 0.69, 0.67, 0.68, 0.69, 
    0.62, 0.68, 0.71, 0.73, 0.72, 0.76, 0.75, 0.85, 0.87, 0.85, 0.82, 0.78, 
    0.82, 0.74, 0.7, 0.66, 0.66, 0.66, 0.66, 0.65, 0.65, 0.6, 0.57, 0.55, 
    0.53, 0.54, 0.53, 0.45, 0.33, 0.38, 0.37, 0.33, 0.37, 0.4, 0.4, 0.43, 
    0.48, 0.47, 0.51, 0.53, 0.55, 0.57, 0.53, 0.57, 0.54, 0.53, 0.52, 0.47, 
    0.46, 0.45, 0.46, 0.44, 0.48, 0.46, 0.5, 0.52, 0.56, 0.51, 0.67, 0.58, 
    0.5, 0.65, 0.59, 0.5, 0.57, 0.53, 0.56, 0.53, 0.59, 0.56, 0.53, 0.47, 
    0.45, 0.47, 0.46, 0.53, 0.47, 0.54, 0.55, 0.56, 0.59, 0.62, 0.66, 0.71, 
    0.75, 0.77, 0.79, 0.81, 0.79, 0.76, 0.74, 0.66, 0.58, 0.57, 0.57, 0.57, 
    0.66, 0.58, 0.55, 0.51, 0.54, 0.69, 0.75, 0.82, 0.88, 0.9, 0.92, 0.93, 
    0.93, 0.92, 0.88, 0.9, 0.89, 0.82, 0.71, 0.68, 0.69, 0.71, 0.68, 0.68, 
    0.68, 0.77, 0.79, 0.88, 0.89, 0.89, 0.9, 0.9, 0.91, 0.92, 0.92, 0.91, 
    0.92, 0.94, 0.94, 0.92, 0.92, 0.87, 0.85, 0.79, 0.83, 0.78, 0.73, 0.64, 
    0.64, 0.58, 0.65, 0.67, 0.65, 0.74, 0.8, 0.79, 0.76, 0.83, 0.82, 0.85, 
    0.84, 0.85, 0.85, 0.87, 0.85, 0.84, 0.84, 0.85, 0.82, 0.81, 0.82, 0.83, 
    0.84, 0.83, 0.82, 0.84, 0.86, 0.87, 0.87, 0.88, 0.89, 0.9, 0.91, 0.9, 
    0.89, 0.88, 0.88, 0.91, 0.92, 0.93, 0.91, 0.86, 0.86, 0.81, 0.79, 0.75, 
    0.73, 0.71, 0.67, 0.71, 0.68, 0.74, 0.79, 0.75, 0.82, 0.81, 0.84, 0.81, 
    0.79, 0.76, 0.75, 0.72, 0.76, 0.78, 0.79, 0.82, 0.75, 0.79, 0.75, 0.76, 
    0.71, 0.7, 0.69, 0.73, 0.83, 0.88, 0.89, 0.77, 0.67, 0.64, 0.6, 0.49, 
    0.55, 0.5, 0.47, 0.42, 0.33, 0.47, 0.46, 0.5, 0.53, 0.5, 0.46, 0.46, 
    0.44, 0.44, 0.45, 0.48, 0.51, 0.47, 0.46, 0.55, 0.52, 0.48, 0.45, 0.52, 
    0.5, 0.53, 0.61, 0.58, 0.6, 0.6, 0.6, 0.59, 0.55, 0.54, 0.53, 0.52, 0.5, 
    0.48, 0.53, 0.52, 0.52, 0.52, 0.57, 0.63, 0.66, 0.58, 0.57, 0.53, 0.55, 
    0.53, 0.51, 0.53, 0.5, 0.48, 0.53, 0.49, 0.45, 0.42, 0.47, 0.51, 0.47, 
    0.56, 0.46, 0.47, 0.49, 0.47, 0.51, 0.39, 0.5, 0.6, 0.64, 0.65, 0.66, 
    0.75, 0.71, 0.7, 0.64, 0.69, 0.71, 0.62, 0.58, 0.63, 0.64, 0.54, 0.61, 
    0.6, 0.59, 0.59, 0.55, 0.5, 0.57, 0.56, 0.58, 0.58, 0.54, 0.6, 0.59, 
    0.64, 0.57, 0.68, 0.62, 0.58, 0.48, 0.51, 0.49, 0.48, 0.45, 0.45, 0.49, 
    0.44, 0.44, 0.45, 0.48, 0.45, 0.46, 0.46, 0.49, 0.52, 0.57, 0.53, 0.57, 
    0.59, 0.62, 0.62, 0.61, 0.61, 0.6, 0.57, 0.54, 0.53, 0.51, 0.53, 0.54, 
    0.55, 0.57, 0.56, 0.56, 0.58, 0.56, 0.55, 0.57, 0.6, 0.63, 0.63, 0.64, 
    0.63, 0.65, 0.62, 0.66, 0.65, 0.63, 0.6, 0.65, 0.66, 0.62, 0.63, 0.6, 
    0.61, 0.58, 0.57, 0.61, 0.62, 0.57, 0.6, 0.61, 0.59, 0.66, 0.66, 0.63, 
    0.65, 0.68, 0.7, 0.66, 0.67, 0.63, 0.61, 0.61, 0.6, 0.61, 0.61, 0.63, 
    0.63, 0.6, 0.58, 0.58, 0.62, 0.6, 0.62, 0.58, 0.6, 0.64, 0.65, 0.68, 
    0.65, 0.68, 0.67, 0.66, 0.6, 0.61, 0.62, 0.63, 0.57, 0.56, 0.72, 0.55, 
    0.53, 0.53, 0.5, 0.5, 0.51, 0.53, 0.53, 0.56, 0.57, 0.5, 0.56, 0.55, 
    0.56, 0.55, 0.56, 0.59, 0.55, 0.51, 0.49, 0.5, 0.49, 0.5, 0.5, 0.52, 
    0.54, 0.51, 0.5, 0.52, 0.54, 0.6, 0.54, 0.52, 0.56, 0.61, 0.57, 0.58, 
    0.63, 0.68, 0.68, 0.69, 0.64, 0.66, 0.64, 0.65, 0.65, 0.64, 0.63, 0.63, 
    0.62, 0.65, 0.62, 0.65, 0.61, 0.65, 0.64, 0.63, 0.63, 0.65, 0.7, 0.7, 
    0.76, 0.77, 0.79, 0.77, 0.66, 0.66, 0.65, 0.59, 0.59, 0.6, 0.62, 0.57, 
    0.56, 0.59, 0.59, 0.66, 0.63, 0.67, 0.66, 0.62, 0.64, 0.71, 0.63, 0.67, 
    0.72, 0.73, 0.72, 0.77, 0.72, 0.72, 0.77, 0.76, 0.7, 0.62, 0.66, 0.68, 
    0.69, 0.72, 0.63, 0.6, 0.66, 0.69, 0.7, 0.71, 0.74, 0.73, 0.73, 0.71, 
    0.72, 0.72, 0.68, 0.66, 0.64, 0.66, 0.66, 0.68, 0.58, 0.57, 0.74, 0.83, 
    0.84, 0.84, 0.64, 0.63, 0.66, 0.72, 0.72, 0.69, 0.66, 0.67, 0.72, 0.66, 
    0.7, 0.7, 0.73, 0.73, 0.76, 0.72, 0.77, 0.75, 0.79, 0.78, 0.77, 0.77, 
    0.89, 0.79, 0.89, 0.87, 0.92, 0.93, 0.93, 0.94, 0.94, 0.94, 0.95, 0.95, 
    0.94, 0.95, 0.96, 0.96, 0.94, 0.92, 0.88, 0.91, 0.88, 0.88, 0.88, 0.88, 
    0.82, 0.72, 0.74, 0.76, 0.76, 0.67, 0.7, 0.65, 0.67, 0.68, 0.64, 0.66, 
    0.65, 0.67, 0.65, 0.66, 0.66, 0.66, 0.65, 0.55, 0.66, 0.68, 0.7, 0.65, 
    0.68, 0.67, 0.64, 0.6, 0.71, 0.66, 0.67, 0.68, 0.69, 0.73, 0.74, 0.75, 
    0.76, 0.78, 0.76, 0.76, 0.76, 0.73, 0.72, 0.71, 0.71, 0.71, 0.71, 0.68, 
    0.68, 0.68, 0.69, 0.69, 0.71, 0.71, 0.7, 0.69, 0.7, 0.72, 0.73, 0.74, 
    0.73, 0.77, 0.78, 0.78, 0.79, 0.77, 0.76, 0.73, 0.74, 0.78, 0.72, 0.72, 
    0.68, 0.72, 0.7, 0.65, 0.67, 0.7, 0.71, 0.73, 0.73, 0.74, 0.78, 0.81, 
    0.78, 0.78, 0.72, 0.75, 0.78, 0.73, 0.75, 0.76, 0.75, 0.73, 0.74, 0.72, 
    0.72, 0.73, 0.71, 0.71, 0.72, 0.71, 0.68, 0.71, 0.7, 0.7, 0.69, 0.67, 
    0.67, 0.68, 0.66, 0.67, 0.67, 0.67, 0.69, 0.67, 0.65, 0.64, 0.65, 0.67, 
    0.68, 0.71, 0.73, 0.72, 0.73, 0.73, 0.72, 0.7, 0.71, 0.7, 0.69, 0.7, 
    0.69, 0.71, 0.73, 0.7, 0.69, 0.71, 0.71, 0.68, 0.66, 0.7, 0.67, 0.65, 
    0.64, 0.62, 0.64, 0.65, 0.64, 0.62, 0.6, 0.61, 0.64, 0.62, 0.64, 0.68, 
    0.63, 0.67, 0.67, 0.66, 0.63, 0.64, 0.65, 0.62, 0.66, 0.64, 0.61, 0.58, 
    0.64, 0.67, 0.7, 0.71, 0.62, 0.62, 0.56, 0.53, 0.58, 0.54, 0.58, 0.63, 
    0.61, 0.63, 0.6, 0.58, 0.58, 0.56, 0.63, 0.59, 0.57, 0.59, 0.57, 0.59, 
    0.62, 0.58, 0.6, 0.56, 0.58, 0.6, 0.66, 0.61, 0.58, 0.58, 0.62, 0.62, 
    0.61, 0.58, 0.63, 0.65, 0.64, 0.69, 0.77, 0.65, 0.61, 0.59, 0.6, 0.59, 
    0.58, 0.64, 0.55, 0.52, 0.48, 0.46, 0.45, 0.49, 0.53, 0.56, 0.55, 0.58, 
    0.55, 0.59, 0.63, 0.6, 0.61, 0.58, 0.57, 0.6, 0.65, 0.66, 0.58, 0.62, 
    0.7, 0.63, 0.61, 0.6, 0.56, 0.65, 0.67, 0.6, 0.59, 0.6, 0.55, 0.52, 0.54, 
    0.53, 0.53, 0.54, 0.5, 0.53, 0.51, 0.77, 0.5, 0.72, 0.51, 0.68, 0.5, 0.5, 
    0.47, 0.47, 0.49, 0.45, 0.47, 0.5, 0.53, 0.55, 0.53, 0.62, 0.61, 0.63, 
    0.67, 0.65, 0.58, 0.59, 0.54, 0.48, 0.48, 0.5, 0.48, 0.52, 0.55, 0.5, 
    0.5, 0.47, 0.48, 0.53, 0.49, 0.53, 0.6, 0.58, 0.61, 0.62, 0.62, 0.6, 
    0.61, 0.66, 0.66, 0.66, 0.66, 0.68, 0.69, 0.66, 0.7, 0.65, 0.67, 0.64, 
    0.66, 0.68, 0.67, 0.75, 0.64, 0.68, 0.69, 0.73, 0.77, 0.9, 0.88, 0.91, 
    0.88, 0.89, 0.89, 0.87, 0.89, 0.92, 0.9, 0.88, 0.86, 0.85, 0.83, 0.7, 
    0.62, 0.64, 0.64, 0.72, 0.67, 0.66, 0.65, 0.66, 0.68, 0.72, 0.65, 0.7, 
    0.71, 0.64, 0.63, 0.56, 0.59, 0.57, 0.57, 0.59, 0.57, 0.53, 0.47, 0.49, 
    0.56, 0.59, 0.58, 0.58, 0.62, 0.65, 0.66, 0.62, 0.61, 0.59, 0.6, 0.61, 
    0.62, 0.57, 0.56, 0.67, 0.64, 0.67, 0.67, 0.66, 0.64, 0.51, 0.59, 0.56, 
    0.55, 0.53, 0.54, 0.54, 0.53, 0.53, 0.48, 0.57, 0.54, 0.44, 0.47, 0.47, 
    0.49, 0.51, 0.55, 0.55, 0.57, 0.57, 0.57, 0.57, 0.55, 0.58, 0.59, 0.56, 
    0.6, 0.57, 0.61, 0.54, 0.51, 0.54, 0.56, 0.63, 0.61, 0.66, 0.7, 0.72, 
    0.72, 0.64, 0.56, 0.58, 0.59, 0.55, 0.55, 0.56, 0.58, 0.59, 0.6, 0.61, 
    0.58, 0.56, 0.58, 0.57, 0.59, 0.64, 0.6, 0.61, 0.64, 0.71, 0.74, 0.73, 
    0.74, 0.75, 0.74, 0.73, 0.72, 0.67, 0.7, 0.69, 0.69, 0.69, 0.67, 0.68, 
    0.68, 0.79, 0.75, 0.72, 0.75, 0.73, 0.69, 0.73, 0.7, 0.72, 0.71, 0.71, 
    0.72, 0.72, 0.71, 0.73, 0.72, 0.72, 0.71, 0.72, 0.73, 0.68, 0.65, 0.64, 
    0.67, 0.66, 0.66, 0.68, 0.69, 0.65, 0.65, 0.67, 0.73, 0.75, 0.75, 0.73, 
    0.72, 0.71, 0.7, 0.67, 0.67, 0.66, 0.63, 0.67, 0.64, 0.65, 0.66, 0.65, 
    0.71, 0.76, 0.67, 0.7, 0.68, 0.63, 0.75, 0.83, 0.83, 0.79, 0.74, 0.74, 
    0.66, 0.74, 0.73, 0.83, 0.67, 0.8, 0.67, 0.67, 0.69, 0.69, 0.67, 0.67, 
    0.68, 0.68, 0.7, 0.69, 0.75, 0.78, 0.78, 0.73, 0.72, 0.67, 0.63, 0.66, 
    0.73, 0.78, 0.71, 0.7, 0.7, 0.68, 0.66, 0.66, 0.65, 0.69, 0.68, 0.67, 
    0.67, 0.68, 0.66, 0.76, 0.73, 0.69, 0.7, 0.67, 0.66, 0.69, 0.7, 0.73, 
    0.73, 0.72, 0.7, 0.65, 0.64, 0.61, 0.59, 0.57, 0.6, 0.62, 0.63, 0.62, 
    0.62, 0.72, 0.67, 0.77, 0.72, 0.71, 0.69, 0.68, 0.64, 0.68, 0.67, 0.63, 
    0.65, 0.6, 0.64, 0.61, 0.65, 0.61, 0.62, 0.64, 0.63, 0.61, 0.6, 0.65, 
    0.62, 0.62, 0.57, 0.59, 0.58, 0.57, 0.57, 0.62, 0.62, 0.68, 0.71, 0.7, 
    0.67, 0.7, 0.63, 0.55, 0.5, 0.5, 0.49, 0.53, 0.53, 0.52, 0.51, 0.38, 
    0.53, 0.5, 0.53, 0.47, 0.51, 0.48, 0.45, 0.48, 0.55, 0.54, 0.59, 0.62, 
    0.63, 0.62, 0.52, 0.56, 0.56, 0.57, 0.51, 0.47, 0.5, 0.48, 0.54, 0.6, 
    0.68, 0.71, 0.84, 0.76, 0.74, 0.79, 0.8, 0.77, 0.68, 0.65, 0.67, 0.69, 
    0.68, 0.67, 0.62, 0.61, 0.59, 0.6, 0.62, 0.72, 0.74, 0.77, 0.7, 0.72, 
    0.73, 0.74, 0.76, 0.76, 0.77, 0.78, 0.83, 0.83, 0.8, 0.79, 0.78, 0.78, 
    0.84, 0.81, 0.81, 0.81, 0.85, 0.76, 0.68, 0.69, 0.71, 0.72, 0.73, 0.74, 
    0.69, 0.69, 0.68, 0.75, 0.79, 0.84, 0.82, 0.87, 0.89, 0.87, 0.89, 0.86, 
    0.85, 0.83, 0.86, 0.87, 0.89, 0.88, 0.86, 0.83, 0.81, 0.79, 0.8, 0.82, 
    0.76, 0.74, 0.8, 0.76, 0.89, 0.89, 0.86, 0.77, 0.83, 0.84, 0.83, 0.87, 
    0.86, 0.82, 0.75, 0.86, 0.85, 0.85, 0.91, 0.84, 0.92, 0.92, 0.78, 0.69, 
    0.62, 0.64, 0.47, 0.53, 0.55, 0.53, 0.53, 0.58, 0.61, 0.61, 0.62, 0.66, 
    0.63, 0.63, 0.62, 0.6, 0.58, 0.85, 0.56, 0.58, 0.54, 0.53, 0.57, 0.56, 
    0.59, 0.54, 0.53, 0.58, 0.6, 0.6, 0.63, 0.62, 0.6, 0.63, 0.61, 0.61, 
    0.59, 0.63, 0.63, 0.65, 0.66, 0.64, 0.62, 0.62, 0.65, 0.71, 0.77, 0.71, 
    0.75, 0.7, 0.63, 0.64, 0.62, 0.64, 0.68, 0.67, 0.67, 0.71, 0.65, 0.65, 
    0.78, 0.71, 0.71, 0.66, 0.66, 0.6, 0.54, 0.58, 0.51, 0.58, 0.56, 0.61, 
    0.6, 0.64, 0.63, 0.59, 0.58, 0.68, 0.7, 0.66, 0.65, 0.65, 0.7, 0.74, 
    0.73, 0.71, 0.68, 0.66, 0.65, 0.63, 0.66, 0.73, 0.66, 0.64, 0.62, 0.62, 
    0.63, 0.62, 0.61, 0.58, 0.59, 0.6, 0.61, 0.6, 0.59, 0.6, 0.64, 0.75, 
    0.73, 0.67, 0.71, 0.66, 0.75, 0.73, 0.71, 0.76, 0.75, 0.73, 0.68, 0.63, 
    0.56, 0.58, 0.72, 0.6, 0.72, 0.77, 0.82, 0.85, 0.86, 0.85, 0.86, 0.87, 
    0.83, 0.82, 0.8, 0.79, 0.8, 0.78, 0.79, 0.76, 0.75, 0.76, 0.76, 0.77, 
    0.81, 0.82, 0.63, 0.74, 0.73, 0.81, 0.76, 0.76, 0.74, 0.75, 0.7, 0.74, 
    0.85, 0.77, 0.79, 0.79, 0.72, 0.69, 0.66, 0.65, 0.64, 0.64, 0.64, 0.65, 
    0.67, 0.66, 0.54, 0.58, 0.55, 0.6, 0.69, 0.67, 0.59, 0.72, 0.67, 0.68, 
    0.69, 0.69, 0.68, 0.67, 0.66, 0.66, 0.72, 0.69, 0.65, 0.67, 0.65, 0.66, 
    0.65, 0.69, 0.75, 0.83, 0.82, 0.79, 0.84, 0.85, 0.85, 0.79, 0.8, 0.75, 
    0.74, 0.77, 0.79, 0.78, 0.79, 0.74, 0.71, 0.69, 0.66, 0.58, 0.41, 0.39, 
    0.51, 0.47, 0.5, 0.54, 0.57, 0.59, 0.7, 0.68, 0.69, 0.72, 0.75, 0.76, 
    0.74, 0.75, 0.78, 0.81, 0.76, 0.68, 0.66, 0.69, 0.71, 0.72, 0.73, 0.64, 
    0.61, 0.63, 0.61, 0.73, 0.76, 0.75, 0.72, 0.77, 0.75, 0.88, 0.74, 0.75, 
    0.75, 0.71, 0.69, 0.68, 0.7, 0.72, 0.7, 0.67, 0.64, 0.65, 0.65, 0.63, 
    0.66, 0.65, 0.65, 0.66, 0.68, 0.68, 0.67, 0.66, 0.68, 0.68, 0.67, 0.66, 
    0.69, 0.7, 0.68, 0.67, 0.66, 0.7, 0.77, 0.75, 0.73, 0.67, 0.63, 0.61, 
    0.61, 0.63, 0.63, 0.62, 0.64, 0.64, 0.66, 0.63, 0.65, 0.73, 0.8, 0.78, 
    0.74, 0.66, 0.64, 0.61, 0.57, 0.58, 0.51, 0.55, 0.53, 0.57, 0.57, 0.56, 
    0.56, 0.57, 0.56, 0.58, 0.56, 0.56, 0.55, 0.59, 0.59, 0.61, 0.63, 0.55, 
    0.59, 0.59, 0.63, 0.57, 0.65, 0.65, 0.69, 0.57, 0.57, 0.57, 0.56, 0.57, 
    0.56, 0.55, 0.54, 0.55, 0.62, 0.52, 0.54, 0.57, 0.72, 0.67, 0.6, 0.63, 
    0.61, 0.55, 0.63, 0.58, 0.57, 0.55, 0.54, 0.59, 0.64, 0.58, 0.56, 0.54, 
    0.52, 0.6, 0.59, 0.57, 0.57, 0.62, 0.49, 0.47, 0.48, 0.47, 0.46, 0.44, 
    0.49, 0.53, 0.6, 0.57, 0.55, 0.54, 0.52, 0.53, 0.57, 0.59, 0.57, 0.55, 
    0.5, 0.47, 0.48, 0.52, 0.48, 0.48, 0.45, 0.51, 0.51, 0.53, 0.52, 0.52, 
    0.53, 0.53, 0.54, 0.55, 0.61, 0.6, 0.62, 0.63, 0.62, 0.63, 0.67, 0.7, 
    0.62, 0.63, 0.67, 0.66, 0.58, 0.56, 0.65, 0.7, 0.68, 0.71, 0.69, 0.67, 
    0.67, 0.75, 0.77, 0.77, 0.77, 0.74, 0.77, 0.79, 0.79, 0.79, 0.75, 0.75, 
    0.77, 0.81, 0.8, 0.79, 0.77, 0.79, 0.81, 0.8, 0.85, 0.86, 0.88, 0.89, 
    0.9, 0.86, 0.83, 0.8, 0.83, 0.79, 0.74, 0.73, 0.73, 0.7, 0.69, 0.71, 
    0.64, 0.7, 0.63, 0.58, 0.62, 0.59, 0.62, 0.63, 0.65, 0.64, 0.64, 0.56, 
    0.53, 0.57, 0.61, 0.57, 0.51, 0.46, 0.49, 0.48, 0.49, 0.56, 0.7, 0.69, 
    0.61, 0.58, 0.63, 0.62, 0.72, 0.72, 0.74, 0.79, 0.78, 0.75, 0.84, 0.88, 
    0.86, 0.89, 0.87, 0.85, 0.83, 0.79, 0.75, 0.72, 0.81, 0.79, 0.78, 0.78, 
    0.78, 0.76, 0.6, 0.67, 0.79, 0.55, 0.62, 0.66, 0.74, 0.75, 0.78, 0.76, 
    0.8, 0.79, 0.76, 0.76, 0.73, 0.72, 0.68, 0.63, 0.63, 0.61, 0.68, 0.69, 
    0.75, 0.71, 0.76, 0.84, 0.83, 0.83, 0.8, 0.76, 0.79, 0.82, 0.78, 0.8, 
    0.8, 0.77, 0.77, 0.79, 0.69, 0.67, 0.65, 0.67, 0.65, 0.63, 0.64, 0.66, 
    0.66, 0.64, 0.65, 0.66, 0.76, 0.78, 0.74, 0.8, 0.84, 0.84, 0.83, 0.84, 
    0.83, 0.86, 0.83, 0.87, 0.85, _, 0.87, 0.86, 0.85, 0.82, 0.83, 0.78, 0.8, 
    0.76, 0.76, 0.78, 0.78, 0.74, 0.77, 0.77, 0.72, 0.78, 0.81, 0.87, 0.85, 
    0.83, 0.84, 0.85, 0.8, 0.85, 0.86, 0.88, 0.89, 0.89, 0.89, 0.89, 0.88, 
    0.86, 0.88, 0.88, 0.9, 0.9, 0.92, 0.92, 0.93, 0.93, 0.93, 0.93, 0.92, 
    0.92, 0.92, 0.92, 0.91, 0.9, 0.91, 0.9, 0.87, 1, 0.87, 0.9, 0.86, 0.81, 
    0.84, 0.84, 0.83, 0.84, 0.85, 0.76, 0.77, 0.77, 0.76, 0.78, 0.8, 0.83, 
    0.81, 0.75, 0.77, 0.74, 0.69, 0.71, 0.72, 0.68, 0.69, 0.68, 0.69, 0.67, 
    0.68, 0.67, 0.66, 0.69, 0.72, 0.71, 0.73, 0.76, 0.76, 0.76, 0.78, 0.78, 
    0.78, 0.73, 0.73, 0.75, 0.77, 0.75, 0.71, 0.72, 0.69, 0.7, 0.67, 0.62, 
    0.66, 0.82, 0.94, 0.82, 0.83, 0.79, 0.79, 0.77, 0.72, 0.72, 0.73, 0.7, 
    0.71, 0.71, 0.66, 0.72, 0.73, 0.79, 0.78, 0.83, 0.84, 0.86, 0.85, 0.75, 
    0.76, 0.8, 0.84, 0.89, 0.91, 0.9, 0.87, 0.86, 0.88, 0.87, 0.87, 0.83, 
    0.84, 0.84, 0.82, 0.81, 0.79, 0.78, 0.77, 0.76, 0.77, 0.78, 0.79, 0.77, 
    0.8, 0.8, 0.79, 0.83, 0.85, 0.86, 0.85, 0.87, 0.88, 0.88, 0.87, 0.86, 
    0.85, 0.84, 0.86, 0.82, 0.84, 0.8, 0.83, 0.79, 0.89, 0.8, 0.78, 0.78, 
    0.74, 0.8, 0.8, 0.82, 0.79, 0.82, 0.83, 0.83, 0.84, 0.84, 0.82, 0.77, 
    0.72, 0.74, 0.72, 0.7, 0.69, 0.66, 0.66, 0.66, 0.68, 0.69, 0.65, 0.68, 
    0.64, 0.64, 0.66, 0.64, 0.67, 0.72, 0.74, 0.75, 0.77, 0.79, 0.79, 0.78, 
    0.76, 0.68, 0.67, 0.67, 0.66, 0.67, 0.68, 0.67, 0.68, 0.7, 0.68, 0.6, 
    0.64, 0.68, 0.67, 0.67, 0.64, 0.64, 0.71, 0.75, 0.71, 0.69, 0.7, 0.7, 
    0.71, 0.72, 0.74, 0.84, 0.76, 0.8, 0.72, 0.75, 0.68, 0.77, 0.7, 0.76, 
    0.77, 0.76, 0.83, 0.82, 0.81, 0.77, 0.81, 0.79, 0.78, 0.77, 0.8, 0.81, 
    0.8, 0.82, 0.79, 0.81, 0.71, 0.71, 0.74, 0.69, 0.69, 0.71, 0.71, 0.68, 
    0.75, 0.8, 0.75, 0.76, 0.73, 0.76, 0.73, 0.69, 0.7, 0.66, 0.66, 0.67, 
    0.74, 0.73, 0.77, 0.72, 0.72, 0.68, 0.66, 0.71, 0.72, 0.81, 0.93, 0.79, 
    0.76, 0.76, 0.75, 0.81, 0.77, 0.77, 0.82, 0.79, 0.84, 0.86, 0.85, 0.83, 
    0.85, 0.86, 0.78, 0.75, 0.7, 0.71, 0.75, 0.92, 0.78, 0.9, 0.81, 0.9, 0.9, 
    0.91, 0.94, 0.93, 0.91, 0.91, 0.9, 0.86, 0.85, 0.86, 0.86, 0.87, 0.84, 
    0.73, 0.75, 0.72, 0.68, 0.66, 0.66, 0.66, 0.66, 0.75, 0.78, 0.75, 0.73, 
    0.72, 0.8, 0.8, 0.78, 0.79, 0.8, 0.84, 0.82, 0.8, 0.78, 0.76, 0.75, 0.75, 
    0.63, 0.62, 0.63, 0.65, 0.62, 0.65, 0.6, 0.59, 0.55, 0.55, 0.54, 0.59, 
    0.58, 0.62, 0.66, 0.63, 0.67, 0.7, 0.68, 0.69, 0.71, 0.72, 0.71, 0.68, 
    0.76, 0.71, 0.7, 0.65, 0.62, 0.61, 0.62, 0.65, 0.72, 0.71, 0.68, 0.78, 
    0.7, 0.82, 0.81, 0.83, 0.81, 0.76, 0.82, 0.82, 0.82, 0.77, 0.78, 0.75, 
    0.74, 0.69, 0.69, 0.67, 0.69, 0.68, 0.63, 0.58, 0.52, 0.54, 0.53, 0.52, 
    0.54, 0.62, 0.7, 0.74, 0.76, 0.75, 0.78, 0.78, 0.78, 0.7, 0.67, 0.62, 
    0.62, 0.59, 0.56, 0.55, 0.56, 0.52, 0.53, 0.53, 0.55, 0.51, 0.54, 0.52, 
    0.51, 0.54, 0.54, 0.6, 0.6, 0.58, 0.61, 0.59, 0.58, 0.56, 0.57, 0.55, 
    0.54, 0.5, 0.46, 0.46, 0.46, 0.45, 0.42, 0.41, 0.41, 0.42, 0.39, 0.39, 
    0.39, 0.38, 0.42, 0.47, 0.45, 0.5, 0.53, 0.63, 0.59, 0.7, 0.67, 0.73, 
    0.69, 0.73, 0.67, 0.67, 0.65, 0.73, 0.69, 0.66, 0.67, 0.74, 0.79, 0.83, 
    0.82, 0.76, 0.79, 0.85, 0.76, 0.78, 0.79, 0.79, 0.79, 0.78, 0.82, 0.82, 
    0.79, 0.79, 0.81, 0.82, 0.83, 0.82, 0.84, 0.84, 0.85, 0.83, 0.84, 0.83, 
    0.81, 0.85, 0.86, 0.86, 0.85, 0.85, 0.87, 0.87, 0.87, 0.87, 0.9, 0.87, 
    0.88, 0.87, 0.83, 0.82, 0.82, 0.82, 0.82, 0.77, 0.72, 0.62, 0.58, 0.53, 
    0.49, 0.5, 0.52, 0.59, 0.63, 0.69, 0.72, 0.74, 0.75, 0.77, 0.69, 0.78, 
    0.74, 0.96, 0.98, 0.96, 0.94, 0.92, 0.91, 0.91, 0.89, 0.88, 0.86, 0.85, 
    0.84, 0.84, 0.84, 0.79, 0.83, 0.76, 0.76, 0.76, 0.78, 0.79, 0.85, 0.86, 
    0.83, 0.78, 0.79, 0.75, 0.72, 0.73, 0.75, 0.71, 0.67, 0.66, 0.6, 0.7, 
    0.69, 0.7, 0.78, 0.8, 0.82, 0.83, 0.82, 0.83, 0.84, 0.83, 0.81, 0.81, 
    0.81, 0.81, 0.8, 0.78, 0.8, 0.75, 0.75, 0.73, 0.72, 0.7, 0.78, 0.86, 
    0.85, 0.88, 0.87, 0.86, 0.87, 0.88, 0.88, 0.88, 0.88, 0.91, 0.89, 0.89, 
    0.87, 0.87, 0.87, 0.88, 0.85, 0.84, 0.83, 0.82, 0.81, 0.8, 0.81, 0.79, 
    0.77, 0.78, 0.79, 0.76, 0.75, 0.71, 0.71, 0.72, 0.73, 0.75, 0.7, 0.66, 
    0.69, 0.7, 0.71, 0.69, 0.69, 0.54, 0.59, 0.54, 0.54, 0.58, 0.55, 0.57, 
    0.65, 0.66, 0.7, 0.74, 0.75, 0.78, 0.76, 0.78, 0.79, 0.84, 0.78, 0.72, 
    0.77, 0.69, 0.63, 0.66, 0.71, 0.65, 0.64, 0.64, 0.58, 0.59, 0.63, 0.67, 
    0.68, 0.68, 0.71, 0.7, 0.67, 0.65, 0.65, 0.64, 0.62, 0.59, 0.55, 0.56, 
    0.54, 0.55, 0.53, 0.52, 0.52, 0.53, 0.53, 0.51, 0.5, 0.55, 0.55, 0.57, 
    0.62, 0.64, 0.67, 0.71, 0.7, 0.69, 0.71, 0.7, 0.7, 0.71, 0.7, 0.72, 0.72, 
    0.71, 0.71, 0.66, 0.59, 0.61, 0.61, 0.57, 0.58, 0.58, 0.58, 0.58, 0.59, 
    0.64, 0.63, 0.63, 0.67, 0.71, 0.73, 0.74, 0.75, 0.74, 0.71, 0.7, 0.68, 
    0.66, 0.64, 0.65, 0.65, 0.67, 0.69, 0.69, 0.65, 0.64, 0.65, 0.64, 0.6, 
    0.61, 0.59, 0.56, 0.58, 0.6, 0.64, 0.68, 0.7, 0.73, 0.75, 0.73, 0.73, 
    0.69, 0.7, 0.68, 0.66, 0.65, 0.66, 0.66, 0.64, 0.65, 0.62, 0.6, 0.59, 
    0.64, 0.57, 0.63, 0.66, 0.64, 0.62, 0.62, 0.62, 0.65, 0.66, 0.63, 0.61, 
    0.58, 0.62, 0.59, 0.59, 0.57, 0.54, 0.54, 0.56, 0.54, 0.58, 0.57, 0.64, 
    0.67, 0.63, 0.67, 0.69, 0.72, 0.74, 0.7, 0.64, 0.5, 0.51, 0.49, 0.51, 
    0.53, 0.51, 0.53, 0.56, 0.58, 0.55, 0.59, 0.57, 0.58, 0.56, 0.56, 0.57, 
    0.58, 0.59, 0.61, 0.61, 0.6, 0.6, 0.6, 0.62, 0.64, 0.63, 0.64, 0.63, 
    0.64, 0.63, 0.6, 0.6, 0.6, 0.55, 0.52, 0.53, 0.54, 0.54, 0.6, 0.64, 0.67, 
    0.52, 0.56, 0.58, 0.61, 0.62, 0.67, 0.71, 0.64, 0.61, 0.63, 0.62, 0.55, 
    0.55, 0.55, 0.53, 0.53, 0.51, 0.5, 0.5, 0.5, 0.51, 0.52, 0.55, 0.61, 
    0.62, 0.61, 0.68, 0.68, 0.67, 0.76, 0.73, 0.73, 0.74, 0.75, 0.74, 0.76, 
    0.78, 0.8, 0.86, 0.87, 0.85, 0.83, 0.84, 0.82, 0.87, 0.87, 0.88, 0.88, 
    0.9, 0.89, 0.93, 0.95, 0.95, 0.94, 0.96, 0.97, 0.91, 0.7, 0.69, 0.66, 
    0.7, 0.67, 0.69, 0.72, 0.67, 0.68, 0.69, 0.66, 0.65, 0.67, 0.62, 0.7, 
    0.72, 0.75, 0.7, 0.72, 0.68, 0.67, 0.67, 0.67, 0.7, 0.66, 0.65, 0.66, 
    0.65, 0.68, 0.64, 0.62, 0.58, 0.6, 0.61, 0.62, 0.63, 0.66, 0.64, 0.72, 
    0.7, 0.71, 0.72, 0.75, 0.77, 0.81, 0.82, 0.8, 0.78, 0.77, 0.75, 0.71, 
    0.71, 0.7, 0.69, 0.66, 0.64, 0.76, 0.76, 0.72, 0.75, 0.75, 0.76, 0.78, 
    0.79, 0.81, 0.83, 0.8, 0.82, 0.82, 0.86, 0.85, 0.83, 0.83, 0.68, 0.61, 
    0.6, 0.58, 0.58, 0.6, 0.6, 0.62, 0.61, 0.65, 0.65, 0.64, 0.62, 0.63, 
    0.64, 0.63, 0.63, 0.63, 0.65, 0.62, 0.63, 0.67, 0.62, 0.64, 0.6, 0.58, 
    0.56, 0.59, 0.55, 0.57, 0.6, 0.58, 0.63, 0.66, 0.69, 0.7, 0.71, 0.68, 
    0.68, 0.68, 0.65, 0.64, 0.63, 0.64, 0.64, 0.6, 0.63, 0.65, 0.66, 0.65, 
    0.62, 0.61, 0.59, 0.52, 0.54, 0.57, 0.52, 0.57, 0.49, 0.52, 0.69, 0.61, 
    0.64, 0.65, 0.64, 0.6, 0.73, 0.74, 0.74, 0.74, 0.74, 0.73, 0.73, 0.67, 
    0.65, 0.65, 0.63, 0.62, 0.6, 0.56, 0.54, 0.48, 0.5, 0.51, 0.55, 0.55, 
    0.59, 0.61, 0.65, 0.72, 0.76, 0.76, 0.74, 0.81, 0.77, 0.63, 0.75, 0.79, 
    0.69, 0.67, 0.67, 0.66, 0.65, 0.65, 0.64, 0.64, 0.64, 0.67, 0.7, 0.72, 
    0.84, 0.85, 0.83, 0.83, 0.81, 0.78, 0.77, 0.78, 0.66, 0.65, 0.76, 0.83, 
    0.74, 0.74, 0.68, 0.72, 0.78, 0.77, 0.8, 0.76, 0.74, 0.71, 0.71, 0.66, 
    0.67, 0.7, 0.73, 0.78, 0.84, 0.89, 0.92, 0.96, 0.96, 0.93, 0.92, 0.71, 
    0.86, 0.85, 0.83, 0.76, 0.72, 0.7, 0.67, 0.68, 0.72, 0.72, 0.76, 0.75, 
    0.79, 0.78, 0.84, 0.85, 0.82, 0.86, 0.86, 0.87, 0.85, 0.81, 0.8, 0.79, 
    0.81, 0.81, 0.79, 0.8, 0.75, 0.69, 0.67, 0.69, 0.58, 0.63, 0.66, 0.74, 
    0.74, 0.69, 0.64, 0.62, 0.63, 0.59, 0.79, 0.76, 0.6, 0.74, 0.72, 0.62, 
    0.6, 0.6, 0.58, 0.54, 0.59, 0.63, 0.64, 0.64, 0.67, 0.67, 0.66, 0.67, 
    0.7, 0.71, 0.69, 0.67, 0.73, 0.71, 0.68, 0.7, 0.71, 0.7, 0.61, 0.67, 0.7, 
    0.72, 0.75, 0.76, 0.79, 0.86, 0.84, 0.81, 0.84, 0.88, 0.94, 0.93, 0.93, 
    0.94, 0.93, 0.95, 0.96, 0.96, 0.97, 0.98, 0.98, 0.93, 0.97, 0.95, 0.95, 
    0.95, 0.94, 0.94, 0.93, 0.91, 0.91, 0.9, 0.89, 0.92, 0.92, 0.89, 0.81, 
    0.81, 0.81, 0.79, 0.83, 0.81, 0.87, 0.91, 0.91, 0.93, 0.92, 0.94, 0.94, 
    0.95, 0.93, 0.85, 0.9, 0.91, 0.83, 0.9, 0.84, 0.89, 0.89, 0.91, 0.87, 
    0.91, 0.91, 0.93, 0.95, 0.91, 0.93, 0.95, 0.95, 0.96, 0.97, 0.98, 0.98, 
    0.98, 0.98, 0.98, 0.98, 0.98, 0.98, 0.96, 0.96, 0.94, 0.92, 0.98, 0.99, 
    0.98, 0.98, 0.98, 0.98, 0.99, 1, 0.99, 0.99, 0.99, 0.99, 0.99, 0.98, 
    0.97, 0.93, 0.92, 0.89, 0.89, 0.84, 0.85, 0.85, 0.84, 0.84, 0.83, 0.83, 
    1, 0.83, 0.83, 0.79, 0.79, 0.77, 0.77, 0.79, 0.8, 0.79, 0.74, 0.74, 0.71, 
    0.66, 0.85, 0.6, 0.66, 0.61, 0.68, 0.67, 0.68, 0.69, 0.7, 0.69, 0.7, 
    0.88, 0.71, 0.82, 0.7, 0.7, 0.68, 0.67, 0.71, 0.7, 0.69, 0.65, 0.63, 
    0.63, 0.66 ;

 surface_air_pressure_2m = _, 100580, 100540, 100540, 100550, 100550, 100540, 
    100530, 100590, 100580, 100600, 100620, 100620, 100620, 100620, 100620, 
    100620, 100630, 100650, 100660, 100560, 100570, 100550, 100550, 100530, 
    100530, 100520, 100510, 100510, 100500, 100500, 100490, 100530, 100530, 
    100520, 100520, 100520, 100510, 100480, 100460, 100450, 100430, 100400, 
    100390, 100340, 100340, 100330, 100320, 100320, 100320, 100290, 100260, 
    100230, 100200, 100180, 100190, 100210, 100200, 100190, 100200, 100200, 
    100200, 100190, 100190, 100170, 100180, 100200, 100210, 100220, 100240, 
    100260, 100140, 100150, 100170, _, 100230, 100260, 100270, 100300, 
    100310, 100360, 100400, 100420, 100460, 100470, 100500, 100500, 100520, 
    100540, 100570, 100560, 100540, 100560, 100560, 100580, 100600, 100620, 
    100600, 100620, 100630, 100630, 100630, 100670, 100670, 100700, 100740, 
    100780, 100810, 100830, 100850, 100860, 100880, 100890, 100900, 100910, 
    100890, 100890, 100900, 100930, 100920, 100930, 100940, 100940, 100920, 
    100910, 100890, 100880, 100860, 100870, 100870, 100870, 100890, 100880, 
    100870, 100890, 100880, 100900, 100930, 100960, 100990, 101040, 101100, 
    101160, 101220, 101280, 101340, 101390, 101450, 101510, 101570, 101610, 
    101650, 101710, 101750, 101760, 101820, 101840, _, _, _, _, _, 101940, 
    101950, _, _, 102120, 102170, 102200, 102230, 102270, 102300, 102310, 
    102310, 102320, 102360, 102380, 102410, 102450, 102490, 102480, 102480, 
    102490, 102520, 102510, 102470, 102450, 102440, 102400, 102450, 102440, 
    102410, 102470, 102460, 102440, 102420, 102420, 102420, 102330, 102310, 
    102290, 102270, 102270, 102270, 102280, 102290, 102300, 102270, 102280, 
    102240, 102230, 102230, 102260, 102300, 102330, 102370, 102390, 102410, 
    102430, 102450, 102430, 102450, 102470, 102510, 102520, 102560, 102590, 
    102640, 102690, 102720, 102740, 102760, 102790, 102830, 102810, 102860, 
    102890, 102910, 102950, 103020, 103040, 103090, 103110, 103130, 101350, 
    103170, 103220, 103220, 103250, 103270, 103310, 103330, 103340, 103370, 
    103350, 103360, 103370, 103380, 103370, 103370, 103350, 103360, 103350, 
    103330, 103320, 103290, 103270, 103290, 103300, 103270, 103260, 103250, 
    103260, 103280, 103270, 103260, 103280, 103280, 103260, 103260, 103250, 
    103220, 103220, 103230, 103220, 103230, 103240, 103270, 103300, 103300, 
    103300, 103300, 103310, 103310, 103320, 103300, 103310, 103320, 103360, 
    103370, 103380, 103350, 103370, 103390, 103390, 103400, 103370, 103370, 
    103360, 103340, 103360, 103360, 103360, 103350, 103350, 103340, 103340, 
    103340, 103340, 103360, 103380, 103380, 103400, 103410, 103450, 103440, 
    103440, 103470, 103470, 103490, 103500, 103510, 103510, 103500, 103550, 
    103580, 103590, 103600, 103610, 103600, 103560, 103550, 103500, 103460, 
    103450, 103430, 103410, 103370, 103340, 103300, 103240, 103200, 103170, 
    103130, 103090, 103050, 102980, 102940, 102910, 102890, 102850, 102830, 
    102780, 102730, 102670, 102630, 102580, 102530, 102480, 102440, 102390, 
    102370, 102310, 102290, 102240, 102230, 102220, 102210, 102180, 102180, 
    102210, 102230, 102250, 102270, 102320, 102330, 102330, 102340, 102350, 
    102350, 102330, 102320, 102320, 102330, 102320, 102340, 102350, 102340, 
    102340, 102330, 102310, 102320, 102320, 102290, 102290, 102260, 102270, 
    102260, 102270, 102260, 102250, 102230, 102200, 102200, 102200, 102180, 
    102180, 102180, 102190, 102190, 102180, 102160, 102150, 102130, 102110, 
    102080, 102060, 102010, 102000, 101970, 101980, 101990, 101990, 101950, 
    101920, 101900, 101880, 101850, 101820, 101810, 101790, 101770, 101750, 
    101720, 101710, 101690, 101650, 101610, 101570, 101560, 101550, 101510, 
    101480, 101480, 101480, 101470, 101450, 101430, 101430, 101390, 101370, 
    101360, 101320, 101310, 101310, 101270, 101240, 101200, 101180, 101130, 
    101070, 101020, 101000, 100970, 100940, 100910, 100890, 100880, 100860, 
    100880, 100870, 100850, 100840, 100830, 100820, 100810, 100810, 100790, 
    100760, 100790, 100840, 100820, 100880, 100900, 100940, 100990, 101050, 
    101100, 101160, 101210, 101240, 101320, 101410, 101480, 101530, 101580, 
    101610, 101640, 101690, 101760, 101830, 101890, 101940, 102010, 102090, 
    102160, 102210, 102270, 102330, 102380, 102440, 102510, 102570, 102630, 
    102690, 102760, 102830, 102900, 102950, 102990, 103020, 103040, 103070, 
    103070, 103020, 103010, 102990, 102930, 102910, 102880, 102820, 102760, 
    102650, 102530, 102450, 102360, 102200, 102080, 101990, 101890, 101840, 
    101810, 101800, 101790, 101790, 101760, 101780, 101780, 101790, 101790, 
    101770, 101790, 101790, 101820, 101850, 101890, 101920, 101960, 101990, 
    102030, 102040, 102050, 102070, 102110, 102100, 102100, 102120, 102140, 
    102130, 102140, 102140, 102170, 102200, 102230, 102210, 102250, 102280, 
    102340, 102390, 102430, 102450, 102460, 102490, 102520, 102540, 102580, 
    102600, 102630, 102680, 102750, 102800, 102820, 102850, 102890, 102930, 
    102940, 102960, 103000, 103030, 103050, 103060, 103090, 103080, 103060, 
    103040, 102990, 102950, 102910, 102870, 102810, 102770, 102740, 102690, 
    102650, 102610, 102590, 102530, 102480, 102440, 102380, 102330, 102290, 
    102250, 102200, 102170, 102170, 102130, 102110, 102070, 102040, 102010, 
    101990, 101980, 101940, 101920, 101910, 101930, 101930, 101900, 101890, 
    101880, 101870, 101870, 101860, 101830, 101830, 101810, 101850, 101890, 
    101900, 101890, 101910, 101910, 101950, 101960, 101970, 101990, 102010, 
    102020, 102040, 102070, 102080, 102080, 102050, 101980, 101940, 101880, 
    101800, 101670, 101550, 101430, 101310, 101180, 101100, 101010, 100920, 
    100840, 100770, 100720, 100640, 100520, 100440, 100380, 100370, 100390, 
    100400, 100420, 100420, 100440, 100440, 100460, 100460, 100470, 100470, 
    100480, 100460, 100450, 100420, 100400, 100370, 100350, 100330, 100340, 
    100320, 100300, 100340, 100390, 100470, 100580, 100670, 100760, 100870, 
    100980, 101110, 101230, 101330, 101420, 101520, 101580, 101690, 101770, 
    101840, 101920, 101940, 102020, 102080, 102130, 102170, 102220, 102280, 
    102330, 102390, 102470, 102540, 102600, 102660, 102710, 102760, 102810, 
    102870, 102910, 102950, 102980, 103010, 103060, 103060, 103070, 103080, 
    103050, 103030, 103010, 102960, 102880, 102810, 102710, 102600, 102460, 
    102320, 102210, 102110, 101970, 101810, 101700, 101620, 101530, 101520, 
    101580, 101680, 101800, 101840, 101920, 102020, 102040, 102160, 102210, 
    102290, 102370, 102380, 102440, 102510, 102580, 102660, 102710, 102730, 
    102760, 102780, 102800, 102850, 102860, 102880, 102900, 102900, 102890, 
    102900, 102900, 102890, 102860, 102840, 102820, 102780, 102750, 102720, 
    102690, 102660, 102630, 102600, 102560, 102470, 102360, 102240, 102150, 
    102020, 101900, 101720, 101600, 101470, 101360, 101280, 101150, 101060, 
    100960, 100870, 100850, 100810, 100770, 100700, 100660, 100600, 100600, 
    100600, 100540, 100530, 100480, 100370, 100280, 100260, 100250, 100260, 
    100320, 100330, 100390, 100470, 100470, 100460, 100560, 100740, 100840, 
    100950, 101070, 101180, 101300, 101410, 101510, 101650, 101790, 101890, 
    101980, 102060, 102130, 102190, 102240, 102290, 102280, 102320, 102360, 
    102340, 102340, 102310, 102270, 102200, 102130, 102070, 102000, 101920, 
    101840, 101770, 101710, 101650, 101570, 101520, 101420, 101350, 101280, 
    101190, 101130, 101060, 100950, 100880, 100820, 100750, 100650, 100590, 
    100520, 100490, 100440, 100400, 100350, 100310, 100240, 100200, 100150, 
    100100, 100020, 99960, 99880, 99810, 99750, 99730, 99710, 99700, 99700, 
    99710, 99730, 99760, 99750, 99760, 99760, 99750, 99760, 99750, 99750, 
    99720, 99710, 99730, 99730, 99720, 99700, 99670, 99620, 99560, 99510, 
    99410, 99370, 99370, 99330, 99250, 99170, 99150, 99130, 99100, 99050, 
    98980, 98940, 98910, 98880, 98840, 98790, 98740, 98710, 98700, 98670, 
    98640, 98580, 98540, 98520, 98530, 98530, 98540, 98550, 98570, 98600, 
    98650, 98700, 98720, 98740, 98760, 98810, 98860, 98920, 98980, 99010, 
    99050, 99120, 99210, 99260, 99320, 99370, 99440, 99530, 99610, 99700, 
    99770, 99860, 99910, 99970, 100030, 100090, 100150, 100200, 100220, 
    100280, 100310, 100320, 100330, 100350, 100380, 100380, 100400, 100390, 
    100380, 100370, 100310, 100270, 100180, 100060, 99960, 99900, 99860, 
    99830, 99810, 99780, 99760, 99750, 99790, 99840, 99890, 99910, 99910, 
    99930, 100010, 100060, 100150, 100230, 100290, 100320, 100350, 100400, 
    100390, 100430, 100460, 100480, 100510, 100520, 100560, 100590, 100580, 
    100570, 100550, 100480, 100380, 100300, 100250, 100220, 100180, 100170, 
    100190, 100180, 100180, 100170, 100100, 100050, 99990, 99980, 99980, 
    99980, 99960, 99950, 99930, 99940, 99920, 99890, 99830, 99820, 99730, 
    99680, 99650, 99610, 99580, 99540, 99500, 99490, 99430, 99400, 99420, 
    99380, 99360, 99370, 99360, 99330, 99300, 99230, 99320, 99270, 99270, 
    99310, 99330, 99340, 99330, 99360, 99400, 99400, 99440, 99460, 99490, 
    99470, 99440, 99420, 99440, 99430, 99430, 99390, 99410, 99400, 99400, 
    99390, 99420, 99420, 99410, 99400, 99370, 99360, 99340, 99290, 99310, 
    99330, 99350, 99370, 99360, 99390, 99370, 99360, 99350, 99310, 99260, 
    99230, 99180, 99130, 99120, 99090, 99080, 99040, 99010, 98970, 98940, 
    98920, 98920, 98900, 98880, 98900, 98930, 98940, 98990, 99060, 99100, 
    99130, 99180, 99230, 99280, 99330, 99390, 99420, 99480, 99530, 99580, 
    99640, 99730, 99790, 99860, 99920, 99990, 100040, 100120, 100180, 100240, 
    100320, 100400, 100460, 100530, 100580, 100630, 100680, 100730, 100790, 
    100850, 100880, 100940, 101010, 101070, 101120, 101160, 101200, 101250, 
    101290, 101340, 101360, 101390, 101400, 101430, 101450, 101450, 101470, 
    101490, 101490, 101470, 101450, 101400, 101360, 101300, 101230, 101160, 
    101070, 100940, 100820, 100700, 100590, 100460, 100300, 100080, 99900, 
    99690, 99590, 99530, 99480, 99440, 99400, 99370, 99350, 99350, 99290, 
    99240, 99190, 99140, 99080, 99050, 99010, 98990, 98960, 98980, 99000, 
    99050, 99080, 99130, 99150, 99160, 99200, 99220, 99230, 99250, 99250, 
    99230, 99210, 99200, 99260, 99310, 99420, 99500, 99540, 99570, 99660, 
    99700, 99770, 99780, 99800, 99800, 99830, 99860, 99880, 99910, 99940, 
    100000, 100040, 100080, 100150, 100200, 100250, 100320, 100380, 100450, 
    100550, 100620, 100670, 100750, 100840, 100880, 100940, 101040, 101070, 
    101120, 101160, 101190, 101190, 101260, 101300, 101340, 101370, 101400, 
    101410, 101400, 101400, 101390, 101330, 101300, 101260, 101220, 101140, 
    101130, 101080, 101060, 101090, 101070, 101050, 101000, 101050, 101060, 
    101050, 101040, 101040, 100990, 100930, 100870, _, 100680, 100580, 
    100460, 100360, 100300, 100180, 100120, 100080, 99960, 99860, 99740, 
    99620, 99460, 99280, 99200, 99180, 99180, 99190, 99170, 99170, 99230, 
    99270, 99360, 99440, 99510, 99590, 99610, 99680, 99720, 99740, 99810, 
    99890, 99940, 100020, 100150, 100250, 100360, 100430, 100550, 100630, 
    100750, 100850, 100920, 101000, 101080, 101160, 101240, 101300, 101350, 
    101390, 101440, 101460, 101490, 101510, 101540, 101550, 101580, 101600, 
    101630, 101650, 101670, 101680, 101690, 101710, 101720, 101760, 101770, 
    101770, 101780, 101800, 101820, 101850, 101890, 101900, 101940, 101940, 
    101970, 101990, 101980, 101960, 101980, 102000, 102010, 102020, 102060, 
    102070, 102090, 102070, 102080, 102080, 102080, 102110, 102100, 102140, 
    102190, 102210, 102230, 102240, 102270, 102280, 102290, 102280, 102290, 
    102290, 102260, 102240, 102230, 102210, 102200, 102180, 102170, 102140, 
    102110, 102060, 102030, 101980, 101940, 101920, 101900, 101870, 101830, 
    101790, 101740, 101690, 101600, 101540, 101490, 101420, 101320, 101230, 
    101150, 101050, 100950, 100810, 100740, 100640, 100560, 100450, 100360, 
    100290, 100240, 100180, 100150, 100150, 100170, 100180, 100180, 100180, 
    100180, 100180, 100170, 100180, 100200, 100210, 100230, 100220, 100230, 
    100230, 100210, 100180, 100160, 100130, 100090, 100090, 100090, 100080, 
    100090, 100080, 100090, 100080, 100050, 100010, 99970, 99990, 99970, 
    99980, 99960, 99930, 99920, 99860, 99850, 99890, 99910, 100000, 100070, 
    100160, 100230, 100280, 100330, 100380, 100440, 100490, 100540, 100610, 
    100640, 100690, 100770, 100820, 100880, 100940, 100990, 101060, 101130, 
    101210, 101280, 101310, 101320, 101360, 101370, 101400, 101420, 101440, 
    101440, 101470, 101500, 101500, 101500, 101500, 101470, 101460, 101440, 
    101430, 101380, 101320, 101270, 101220, 101190, 101120, 101040, 100970, 
    100900, 100810, 100700, 100620, 100530, 100430, 100320, 100200, 100120, 
    100000, 99850, 99790, 99690, 99560, 99480, 99430, 99390, 99360, 99340, 
    99370, 99400, 99450, 99480, 99540, 99600, 99660, 99730, 99810, 99930, 
    100060, 100150, 100230, 100360, 100470, 100570, 100660, 100760, 100910, 
    101000, 101030, 101090, 101160, 101220, 101270, 101340, 101380, 101370, 
    101380, 101400, 101410, 101430, 101390, 101390, 101370, 101360, 101360, 
    101350, 101350, 101340, 101310, 101300, 101280, 101280, 101260, 101270, 
    101330, 101360, 101400, 101430, 101450, 101470, 101500, 101560, 101590, 
    101630, 101600, 101610, 101630, 101650, 101710, 101770, 101850, 101900, 
    101960, 101990, 101990, 102010, 102010, 102020, 102040, 102070, 102070, 
    102080, 102090, 102100, 102100, 102070, 102040, 102030, 102040, 102020, 
    101970, 101950, 101920, 101860, 101810, 101790, 101740, 101660, 101640, 
    101570, 101490, 101440, 101390, 101320, 101270, 101240, 101210, 101180, 
    101160, 101130, 101100, 101070, 101060, 101060, 101060, 101050, 101050, 
    101030, 101010, 100980, 100970, 100950, 100910, 100900, 100890, 100880, 
    100870, 100850, 100840, 100810, 100770, 100770, 100770, 100750, 100750, 
    100780, 100790, 100780, 100760, 100750, 100750, 100750, 100740, 100740, 
    100730, 100720, 100730, 100750, 100730, 100710, 100690, 100680, 100670, 
    100660, 100660, 100640, 100630, 100620, 100630, 100600, 100580, 100560, 
    100550, 100560, 100570, 100560, 100570, 100580, 100580, 100580, 100550, 
    100530, 100520, 100510, 100500, 100490, 100500, 100500, 100500, 100500, 
    100480, 100470, 100480, 100480, 100470, 100460, 100470, 100470, 100470, 
    100470, 100490, 100490, 100500, 100490, 100490, 100490, 100490, 100480, 
    100460, 100450, 100450, 100450, 100460, 100450, 100450, 100450, 100440, 
    100440, 100440, 100440, 100440, 100440, 100470, 100500, 100510, 100520, 
    100510, 100490, 100510, 100500, 100470, 100480, 100480, 100470, 100460, 
    100440, 100410, 100400, 100390, 100370, 100350, 100320, 100280, 100240, 
    100210, 100200, 100190, 100180, 100170, 100150, 100110, 100090, 100080, 
    100060, 100050, 100030, 100030, 100030, 100040, 100050, 100050, 100040, 
    100040, 100040, 100040, 100070, 100060, 100020, 99960, 99940, 99950, 
    99960, 99970, 99970, 99980, 99980, 100000, 100040, 100040, 100040, 
    100050, 100080, 100100, 100150, 100180, 100200, 100210, 100190, 100200, 
    100220, 100220, 100190, 100180, 100210, 100220, 100250, 100280, 100310, 
    100350, 100340, 100370, 100360, 100340, 100350, 100330, 100320, 100320, 
    100320, 100320, 100320, 100320, 100340, 100340, 100330, 100310, 100320, 
    100310, 100310, 100280, 100280, 100230, 100210, 100200, 100180, 100150, 
    100140, 100130, 100120, 100120, 100080, 100090, 100090, 100090, 100070, 
    100050, 100060, 100080, 100080, 100040, 100050, 100050, 100060, 100090, 
    100110, 100120, 100130, 100150, 100140, 100160, 100170, 100170, 100150, 
    100170, 100160, 100170, 100190, 100210, 100200, 100190, 100190, 100180, 
    100170, 100150, 100140, 100150, 100140, 100140, 100120, 100110, 100110, 
    100090, 100080, 100090, 100090, 100090, 100080, 100090, 100100, 100100, 
    100130, 100180, 100220, 100260, 100280, 100320, 100370, 100420, 100450, 
    100490, 100540, 100590, 100650, 100690, 100720, 100760, 100790, 100820, 
    100860, 100930, 100980, 101030, 101070, 101120, 101170, 101220, 101230, 
    101270, 101300, 101330, 101370, 101410, 101430, 101450, 101450, 101490, 
    101490, 101510, 101490, 101490, 101460, 101450, 101460, 101450, 101460, 
    101450, 101430, 101420, 101420, 101400, 101390, 101370, 101360, 101340, 
    101310, 101290, 101270, 101250, 101260, 101260, 101260, 101260, 101270, 
    101270, 101280, 101280, 101290, 101280, 101260, 101250, 101220, 101210, 
    101210, 101210, 101230, 101240, 101240, 101220, 101200, 101160, 101160, 
    101170, 101110, 101120, 101130, 101100, 101130, 101120, 101110, 101100, 
    101090, 101070, 101070, 101060, 101050, 101050, 101050, 101030, 101020, 
    101020, 101000, 100980, 100950, 100910, 100880, 100860, 100870, 100870, 
    100860, 100840, 100800, 100790, 100790, 100810, 100850, 100900, 100950, 
    100970, 101020, 101060, 101120, 101160, 101210, 101250, 101330, 101400, 
    101450, 101490, 101510, 101500, 101520, 101520, 101500, 101530, 101460, 
    101400, 101310, 101210, 101080, 100990, 100960, 101000, 101030, 101040, 
    101130, 101220, 101300, 101370, 101470, 101550, 101610, _, 101740, 
    101780, 101820, 101860, 101890, 101920, 101920, 101940, 101930, 101920, 
    101930, 101930, 101930, 101910, 101930, 101940, 101980, 102010, 102020, 
    102040, 102080, 102160, 102200, 102220, 102220, 102240, 102290, 102330, 
    102400, 102440, 102460, 102500, 102500, 102510, 102500, 102510, 102500, 
    102500, 102500, 102470, 102470, 102440, 102380, 102330, 102270, 102200, 
    102180, 102150, 102120, 102120, 102100, 102070, 102100, 102110, 102100, 
    102100, 102060, 102030, 102010, 101970, 101920, 101880, 101830, 101760, 
    101710, 101660, 101620, 101520, 101440, 101370, 101280, 101210, 101140, 
    101070, 101030, 100990, 100960, 100910, 100860, 100810, 100770, 100740, 
    100710, 100670, 100660, 100660, 100650, 100680, 100710, 100760, _, 
    100810, 100800, 100810, 100810, 100820, 100820, 100880, 100930, 101010, 
    101120, 101220, 101360, 101430, 101510, 101570, 101640, 101700, 101720, 
    101770, 101810, 101890, 101940, 101970, 101990, 101980, 101980, 102010, 
    102040, 102060, 102070, 102070, 102050, 102070, 102090, 102120, 102130, 
    102110, 102070, 102020, 101920, 101860, 101840, 101850, 101850, 101830, 
    101800, 101780, 101740, 101680, 101640, 101620, 101610, 101580, 101550, 
    101540, 101530, 101530, 101520, 101520, 101490, 101470, 101470, 101450, 
    101450, 101480, 101500, 101510, 101550, 101610, 101640, 101700, 101750, 
    101790, 101830, 101850, 101850, 101890, 101930, 101980, 102030, 102090, 
    102140, 102190, 102230, 102240, 102260, 102290, 102290, 102300, 102290, 
    102270, 102260, 102240, 102210, 102190, 102170, 102110, 102120, 102100, 
    102080, 102100, 102100, 102120, 102140, 102160, 102190, 102200, 102190, 
    102190, 102190, 102190, 102140, 102120, 102070, 102060, 102050, 102020, 
    101990, 101940, 101910, 101840, 101760, 101730, 101680, 101610, 101530, 
    101440, 101360, 101320, 101250, 101190, 101120, 101070, 101050, 101050, 
    101090, 101140, 101220, 101300, 101380, 101460, 101560, 101630, 101710, 
    101790, 101830, 101980, 101940, 101980, 102020, 102090, 102150, 102220, 
    102260, 102310, 102360, 102390, 102430, 102470, 102510, 102530, 102530, 
    102560, 102580, 102580, 102560, 102560, 102500, 102420, 102340, 102310, 
    102300, 102240, 102150, 102050, 101960, 101870, 101790, 101750, 101710, 
    101690, 101710, 101680, 101670, 101690, 101700, 101730, 101750, 101770, 
    101790, 101840, 101860, 101870, 101920, 101960, 101970, 101990, 102000, 
    102020, 102020, 102020, 102020, 102030, 102040, 102030, 102000, 101960, 
    101950, 101920, 101880, 101810, 101780, 101770, 101770, 101720, 101700, 
    101670, 101670, 101670, 101650, 101660, 101670, 101680, 101710, 101750, 
    101810, 101840, 101880, 101910, 101930, 101940, 101940, 101940, 101920, 
    101900, 101890, 101860, 101810, 101780, 101720, 101670, 101590, 101500, 
    101410, 101310, 101190, 101090, 100980, 100860, 100790, 100770, 100690, 
    100610, 100540, 100520, 100500, 100510, 100520, 100500, 100500, 100530, 
    100570, 100660, 100730, 100790, 100840, 100870, 100940, 101020, 101120, 
    101210, 101290, 101400, 101490, 101580, 101670, 101750, 101820, 101910, 
    101960, 102010, 102070, 102080, 102110, 102130, 102140, 102140, 102120, 
    102110, 102070, 102000, 101930, 101870, 101790, 101770, 101730, 101690, 
    101690, 101720, 101700, 101700, 101690, 101670, 101690, 101690, 101720, 
    101740, 101780, 101830, 101860, 101890, 101890, 101910, 101890, 101890, 
    101890, 101910, 101900, 101890, 101900, 101920, 101950, 101990, 101980, 
    101990, 101990, 102000, 102020, 102010, 101980, 101950, 101930, 101940, 
    101940, 101900, 101880, 101880, _, 101830, 101810, 101780, 101760, 
    101740, 101740, 101710, 101710, 101690, 101670, 101640, 101670, 101640, 
    101620, 101620, 101590, 101540, 101500, 101460, 101460, 101450, 101430, 
    101410, 101380, 101370, 101360, _, 101350, 101350, 101340, 101350, 
    101390, 101410, 101420, 101450, 101450, 101440, 101450, 101460, 101470, 
    101480, 101490, 101510, 101530, 101540, 101570, 101580, 101570, 101570, 
    101590, 101590, 101570, 101550, 101540, 101550, 101570, 101600, 101610, 
    101640, 101660, 101710, 101720, 101750, 101760, 101790, 101810, 101810, 
    101840, 101840, 101830, 101830, _, 101780, 101760, 101750, 101730, 
    101740, 101740, 101780, 101800, 101830, 101830, 101830, 101830, 101830, 
    101840, 101840, 101840, 101820, 101800, 101780, 101730, 101700, 101680, 
    101680, 101700, 101650, 101730, 101770, 101910, 102010, 101990, 102050, 
    102100, 102190, 102190, 102210, 102280, 102370, 102440, 102480, 102520, 
    102600, 102670, 102690, 102730, 102790, 102780, 102810, 102780, 102820, 
    102820, 102770, 102740, 102710, 102710, 102730, 102760, 102770, 102750, 
    102720, 102690, 102660, 102640, 102610, 102600, 102580, 102560, 102530, 
    102530, 102510, 102480, 102430, 102400, _, 102330, 102320, 102300, 
    102280, 102300, 102320, 102330, 102330, 102360, 102400, 102410, 102440, 
    102450, 102500, 102520, 102560, 102600, 102650, 102680, 102710, 102770, 
    102810, 102810, 102850, 102870, 102890, 102900, 102910, 102940, 102940, 
    102960, 102980, 102970, 102950, 102920, 102880, 102820, 102790, 102720, 
    102660, 102620, 102580, 102550, 102500, 102480, 102480, 102450, 102440, 
    102410, 102380, 102340, 102330, 102270, 102250, 102260, 102230, 102190, 
    102220, 102190, 102180, 102130, 102110, 102110, 102160, 102160, 102170, 
    102150, 102120, 102090, 102080, 102070, 102050, 102020, 101970, 101960, 
    101930, 101950, 101970, 101970, 101960, 101990, 102050, 102110, 102160, 
    102210, 102240, 102260, 102260, 102280, 102310, 102350, 102360, 102370, 
    102380, _, _, 102420, _, 102430, _, _, _, _, _, 102480, 102480, 102460, 
    102440, 102410, _, 102380, 102350, 102280, 102270, 102220, 102220, 
    102180, 102110, _, 102120, 102150, 102110, 102100, 102080, 102080, 
    102090, 102090, 102130, 102130, 102140, 102110, 102090, 102090, 102090, 
    102050, 102050, 102010, 101970, 101960, 101940, 101900, 101850, 101810, 
    101770, 101720, 101670, 101600, 101540, 101490, 101450, 101400, 101350, 
    101320, 101270, 101210, 101160, 101120, 101090, 101030, 101000, 100940, 
    100920, 100900, 100870, 100830, 100790, 100750, 100720, 100680, _, 
    100580, 100540, 100490, 100470, 100440, _, 100340, 100310, 100270, 
    100240, 100210, 100200, 100210, 100220, 100250, 100260, 100250, 100240, 
    100280, 100360, _, 100420, 100430, 100460, 100460, 100490, 100550, 
    100620, 100680, 100730, 100770, 100800, 100810, 100820, 100830, 100830, 
    100850, 100870, 100900, 100940, 100970, 100990, 100990, 100980, _, 
    100980, 101010, 101070, 101110, 101140, 101190, 101220, 101280, 101330, 
    101390, 101460, 101520, 101600, 101650, 101720, 101770, 101850, 101970, 
    102080, 102180, 102290, 102340, 102410, 102480, 102540, 102580, _, 
    102690, 102750, 102810, 102880, 102930, 102960, 102980, 103020, 103060, 
    103090, 103130, 103140, 103170, 103200, 103250, 103310, 103400, 103450, 
    103520, 103580, _, 103680, 103760, 103810, 103900, 103980, 104060, 
    104130, 104190, 104280, 104300, 104360, 104450, 104490, 104500, 104540, 
    104570, 104600, 104610, 104630, 104680, 104750, 104780, 104840, _, 
    104980, 105010, 105050, 105090, 105120, 105140, 105160, 105160, 105150, 
    105140, 105130, 105140, 105150, 105180, 105170, 105170, 105180, 105230, 
    105280, 105310, 105340, 105360, 105370, 105370, 105420, 105430, 105450, 
    105440, 105450, 105460, 105490, 105540, 105570, 105580, 105590, 105590, 
    105590, 105590, 105560, 105550, 105550, 105550, 105540, 105520, 105520, 
    105500, 105470, _, 105420, 105390, 105370, 105310, 105310, 105290, 
    105260, 105230, 105190, 105160, 105120, 105080, 105020, 104960, 104920, 
    104870, 104800, 104750, 104730, 104680, 104660, 104610, 104540, _, _, 
    104320, 104240, 104190, 104120, 104060, 104010, 103950, 103890, 103830, 
    103750, 103690, 103640, 103620, 103560, 103560, 103490, 103460, 103460, 
    103440, 103400, 103360, 103320, 103310, 103290, 103240, 103250, 103210, 
    103160, 103180, 103210, 103240, 103240, 103260, 103240, 103210, 103190, 
    103160, 103160, 103140, _, 103070, 102980, 102960, 102940, 102890, 
    102850, _, 102750, 102740, 102720, 102710, 102730, 102740, 102760, 
    102790, 102810, 102830, 102830, 102820, 102830, 102860, 102880, 102890, 
    102880, 102900, 102930, 102950, 102950, 102920, _, _, _, 102880, 102870, 
    102850, 102820, 102810, 102810, 102790, 102790, 102750, 102730, 102700, 
    102660, 102640, 102600, 102560, 102520, 102490, 102490, 102480, 102460, 
    102430, 102380, 102350, 102340, 102300, 102290, _, _, 102190, 102170, 
    102120, 102100, 102060, 102020, 101970, 101920, 101860, 101810, 101760, 
    101730, 101670, 101610, 101570, 101490, 101420, 101330, _, 101170, 
    101070, 101050, 100980, 100980, 101010, 101060, 101010, 101060, 101100, 
    101140, 101150, 101160, 101100, 101190, 101220, 101190, 101170, 101180, 
    101130, 101070, 101070, 101040, 101070, 101080, 101120, 101160, 101220, 
    101250, 101310, 101370, 101420, 101480, 101520, 101550, 101600, 101620, 
    101640, 101660, 101680, 101690, 101700, 101720, 101710, 101710, 101690, 
    101670, 101660, 101650, 101610, 101610, 101610, 101590, 101560, 101550, 
    101540, 101530, 101510, 101480, 101450, 101410, 101400, 101370, 101330, 
    101310, 101300, 101260, 101240, 101220, 101210, 101210, 101170, 101130, 
    101090, 101060, 101020, 100990, 100950, 100930, 100900, 100860, 100860, 
    100830, 100780, 100750, 100720, 100690, 100650, 100610, 100550, 100510, 
    100470, 100450, 100420, 100380, 100340, 100300, 100250, 100220, 100200, 
    100140, 100110, 100110, 100100, 100090, 100060, 100060, 100040, 100040, 
    _, 100060, 100060, 100040, 100040, 100040, 100040, 100050, 100060, 
    100070, 100070, 100080, 100080, 100070, 100090, 100100, 100120, 100160, 
    100180, 100210, 100240, 100290, 100310, 100320, 100350, 100370, 100400, 
    100450, 100500, 100540, 100590, 100640, 100680, 100720, 100950, 100780, 
    100810, 100870, 100890, 100930, 100980, 101020, 101080, 101120, 101140, 
    101170, 101220, 101230, 101240, 101260, 101280, 101280, 101300, 101330, 
    101360, 101350, 101360, 101440, 101400, 101410, 101400, 101410, 101410, 
    101410, 101440, 101450, 101470, 101510, 101530, 101540, 101550, 101560, 
    101570, 101590, 101630, 101650, 101680, 101710, 101770, 101810, 101820, 
    101850, 101860, 101880, 101900, 101930, 101970, 102000, 102010, 102030, 
    102060, 102060, 102070, 102130, 102140, 102150, 102140, 102130, 102080, 
    102150, 102210, 102200, 102250, 102290, 102310, 102300, _, 102380, 
    102400, 102390, 102400, 102400, 102400, 102380, 102430, 102420, 102410, 
    102380, 102340, 102320, 102310, 102320, 102450, 102540, 102610, 102650, 
    102670, 102680, 102680, 102660, 102640, 102620, 102580, 102500, 102470, 
    102430, 102410, 102350, 102300, 102240, 102180, 102090, 102010, 101940, 
    101850, 101760, 101690, 101650, 101600, 101570, 101590, 101570, 101560, 
    101560, 101570, 101580, 101570, 101570, 101590, 101630, 101690, 101720, 
    101740, 101740, 101750, 101740, 101700, 101690, 101650, 101630, 101580, 
    101540, 101530, 101520, 101490, 101440, 101420, 101380, _, 101350, 
    101310, 101250, _, 101150, 101120, 101100, 101060, 101030, 101000, 
    100970, 100940, 100930, 100910, 100890, 100890, 100850, 100860, 100870, 
    100880, 100910, _, 100920, 100930, 100930, 100920, 100940, 100940, 
    100950, 100950, 100970, 100980, 100980, 100970, 100970, 100970, 100970, 
    100950, 100940, 100930, 100940, 100950, 100960, 100970, 100950, 100950, 
    100940, 100910, 100910, 100900, 100910, 100910, 100900, 100900, 100910, 
    100920, 100910, 100910, 100910, 100920, 100930, 100910, 100890, 100900, 
    100920, 100960, 100990, 101020, 101010, 101000, 101030, 101030, 101050, 
    101020, 101060, 101090, 101110, 101140, 101160, 101200, 101250, 101280, 
    101290, 101310, 101350, 101380, 101380, 101390, 101440, 101470, 101510, 
    101520, 101520, 101510, 101510, 101510, 101530, 101540, 101520, 101490, 
    101470, 101480, 101470, 101460, 101440, 101410, 101390, 101370, 101370, 
    101360, 101320, 101310, 101300, 101300, 101300, _, 101310, _, 101300, 
    101290, 101290, 101270, 101270, 101250, 101250, 101270, 101290, 101290, 
    101280, 101270, 101240, 101220, 101220, 101200, 101190, 101180, 101160, 
    101130, 101130, 101120, 101100, 101080, 101070, 101050, 101040, 101020, 
    101010, 100990, 100970, 100960, 100960, 100940, 100940, 100940, 100920, 
    100910, 100900, 100900, 100870, 100870, 100850, 100860, 100850, 100850, 
    100840, 100820, 100820, 100810, 100800, 100820, 100810, 100800, 100800, 
    100800, 100800, 100810, 100820, 100830, 100830, 100840, 100870, 100890, 
    100900, 100930, 100940, 100950, 100970, 100980, 101000, 101030, 101050, 
    101040, 101040, 101060, 101040, 101030, 101050, 101050, 101060, 101030, 
    101030, 101000, 100980, 100970, 100930, 100880, 100840, 100790, 100750, 
    100710, 100660, 100630, 100580, 100540, 100490, 100450, 100410, 100350, 
    100310, 100280, 100240, 100230, 100210, 100190, 100190, 100170, 100170, 
    100170, 100170, 100170, 100200, 100180, 100210, 100220, 100250, 100250, 
    100280, 100300, 100330, 100350, 100360, 100360, 100340, 100320, 100340, 
    100350, 100350, 100340, 100340, 100340, 100370, 100350, 100350, 100330, 
    100330, _, 100330, 100330, 100340, _, 100310, 100300, 100300, 100300, 
    100270, 100250, 100240, 100250, 100260, 100280, 100320, 100340, 100340, 
    100380, 100390, 100420, 100440, 100500, 100540, 100560, _, _, _, 100740, 
    100770, 100800, 100850, 100900, 100940, 100970, 101020, 101080, 101110, 
    101150, 101210, 101260, 101300, 101340, 101380, 101400, 101450, 101450, 
    101470, 101510, 101530, 101540, _, 101600, 101620, 101610, 101620, 
    101620, 101610, 101610, 101600, 101580, 101570, 101560, 101540, 101490, 
    101450, 101410, 101380, 101340, 101300, 101220, 101110, 101030, 100950, 
    100830, 100680, 100540, 100330, _, _, 99870, 99690, 99590, 99510, 99470, 
    99460, 99450, 99460, 99480, 99520, _, 99520, 99490, 99470, 99430, 99390, 
    99360, 99320, 99270, 99220, 99170, 99140, 99100, 99050, 99030, 99010, 
    99000, 98990, 98990, 98990, _, 99010, 99030, 99070, 99090, 99110, 99130, 
    99160, 99140, 99150, 99160, 99170, 99200, _, 99190, 99190, 99180, 99140, 
    99120, 99070, 99080, 99040, 99010, 98990, 98940, 98930, 98900, 98880, 
    98880, 98890, 98890, 98910, 98930, 98940, 98970, 99010, 99040, 99070, 
    99110, 99150, _, 99210, 99230, 99270, 99300, 99330, 99380, 99410, 99440, 
    99460, 99480, 99500, 99530, 99560, 99590, 99600, 99630, 99660, 99710, 
    99740, 99780, 99820, 99840, 99870, 99890, 99920, 99940, 99940, 99950, 
    99970, 99980, 100010, 100020, 100010, 100010, 100000, 99980, 99960, 
    99960, 99960, 99960, 99960, 99980, 100010, 100030, 100060, 100080, 
    100130, 100150, 100180, 100220, 100230, 100260, 100290, 100330, 100360, 
    100420, 100450, 100490, 100540, 100610, 100660, 100700, 100740, 100780, 
    100820, 100840, 100880, 100920, 100960, 100990, 101000, 101030, 101060, 
    101060, 101060, 101050, 101030, 101010, 101000, 100980, 100990, 100980, 
    100950, 100940, 100920, 100930, 100890, 100850, 100820, 100780, 100740, 
    100680, 100630, 100610, 100580, 100520, 100510, 100480, 100450, 100440, 
    100430, 100400, 100410, 100420, 100430, 100430, 100460, 100490, 100510, 
    100550, 100560, 100590, 100580, 100600, 100630, 100640, 100660, 100690, 
    100700, 100720, 100730, 100720, 100720, 100750, 100750, 100750, 100740, 
    100770, 100800, 100820, 100830, 100860, 100880, 100900, 100920, 100910, 
    100910, 100930, 100960, _, 101000, 101030, 101060, _, 101060, 101060, 
    101070, 101090, 101080, 101090, 101110, 101100, 101120, 101150, 101150, 
    101140, 101130, 101100, 101100, 101070, _, 101050, 101020, 101010, 
    100990, 100980, 100950, 100930, 100910, 100880, 100860, 100830, 100810, 
    100800, 100820, 100820, 100820, 100810, 100790, 100770, 100760, 100750, 
    100730, 100710, 100670, 100640, 100580, 100580, 100550, 100500, 100500, 
    100460, 100420, 100390, 100370, 100330, 100320, 100340, 100340, 100340, 
    100360, 100390, 100400, 100410, 100430, 100440, 100470, 100490, 100490, 
    100510, 100530, 100530, 100580, 100620, 100650, 100690, 100730, 100750, 
    100780, 100800, 100840, 100870, 100880, 100910, 100960, 101010, 101030, 
    101040, 101070, 101080, 101090, 101120, 101120, 101110, 101160, 101190, 
    101200, 101240, 101270, 101280, 101290, 101300, 101280, 101280, 101280, 
    101280, 101290, 101310, 101330, 101330, 101350, 101380, 101380, 101420, 
    101450, 101450, 101450, 101460, 101460, 101480, 101490, 101510, 101530, 
    101510, 101500, 101460, 101440, 101420, 101410, 101390, 101350, 101330, 
    101310, 101300, 101290, 101260, 101230, 101200, 101160, 101100, 101060, 
    101030, 100990, 100970, 100950, 100910, 100870, 100830, 100810, 100780, 
    100760, 100730, 100690, 100630, 100600, 100550, 100530, 100480, 100460, 
    100430, 100420, 100410, 100390, 100380, 100390, 100390, 100420, 100450, 
    _, 100510, 100530, 100560, 100590, 100620, 100640, 100670, 100700, 
    100730, 100800, 100830, 100890, 100930, 100970, 101030, 101050, 101090, 
    101120, 101140, 101170, 101180, 101230, 101270, 101310, 101350, 101390, 
    101400, 101430, 101470, 101470, 101460, 101480, 101490, 101500, 101500, 
    _, 101500, 101490, 101490, 101470, 101460, 101430, 101420, 101400, 
    101370, 101360, 101330, 101330, 101320, 101300, 101270, 101250, 101200, 
    101150, 101120, 101010, 100990, 100920, 100890, 100860, 100850, 100850, 
    100840, 100850, 100860, 100840, 100830, 100820, 100820, 100820, 100850, 
    _, 100890, 100930, 100950, 100980, 100990, 101010, 101020, 101060, _, _, 
    _, 101200, 101250, 101300, 101340, 101370, 101420, 101470, 101510, 
    101530, 101570, 101620, 101670, _, 101770, 101800, 101810, 101850, 
    101880, 101890, 101910, 101930, 101950, 101980, 102020, 102040, 102060, 
    102070, 102120, 102150, 102170, 102200, 102210, 102260, 102280, 102300, 
    102350, 102390, 102450, 102480, 102520, 102540, 102580, 102610, 102650, 
    102670, 102690, 102720, 102750, 102770, 102800, 102830, 102830, 102830, 
    102840, 102840, 102830, 102830, 102810, 102830, 102830, _, 102830, 
    102820, 102800, 102790, 102760, 102730, 102700, 102680, 102680, 102660, 
    102650, 102650, 102630, 102620, 102600, 102590, 102570, 102560, 102540, 
    102500, 102490, 102470, 102460, _, 102460, 102450, 102420, 102390, 
    102370, 102350, 102320, 102300, 102300, 102310, 102320, 102310, 102300, 
    102290, 102300, 102310, 102290, 102310, 102310, 102300, 102320, 102350, 
    102380, 102410, 102440, 102460, 102480, 102510, 102540, 102590, 102630, 
    102660, 102690, 102730, 102770, 102810, 102840, 102880, 102910, 102930, 
    102920, 102940, 102960, 102980, 102980, 102990, 102980, _, 102970, 
    103000, 102980, 102920, 102920, 102890, 102820, 102750, 102720, 102680, 
    102630, 102600, 102530, 102440, 102410, 102300, 102140, 102050, 101940, 
    101800, 101680, 101580, 101470, _, 101300, 101220, 101140, 101070, 
    101020, 100940, 100880, 100850, 100830, 100840, 100860, 100870, 100930, 
    100980, 101040, 101070, 101150, 101210, 101260, 101320, 101350, 101410, 
    101460, 101540, 101620, 101700, 101780, 101870, 101930, 102000, 102060, 
    102130, 102170, 102210, 102230, 102300, 102360, 102400, 102440, 102430, 
    102450, 102470, 102460, 102450, 102440, 102430, 102430, _, 102400, 
    102390, 102390, 102360, 102360, 102320, 102290, 102250, 102220, 102200, 
    102200, 102200, 102210, 102220, 102210, 102210, 102190, 102170, 102130, 
    102110, 102090, _, 102020, _, 102020, 102000, 101970, 101940, 101910, 
    101870, 101860, 101840, 101810, 101790, 101810, 101800, 101820, 101830, 
    101830, 101820, 101800, 101800, 101810, 101830, 101870, 101880, 101910, 
    101970, 101990, 102030, 102030, 102050, 102040, 102070, 102070, 102070, 
    102070, 102100, 102100, 102130, 102150, 102170, 102190, 102170, 102180, 
    102190, 102210, 102220, 102200, 102200, 102230, _, 102260, 102240, 
    102210, 102190, 102130, 102090, 102030, 102010, 101950, 101920, 101880, 
    101840, 101790, 101750, 101710, 101630, 101560, 101470, 101360, 101270, 
    101180, _, 101020, _, _, 100820, 100760, 100670, 100630, 100550, 100450, 
    100350, 100290, 100220, 100140, 100090, 100070, 100040, 100000, 99970, 
    99930, 99960, 99970, 99990, 100020, 100030, 100100, 100170, 100240, 
    100300, 100430, 100520, 100610, 100690, 100760, 100820, 100890, 100990, 
    101090, 101190, 101280, 101370, 101450, 101520, 101600, 101670, 101730, 
    101790, 101850, 101920, 101970, _, 102010, 102040, 102070, 102090, 
    102070, 102090, 102070, 102050, 102030, 102050, 102040, 102030, 102040, 
    102030, 102020, _, 102010, 101980, 101950, 101950, _, _, 101890, _, 
    101870, 101860, 101850, 101830, 101780, 101770, 101740, 101710, 101680, 
    101670, 101660, 101640, 101650, 101660, 101670, 101670, 101650, 101620, 
    101610, 101610, 101610, 101610, 101640, 101680, 101730, 101780, 101860, 
    101930, 101950, 102000, 102030, 102060, 102120, 102170, 102210, 102250, 
    102290, 102330, 102370, 102380, 102380, 102390, 102410, 102430, 102410, 
    102400, 102410, _, 102340, 102280, 102220, 102100, 102030, 102010, 
    101960, 101910, 101920, 101970, 102010, 102050, _, 102150, 102180, 
    102200, 102250, 102270, 102250, 102210, 102190, 102170, 102170, 102170, 
    102160, 102130, 102100, 102060, 102020, 101960, 101930, 101880, 101820, 
    101770, 101720, 101680, 101640, _, _, 101580, 101520, 101500, 101470, 
    101440, 101420, 101440, 101420, 101420, 101430, 101440, 101450, 101480, 
    101460, 101490, 101500, 101520, 101530, 101570, 101620, 101670, 101700, 
    101740, 101760, 101800, 101830, 101850, 101880, 101910, 101950, 101970, 
    102010, _, 102080, 102130, 102140, _, 102200, 102230, 102250, 102270, 
    102290, 102320, 102350, _, 102410, 102440, 102440, 102450, 102430, 
    102430, 102410, 102420, 102420, _, 102410, 102420, 102430, 102420, 
    102420, 102410, 102380, 102370, 102330, 102290, 102250, 102210, 102200, 
    102230, 102220, 102160, 102140, 102110, 102060, 102010, 102000, _, 
    101900, 101880, 101840, 101830, 101790, 101720, 101660, 101580, 101510, 
    101490, 101400, 101330, 101310, 101270, 101300, 101300, 101310, 101310, 
    101300, 101260, 101210, 101100, 101020, 100940, 100910, 100890, 100860, 
    _, 100940, 101000, 101020, 101060, 101060, 101150, 101170, 101260, 
    101310, 101340, 101420, 101460, 101530, 101570, 101590, 101590, 101610, 
    101660, 101710, 101720, 101780, _, _, _, 101850, 101840, 101790, 101720, 
    101630, 101570, 101520, 101460, 101430, 101410, 101340, 101300, 101310, 
    101320, 101280, 101270, 101220, 101180, _, _, 101140, _, 101140, 101150, 
    101180, 101170, 101170, 101150, 101150, 101160, 101160, 101180, 101190, 
    101210, 101270, 101280, 101290, 101300, 101280, 101320, 101290, 101280, 
    101300, 101270, 101230, 101190, 101150, 101150, 101080, 101010, 100940, 
    100860, 100780, 100680, 100630, 100600, 100550, 100600, 100640, 100690, 
    100760, 100890, 101000, 101080, 101170, 101230, 101310, 101340, 101370, 
    _, 101410, 101450, 101480, 101510, 101520, 101530, 101540, 101540, 
    101530, 101530, 101520, 101540, 101520, 101520, 101550, 101530, 101520, 
    101480, 101450, _, 101400, _, 101300, _, 101200, 101170, 101140, 101070, 
    101010, 100960, 100890, 100820, 100760, 100700, 100640, 100630, 100620, 
    100610, 100600, 100600, 100620, 100650, _, 100670, 100680, 100700, 
    100710, 100720, 100780, 100820, 100870, 100920, 100960, 100970, 100970, 
    101000, 101010, 100990, 101010, 101020, 101020, 101000, 101030, 101030, 
    101010, 101010, 101010, 101040, 101060, 101080, 101060, 101110, 101130, 
    101160, 101180, 101220, 101240, 101260, 101280, 101290, 101290, 101300, 
    101300, 101300, 101310, 101320, 101330, 101340, 101330, 101320, 101280, 
    101250, 101200, _, 101100, _, 101050, 101030, 101010, 100970, 100940, 
    100880, 100840, 100780, 100750, 100710, 100670, 100670, 100660, 100660, 
    100670, _, 100670, 100650, 100640, 100650, 100680, 100690, 100720, 
    100730, 100740, 100780, 100790, 100800, 100810, 100810, 100790, 100760, 
    100750, 100720, 100700, 100680, 100660, 100650, 100610, 100600, 100530, 
    100490, 100470, 100460, 100420, 100390, 100350, 100280, 100230, 100240, 
    100220, 100190, 100140, 100110, 100100, 100060, 100020, 99970, 99950, 
    99930, 99930, 99960, 99970, 99980, 100000, 100000, 100000, 100010, 
    100010, 100020, 100010, _, 99980, 99990, 99980, 99990, 100010, 100030, 
    100060, 100070, 100090, 100090, 100090, 100130, 100160, 100200, 100220, 
    _, 100290, 100320, 100340, 100360, 100370, 100390, 100400, 100400, 
    100410, 100420, _, 100450, 100450, 100460, 100460, 100460, 100440, 
    100440, 100430, 100430, 100410, 100420, 100400, 100400, 100410, 100420, 
    100420, 100400, 100360, 100320, 100280, 100260, 100250, 100260, 100250, 
    100250, 100240, 100230, 100200, 100160, 100120, 100110, 100080, 100040, 
    100030, 100040, 100060, 100080, 100110, 100110, 100140, 100170, 100160, 
    100130, 100150, _, 100190, 100210, 100220, 100230, 100260, 100290, 
    100310, 100350, 100370, 100370, 100380, 100400, 100450, 100460, 100490, 
    100480, 100500, 100520, 100550, 100580, 100570, 100610, 100610, 100620, 
    100620, 100630, 100660, 100700, 100740, 100800, 100820, 100850, 100870, 
    100880, 100890, 100900, 100910, 100930, 100950, 100980, 100970, 100990, 
    100980, 100970, 100930, 100940, 100890, 100850, 100840, 100820, _, 
    100850, 100840, 100830, 100810, 100800, 100800, 100800, 100790, 100800, 
    100790, 100790, 100800, 100780, 100770, 100730, 100720, 100700, 100700, 
    100670, 100660, _, 100660, 100660, 100670, 100660, 100640, 100640, 
    100660, 100670, 100660, 100660, 100680, 100680, 100670, 100700, 100710, 
    100740, 100750, 100760, 100770, 100770, 100800, 100800, 100840, 100870, 
    100910, 100950, 100980, 101000, 101010, 101000, 100990, 100970, 100970, 
    100960, 100930, 100880, 100850, 100840, 100820, 100800, 100750, 100720, 
    100700, 100640, 100590, 100540, 100470, 100400, 100360, 100320, 100240, 
    100200, 100140, 100100, 100040, 100000, 99960, 99910, 99890, 99880, 
    99850, 99860, 99850, 99840, 99830, 99830, 99830, 99830, 99830, 99870, 
    99890, _, 99950, 99990, 100050, 100120, 100140, 100160, 100240, 100290, 
    100350, 100390, 100420, 100480, 100590, 100670, 100760, 100840, 100920, 
    100980, 101060, 101120, 101160, 101220, _, _, _, _, _, 101430, 101440, 
    101460, 101450, _, 101460, 101460, 101470, 101460, 101450, 101440, 
    101420, 101420, 101420, 101410, 101400, 101370, 101360, 101330, 101290, 
    101250, 101240, 101230, _, 101210, 101190, 101180, 101170, 101160, 
    101150, 101120, 101100, 101100, 101100, 101130, 101150, 101130, 101110, 
    101090, 101080, 101030, 101000, 100980, _, 101020, _, 101070, 101100, 
    101130, 101150, 101160, 101190, 101210, 101190, 101190, 101210, 101210, 
    101220, 101250, 101280, 101310, 101340, 101360, 101390, 101400, 101390, 
    101380, 101360, 101370, 101360, 101350, 101330, 101300, 101260, 101270, 
    101260, 101250, 101210, 101180, 101190, 101180, 101200, 101250, 101310, 
    101370, 101430, _, 101470, 101470, 101450, 101430, 101410, 101380, 
    101380, 101340, 101300, 101290, 101250, 101200, 101150, 101070, 101000, 
    100930, 100870, 100830, 100780, 100730, 100690, 100660, 100630, 100640, 
    100630, 100630, 100620, 100650, 100670, 100700, 100780, 100820, 100880, 
    100900, 100920, 100960, 100930, 100910, 100880, 100880, 100820, 100780, 
    100710, 100650, 100650, 100600, 100510, 100490, 100440, 100430, _, 
    100370, 100360, 100350, 100440, 100500, 100580, 100590, _, 100630, 
    100600, 100600, 100600, 100600, 100580, 100570, 100570, 100590, 100600, 
    100600, 100590, 100570, 100570, 100590, 100570, 100530, 100480, 100460, 
    100460, 100490, 100560, 100610, 100650, 100700, 100730, 100740, 100780, 
    100800, 100850, 100880, 100880, 100910, 100930, 100950, 100950, 100950, 
    100950, 100950, 100940, 100950, 100980, 100970, 101010, 101060, 101090, 
    101090, 101060, 101060, 101060, 101040, 101020, 101020, 101000, 100990, 
    100980, 100980, 100980, 100940, 100890, 100870, 100820, 100810, _, 
    100740, 100700, 100660, 100620, 100600, 100610, 100570, 100550, 100520, 
    100460, 100430, 100410, 100370, 100340, 100290, 100260, 100270, 100240, 
    100210, 100220, 100200, _, 100210, _, 100190, 100190, 100190, 100190, 
    100190, 100210, 100210, 100210, 100200, 100210, 100220, 100240, 100250, 
    100250, 100280, 100330, 100360, 100400, 100430, 100470, 100510, 100520, 
    100530, 100540, 100550, 100570, 100590, 100580, 100560, 100540, 100530, 
    100520, 100490, 100450, 100440, 100420, 100400, 100380, 100390, 100430, 
    100480, 100500, 100540, 100560, 100550, 100520, 100490, _, 100450, 
    100460, 100450, 100450, 100470, 100490, 100490, 100480, 100490, 100460, 
    100430, 100390, 100330, 100290, 100260, 100210, 100190, 100160, 100130, 
    100110, 100070, 100050, 100000, _, 99860, 99860, 99880, 99930, 100000, 
    100040, 100060, 100090, 100100, 100070, 100040, 100010, 100000, 99970, 
    99950, 99950, 99920, 99910, 99920, 99900, 99870, 99850, 99830, 99830, 
    99810, 99800, 99790, 99780, 99780, 99780, 99790, 99780, 99770, 99760, 
    99770, 99770, 99760, 99750, 99750, 99750, _, 99780, 99780, 99770, 99750, 
    99720, 99700, _, 99650, 99650, 99630, 99600, 99590, 99590, 99590, 99550, 
    99530, 99520, 99510, 99490, 99480, 99480, 99470, 99470, 99490, 99490, 
    99510, 99540, 99550, 99570, 99570, 99580, 99610, 99620, 99650, 99680, 
    99720, 99780, 99790, 99830, 99860, 99910, 99940, 99980, 100010, 100050, 
    100090, 100130, 100170, 100200, 100250, 100290, 100340, 100370, 100410, 
    100450, 100480, 100490, 100540, 100580, 100640, 100690, 100750, 100800, 
    100860, 100900, 100940, 100990, 101020, 101060, 101100, 101150, 101190, 
    101250, 101290, 101340, 101380, 101400, 101420, 101440, 101460, 101480, 
    101480, 101480, 101500, 101500, 101500, 101490, 101490, 101490, 101470, 
    101460, 101440, 101420, 101410, 101390, 101340, 101310, 101280, 101270, 
    101230, 101200, 101160, 101120, 101080, 101040, 101030, 101000, 100970, 
    100980, 100950, 100910, 100890, 100840, 100830, 100800, 100760, 100710, 
    100670, 100630, 100600, 100570, 100550, 100520, 100490, 100480, 100400, 
    _, 100350, 100330, 100290, 100270, 100210, 100180, 100130, 100110, 
    100140, 100080, 100040, 100010, 99980, 99960, 99890, 99880, 99850, 99820, 
    99790, 99790, 99750, 99720, 99670, _, 99630, 99600, 99570, 99580, 99550, 
    99570, 99580, 99570, 99600, 99640, 99670, 99670, 99690, 99710, 99700, 
    99700, 99730, 99760, 99800, 99840, _, _, 99950, _, 100020, 100040, 
    100100, 100160, 100210, 100240, 100300, 100330, _, 100420, 100440, 
    100470, 100500, 100520, 100560, 100590, 100650, 100670, 100720, 100760, 
    100800, 100840, 100870, 100890, 100910, 100940, 100950, 100970, 100980, 
    101020, 101040, 101060, 101070, 101080, 101090, 101090, 101090, 101120, 
    101150, 101170, 101190, 101200, 101220, 101250, 101260, 101280, 101290, 
    101300, 101320, 101350, 101370, 101410, 101440, 101470, 101500, 101540, 
    101570, 101570, 101600, 101610, 101590, 101600, 101620, 101640, 101670, 
    101650, 101670, 101660, 101660, 101660, 101660, 101650, 101640, 101610, 
    101550, 101510, 101480, 101420, 101390, 101310, 101240, 101180, 101120, 
    101020, 100920, 100820, 100770, 100650, 100570, 100520, 100480, 100390, 
    100340, 100300, 100190, 100110, 100040, 99990, 99920, 99860, 99830, 
    99810, 99800, 99800, 99810, 99810, 99830, 99860, 99870, 99880, 99890, 
    99960, 100030, 100140, 100190, 100250, 100310, 100380, 100430, 100480, 
    100550, 100600, 100630, 100630, 100670, 100720, 100750, 100770, 100790, 
    100810, 100840, 100850, 100880, 100930, 100970, 101000, 100990, 101000, 
    101020, 101030, 101030, 101040, 101050, 101060, 101080, 101100, 101140, 
    101180, 101200, _, 101260, 101300, 101310, 101320, 101340, 101350, 
    101370, _, _, 101380, 101400, 101430, 101440, 101430, 101450, _, 101470, 
    101450, 101480, 101500, 101510, 101520, 101550, 101570, 101580, 101600, 
    101610, 101620, 101600, 101600, 101620, 101630, 101620, 101620, 101590, 
    101590, 101580, 101580, 101600, 101620, 101590, 101570, 101540, 101540, 
    101540, 101540, 101520, 101520, 101510, 101510, 101510, 101500, 101490, 
    101460, 101440, 101440, 101430, 101410, 101390, 101380, 101360, 101360, 
    101360, 101350, 101350, 101340, 101340, 101350, 101340, 101340, 101350, 
    101350, 101340, 101340, 101340, 101330, 101310, 101280, 101240, 101210, 
    101180, 101150, 101120, 101100, 101090, 101080, 101060, 101010, 100970, 
    100930, 100920, 100890, 100840, 100830, 100820, 100810, 100800, 100770, 
    100770, 100760, 100770, 100750, 100740, 100750, 100750, 100770, 100780, 
    100780, 100780, 100820, 100840, 100840, 100860, 100860, 100860, 100870, 
    100900, 100950, 101000, 101030, 101050, 101100, 101130, 101160, 101200, 
    101220, 101250, 101250, 101270, 101310, 101330, 101340, 101340, 101350, 
    101340, 101330, 101310, 101310, 101300, 101310, 101300, 101310, 101300, 
    101320, 101320, 101340, 101320, 101320, 101330, 101330, 101310, 101300, 
    101320, 101330, 101340, 101370, 101380, 101380, 101370, 101360, 101360, 
    101360, 101350, 101360, 101360, 101390, 101390, 101390, 101390, 101390, 
    101380, 101370, 101360, 101320, 101300, 101310, 101310, 101290, 101280, 
    101280, 101270, 101230, 101220, 101190, 101180, 101150, 101140, 101140, 
    101120, 101100, 101100, 101100, 101110, 101120, 101120, 101120, 101080, 
    101070, 101050, 101040, 101020, 101030, 101010, 101020, 101020, 101020, 
    101030, 101030, 101040, 101030, 101000, 100980, 100960, 100970, 100910, 
    100900, 100900, 100880, 100840, 100800, 100750, 100710, 100670, 100630, 
    100560, 100520, 100450, 100420, 100340, 100230, 100120, 100070, 100020, 
    99980, 99950, 99970, 99920, 99920, 99940, 100010, 100030, 100060, 100080, 
    100140, 100200, 100250, 100310, 100360, 100420, 100490, 100550, 100610, 
    100660, 100720, 100760, 100810, 100850, 100900, 100940, 100990, 101030, 
    101070, 101130, 101170, 101240, 101290, 101350, 101370, 101400, 101400, 
    101430, 101440, 101460, 101470, 101480, 101510, 101510, 101520, 101530, 
    101520, 101510, 101510, 101500, 101500, 101500, 101490, 101490, 101530, 
    101550, 101560, 101530, 101520, 101460, 101470, 101460, 101470, 101500, 
    101500, 101480, 101510, 101490, 101490, 101490, 101460, 101440, 101440, 
    101410, 101400, 101390, 101390, 101340, 101320, 101300, 101300, 101310, 
    101280, 101260, 101220, 101220, 101220, 101210, 101230, 101240, 101250, 
    101240, 101240, 101250, 101240, 101250, 101280, 101300, 101310, 101320, 
    101340, 101360, 101370, 101390, 101400, 101400, 101410, 101400, 101390, 
    101390, 101370, 101380, 101390, 101370, 101370, 101380, 101360, 101320, 
    101300, 101270, 101230, 101200, 101190, 101170, 101140, 101110, 101110, 
    101080, 101080, 101020, 100970, 100940, 100900, 100840, 100780, 100710, 
    100680, 100640, 100620, 100550, 100490, 100440, 100420, 100380, 100370, 
    100370, 100350, 100350, 100370, 100390, 100410, 100450, 100460, 100500, 
    100500, 100520, 100560, 100560, 100580, 100600, 100630, 100650, 100670, 
    100680, 100670, 100690, 100670, 100670, 100670, 100670, 100660, 100680, 
    100670, 100670, 100670, 100670, 100670, 100660, 100650, 100650, 100630, 
    100650, 100650, 100660, 100650, 100670, 100680, 100680, 100680, 100670, 
    100670, 100670, 100640, 100640, 100640, 100590, 100550, 100520, 100500, 
    100470, 100440, 100390, 100360, 100300, 100190, 100140, 100050, 100010, 
    99960, 99940, 99940, 99970, 99990, 99990, 100020, 100050, 100080, 100130, 
    100180, 100250, 100290, 100340, 100350, 100390, 100420, 100410, 100410, 
    100380, 100340, 100310, 100270, 100220, 100200, 100170, 100150, 100100, 
    100050, 100010, 99980, 99910, 99840, 99780, 99730, 99680, 99640, 99600, 
    99570, 99560, 99520, 99440, 99370, 99320, 99290, 99280, 99260, 99250, 
    99260, 99270, 99280, 99300, 99310, 99340, 99360, 99380, 99380, 99430, 
    99450, 99500, 99530, 99540, 99550, 99570, 99580, 99590, 99580, 99570, 
    99550, 99530, 99490, 99480, 99490, 99480, 99490, 99500, 99510, 99530, 
    99570, 99610, 99640, 99730, 99800, 99870, 99930, 100010, 100060, 100120, 
    100160, 100230, 100270, 100310, 100340, 100370, 100390, 100410, 100400, 
    100410, 100390, 100310, 100240, 100140, 100040, 99930, 99870, 99790, 
    99720, 99660, 99640, 99630, 99640, 99670, 99720, 99810, 99860, 99910, 
    99970, 100020, 100030, 100060, 100090, 100140, 100170, 100190, 100210, 
    100210, 100200, 100210, 100220, 100210, 100200, 100190, 100180, 100180, 
    100160, 100180, 100170, 100190, 100170, 100150, 100140, 100120, 100130, 
    100160, 100170, 100190, 100200, 100220, 100230, 100250, 100280, 100310, 
    100320, 100350, 100370, 100390, 100410, 100430, 100460, 100480, 100490, 
    100520, 100520, 100510, 100480, 100480, 100490, 100520, 100510, 100550, 
    100540, 100510, 100490, 100450, 100450, 100430, 100410, 100370, 100390, 
    100380, 100420, 100440, 100410, 100450, 100470, 100500, 100460, 100440, 
    100450, 100430, 100390, 100390, 100410, 100370, 100360, 100340, 100300, 
    100280, 100270, 100270, 100270, 100270, 100280, 100250, 100270, 100290, 
    100280, 100270, 100250, 100260, 100280, 100320, 100320, 100280, 100250, 
    100270, 100290, 100290, 100280, 100250, 100200, 100170, 100120, 100070, 
    100080, 100080, 100060, 100040, 100060, 100080, 100090, 100050, 100030, 
    100020, 99970, 99930, 99890, 99870, 99830, 99810, 99790, 99760, 99760, 
    99750, 99740, 99740, 99740, 99730, 99740, 99740, 99760, 99740, 99750, 
    99770, 99800, 99810, 99810, 99850, 99860, 99860, 99860, 99880, 99870, 
    99880, 99880, 99890, 99940, 99940, 99980, 99990, 100000, 100010, 100030, 
    100030, 100050, 100050, 100060, 100090, 100110, 100130, 100140, 100170, 
    100210, 100230, 100250, 100250, 100240, 100260, 100300, 100340, 100350, 
    100380, 100420, 100440, 100470, 100490, 100520, 100540, 100540, 100570, 
    100590, 100600, 100630, 100640, 100650, 100670, 100670, 100660, 100650, 
    100620, 100590, 100550, 100530, 100530, 100480, 100440, 100410, 100340, 
    100260, 100190, 100140, 100080, 100020, 100000, 100000, 100000, 99980, 
    100090, 100190, 100320, 100440, 100560, 100660, 100760, 100860, 100930, 
    101020, 101110, 101200, 101270, 101310, 101360, 101420, 101450, 101480, 
    101520, 101540, 101580, 101600, 101650, 101670, 101700, 101720, 101720, 
    101720, 101720, 101730, 101700, 101700, 101690, 101680, 101660, 101640, 
    101610, 101540, 101490, 101450, 101400, 101330, 101250, 101180, 101090, 
    101040, 100960, 100870, 100800, 100740, 100720, 100680, 100590, 100460, 
    100370, 100310, 100270, 100230, 100180, 100150, 100090, 100010, 99910, 
    99810, 99670, 99550, 99500, 99440, 99350, 99280, 99230, 99200, 99140, 
    99130, 99110, 99100, 99110, 99130, 99140, 99160, 99140, 99200, 99230, 
    99250, 99280, 99300, 99320, 99350, 99370, 99380, 99380, 99390, 99400, 
    99400, 99410, 99400, 99420, 99420, 99430, 99430, 99410, 99410, 99410, 
    99420, 99420, 99400, 99400, 99400, 99390, 99350, 99340, 99320, 99290, 
    99270, 99260, 99230, 99200, 99180, 99160, 99130, 99110, 99060, 99060, 
    99040, 99010, 98980, 98960, 98990, 98980, 98960, 98920, 98920, 98900, 
    98900, 98920, 98940, 98960, 98980, 99000, 99070, 99110, 99150, 99190, 
    99210, 99250, 99340, 99370, 99460, 99510, 99590, 99600, 99690, 99780, 
    99840, 99920, 99980, 100030, 100110, 100160, 100240, 100280, 100330, 
    100370, 100440, 100500, 100550, 100600, 100660, 100710, 100770, 100810, 
    100830, 100880, 100920, 100940, 100970, 100990, 101020, 101030, 101070, 
    101120, 101150, 101180, 101210, 101220, 101260, 101260, 101280, 101310, 
    101330, 101350, 101380, 101400, 101420, 101420, 101430, 101440, 101430, 
    101460, 101430, 101460, 101450, 101480, 101480, 101490, 101490, 101490, 
    101480, 101470, 101450, 101450, 101440, 101440, 101430, 101430, 101430, 
    101440, 101430, 101410, 101400, 101390, 101390, 101380, 101370, 101360, 
    101370, 101370, 101390, 101380, 101370, 101380, 101370, 101370, 101370, 
    101380, 101360, 101340, 101330, 101350, 101360, 101360, 101370, 101360, 
    101320, 101270, 101250, 101230, 101220, 101190, 101170, 101160, 101170, 
    101190, 101190, 101180, 101130, 101090, 101050, 100990, 100960, 100900, 
    100850, 100850, 100820, 100800, 100740, 100700, 100670, 100650, 100640, 
    100630, 100620, 100620, 100600, 100600, 100610, 100600, 100590, 100580, 
    100520, 100480, 100430, 100400, 100380, 100370, 100370, 100370, 100330, 
    100340, 100330, 100280, 100230, 100190, 100130, 100100, 100130, 100150, 
    100160, 100160, 100140, 100130, 100070, 100060, 100010, 100000, 99970, 
    99960, 99940, 99940, 99920, 99890, 99850, 99870, 99870, 99880, 99910, 
    99930, 99930, 99940, 99950, 99960, 99960, 99990, 100000, 100020, 100010, 
    100010, 100030, 100060, 100060, 100060, 100030, 100010, 100000, 99990, 
    99960, 99940, 99910, 99870, 99810, 99770, 99730, 99720, 99730, 99750, 
    99810, 99840, 99890, 99950, 100030, 100090, 100120, 100160, 100190, 
    100200, 100240, 100250, 100240, 100210, 100160, 100060, 99970, 99920, 
    99890, 99800, 99780, 99760, 99740, 99790, 99840, 99900, 99970, 100070, 
    100160, 100240, 100300, 100340, 100390, 100440, 100490, 100510, 100560, 
    100570, 100590, 100600, 100570, 100560, 100540, 100490, 100480, 100480, 
    100470, 100490, 100500, 100570, 100620, 100690, 100760, 100790, 100870, 
    100900, 100990, 101000, 101110, 101180, 101230, 101270, 101320, 101360, 
    101380, 101420, 101440, 101440, 101440, 101460, 101440, 101480, 101450, 
    101410, 101420, 101370, 101360, 101350, 101300, 101230, 101180, 101130, 
    101080, 101050, 100990, 100920, 100830, 100770, 100710, 100630, 100550, 
    100500, 100440, 100380, 100330, 100300, 100280, 100280, 100240, 100240, 
    100240, 100260, 100280, 100280, 100270, 100270, 100260, 100250, 100250, 
    100270, 100270, 100310, 100340, 100360, 100350, 100350, 100330, 100330, 
    100330, 100340, 100320, 100350, 100350, 100360, 100400, 100460, 100480, 
    100510, 100560, 100580, 100610, 100630, 100660, 100670, 100670, 100720, 
    100730, 100730, 100690, 100640, 100610, 100570, 100580, 100560, 100540, 
    100510, 100490, 100470, 100440, 100410, 100340, 100240, 100200, 100150, 
    100130, 100150, 100100, 100080, 100080, 100070, 100040, 100030, 100000, 
    100030, 100020, 100000, 100020, 100050, 100090, 100130, 100180, 100230, 
    100280, 100270, 100260, 100270, 100290, 100270, 100260, 100230, 100240, 
    100250, 100280, 100320, 100360, 100410, 100450, 100460, 100470, 100500, 
    100520, 100550, 100590, 100610, 100610, 100630, 100640, 100660, 100680, 
    100710, 100730, 100780, 100810, 100860, 100930, 101000, 101040, 101090, 
    101150, 101190, 101230, 101230, 101270, 101290, 101330, 101370, 101410, 
    101440, 101450, 101460, 101490, 101500, 101490, 101480, 101490, 101490, 
    101480, 101480, 101500, 101490, 101470, 101410, 101380, 101350, 101340, 
    101300, 101280, 101230, 101200, 101190, 101170, 101180, 101190, 101160, 
    101110, 101080, 101070, 101070, 101030, 101030, 101050, 101010, 101010, 
    101060, 101110, 101120, 101090, 101070, 101050, 101110, 101120, 101130, 
    101160, 101190, 101210, 101210, 101230, 101230, 101210, 101230, 101250, 
    101270, 101260, 101270, 101310, 101350, 101370, 101380, 101430, 101480, 
    101480, 101510, 101520, 101540, 101580, 101600, 101620, 101660, 101690, 
    101690, 101700, 101720, 101740, 101760, 101780, 101790, 101800, 101820, 
    101830, 101850, 101870, 101890, 101910, 101910, 101910, 101910, 101910, 
    101920, 101930, 101940, 101960, 101970, 101980, 101980, 101990, 101990, 
    102010, 102020, 102040, 102040, 102040, 102080, 102080, 102100, 102100, 
    102110, 102130, 102140, 102100, 102110, 102100, 102090, 102100, 102120, 
    102100, 102140, 102140, 102150, 102170, _, 102210, 102220, 102230, 
    102230, 102250, 102270, 102330, 102360, 102400, 102420, 102400, 102400, 
    102420, 102420, 102420, _, 102400, 102440, 102450, 102470, 102470, 
    102490, 102500, 102510, 102540, 102590, 102600, 102620, 102630, 102640, 
    102670, 102690, 102760, 102800, 102820, 102860, 102910, 102940, 102970, 
    103000, 103040, 103050, 103080, 103120, 103160, _, _, 103260, 103280, 
    103300, 103320, 103320, 103340, 103330, 103320, 103340, 103360, 103360, 
    103370, 103390, 103380, 103380, 103390, 103370, 103380, 103360, 103350, 
    _, 103350, 103350, 103360, 103360, 103340, 103320, 103290, 103280, 
    103270, 103260, 103240, 103210, 103190, 103180, 103190, 103180, 103180, 
    103160, 103160, _, 103140, 103130, 103140, 103140, 103120, 103120, 
    103130, 103130, 103120, 103110, 103100, 103090, 103080, 103060, _, 
    103050, 103060, 103030, 103020, 103010, 103000, 102990, 102980, 102990, 
    102980, 102960, 102960, 102970, 102960, 102980, 102970, 102990, 102990, 
    102980, 102970, 102960, 102950, 102970, 102980, 102990, 102970, 102980, 
    102990, 102980, 102970, 102940, 102960, 102950, 102940, 102900, 102870, 
    102870, 102850, 102880, 102910, 102900, 102930, 102940, 102930, 102920, 
    102890, 102890, 102870, 102870, 102870, 102850, 102830, 102830, 102840, 
    102820, 102800, 102790, 102770, 102750, 102730, 102730, 102720, 102720, 
    102720, 102720, _, _, _, _, _, _, _, 102590, _, _, _, _, 102520, _, _, _, 
    _, _, _, 102390, _, _, _, _, 102290, 102280, 102270, 102290, 102260, 
    102230, 102230, 102230, 102230, 102210, 102220, 102220, 102210, 102200, 
    102180, 102130, 102110, 102070, 102040, 102000, 101950, 101900, 101860, 
    101820, 101760, 101700, 101610, 101480, 101350, 101250, 101130, 100980, 
    100870, 100750, 100630, 100540, 100440, 100310, 100190, 100080, 100000, 
    99920, 99880, 99800, 99740, 99680, 99580, 99500, 99440, 99370, 99390, 
    99410, 99410, 99390, 99390, 99420, 99480, 99530, 99590, 99630, 99680, 
    99700, 99720, 99700, 99650, 99600, 99530, 99500, 99470, 99420, 99360, 
    99280, 99180, 99080, 98960, 98900, 98890, 98910, 98910, 98930, 99000, 
    99070, 99130, 99190, 99220, 99280, 99360, 99420, 99490, 99540, 99610, 
    99680, 99770, 99820, 99870, 99920, 99960, 100030, 100050, 100070, 100080, 
    100130, 100140, 100140, 100190, 100220, 100250, 100310, 100340, 100370, 
    100400, 100430, 100430, 100480, 100500, 100500, 100530, 100560, 100590, 
    100620, 100640, 100680, 100680, 100680, 100700, 100700, 100700, 100710, 
    100720, 100760, 100760, 100770, 100780, 100770, 100760, 100780, 100830, 
    100820, 100860, 100890, 100950, 100950, 100970, 100980, 100990, 101000, 
    101040, 101020, 101030, 101020, 101040, 101020, 101020, 101050, 101010, 
    101000, 101000, 100970, 100960, 100940, 100940, 100910, 100900, 100910, 
    100900, 100920, 100950, 100970, 100990, 101020, 101050, 101080, 101060, 
    101090, 101080, 101130, 101130, 101130, 101160, 101200, 101220, 101250, 
    101240, 101290, 101300, 101330, 101350, 101390, 101420, 101440, 101480, 
    101500, 101500, 101520, 101520, 101520, 101520, 101510, 101520, 101520, 
    101520, 101510, 101510, 101500, 101480, 101480, 101470, 101440, 101410, 
    101400, 101400, 101410, 101410, 101410, 101420, 101410, 101400, 101390, 
    101360, 101310, 101300, 101270, 101230, 101200, 101170, 101120, 101090, 
    101060, 101020, 101000, 100940, 100880, 100840, 100810, 100770, 100730, 
    100690, 100680, 100660, 100630, 100600, 100550, 100500, 100440, 100410, 
    100390, 100360, 100320, 100300, 100270, 100210, 100170, 100120, 100080, 
    100020, 99970, _, 99860, 99800, 99730, 99670, 99630, 99580, 99490, 99420, 
    _, _, 99330, 99300, 99290, _, 99300, 99330, 99330, 99360, 99370, 99390, 
    99440, 99480, 99490, 99550, 99610, 99690, 99780, 99880, 99980, 100120, 
    100230, 100360, 100480, 100560, 100650, 100740, 100830, 100890, 100980, 
    101010, 101070, 101120, 101160, 101180, 101140, 101170, 101140, 101110, 
    101090, 101070, 101080, 101030, 101010, 101010, 101040, 101060, 101050, 
    101080, 101120, 101190, 101270, 101380, 101500, 101610, 101770, 101900, 
    102020, 102070, 102170, 102240, 102290, 102290, 102330, 102330, 102310, 
    102270, 102260, 102270, 102220, 102180, 102110, 102040, 101980, 101920, 
    101860, 101790, 101750, 101710, 101690, 101650, 101600, 101540, 101480, 
    101430, 101360, 101290, 101250, 101190, 101110, 101070, 101020, 100980, 
    100980, 100980, 100980, 100960, 100950, 100950, 100960, 101010, 101070, 
    101140, 101240, 101360, 101400, 101450, 101500, 101550, 101590, 101640, 
    101690, 101710, 101740, 101800, 101850, 101900, 101930, 101950, 101950, 
    101970, 101970, 101990, 101980, 101970, 101950, 101960, 101960, 101950, 
    101910, 101870, 101840, 101820, 101790, 101760, 101710, 101670, 101640, 
    101600, 101580, 101550, 101490, 101420, 101350, 101310, 101240, 101170, 
    101120, 101050, 101010, 100970, 100930, 100890, 100860, 100810, 100790, 
    100750, 100730, 100670, 100650, 100630, 100630, 100620, 100630, 100630, 
    100660, 100650, 100640, 100640, 100640, 100670, 100720, 100720, 100740, 
    100760, 100810, 100830, 100850, 100890, 100920, 100920, 100960, 100980, 
    101020, 101050, 101070, 101130, 101140, 101180, 101230, 101270, 101300, 
    101340, 101380, 101420, 101440, 101450, 101480, 101510, 101540, 101580, 
    101590, 101610, 101610, 101620, 101630, 101650, 101660, 101680, 101680, 
    101670, 101700, 101710, 101730, 101750, 101750, 101750, 101750, 101760, 
    101770, 101790, 101800, 101820, 101850, 101850, 101840, 101840, 101830, 
    101820, 101820, 101790, 101770, 101740, 101720, 101690, 101680, 101660, 
    101630, 101600, 101570, 101520, 101480, 101450, 101420, 101370, 101320, 
    101280, 101240, 101200, 101150, 101110, 101070, 101020, 100990, 100950, 
    100930, 100910, 100890, 100880, 100880, 100870, 100810, 100780, 100760, 
    100760, 100720, 100660, 100610, 100570, 100550, 100530, 100530, 100520, 
    100500, 100500, 100470, 100440, 100440, 100430, 100430, 100400, 100400, 
    100390, 100390, 100400, 100400, 100380, 100350, 100330, 100300, 100260, 
    100250, 100240, 100200, 100200, 100170, 100150, 100150, 100130, 100110, 
    100110, 100100, 100090, 100080, 100080, 100080, 100100, 100130, 100160, 
    100160, 100170, 100180, 100180, 100200, 100210, 100220, 100220, 100240, 
    100240, 100240, 100260, 100270, 100260, 100260, 100260, 100260, 100250, 
    100230, 100230, 100250, 100260, 100290, 100320, 100330, 100320, 100340, 
    100340, 100320, 100320, 100300, 100290, 100290, 100280, 100270, 100260, 
    100240, 100170, 100140, 100110, 100060, 100020, 100000, 100000, 100000, 
    100010, 100020, 100030, 100030, 100050, 100050, 100060, 100080, _, 
    100140, 100170, 100170, 100190, 100180, 100210, 100220, 100230, 100240, 
    100240, 100230, 100230, 100220, 100220, 100210, 100210, 100220, 100230, 
    100240, 100230, 100220, 100210, 100200, 100200, 100200, 100190, 100180, 
    100170, 100170, 100160, 100150, 100150, 100130, 100120, 100090, 100080, 
    100060, 100050, 100040, 100040, 100040, 100040, 100050, 100050, 100050, 
    100040, 100040, 100030, 100010, 100020, 100020, 100010, 100010, 100000, 
    99990, 99980, 99970, 99960, 99950, 99940, 99920, 99920, 99920, 99950, 
    99960, 99980, 99970, 99980, 100010, 100020, 100010, 100020, 100030, 
    100040, 100060, 100080, 100100, 100110, 100110, 100140, 100150, 100170, 
    100170, 100200, 100220, 100230, 100260, 100310, 100320, 100350, 100370, 
    100370, 100420, 100420, 100420, 100410, 100440, 100430, 100460, 100460, 
    100450, 100440, 100450, 100450, 100420, 100380, 100370, 100340, 100300, 
    100290, 100290, 100290, 100280, 100290, 100280, 100290, 100280, 100270, 
    100300, 100330, 100350, 100400, 100440, 100480, 100520, _, 100610, 
    100660, 100670, 100700, 100730, 100720, 100730, _, 100760, 100790, 
    100810, 100820, 100860, 100890, 100890, 100880, 100880, 100860, 100860, 
    100860, 100840, 100840, 100850, 100850, 100830, 100850, 100840, 100840, 
    100830, 100800, 100770, 100740, 100740, 100730, 100740, 100760, 100760, 
    100760, 100760, 100710, 100690, 100690, 100660, 100630, 100620, 100600, 
    100590, 100600, 100580, 100570, 100550, 100520, 100480, _, 100350, 
    100300, 100260, 100210, 100190, 100160, 100110, 100090, _, 100030, 99970, 
    99880, 99800, 99770, 99730, 99650, 99610, _, 99520, 99470, 99410, 99370, 
    99340, 99320, 99290, _, 99200, 99170, 99140, 99100, 99090, 99060, 99030, 
    99040, 99050, 99030, 99040, 99070, 99100, 99140, 99160, 99200, 99240, 
    99260, 99270, 99280, 99330, _, 99370, 99390, 99410, 99440, 99460, 99460, 
    99440, 99430, 99420, 99370, 99330, 99290, 99230, 99140, 99030, 98960, 
    98860, 98750, 98720, 98600, 98430, 98280, 98150, _, 98000, 97930, 97860, 
    97790, 97760, 97770, 97770, 97760, 97740, 97710, 97690, 97660, 97640, 
    97580, 97570, 97550, 97580, 97600, _, 97670, 97650, 97680, 97670, 97660, 
    97670, 97710, 97720, 97780, 97870, 97940, 98030, 98070, 98120, 98140, 
    98180, 98200, 98230, 98250, 98250, 98250, 98230, 98220, 98200, 98220, 
    98180, 98160, 98150, _, 98130, 98100, 98090, 98060, 98070, 98070, 98060, 
    98040, 98030, 98010, 97970, 97980, 98030, 98020, 98000, 98000, 98040, 
    98140, 98240, 98370, 98490, 98570, 98660, 98730, 98810, 98900, 98950, 
    99040, 99120, 99200, 99280, 99350, 99410, 99500, 99560, 99630, 99680, 
    99730, 99780, 99830, 99880, _, 99960, 99980, _, _, _, 99970, 99960, _, 
    99950, 99920, 99930, 99920, 99870, 99860, 99830, 99850, 99830, 99730, 
    99690, 99650, 99580, 99510, 99470, 99410, 99410, 99380, 99350, 99310, 
    99290, _, 99240, 99200, 99190, 99170, 99150, 99130, 99130, 99100, 99080, 
    99060, 99030, 98990, 98940, 98900, 98840, 98780, 98760, 98730, 98710, 
    98680, 98650, 98650, 98680, 98720, 98730, 98750, 98800, 98830, 98860, 
    98930, 98980, 99040, 99090, 99140, 99150, 99160, 99190, 99220, 99270, 
    99320, 99350, 99390, 99410, 99450, 99480, 99480, 99490, 99470, 99450, 
    99450, 99430, 99420, 99400, 99410, 99400, 99380, 99340, 99310, 99280, 
    99270, 99250, 99210, 99200, 99190, 99220, 99230, 99240, 99260, 99280, 
    99280, 99270, 99310, 99330, 99360, 99420, 99500, 99580, 99650, 99760, 
    99820, 99860, 99890, 99960, 100000, 100030, 100090, 100140, 100150, 
    100220, 100260, 100320, 100340, 100380, 100430, 100460, 100490, 100500, 
    100520, 100550, 100550, 100600, 100640, 100610, 100620, 100590, 100560, 
    100460, 100390, 100300, 100190, 100130, 100020, 99930, 99840, 99710, 
    99550, 99400, 99230, 98860, 98750, 98450, 98030, 97680, 97260, 96930, 
    96690, 96480, 96320, 96190, 96090, 96020, 95940, 95860, 95850, 95850, 
    95870, 95940, 96020, 96110, 96180, 96250, 96350, 96420, 96480, 96580, 
    96670, 96790, 96830, 96930, 97020, 97080, 97130, 97190, 97240, 97270, 
    97260, 97260, 97270, 97290, 97280, 97320, 97300, 97320, 97300, 97310, 
    97360, 97350, 97390, 97450, 97480, 97570, 97590, 97630, 97690, 97720, 
    97790, 97850, 97910, 97980, 98040, 98080, 98150, 98210, 98290, 98360, 
    98420, 98470, 98510, 98530, 98540, 98580, 98580, 98660, 98700, 98710, 
    98720, 98780, 98820, 98850, 98850, 98900, 98910, 98930, 98940, 98950, 
    98970, 98980, 98980, 98990, 98990, 98960, 98930, 98910, 98890, 98870, 
    98850, 98840, 98830, 98820, 98830, 98860, 98870, 98890, 98890, 98920, 
    98970, 99000, 99020, 99050, 99080, 99100, 99140, 99160, 99180, 99230, 
    99230, 99260, 99290, 99340, 99400, 99410, 99440, 99480, 99480, 99540, 
    99580, 99580, 99590, 99590, 99620, 99660, 99680, 99700, 99720, 99750, 
    99800, 99820, 99850, 99880, 99920, 99930, 99930, 99960, 99950, 99930, 
    99920, 99930, 99940, 99960, 99980, 100010, 100010, 99970, 99950, 99910, 
    99890, 99880, 99810, 99750, 99670, 99630, 99600, 99530, 99470, 99370, 
    99320, 99250, 99200, 99110, 99050, 99000, 98890, 98840, 98720, 98640, 
    98520, 98360, 98260, 98140, 98100, 98030, 98030, 98050, 98100, 98050, 
    98030, 98040, 98040, 98040, 97990, 98030, 98050, 98040, 98010, 97930, 
    97870, 97750, 97780, 97690, 97760, 97840, 97970, 98150, 98320, 98480, 
    98600, 98650, 98710, 98780, 98830, 98850, 98860, 98850, 98850, 98880, 
    98930, 98980, 99060, 99130, 99210, 99340, 99430, 99530, 99590, 99670, 
    99710, 99830, 99910, 100000, 100080, 100140, 100210, 100280, 100320, 
    100390, 100400, 100430, 100400, 100420, 100460, 100490, 100490, 100510, 
    100530, 100560, 100550, 100600, 100630, 100640, 100640, 100660, 100680, 
    100720, 100730, 100740, 100740, 100750, 100780, 100770, 100760, 100760, 
    100730, 100680, 100650, 100600, 100540, 100530, 100510, 100460, 100420, 
    100430, 100390, 100360, 100340, 100320, 100290, 100280, 100260, 100270, 
    100290, 100270, 100280, 100260, 100210, 100150, 100090, 100060, 100020, 
    99960, 99910, 99890, 99870, 99860, 99850, 99810, 99790, 99780, 99800, 
    99830, 99850, 99870, 99920, 99960, 100000, 100040, 100080, 100120, 
    100150, 100200, 100250, 100290, 100310, 100350, 100350, 100390, 100430, 
    100460, 100470, 100460, 100450, 100450, 100450, 100440, 100410, 100360, 
    100340, 100310, 100270, 100250, 100220, 100180, 100120, 100070, 100040, 
    100010, 99950, 99900, 99840, 99790, 99790, 99730, 99700, 99650, 99610, 
    99540, 99500, 99440, 99400, 99360, 99320, 99270, 99220, 99170, 99100, 
    99060, 99050, 99020, 99000, 98960, 98920, 98850, 98840, 98840, 98840, 
    98850, 98820, 98810, 98790, 98780, 98810, 98840, 98820, 98850, 98880, 
    98860, 98880, 98940, 98970, 98960, 99030, 99070, 99130, 99180, 99220, 
    99270, 99330, 99360, 99410, 99460, 99510, 99570, 99620, 99640, 99650, 
    99650, 99670, 99680, 99730, 99770, 99810, 99840, 99870, 99930, 99930, 
    99940, 99960, 99910, 99920, 99960, 99950, 99940, 99900, 99870, 99830, 
    99820, 99780, 99760, 99720, 99660, 99580, 99510, 99420, 99350, 99310, 
    99270, 99230, 99160, 99120, 99060, 99020, 99000, 98960, 98920, 98890, 
    98860, 98840, 98830, 98840, 98850, 98840, 98840, 98860, 98870, 98890, 
    98890, 98890, 98900, 98920, 98950, 98990, 99020, 99040, 99030, 99070, 
    99080, 99100, 99120, 99110, 99130, 99170, 99210, 99250, 99260, 99280, 
    99310, 99320, 99320, 99330, 99350, 99340, 99330, 99360, 99390, 99420, 
    99480, 99520, 99520, 99550, 99550, 99600, 99620, 99620, 99640, 99720, 
    99800, 99880, 99930, 100010, 100080, 100100, 100150, 100190, 100220, 
    100270, 100270, 100300, 100330, 100390, 100440, 100460, 100470, 100510, 
    100530, 100530, 100520, 100520, 100510, 100510, 100540, 100540, 100560, 
    100550, 100540, 100540, 100570, 100580, 100580, 100590, 100600, 100620, 
    100660, 100690, 100680, 100700, 100710, 100730, 100730, 100750, 100740, 
    100740, 100740, 100740, 100760, 100770, 100790, 100790, 100770, 100760, 
    100750, 100730, 100720, 100710, 100700, 100710, 100710, 100730, 100740, 
    100790, 100790, 100800, 100840, 100860, 100840, 100810, 100850, 100870, 
    100900, 100880, 100900, 100910, 100910, 100930, 100940, 100960, 100960, 
    100930, 100930, 100950, 100970, 100970, 100960, 100920, 100900, 100910, 
    100900, 100890, 100890, 100910, 100940, 100950, 100960, 101010, 101020, 
    101030, 101070, 101080, 101100, 101100, 101100, 101080, 101090, 101090, 
    101100, 101080, 101070, 101080, 101100, 101070, 101080, 101050, 101020, 
    101000, 100970, 100950, 100940, 100940, 100940, 100900, 100880, 100870, 
    100880, 100850, 100830, 100790, 100740, 100710, 100670, 100630, 100570, 
    100520, 100440, 100370, 100290, 100190, 100080, 99970, 99870, 99800, 
    99730, 99670, 99590, 99510, 99430, 99370, 99340, 99300, 99310, 99360, 
    99360, 99390, 99380, 99370, 99390, 99400, 99400, 99430, 99420, 99390, 
    99370, 99410, 99440, 99460, 99470, 99470, 99490, 99490, 99520, 99520, 
    99540, 99580, 99600, 99680, 99780, 99860, 99950, 100020, 100130, 100210, 
    100290, 100370, 100430, 100490, 100540, 100580, 100640, 100670, 100700, 
    100740, 100760, 100800, 100810, 100860, 100890, 100870, 100870, 100850, 
    100850, 100840, 100770, 100710, 100670, 100610, 100580, 100570, 100550, 
    100500, 100420, 100310, 100210, 100160, 100160, 100180, 100200, 100220, 
    100250, 100240, 100190, 100140, 100210, 100210, 100210, 100220, 100120, 
    100140, 100140, 100120, 100080, 100040, 99970, 99920, 99850, 99810, 
    99730, 99680, 99660, 99620, 99540, 99450, 99400, 99320, 99240, 99150, 
    99080, 98990, 98890, 98860, 98780, 98680, 98610, 98520, 98420, 98390, 
    98330, 98230, 98200, 98250, 98320, 98320, 98350, 98320, 98310, 98260, 
    98210, 98180, 98140, 98040, 97970, 97830, 97720, 97660, 97610, 97600, 
    97530, 97400, 97360, 97360, 97330, 97360, 97370, 97400, 97410, 97460, 
    97430, 97400, 97370, 97350, 97400, 97460, 97580, 97680, 97840, 97960, 
    98040, 98160, 98280, 98340, 98410, 98540, 98680, 98820, 98930, 99030, 
    99120, 99200, 99310, 99430, 99510, 99620, 99710, 99800, 99870, 99920, 
    99980, 99980, 100000, 99990, 99980, 100010, 100030, 100060, 100090, 
    100130, 100120, 100120, 100150, 100140, 100140, 100130, 100120, 100120, 
    100120, 100120, 100140, 100100, 100060, 100040, 100020, 100010, 100010, 
    100030, 100050, 100070, 100080, 100090, 100140, 100150, 100170, 100140, 
    100150, 100140, 100120, 100100, 100090, 100090, 100060, 100050, 100030, 
    100030, 100030, 100020, 100020, 100030, 100020, 100020, 100020, 100060, 
    100070, 100100, 100100, 100090, 100100, 100100, 100120, 100120, 100100, 
    100080, 100110, 100130, 100150, 100160, 100180, 100200, 100220, 100220, 
    100230, 100250, 100230, 100260, 100260, 100270, 100290, 100320, 100330, 
    100360, 100370, 100440, 100470, 100480, 100490, 100490, 100480, 100510, 
    100530, 100560, 100590, 100600, 100610, 100600, 100630, 100700, 100720, 
    100730, 100730, 100750, 100770, 100750, 100720, 100720, 100760, 100730, 
    100710, 100740, 100710, 100720, 100710, 100700, 100750, 100770, 100760, 
    100760, 100770, 100800, 100820, 100830, 100830, 100830, 100850, 100880, 
    100890, 100940, 100970, 101020, 101040, 101070, 101100, 101130, 101130, 
    101140, 101190, 101180, 101220, 101230, 101300, 101330, 101360, 101350, 
    101330, 101330, 101310, 101330, 101320, 101310, 101340, 101330, 101350, 
    101350, 101310, 101280, 101290, 101240, 101190, 101220, 101210, 101180, 
    101160, 101160, 101130, 101100, 101050, 101010, 100960, 100920, 100890, 
    100850, 100840, 100830, 100810, 100800, 100790, 100740, 100720, 100690, 
    100660, 100620, 100610, 100580, 100540, 100560, 100530, 100530, 100530, 
    100500, 100450, 100430, 100410, 100410, 100390, 100380, 100370, 100340, 
    100350, 100360, 100380, 100380, 100360, 100350, 100380, 100360, 100420, 
    100430, 100460, 100480, 100470, 100500, 100520, 100530, 100520, 100550, 
    100530, 100560, 100530, 100540, 100530, 100540, 100550, 100530, 100530, 
    100510, 100460, 100450, 100430, 100400, 100370, 100360, 100360, 100330, 
    100320, 100350, 100360, 100370, 100310, 100280, 100280, 100300, 100320, 
    100330, 100340, 100360, 100390, 100420, 100470, 100490, 100530, 100570, 
    100590, 100630, 100660, 100690, 100690, 100740, 100800, 100840, 100870, 
    100890, 100920, 100940, 100950, 100990, 101010, 101020, 101060, 101080, 
    101110, 101130, 101160, 101210, 101230, 101250, 101290, 101320, 101330, 
    101350, 101400, 101430, 101480, 101530, 101570, 101600, 101620, 101630, 
    101650, 101650, 101660, 101690, 101740, 101760, 101790, 101820, 101830, 
    101860, 101900, 101900, 101900, 101900, 101930, 101930, 101950, 101980, 
    102030, 102070, 102100, 102120, 102150, 102140, 102160, 102160, 102160, 
    102170, 102170, 102170, 102180, 102180, 102150, 102100, 102060, 102020, 
    101970, 101910, 101850, 101800, 101730, 101670, 101640, 101640, 101610, 
    101590, 101560, 101530, 101520, 101510, 101500, 101510, 101540, 101550, 
    101590, 101610, 101640, 101670, 101690, 101700, 101700, 101710, 101720, 
    101730, 101730, 101730, 101770, 101810, 101820, 101820, 101790, 101770, 
    101730, 101720, 101710, 101700, 101680, 101720, 101730, 101740, 101760, 
    101750, 101720, 101710, 101650, 101620, 101620, 101600, 101590, 101580, 
    101580, 101610, 101600, 101600, 101590, 101580, 101560, 101530, 101500, 
    101460, 101460, 101460, 101440, 101420, 101390, 101370, 101360, 101350, 
    101330, 101310, 101300, 101310, 101280, 101280, 101300, 101340, 101350, 
    101360, 101370, 101400, 101420, 101420, 101440, 101450, 101470, 101500, 
    101510, 101520, 101540, 101540, 101560, 101570, 101580, 101610, 101600, 
    101610, 101620, 101620, 101660, 101670, 101680, 101690, 101710, 101750, 
    101780, 101780, 101810, 101810, 101820, 101840, 101860, 101880, 101910, 
    101920, 101910, 101920, 101950, 101950, 101940, 101950, 101970, 102000, 
    102010, 102040, 102050, 102080, 102090, 102100, 102100, 102080, 102080, 
    102090, 102090, 102090, 102100, 102120, 102130, 102160, 102140, 102150, 
    102160, 102150, 102140, 102130, 102130, 102130, 102140, 102150, 102170, 
    102200, 102210, 102210, 102220, 102230, 102240, 102250, 102270, 102300, 
    102320, 102350, 102370, 102390, 102380, 102390, 102390, 102380, 102370, 
    102380, 102370, 102360, 102380, 102380, 102370, 102390, 102370, 102370, 
    102360, 102310, 102270, 102270, 102260, 102280, 102230, 102230, 102200, 
    102190, 102190, 102160, 102080, 102060, 101990, 101980, 101980, 101950, 
    101920, 101890, 101860, 101830, 101760, 101670, 101600, 101520, 101440, 
    101370, 101320, 101210, 101080, 101010, 100980, 100920, 100870, 100780, 
    100700, 100640, 100540, 100500, 100460, 100470, 100470, 100460, 100460, 
    100450, 100480, 100460, 100480, 100490, 100510, 100520, 100520, 100550, 
    100590, 100610, 100620, 100640, 100660, 100600, 100670, 100670, 100670, 
    100670, 100680, 100700, 100730, 100750, 100780, 100780, 100780, 100780, 
    100790, 100800, 100820, 100840, 100870, 100910, 100960, 101010, 101060, 
    101100, 101140, 101200, 101220, 101250, 101250, 101250, 101270, 101320, 
    101360, 101410, 101450, 101510, 101540, 101560, 101570, 101600, 101620, 
    101650, 101690, 101710, 101760, 101800, 101820, 101840, 101850, 101860, 
    101890, 101910, 101920, 101920, 101910, 101900, 101910, 101900, 101870, 
    101850, 101810, 101820, 101800, 101790, 101800, 101810, 101840, 101880, 
    101940, 101970, 102060, 102150, 102220, 102270, 102300, 102320, 102330, 
    102310, 102300, 102320, 102360, 102400, 102410, 102430, 102430, 102420, 
    102410, 102430, 102430, 102420, 102360, 102320, 102310, 102270, 102240, 
    102210, 102170, 102140, 102090, 102050, 102000, 101960, 101930, 101920, 
    101900, 101900, 101920, 101900, 101850, 101830, 101820, 101790, 101790, 
    101780, 101740, 101720, 101720, 101740, 101720, 101710, 101670, 101640, 
    101620, 101610, 101600, 101570, 101530, 101520, 101510, 101540, 101540, 
    101510, 101450, 101390, 101320, 101290, 101260, 101250, 101210, 101190, 
    101150, 101150, 101160, 101120, 101090, 101090, 101080, 101070, 101080, 
    101120, 101160, 101150, 101150, 101170, 101180, 101160, 101140, 101130, 
    101110, 101100, 101110, 101100, 101100, 101070, 101030, 101030, 101010, 
    100970, 100950, 100950, 100900, 100870, 100890, 100840, 100830, 100810, 
    100800, 100780, 100810, 100870, 100950, 101040, 101070, 101160, 101280, 
    101390, 101440, 101530, 101610, 101680, 101730, 101770, 101800, 101860, 
    101900, 101920, 101950, 102000, 102010, 102040, 102080, 102120, 102160, 
    102190, 102210, 102220, 102200, 102200, 102200, 102180, 102140, 102180, 
    102210, 102210, 102140, 102100, 102090, 102050, 102030, 101970, 101930, 
    101890, 101860, 101830, 101780, 101750, 101720, 101680, 101590, 101500, 
    101450, 101380, 101320, 101290, 101280, 101310, 101370, 101410, 101410, 
    101410, 101410, 101390, 101350, 101350, 101390, 101410, 101420, 101420, 
    101470, 101510, 101570, 101590, 101610, 101640, 101640, 101650, 101690, 
    101700, 101710, 101710, 101700, 101720, 101700, 101670, 101640, 101610, 
    101530, 101470, 101420, 101380, 101320, 101260, 101200, 101150, 101070, 
    101020, 100950, 100900, 100850, 100800, 100780, 100750, 100710, 100670, 
    100660, 100640, 100620, 100600, 100600, 100630, 100660, 100680, 100670, 
    100690, 100700, 100730, 100750, 100800, 100870, 100910, 100930, 100970, 
    101020, 101050, 101090, 101120, 101170, 101230, 101270, 101300, 101320, 
    101350, 101390, 101410, 101430, 101470, 101480, 101490, 101500, 101540, 
    101550, 101570, 101580, 101580, 101560, 101560, 101580, 101570, 101570, 
    101570, 101530, 101530, 101560, 101530, 101540, 101540, 101500, 101510, 
    101500, 101490, 101490, 101480, 101490, 101520, 101540, 101590, 101640, 
    101660, 101690, 101710, 101730, 101760, 101810, 101860, 101890, 101940, 
    102030, 102050, 102090, 102140, 102220, 102250, 102250, 102310, 102340, 
    102420, 102410, 102510, 102600, 102660, 102680, 102760, 102820, 102830, 
    102860, 102900, 102960, 103010, 103060, 103080, 103130, 103190, 103230, 
    103260, 103270, 103280, 103310, 103320, 103320, 103330, 103330, 103340, 
    103350, 103340, 103310, 103310, 103260, 103230, 103210, 103180, 103150, 
    103120, 103080, 103040, 103030, 103000, 102950, 102900, 102860, 102800, 
    102730, 102690, 102650, 102590, 102560, 102520, 102490, 102470, 102450, 
    102400, 102360, 102310, 102260, 102190, 102140, 102080, 102030, 101980, 
    101930, 101880, 101840, 101780, 101710, 101680, 101620, 101580, 101520, 
    101450, 101400, 101370, 101330, 101310, 101300, 101250, 101220, 101190, 
    101150, 101120, 101090, 101080, 101070, 101070, 101060, 101090, 101080, 
    101100, 101110, 101080, 101050, 101060, 101060, 101050, 101070, 101090, 
    101150, 101200, 101260, 101280, 101290, 101360, 101410, 101460, 101500, 
    101510, 101540, 101610, 101620, 101650, 101700, 101730, 101720, 101710, 
    101740, 101760, 101760, 101750, 101780, 101790, 101790, 101820, 101850, 
    101850, 101850, 101890, 101920, 101950, 101950, 101970, 102010, 101990, 
    102010, 102020, 102040, 102030, 102030, 102010, 102010, 101980, 101970, 
    101980, 101940, 101940, 101940, 101980, 102010, 102030, 102040, 102030, 
    102020, 101990, 101970, 101950, 101930, 101920, 101900, 101890, 101880, 
    101880, 101830, 101800, 101780, 101740, 101700, 101650, 101620, 101600, 
    101590, 101590, 101550, 101490, 101450, 101420, 101380, 101300, 101230, 
    101190, 101140, 101110, 101070, 101020, 100940, 100860, 100730, 100610, 
    100490, 100400, 100290, 100210, 100140, 100090, 100050, 100050, 100030, 
    100020, 100020, 100000, 99990, 99980, 99960, 99940, 99930, 99960, 99980, 
    100000, 100010, 100020, 100000, 100010, 100020, 100030, 100020, 100020, 
    100050, 100070, 100110, 100160, 100200, 100230, 100230, 100230, 100240, 
    100240, 100230, 100240, 100260, 100280, 100290, 100270, 100270, 100270, 
    100270, 100270, 100290, 100320, 100330, 100370, 100360, 100400, 100450, 
    100470, 100500, 100520, 100540, 100570, 100580, 100580, 100610, 100650, 
    100670, 100680, 100720, 100750, 100760, 100780, 100790, 100790, 100800, 
    100820, 100800, 100800, 100800, 100800, 100800, 100790, 100810, 100780, 
    100750, 100720, 100710, 100680, 100650, 100610, 100630, 100600, 100580, 
    100590, 100570, 100560, 100530, 100530, 100530, 100500, 100490, 100470, 
    100450, 100450, 100440, 100440, 100440, 100430, 100410, 100410, 100430, 
    100450, 100410, 100390, 100330, 100290, 100270, 100230, 100220, 100180, 
    100160, 100140, 100120, 100090, 100060, 100030, 100000, 99990, 99970, 
    99960, 99960, 99930, 99920, 99910, 99880, 99850, 99810, 99790, 99760, 
    99760, 99780, 99800, 99770, 99740, 99710, 99680, 99680, 99660, 99630, 
    99600, 99570, 99550, 99540, 99530, 99530, 99520, 99510, 99480, 99470, 
    99450, 99380, 99340, 99310, 99280, 99230, 99190, 99160, 99080, 99020, 
    99000, 98970, 98950, 98900, 98870, 98880, 98830, 98820, 98780, 98760, 
    98720, 98640, 98610, 98530, 98470, 98450, 98430, 98350, 98310, 98290, 
    98260, 98230, 98230, 98240, 98280, 98340, 98410, 98490, 98600, 98680, 
    98770, 98840, 98880, 98930, 98940, 98950, 98990, 99030, 99100, 99130, 
    99190, 99260, 99340, 99400, 99450, 99480, 99520, 99550, 99540, 99590, 
    99630, 99670, 99700, 99780, 99850, 99900, 100000, 100080, 100150, 100230, 
    100290, 100290, 100310, 100340, 100440, 100450, 100470, 100510, 100520, 
    100550, 100600, 100630, 100640, 100640, 100640, 100630, 100650, 100650, 
    100630, 100610, 100610, 100640, 100610, 100560, 100550, 100530, 100460, 
    100370, 100340, 100290, 100210, 100200, 100140, 100130, 100200, 100200, 
    100140, 100150, 100170, 100240, 100300, 100340, 100350, 100440, 100480, 
    100500, 100510, 100500, 100480, 100460, 100440, 100410, 100370, 100350, 
    100310, 100300, 100290, 100280, 100250, 100220, 100200, 100190, 100170, 
    100140, 100130, 100110, 100130, 100130, 100140, 100140, 100130, 100120, 
    100100, 100090, 100070, 100070, 100060, 100040, 100040, 100040, 100040, 
    100030, 100010, 99980, 99950, 99920, 99900, 99880, 99870, 99840, 99820, 
    99810, 99800, 99830, 99830, 99830, 99840, 99820, 99820, 99800, 99820, 
    99820, 99810, 99830, 99870, 99860, 99870, 99880, 99900, 99910, 99940, 
    99960, 100000, 100040, 100090, 100140, 100210, 100270, 100330, 100400, 
    100450, 100510, 100570, 100600, 100640, 100700, 100780, 100820, 100870, 
    100930, 100990, 101040, 101090, 101130, 101180, 101190, 101200, 101200, 
    101250, 101270, 101310, 101390, 101450, 101500, 101580, 101590, 101620, 
    101640, 101670, 101710, 101740, 101750, 101770, 101800, 101790, 101810, 
    101800, 101790, 101810, 101790, 101760, 101770, 101790, 101780, 101800, 
    101810, 101820, 101810, 101790, 101800, 101780, 101750, 101720, 101690, 
    101680, 101660, 101640, 101620, 101590, 101580, 101540, 101500, 101470, 
    101410, 101360, 101330, 101310, 101260, 101250, 101210, 101190, 101160, 
    101100, 101030, 101010, 100960, 100950, 100930, 100910, 100900, 100880, 
    100880, 100860, 100820, 100790, 100750, 100710, 100650, 100600, 100580, 
    100550, 100580, 100550, 100500, 100530, 100490, 100470, 100450, 100440, 
    100430, 100380, 100350, 100350, 100330, 100330, 100330, 100310, 100300, 
    100280, 100240, 100210, 100170, 100140, 100130, 100100, 100090, 100080, 
    100060, 100030, 100000, 99970, 99940, 99900, 99880, 99850, 99800, 99750, 
    99730, 99700, 99670, 99610, 99580, 99530, 99500, 99450, 99420, 99390, 
    99340, 99320, 99310, 99290, 99290, 99270, 99280, 99280, 99270, 99240, 
    99210, 99190, 99190, 99170, 99170, 99150, 99160, 99160, 99140, 99140, 
    99110, 99070, 99040, 99030, 99000, 98940, 98990, 98970, 98970, 98970, 
    98960, 98950, 98910, 98950, 98990, 99010, 99020, 99050, 99060, 99070, 
    99140, 99200, 99200, 99180, 99160, 99130, 99140, 99150, 99180, 99220, 
    99280, 99350, 99420, 99500, 99580, 99650, 99710, 99790, 99870, 99940, 
    100020, 100110, 100200, 100310, 100420, 100510, 100610, 100700, 100780, 
    100860, 100930, 100970, 101040, 101080, 101150, 101240, 101300, 101390, 
    101450, 101520, 101560, 101590, 101620, 101640, 101670, 101660, 101610, 
    101590, 101560, 101500, 101460, 101430, 101380, 101320, 101280, 101250, 
    101220, 101230, 101230, 101230, 101220, 101230, 101220, 101230, 101200, 
    101190, 101190, 101170, 101170, 101170, 101160, 101150, 101130, 101110, 
    101090, 101110, 101120, 101130, 101190, 101210, 101220, 101260, 101300, 
    101330, 101330, 101380, 101430, 101440, 101460, 101510, 101550, 101610, 
    101650, 101690, 101740, 101770, 101800, 101850, 101860, 101870, 101900, 
    101900, 101910, 101940, 101940, 101960, 102000, 102030, 102070, 102090, 
    102090, 102080, 102080, 102080, 102070, 102050, 102040, 101970, 101900, 
    101870, 101850, 101820, 101760, 101690, 101620, 101560, 101480, 101400, 
    101340, 101280, 101220, 101190, 101140, 101100, 101050, 100990, 100920, 
    100860, 100810, 100740, 100640, 100550, 100460, 100300, 100190, 100060, 
    99950, 99840, 99720, 99580, 99390, 99250, 99130, 99090, 99090, 99180, 
    99200, 99180, 99180, 99170, 99170, 99290, 99300, 99340, 99390, 99240, 
    99260, 99310, 99340, 99370, 99380, 99420, 99470, 99510, 99540, 99610, 
    99680, 99760, 99860, 99940, 100030, 100110, 100200, 100300, 100330, 
    100390, 100440, 100490, 100540, 100580, 100620, 100640, 100650, 100610, 
    100550, 100520, 100500, 100500, 100530, 100570, 100610, 100650, 100680, 
    100730, 100790, 100940, 100800, 100830, 100840, 100830, 100800, 100760, 
    100690, 100640, 100610, 100560, 100530, 100480, 100420, 100360, 100300, 
    100210, 100080, 99960, 99840, 99740, 99630, 99530, 99400, 99290, 99140, 
    98970, 98860, 98770, 98650, 98520, 98370, 98220, 98130, 98040, 97950, 
    97910, 97910, 97890, 97850, 97810, 97840, 97780, 97730, 97710, 97690, 
    97690, 97640, 97700, 97690, 97640, 97600, 97570, 97600, 97600, 97590, 
    97590, 97630, 97660, 97670, 97660, 97650, 97710, 97660, 97680, 97670, 
    97700, 97750, 97810, 97850, 97920, 97990, 98040, 98070, 98130, 98140, 
    98230, 98240, 98260, 98270, 98320, 98360, 98390, 98430, 98450, 98490, 
    98490, 98500, 98500, 98490, 98470, 98460, 98460, 98470, 98500, 98500, 
    98480, 98490, 98480, 98490, 98500, 98510, 98500, 98490, 98490, 98500, 
    98520, 98520, 98540, 98560, 98560, 98590, 98600, 98610, 98620, 98670, 
    98730, 98780, 98860, 98890, 98950, 98990, 99060, 99120, 99170, 99250, 
    99300, 99340, 99400, 99450, 99490, 99550, 99580, 99610, 99640, 99680, 
    99700, 99720, 99730, 99710, 99700, 99680, 99680, 99700, 99690, 99670, 
    99660, 99650, 99620, 99570, 99510, 99470, 99460, 99460, 99460, 99490, 
    99500, 99530, 99560, 99580, 99640, 99710, 99770, 99840, 99910, 100000, 
    100110, 100170, 100250, 100320, 100380, 100450, 100500, 100540, 100560, 
    100580, 100610, 100630, 100660, 100700, 100770, 100780, 100780, 100800, 
    100800, 100770, 100700, 100670, 100650, 100650, 100640, 100580, 100550, 
    100490, 100440, 100370, 100310, 100270, 100270, 100260, 100240, 100240, 
    100240, 100240, 100230, 100240, 100240, 100260, 100250, 100260, 100270, 
    100270, 100280, 100310, 100350, 100400, 100450, 100460, 100430, 100420, 
    100440, 100460, 100450, 100430, 100420, 100430, 100440, 100440, 100460, 
    100470, 100470, 100480, 100480, 100490, 100480, 100480, 100480, 100530, 
    100540, 100560, 100560, 100560, 100590, 100580, 100590, 100590, 100580, 
    100580, 100590, 100590, 100610, 100630, 100640, 100640, 100630, 100630, 
    100620, 100630, 100620, 100650, 100660, 100680, 100690, 100710, 100700, 
    100720, 100730, 100750, 100750, 100760, 100740, 100730, 100720, 100730, 
    100730, 100760, 100770, 100720, 100680, 100680, 100630, 100610, 100570, 
    100520, 100510, 100460, 100420, 100400, 100380, 100390, 100360, 100370, 
    100310, 100330, 100310, 100300, 100270, 100270, 100250, 100230, 100240, 
    100220, 100180, 100130, 100120, 100090, 100060, 100010, 100020, 100040, 
    100050, 100100, 100150, 100190, 100220, 100210, 100210, 100180, 100180, 
    100170, 100170, 100160, 100180, 100200, 100190, 100180, 100160, 100150, 
    100170, 100160, 100170, 100190, 100200, 100200, 100220, 100250, 100270, 
    100290, 100300, 100310, 100330, 100370, 100360, 100370, 100400, 100410, 
    100440, 100460, 100450, 100450, 100440, 100430, 100440, 100420, 100390, 
    100370, 100340, 100330, 100310, 100270, 100210, 100160, 100120, 100060, 
    100000, 99950, 99870, 99810, 99720, 99650, 99570, 99510, 99450, 99380, 
    99300, 99220, 99120, 99040, 98940, 98880, 98820, 98780, 98760, 98740, 
    98730, 98720, 98700, 98670, 98680, 98690, 98690, 98700, 98720, 98740, 
    98760, 98780, 98780, 98800, 98800, 98800, 98810, 98810, 98830, 98840, 
    98890, 98910, 98950, 98990, 99000, 99040, 99080, 99110, 99140, 99170, 
    99210, 99240, 99280, 99310, 99340, 99390, 99400, 99440, 99460, 99500, 
    99540, 99570, 99610, 99630, 99660, 99700, 99730, 99750, 99750, 99740, 
    99740, 99710, 99670, 99650, 99630, 99640, 99630, 99620, 99630, 99640, 
    99620, 99630, 99620, 99620, 99640, 99660, 99670, 99680, 99700, 99720, 
    99740, 99770, 99780, 99810, 99820, 99850, 99880, 99930, 99980, 100050, 
    100140, 100230, 100310, 100380, 100460, 100540, 100600, 100680, 100740, 
    100800, 100850, 100890, 100910, 100900, 100880, 100840, 100860, 100820, 
    100840, 100890, 100980, 101080, 101200, 101290, 101390, 101530, 101610, 
    101650, 101690, 101720, 101740, 101750, 101690, 101680, 101560, 101510, 
    101470, 101390, 101340, 101270, 101230, 101210, 101210, 101220, 101250, 
    101290, 101350, 101440, 101520, 101610, 101710, 101820, 101870, 101890, 
    102020, 102060, 102080, 102100, 102090, 102090, 102100, 102090, 102090, 
    102010, 101950, 101890, 101780, 101730, 101590, 101460, 101340, 101210, 
    101060, 100850, 100710, 100660, 100620, 100630, 100660, 100650, 100620, 
    100600, 100600, 100600, 100560, 100530, 100510, 100540, 100530, 100530, 
    100540, 100460, 100400, 100360, 100310, 100320, 100350, 100410, 100450, 
    100520, 100560, 100600, 100660, 100690, 100750, 100810, 100860, 100940, 
    100980, 101080, 101120, 101200, 101220, 101240, 101280, 101320, 101320, 
    101370, 101340, 101350, 101410, 101420, 101470, 101470, 101450, 101490, 
    101480, 101510, 101520, 101540, 101520, 101510, 101540, 101560, 101580, 
    101580, 101580, 101590, 101560, 101550, 101530, 101530, 101520, 101510, 
    101530, 101560, 101560, 101570, 101530, 101510, 101530, 101540, 101530, 
    101510, 101480, 101460, 101440, 101440, 101450, 101460, 101430, 101410, 
    101400, 101380, 101360, 101370, 101370, 101320, 101330, 101350, 101400, 
    101390, 101360, 101300, 101280, 101270, 101240, 101200, 101130, 101040, 
    100960, 100900, 100840, 100790, 100740, 100650, 100610, 100560, 100500, 
    100450, 100390, 100350, 100340, 100330, 100290, 100250, 100270, 100270, 
    100280, 100280, 100310, 100340, 100330, 100300, 100290, 100340, 100360, 
    100400, 100410, 100410, 100430, 100450, 100470, 100480, 100500, 100500, 
    100500, 100510, 100540, 100580, 100600, 100600, 100570, 100570, 100580, 
    100590, 100580, 100580, 100570, 100580, 100600, 100600, 100580, 100580, 
    100570, 100560, 100560, 100540, 100510, 100450, 100430, 100400, 100370, 
    100350, 100320, 100290, 100230, 100200, 100150, 100070, 100020, 99950, 
    99880, 99810, 99750, 99670, 99580, 99510, 99440, 99400, 99390, 99370, 
    99360, 99370, 99400, 99410, 99440, 99500, 99520, 99540, 99590, 99640, 
    99670, 99700, 99700, 99720, 99740, 99800, 99830, 99870, 99910, 99950, 
    99990, 100020, 100060, 100100, 100120, 100160, 100200, 100240, 100270, 
    100320, 100360, 100420, 100450, 100480, 100520, 100580, 100610, 100650, 
    100670, 100740, 100780, 100860, 100930, 100990, 101030, 101080, 101110, 
    101150, 101180, 101220, 101250, 101290, 101350, 101390, 101470, 101510, 
    101570, 101610, 101640, 101650, 101680, 101710, 101750, 101800, 101850, 
    101880, 101890, 101920, 101960, 101980, 101990, 101990, 102010, 102000, 
    102010, 102010, 102030, 102050, 102060, 102080, 102030, 102000, 101990, 
    101990, 101960, 101940, 101930, 101950, 101950, 101930, 101940, 101940, 
    101920, 101910, 101880, 101830, 101770, 101740, 101660, 101620, 101580, 
    101530, 101470, 101450, 101430, 101400, 101360, 101310, 101270, 101240, 
    101190, 101140, 101120, 101080, 101040, 100970, 100900, 100830, 100740, 
    100670, 100580, 100500, 100430, 100380, 100310, 100230, 100120, 100020, 
    99940, 99840, 99770, 99680, 99600, 99520, 99450, 99390, 99330, 99290, 
    99250, 99180, 99160, 99140, 99130, 99140, 99130, 99140, 99180, 99210, 
    99230, 99250, 99250, 99280, 99280, 99270, 99240, 99190, 99140, 99110, 
    99110, 99120, 99100, 99110, 99110, 99130, 99160, 99190, 99230, 99280, 
    99310, 99360, 99390, 99430, 99470, 99480, 99510, 99520, 99520, 99540, 
    99560, 99570, 99590, 99600, 99630, 99640, 99690, 99730, 99770, 99810, 
    99830, 99870, 99860, 99890, 99950, 99970, 100000, 100030, 100070, 100110, 
    100130, 100110, 100080, 100070, 100100, 100090, 100100, 100080, 100070, 
    100070, 100070, 100070, 100060, 100070, 100070, 100050, 100050, 100040, 
    100040, 100030, 100040, 100060, 100090, 100090, 100090, 100080, 100120, 
    100130, 100150, 100180, 100220, 100240, 100240, 100270, 100300, 100310, 
    100300, 100340, 100350, 100360, 100360, 100380, 100390, 100410, 100440, 
    100470, 100490, 100480, 100500, 100540, 100570, 100600, 100630, 100650, 
    100680, 100700, 100690, 100680, 100690, 100720, 100750, 100730, 100670, 
    100680, 100660, 100670, 100660, 100660, 100650, 100630, 100600, 100580, 
    100550, 100490, 100440, 100360, 100280, 100190, 100080, 99960, 99830, 
    99720, 99600, 99460, 99290, 99170, 98980, 98830, 98670, 98580, 98460, 
    98340, 98210, 98090, 98000, 97870, 97750, 97660, 97540, 97380, 97320, 
    97270, 97290, 97310, 97360, 97400, 97450, 97510, 97550, 97610, 97610, 
    97770, 97840, 97900, 97990, 98070, 98180, 98270, 98370, 98440, 98510, 
    98620, 98710, 98780, 98850, 98910, 98980, 99020, 99080, 99130, 99190, 
    99240, 99260, 99270, 99290, 99300, 99300, 99300, 99270, 99230, 99180, 
    99140, 99100, 99090, 99060, 99020, 98980, 98950, 98920, 98870, 98860, 
    98880, 98900, 98910, 98930, 98980, 99030, 99100, 99180, 99270, 99360, 
    99440, 99530, 99640, 99760, 99860, 99970, 100060, 100190, 100300, 100400, 
    100490, 100600, 100670, 100700, 100700, 100720, 100730, 100730, 100730, 
    100700, 100660, 100640, 100620, 100550, 100470, 100420, 100370, 100340, 
    100340, 100350, 100330, 100360, 100380, 100410, 100410, 100360, 100350, 
    100320, 100290, 100240, 100200, 100160, 100110, 100060, 100000, 99940, 
    99880, 99830, 99770, 99760, 99780, 99800, 99870, 99940, 100050, 100150, 
    100260, 100310, 100430, 100530, 100630, 100770, 100890, 100970, 101110, 
    101210, 101310, 101400, 101490, 101560, 101630, 101680, 101700, 101740, 
    101750, 101770, 101810, 101830, 101830, 101840, 101840, 101840, 101850, 
    101840, 101850, 101830, 101790, 101790, 101790, 101780, 101750, 101700, 
    101690, 101650, 101640, 101590, 101510, 101520, 101520, 101520, 101540, 
    101560, 101570, 101600, 101630, 101680, 101700, 101740, 101810, 101860, 
    101910, 101950, 102030, 102080, 102110, 102160, 102230, 102280, 102320, 
    102340, 102350, 102380, 102390, 102400, 102430, 102460, 102460, 102450, 
    102440, 102430, 102410, 102380, 102360, 102320, 102320, 102310, 102280, 
    102260, 102260, 102250, 102230, 102200, 102180, 102160, 102150, 102120, 
    102110, 102120, 102140, 102150, 102150, 102150, 102160, 102160, 102160, 
    102150, 102150, 102150, 102150, 102160, 102160, 102150, 102130, 102130, 
    102110, 102120, 102100, 102020, 101980, 102020, 102000, 101990, 101970, 
    101950, 101920, 101880, 101840, 101800, 101760, 101730, 101690, 101610, 
    101600, 101570, 101540, 101520, 101520, 101500, 101510, 101520, 101500, 
    101490, 101490, 101490, 101510, 101530, 101560, 101610, 101660, 101690, 
    101740, 101760, 101780, 101800, 101840, 101860, 101910, 101970, 102020, 
    102050, 102110, 102130, 102180, 102250, 102280, 102310, 102320, 102330, 
    102350, 102380, 102400, 102390, 102400, 102400, 102390, 102360, 102330, 
    102280, 102220, 102180, 102110, 102060, 102030, 102000, 101990, 102000, 
    102010, 102000, 101980, 102000, 101990, 101970, 101970, 101970, 102000, 
    102020, 101990, 101960, 101940, 101940, 101920, 101910, 101890, 101880, 
    101880, 101880, 101890, 101880, 101880, 101860, 101870, 101860, 101840, 
    101830, 101810, 101790, 101770, 101760, 101750, 101740, 101750, 101700, 
    101690, 101690, 101670, 101650, 101670, 101670, 101670, 101690, 101680, 
    101700, 101690, 101720, 101710, 101710, 101730, 101750, 101790, 101800, 
    101810, 101830, 101880, 101900, 101930, 101950, 101970, 102000, 102020, 
    102050, 102080, 102100, 102130, 102140, 102180, 102220, 102220, 102260, 
    102280, 102300, 102320, 102320, 102340, 102350, 102360, 102370, 102380, 
    102390, 102400, 102420, 102420, 102410, 102400, 102410, 102380, 102380, 
    102360, 102350, 102360, 102360, 102350, 102330, 102310, 102290, 102290, 
    102260, 102230, 102230, 102210, 102200, 102190, 102180, 102160, 102150, 
    102130, 102120, 102110, 102080, 102070, 102060, 102070, 102070, 102060, 
    102060, 102070, 102090, 102090, 102100, 102110, 102120, 102130, 102130, 
    102150, 102140, 102140, 102170, 102190, 102190, 102190, 102170, 102160, 
    102180, 102170, 102160, 102180, 102180, 102180, 102200, 102190, 102200, 
    102200, 102200, 102200, 102230, 102240, 102230, 102220, 102220, 102220, 
    102220, 102240, 102270, 102290, 102340, 102350, 102370, 102400, 102430, 
    102450, 102470, 102490, 102490, 102520, 102550, 102550, 102530, 102510, 
    102520, 102540, 102560, 102560, 102560, 102560, 102540, 102530, 102480, 
    102450, 102420, 102410, 102360, 102310, 102280, 102240, 102200, 102170, 
    102140, 102110, 102080, 102030, 101990, 101950, 101900, 101860, 101810, 
    101750, 101690, 101620, 101540, 101490, 101410, 101330, 101290, 101240, 
    101210, 101180, 101150, 101160, 101230, 101250, 101290, 101320, 101340, 
    101350, 101350, 101330, 101300, 101300, 101280, 101250, 101220, 101170, 
    101130, 101080, 101050, 100990, 100950, 100890, 100830, 100780, 100760, 
    100740, 100730, 100710, 100690, 100680, 100680, 100670, 100650, 100630, 
    100610, 100600, 100590, 100600, 100600, 100620, 100610, 100630, 100620, 
    100630, 100630, 100630, 100620, 100600, 100610, 100610, 100630, 100650, 
    100640, 100620, 100610, 100600, 100560, 100570, 100580, 100580, 100580, 
    100590, 100610, 100600, 100610, 100600, 100610, 100610, 100620, 100600, 
    100590, 100560, 100560, 100560, 100570, 100570, 100560, 100530, 100540, 
    100530, 100530, 100530, 100510, 100500, 100490, 100500, 100510, 100540, 
    100540, 100560, 100560, 100580, 100580, 100580, 100580, 100590, 100590, 
    100590, 100620, 100640, 100660, 100690, 100720, 100730, 100760, 100760, 
    100770, 100790, 100790, 100810, 100830, 100860, 100880, 100890, 100890, 
    100900, 100890, 100890, 100880, 100850, 100860, 100860, 100860, 100860, 
    100870, 100890, 100900, 100900, 100910, 100900, 100910, 100920, 100940, 
    100970, 100990, 101010, 101040, 101050, 101060, 101080, 101080, 101100, 
    101120, 101110, 101130, 101140, 101160, 101190, 101220, 101240, 101270, 
    101270, 101280, 101290, 101300, 101300, 101320, 101330, 101340, 101360, 
    101360, 101380, 101390, 101380, 101380, 101360, 101350, 101360, 101340, 
    101330, 101330, 101330, 101310, 101300, 101290, 101310, 101300, 101280, 
    101220, 101190, 101130, 101100, 101030, 100990, 100950, 100890, 100830, 
    100830, 100800, 100790, 100770, 100730, 100700, 100670, 100640, 100590, 
    100550, 100500, 100450, 100390, 100310, 100210, 100100, 99990, 99880, 
    99790, 99690, 99590, 99510, 99440, 99400, 99360, 99340, 99300, 99270, 
    99200, 99260, 99280, 99390, 99520, 99580, 99580, 99610, 99680, 99690, 
    99670, 99710, 99720, 99760, 99770, 99790, 99820, 99870, 99930, 99970, 
    100040, 100100, 100170, 100260, 100330, 100380, 100460, 100560, 100650, 
    100730, 100800, 100870, 100950, 101010, 101060, 101090, 101140, 101180, 
    101220, 101290, 101340, 101390, 101410, 101440, 101450, 101460, 101470, 
    101450, 101430, 101410, 101400, 101400, 101370, 101360, 101340, 101310, 
    101280, 101260, 101230, 101200, 101160, 101140, 101130, 101130, 101110, 
    101110, 101110, 101130, 101110, 101110, 101090, 101060, 101040, 101030, 
    101030, 101040, 101050, 101030, 101010, 101010, 101010, 100990, 100960, 
    100980, 101010, 100990, 100970, 100980, 100980, 100950, 100910, 100850, 
    100820, 100780, 100780, 100740, 100680, 100620, 100580, 100580, 100570, 
    100570, 100630, 100650, 100700, 100760, 100820, 100860, 100900, 100970, 
    101030, 101100, 101170, 101240, 101310, 101360, 101430, 101460, 101500, 
    101520, 101570, 101590, 101630, 101660, 101720, 101760, 101820, 101870, 
    101900, 101950, 101970, 101990, 102020, 102040, 102070, 102120, 102160, 
    102210, 102260, 102270, 102300, 102330, 102340, 102370, 102340, 102370, 
    102380, 102400, 102400, 102430, 102470, 102490, 102500, 102490, 102500, 
    102490, 102470, 102450, 102430, 102430, 102430, 102440, 102430, 102420, 
    102420, 102420, 102400, 102400, 102400, 102410, 102420, 102440, 102460, 
    102490, 102500, 102510, 102530, 102560, 102590, 102620, 102640, 102660, 
    102680, 102710, 102740, 102780, 102830, 102870, 102900, 102940, 102970, 
    102990, 103000, 103030, 103050, 103080, 103100, 103130, 103150, 103170, 
    103210, 103230, 103230, 103230, 103260, 103250, 103250, 103260, 103290, 
    103290, 103320, 103350, 103340, 103330, 103360, 103350, 103340, 103340, 
    103350, 103360, 103350, 103360, 103370, 103350, 103350, 103340, 103340, 
    103300, 103260, 103240, 103210, 103180, 103160, 103140, 103120, 103080, 
    103060, 103060, 103040, 103020, 103010, 102980, 102950, 102940, 102940, 
    102940, 102910, 102940, 102900, 102870, 102820, 102760, 102710, 102660, 
    102610, 102560, 102570, 102600, 102600, 102590, 102600, 102590, 102570, 
    102580, 102560, 102550, 102540, 102530, 102480, 102450, 102420, 102400, 
    102370, 102360, 102310, 102260, 102210, 102190, 102170, 102150, 102150, 
    102130, 102110, 102120, 102130, 102100, 102090, 102080, 102070, 102090, 
    102090, 102110, 102150, 102180, 102180, 102190, 102190, 102180, 102130, 
    102120, 102110, 102080, 102060, 102040, 102020, 102000, 101960, 101950, 
    101920, 101880, 101870, 101850, 101820, 101780, 101780, 101770, 101760, 
    101740, 101720, 101700, 101650, 101630, 101580, 101550, 101510, 101450, 
    101420, 101390, 101380, 101350, 101330, 101310, 101310, 101290, 101270, 
    101250, 101250, 101270, 101280, 101270, 101290, 101290, 101290, 101300, 
    101290, 101300, 101310, 101320, 101330, 101330, 101310, 101320, 101350, 
    101360, 101370, 101380, 101400, 101390, 101410, 101410, 101420, 101420, 
    101440, 101450, 101510, 101550, 101560, 101590, 101610, 101630, 101650, 
    101640, 101650, 101640, 101670, 101680, 101690, 101700, 101700, 101700, 
    101710, 101710, 101720, 101690, 101690, 101670, 101650, 101640, 101640, 
    101660, 101610, 101590, 101550, 101530, 101500, 101470, 101440, 101420, 
    101410, 101380, 101360, 101350, 101330, 101290, 101260, 101250, 101250, 
    101240, 101230, 101240, 101280, 101320, 101390, 101420, 101470, 101510, 
    101570, 101620, 101670, 101710, 101760, 101810, 101860, 101890, 101930, 
    101980, 102050, 102070, 102120, 102160, 102180, 102200, 102210, 102250, 
    102290, 102330, 102360, 102380, 102400, 102430, 102440, 102440, 102440, 
    102440, 102420, 102400, 102370, 102360, 102360, 102340, 102320, 102320, 
    102300, 102270, 102260, 102230, 102190, 102170, 102140, 102110, 102080, 
    102040, 102030, 102010, 101990, 101970, 101940, 101910, 101910, 101880, 
    101850, 101820, 101820, 101810, 101810, 101780, 101780, 101760, 101730, 
    101740, 101710, 101700, 101700, 101680, 101680, 101690, 101670, 101650, 
    101660, 101680, 101680, 101670, 101640, 101640, 101630, 101640, 101660, 
    101680, 101690, 101690, 101710, 101720, 101720, 101730, 101730, 101730, 
    101720, 101740, 101730, 101730, 101710, 101710, 101690, 101670, 101630, 
    101620, 101610, 101560, 101540, 101530, 101520, 101500, 101470, 101460, 
    101460, 101460, 101450, 101430, 101440, 101410, 101420, 101400, 101400, 
    101430, 101440, 101450, 101470, 101500, 101510, 101540, 101540, 101550, 
    101580, 101610, 101630, 101690, 101740, 101770, 101780, 101800, 101830, 
    101870, 101880, 101910, 101920, 101960, 101990, 102020, 102040, 102050, 
    102060, 102070, 102080, 102090, 102080, 102070, 102060, 102050, 102050, 
    102070, 102030, 102000, 101970, 101930, 101930, 101890, 101840, 101810, 
    101760, 101730, 101700, 101650, 101630, 101600, 101560, 101540, 101520, 
    101510, 101470, 101430, 101420, 101420, 101440, 101460, 101450, 101460, 
    101450, 101460, 101470, 101450, 101450, 101430, 101440, 101440, 101450, 
    101460, 101460, 101430, 101420, 101410, 101400, 101380, 101350, 101330, 
    101290, 101280, 101290, 101270, 101270, 101260, 101250, 101220, 101210, 
    101220, 101230, 101230, 101230, 101260, 101280, 101300, 101320, 101340, 
    101360, 101370, 101390, 101380, 101400, 101420, 101440, 101460, 101480, 
    101520, 101500, 101500, 101500, 101510, 101500, 101500, 101480, 101460, 
    101430, 101400, 101370, 101350, 101280, 101240, 101210, 101150, 101090, 
    101020, 101000, 100950, 100880, 100840, 100790, 100770, 100710, 100650, 
    100610, 100590, 100530, 100510, 100490, 100480, 100460, 100440, 100420, 
    100360, 100280, 100240, 100190, 100220, 100300, 100320, 100370, 100350, 
    100320, 100290, 100300, 100290, 100360, 100410, 100440, 100450, 100480, 
    100510, 100580, 100620, 100630, 100720, 100780, 100830, 100890, 100940, 
    101010, 101010, 101090, 101140, 101180, 101200, 101240, 101280, 101360, 
    101370, 101460, 101420, 101450, 101470, 101500, 101480, 101470, 101460, 
    101450, 101420, 101390, 101360, 101320, 101280, 101230, 101180, 101130, 
    101060, 101010, 100970, 100930, 100850, 100780, 100740, 100680, 100640, 
    100590, 100560, 100550, 100530, 100510, 100510, 100520, 100520, 100540, 
    100560, 100610, 100630, 100660, 100700, 100740, 100780, 100780, 100800, 
    100800, 100800, 100800, 100830, 100850, 100870, 100890, 100920, 100940, 
    100960, 100960, 100990, 101000, 101030, 101030, 101030, 101060, 101100, 
    101150, 101180, 101230, 101240, 101260, 101240, 101260, 101260, 101260, 
    101250, 101250, 101280, 101250, 101230, 101240, 101260, 101240, 101240, 
    101230, 101230, 101230, 101230, 101260, 101280, 101300, 101330, 101360, 
    101380, 101400, 101460, 101460, 101510, 101550, 101560, 101590, 101610, 
    101660, 101690, 101690, 101690, 101720, 101750, 101750, 101760, 101780, 
    101810, 101800, 101820, 101820, 101830, 101810, 101810, 101790, 101780, 
    101770, 101770, 101770, 101760, 101740, 101740, 101720, 101700, 101690, 
    101670, 101650, 101650, 101650, 101650, 101650, 101630, 101620, 101640, 
    101640, 101650, 101660, 101660, 101660, 101680, 101700, 101710, 101730, 
    101750, 101770, 101790, 101810, 101850, 101870, 101900, 101930, 101950, 
    101980, 102020, 102040, 102080, 102100, 102110, 102140, 102140, 102150, 
    102150, 102160, 102160, 102180, 102210, 102230, 102220, 102230, 102240, 
    102250, 102260, 102250, 102260, 102260, 102280, 102290, 102310, 102320, 
    102330, 102330, 102350, 102340, 102360, 102340, 102340, 102340, 102330, 
    102340, 102340, 102340, 102340, 102340, 102340, 102340, 102340, 102340, 
    102340, 102330, 102330, 102330, 102350, 102370, 102370, 102370, 102360, 
    102360, 102360, 102340, 102320, 102330, 102330, 102320, 102300, 102280, 
    102270, 102260, 102230, 102220, 102190, 102190, 102170, 102140, 102110, 
    102090, 102090, 102060, 102040, 102020, 102000, 101990, 101970, 101970, 
    101940, 101920, 101900, 101900, 101850, 101820, 101810, 101780, 101760, 
    101740, 101720, 101700, 101700, 101670, 101650, 101620, 101610, 101600, 
    101570, 101550, 101540, 101550, 101550, 101550, 101550, 101550, 101550, 
    101540, 101540, 101540, 101530, 101530, 101530, 101520, 101530, 101550, 
    101530, 101550, 101540, 101560, 101560, 101560, 101570, 101590, 101590, 
    101590, 101580, 101570, 101580, 101570, 101560, 101560, 101580, 101580, 
    101580, 101590, 101580, 101580, 101580, 101570, 101580, 101580, 101580, 
    101570, 101570, 101570, 101570, 101560, 101560, 101540, 101530, 101500, 
    101480, 101430, 101400, 101370, 101350, 101320, 101300, 101270, 101230, 
    101190, 101170, 101150, 101120, 101090, 101050, 101020, 101000, 100980, 
    100940, 100920, 100920, 100910, 100890, 100860, 100830, 100810, 100800, 
    100790, 100770, 100750, 100740, 100720, 100710, 100680, 100660, 100650, 
    100650, 100620, 100600, 100610, 100610, 100620, 100610, 100610, 100610, 
    100620, 100640, 100650, 100650, 100640, 100620, 100630, 100640, 100660, 
    100660, 100670, 100680, 100690, 100710, 100710, 100740, 100760, 100780, 
    100800, 100820, 100850, 100870, 100880, 100920, 100950, 100970, 100990, 
    101030, 101070, 101110, 101130, 101190, 101240, 101270, 101310, 101340, 
    101340, 101360, 101420, 101460, 101480, 101470, 101500, 101500, 101540, 
    101540, 101570, 101590, 101600, 101610, 101610, 101600, 101600, 101600, 
    101580, 101590, 101580, 101570, 101570, 101560, 101550, 101520, 101510, 
    101490, 101490, 101470, 101460, 101480, 101510, 101510, 101530, 101530, 
    101540, 101540, 101540, 101550, 101530, 101540, 101530, 101510, 101510, 
    101530, 101520, 101500, 101490, 101480, 101490, 101460, 101450, 101450, 
    101450, 101460, 101450, 101480, 101500, 101520, 101520, 101530, 101540, 
    101540, 101560, 101560, 101550, 101570, 101600, 101620, 101630, 101660, 
    101670, 101690, 101710, 101700, 101700, 101700, 101700, 101730, 101750, 
    101760, 101780, 101800, 101780, 101790, 101790, 101790, 101780, 101780, 
    101780, 101780, 101810, 101810, 101810, 101810, 101800, 101780, 101800, 
    101810, 101770, 101780, 101770, 101760, 101750, 101770, 101770, 101790, 
    101800, 101800, 101810, 101820, 101830, 101840, 101860, 101880, 101900, 
    101920, 101980, 102010, 102040, 102050, 102080, 102110, 102140, 102160, 
    102210, 102250, 102290, 102340, 102370, 102380, 102410, 102410, 102410, 
    102430, 102430, 102440, 102450, 102460, 102470, 102490, 102510, 102530, 
    102550, 102580, 102600, 102600, 102600, 102590, 102600, 102630, 102650, 
    102680, 102710, 102690, 102700, 102710, 102700, 102710, 102700, 102690, 
    102680, 102680, 102670, 102710, 102700, 102690, 102690, 102660, 102630, 
    102580, 102560, 102510, 102480, 102420, 102390, 102360, 102340, 102300, 
    102270, 102240, 102180, 102140, 102120, 102070, 102060, 102020, 101990, 
    102000, 101930, 101870, 101840, 101780, 101700, 101630, 101550, 101490, 
    101420, 101350, 101300, 101210, 101130, 101060, 101020, 100980, 100950, 
    100910, 100870, 100830, 100810, 100810, 100800, 100830, 100850, 100860, 
    100910, 100920, 100920, 100940, 100940, 100950, 100950, 100930, 100930, 
    100930, 100880, 100850, 100800, 100760, 100700, 100650, 100620, 100580, 
    100550, 100510, 100490, 100470, 100500, 100500, 100530, 100580, 100600, 
    100650, 100690, 100690, 100760, 100800, 100850, 100920, 100960, 101030, 
    101040, 101080, 101120, 101160, 101180, 101220, 101230, 101270, 101300, 
    101350, 101380, 101430, 101460, 101490, 101520, 101540, 101540, 101540, 
    101550, 101570, 101590, 101620, 101660, 101670, 101670, 101700, 101700, 
    101710, 101720, 101710, 101720, 101750, 101770, 101780, 101790, 101830, 
    101850, 101850, 101860, 101860, 101850, 101860, 101850, 101840, 101840, 
    101860, 101890, 101910, 101920, 101930, 101920, 101900, 101910, 101900, 
    101910, 101920, 101930, 101940, 101970, 101980, 102000, 102000, 102030, 
    102040, 102040, 102040, 102040, 102030, 102050, 102070, 102090, 102110, 
    102100, 102100, 102100, 102090, 102080, 102060, 102050, 102060, 102060, 
    102050, 102050, 102040, 102050, 102030, 101980, 101950, 101880, 101810, 
    101770, 101730, 101720, 101710, 101660, 101600, 101580, 101570, 101540, 
    101490, 101430, 101380, 101370, 101340, 101300, 101280, 101250, 101230, 
    101230, 101250, 101240, 101210, 101210, 101180, 101190, 101190, 101190, 
    101200, 101200, 101220, 101220, 101240, 101230, 101220, 101230, 101230, 
    101230, 101240, 101270, 101300, 101330, 101340, 101370, 101380, 101400, 
    101430, 101460, 101460, 101480, 101510, 101540, 101580, 101600, 101630, 
    101620, 101620, 101620, 101620, 101630, 101650, 101650, 101670, 101700, 
    101750, 101760, 101770, 101800, 101830, 101850, 101850, 101850, 101850, 
    101870, 101850, 101850, 101850, 101800, 101780, 101750, 101720, 101640, 
    101570, 101490, 101470, 101460, 101470, 101490, 101510, 101500, 101470, 
    101470, 101460, 101430, 101420, 101380, 101360, 101320, 101300, 101310, 
    101320, 101310, 101320, 101330, 101350, 101360, 101360, 101380, 101400, 
    101410, 101430, 101470, 101480, 101500, 101500, 101470, 101460, 101450, 
    101450, 101420, 101380, 101380, 101360, 101350, 101350, 101350, 101370, 
    101370, 101390, 101380, 101410, 101450, 101470, 101490, 101530, 101570, 
    101620, 101650, 101670, 101690, 101720, 101760, 101790, 101810, 101820, 
    101850, 101870, 101890, 101910, 101930, 101940, 101930, 101910, 101870, 
    101830, 101780, 101750, 101690, 101660, 101620, 101570, 101520, 101460, 
    101410, 101350, 101300, 101240, 101180, 101110, 101090, 101050, 101020, 
    100970, 100920, 100890, 100840, 100810, 100780, 100760, 100740, 100730, 
    100720, 100690, 100690, 100680, 100660, 100640, 100640, 100600, 100560, 
    100520, 100460, 100400, 100360, 100360, 100350, 100340, 100310, 100290, 
    100300, 100310, 100300, 100300, 100340, 100340, 100380, 100390, 100460, 
    100520, 100570, 100620, 100680, 100760, 100830, 100890, 100940, 100980, 
    101000, 101050, 101070, 101080, 101070, 101110, 101090, 101070, 101040, 
    101010, 101000, 100970, 100940, 100930, 100910, 100880, 100860, 100840, 
    100830, 100820, 100800, 100780, 100770, 100760, 100740, 100730, 100730, 
    100740, 100750, 100750, 100760, 100780, 100790, 100810, 100810, 100800, 
    100800, 100810, 100850, 100870, 100890, 100910, 100920, 100930, 100910, 
    100930, 100930, 100930, 100930, 100940, 100950, 100970, 100980, 101010, 
    101040, 101050, 101030, 101010, 101010, 101020, 101030, 101020, 101040, 
    101030, 101040, 101030, 101020, 101020, 101010, 101010, 101010, 101010, 
    101020, 101040, 101060, 101080, 101110, 101140, 101150, 101170, 101170, 
    101170, 101190, 101210, 101220, 101230, 101250, 101270, 101300, 101310, 
    101320, 101340, 101330, 101330, 101330, 101320, 101320, 101340, 101350, 
    101360, 101360, 101380, 101360, 101360, 101350, 101330, 101330, 101300, 
    101290, 101280, 101290, 101290, 101290, 101290, 101300, 101270, 101270, 
    101260, 101250, 101240, 101230, 101210, 101220, 101200, 101190, 101180, 
    101140, 101100, 101060, 101030, 100990, 100960, 100880, 100810, 100770, 
    100750, 100720, 100690, 100670, 100630, 100590, 100560, 100500, 100450, 
    100400, 100360, 100310, 100270, 100240, 100190, 100150, 100120, 100080, 
    100030, 100000, 99980, 99930, 99910, 99890, 99870, 99850, 99860, 99860, 
    99880, 99850, 99840, 99830, 99830, 99850, 99850, 99860, 99870, 99880, 
    99890, 99920, 99930, 99950, 99960, 99970, 99980, 100000, 100020, 100050, 
    100060, 100080, 100120, 100140, 100160, 100180, 100220, 100230, 100270, 
    100300, 100310, 100380, 100430, 100480, 100500, 100560, 100650, 100700, 
    100750, 100790, 100840, 100870, 100920, 100960, 101000, 101050, 101100, 
    101130, 101140, 101140, 101150, 101140, 101140, 101140, 101130, 101140, 
    101180, 101210, 101220, 101230, 101240, 101260, 101270, 101280, 101280, 
    101230, 101250, 101270, 101300, 101330, 101350, 101370, 101380, 101400, 
    101400, 101400, 101400, 101490, 101500, 101460, 101460, 101510, 101460, 
    101450, 101520, 101540, 101530, 101530, 101530, 101550, 101570, 101590, 
    101610, 101640, 101680, 101700, 101710, 101720, 101730, 101750, 101760, 
    101800, 101820, 101720, 101740, 101750, 101790, 101800, 101810, 101810, 
    101790, 101780, 101790, 101790, 101770, 101770, 101780, 101790, 101790, 
    101760, 101760, 101760, 101760, 101740, 101730, 101720, 101710, 101710, 
    101730, 101740, 101760, 101750, 101720, 101710, 101670, 101640, 101610, 
    101600, 101630, 101660, 101670, 101690, 101700, 101720, 101730, 101740, 
    101740, 101750, 101780, 101820, 101860, 101890, 101920, 101940, 101970, 
    101970, 101970, 101970, 101970, 101960, 101940, 101920, 101910, 101930, 
    101920, 101910, 101900, 101970, 101960, 101830, 101800, 101770, 101740, 
    101720, 101710, 101710, 101700, 101680, 101650, 101630, 101610, 101600, 
    101580, 101560, 101540, 101540, 101540, 101550, 101540, 101530, 101540, 
    101540, 101560, 101570, 101590, 101640, 101630, 101650, 101680, 101700, 
    _, _, _, _, _, _, _, _, _, _, _, 101960, 101980, 102000, 102020, 102000, 
    101970, 101960, 101950, 101940, 101930, 101910, 101900, 101870, 101870, 
    101850, 101820, 101810, 101790, 101770, 101730, 101680, 101650, 101620, 
    101600, 101600, 101590, 101590, 101590, 101590, 101530, 101520, 101500, 
    101480, 101460, 101460, 101450, 101430, 101420, 101370, 101350, 101340, 
    101350, 101320, 101290, 101260, 101230, 101220, 101220, 101200, 101190, 
    101190, 101180, 101160, 101120, 101090, 101080, 101070, 101040, 101040, 
    101030, 101020, 101010, 101030, 101000, 100970, 100970, 100960, 100940, 
    100920, 100890, 100890, 100880, 100890, 100890, 100870, 100830, _, _, _, 
    _, _, _, _, _, 100680, 100680, 100640, 100640, 100620, 100600, 100580, 
    100570, 100550, 100550, 100540, 100540, 100540, 100520, 100550, 100550, 
    100550, 100550, 100560, 100570, 100570, 100560, 100560, 100560, 100580, 
    100580, 100580, 100580, 100580, 100570, 100570, 100590, 100600, 100610, 
    100610, 100630, 100660, 100660, 100650, 100650, 100630, 100630, 100630, 
    100640, 100640, 100650, 100660, 100670, 100670, 100700, 100720, 100730, 
    100740, 100740, 100760, 100770, 100790, 100810, 100840, 100860, 100880, 
    100890, 100880, 100900, 100930, 100920, 100960, 100990, 101010, 101040, 
    101050, 101050, 101030, 101030, 101030, 101060, 101060, 101040, 101020, 
    101020, 101010, 100990, 101000, 101000, 101000, 101030, 101030, 101010, 
    101050, 101020, 101000, 101000, 100960, 100930, 100910, 100920, 100910, 
    100880, 100870, 100840, 100830, 100830, 100830, 100830, 100840, 100810, 
    100810, 100800, 100800, 100790, 100790, 100780, 100750, 100730, 100730, 
    100720, 100700, 100700, 100660, 100650, 100650, 100640, 100670, 100670, 
    100650, 100640, 100630, 100610, 100610, _, 100680, _, _, _, _, 100790, _, 
    100730, 100740, 100750, 100770, 100800, 100830, 100860, 100890, 100910, 
    100930, 100960, 101000, 101020, 101060, 101060, 101060, 101110, 101170, 
    101200, _, _, _, 101430, _, 101340, 101340, 101330, 101330, 101320, 
    101320, 101320, 101310, 101310, 101290, 101280, 101250, 101230, 101240, 
    101220, 101200, 101160, 101160, 101170, 101170, 101160, 101160, 101150, 
    101160, 101150, 101110, 101070, 101170, 101120, 101080, 100980, 100970, 
    101030, 100940, 100930, 100910, 100870, 100840, 100820, _, _, 100750, _, 
    _, _, _, _, _, _, _, _, 100650, 100590, 100570, 100560, 100560, 100570, 
    100570, 100540, 100520, 100520, 100520, _, _, _, 100540, _, _, 100560, 
    100550, 100540, 100530, 100540, 100560, 100550, 100570, 100590, 100620, 
    100660, 100680, 100700, 100710, 100720, 100740, 100730, 100740, 100760, 
    _, _, _, _, _, 100900, 100930, 100960, 100990, 101010, 101020, 101050, 
    101070, 101070, 101090, 101110, 101130, 101140, 101160, 101180, 101200, 
    101210, 101230, 101270, 101290, 101310, 101360, 101390, 101430, 101460, 
    101490, 101510, 101550, 101580, 101590, 101590, 101590, 101620, 101640, 
    101660, 101670, 101690, 101700, 101720, 101730, 101730, 101710, 101710, 
    101710, 101710, 101720, 101730, 101750, 101780, 101760, 101760, 101780, 
    101770, 101760, 101750, 101740, 101730, 101720, 101730, 101740, 101740, 
    101730, 101730, 101720, 101700, 101680, 101650, 101620, 101610, 101600, 
    101610, 101610, 101610, 101610, 101700, _, 101590, 101570, 101550, 
    101530, 101510, 101490, 101470, 101460, 101440, 101420, 101390, 101360, 
    101340, 101300, 101260, 101210, 101180, 101150, 101100, 101050, 101000, 
    100960, 100920, 100890, 100870, 100790, 100760, 100750, 100680, 100660, 
    100640, 100610, 100560, 100550, 100540, 100500, 100480, 100460, 100430, 
    100400, 100430, 100440, 100420, _, 100380, 100350, 100360, 100340, _, 
    100360, 100360, 100390, 100430, 100500, 100540, 100560, 100580, _, 
    100620, 100650, 100650, 100670, 100690, 100730, 100770, 100810, _, 
    100930, 101010, 101050, 101110, 101190, 101230, 101260, 101300, 101320, 
    _, 101320, 101320, 101310, 101310, 101280, 101250, 101180, 101110, 
    101050, 100960, 100870, 100790, 100690, 100630, 100620, 100510, 100560, 
    100600, 100640, 100680, 100720, 100730, 100770, 100770, 100810, 100840, 
    100900, 100920, 100930, 100930, 100950, 100950, 100950, 100940, 100950, 
    100930, 100910, 100880, _, 100880, 100890, 100890, 100880, 100900, 
    100890, 100890, 100920, 100910, 100920, 100960, 100980, 100990, 101010, 
    101040, 101060, 101070, 101090, 101080, 101100, 101090, 101110, 101120, 
    101130, 101130, 101170, 101170, 101180, 101180, 101160, 101140, 101130, 
    101120, 101100, 101100, _, 101090, 101110, 101100, 101090, 101070, 
    101020, 100980, 100970, 100980, 100940, _, _, 100910, 100890, 100870, 
    100860, 100860, 100850, 100850, 100820, 100820, 100810, _, 100780, 
    100770, 100770, 100780, 100780, 100770, 100760, 100750, 100740, 100730, 
    _, _, _, _, _, 100750, _, _, 100630, 100620, 100620, 100610, 100610, 
    100620, 100640, 100660, 100700, _, _, _, _, _, _, _, _, _, 100820, 
    100860, 100880, 100900, 100920, 100930, 100950, 100960, 100980, 100990, 
    100990, 101010, 101020, 101050, 101070, 101070, 101070, 101050, 101030, 
    _, _, _, 101000, 100950, 100920, 100890, 100860, 100850, 100820, 100760, 
    100700, 100630, 100570, 100520, 100450, _, 100390, 100350, 100320, 
    100260, 100180, 100110, 100040, 99980, 99900, 99840, 99810, _, 99770, 
    99760, 99760, 99790, 99800, 99820, 99850, 99930, 99990, 100070, 100210, 
    _, _, _, 100570, 100650, 100700, 100800, 100870, 100920, 100970, 101010, 
    101070, 101130, 101180, _, 101250, 101270, 101290, 101290, 101270, 
    101270, 101280, 101260, 101260, 101250, 101230, 101200, 101200, 101160, 
    101130, 101080, 101010, 100970, 100930, 100870, 100800, 100720, 100660, 
    100560, 100480, 100390, 100270, 100150, 100030, 99920, 99840, 99790, 
    99750, 99720, 99700, 99680, 99670, 99660, 99650, 99650, 99650, 99640, 
    99660, 99690, 99710, 99730, 99750, _, _, 99830, _, _, 99850, 99870, 
    99890, 99900, 99900, 99880, 99890, 99900, 99900, 99890, 99880, 99870, 
    99860, 99840, 99840, 99840, 99840, 99840, 99840, _, _, 99920, _, _, _, 
    99730, 99700, 99670, 99640, 99610, 99600, 99550, 99550, 99550, 99560, 
    99580, 99610, 99650, 99710, 99750, 99790, 99830, 99890, 99950, 100020, 
    100240, 100220, 100310, 100390, 100470, 100550, 100590, 100660, 100690, 
    100740, 100770, 100810, 100840, 100870, 100880, 100890, 100890, 100830, 
    100740, 100690, _, 100610, 100540, 100470, 100390, 100280, 100140, 
    100030, 99930, 99790, 99660, _, 99400, 99270, 99080, 98920, 98720, 98530, 
    98330, 98180, 98130, 98120, 98110, 98100, 98090, 98110, 98130, 98210, 
    98270, 98350, 98420, 98550, 98670, 98820, 98970, 99060, 99240, 99470, 
    99650, 99830, 99960, 100080, 100170, 100240, 100320, 100380, 100460, 
    100550, 100600, 100690, 100760, 100820, 100890, 100990, 101060, 101060, 
    101140, 101180, 101230, 101330, 101380, 101490, 101520, 101540, 101600, 
    101620, 101640, 101640, 101650, 101630, 101620, 101610, _, _, 101530, 
    101490, 101460, 101400, 101310, 101230, 101180, 101100, 101030, 101000, 
    100960, 100910, 100860, 100790, 100730, 100650, 100560, 100510, 100440, 
    100390, 100380, 100360, 100340, 100320, 100260, 100170, 100090, 100010, 
    99940, 99850, 99850, 99800, 99790, 99770, 99770, 99770, 99720, 99760, 
    99820, 99770, 99740, 99750, 99790, 99830, 99870, 99910, 99950, 99920, 
    100000, 100050, 100040, 100020, 100010, 100000, 99980, 99980, 99980, 
    100000, 100040, 100070, 100100, 100110, 100080, 100080, 100020, 100000, 
    _, _, _, 100390, _, _, 99940, 99910, 99880, 99850, 99820, 99800, 99780, 
    99760, 99730, 99720, 99750, 99770, 99800, 99840, 99850, 99850, 99880, 
    99890, 99930, 99940, 99970, 100030, _, _, 100080, 100100, 100130, 100160, 
    100190, 100220, 100250, _, 100320, 100350, 100370, 100380, 100440, 
    100460, 100480, 100570, 100630, 100670, 100700, 100720, 100730, 100720, 
    100730, 100770, 100790, 100830, 100870, 100930, 100950, 100960, 101050, 
    101040, 101060, 101100, 101150, 101190, _, _, _, _, _, 101430, 101460, 
    101510, 101560, 101590, 101640, 101690, 101750, 101810, 101860, 102030, 
    102050, 102050, 102010, 102040, 102060, 102030, 102070, 102100, 102100, 
    102120, 102110, _, _, 102090, 102070, 102060, 102060, 102010, 101990, 
    101970, 101950, 101950, 101930, 101890, 101850, 101850, 101810, 101800, 
    101800, 101820, 101840, 101850, 101870, 101880, 101900, 101910, 101880, 
    101870, 101860, 101850, 101830, 101810, 101810, 101810, 101800, 101780, 
    101760, 101730, 101700, 101670, _, 101620, 101590, 101560, 101560, 
    101550, 101550, 101540, 101510, 101470, 101390, 101340, 101260, 101240, 
    101220, 101150, 101120, 101080, _, _, 101010, 100920, 100870, 100810, 
    100780, 100750, 100700, 100650, 100610, 100590, 100580, 100540, 100490, 
    100420, 100390, 100340, 100270, 100190, 100110, 100040, 99950, 99880, 
    99790, 99710, 99620, 99520, _, 99310, 99210, 99140, 99040, 98940, 98880, 
    98800, 98730, 98700, 98670, 98630, 98590, 98580, 98530, 98480, 98460, 
    98440, 98430, 98410, 98390, 98380, 98360, 98350, 98350, 98380, 98420, 
    98460, 98500, 98520, 98570, 98580, 98590, 98660, 98750, 98800, 98830, 
    98870, _, 98950, 99000, 99050, 99100, 99140, 99180, 99210, 99240, 99280, 
    99320, 99330, 99360, 99380, 99390, 99410, 99420, 99450, 99480, _, 99550, 
    99580, 99570, 99590, 99600, 99640, 99650, 99660, 99660, 99690, _, 99750, 
    99780, 99790, 99790, 99820, 99840, 99860, 99890, 99930, 99980, 100020, 
    100070, 100110, 100160, 100210, 100270, 100320, 100380, 100420, 100460, 
    100510, 100570, 100620, 100670, 100740, 100810, 100850, 100920, 100990, 
    101050, _, 101170, 101200, 101220, 101200, 101210, 101200, 101160, 
    101140, 101140, 101170, _, 101280, 101330, 101350, 101380, 101410, 
    101440, 101480, 101480, 101490, 101500, _, _, _, _, 101570, 101500, 
    101490, 101450, 101410, 101370, 101320, 101280, 101180, 101130, 101060, 
    100970, 100890, 100800, 100720, 100630, 100540, 100440, 100340, 100230, 
    100120, 100020, 99960, 99920, 99910, 99940, 99970, 99960, 100000, 100050, 
    100100, 100130, 100160, 100190, _, 100260, 100300, 100350, _, 100490, 
    100570, 100660, 100740, 100820, _, 100970, 101050, 101130, 101210, 
    101280, 101340, 101440, 101500, 101550, 101590, 101640, 101660, 101630, 
    101610, 101620, 101610, 101600, 101610, 101620, 101620, 101560, 101490, 
    101460, 101420, 101350, 101270, 101220, 101140, 101160, 101200, 101160, 
    101170, 101160, 101140, 101150, 101120, 101160, 101140, 101150, 101160, 
    101180, 101200, 101230, 101250, 101260, 101330, 101410, 101470, 101520, 
    _, _, 101640, _, _, _, _, _, 101560, 101510, 101380, 101210, 101120, 
    101060, 101040, 101110, 101230, 101320, 101440, 101560, 101680, 101780, 
    101860, 101960, 102050, 102140, 102190, _, _, 102450, 102530, 102600, 
    102660, 102690, 102720, 102760, 102820, 102890, 102930, 102990, 103050, 
    103110, 103140, 103170, 103210, 103250, 103260, 103240, 103240, 103280, 
    103320, 103350, 103380, 103400, 103420, 103450, 103490, 103520, 103530, 
    103520, 103560, 103570, 103550, 103630, 103610, _, _, 103570, 103570, 
    103570, 103550, 103550, 103530, 103510, 103510, 103510, 103500, 103510, 
    103490, 103460, 103450, 103440, 103410, 103390, 103380, 103350, 103320, 
    103280, 103260, 103240, 103200, 103170, 103140, 103090, 103030, 102980, 
    102940, _, 102860, 102830, 102800, 102760, 102720, 102690, 102640, 
    102580, 102530, 102470, 102420, 102380, 102350, 102350, 102320, 102240, 
    102200, 102160, 102120, 102060, 102000, 101950, 101900, 101870, 101870, 
    101860, 101830, 101820, 101830, 101830, 101810, 101780, 101790, 101790, 
    101770, 101800, 101820, 101840, 101840, 101880, 101910, 101910, 101890, 
    101880, 101880, 101860, 101850, 101860, 101860, 101840, 101840, 101840, 
    101840, 101820, 101820, 101800, 101790, 101770, 101770, 101760, 101760, 
    101740, 101720, 101710, 101680, 101630, 101600, 101600, 101540, 101500, 
    101470, 101430, 101410, 101360, 101330, 101290, 101280, 101290, 101270, 
    101280, 101270, 101300, 101320, 101340, 101360, 101400, 101430, 101450, 
    101450, 101470, 101500, 101500, 101500, 101490, 101490, 101480, 101470, 
    101480, 101510, 101520, 101540, 101560, 101590, 101600, 101630, 101640, 
    101670, 101700, 101720, 101740, 101760, 101780, 101790, 101810, 101800, 
    101800, 101790, _, 101790, 101790, 101790, 101790, 101810, 101830, 
    101840, 101850, 101850, 101850, 101850, 101850, 101860, 101880, 101900, 
    101920, 101940, 102010, 102060, 102130, 102180, 102200, 102220, 102250, 
    102270, 102270, 102270, 102280, 102300, 102290, 102300, 102300, 102280, 
    102250, 102230, 102200, 102160, 102120, 102110, 102100, 102060, 102020, 
    _, 102060, 101920, 101880, 101850, 101820, 101770, 101740, 101720, 
    101690, 101670, 101660, 101630, 101600, 101580, 101560, 101500, 101480, 
    101450, 101420, 101410, 101370, _, 101300, 101260, 101230, 101170, 
    101140, 101090, 101070, 101060, 101040, 101030, 101040, 101060, 101100, 
    101120, 101150, 101190, 101240, 101260, 101280, 101300, _, 101350, 
    101380, 101410, 101440, 101460, 101470, 101490, 101520, 101540, 101560, 
    101570, _, 101620, 101640, 101670, 101690, 101730, 101750, 101770, 
    101790, 101800, 101800, _, _, 101980, _, _, _, _, 101690, 101670, 101650, 
    101630, 101580, 101530, 101500, 101480, 101450, 101460, 101440, 101440, 
    101430, 101420, 101400, 101400, 101400, 101400, _, 101560, _, _, 101390, 
    101400, 101400, 101390, 101380, 101350, 101330, 101320, 101310, 101310, 
    101300, 101300, 101340, 101370, 101380, 101390, 101390, 101400, 101420, 
    101420, 101430, 101440, 101450, 101470, 101480, 101500, 101520, 101520, 
    101500, 101480, 101510, 101510, 101500, 101480, 101510, 101540, 101560, 
    101590, 101610, 101640, 101650, 101630, _, 101590, 101570, 101530, _, _, 
    101460, 101430, 101430, 101390, 101360, 101320, 101260, 101240, 101200, 
    101160, 101130, _, _, 101070, 101050, 101020, 100980, 100920, 100880, 
    100840, 100790, 100750, 100720, _, _, _, 100740, _, _, _, 100510, 100490, 
    100470, 100440, 100390, 100450, 100460, 100490, 100540, 100580, 100580, 
    100570, 100570, 100570, 100570, 100590, 100580, 100560, 100530, 100530, 
    100480, _, _, 100340, 100290, 100240, 100220, 100190, 100170, 100180, 
    100220, 100220, 100210, 100190, 100170, 100170, _, 100180, 100190, 
    100210, 100210, 100220, 100240, 100230, 100200, 100180, 100170, 100100, 
    100110, 100040, 100010, 100060, 100070, 100070, 100080, 100090, 100100, 
    100140, 100150, 100190, 100230, 100270, 100280, 100350, 100370, 100390, 
    100400, 100410, 100410, 100410, 100350, 100290, 100230, 100180, 100100, 
    100030, 99980, 99930, 99880, 99880, 99810, 99780, 99750, 99710, 99690, 
    99650, 99620, _, 99570, 99530, 99490, 99450, 99400, 99370, 99360, 99330, 
    99290, 99270, _, 99250, 99240, 99230, 99220, 99220, 99220, 99250, 99280, 
    99290, 99300, _, _, 99530, 99410, 99450, 99510, 99550, 99600, 99650, 
    99700, 99770, 99820, 99860, 99890, 99960, 100040, 100120, 100190, 100240, 
    100300, 100330, 100380, 100400, 100420, 100470, 100480, 100540, 100590, 
    100620, 100680, 100700, 100790, _, _, 100730, 100730, 100720, 100710, 
    100700, 100730, 100760, 100770, 100800, 100800, 100830, 100840, 100840, 
    100880, 100880, 100870, 100890, 100910, 100930, 100940, 100960, 101000, 
    101030, 101050, 101070, 101080, 101100, 101140, 101190, 101230, 101280, 
    101340, 101400, 101420, 101460, 101480, 101510, 101530, 101540, 101550, 
    101580, 101590, 101610, 101640, 101660, 101660, 101660, 101680, 101680, 
    101680, 101680, 101680, 101700, 101700, 101730, 101740, 101730, 101720, 
    101720, 101690, 101660, 101620, 101590, 101560, 101540, 101510, 101500, 
    101480, 101430, 101390, 101360, 101320, 101290, 101260, 101230, 101210, 
    101190, 101190, 101180, 101150, 101110, 101120, 101080, 101050, 101030, 
    100980, 100930, 100900, 100860, 100840, 100810, 100780, 100740, 100710, 
    100650, 100610, 100570, 100530, 100490, 100460, 100430, 100380, 100380, 
    100360, 100350, 100320, 100290, 100250, 100230, 100230, 100230, 100210, 
    100200, 100210, 100200, 100190, 100160, 100150, 100140, 100120, 100120, 
    100110, 100100, 100100, 100130, 100130, 100150, 100140, 100160, 100150, 
    100170, 100190, 100200, 100210, 100230, 100250, 100310, 100360, 100400, 
    100430, 100460, 100480, 100480, 100480, 100500, 100520, 100550, 100550, 
    100520, 100540, 100530, 100530, 100510, 100490, 100470, 100470, 100440, 
    100400, 100400, 100370, 100340, 100280, 100250, 100200, 100150, 100110, 
    100060, 100010, 99970, 99900, 99870, 99860, 99830, 99840, 99850, 99870, 
    99880, 99860, 99890, 99900, 99910, 99970, 100040, 100080, 100150, 100230, 
    100280, 100330, 100400, 100490, 100530, 100570, 100610, 100620, 100670, 
    100690, 100730, 100760, 100780, 100830, 100830, 100870, 100860, 100860, 
    100880, 100880, 100860, 100850, 100840, 100810, 100780, 100720, 100640, 
    100550, 100520, 100490, 100430, 100360, 100320, 100290, 100220, 100160, 
    100110, 100060, 99990, 99930, 99860, 99770, 99640, 99520, 99420, 99330, 
    99220, 99150, 99070, 98960, 98850, 98730, 98640, 98570, 98480, 98420, 
    98330, 98270, 98290, 98300, 98290, 98410, 98500, 98570, 98610, 98690, 
    98760, 98820, 98880, 98890, 98920, 99020, 99090, 99170, 99250, 99320, 
    99390, 99450, 99560, 99650, 99720, 99790, 99900, 99970, 100000, 100060, 
    100110, 100170, 100160, 100160, 100200, 100220, 100240, 100250, 100240, 
    100250, 100280, 100300, 100320, 100350, 100360, 100380, 100390, 100410, 
    100420, 100460, 100490, 100530, 100580, 100630, 100690, 100760, 100810, 
    100860, 100910, 100950, 100990, 101020, 101040, 101020, 101020, 101040, 
    101050, 101070, 101060, 101070, 101070, 101090, 101120, 101160, 101200, 
    101230, 101300, 101360, 101410, 101470, 101490, 101510, 101530, 101570, 
    101600, 101630, 101670, 101710, 101740, 101760, 101810, 101870, 101900, 
    101910, 101940, 101980, 102020, 102060, 102110, 102180, 102230, 102290, 
    102340, 102380, 102410, 102430, 102470, 102500, 102530, 102560, 102550, 
    102570, 102570, 102610, 102620, 102640, 102640, 102610, 102650, 102630, 
    102660, 102680, 102690, 102720, 102750, 102800, 102850, 102870, 102890, 
    102880, 102910, 102920, 102920, 102940, 102980, 103000, 103040, 103060, 
    103100, 103120, 103130, 103140, 103140, 103130, 103140, 103130, 103130, 
    103140, 103110, 103070, 103060, 103050, 102990, 102930, 102880, 102840, 
    102760, 102700, 102620, 102520, 102410, 102310, 102200, 102060, 101920, 
    101760, 101570, 101400, 101200, 101050, 100970, 100820, 100640, 100560, 
    100450, 100450, 100430, 100440, 100400, 100400, 100450, 100570, 100620, 
    100660, 100750, 100800, 100840, 100900, 101000, 101060, 101090, 101130, 
    101210, 101250, 101290, 101370, 101410, 101410, 101400, 101410, 101420, 
    101400, 101340, 101340, 101340, 101320, 101280, 101260, 101240, 101180, 
    101120, 101000, 100880, 100830, 100730, 100620, 100480, 100360, 100210, 
    100110, 99990, 99930, 99880, 99820, 99820, 99830, 99850, 99840, 99860, 
    99870, 99900, 99950, 99940, 99980, 99980, 99980, 99970, 99990, 99980, 
    99980, 99980, 100020, 100060, 100040, 100070, 100110, 100140, 100170, 
    100200, 100200, 100260, 100280, 100320, 100380, 100410, 100450, 100490, 
    100490, 100520, 100520, 100510, 100530, 100510, 100480, 100490, 100510, 
    100540, 100570, 100600, 100700, 100770, 100890, 101000, 101100, 101200, 
    101350, 101440, 101540, 101630, 101730, 101760, 101860, 101910, 101980, 
    101970, 102000, 102020, 101980, 102000, 101950, 101930, 101860, 101880, 
    101850, 101760, 101710, 101640, 101560, 101470, 101430, 101420, 101400, 
    101360, 101300, 101290, 101230, 101200, 101130, 101040, 100980, 100910, 
    100860, 100770, 100740, 100660, 100640, 100680, 100670, 100760, 100830, 
    100840, 100860, 100910, 100930, 100980, 101000, 101040, 101060, 101120, 
    101150, 101170, 101180, 101180, 101140, 101150, 101120, 101090, 101030, 
    101010, 101000, 100980, 101010, 100960, 100920, 100910, 100990, 100960, 
    100980, 101010, 101030, 101070, 101050, 101040, 101030, 101000, 100990, 
    100950, 100900, 100910, 100920, 100880, 100860, 100860, 100850, 100800, 
    100790, 100720, 100710, 100610, 100490, 100390, 100290, 100200, 100080, 
    99950, 99830, 99780, 99680, 99790, 99900, 99980, 100090, 100200, 100360, 
    100510, 100470, 100540, 100630, 100720, 100730, 100760, 100790, 100800, 
    100820, 100790, 100750, 100720, 100670, 100660, 100690, 100670, 100660, 
    100660, 100620, 100620, 100620, 100630, 100640, 100640, 100650, 100660, 
    100690, 100740, 100770, 100760, 100740, 100780, 100780, 100790, 100790, 
    100770, 100790, 100800, 100780, 100780, 100790, 100800, 100790, 100790, 
    100750, 100720, 100650, 100610, 100610, 100620, 100550, 100530, 100480, 
    100410, 100400, 100340, 100250, 100150, 100090, 100060, 100040, 100000, 
    99980, 99940, 99950, 99930, 99880, 99790, 99710, 99640, 99560, 99500, 
    99450, 99430, 99420, 99350, 99250, 99190, 99150, 99090, 99050, 99050, 
    99100, 99150, 99190, 99260, 99350, 99420, 99510, 99570, 99620, 99630, 
    99650, 99660, 99670, 99610, 99610, 99550, 99540, 99490, 99450, 99460, 
    99560, 99680, 99810, 99980, 100110, 100290, 100470, 100690, 100930, 
    101180, 101380, 101560, 101730, 101870, 101980, 102090, 102170, 102260, 
    102320, 102400, 102470, 102560, 102590, 102670, 102690, 102730, 102740, 
    102740, 102780, 102810, 102840, 102870, 102890, 102890, 102910, 102940, 
    102950, 102970, 102960, 102950, 102970, 102970, 102990, 102990, 103000, 
    103000, 103000, 102980, 102970, 102970, 102950, 102940, 102920, 102860, 
    102840, 102780, 102740, 102690, 102650, 102610, 102570, 102550, 102510, 
    102470, 102410, 102380, 102350, 102340, 102330, 102300, 102280, 102270, 
    102230, 102190, 102160, 102090, 102070, 102070, 102020, 102020, 102090, 
    102060, 101990, 101990, 101960, 101900, 101880, 101830, 101760, 101690, 
    101670, 101680, 101680, 101630, 101640, 101590, 101530, 101460, 101430, 
    101390, 101340, 101280, 101240, 101220, 101200, 101170, 101150, 101170, 
    101100, 101020, 101010, 100980, 100930, 100930, 100910, 100890, 100860, 
    100860, 100910, 100900, 100890, 100910, 100920, 100950, 100970, 101020, 
    100950, 100970, 101030, 101110, 101170, 101230, 101260, 101310, 101410, 
    101470, 101510, 101590, 101580, 101580, 101630, 101640, 101650, 101650, 
    101650, 101640, 101630, 101630, 101590, 101560, 101520, 101490, 101460, 
    101420, 101400, 101370, 101320, 101270, 101190, 101130, 101040, 100940, 
    100860, 100790, 100650, 100570, 100510, 100390, 100250, 100130, 100010, 
    99890, 99760, 99670, 99510, 99390, 99290, 99190, 99110, 99000, 98920, 
    98840, 98760, 98640, 98540, 98450, 98360, 98340, 98220, 98120, 98090, 
    98040, 97980, 97890, 97840, 97760, 97710, 97660, 97600, 97500, 97450, 
    97410, 97340, 97290, 97260, 97210, 97180, 97120, 97040, 97030, 97030, 
    97010, 97070, 97090, 97100, 97130, 97200, 97240, 97300, 97390, 97400, 
    97510, 97550, 97660, 97750, 97850, 97920, 98020, 98090, 98170, 98200, 
    98200, 98240, 98300, 98390, 98390, 98420, 98450, 98500, 98560, 98610, 
    98620, 98600, 98650, 98650, 98680, 98690, 98670, 98700, 98740, 98750, 
    98770, 98780, 98760, 98760, 98770, 98750, 98740, 98720, 98710, 98720, 
    98720, 98730, 98750, 98760, 98750, 98750, 98750, 98760, 98790, 98800, 
    98800, 98840, 98880, 98890, 98900, 98910, 98930, 98920, 98920, 98890, 
    98890, 98900, 98910, 98940, 98990, 99040, 99090, 99130, 99130, 99150, 
    99150, 99150, 99180, 99210, 99200, 99210, 99240, 99240, 99220, 99190, 
    99190, 99150, 99080, 99040, 98990, 98940, 98880, 98860, 98790, 98720, 
    98640, 98520, 98440, 98350, 98280, 98150, 98020, 97870, 97740, 97720, 
    97680, 97660, 97560, 97520, 97470, 97400, 97400, 97370, 97360, 97350, 
    97350, 97350, 97360, 97370, 97380, 97390, 97380, 97360, 97400, 97400, 
    97380, 97390, 97390, 97400, 97380, 97370, 97380, 97360, 97330, 97320, 
    97330, 97350, 97350, 97340, 97330, 97370, 97420, 97450, 97510, 97580, 
    97660, 97740, 97810, 97870, 97920, 97970, 98040, 98100, 98150, 98200, 
    98220, 98240, 98260, 98280, 98280, 98310, 98340, 98390, 98400, 98450, 
    98530, 98580, 98610, 98620, 98650, 98690, 98690, 98690, 98700, 98690, 
    98680, 98680, 98690, 98690, 98650, 98650, 98640, 98640, 98600, 98580, 
    98570, 98560, 98570, 98540, 98530, 98510, 98500, 98480, 98460, 98450, 
    98410, 98390, 98370, 98330, 98310, 98270, 98260, 98220, 98210, 98210, 
    98210, 98190, 98200, 98190, 98180, 98180, 98180, 98190, 98190, 98170, 
    98150, 98150, 98140, 98160, 98170, 98170, 98210, 98230, 98260, 98300, 
    98340, 98380, 98450, 98520, 98570, 98600, 98610, 98640, 98670, 98720, 
    98740, 98800, 98900, 98990, 99040, 99100, 99130, 99190, 99220, 99260, 
    99310, 99390, 99400, 99460, 99510, 99540, 99590, 99620, 99610, 99660, 
    99670, 99690, 99710, 99730, 99730, 99760, 99760, 99780, 99750, 99740, 
    99730, 99680, 99660, 99650, 99590, 99550, 99520, 99510, 99450, 99430, 
    99390, 99330, 99250, 99220, 99160, 99120, 99070, 99040, 99020, 99050, 
    99090, 99190, 99230, 99270, 99280, 99290, 99310, 99320, 99350, 99360, 
    99340, 99310, 99330, 99340, 99350, 99380, 99420, 99430, 99460, 99470, 
    99490, 99520, 99560, 99600, 99670, 99730, 99810, 99820, 99840, 99880, 
    99930, 99970, 100000, 100040, 100080, 100100, 100160, 100200, 100220, 
    100260, 100290, 100330, 100350, 100360, 100390, 100380, 100400, 100430, 
    100460, 100460, 100500, 100480, 100490, 100490, 100490, 100520, 100520, 
    100530, 100510, 100490, 100490, 100500, 100490, 100480, 100480, 100490, 
    100460, 100450, 100440, 100420, 100410, 100430, 100460, 100470, 100450, 
    100420, 100410, 100390, 100400, 100400, 100420, 100420, 100420, 100420, 
    100440, 100410, 100400, 100390, 100430, 100420, 100450, 100440, 100430, 
    100450, 100450, 100450, 100490, 100510, 100530, 100500, 100500, 100510, 
    100520, 100510, 100530, 100520, 100540, 100560, 100570, 100580, 100600, 
    100590, 100610, 100600, 100610, 100610, 100600, 100590, 100590, 100630, 
    100640, 100680, 100690, 100710, 100730, 100740, 100750, 100770, 100780, 
    100790, 100800, 100810, 100810, 100870, 100910, 100920, 100960, 100990, 
    101020, 101050, 101060, 101070, 101070, 101130, 101160, 101220, 101260, 
    101280, 101340, 101370, 101400, 101440, 101460, 101490, 101490, 101520, 
    101530, 101570, 101610, 101610, 101600, 101630, 101660, 101650, 101670, 
    101720, 101720, 101720, 101760, 101800, 101800, 101840, 101870, 101890, 
    101910, 101940, 101950, 101960, 101980, 102000, 102030, 102050, 102080, 
    102080, 102110, 102140, 102120, 102150, 102160, 102160, 102140, 102130, 
    102150, 102150, 102140, 102130, 102090, 102050, 102020, 102000, 102000, 
    101960, 101930, 101890, 101860, 101850, 101820, 101770, 101710, 101670, 
    101640, 101580, 101490, 101400, 101350, 101270, 101190, 101140, 101100, 
    101070, 101010, 100930, 100880, 100820, 100780, 100690, 100650, 100560, 
    100490, 100440, 100360, 100260, 100180, 100120, 100040, 99960, 99870, 
    99870, 99770, 99750, 99810, 99850, 99890, 99910, 99940, 99890, 99900, 
    99950, 99980, 99940, 99930, 99910, 99910, 99910, 99910, 99880, 99840, 
    99790, 99670, 99580, 99470, 99380, 99180, 99030, 98870, 98760, 98670, 
    98580, 98400, 98280, 98090, 97980, 97830, 97750, 97650, 97620, 97550, 
    97510, 97490, 97490, 97540, 97600, 97650, 97720, 97740, 97750, 97780, 
    97850, 97960, 98040, 98130, 98160, 98230, 98250, 98310, 98360, 98400, 
    98430, 98450, 98470, 98510, 98520, 98530, 98540, 98540, 98530, 98530, 
    98520, 98490, 98450, 98450, 98450, 98450, 98440, 98430, 98390, 98360, 
    98320, 98300, 98260, 98230, 98180, 98150, 98130, 98090, 98060, 98040, 
    98000, 97960, 97950, 97940, 97900, 97880, 97830, 97810, 97800, 97810, 
    97810, 97800, 97790, 97780, 97760, 97760, 97780, 97800, 97790, 97820, 
    97850, 97890, 97970, 98050, 98110, 98180, 98250, 98330, 98400, 98510, 
    98620, 98720, 98870, 98990, 99120, 99210, 99300, 99410, 99510, 99630, 
    99720, 99800, 99890, 99940, 100010, 100110, 100190, 100280, 100350, 
    100410, 100490, 100570, 100650, 100700, 100770, 100840, 100910, 100980, 
    101060, 101100, 101150, 101210, 101260, 101310, 101350, 101380, 101430, 
    101470, 101520, 101560, 101600, 101650, 101700, 101720, 101750, 101790, 
    101790, 101810, 101820, 101830, 101870, 101900, 101890, 101900, 101890, 
    101910, 101910, 101900, 101880, 101900, 101860, 101810, 101820, 101780, 
    101740, 101700, 101680, 101600, 101540, 101480, 101370, 101290, 101150, 
    101030, 100960, 100880, 100780, 100680, 100600, 100510, 100400, 100280, 
    100180, 100120, 100030, 99950, 99920, 99870, 99800, 99740, 99690, 99630, 
    99590, 99540, 99510, 99450, 99410, 99380, 99360, 99310, 99310, 99300, 
    99240, 99210, 99140, 99050, 98970, 98950, 98920, 98920, 98940, 98980, 
    99030, 99120, 99200, 99220, 99280, 99300, 99360, 99400, 99430, 99470, 
    99490, 99470, 99500, 99530, 99520, 99510, 99540, 99560, 99540, 99550, 
    99560, 99550, 99540, 99480, 99410, 99410, 99410, 99380, 99340, 99320, 
    99320, 99280, 99390, 99460, 99510, 99550, 99630, 99660, 99690, 99780, 
    99840, 99860, 99880, 99920, 99970, 100050, 100080, 100160, 100210, 
    100260, 100320, 100340, 100380, 100420, 100440, 100460, 100480, 100500, 
    100510, 100520, 100490, 100500, 100480, 100460, 100450, 100420, 100410, 
    100410, 100410, 100390, 100390, 100410, 100420, 100450, 100430, 100430, 
    100460, 100460, 100470, 100480, 100490, 100550, 100580, 100600, 100630, 
    100640, 100690, 100700, 100720, 100750, 100760, 100790, 100820, 100840, 
    100860, 100860, 100870, 100890, 100920, 100920, 100940, 100940, 100920, 
    100890, 100890, 100880, 100890, 100890, 100900, 100890, 100860, 100830, 
    100790, 100760, 100740, 100720, 100690, 100670, 100640, 100600, 100560, 
    100510, 100460, 100400, 100360, 100290, 100240, 100200, 100160, 100130, 
    100130, 100160, 100200, 100220, 100250, 100330, 100360, 100410, 100390, 
    100400, 100360, 100360, 100350, 100370, 100370, 100390, 100410, 100390, 
    100390, 100380, 100370, 100370, 100320, 100300, 100330, 100400, 100370, 
    100380, 100410, 100410, 100430, 100450, 100460, 100450, 100440, 100440, 
    100450, 100460, 100460, 100470, 100470, 100480, 100490, 100480, 100480, 
    100460, 100440, 100450, 100430, 100440, 100430, 100410, 100410, 100420, 
    100400, 100410, 100430, 100440, 100460, 100520, 100570, 100620, 100670, 
    100710, 100740, 100790, 100800, 100820, 100830, 100840, 100840, 100860, 
    100900, 100930, 100950, 100970, 100980, 100970, 100950, 100970, 100960, 
    100950, 100960, 100990, 100950, 100970, 100990, 101010, 101030, 101040, 
    101060, 101090, 101100, 101100, 101120, 101140, 101180, 101220, 101270, 
    101300, 101330, 101360, 101370, 101390, 101410, 101430, 101460, 101470, 
    101510, 101560, 101600, 101650, 101660, 101660, 101660, 101680, 101670, 
    101650, 101630, 101620, 101590, 101530, 101480, 101380, 101320, 101200, 
    101080, 101010, 100960, 100910, 100900, 100910, 100970, 101050, 101180, 
    101190, 101300, 101330, 101350, 101300, 101260, 101190, 101090, 100960, 
    100850, 100730, 100590, 100470, 100330, 100220, 100110, 100000, 99910, 
    99920, 99870, 99860, 99890, 99940, 99970, 100020, 100060, 100040, 100060, 
    100090, 100110, 100150, 100100, 100240, 100340, 100400, 100490, 100590, 
    100680, 100780, 100840, 100910, 101030, 101110, 101180, 101250, 101330, 
    101400, 101460, 101530, 101600, 101650, 101700, 101720, 101780, 101810, 
    101860, 101900, 101940, 101950, 101950, 101950, 101940, 101880, 101820, 
    101720, 101610, 101490, 101400, 101260, 101080, 100900, 100720, 100620, 
    100570, 100480, 100440, 100380, 100280, 100220, 100130, 100070, 100110, 
    100120, 100170, 100170, 100180, 100140, 100100, 100080, 100100, 100080, 
    100110, 100110, 100050, 100050, 100070, 100040, 100040, 100040, 100030, 
    100070, 100060, 100070, 100110, 100130, 100140, 100150, 100170, 100210, 
    100250, 100130, 100120, 100130, 100160, 100170, 100160, 100140, 100130, 
    100120, 100090, 100080, 100080, 100040, 100000, 99980, 99960, 99950, 
    99970, 99970, 99960, 99990, 100010, 100060, 100090, 100100, 100090, 
    100120, 100160, 100190, 100210, 100260, 100300, 100320, 100350, 100390, 
    100420, 100440, 100470, 100490, 100500, 100540, 100560, 100590, 100630, 
    100690, 100720, 100740, 100770, 100780, 100810, 100810, 100810, 100770, 
    100790, 100780, 100770, 100760, 100730, 100750, 100690, 100690, 100670, 
    100620, 100610, 100610, 100570, 100560, 100570, 100540, 100570, 100560, 
    100570, 100540, 100580, 100580, 100620, 100670, 100700, 100690, 100730, 
    100750, 100750, 100780, 100830, 100810, 100860, 100850, 100840, 100880, 
    100920, 100920, 100990, 100970, 101030, 101080, 101070, 101080, 101110, 
    101120, 101190, 101190, 101200, 101190, 101160, 101170, 101230, 101250, 
    101250, 101240, 101230, 101270, 101280, 101320, 101310, 101330, 101380, 
    101400, 101440, 101480, 101490, 101490, 101500, 101490, 101510, 101480, 
    101420, 101380, 101370, 101360, 101320, 101340, 101330, 101290, 101250, 
    101220, 101170, 101170, 101160, 101140, 101140, 101180, 101200, 101240, 
    101230, 101250, 101270, 101260, 101280, 101300, 101310, 101320, 101330, 
    101350, 101380, 101410, 101410, 101420, 101470, 101470, 101480, 101510, 
    101520, 101540, 101580, 101640, 101640, 101640, 101680, 101650, 101640, 
    101650, 101680, 101680, 101660, 101650, 101650, 101640, 101690, 101690, 
    101700, 101690, 101690, 101690, 101690, 101690, 101710, 101710, 101730, 
    101750, 101790, 101810, 101820, 101840, 101860, 101870, 101890, 101920, 
    101920, 101940, 101950, 101980, 102000, 102040, 102040, 102020, 102030, 
    102020, 101990, 102000, 101990, 102010, 102030, 102040, 102080, 102090, 
    102110, 102130, 102130, 102140, 102140, 102170, 102220, 102210, 102230, 
    102240, 102230, 102270, 102290, 102280, 102280, 102290, 102290, 102300, 
    102340, 102360, 102410, 102450, 102490, 102510, 102490, 102490, 102510, 
    102520, 102560, 102550, 102540, 102530, 102470, 102490, 102460, 102420, 
    102390, 102350, 102320, 102270, 102190, 102110, 102070, 102020, 101960, 
    101900, 101840, 101790, 101710, 101640, 101580, 101480, 101440, 101380, 
    101340, 101250, 101160, 101120, 101080, 101020, 100970, 100870, 100790, 
    100730, 100680, 100590, 100550, 100500, 100440, 100400, 100310, 100230, 
    100110, 100000, 99870, 99730, 99580, 99420, 99270, 99070, 98880, 98740, 
    98580, 98390, 98240, 98060, 97840, 97610, 97390, 97160, 96970, 96770, 
    96630, 96510, 96460, 96450, 96500, 96550, 96610, 96620, 96650, 96750, 
    96840, 96970, 97130, 97370, 97540, 97720, 97930, 98090, 98240, 98360, 
    98460, 98550, 98610, 98630, 98680, 98730, 98760, 98790, _, _, _, 98880, 
    98870, 98870, 98870, 98840, 98850, 98840, 98820, 98790, 98780, 98670, 
    98630, 98610, 98580, 98560, 98520, 98500, 98500, 98500, 98500, 98490, 
    98470, 98480, 98500, 98520, 98560, 98610, 98600, 98620, 98670, 98730, 
    98780, 98860, 98920, 98960, 98980, 98960, 98960, 98980, 99000, 99040, 
    99080, 99080, 99110, 99110, 99110, 99120, 99130, 99170, 99170, 99160, 
    99140, 99150, 99160, 99190, 99210, 99250, 99260, 99230, 99170, 99140, 
    99100, 99070, _, 99000, 98960, 98860, 98790, 98750, 98670, 98600, 98510, 
    98420, 98320, 98270, 98260, 98220, 98160, 98100, 98090, 98120, 98140, 
    98150, 98140, 98170, 98200, 98220, 98230, 98260, 98300, 98360, 98440, 
    98500, 98540, 98580, 98600, 98600, 98640, 98670, 98680, 98670, 98680, 
    98690, 98700, 98730, 98730, 98730, 98700, 98700, 98680, 98650, 98670, 
    98670, 98650, 98610, 98580, 98580, 98560, 98530, 98520, 98490, 98460, 
    98450, 98420, 98450, 98430, 98440, 98450, 98460, 98450, 98450, 98460, 
    98480, 98500, 98520, 98530, 98530, 98540, 98600, 98640, 98680, 98710, 
    98710, 98750, 98790, 98840, 98880, 98920, 98940, 98980, 99020, 99050, 
    99080, 99120, 99140, 99170, 99200, 99240, 99250, 99290, 99330, 99370, 
    99450, 99520, 99590, 99640, 99720, 99790, 99860, 99940, 100020, 100070, 
    100130, 100220, 100330, 100420, 100490, 100570, 100600, 100650, 100670, 
    100730, 100740, 100760, 100780, 100800, 100870, 100890, 100890, 100940, 
    101000, 101030, 101060, 101130, 101210, 101240, 101330, 101370, 101450, 
    101500, 101560, 101580, 101600, 101650, 101640, 101600, 101600, 101510, 
    101390, 101260, 101130, 100930, 100730, 100550, 100310, 100080, 99820, 
    99540, 99290, 99040, 98750, 98560, 98400, 98320, 98260, 98240, 98240, 
    98210, 98180, 98160, 98150, 98120, 98100, 98060, 98030, 98010, 98000, 
    97980, 98010, 98030, 98040, 98030, 97950, 97910, 97860, 97950, 97970, 
    98050, 98190, 98250, 98320, 98320, 98350, 98340, 98300, 98290, 98250, 
    98230, 98260, 98210, 98200, 98160, 98110, 98030, 97980, 97890, 97910, 
    97890, 97910, 97950, 98000, 98080, 98110, 98120, 98140, 98160, 98180, 
    98210, 98270, 98290, 98360, 98380, 98420, 98490, 98530, 98570, 98650, 
    98680, 98730, 98770, 98800, 98810, 98800, 98830, 98860, 98890, 98920, 
    98940, 98970, 98980, 98960, 98970, 98980, 98990, 99020, 99040, 99040, 
    99060, 99100, 99160, 99190, 99150, 99160, 99190, 99190, 99180, 99160, 
    99180, 99200, 99220, 99200, 99200, 99210, 99210, 99190, 99200, 99240, 
    99240, 99260, 99250, 99280, 99320, 99340, 99340, 99330, 99320, 99310, 
    99280, 99230, 99200, 99180, 99170, 99150, 99140, 99120, 99100, 99090, 
    99060, 99030, 99010, 98990, 98990, 98990, 98970, 98950, 98970, 98970, 
    98950, 98940, 98930, 98910, 98910, 98890, 98880, 98870, 98850, 98860, 
    98860, 98840, 98800, 98770, 98730, 98730, 98700, 98660, 98670, 98660, 
    98640, 98650, 98650, 98640, 98660, 98700, 98700, 98680, 98700, 98740, 
    98760, 98810, 98840, 98880, 98920, 98970, 98980, 99040, 99090, 99130, 
    99160, 99240, 99300, 99340, 99410, 99450, 99520, 99580, 99630, 99680, 
    99690, 99730, 99760, 99780, 99830, 99870, 99900, 99950, 100010, 100050, 
    100090, 100100, 100120, 100150, 100180, 100210, 100200, 100220, 100260, 
    100290, 100300, 100340, 100320, 100310, 100300, 100240, 100270, 100250, 
    100240, 100250, 100190, 100150, 100140, 100130, 100080, 99970, 99870, 
    99740, 99700, 99630, 99560, 99550, 99550, 99530, 99510, 99510, 99460, 
    99400, 99380, 99380, 99370, 99350, 99340, 99370, 99430, 99460, 99490, 
    99530, 99610, 99670, 99740, 99800, 99860, 99910, 99970, 100020, 100110, 
    100180, 100280, 100390, 100470, 100550, 100630, 100690, 100770, 100830, 
    100880, 100970, 101000, 101040, 101130, 101180, 101230, 101240, 101260, 
    101280, 101250, 101240, 101230, 101240, 101230, 101220, 101230, 101270, 
    101200, 101080, 101060, 101100, 101050, 100970, 100950, 100870, 100840, 
    100770, 100710, 100680, 100620, 100560, 100540, 100500, 100410, 100370, 
    100330, 100270, 100250, 100240, 100220, 100230, 100180, 100160, 100150, 
    100110, 100070, 100050, 100030, 99990, 99930, 99940, 99880, 99880, 99830, 
    99760, 99730, 99740, 99700, 99660, 99580, 99550, 99540, 99540, 99540, 
    99510, 99490, 99450, 99480, 99440, 99440, 99410, 99440, 99380, 99340, 
    99370, 99410, 99450, 99460, 99450, 99480, 99480, 99480, 99480, 99460, 
    99460, 99460, 99500, 99520, 99550, 99550, 99530, 99530, 99510, 99470, 
    99460, 99420, 99380, 99350, 99270, 99300, 99200, 99170, 99120, 99070, 
    99020, 98980, 98960, 98970, 98970, 99000, 99040, 99090, 99110, 99180, 
    99210, 99250, 99290, 99310, 99370, 99440, 99510, 99580, 99660, 99710, 
    99740, 99800, 99850, 99990, 100040, 100080, 100110, 100140, 100210, 
    100250, 100260, 100270, 100280, 100280, 100260, 100260, 100270, 100260, 
    100220, 100180, 100210, 100170, 100130, 100100, 100070, 100040, 99950, 
    99910, 99860, 99800, 99770, 99740, 99750, 99730, 99710, 99690, 99700, 
    99750, 99750, 99740, 99780, 99790, 99790, 99810, 99790, 99770, 99770, 
    99750, 99700, 99630, 99530, 99450, 99410, 99330, 99230, 99160, 99050, 
    99000, 98930, 98840, 98800, 98740, 98630, 98570, 98510, 98450, 98400, 
    98370, 98380, 98320, 98280, 98230, 98190, 98160, 98120, 98080, 98040, 
    97980, 97930, 97850, 97820, 97780, 97760, 97710, 97650, 97560, 97390, 
    97250, 97120, 96980, 96770, 96570, 96840, 96650, 96530, 96390, 96220, 
    96070, 95950, 95830, 95710, 95580, 95470, 95370, 95250, 95150, 95090, 
    95070, 95050, 95050, 95080, 95130, 95180, 95180, 95170, 95160, 95400, 
    95390, 95390, 95380, 95400, 95410, 95430, 95460, 95500, 95520, 95560, 
    95590, 95780, 95830, 95890, 95950, 96040, 96100, 96170, 96260, 96350, 
    96430, 96520, 96620, 96750, 96820, 96900, 97000, 97070, 97160, 97250, 
    97320, 97400, 97460, 97510, 97580, 97640, 97720, 97780, 97960, 98050, 
    98110, 98210, 98320, 98420, 98500, 98570, 98520, 98590, 98690, 98790, 
    98900, 98980, 99040, 99120, 99210, 99290, 99350, 99430, 99390, 99470, 
    99540, 99640, 99740, 99830, 99900, 99970, 100040, 100080, 100120, 100110, 
    100150, 100170, 100220, 100250, 100220, 100230, 100210, 100180, 100170, 
    100120, 100080, 100020, 100060, 99950, 99890, 99820, 99700, 99500, 99310, 
    99170, 98990, 98780, 98610, 98490, 98500, 98470, 98520, 98640, 98800, 
    98960, 99140, 99320, 99510, 99730, 99800, 100040, 100100, 100190, 100330, 
    100390, 100390, 100370, 100330, 100230, 100140, 100060, 100010, 99940, 
    99930, 99900, 99870, 99870, 99920, 99990, 100100, 100240, 100450, 100670, 
    100820, 101000, 101320, 101440, 101530, 101700, 101770, 101790, 101810, 
    101870, 101850, 101840, 101730, 101670, 101550, 101400, 101220, 101060, 
    100860, 100690, 100500, 100310, 100070, 99920, 99730, 99630, 99550, 
    99480, 99450, 99410, 99360, 99290, 99200, 98990, 98720, 98440, 98070, 
    97820, 97650, 97950, 98040, 98020, 98060, 98150, 98340, 98550, 98800, 
    99110, 99550, 99870, 100090, 100360, 100580, 100810, 101010, _, 101330, 
    _, 101420, 101510, 101480, 101450, 101310, 101370, 101370, 101330, 
    101320, 101300, 101280, 101270, 101230, 101230, 101250, _, 101220, 
    101290, 101350, 101390, 101450, 101520, 101540, 101570, 101550, 101540, 
    101560, 101560, 101590, 101620, 101660, 101690, 101710, 101760, 101870, 
    101770, 101770, 101770, 101770, 101790, 101790, 101790, 101790, 101820, 
    101810, 101790, 101750, 101740, 101730, 101710, 101670, 101650, 101660, 
    101690, 101730, 101740, 101780, 101800, 101810, 101830, 101830, 101850, 
    102040, 102050, 101910, 101950, 101970, 102030, 102080, 102110, 102100, 
    102130, 102150, 102150, 102170, 102220, 102220, 102190, 102210, 102230, 
    102250, 102240, 102250, 102380, 102270, 102300, 102250, 102290, 102310, 
    102330, 102350, 102430, 102450, 102430, 102410, 102400, 102400, 102360, 
    102340, 102320, 102330, 102310, 102280, 102270, 102250, 102280, 102260, 
    102150, 102140, 102100, 102050, 102030, 102010, 101980, 101970, 101940, 
    101930, 101860, 101810, 101750, 101670, 101640, 101560, 101490, 101410, 
    101350, 101310, 101400, 101140, 101310, 101000, 100970, 100920, 100840, 
    101070, 101030, 100740, 100730, 100980, 100960, 100950, 100730, 100740, 
    100750, 100780, 100790, 100800, 100800, 101040, 100870, 100880, 101080, 
    100950, 100990, 101030, 101210, 101080, 101080, 101260, 101150, 101190, 
    101390, 101260, 101440, 101340, 101370, 101390, 101410, 101440, 101480, 
    101510, 101520, 101490, 101610, 101540, 101580, 101580, 101660, 101580, 
    101590, 101590, 101590, 101590, 101600, 101570, 101550, 101550, 101550, 
    101530, 101530, 101530, 101530, 101510, 101490, 101480, 101460, 101440, 
    101440, 101430, 101420, 101410, 101380, 101310, 101320, 101290, 101290, 
    101280, 101310, 101260, 101220, 101150, 101100, 101070, 101040, 100980, 
    100870, 100790, 100690, 100650, 100580, 100510, 100450, 100400, 100510, 
    100360, 100300, 100210, 100110, 100030, 99970, 99960, 99960, 99920, 
    99890, 99830, 99790, 99810, 99830, 99860, 99880, 99890, 99950, 99980, 
    100010, 100010, 100060, 100020, 100050, 99990, 99910, 99880, 99820, 
    99770, 99700, 99660, 99620, 99580, 99530, 99490, 99320, 99280, 99200, 
    99100, 99030, 98970, 98950, 98910, 98870, 98830, 98810, 98800, 98790, 
    98780, 98770, 98770, 98870, 98760, 98780, 98800, 98810, 98840, 98860, 
    98880, 98900, 98930, 98950, 99020, 99080, 99130, 99190, 99240, 99300, 
    99360, 99410, 99450, 99470, 99490, 99520, 99520, 99520, 99550, 99580, 
    99610, 99710, 99760, 99780, 99770, 99760, 99770, 99760, 99720, 99700, 
    99910, 99880, 99930, 99960, 99950, 99950, 99910, 99870, 99840, 99770, 
    99680, 99680, 99770, 99700, 99670, 99620, 99570, 99550, 99500, 99460, 
    99360, 99330, 99300, 99290, 99240, 99190, 99090, 99080, 99120, 99050, 
    99070, 99130, 99020, 99010, 99240, 99250, 99210, 99170, 99310, 99300, 
    99400, 99370, 99430, 99450, 99570, 99620, 99630, 99710, 99760, 99780, 
    99820, 99870, 99920, 99950, 100010, 100100, 100050, 100070, 100070, 
    100100, 100130, 100160, 100170, 100140, 100160, 100150, 100130, 100090, 
    100080, 100100, 100090, 100040, 100000, 100000, 100010, 100060, 100040, 
    99960, 100000, 100020, 100040, 100080, 100090, 100090, 100150, 100140, 
    100220, 100280, 100360, 100390, 100460, 100530, 100560, 100650, 100730, 
    100800, 100900, 100960, 101050, 101120, 101190, 101220, 101340, 101390, 
    101450, 101490, 101570, 101570, 101630, 101720, 101740, 101800, 101830, 
    101860, 101860, 101870, 101890, 101930, 101970, 102000, 102030, 102030, 
    102060, 102100, 102130, 102170, 102200, 102230, 102280, 102300, 102290, 
    102300, 102310, 102310, 102340, 102360, 102400, 102460, 102480, 102490, 
    102500, 102480, 102510, 102510, 102550, 102560, 102580, 102560, 102630, 
    102540, 102520, 102620, 102450, 102420, 102440, 102450, 102460, 102400, 
    102370, 102340, 102320, 102260, 102200, 102180, 102120, 102110, 102050, 
    101960, 101940, 101920, 101830, 101770, 101640, 101680, 101460, 101380, 
    101270, 101180, 101100, 101020, 101110, 100860, 100810, 100730, 100640, 
    100550, 100480, 100410, 100290, 100220, 100130, 100070, 100040, 99980, 
    99910, 99840, 99770, 99710, 99660, 99760, 99550, 99510, 99580, 99440, 
    99400, 99350, 99310, 99230, 99130, 99070, 98980, 98920, 98840, 98810, 
    98770, 98730, 98700, 98680, 98660, 98630, 98690, 98670, 98680, 98740, 
    98710, 98720, 98770, 98830, 98890, 98930, 98990, 99040, 99100, 99160, 
    99210, 99250, 99300, 99350, 99410, 99440, 99470, 99490, 99500, 99530, 
    99520, 99600, 99630, 99550, 99580, 99580, 99570, 99570, 99670, 99560, 
    99560, 99550, 99560, 99570, 99590, 99600, 99600, 99580, 99560, 99540, 
    99530, 99520, 99510, 99510, 99460, 99410, 99370, 99330, 99280, 99230, 
    99220, 99160, 99090, 99080, 99050, 99040, 99040, 99050, 99040, 99060, 
    99080, 99090, 99120, 99150, 99180, 99220, 99280, 99330, 99360, 99410, 
    99550, 99590, 99640, 99650, 99700, 99730, 99780, 99820, 99870, 99890, 
    99960, 99980, 100010, 100010, 100010, 100030, 100040, 100080, 100100, 
    100100, 100110, 100130, 100110, 100130, 100120, 100120, 100120, 100110, 
    100130, 100120, 100130, 100130, 100100, 100110, 100120, 100090, 100080, 
    100060, 100040, 100040, 100040, 100010, 99980, 99940, 99930, 99900, 
    99870, 99830, 99810, 99790, 99770, 99750, 99700, 99690, 99650, 99600, 
    99590, 99500, 99450, 99390, 99360, 99350, 99340, 99350, 99360, 99540, 
    99580, 99650, 99720, 99800, 99850, 99900, 99950, 99990, 100030, 100060, 
    100100, 100120, 100140, 100180, 100190, 100210, 100230, 100230, 100240, 
    100240, 100230, 100250, 100250, 100230, 100210, 100220, 100210, 100170, 
    100150, 100140, 99870, 99820, 99780, 99740, 99670, 99610, 99520, 99440, 
    99340, 99240, 99270, 99250, 99290, 99340, 99430, 99500, 99590, 99730, 
    99880, 99990, 100130, 100290, 100410, 100520, 100630, 100700, 100730, 
    100780, 100830, 100880, 100930, 100940, 100900, 100810, 100690, 100630, 
    100520, 100400, 100230, 100110, 100020, 99950, 99880, 99770, 99680, 
    99580, 99480, 99410, 99340, 99280, 99230, 99190, 99190, 99190, 99230, 
    99260, 99300, 99370, 99460, 99550, 99630, 99700, 99780, 99830, 99920, 
    100000, 100070, 100150, 100220, 100270, 100350, 100430, 100490, 100560, 
    100590, 100630, 100650, 100670, 100680, 100690, 100690, 100660, 100630, 
    100610, 100590, 100580, 100540, 100520, 100530, 100550, 100580, 100620, 
    100640, 100700, 100730, 100770, 100810, 100870, 100940, 100980, 101010, 
    101060, 101110, 101120, 101180, 101170, 101160, 101180, 101190, 101190, 
    101170, 101190, 101170, 101140, 101110, 101060, 101010, 100880, 100710, 
    100650, 100540, 100470, 100410, 100360, 100310, 100260, 100200, 100190, 
    100220, 100200, 100180, 100210, 100200, 100190, 100180, 100180, 100200, 
    100210, 100260, 100250, 100240, 100210, 100180, 100180, 100140, 100140, 
    100100, 100110, 100120, 100060, 100070, 100090, 100200, 100240, 100300, 
    100320, 100350, 100580, 100700, 100760, 100850, 100890, 100970, 101070, 
    101160, 101260, 101380, 101690, 101800, 101910, 101970, 102070, 102290, 
    102360, 102470, 102490, 102560, 102600, 102610, 102600, 102550, 102530, 
    102470, 102440, 102380, 102350, 102320, 102290, 102300, 102250, 102280, 
    102250, 102200, 102130, 102060, 101880, 101840, 101780, 101760, 101690, 
    101730, 101740, 101770, 101820, 101880, 101880, 101860, 101840, 101790, 
    101830, 101840, 101830, 101830, 101850, 101820, 101820, 101820, 101800, 
    101730, 101710, 101700, 101660, 101670, 101640, 101600, 101540, 101570, 
    101560, 101550, 101580, 101580, 101570, 101540, 101510, 101530, 101530, 
    101570, 101560, 101580, 101580, 101590, 101590, 101600, 101600, 101600, 
    101610, 101630, 101650, 101690, 101690, 101670, 101700, 101720, 101750, 
    101750, 101760, 101770, 101740, 101740, 101730, 101740, 101730, 101700, 
    101700, 101680, 101680, 101680, 101670, 101680, 101680, 101680, 101670, 
    101680, 101680, 101700, 101720, 101750, 101760, 101770, 101770, 101770, 
    101760, 101760, 101760, 101790, 101800, 101810, 101750, 101770, 101770, 
    101770, 101760, 101750, 101750, 101750, 101740, 101730, 101710, 101720, 
    101720, 101720, 101710, 101720, 101720, 101700, 101690, 101670, 101670, 
    101670, 101660, 101660, 101640, 101620, 101600, 101590, 101570, 101540, 
    101510, 101500, 101470, 101400, 101090, 101120, 101130, 101120, 101120, 
    101140, 101160, 101170, 101200, 101200, 101200, 101220, 101240, 101260, 
    101270, 101310, 101310, 101320, 101350, 101370, 101390, 101430, 101470, 
    101500, 101540, 101560, 101570, 101590, 101600, 101580, 101560, 101570, 
    101560, 101550, 101510, 101490, 101480, 101510, 101510, 101510, 101510, 
    101520, 101520, 101530, 101540, 101500, 101500, 101510, 101520, 101480, 
    101480, 101480, 101490, 101490, 101490, 101480, 101470, 101470, 101420, 
    101400, 101400, 101410, 101390, 101390, 101350, 101340, 101330, 101320, 
    101320, 101300, 101310, 101310, 101290, 101290, 101310, 101330, 101340, 
    101340, 101350, 101380, 101380, 101410, 101420, 101460, 101470, 101470, 
    101500, 101520, 101530, 101560, 101600, 101620, 101600, 101630, 101660, 
    101690, 101730, 101760, 101770, 101770, 101780, 101780, 101800, 101830, 
    101840, 101840, 101830, 101810, 101810, 101800, 101790, 101770, 101790, 
    101770, 101770, 101740, 101720, 101700, 101680, 101670, 101660, 101570, 
    101530, 101510, 101490, 101480, 101460, 101430, 101400, 101380, 101340, 
    101310, 101280, 101250, 101240, 101200, 101190, 101170, 101150, 101140, 
    101110, 101080, 101020, 100980, 100940, 100900, 100870, 100840, 100810, 
    100770, 100740, 100710, 100610, 100580, 100550, 100550, 100530, 100520, 
    100510, 100510, 100510, 100500, 100490, 100490, 100480, 100440, 100420, 
    100420, 100450, 100460, 100470, 100460, 100480, 100470, 100470, 100480, 
    100500, 100520, 100540, 100580, 100600, 100630, 100650, 100670, 100680, 
    100700, 100690, 100700, 100710, 100730, 100750, 100770, 100790, 100790, 
    100790, 100820, 100840, 100850, 100850, 100860, 100880, 100890, 100930, 
    100960, 100970, 100980, 101000, 101030, 101050, 101070, 101080, 101110, 
    101150, 101280, 101280, 101320, 101350, 101390, 101400, 101420, 101430, 
    101470, 101510, 101530, 101580, 101610, 101620, 101650, 101660, 101680, 
    101690, 101680, 101690, 101690, 101700, 101710, 101710, 101710, 101690, 
    101630, 101610, 101590, 101580, 101590, 101590, 101590, 101590, 101570, 
    101560, 101550, 101530, 101500, 101490, 101480, 101440, 101420, 101410, 
    101390, 101360, 101320, 101300, 101300, 101290, 101280, 101240, 101220, 
    101190, 101140, 101100, 101090, 101060, 101020, 101010, 100970, 100950, 
    100940, 100950, 100940, 100940, 100890, 100880, 100900, 100920, 100950, 
    100980, 100990, 101020, 101040, 101090, 101120, 101160, 101190, 101220, 
    101250, 101280, 101310, 101330, 101350, 101350, 101370, 101380, 101400, 
    101430, 101450, 101470, 101500, 101500, 101500, 101490, 101480, 101500, 
    101500, 101500, 101520, 101510, 101520, 101510, 101480, 101460, 101440, 
    101430, 101420, 101410, 101390, 101380, 101370, 101350, 101340, 101300, 
    101280, 101270, 101250, 101250, 101230, 101210, 101210, 101200, 101220, 
    101230, 101210, 101210, 101210, 101200, 101200, 101190, 101220, 101230, 
    101230, 101220, 101180, 101180, 101140, 101070, 101050, 101050, 101040, 
    101000, 100960, 100930, 100900, 100850, 100790, 100790, 100770, 100760, 
    100730, 100720, 100700, 100660, 100600, 100580, 100510, 100480, 100440, 
    100400, 100370, 100340, 100310, 100290, 100250, 100220, 100180, 100140, 
    100090, 100040, 99970, 99930, 99870, 99820, 99790, 99680, 99620, 99600, 
    99580, 99570, 99530, 99500, 99500, 99500, 99510, 99520, 99550, 99570, 
    99570, 99590, 99600, 99590, 99600, 99620, 99630, 99670, 99730, 99740, 
    99770, 99810, 99790, 99820, 99820, 99850, 99850, 99890, 99930, 99960, 
    99990, 100030, 100060, 100090, 100120, 100150, 100170, 100350, 100390, 
    100420, 100470, 100570, 100600, 100800, 100810, 100820, 100840, 100870, 
    100890, 100900, 100900, 100960, 100980, 101000, 101000, 101010, 101050, 
    101080, 101110, 101140, 101160, 101170, 101220, 101240, 101250, 101280, 
    101290, 101290, 101340, 101400, 101440, 101450, 101470, 101490, 101510, 
    101540, 101600, 101620, 101700, 101720, 101770, 101790, 101810, 101840, 
    101870, 101870, 101890, 101890, 101930, 101960, 101990, 102010, 102020, 
    102060, 102060, 102050, 102050, 102060, 102060, 102060, 102060, 102050, 
    102060, 102050, 102030, 102020, 101990, 101960, 101940, 101920, 101900, 
    101860, 101850, 101850, 101830, 101810, 101790, 101750, 101720, 101690, 
    101670, 101650, 101640, 101620, 101600, 101570, 101550, 101530, 101510, 
    101490, 101460, 101450, 101430, 101400, 101400, 101380, 101350, 101330, 
    101320, 101290, 101280, 101240, 101210, 101170, 101180, 101210, 101220, 
    101230, 101240, 101230, 101210, 101200, 101180, 101170, 101170, 101150, 
    101150, 101130, 101120, 101130, 101130, 101110, 101080, 101060, 101050, 
    101020, 101000, 101000, 101000, 101000, 100990, 101000, 101020, 101020, 
    101010, 101010, 101020, 101020, 101000, 101010, 101010, 101030, _, 
    101090, 101110, 101110, 101140, 101170, 101160, 101200, 101200, 101230, 
    101240, _, 101300, 101320, 101360, 101380, 101420, _, 101490, 101530, _, 
    _, _, 101610, 101640, _, _, 101720, 101730, 101750, 101750, 101740, 
    101740, 101740, 101730, 101740, 101730, 101710, 101690, 101660, 101640, 
    101680, 101640, 101600, 101580, 101550, 101520, 101490, 101420, 101400, 
    101380, 101380, 101320, 101280, 101250, 101230, 101230, 101180, 101130, 
    101110, 101090, 101040, 101000, 100980, 100950, 100950, 100900, 100850, 
    100830, 100760, 100850, 100680, 100650, 100580, 100510, 100470, 100410, 
    100330, 100250, 100200, 100100, 100060, 100000, 99970, 99890, 99850, 
    99810, 99780, 99740, 99720, 99650, 99670, 99670, 99640, 99630, 99630, 
    99610, 99600, 99610, 99580, 99560, 99540, 99510, 99500, 99450, 99460, 
    99480, 99450, 99420, 99430, 99410, 99450, 99470, 99480, 99490, 99440, 
    99510, 99500, 99490, 99460, 99380, 99370, 99450, 99470, 99500, 99470, 
    99510, 99500, 99490, 99460, 99480, 99510, 99530, 99560, 99610, 99630, 
    99660, 99690, 99730, 99750, 99790, 99810, 99860, 99890, 99960, 99990, 
    100020, 100070, 100100, 100140, 100170, 100210, 100230, 100260, 100260, 
    100320, 100350, 100390, 100400, 100440, 100460, 100480, 100510, 100530, 
    100520, 100530, 100530, 100550, 100550, 100550, 100560, 100560, 100580, 
    100590, 100570, 100570, 100560, 100560, 100560, 100580, 100610, 100630, 
    100650, 100660, 100670, 100680, 100670, 100660, 100660, 100640, 100620, 
    100610, 100610, 100610, 100590, 100570, 100560, 100530, 100510, 100490, 
    100460, 100410, 100380, 100370, 100350, 100340, 100320, 100280, 100280, 
    100250, 100200, 100180, 100160, 100140, 100140, 100120, 100100, 100080, 
    100090, 100080, 100060, 100040, 100020, 100010, 100000, 99980, 99970, 
    99960, 99960, 99980, 99980, 99960, 99950, 99940, 99910, 99910, 99880, 
    99870, 99850, 99820, 99790, 99760, 99750, 99750, 99740, 99730, 99720, 
    99750, 99760, 99780, 99780, 99790, 99820, 99840, 99880, 99890, 99920, 
    99950, 99990, 100030, 100050, 100070, 100080, 100090, 100120, 100150, 
    100160, 100180, 100170, 100210, 100190, 100170, 100160, 100170, 100170, 
    100140, 100090, 100120, 100120, 100120, 100100, 100070, 99980, 99900, 
    99820, 99740, 99590, 99500, 99490, 99420, 99470, 99470, 99440, 99410, 
    99430, 99370, 99320, 99320, 99380, 99300, 99290, 99320, 99370, 99340, 
    99400, 99400, 99320, 99270, 99240, 99280, 99240, 99270, 99310, 99280, 
    99350, 99400, 99410, 99450, 99430, 99450, 99440, 99440, 99480, 99510, 
    99470, 99490, 99450, 99480, 99520, 99560, 99570, 99600, 99610, 99630, 
    99670, 99670, 99700, 99740, 99740, 99780, 99820, 99810, 99820, 99830, 
    99840, 99870, 99890, 99910, 99890, 99900, 99910, 99990, 100030, 100100, 
    100160, 100210, 100270, 100300, 100350, 100400, 100430, 100490, 100510, 
    100530, 100550, 100580, 100590, 100650, 100700, 100720, 100780, 100830, 
    100850, 100890, 100940, 100980, 101010, 101030, 101030, 101030, 101030, 
    101020, 101010, 100990, 100970, 100940, 100930, 100910, 100900, 100900, 
    100880, 100860, 100860, 100840, 100830, 100810, 100800, 100800, 100810, 
    100800, 100780, 100770, 100770, 100760, 100750, 100720, 100700, 100690, 
    100680, 100670, 100670, 100660, 100640, 100630, 100620, 100600, 100600, 
    100590, 100570, 100550, 100530, 100520, 100500, 100510, 100510, 100510, 
    100490, 100470, 100460, 100430, 100400, 100380, 100370, 100370, 100360, 
    100360, 100360, 100350, 100360, 100360, 100350, 100360, 100370, 100380, 
    100400, 100430, 100450, 100480, 100500, 100530, 100560, 100560, 100580, 
    100600, 100620, 100630, 100650, 100680, 100700, 100720, 100750, 100760, 
    100790, 100800, 100820, 100840, 100860, 100880, 100900, 100930, 100950, 
    100970, 100990, 101000, 101000, 101000, 101020, 101030, 101020, 101030, 
    101040, 101060, 101070, 101070, 101080, 101100, 101120, 101130, 101130, 
    101120, 101110, 101110, 101120, 101120, 101120, 101130, 101140, 101130, 
    101130, 101130, 101120, 101130, 101130, 101150, 101170, 101190, 101210, 
    101230, 101250, 101270, 101290, 101300, 101340, 101340, 101380, 101390, 
    101420, 101460, 101500, 101520, 101550, 101600, 101630, 101640, 101680, 
    101690, 101710, 101740, 101790, 101820, 101870, 101890, 101910, 101930, 
    101960, 101960, 101970, 101980, 101980, 102000, 102020, 102010, 102010, 
    102010, 102020, 102020, 102040, 102050, 102030, 102010, 102010, 102000, 
    102010, 102030, 102060, 102060, 102070, 102090, 102070, 102090, 102080, 
    102070, 102060, 102060, 102060, 102060, 102050, 102060, 102040, 102030, 
    102010, 101980, 101940, 101920, 101930, 101920, 101920, 101920, 101910, 
    101910, 101910, 101930, 101910, 101880, 101870, 101850, 101820, 101820, 
    101810, 101790, 101790, 101780, 101770, 101740, 101720, 101710, 101710, 
    101690, 101690, 101670, 101660, 101660, 101660, 101650, 101620, 101600, 
    101580, 101590, 101570, 101530, 101500, 101500, 101490, 101470, 101460, 
    101450, 101430, 101420, 101410, 101380, 101370, 101350, 101310, 101290, 
    101310, 101290, 101290, 101300, 101300, 101290, 101290, 101270, 101280, 
    101260, 101270, 101280, 101290, 101270, 101290, 101270, 101230, 101240, 
    101250, 101230, 101230, 101220, 101200, 101190, 101180, 101140, 101130, 
    101120, 101110, 101080, 101070, 101070, 101050, 101020, 101010, 100980, 
    100990, 100980, 100980, 100980, 100970, 100970, 100960, 100960, 100960, 
    100970, 100980, 101000, 101030, 101050, 101070, 101090, 101120, 101160, 
    101190, 101220, 101230, 101260, 101280, 101310, 101340, 101360, 101410, 
    101430, 101470, 101500, 101520, 101540, 101570, 101580, 101590, 101590, 
    101600, 101630, 101640, 101660, 101650, 101650, 101640, 101630, 101620, 
    101630, 101620, 101620, 101640, 101630, 101650, 101650, 101660, 101670, 
    101670, 101660, 101650, 101630, 101620, 101600, 101590, 101580, 101590, 
    101600, 101610, 101580, 101550, 101540, 101550, 101540, 101560, 101560, 
    101570, 101600, 101650, 101670, 101680, 101690, 101720, 101720, 101750, 
    101750, 101760, 101760, 101760, 101760, 101780, 101810, 101810, 101820, 
    101840, 101850, 101850, 101850, 101860, 101870, 101900, 101890, 101900, 
    101910, 101920, 101900, 101870, 101840, 101820, 101770, 101730, 101720, 
    101720, 101690, 101670, 101650, 101630, 101600, 101590, 101550, 101520, 
    101480, 101460, 101430, 101410, 101410, 101390, 101370, 101370, 101330, 
    101300, 101300, 101280, 101290, 101280, 101290, 101310, 101340, 101340, 
    101370, 101390, 101390, 101400, 101400, 101430, 101450, 101480, 101480, 
    101530, 101550, 101590, 101620, 101650, 101660, 101690, 101740, 101770, 
    101770, 101780, 101810, 101840, 101880, 101900, 101930, 101930, 101940, 
    101940, 101950, 101940, 101940, 101940, 101940, 101960, 101980, 102020, 
    102020, 102040, 102060, 102060, 102080, 102100, 102120, 102130, 102150, 
    102150, 102160, 102170, 102170, 102180, 102190, 102230, 102240, 102240, 
    102260, 102260, 102300, 102320, 102350, 102380, 102390, 102410, 102430, 
    102450, 102450, 102480, 102490, 102500, 102520, 102510, 102510, 102520, 
    102530, 102530, 102540, 102550, 102560, 102550, 102530, 102530, 102520, 
    102500, 102480, 102470, 102450, 102470, 102460, 102430, 102380, 102380, 
    102360, 102360, 102300, 102290, 102280, 102280, 102270, 102260, 102220, 
    102210, 102200, 102140, 102110, 102070, 102000, 101950, 101900, 101870, 
    101840, 101820, 101810, 101800, 101760, 101770, 101750, 101740, 101750, 
    101720, 101760, 101760, 101770, 101800, 101810, 101820, 101840, 101870, 
    101880, 101890, 101940, 101950, 101950, 102010, 102050, 102050, 102090, 
    102120, 102130, 102120, 102130, 102110, 102120, 102130, 102130, 102140, 
    102130, 102140, 102140, 102150, 102160, 102150, 102140, 102160, 102170, 
    102180, 102170, 102170, 102150, 102150, 102140, 102130, 102130, 102120, 
    102130, 102110, 102110, 102080, 102100, 102080, 102080, 102100, 102080, 
    102070, 102080, 102070, 102050, 102040, 102010, 102020, 102030, 102050, 
    102040, 102010, 102000, 101990, 101990, 101970, 101950, 101950, 101950, 
    101960, 101980, 101970, 101990, 102000, 102000, 101980, 101960, 101970, 
    102000, 102040, 102050, 102060, 102070, 102080, 102090, 102090, 102110, 
    102120, 102120, 102110, 102130, 102150, 102170, 102190, 102210, 102220, 
    102230, 102230, 102230, 102230, 102230, 102230, 102230, 102230, 102230, 
    102230, 102250, 102250, 102230, 102220, 102210, 102200, 102200, 102200, 
    102190, 102190, 102190, 102170, 102150, 102130, 102120, 102110, 102100, 
    102090, 102060, 102030, 102000, 101980, 101950, 101930, 101920, 101890, 
    101870, 101850, 101830, 101800, 101760, 101740, 101730, 101680, 101650, 
    101620, 101610, 101590, 101560, 101530, 101500, 101470, 101460, 101430, 
    101400, 101390, 101360, 101350, 101320, 101300, 101290, 101290, 101290, 
    101280, 101270, 101260, 101250, 101230, 101210, 101200, 101200, 101210, 
    101210, 101200, 101200, 101180, 101160, 101120, 101080, 101060, 101010, 
    101030, 101030, 101020, 100990, 100970, 100940, 100910, 100870, 100780, 
    100700, 100630, 100600, 100590, 100580, 100630, 100590, 100690, 100710, 
    100760, 100770, 100800, 100780, 100820, 100810, 100850, 100820, 100820, 
    100790, 100830, 100910, 100930, 100960, 100940, 100970, 100980, 101010, 
    101070, 101080, 101130, 101120, 101140, 101150, 101130, 101150, 101170, 
    101180, 101210, 101230, 101260, 101260, 101270, 101260, 101270, 101260, 
    101260, 101260, 101260, 101260, 101270, 101290, 101310, 101320, 101330, 
    101350, 101350, 101370, 101390, 101400, 101380, 101350, 101350, 101310, 
    101300, 101260, 101250, 101240, 101240, 101250, 101240, 101270, 101260, 
    101250, 101230, 101260, 101270, 101270, 101270, 101300, 101310, 101330, 
    101350, 101360, 101360, 101360, 101350, 101350, 101370, 101410, 101420, 
    101430, 101450, 101470, 101470, 101500, 101480, 101480, 101490, 101500, 
    101510, 101500, 101510, 101540, 101550, 101550, 101530, 101530, 101540, 
    101520, 101510, 101510, 101510, 101540, 101550, 101560, 101570, 101570, 
    101560, 101560, 101550, 101530, 101540, 101530, 101500, 101490, 101490, 
    101490, 101490, 101490, 101490, 101480, 101480, 101460, 101440, 101410, 
    101400, 101390, 101360, 101350, 101350, 101350, 101350, 101360, 101360, 
    101340, 101340, 101330, 101340, 101330, 101340, 101340, 101340, 101340, 
    101350, 101340, 101340, 101310, 101290, 101270, 101260, 101270, 101240, 
    101230, 101200, 101190, 101130, 101110, 101080, 101040, 100980, 100970, 
    100920, 100920, 100880, 100830, 100780, 100750, 100730, 100700, 100640, 
    100570, 100530, 100470, 100510, 100450, 100430, 100400, 100380, 100390, 
    100360, 100330, 100310, 100280, 100260, 100250, 100220, 100270, 100270, 
    100250, 100240, 100230, 100220, 100210, 100210, 100180, 100180, 100180, 
    100170, 100140, 100140, 100140, 100140, 100140, 100140, 100130, 100140, 
    100140, 100150, 100160, 100170, 100210, 100220, 100230, 100250, 100270, 
    100290, 100320, 100350, 100390, 100400, 100440, 100470, 100490, 100530, 
    100570, 100600, 100640, 100680, 100710, 100760, 100810, 100840, 100880, 
    100940, 101000, 101050, 101100, 101150, 101220, 101270, 101310, 101350, 
    101400, 101450, 101480, 101510, 101550, 101600, 101630, 101660, 101690, 
    101720, 101760, 101790, 101810, 101840, 101860, 101880, 101900, 101930, 
    101970, 101990, 101990, 102000, 102000, 101990, 102000, 102010, 102010, 
    102030, 102040, 102050, 102050, 102050, 102050, 102030, 102030, 102000, 
    101970, 101960, 101950, 101940, 101910, 101910, 101860, 101820, 101850, 
    101820, 101800, 101810, 101750, 101720, 101700, 101670, 101640, 101580, 
    101560, 101480, 101390, 101370, 101400, 101400, 101320, 101250, 101210, 
    101190, 101170, 101140, 101130, 101140, 101100, 101150, 101150, 101160, 
    101180, 101200, 101230, 101220, 101250, 101250, 101270, 101290, 101310, 
    101320, 101330, 101350, 101360, 101400, 101440, 101470, 101510, 101540, 
    101560, 101580, 101620, 101650, 101680, 101710, 101740, 101770, 101790, 
    101810, 101850, 101870, 101890, 101900, 101890, 101910, 101920, 101920, 
    101920, 101910, 101920, 101940, 101960, 101960, 101980, 101990, 101990, 
    101970, 101970, 101980, 101960, 101950, 101930, 101900, 101890, 101910, 
    101900, 101890, 101850, 101860, 101840, 101820, 101820, 101820, 101780, 
    101790, 101840, 101850, 101860, 101880, 101910, 101910, 101930, 101910, 
    101900, 101910, 101940, 101970, 101980, 101990, 101990, 102000, 102020, 
    102020, 102020, 102030, 102010, 102000, 101990, 102010, 102030, 102060, 
    102070, 102070, 102050, 102040, 102020, 102020, 102000, 101990, 101960, 
    101950, 101950, 101960, 101950, 101960, 101950, 101950, 101930, 101890, 
    101840, 101830, 101820, 101820, 101840, 101840, 101840, 101820, 101800, 
    101780, 101760, 101750, 101770, 101750, 101740, 101750, 101750, 101760, 
    101770, 101770, 101770, 101790, 101800, 101810, 101820, 101840, 101890, 
    101920, 101940, 101970, 101990, 102000, 102020, 102040, 102050, 102070, 
    102080, 102100, 102110, 102120, 102150, 102160, 102160, 102170, 102160, 
    102160, 102160, 102160, 102150, 102130, 102100, 102080, 102070, 102050, 
    102000, 102000, 101970, 101940, 101900, 101860, 101850, 101790, 101740, 
    101680, 101660, 101650, 101610, 101570, 101540, 101430, 101410, 101340, 
    101290, 101250, 101220, 101200, 101190, 101180, 101160, 101140, 101120, 
    101120, 101100, 101090, 101060, 101040, 101020, 101010, 100980, 100960, 
    100960, 100940, 100920, 100920, 100890, 100890, 100880, 100880, 100870, 
    100870, 100870, 100880, 100900, 100880, 100880, 100890, 100890, 100890, 
    100890, 100880, 100890, 100900, 100900, 100930, 100950, 100970, 100980, 
    101000, 101010, 100990, 101010, 101020, 101020, 101020, 101040, 101050, 
    101060, 101060, 101060, 101070, 101080, 101060, 101040, 101020, 101040, 
    101050, 101050, 101040, 101040, 101050, 101040, 101020, 101010, 100990, 
    100990, 100980, 100960, 100960, 100970, 100970, 100960, 100980, 100980, 
    100980, 100990, 100980, 100990, 100980, 100990, 101000, 101000, 101000, 
    101030, 101040, 101050, 101060, 101050, 101050, 101050, 101050, 101050, 
    101070, 101090, 101110, 101140, 101160, 101170, 101180, 101210, 101220, 
    101240, 101250, 101260, 101280, 101290, 101310, 101340, 101350, 101360, 
    101380, 101380, 101380, 101380, 101380, 101370, 101380, 101380, 101380, 
    101390, 101390, 101390, 101370, 101390, 101390, 101370, 101350, 101360, 
    101380, 101370, 101370, 101360, 101350, 101350, 101330, 101300, 101280, 
    101290, 101290, 101310, 101320, 101330, 101330, 101330, 101330, 101320, 
    101300, 101280, 101270, 101250, 101230, 101210, 101190, 101180, 101160, 
    101160, 101140, 101120, 101090, 101060, 101030, 100990, 100960, 100950, 
    100940, 100940, 100930, 100910, 100890, 100890, 100880, 100880, 100900, 
    100890, 100880, 100890, 100900, 100910, 100900, 100920, 100930, 100950, 
    100980, 101010, 101030, 101060, 101090, 101120, 101170, 101210, 101270, 
    101340, 101400, 101450, 101520, 101570, 101620, 101660, 101690, 101730, 
    101800, 101840, 101910, 101990, 102050, 102080, 102130, 102180, 102220, 
    102250, 102270, 102300, 102320, 102370, 102400, 102420, 102450, 102490, 
    102490, 102470, 102480, 102500, 102510, 102540, 102540, 102580, 102600, 
    102630, 102650, 102660, 102660, 102670, 102670, 102670, 102660, 102650, 
    102620, 102600, 102590, 102570, 102580, 102550, 102520, 102460, 102430, 
    102430, 102410, 102370, 102360, 102360, 102360, 102350, 102320, 102320, 
    102280, 102240, 102200, 102150, 102110, 102050, 102020, 101970, 101920, 
    101890, 101880, 101840, 101830, 101780, 101750, 101710, 101640, 101560, 
    101480, 101450, 101400, 101390, 101360, 101350, 101300, 101280, 101210, 
    101200, 101200, 101190, 101150, 101150, 101170, 101160, 101140, 101190, 
    101190, 101170, 101190, 101180, 101150, 101130, 101110, 101110, 101100, 
    101110, 101100, 101100, 101130, 101130, 101120, 101110, 101110, 101130, 
    101150, 101160, 101180, 101180, 101170, 101170, 101190, 101100, 101020, 
    100950, 100890, 100920, 100910, 100940, 100920, 100930, 100980, 100980, 
    101000, 101030, 101050, 101050, 101070, 101070, 101070, 101100, 101130, 
    101140, 101140, 101120, 101110, 101100, 101130, 101110, 101120, 101130, 
    101130, 101150, 101190, 101210, 101230, 101250, 101290, 101350, 101410, 
    101440, 101490, 101550, 101600, 101670, 101690, 101740, 101780, 101810, 
    101850, 101900, 101920, 101950, 101990, 102020, 102060, 102120, 102150, 
    102170, 102210, 102220, 102260, 102280, 102290, 102310, 102320, 102340, 
    102380, 102420, 102430, 102470, 102490, 102490, 102520, 102540, 102540, 
    102540, 102540, 102560, 102550, 102580, 102580, 102570, 102580, 102570, 
    102530, 102500, 102460, 102440, 102370, 102330, 102240, 102210, 102180, 
    102060, 101980, 101900, 101810, 101720, 101650, 101550, 101460, 101400, 
    101370, 101360, 101350, 101330, 101300, 101290, 101290, 101280, 101260, 
    101290, 101290, 101280, 101290, 101300, 101320, 101320, 101350, 101350, 
    101350, 101360, 101380, 101370, 101370, 101390, 101400, 101430, 101460, 
    101480, 101500, 101530, 101540, 101550, 101560, 101600, 101600, 101620, 
    101630, 101650, 101660, 101700, 101690, 101690, 101680, 101690, 101710, 
    101710, 101720, 101700, 101720, 101750, 101750, 101750, 101780, 101790, 
    101780, 101780, 101790, 101790, 101780, 101780, 101770, 101770, 101770, 
    101760, 101760, 101760, 101760, 101740, 101720, 101710, 101690, 101660, 
    101640, 101620, 101610, 101590, 101580, 101560, 101540, 101540, 101540, 
    101540, 101520, 101510, 101510, 101520, 101520, 101540, 101560, 101560, 
    101590, 101600, 101590, 101590, 101600, 101610, 101620, 101620, 101640, 
    101660, 101670, 101680, 101690, 101690, 101680, 101670, 101660, 101650, 
    101660, 101690, 101680, 101700, 101720, 101740, 101710, 101690, 101690, 
    101670, 101670, 101670, 101650, 101660, 101650, 101630, 101590, 101610, 
    101590, 101530, 101490, 101440, 101370, 101320, 101290, 101290, 101230, 
    101190, 101120, 101080, 101070, 101050, 100990, 100920, 100920, 100910, 
    100870, 100860, 100830, 100810, 100770, 100760, 100750, 100750, 100750, 
    100790, 100780, 100780, 100800, 100810, 100850, 100860, 100870, 100900, 
    100890, 100910, 100900, 100890, 100880, 100860, 100850, 100840, 100850, 
    100820, 100800, 100790, 100770, 100750, 100740, 100710, 100670, 100680, 
    100680, 100680, 100670, 100650, 100630, 100600, 100600, 100590, 100610, 
    100620, 100600, 100590, 100640, 100650, 100650, 100690, 100710, 100750, 
    100780, 100780, 100820, 100850, 100890, 100950, 100970, 101060, 101070, 
    101110, 101200, 101240, 101300, 101360, 101400, 101430, 101500, 101520, 
    101540, 101570, 101620, 101650, 101700, 101710, 101750, 101770, 101800, 
    101840, 101860, 101890, 101910, 101930, 101930, 101930, 101940, 101940, 
    101940, 101930, 101920, 101890, 101880, 101850, 101830, 101810, 101820, 
    101800, 101780, 101750, 101730, 101690, 101670, 101630, 101570, 101530, 
    101500, 101460, 101400, 101360, 101330, 101280, 101250, 101210, 101190, 
    101150, 101090, 101050, 101010, 101000, 100980, 100960, 100950, 100930, 
    100920, 100900, 100900, 100910, 100880, 100870, 100840, 100850, 100860, 
    100870, 100820, 100830, 100830, 100800, 100760, 100710, 100670, 100630, 
    100600, 100590, 100560, 100530, 100510, 100490, 100480, 100480, 100470, 
    100450, 100440, 100430, 100440, 100440, 100450, 100470, 100490, 100500, 
    100510, 100530, 100550, 100570, 100580, 100610, 100650, 100680, 100730, 
    100770, 100790, 100820, 100850, 100870, 100900, 100910, 100930, 100940, 
    100960, 100980, 101000, 101000, 101010, 101010, 101000, 100990, 101000, 
    100990, 100970, 100970, 100960, 100950, 100960, 100950, 100940, 100930, 
    100910, 100890, 100870, 100870, 100860, 100830, 100810, 100780, 100770, 
    100720, 100670, 100610, 100580, 100550, 100510, 100440, 100410, 100340, 
    100260, 100180, 100110, 100070, 99950, 99850, 99730, 99650, 99590, 99590, 
    99610, 99640, 99690, 99760, 99790, 99840, 99880, 99900, 99930, 99970, 
    99990, 99980, 100020, 100070, 100110, 100110, 100130, 100170, 100210, 
    100220, 100220, 100210, 100250, 100260, 100270, 100280, 100320, 100350, 
    100390, 100400, 100410, 100440, 100450, 100480, 100480, 100460, 100500, 
    100530, 100560, 100610, 100690, 100740, 100800, 100860, 100940, 100990, 
    101040, 101080, 101100, 101130, 101160, 101120, 101200, 101170, 101140, 
    101150, 101090, 101030, 100950, 100910, 100840, 100780, 100750, 100740, 
    100740, 100730, 100730, 100740, 100760, 100780, 100790, 100760, 100760, 
    100780, 100810, 100810, 100850, 100880, 100880, 100880, 100860, 100850, 
    100820, 100770, 100720, 100690, 100610, 100590, 100550, 100490, 100390, 
    100330, 100300, 100280, 100290, 100330, 100320, 100390, 100420, 100540, 
    100580, 100650, 100700, 100740, 100790, 100850, 100920, 101000, 101100, 
    101160, 101230, 101270, 101290, 101300, 101320, 101360, 101340, 101320, 
    101290, 101290, 101270, 101250, 101230, 101200, 101180, 101170, 101160, 
    101140, 101120, 101140, 101210, 101230, 101260, 101270, 101340, 101380, 
    101420, 101410, 101470, 101490, 101510, 101550, 101560, 101560, 101570, 
    101590, 101600, 101590, 101610, 101590, 101580, 101560, 101540, 101500, 
    101460, 101420, 101360, 101320, 101260, 101230, 101220, 101180, 101140, 
    101080, 101030, 101000, 100980, 100960, 100940, 100940, 100920, 100930, 
    100960, 100970, 100980, 101000, 101010, 101060, 101090, 101140, 101230, 
    101270, 101320, 101380, 101440, 101500, 101530, 101600, 101620, 101650, 
    101670, 101690, 101700, 101740, 101760, 101780, 101780, 101790, 101800, 
    101780, 101780, 101750, 101730, 101710, 101710, 101720, 101700, 101680, 
    101660, 101650, 101620, 101610, 101580, 101540, 101530, 101500, 101460, 
    101400, 101360, 101340, 101310, 101260, 101220, 101200, 101170, 101160, 
    101130, 101140, 101120, 101120, 101130, 101140, 101170, 101170, 101170, 
    101190, 101220, 101220, 101230, 101260, 101260, 101270, 101270, 101290, 
    101300, 101310, 101330, 101330, 101370, 101370, 101360, 101370, 101390, 
    101370, 101360, 101360, 101370, 101380, 101390, 101410, 101420, 101400, 
    101380, 101360, 101320, 101290, 101310, 101300, 101310, 101310, 101300, 
    101260, 101240, 101210, 101210, 101220, 101220, 101230, 101250, 101290, 
    101300, 101300, 101280, 101280, 101290, 101280, 101270, 101270, 101230, 
    101200, 101200, 101220, 101220, 101190, 101210, 101210, 101220, 101210, 
    101190, 101170, 101160, 101160, 101150, 101150, 101150, 101160, 101160, 
    101170, 101180, 101180, 101190, 101200, 101180, 101210, 101260, 101300, 
    101340, 101360, 101400, 101450, 101490, 101530, 101530, 101530, 101550, 
    101550, 101600, 101660, 101710, 101730, 101770, 101780, 101770, 101750, 
    101750, 101740, 101720, 101700, 101670, 101650, 101630, 101590, 101550, 
    101500, 101460, 101400, 101340, 101300, 101260, 101220, 101160, 101140, 
    101140, 101080, 101060, 101030, 100990, 100940, 100900, 100890, 100860, 
    100840, 100870, 100890, 100870, 100870, 100840, 100840, 100840, 100850, 
    100850, 100850, 100880, 100920, 100930, 100920, 100930, 100940, 100980, 
    101010, 101020, 101030, 101030, 101050, 101050, 101090, 101100, 101120, 
    101130, 101130, 101120, 101120, 101110, 101110, 101110, 101120, 101140, 
    101150, 101140, 101150, 101160, 101160, 101160, 101160, 101150, 101150, 
    101140, 101150, 101140, 101140, 101130, 101130, 101150, 101150, 101140, 
    101140, 101140, 101130, 101130, 101130, 101140, 101170, 101170, 101200, 
    101230, 101240, 101260, 101260, 101280, 101300, 101310, 101330, 101360, 
    101400, 101400, 101430, 101460, 101480, 101510, 101520, 101540, 101570, 
    101600, 101630, 101660, 101680, 101730, 101790, 101820, 101860, 101900, 
    101920, 101940, 101970, 102010, 102050, 102100, 102150, 102170, 102200, 
    102210, 102250, 102270, 102300, 102330, 102350, 102390, 102430, 102450, 
    102470, 102510, 102550, 102580, 102600, 102630, 102650, 102670, 102680, 
    102710, 102710, 102710, 102690, 102650, 102640, 102630, 102630, 102590, 
    102530, 102470, 102400, 102330, 102240, 102170, 102070, 101990, 101910, 
    101820, 101710, 101610, 101520, 101400, 101300, 101180, 101070, 100980, 
    100930, 100870, 100820, 100800, 100750, 100680, 100600, 100510, 100400, 
    100310, 100180, 100110, 99980, 99850, 99680, 99500, 99300, 99060, 98750, 
    98410, 98060, 97760, 97410, 97110, 96900, 96670, 96540, 96490, 96490, 
    96470, 96470, 96500, 96510, 96580, 96660, 96760, 96890, 97030, 97190, 
    97370, 97540, 97700, 97820, 97970, 98120, 98230, 98330, 98440, 98550, 
    98660, 98730, 98820, 98900, 98950, 99010, 99060, 99080, 99140, 99190, 
    99230, 99270, 99280, 99330, 99370, 99410, 99430, 99440, 99460, 99480, 
    99490, 99520, 99540, 99540, 99530, 99540, 99570, 99570, 99570, 99600, 
    99570, 99580, 99590, 99600, 99590, 99600, 99600, 99630, 99660, 99670, 
    99690, 99720, 99740, 99750, 99760, 99790, 99810, 99810, 99840, 99840, 
    99870, 99890, 99900, 99930, 99960, 99980, 100010, 100040, 100060, 100100, 
    100140, 100180, 100220, 100270, 100320, 100340, 100370, 100400, 100430, 
    100450, 100480, 100500, 100510, 100530, 100550, 100600, 100610, 100630, 
    100670, 100700, 100740, 100740, 100760, 100810, 100830, 100880, 100940, 
    100980, 101020, 101060, 101110, 101160, 101200, 101240, 101280, 101330, 
    101360, 101420, 101480, 101530, 101570, 101620, 101680, 101740, 101790, 
    101860, 101910, 101970, 102020, 102080, 102130, 102180, 102230, 102300, 
    102380, 102400, 102410, 102430, 102490, 102490, 102530, 102550, 102590, 
    102600, 102620, 102630, 102650, 102660, 102610, 102610, 102590, 102570, 
    102570, 102580, 102590, 102600, 102610, 102620, 102620, 102640, 102680, 
    102660, 102660, 102690, 102710, 102740, 102760, 102760, 102770, 102760, 
    102780, 102820, 102820, 102820, 102850, 102870, 102920, 102940, 102990, 
    103030, 103020, 103030, 103040, 103060, 103070, 103080, 103050, 103050, 
    103040, 103040, 103070, 103060, 103030, 102990, 102980, 102970, 102960, 
    102950, 102940, 102920, 102910, 102910, 102910, 102900, 102890, 102870, 
    102840, 102810, 102800, 102770, 102730, 102720, 102730, 102690, 102680, 
    102660, 102650, 102630, 102590, 102570, 102530, 102490, 102430, 102400, 
    102410, 102410, 102410, 102410, 102380, 102360, 102370, 102380, 102370, 
    102330, 102320, 102280, 102240, 102210, 102190, 102140, 102110, 102090, 
    102040, 102000, 101960, 101920, 101890, 101860, 101820, 101790, 101750, 
    101720, 101670, 101610, 101550, 101490, 101430, 101370, 101270, 101190, 
    101110, 101030, 100950, 100920, 100860, 100810, 100810, 100780, 100750, 
    100710, 100670, 100640, 100600, 100560, 100540, 100500, 100440, 100400, 
    100370, 100320, 100300, 100280, 100240, 100230, 100220, 100210, 100210, 
    100220, 100210, 100230, 100260, 100290, 100320, 100360, 100400, 100430, 
    100470, 100510, 100550, 100590, 100610, 100630, 100650, 100650, 100680, 
    100690, 100710, 100730, 100740, 100740, 100740, 100750, 100760, 100760, 
    100760, 100770, 100770, 100780, 100780, 100800, 100800, 100820, 100830, 
    100860, 100890, 100920, 100930, 100970, 100980, 100990, 100990, 101030, 
    101050, 101070, 101100, 101130, 101140, 101130, 101140, 101110, 101060, 
    101030, 100990, 100930, 100860, 100830, 100760, 100720, 100660, 100590, 
    100510, 100440, 100400, 100380, 100330, 100330, 100320, 100290, 100270, 
    100220, 100200, 100180, 100140, 100050, 99960, 99930, 99860, 99730, 
    99600, 99460, 99380, 99280, 99170, 99050, 98940, 98840, 98750, 98640, 
    98530, 98410, 98330, 98250, 98190, 98130, 98050, 97990, 97990, 98020, 
    98010, 98060, 98130, 98180, 98250, 98340, 98420, 98500, 98580, 98650, 
    98700, 98780, 98850, 98900, 98980, 99040, 99100, 99170, 99240, 99310, 
    99370, 99430, 99480, 99560, 99620, 99680, 99740, 99800, 99860, 99940, 
    100020, 100090, 100160, 100210, 100250, 100300, 100360, 100390, 100380, 
    100430, 100430, 100460, 100510, 100500, 100520, 100520, 100540, 100530, 
    100520, 100560, 100520, 100510, 100510, 100490, 100470, 100430, 100380, 
    100330, 100250, 100180, 100080, 100010, 99920, 99860, 99770, 99720, 
    99670, 99600, 99510, 99420, 99410, 99370, 99330, 99280, 99250, 99190, 
    99170, 99130, 99100, 99100, 99100, 99070, 99080, 99140, 99140, 99170, 
    99190, 99210, 99260, 99360, 99440, 99480, 99570, 99630, 99740, 99820, 
    99930, 100020, 100100, 100210, 100300, 100380, 100450, 100530, 100580, 
    100610, 100650, 100660, 100700, 100710, 100730, 100710, 100700, 100670, 
    100640, 100610, 100590, 100570, 100550, 100500, 100440, 100390, 100360, 
    100340, 100300, 100260, 100220, 100170, 100130, 100060, 100010, 99960, 
    99940, 99910, 99870, 99840, 99800, 99750, 99710, 99700, 99670, 99610, 
    99560, 99510, 99490, 99500, 99480, 99450, 99400, 99410, 99420, 99430, 
    99440, 99420, 99400, 99400, 99390, 99400, 99380, 99380, 99370, 99350, 
    99360, 99350, 99350, 99350, 99360, 99370, 99370, 99360, 99380, 99370, 
    99380, 99410, 99400, 99410, 99400, 99380, 99380, 99340, 99330, 99280, 
    99260, 99260, 99240, 99210, 99210, 99130, 99090, 99080, 99050, 98980, 
    98950, 98950, 98910, 98890, 98920, 98910, 98880, 98860, 98790, 98720, 
    98630, 98530, 98410, 98310, 98220, 98130, 98030, 97940, 97890, 97880, 
    97790, 97710, 97650, 97620, 97580, 97530, 97500, 97500, 97510, 97570, 
    97580, 97650, 97710, 97770, 97860, 97920, 98000, 98090, 98190, 98270, 
    98370, 98440, 98540, 98650, 98730, 98820, 98910, 98980, 99040, 99120, 
    99170, 99240, 99330, 99410, 99510, 99610, 99680, 99730, 99800, 99880, 
    99980, 100050, 100120, 100170, 100250, 100320, 100370, 100440, 100490, 
    100540, 100570, 100610, 100640, 100640, 100670, 100680, 100710, 100730, 
    100760, 100780, 100800, 100810, 100810, 100800, 100790, 100800, 100810, 
    100820, 100840, 100850, 100900, 100920, 100950, 101000, 101060, 101110, 
    101150, 101190, 101230, 101310, 101390, 101440, 101470, 101520, 101580, 
    101660, 101710, 101760, 101800, 101850, 101890, 101910, 101910, 101960, 
    101970, 102010, 102020, 102010, 101990, 101940, 101890, 101850, 101830, 
    101800, 101800, 101790, 101780, 101760, 101770, 101750, 101740, 101710, 
    101700, 101690, 101690, 101640, 101620, 101560, 101480, 101440, 101350, 
    101280, 101200, 101130, 101080, 101010, 100920, 100810, 100740, 100700, 
    100700, 100700, 100700, 100700, 100690, 100700, 100760, 100780, 100800, 
    100790, 100770, 100790, 100720, 100710, 100710, 100710, 100680, 100650, 
    100610, 100570, 100540, 100530, 100560, 100580, 100590, 100610, 100570, 
    100540, 100510, 100460, 100380, 100310, 100180, 100110, 99970, 99910, 
    99780, 99580, 99440, 99350, 99220, 99070, 98960, 98850, 98730, 98600, 
    98540, 98460, 98400, 98360, 98330, 98280, 98270, 98270, 98280, 98260, 
    98270, 98270, 98270, 98290, 98320, 98330, 98340, 98340, 98360, 98410, 
    98450, 98440, 98440, 98440, 98480, 98520, 98570, 98570, 98600, 98650, 
    98710, 98730, 98760, 98810, 98880, 98920, 99000, 99070, 99130, 99190, 
    99260, 99310, 99360, 99400, 99450, 99460, 99490, 99520, 99540, 99570, 
    99610, 99640, 99630, 99610, 99610, 99590, 99610, 99610, 99590, 99550, 
    99540, 99530, 99520, 99490, 99500, 99500, 99520, 99520, 99520, 99550, 
    99560, 99570, 99620, 99670, 99720, 99750, 99800, 99850, 99940, 99980, 
    100050, 100080, 100120, 100180, 100250, 100300, 100350, 100410, 100480, 
    100550, 100610, 100680, 100710, 100750, 100820, 100870, 100940, 100990, 
    101050, 101110, 101160, 101230, 101240, 101320, 101380, 101420, 101450, 
    101480, 101500, 101550, 101580, 101590, 101640, 101680, 101690, 101670, 
    101700, 101720, 101720, 101710, 101710, 101700, 101710, 101680, 101660, 
    101650, 101650, 101580, 101570, 101520, 101480, 101440, 101420, 101400, 
    101380, 101340, 101330, 101310, 101250, 101200, 101130, 101090, 101030, 
    100980, 100960, 100960, 100940, 100910, 100840, 100800, 100790, 100740, 
    100700, 100630, 100570, 100520, 100480, 100430, 100360, 100380, 100340, 
    100240, 100150, 100030, 99950, 99880, 99790, 99720, 99650, 99570, 99490, 
    99400, 99310, 99240, 99190, 99120, 99070, 99040, 99000, 98960, 98970, 
    98960, 98970, 98960, 98940, 98930, 98920, 98960, 98950, 98920, 98910, 
    98900, 98930, 98970, 98990, 99050, 99110, 99130, 99130, 99150, 99170, 
    99200, 99230, 99220, 99230, 99260, 99280, 99310, 99290, 99260, 99240, 
    99230, 99210, 99180, 99180, 99170, 99160, 99170, 99180, 99200, 99150, 
    99200, 99170, 99110, 99170, 99150, 99070, 99060, 99030, 99090, 99140, 
    99160, 99190, 99240, 99330, 99350, 99390, 99440, 99480, 99590, 99670, 
    99750, 99810, 99910, 99980, 100000, 100080, 100130, 100190, 100250, 
    100330, 100380, 100430, 100490, 100560, 100630, 100680, 100720, 100760, 
    100790, 100860, 100910, 100950, 101010, 101050, 101120, 101220, 101270, 
    101350, 101420, 101460, 101510, 101570, 101610, 101640, 101720, 101760, 
    101820, 101880, 101920, 101950, 101970, 102000, 102050, 102070, 102080, 
    102080, 102100, 102080, 102090, 102110, 102090, 102110, 102100, 102050, 
    102020, 101990, 101940, 101930, 101900, 101880, 101850, 101830, 101780, 
    101750, 101720, 101690, 101570, 101480, 101420, 101380, 101260, 101240, 
    101190, 101140, 101100, 101040, 101000, 100940, 100900, 100850, 100780, 
    100720, 100600, 100520, 100470, 100400, 100290, 100240, 100130, 100020, 
    99930, 99790, 99660, 99500, 99370, 99290, 99210, 99120, 99060, 99010, 
    98960, 98910, 98880, 98890, 98910, 98910, 98900, 98900, 98890, 98890, 
    98900, 98930, 98900, 98900, 98890, 98900, 98880, 98900, 98890, 98930, 
    98950, 98950, 98930, 98950, 98950, 98920, 98900, 98880, 98870, 98870, 
    98880, 98870, 98890, 98910, 98930, 98960, 98980, 98980, 99010, 99020, 
    99020, 99030, 99030, 99060, 99090, 99110, 99120, 99120, 99110, 99110, 
    99120, 99140, 99160, 99180, 99210, 99260, 99300, 99360, 99410, 99470, 
    99500, 99520, 99560, 99600, 99610, 99650, 99710, 99740, 99790, 99830, 
    99900, 99920, 99930, 99970, 99990, 100030, 100040, 100040, 100060, 
    100070, 100060, 100090, 100080, 100050, 100050, 100030, 100030, 100010, 
    100000, 99970, 99960, 99960, 99960, 99940, 99940, 99900, 99860, 99810, 
    99770, 99720, 99670, 99610, 99580, 99550, 99510, 99480, 99480, 99440, 
    99410, 99390, 99400, 99390, 99380, 99350, 99330, 99350, 99320, 99330, 
    99330, 99330, 99330, 99340, 99340, 99370, 99360, 99380, 99380, 99410, 
    99430, 99470, 99500, 99520, 99540, 99550, 99560, 99580, 99600, 99620, 
    99680, 99720, 99760, 99800, 99830, 99840, 99830, 99860, 99870, 99890, 
    99930, 99900, 99920, 99870, 99860, 99860, 99830, 99790, 99720, 99630, 
    99560, 99440, 99270, 99170, 99070, 98970, 98870, 98750, 98660, 98660, 
    98640, 98670, 98750, 98830, 98920, 98980, 99040, 99090, 99110, 99100, 
    99080, 99070, 99080, 99080, 99070, 99090, 99130, 99150, 99150, 99220, 
    99260, 99300, 99340, 99340, 99380, 99390, 99410, 99430, 99440, 99510, 
    99520, 99530, 99520, 99590, 99600, 99660, 99660, 99670, 99680, 99680, 
    99730, 99730, 99730, 99800, 99780, 99770, 99800, 99800, 99800, 99770, 
    99820, 99820, 99790, 99740, 99730, 99710, 99740, 99750, 99770, 99770, 
    99770, 99770, 99720, 99730, 99720, 99690, 99690, 99690, 99670, 99670, 
    99690, 99670, 99650, 99600, 99610, 99580, 99550, 99530, 99500, 99480, 
    99450, 99430, 99400, 99350, 99300, 99270, 99230, 99190, 99140, 99100, 
    99050, 99000, 98970, 98890, 98860, 98820, 98770, 98730, 98690, 98650, 
    98610, 98530, 98460, 98430, 98410, 98380, 98410, 98360, 98340, 98310, 
    98280, 98260, 98280, 98270, 98270, 98340, 98340, 98360, 98380, 98390, 
    98440, 98470, 98520, 98560, 98620, 98670, 98720, 98740, 98780, 98820, 
    98810, 98840, 98840, 98880, 98890, 98950, 98940, 98950, 98960, 98970, 
    99030, 99070, 99100, 99120, 99130, 99130, 99110, 99120, 99120, 99120, 
    99090, 99070, 99070, 99060, 99070, 99040, 99000, 98970, 98930, 98890, _, 
    98810, 98770, 98780, 98850, 98780, 98870, 98860, 98880, 98890, 98860, 
    98890, 98900, 98920, 98940, 98920, 98920, 98940, 98980, 99010, _, 99060, 
    99070, 99080, 99080, 99080, 99120, 99140, 99170, _, 99180, 99180, 99160, 
    99150, 99170, 99210, 99250, 99300, 99350, 99420, 99440, 99480, 99500, 
    99490, 99490, 99480, 99470, 99450, 99480, 99500, 99520, 99560, 99620, 
    99660, 99700, 99760, 99770, 99780, 99830, 99860, 99890, 99900, 99930, 
    99960, 100010, 100020, 100050, 100070, 100100, 100120, 100120, 100130, 
    100130, 100140, 100130, 100140, 100150, 100150, 100130, 100100, 100080, 
    100030, 99970, 99930, 99890, 99850, 99790, 99720, 99650, 99580, 99510, 
    99440, 99380, 99330, 99280, 99200, 99120, 99050, 98980, 98900, 98850, 
    98790, 98720, 98650, 98610, 98550, 98500, 98480, 98420, 98390, 98350, 
    98320, 98320, 98300, 98250, 98220, 98180, 98170, 98130, 98130, 98110, 
    98060, 98060, 98030, 98000, 97980, 98000, 97990, 98020, 98000, 98000, 
    97990, 97950, 97970, 97960, 97940, 97950, 97940, 97930, 97910, 97890, 
    97860, 97840, 97800, 97760, 97720, 97700, 97650, 97550, 97460, 97410, 
    97390, 97400, 97470, 97520, 97540, 97540, 97600, 97700, 97790, 97790, 
    97860, 97870, 97910, 97940, 97970, 98010, 98050, 98090, 98100, 98160, 
    98210, 98230, 98260, 98290, 98270, 98280, 98300, 98290, 98350, 98380, 
    98430, 98490, 98560, 98630, 98660, 98710, 98770, 98820, 98870, 98940, 
    98980, 99040, 99080, 99140, 99230, 99310, 99380, 99430, 99510, 99570, 
    99640, 99720, 99790, 99820, 99920, 99990, 100060, 100110, 100210, 100300, 
    100380, 100430, 100510, 100570, 100610, 100660, 100710, 100760, 100790, 
    100870, 100910, 100940, 100980, 100990, 101010, 101000, 100980, 100960, 
    100940, 100930, 100910, 100890, 100870, 100820, 100790, 100750, 100690, 
    100670, 100650, 100610, 100570, 100560, 100550, 100530, 100550, 100550, 
    100550, 100550, 100520, 100520, 100490, 100490, 100450, 100420, 100400, 
    100400, 100390, 100350, 100340, 100300, 100280, 100220, 100150, 100060, 
    99970, 99870, 99780, 99690, 99600, 99480, 99360, 99300, 99200, 99100, 
    99080, 99060, 99070, 99080, 99050, 99060, 99080, 99150, 99190, 99230, 
    99230, 99250, 99260, 99260, 99280, 99280, 99330, 99350, 99380, 99430, 
    99450, 99410, 99470, 99490, 99510, 99540, 99530, 99530, 99580, 99610, 
    99630, 99670, 99700, 99680, 99710, 99750, 99750, 99750, 99760, 99790, 
    99790, 99830, 99880, 99910, 99940, 99940, 99960, 99970, 99990, 99970, 
    99940, 99970, 99990, 99990, 99980, 99990, 99990, 99990, 99970, 99950, 
    99950, 99920, 99910, 99890, 99900, 99930, 99940, 99940, 99940, 99940, 
    99920, 99940, 99940, 99930, 99910, 99900, 99890, 99900, 99900, 99880, 
    99860, 99840, 99830, 99840, 99830, 99820, 99810, 99800, 99800, 99780, 
    99780, 99750, 99750, 99740, 99700, 99710, 99720, 99720, 99740, 99770, 
    99780, 99820, 99880, 99920, 99960, 99960, 100010, 100060, 100130, 100190, 
    100240, 100270, 100310, 100370, 100400, 100400, 100420, 100410, 100470, 
    100500, 100540, 100600, 100650, 100720, 100780, 100840, 100910, 100990, 
    101130, 101150, 101230, 101260, 101360, 101420, 101470, 101530, 101580, 
    101630, 101690, 101740, 101770, 101800, 101830, 101890, 101890, 101910, 
    101920, 101920, 101940, 101950, 101980, 101980, 101990, 101980, 101970, 
    101960, 101920, 101910, 101890, 101850, 101820, 101830, 101810, 101770, 
    101710, 101630, 101600, 101520, 101460, 101410, 101290, 101220, 101100, 
    101030, 100970, 100880, 100790, 100660, 100560, 100450, 100280, 100160, 
    100030, 99930, 99800, 99710, 99570, 99510, 99380, 99200, 99050, 98900, 
    98750, 98600, 98440, 98310, 98190, 98120, 98030, 97880, 97770, 97660, 
    97610, 97500, 97390, 97360, 97340, 97260, 97200, 97060, 96940, 97130, 
    97160, 97240, 97310, 97290, 97250, 97210, 97150, 97200, 97160, 97090, 
    97110, 97060, 97060, 97060, 97120, 97090, 97030, 97010, 96990, 96930, 
    96910, 96950, 96970, 96970, 96950, 96940, 96950, 96950, 96920, 96900, 
    96900, 96840, 96860, 96860, 96830, 96810, 96770, 96770, 96760, 96750, 
    96730, 96710, 96700, 96700, 96720, 96740, 96760, 96770, 96790, 96800, 
    96810, 96840, 96870, 96900, 96930, 96970, 97030, 97090, 97170, 97230, 
    97280, 97350, 97420, 97500, 97570, 97660, 97760, 97880, 98000, 98130, 
    98230, 98330, 98410, 98520, 98590, 98650, 98710, 98720, 98790, 98840, 
    98890, 98950, 98980, 98990, 99000, 99030, 99090, 99080, 99070, 99030, 
    98990, 98980, 98970, 98910, 98890, 98840, 98790, 98740, 98680, 98610, 
    98500, 98420, 98350, 98260, 98240, 98250, 98250, 98220, 98200, 98180, 
    98160, 98110, 98080, 98040, 97980, 97930, 97900, 97890, 97860, 97830, 
    97790, 97760, 97740, 97730, 97680, 97640, 97610, 97580, 97540, 97520, 
    97490, 97450, 97410, 97440, 97440, 97440, 97440, 97450, 97440, 97450, 
    97490, 97520, 97560, 97610, 97610, 97580, 97580, 97600, 97640, 97690, 
    97720, 97730, 97800, 97820, 97900, 97950, 97990, 98050, 98120, 98200, 
    98260, 98290, 98320, 98390, 98440, 98480, 98560, 98600, 98680, 98750, 
    98780, 98800, 98840, 98860, 98920, 98990, 99040, 99110, 99180, 99250, 
    99340, 99400, 99470, 99550, 99630, 99720, 99790, 99860, 99910, 100000, 
    100070, 100150, 100250, 100330, 100420, 100510, 100530, 100590, 100640, 
    100650, 100680, 100680, 100540, 100390, 100350, 100310, 100280, 100270, 
    100300, 100310, 100350, 100390, 100490, 100600, 100730, 100840, 100900, 
    101050, 101140, 101240, 101330, 101350, 101340, 101380, 101400, 101420, 
    101490, 101500, 101490, 101510, 101510, 101460, 101420, 101360, 101300, 
    101240, 101230, 101230, 101150, 101100, 101060, 101010, 100940, 100850, 
    100710, 100620, 100590, 100490, 100410, 100350, 100280, 100240, 100210, 
    100120, 100010, 99900, 99820, 99710, 99580, 99550, 99570, 99580, 99610, 
    99640, 99770, 99860, 99960, 100020, 100100, 100110, 100150, 100150, 
    100110, 100150, 100130, 100140, 100130, 100120, 100010, 99920, 99810, 
    99690, 99530, 99490, 99330, 99350, 99360, 99440, 99470, 99510, 99540, 
    99560, 99570, 99660, 99760, 99880, 99990, 100100, 100220, 100340, 100450, 
    100550, 100630, 100680, 100760, 100710, 100710, 100710, 100710, 100700, 
    100680, 100600, 100550, 100490, 100380, 100260, 100190, 100150, 100200, 
    100180, 100210, 100300, 100330, 100440, 100540, 100570, 100600, 100630, 
    100590, 100540, 100480, 100490, 100400, 100260, 100220, 100200, 100200, 
    100230, 100380, 100540, 100720, 100910, 101070, 101260, 101430, 101580, 
    101760, 101930, 102010, 102000, 101960, 101890, 101880, 101760, 101670, 
    101610, 101560, 101450, 101400, 101330, 101270, 101190, 101120, 101100, 
    101030, 101070, 101170, 101160, 101210, 101220, 101240, 101280, 101310, 
    101280, 101310, 101300, 101280, 101270, 101290, 101320, 101340, 101370, 
    101400, 101390, 101400, 101430, 101480, 101470, 101500, 101550, 101570, 
    101600, 101650, 101690, 101750, 101790, 101830, 101870, 101920, 101960, 
    101980, 102010, 102030, 102070, 102080, 102110, 102130, 102130, 102130, 
    102100, 102100, 102110, 102110, 102090, 102070, 102060, 102050, 102030, 
    102020, 102000, 101960, 101950, 101920, 101900, 101900, 101860, 101810, 
    101800, 101800, 101820, 101810, 101800, 101790, 101780, 101770, 101770, 
    101790, 101810, 101820, 101850, 101870, 101900, 101920, 101930, 101950, 
    101960, 101980, 102000, 102010, 102020, 102030, 102070, 102090, 102130, 
    102160, 102180, 102190, 102180, 102200, 102200, 102190, 102200, 102190, 
    102190, 102200, 102200, 102150, 102120, 102100, 102060, 102050, 102010, 
    101970, 101930, 101870, 101840, 101820, 101820, 101830, 101810, 101800, 
    101800, 101800, 101810, 101810, 101820, 101820, 101840, 101870, 101890, 
    101910, 101920, 101940, 101940, 101960, 101970, 101990, 102000, 102020, 
    102020, 102030, 102050, 102050, 102040, 102040, 102050, 102050, 102030, 
    102040, 102030, 102030, 102030, 102030, 102050, 102060, 102060, 102050, 
    102050, 102070, 102070, 102060, 102040, 102030, 102050, 102080, 102110, 
    102140, 102140, 102130, 102150, 102140, 102130, 102120, 102150, 102160, 
    102180, 102200, 102250, 102290, 102310, 102340, 102350, 102350, 102380, 
    102400, 102420, 102450, 102490, 102550, 102610, 102650, 102690, 102730, 
    102780, 102820, 102850, 102880, 102910, 102950, 102990, 103030, 103090, 
    103110, 103130, 103160, 103160, 103190, 103210, 103240, 103240, 103230, 
    103240, 103260, 103280, 103270, 103280, 103260, 103240, 103230, 103200, 
    103160, 103110, 103100, 103030, 102990, 102950, 102890, 102840, 102770, 
    102690, 102620, 102550, 102470, 102410, 102330, 102260, 102230, 102200, 
    102190, 102150, 102110, 102060, 102020, 101960, 101920, 101890, 101850, 
    101790, 101730, 101680, 101630, 101550, 101460, 101410, 101320, 101250, 
    101150, 101040, 100920, 100840, 100800, 100780, 100810, 100800, 100760, 
    100720, 100730, 100740, 100760, 100780, 100810, 100820, 100860, 100900, 
    100940, 101010, 101030, 101060, 101080, 101120, 101170, 101170, 101190, 
    101220, 101230, 101270, 101310, 101340, 101350, 101330, 101330, 101360, 
    101380, 101370, 101370, 101390, 101370, 101390, 101390, 101400, 101410, 
    101400, 101400, 101390, 101390, 101390, 101380, 101380, 101400, 101460, 
    101520, 101530, 101530, 101570, 101600, 101580, 101610, 101590, 101590, 
    101600, 101600, 101640, 101680, 101730, 101770, 101790, 101780, 101780, 
    101780, 101800, 101790, 101790, 101740, 101740, 101750, 101730, 101740, 
    101690, 101660, 101630, 101590, 101570, 101530, 101480, 101460, 101440, 
    101400, 101340, 101290, 101220, 101190, 101130, 101080, 101050, 101040, 
    101040, 101000, 100990, 100990, 101000, 100980, 101020, 101030, 101040, 
    101050, 101050, 101070, 101050, 101040, 101050, 101050, 101050, 101040, 
    101040, 101020, 101010, 101010, 100980, 100960, 100970, 100950, 100940, 
    100940, 100930, 100920, 100890, 100890, 100860, 100840, 100820, 100790, 
    100780, 100750, 100740, 100720, 100670, 100650, 100630, 100610, 100580, 
    100550, 100520, 100520, 100510, 100490, 100490, 100520, 100520, 100500, 
    100470, 100450, 100460, 100500, 100520, 100520, 100520, 100560, 100590, 
    100590, 100610, 100620, 100630, 100630, 100640, 100630, 100600, 100570, 
    100570, 100560, 100550, 100540, 100480, 100420, 100320, 100300, 100280, 
    100250, 100170, 100140, 100100, 100060, 100030, 100000, 99950, 99900, 
    99890, 99840, 99840, 99830, 99810, 99800, 99810, 99820, 99880, 99910, 
    99920, 99940, 99950, 99970, 99990, 99990, 99970, 99960, 99950, 99970, 
    99980, 99960, 99970, 99990, 100000, 100030, 100060, 100120, 100140, 
    100180, 100240, 100260, 100350, 100430, 100470, 100520, 100550, 100560, 
    100610, 100630, 100680, 100720, 100720, 100770, 100750, 100810, 100810, 
    100810, 100820, 100830, 100820, 100840, 100790, 100760, 100740, 100730, 
    100730, 100730, 100720, 100730, 100750, 100730, 100720, 100730, 100740, 
    100730, 100720, 100740, 100780, 100770, 100790, 100820, 100830, 100860, 
    100870, 100860, 100850, 100840, 100850, 100860, 100910, 100960, 101010, 
    101020, 101040, 101060, 101100, 101130, 101140, 101170, 101140, 101140, 
    101150, 101140, 101110, 101060, 100990, 100930, 100870, 100780, 100730, 
    100660, 100570, 100500, 100480, 100410, 100350, 100310, 100280, 100220, 
    100150, 100080, 100000, 99930, 99850, 99820, 99750, 99700, 99630, 99560, 
    99490, 99420, 99370, 99310, 99240, 99190, 99130, 99070, 99040, 99030, 
    98990, 98950, 98930, 98900, 98830, 98800, 98770, 98740, 98690, 98660, 
    98660, 98630, 98610, 98600, 98570, 98560, 98520, 98490, 98450, 98400, 
    98380, 98350, 98400, 98350, 98310, 98260, 98220, 98200, 98190, 98200, 
    98160, 98170, 98150, 98110, 98090, 98060, 98010, 97970, 97930, 97880, 
    97840, 97800, 97790, 97780, 97770, 97790, 97810, 97830, 97830, 97830, 
    97850, 97820, 97790, 97800, 97820, 97810, 97810, 97830, 97850, 97840, 
    97830, 97860, 97830, 97840, 97830, 97870, 97920, 97970, 97970, 98010, 
    98090, 98160, 98260, 98300, 98350, 98400, 98420, 98480, 98530, 98620, 
    98630, 98670, 98710, 98740, 98750, 98790, 98830, 98830, 98840, 98880, 
    98860, 98830, 98840, 98850, 98900, 98930, 98910, 98920, 98890, 98850, 
    98830, 98850, 98870, 98880, 98870, 98900, 98900, 98920, 98910, 98960, 
    98890, 98970, 99000, 99000, 99010, 99060, 99070, 99100, 99120, 99160, 
    99130, 99190, 99180, 99180, 99170, 99170, 99140, 99170, 99180, 99180, 
    99240, 99290, 99270, 99320, 99360, 99330, 99320, 99340, 99420, 99390, 
    99390, 99420, 99350, 99380, 99430, 99510, 99540, 99590, 99620, 99700, 
    99750, 99730, 99750, 99780, 99840, 99870, 99880, 99910, 99950, 99980, 
    99980, 100000, 100070, 100090, 100090, 100130, 100180, 100220, 100250, 
    100240, 100320, 100380, 100410, 100410, 100400, 100420, 100430, 100460, 
    100560, 100560, 100580, 100680, 100770, 100830, 100840, 100900, 100960, 
    101020, 101030, 101040, 101090, 101080, 101130, 101140, 101190, 101220, 
    101240, 101270, 101300, 101280, 101250, 101230, 101220, 101230, 101220, 
    101180, 101140, 101120, 101090, 101050, 101010, 100950, 100890, 100860, 
    100850, 100840, 100810, 100770, 100730, 100690, 100650, 100630, 100600, 
    100550, 100510, 100510, 100490, 100470, 100450, 100450, 100410, 100400, 
    100400, 100400, 100390, 100370, 100360, 100350, 100380, 100380, 100400, 
    100410, 100400, 100370, 100390, 100370, 100360, 100350, 100360, 100360, 
    100390, 100380, 100360, 100360, 100340, 100320, 100320, 100320, 100310, 
    100300, 100300, 100320, 100330, 100310, 100290, 100280, 100260, 100250, 
    100220, 100200, 100180, 100160, 100170, 100140, 100150, 100130, 100100, 
    100060, 100030, 99990, 99960, 99940, 99900, 99880, 99840, 99830, 99820, 
    99800, 99780, 99740, 99680, 99640, 99610, 99600, 99570, 99520, 99490, 
    99460, 99430, 99390, 99290, 99190, 99130, 99060, 98970, 98910, 98830, 
    98750, 98770, 98640, 98650, 98640, 98650, 98570, 98560, 98500, 98460, 
    98430, 98400, 98400, 98370, 98390, 98390, 98390, 98400, 98450, 98470, 
    98460, 98490, 98540, 98540, 98570, 98580, 98590, 98620, 98640, 98700, 
    98710, 98720, 98720, 98750, 98770, 98790, 98790, 98800, 98820, 98840, 
    98860, 98880, 98890, 98900, 98940, 98970, 98990, 99000, 99000, 99020, 
    99050, 99100, 99130, 99150, 99170, 99190, 99210, 99220, 99240, 99260, 
    99280, 99300, 99320, 99350, 99370, 99410, 99420, 99490, 99540, 99580, 
    99630, 99660, 99700, 99770, 99850, 99920, 100000, 100060, 100110, 100170, 
    100210, 100250, 100290, 100310, 100330, 100340, 100350, 100360, 100400, 
    100410, 100420, 100420, 100420, 100430, 100450, 100450, 100450, 100460, 
    100450, 100510, 100530, 100540, 100550, 100560, 100560, 100560, 100550, 
    100500, 100460, 100410, 100370, 100340, 100300, 100300, 100320, 100330, 
    100340, 100350, 100410, 100420, 100450, 100480, 100530, 100600, 100650, 
    100700, 100720, 100720, 100740, 100770, 100770, 100780, 100770, 100770, 
    100780, 100800, 100840, 100770, 100780, 100710, 100640, 100570, 100570, 
    100540, 100500, 100470, 100450, 100430, 100430, 100450, 100480, 100510, 
    100530, 100560, 100580, 100610, 100610, 100610, 100640, 100660, 100650, 
    100620, 100600, 100580, 100560, 100550, 100530, 100520, 100490, 100480, 
    100480, 100490, 100500, 100500, 100520, 100540, 100550, 100540, 100550, 
    100560, 100570, 100570, 100600, 100630, 100620, 100650, 100670, 100660, 
    100660, 100640, 100600, 100540, 100510, 100470, 100440, 100410, 100350, 
    100320, 100310, 100240, 100160, 100110, 100100, 100050, 99990, 99950, 
    99930, 99920, 99930, 99950, 99950, 99960, 99960, 100010, 100020, 100040, 
    100060, 100090, 100140, 100190, 100220, 100250, 100280, 100280, 100260, 
    100230, 100180, 100150, 100100, 100040, 100040, 100040, 100020, 99970, 
    99910, 99830, 99750, 99690, 99610, 99530, 99450, 99430, 99400, 99390, 
    99350, 99310, 99270, 99230, 99150, 99110, 99060, 99060, 99010, 98970, 
    98940, 98930, 98930, 98900, 98870, 98860, 98850, 98830, 98810, 98800, 
    98760, 98790, 98840, 98860, 98910, 98960, 99020, 99030, 99050, 99090, 
    99130, 99190, 99240, 99290, 99350, 99410, 99500, 99560, 99620, 99670, 
    99710, 99750, 99810, 99840, 99890, 99900, 99920, 99960, 99980, 99990, 
    100010, 100030, 100000, 100000, 99980, 99960, 99910, 99870, 99860, 99800, 
    99760, 99750, 99710, 99700, 99650, 99590, 99530, 99550, 99560, 99580, 
    99580, 99560, 99600, 99620, 99670, 99700, 99700, 99720, 99800, 99840, 
    99890, 99950, 100020, 100060, 100110, 100170, 100220, 100250, 100300, 
    100340, 100390, 100430, 100460, 100480, 100500, 100540, 100590, 100580, 
    100580, 100580, 100520, 100520, 100540, 100600, 100610, 100650, 100690, 
    100710, 100760, 100810, 100860, 100920, 100990, 101060, 101110, 101160, 
    101200, 101220, 101260, 101310, 101360, 101400, 101410, 101390, 101420, 
    101450, 101470, 101470, 101450, 101450, 101580, 101450, 101460, 101460, 
    101450, 101450, 101430, 101410, 101420, 101390, 101350, 101340, 101370, 
    101360, 101340, 101350, 101330, 101300, 101270, 101270, 101250, 101250, 
    101270, 101270, 101270, 101290, 101300, 101280, 101270, 101270, 101250, 
    101260, 101270, 101260, 101270, 101280, 101320, 101300, 101310, 101350, 
    101370, 101380, 101360, 101330, 101340, 101350, 101340, 101350, 101370, 
    101370, 101350, 101320, 101300, 101270, 101220, 101180, 101160, 101150, 
    101110, 101080, 101050, 101050, 101040, 101000, 100960, 100930, 100910, 
    100890, 100870, 100830, 100780, 100760, 100750, 100710, 100700, 100680, 
    100650, 100630, 100610, 100600, 100590, 100580, 100570, 100570, 100560, 
    100570, 100580, 100580, 100570, 100570, 100550, 100540, 100530, 100530, 
    100510, 100510, 100500, 100500, 100500, 100500, 100460, 100450, 100420, 
    100400, 100390, 100370, 100340, 100330, 100310, 100320, 100310, 100320, 
    100310, 100320, 100320, 100310, 100300, 100300, 100280, 100260, 100240, 
    100190, 100160, 100140, 100100, 100090, 100050, 100020, 100020, 99980, 
    99980, 99960, 99940, 99940, 99960, 99990, 99990, 100020, 100030, 100030, 
    100020, 100030, 100050, 100020, 99990, 99950, 99910, 99860, 99810, 99740, 
    99660, 99560, 99450, 99370, 99340, 99260, 99240, 99220, 99240, 99300, 
    99350, 99390, 99370, 99360, 99400, 99390, 99420, 99450, 99470, 99510, 
    99530, 99590, 99650, 99690, 99720, 99730, 99730, 99730, 99730, 99740, 
    99730, 99760, 99790, 99820, 99840, 99870, 99860, 99860, 99860, 99870, 
    99870, 99880, 99900, 99940, 99950, 99970, 100000, 100000, 99990, 100030, 
    100040, 100050, 100070, 100100, 100110, 100100, 100140, 100160, 100160, 
    100180, 100160, 100140, 100140, 100130, 100140, 100110, 100080, 100080, 
    100080, 100090, 100090, 100080, 100060, 100040, 100020, 100010, 100010, 
    99980, 100000, 99950, 99960, 99950, 99950, 99950, 99980, 100040, 100080, 
    100100, 100150, 100190, 100250, 100290, 100330, 100360, 100350, 100360, 
    100380, 100370, 100390, 100390, 100410, 100430, 100440, 100470, 100480, 
    100530, 100530, 100550, 100580, 100590, 100620, 100650, 100670, 100700, 
    100730, 100770, 100810, 100840, 100880, 100900, 100910, 100910, 100920, 
    100910, 100940, 100940, 100940, 100960, 100970, 101010, 101000, 100970, 
    100970, 100970, 100950, 100950, 100950, 100950, 100960, 100950, 100950, 
    100970, 100970, 100970, 100970, 100990, 101010, 101030, 101050, 101080, 
    101100, 101120, 101150, 101180, 101200, 101210, 101220, 101230, 101270, 
    101270, 101310, 101330, 101350, 101380, 101400, 101420, 101450, 101460, 
    101440, 101440, 101440, 101440, 101430, 101430, 101420, 101440, 101450, 
    101440, 101450, 101420, 101400, 101390, 101370, 101380, 101380, 101380, 
    101350, 101330, 101300, 101280, 101270, 101270, 101270, 101280, 101270, 
    101270, 101250, 101280, 101260, 101270, 101280, 101300, 101320, 101340, 
    101330, 101330, 101340, 101320, 101300, 101310, 101300, 101270, 101240, 
    101210, 101180, 101160, 101180, 101170, 101130, 101100, 101050, 101020, 
    101010, 100980, 100950, 100910, 100930, 100860, 100810, 100730, 100620, 
    100560, 100480, 100380, 100280, 100240, 100190, 100170, 100150, 100220, 
    100250, 100280, 100300, 100350, 100380, 100410, 100380, 100370, 100390, 
    100390, 100390, 100400, 100370, 100400, 100370, 100370, 100330, 100340, 
    100340, 100310, 100250, 100230, 100180, 100130, 100080, 100020, 99910, 
    99770, 99590, 99410, 99260, 99120, 99040, 99090, 99100, 99110, 99130, 
    99100, 99050, 99050, 99040, 98980, 98940, 98990, 99020, 99210, 99440, 
    99600, 99820, 99990, 100180, 100310, 100450, 100550, 100590, 100600, 
    100610, 100570, 100530, 100360, 100210, 100050, 99800, 99520, 99250, 
    98920, 98620, 98380, 98140, 97980, 97850, 97770, 97750, 97780, 97840, 
    97930, 98050, 98170, 98340, 98520, 98720, 98940, 99130, 99320, 99470, 
    99590, 99720, 99810, 99930, 100070, 100140, 100260, 100340, 100420, 
    100450, 100490, 100480, 100510, 100520, 100540, 100590, 100610, 100660, 
    100660, 100720, 100750, 100750, 100740, 100760, 100760, 100790, 100830, 
    100860, 100890, 100920, 101020, 101090, 101140, 101200, 101230, 101290, 
    101350, 101370, 101390, 101420, 101440, 101480, 101500, 101540, 101600, 
    101630, 101650, 101650, 101670, 101680, 101670, 101680, 101660, 101680, 
    101700, 101700, 101720, 101740, 101730, 101720, 101690, 101680, 101650, 
    101650, 101600, 101570, 101560, 101570, 101530, 101600, 101560, 101550, 
    101520, 101490, 101460, 101380, 101390, 101380, 101380, 101360, 101350, 
    101350, 101320, 101280, 101260, 101230, 101200, 101160, 101140, 101120, 
    101100, 101080, 101080, 101070, 101050, 101020, 101020, 101050, 101030, 
    101030, 101000, 100980, 100990, 101000, 101010, 101000, 101000, 101000, 
    100990, 101000, 101030, 100990, 100990, 101010, 101050, 101070, 101090, 
    101100, 101100, 101090, 101100, 101080, 101090, 101070, 101070, 101050, 
    101040, 101020, 101020, 101020, 101000, 100950, 100910, 100900, 100880, 
    100850, 100840, 100810, 100790, 100800, 100780, 100770, 100750, 100720, 
    100690, 100670, 100670, 100640, 100620, 100620, 100600, 100580, 100590, 
    100570, 100560, 100550, 100530, 100520, 100510, 100500, 100500, 100500, 
    100510, 100510, 100520, 100550, 100550, 100570, 100600, 100600, 100640, 
    100630, 100670, 100690, 100700, 100730, 100760, 100770, 100790, 100810, 
    100800, 100810, 100830, 100830, 100840, 100840, 100870, 100880, 100910, 
    100920, 100930, 100960, 100970, 100990, 100970, 100960, 100960, 100930, 
    100910, 100890, 100870, 100880, 100860, 100840, 100800, 100790, 100770, 
    100740, 100730, 100720, 100720, 100720, 100720, 100710, 100710, 100680, 
    100670, 100670, 100670, 100660, 100650, 100650, 100650, 100650, 100620, 
    100610, 100600, 100580, 100590, 100570, 100550, 100530, 100530, 100500, 
    100470, 100450, 100450, 100430, 100410, 100410, 100410, 100390, 100400, 
    100390, 100380, 100390, 100410, 100430, 100430, 100420, 100420, 100420, 
    100420, 100410, 100400, 100380, 100370, 100350, 100330, 100320, 100300, 
    100290, 100250, 100220, 100190, 100150, 100100, 100050, 100040, 100010, 
    99950, 99910, 99850, 99820, 99740, 99660, 99620, 99580, 99510, 99450, 
    99370, 99320, 99250, 99200, 99140, 99090, 98970, 98860, 98790, 98620, 
    98500, 98380, 98290, 98210, 98140, 98050, 98000, 97940, 97860, 97800, 
    97710, 97630, 97560, 97530, 97470, 97410, 97370, 97320, 97260, 97210, 
    97180, 97190, 97190, 97180, 97220, 97250, 97290, 97360, 97450, 97550, 
    97660, 97770, 97890, 98000, 98100, 98190, 98250, 98290, 98360, 98430, 
    98520, 98610, 98660, 98710, 98750, 98790, 98830, 98850, 98860, 98890, 
    98910, 98920, 98960, 98950, 98980, 98970, 98980, 98990, 99010, 99030, 
    99030, 99040, 99070, 99120, 99110, 99160, 99170, 99180, 99190, 99210, 
    99210, 99210, 99220, 99200, 99200, 99220, 99220, 99210, 99240, 99270, 
    99270, 99300, 99320, 99330, 99380, 99400, 99450, 99500, 99530, 99570, 
    99620, 99680, 99740, 99770, 99840, 99880, 99960, 99990, 100020, 100070, 
    100120, 100180, 100250, 100300, 100380, 100440, 100490, 100520, 100550, 
    100600, 100650, 100690, 100740, 100800, 100850, 100890, 100930, 100950, 
    101010, 101030, 101050, 101110, 101150, 101190, 101210, 101270, 101290, 
    101290, 101310, 101350, 101350, 101380, 101390, 101400, 101400, 101420, 
    101440, 101450, 101470, 101490, 101500, 101520, 101510, 101520, 101540, 
    101550, 101560, 101560, 101560, 101580, 101590, 101590, 101570, 101570, 
    101560, 101560, 101570, 101570, 101580, 101600, 101620, 101620, 101640, 
    101640, 101630, 101610, 101600, 101570, 101570, 101580, 101580, 101610, 
    101610, 101620, 101640, 101650, 101650, 101630, 101630, 101620, 101600, 
    101610, 101610, 101610, 101640, 101670, 101700, 101690, 101710, 101720, 
    101720, 101730, 101730, 101740, 101740, 101760, 101780, 101780, 101780, 
    101770, 101740, 101720, 101710, 101700, 101680, 101680, 101680, 101680, 
    101670, 101670, 101670, 101660, 101640, 101630, 101600, 101570, 101540, 
    101530, 101520, 101520, 101510, 101510, 101510, 101490, 101460, 101430, 
    101390, 101390, 101380, 101380, 101370, 101370, 101380, 101390, 101390, 
    101380, 101370, 101340, 101340, 101340, 101340, 101340, 101340, 101330, 
    101320, 101340, 101350, 101360, 101380, 101400, 101410, 101430, 101450, 
    101490, 101510, 101530, 101550, 101560, 101580, 101590, 101600, 101600, 
    101590, 101580, 101580, 101600, 101600, 101600, 101610, 101610, 101620, 
    101620, 101600, 101570, 101580, 101580, 101580, 101570, 101570, 101570, 
    101560, 101570, 101560, 101530, 101520, 101500, 101480, 101480, 101480, 
    101460, 101460, 101440, 101420, 101430, 101410, 101400, 101350, 101310, 
    101290, 101250, 101230, 101200, 101190, 101160, 101120, 101100, 101090, 
    101080, 101060, 101060, 101050, 101080, 101110, 101130, 101170, 101220, 
    101260, 101280, 101270, 101290, 101350, 101350, 101390, 101410, 101440, 
    101460, 101510, 101520, 101530, 101570, 101580, 101560, 101590, 101630, 
    101630, 101670, 101650, 101670, 101670, 101700, 101720, 101740, 101740, 
    101750, 101780, 101790, 101810, 101820, 101840, 101790, 101810, 101830, 
    101870, 101880, 101850, 101880, 101880, 101890, 101880, 101860, 101850, 
    101860, 101860, 101880, 101930, 101920, 101970, 101960, 102000, 102040, 
    102050, 102070, 102060, 102050, 102060, 102040, 102050, 102070, 102080, 
    102070, 102060, 102080, 102060, 102040, 102010, 101990, 101970, 101950, 
    101960, 101940, 101900, 101870, 101830, 101790, 101730, 101720, 101630, 
    101590, 101540, 101470, 101420, 101370, 101290, 101260, 101230, 101160, 
    101120, 101090, 101080, 101050, 101040, 101020, 101010, 101010, 101000, 
    100990, 100990, 100980, 100990, 100980, 100960, 100950, 100930, 100900, 
    100980, 100980, 101000, 101000, 101060, 101060, 101050, 101080, 101090, 
    101110, 101100, 101100, 101140, 101130, 101150, 101200, 101180, 101190, 
    101210, 101180, 101200, 101200, 101220, 101200, 101230, 101250, 101270, 
    101260, 101290, 101310, 101300, 101310, 101290, 101290, 101290, 101300, 
    101320, 101330, 101330, 101330, 101330, 101330, 101340, 101360, 101340, 
    101350, 101350, 101370, 101380, 101390, 101400, 101410, 101410, 101410, 
    101420, 101400, 101410, 101430, 101440, 101450, 101470, 101470, 101460, 
    101430, 101430, 101430, 101420, 101390, 101370, 101350, 101330, 101320, 
    101320, 101270, 101280, 101250, 101220, 101210, 101180, 101170, 101140, 
    101120, 101090, 101070, 101050, 101020, 101030, 101020, 101000, 100970, 
    100950, 100930, 100920, 100880, 100870, 100860, 100840, 100810, 100780, 
    100760, 100740, 100720, 100690, 100670, 100650, 100640, 100650, 100620, 
    100630, 100640, 100660, 100670, 100680, 100700, 100720, 100730, 100740, 
    100760, 100770, 100770, 100800, 100810, 100840, 100880, 100900, 100920, 
    100920, 100930, 100940, 100960, 100960, 100970, 100970, 100980, 100980, 
    101000, 101000, 101000, 101010, 100990, 100990, 101000, 101000, 101000, 
    101000, 101020, 101030, 101050, 101080, 101090, 101090, 101100, 101110, 
    101110, 101120, 101130, 101140, 101160, 101190, 101210, 101220, 101240, 
    101260, 101270, 101280, 101310, 101330, 101360, 101400, 101410, 101440, 
    101450, 101460, 101490, 101510, 101500, 101500, 101490, 101490, 101480, 
    101460, 101460, 101440, 101410, 101390, 101360, 101340, 101320, 101310, 
    101290, 101290, 101280, 101290, 101280, 101280, 101270, 101240, 101250, 
    101240, 101230, 101210, 101180, 101190, 101200, 101200, 101200, 101190, 
    101200, 101190, 101190, 101170, 101160, 101130, 101120, 101120, 101120, 
    101110, 101110, 101090, 101070, 101060, 101030, 101030, 101020, 101020, 
    101040, 101040, 101060, 101090, 101130, 101140, 101170, 101190, 101200, 
    101220, 101260, 101310, 101330, 101380, 101440, 101500, 101540, 101580, 
    101640, 101690, 101730, 101780, 101820, 101840, 101880, 101910, 101960, 
    102010, 102040, 102080, 102120, 102150, 102180, 102190, 102210, 102220, 
    102250, 102290, 102320, 102350, 102400, 102450, 102500, 102550, 102590, 
    102610, 102640, 102690, 102720, 102760, 102820, 102880, 102930, 102970, 
    103020, 103060, 103090, 103130, 103170, 103210, 103250, 103300, 103350, 
    103400, 103430, 103450, 103470, 103460, 103480, 103440, 103440, 103480, 
    103470, 103470, 103460, 103460, 103440, 103460, 103410, 103420, 103440, 
    103390, 103350, 103330, 103330, 103330, 103360, 103370, 103360, 103360, 
    103340, 103360, 103340, 103310, 103300, 103270, 103270, 103240, 103230, 
    103220, 103230, 103220, 103180, 103150, 103120, 103070, 103020, 102980, 
    102960, 102950, 102940, 102920, 102890, 102870, 102880, 102890, 102870, 
    102880, 102880, 102900, 102930, 102980, 103030, 103060, 103110, 103170, 
    103210, 103230, 103260, 103290, 103320, 103340, 103380, 103410, 103430, 
    103450, 103470, 103480, 103510, 103530, 103540, 103530, 103490, 103480, 
    103450, 103430, 103410, 103410, 103380, 103370, 103350, 103340, 103310, 
    103290, 103270, 103240, 103230, 103200, 103170, 103150, 103130, 103080, 
    103040, 102990, 102970, 102920, 102860, 102800, 102720, 102670, 102640, 
    102600, 102540, 102490, 102460, 102400, 102350, 102310, 102270, 102210, 
    102140, 102090, 102050, 102000, 102000, 102000, 101970, 101970, 101940, 
    101910, 101900, 101880, 101860, 101850, 101830, 101820, 101820, 101810, 
    101820, 101840, 101850, 101840, 101830, 101800, 101780, 101790, 101800, 
    101800, 101830, 101850, 101850, 101860, 101840, 101850, 101850, 101840, 
    101830, 101810, 101820, 101830, 101840, 101870, 101880, 101900, 101900, 
    101900, 101890, 101910, 101930, 101950, 101990, 102030, 102080, 102100, 
    102120, 102150, 102180, 102200, 102210, 102210, 102220, 102250, 102270, 
    102290, 102320, 102330, 102350, 102340, 102340, 102340, 102350, 102340, 
    102310, 102310, 102330, 102340, 102330, 102310, 102300, 102290, 102280, 
    102240, 102200, 102160, 102160, 102120, 102090, 102080, 102060, 102050, 
    102020, 102000, 101990, 101970, 101950, 101930, 101920, 101950, 101970, 
    102010, 102030, 102050, 102060, 102080, 102090, 102110, 102110, 102140, 
    102150, 102150, 102160, 102150, 102160, 102170, 102150, 102130, 102120, 
    102080, 102050, 102020, 102000, 102000, 101990, 101990, 102010, 101980, 
    101980, 101970, 101950, 101940, 101920, 101890, 101860, 101840, 101810, 
    101780, 101780, 101780, 101760, 101750, 101720, 101700, 101680, 101680, 
    101670, 101650, 101660, 101650, 101640, 101630, 101620, 101630, 101620, 
    101580, 101540, 101520, 101490, 101480, 101470, 101440, 101430, 101410, 
    101370, 101340, 101320, 101310, 101300, 101280, 101280, 101280, 101270, 
    101300, 101310, 101340, 101350, 101370, 101400, 101410, 101420, 101420, 
    101440, 101490, 101490, 101520, 101560, 101590, 101620, 101660, 101680, 
    101700, 101710, 101720, 101740, 101770, 101790, 101810, 101820, 101840, 
    101840, 101850, 101860, 101850, 101860, 101840, 101820, 101820, 101790, 
    101790, 101800, 101790, 101790, 101770, 101770, 101760, 101750, 101730, 
    101750, 101750, 101760, 101760, 101770, 101770, 101760, 101770, 101770, 
    101760, 101730, 101710, 101670, 101690, 101680, 101670, 101610, 101580, 
    101590, 101580, 101570, 101570, 101530, 101490, 101440, 101400, 101380, 
    101330, 101320, 101290, 101220, 101130, 101100, 101040, 101000, 101000, 
    100970, 100950, 100940, 100910, 100910, 100890, 100800, 100720, 100680, 
    100600, 100550, 100530, 100460, 100470, 100460, 100480, 100500, 100540, 
    100580, 100630, 100700, 100770, 100810, 100860, 100920, 100970, 100990, 
    101040, 101080, 101110, 101150, 101210, 101230, 101260, 101280, 101280, 
    101290, 101320, 101340, 101350, 101360, 101390, 101400, 101400, 101410, 
    101420, 101400, 101390, 101390, 101360, 101340, 101310, 101310, 101290, 
    101290, 101260, 101250, 101210, 101180, 101110, 101080, 101010, 100960, 
    100900, 100880, 100860, 100810, 100750, 100690, 100640, 100590, 100530, 
    100440, 100400, 100340, 100260, 100190, 100120, 100070, 100020, 99980, 
    99930, 99890, 99860, 99860, 99840, 99820, 99800, 99780, 99780, 99780, 
    99790, 99780, 99770, 99760, 99760, 99750, 99760, 99770, 99780, 99780, 
    99790, 99800, 99800, 99810, 99800, 99790, 99790, 99800, 99800, 99820, 
    99850, 99860, 99890, 99910, 99920, 99910, 99920, 99910, 99910, 99910, 
    99900, 99910, 99910, 99920, 99920, 99910, 99900, 99890, 99870, 99840, 
    99810, 99800, 99820, 99820, 99840, 99860, 99870, 99880, 99860, 99830, 
    99800, 99800, 99750, 99740, 99730, 99710, 99700, 99670, 99640, 99620, 
    99610, 99600, 99570, 99520, 99490, 99400, 99420, 99470, 99480, 99500, 
    99550, 99550, 99580, 99590, 99580, 99570, 99570, 99570, 99570, 99560, 
    99560, 99580, 99570, 99550, 99570, 99570, 99560, 99570, 99600, 99650, 
    99700, 99710, 99740, 99780, 99830, 99860, 99900, 99940, 99970, 100000, 
    100030, 100060, 100100, 100140, 100160, 100200, 100250, 100280, 100300, 
    100320, 100350, 100370, 100390, 100420, 100440, 100480, 100510, 100540, 
    100570, 100610, 100640, 100680, 100720, 100760, 100800, 100830, 100890, 
    100930, 100960, 101040, 101090, 101150, 101190, 101220, 101270, 101290, 
    101310, 101340, 101340, 101360, 101390, 101400, 101390, 101420, 101460, 
    101500, 101530, 101540, 101570, 101590, 101610, 101650, 101670, 101700, 
    101730, 101760, 101780, 101800, 101820, 101830, 101840, 101850, 101860, 
    101890, 101900, 101910, 101920, 101920, 101880, 101860, 101820, 101790, 
    101760, 101740, 101730, 101690, 101670, 101650, 101630, 101610, 101560, 
    101520, 101500, 101450, 101440, 101450, 101450, 101460, 101470, 101480, 
    101490, 101500, 101480, 101480, 101450, 101450, 101430, 101420, 101440, 
    101450, 101460, 101460, 101430, 101440, 101430, 101430, 101420, 101420, 
    101410, 101410, 101430, 101420, 101410, 101400, 101400, 101400, 101400, 
    101390, 101380, 101370, 101390, 101380, 101400, 101410, 101420, 101420, 
    101420, 101440, 101450, 101470, 101490, 101480, 101490, 101510, 101520, 
    101540, 101560, 101560, 101560, 101570, 101590, 101600, 101590, 101590, 
    101590, 101590, 101590, 101570, 101560, 101560, 101570, 101560, 101560, 
    101550, 101540, 101490, 101450, 101410, 101380, 101360, 101340, 101300, 
    101260, 101230, 101200, 101160, 101130, 101110, 101080, 101040, 101010, 
    100990, 100980, 100980, 100980, 100930, 100910, 100870, 100850, 100800, 
    100730, 100640, 100590, 100480, 100400, 100350, 100300, 100300, 100360, 
    100390, 100390, 100390, 100390, 100430, 100440, 100460, 100470, 100490, 
    100510, 100510, 100510, 100500, 100520, 100490, 100470, 100480, 100490, 
    100560, 100620, 100710, 100820, 100910, 101030, 101130, 101260, 101320, 
    101430, 101490, 101620, 101720, 101830, 101940, 102030, 102120, 102240, 
    102350, 102370, 102430, 102530, 102580, 102630, 102690, 102750, 102810, 
    102880, 102920, 102950, 102990, 103030, 103060, 103070, 103080, 103100, 
    103120, 103140, 103140, 103150, 103160, 103150, 103140, 103120, 103090, 
    103080, 103050, 103010, 103000, 102980, 102950, 102930, 102900, 102860, 
    102820, 102790, 102730, 102680, 102640, 102580, 102530, 102490, 102440, 
    102380, 102330, 102270, 102200, 102140, 102080, 102020, 101980, 101910, 
    101860, 101810, 101760, 101710, 101680, 101640, 101620, 101590, 101560, 
    101510, 101490, 101460, 101450, 101440, 101420, 101420, 101420, 101410, 
    101410, 101410, 101430, 101460, 101490, 101530, 101590, 101660, 101740, 
    101790, 101830, 101890, 101940, 101970, 102010, 101990, 102010, 102000, 
    102020, 102000, 102000, 102000, 101950, 101910, 101870, 101830, 101760, 
    101700, 101640, 101590, 101510, 101480, 101450, 101370, 101310, 101250, 
    101190, 101130, 101100, 101080, 101040, 101070, 101050, 101090, 101090, 
    101110, 101130, 101120, 101150, 101190, 101210, 101200, 101220, 101260, 
    101280, 101310, 101330, 101360, 101370, 101390, 101410, 101400, 101430, 
    101420, 101400, 101440, 101430, 101400, 101430, 101440, 101400, 101420, 
    101440, 101430, 101440, 101430, 101420, 101440, 101440, 101450, 101460, 
    101520, 101570, 101600, 101620, 101640, 101670, 101690, 101730, 101760, 
    101800, 101860, 101900, 101940, 101960, 101980, 102010, 102020, 102030, 
    102030, 102040, 102060, 102080, 102120, 102120, 102120, 102140, 102160, 
    102180, 102170, 102150, 102130, 102110, 102090, 102080, 102070, 102050, 
    102010, 101990, 101980, 101950, 101930, 101880, 101850, 101830, 101800, 
    101790, 101770, 101760, 101720, 101710, 101690, 101640, 101630, 101620, 
    101590, 101550, 101520, 101500, 101490, 101450, 101440, 101430, 101410, 
    101380, 101360, 101340, 101310, 101290, 101280, 101270, 101260, 101250, 
    101230, 101230, 101210, 101210, 101190, 101180, 101170, 101170, 101180, 
    101190, 101190, 101210, 101220, 101250, 101270, 101280, 101280, 101290, 
    101290, 101280, 101300, 101320, 101350, 101400, 101420, 101430, 101440, 
    101440, 101420, 101430, 101430, 101430, 101440, 101450, 101450, 101430, 
    101420, 101410, 101380, 101370, 101360, 101340, 101320, 101320, 101320, 
    101330, 101310, 101300, 101290, 101320, 101320, 101270, 101270, 101270, 
    101270, 101260, 101240, 101260, 101280, 101280, 101280, 101270, 101250, 
    101240, 101210, 101190, 101160, 101130, 101100, 101060, 101030, 100990, 
    100950, 100910, 100850, 100810, 100780, 100740, 100690, 100660, 100630, 
    100570, 100540, 100500, 100490, 100490, 100490, 100500, 100520, 100520, 
    100510, 100520, 100550, 100580, 100600, 100630, 100660, 100700, 100710, 
    100730, 100720, 100730, 100750, 100760, 100770, 100800, 100820, 100840, 
    100880, 100890, 100900, 100910, 100910, 100920, 100910, 100910, 100910, 
    100920, 100940, 100940, 100940, 100940, 100940, 100940, 100940, 100960, 
    100950, 100950, 100980, 101000, 101010, 101030, 101040, 101050, 101090, 
    101110, 101110, 101120, 101130, 101140, 101170, 101210, 101230, 101250, 
    101270, 101310, 101320, 101330, 101330, 101370, 101400, 101420, 101440, 
    101470, 101510, 101530, 101560, 101570, 101600, 101620, 101630, 101640, 
    101680, 101670, 101700, 101710, 101750, 101740, 101740, 101740, 101760, 
    101760, 101760, 101760, 101770, 101740, 101700, 101700, 101670, 101660, 
    101640, 101620, 101580, 101540, 101450, 101390, 101380, 101350, 101270, 
    101190, 101080, 101050, 101000, 100900, 100820, 100740, 100660, 100610, 
    100520, 100510, 100480, 100460, 100450, 100430, 100460, 100430, 100400, 
    100390, 100340, 100320, 100310, 100310, 100280, 100280, 100280, 100300, 
    100320, 100370, 100360, 100380, 100390, 100390, 100400, 100420, 100440, 
    100480, 100510, 100530, 100550, 100540, 100550, 100560, 100580, 100610, 
    100630, 100640, 100640, 100670, 100670, 100690, 100720, 100730, 100740, 
    100760, 100770, 100800, 100810, 100840, 100830, 100840, 100900, 100950, 
    100940, 100930, 100910, 100900, 100850, 100820, 100790, 100770, 100750, 
    100740, 100730, 100730, 100720, 100700, 100690, 100670, 100650, 100630, 
    100620, 100610, 100600, 100600, 100590, 100610, 100600, 100600, 100590, 
    100570, 100550, 100520, 100490, 100490, 100470, 100460, 100450, 100440, 
    100440, 100420, 100420, 100420, 100420, 100420, 100390, 100390, 100380, 
    100370, 100370, 100370, 100360, 100330, 100340, 100300, 100300, 100300, 
    100290, 100270, 100280, 100290, 100290, 100310, 100330, 100360, 100400, 
    100440, 100470, 100470, 100490, 100470, 100510, 100530, 100540, 100570, 
    100580, 100580, 100600, 100620, 100620, 100620, 100640, 100660, 100680, 
    100700, 100730, 100730, 100750, 100750, 100760, 100760, 100780, 100780, 
    100770, 100740, 100710, 100710, 100710, 100710, 100690, 100700, 100700, 
    100680, 100670, 100660, 100640, 100620, 100630, 100630, 100640, 100600, 
    100610, 100600, 100620, 100620, 100600, 100600, 100580, 100570, 100550, 
    100520, 100520, 100500, 100490, 100460, 100430, 100410, 100390, 100370, 
    100360, 100370, 100340, 100350, 100360, 100400, 100450, 100460, 100500, 
    100520, 100510, 100550, 100560, 100580, 100600, 100620, 100640, 100670, 
    100650, 100660, 100650, 100650, 100650, 100650, 100640, 100630, 100640, 
    100630, 100660, 100680, 100710, 100720, 100760, 100760, 100790, 100820, 
    100830, 100840, 100870, 100900, 100950, 100990, 101010, 101050, 101070, 
    101100, 101130, 101150, 101160, 101180, 101220, 101260, 101290, 101330, 
    101350, 101380, 101410, 101430, 101440, 101450, 101450, 101470, 101480, 
    101490, 101490, 101500, 101520, 101510, 101520, 101510, 101490, 101480, 
    101490, 101460, 101440, 101420, 101420, 101430, 101400, 101390, 101380, 
    101360, 101300, 101260, 101240, 101200, 101160, 101140, 101130, 101100, 
    101040, 101010, 101000, 100960, 100930, 100890, 100850, 100810, 100790, 
    100790, 100810, 100840, 100860, 100890, 100880, 100880, 100890, 100890, 
    100910, 100920, 100940, 100960, 100980, 101010, 101020, 101030, 101020, 
    101030, 101010, 101020, 101000, 101010, 101030, 101010, 101020, 101030, 
    101020, 101030, 101020, 101040, 101030, 101030, 101030, 101040, 101050, 
    101060, 101080, 101110, 101140, 101150, 101160, 101180, 101190, 101220, 
    101250, 101250, 101270, 101290, 101320, 101330, 101350, 101380, 101380, 
    101390, 101390, 101410, 101420, 101430, 101460, 101450, 101470, 101480, 
    101490, 101510, 101510, 101520, 101530, 101530, 101510, 101500, 101500, 
    101510, 101520, 101500, 101510, 101510, 101480, 101480, 101460, 101430, 
    101410, 101370, 101350, 101350, 101330, 101340, 101340, 101310, 101290, 
    101270, 101250, 101240, 101240, 101240, 101240, 101240, 101230, 101240, 
    101250, 101250, 101250, 101240, 101220, 101220, 101220, 101200, 101200, 
    101220, 101210, 101210, 101200, 101190, 101180, 101170, 101160, 101120, 
    101090, 101080, 101040, 101010, 100960, 100960, 100930, 100900, 100870, 
    100840, 100820, 100790, 100760, 100750, 100720, 100720, 100700, 100720, 
    100720, 100710, 100690, 100670, 100630, 100570, 100520, 100510, 100470, 
    100420, 100390, 100330, 100280, 100220, 100180, 100120, 100070, 100020, 
    99890, 99840, 99780, 99670, 99530, 99370, 99190, 99050, 99090, 98900, 
    98960, 98990, 98980, 98930, 98920, 98980, 99030, 99100, 99200, 99320, 
    99420, 99520, 99600, 99690, 99800, 99860, 99950, 100030, 100110, 100180, 
    100280, 100360, 100410, 100470, 100540, 100570, 100620, 100690, 100730, 
    100800, 100870, 100960, 101020, 101080, 101150, 101220, 101250, 101300, 
    101340, 101370, 101420, 101460, 101500, 101570, 101610, 101640, 101660, 
    101680, 101720, 101740, 101720, 101720, 101740, 101760, 101780, 101800, 
    101800, 101810, 101810, 101800, 101780, 101800, 101790, 101790, 101770, 
    101790, 101810, 101810, 101800, 101770, 101760, 101770, 101760, 101740, 
    101710, 101690, 101690, 101720, 101690, 101690, 101700, 101720, 101710, 
    101720, 101710, 101670, 101660, 101670, 101690, 101700, 101720, 101720, 
    101740, 101750, 101760, 101780, 101760, 101770, 101790, 101810, 101840, 
    101880, 101900, 101930, 101960, 101990, 102010, 102040, 102030, 102030, 
    102040, 102050, 102070, 102110, 102110, 102120, 102110, 102120, 102100, 
    102120, 102110, 102110, 102090, 102060, 102070, 102060, 102060, 102040, 
    102030, 102040, 102030, 102010, 102000, 101970, 101910, 101880, 101870, 
    101850, 101830, 101810, 101800, 101780, 101760, 101740, 101710, 101700, 
    101650, 101620, 101610, 101610, 101630, 101600, 101620, 101590, 101560, 
    101550, 101530, 101500, 101480, 101470, 101440, 101440, 101400, 101390, 
    101430, 101430, 101430, 101420, 101370, 101350, 101310, 101260, 101250, 
    101280, 101240, 101250, 101210, 101190, 101150, 101110, 101050, 100990, 
    100990, 100980, 100960, 100960, 100980, 101000, 100950, 100940, 100930, 
    100940, 100920, 100900, 100870, 100890, 100900, 100920, 100980, 101000, 
    101040, 101040, 101040, 101050, 101020, 101010, 100990, 100970, 100960, 
    100950, 100940, 100930, 100870, 100840, 100860, 100790, 100770, 100780, 
    100780, 100780, 100800, 100820, 100830, 100840, 100880, 100880, 100910, 
    100940, 100950, 100930, 100890, 100880, 100900, 100920, 100900, 100880, 
    100880, 100880, 100840, 100810, 100770, 100750, 100750, 100760, 100750, 
    100700, 100670, 100650, 100650, 100640, 100630, 100620, 100600, 100590, 
    100570, 100580, 100600, 100600, 100600, 100610, 100620, 100620, 100610, 
    100620, 100610, 100600, 100590, 100580, 100590, 100580, 100590, 100600, 
    100600, 100620, 100620, 100610, 100610, 100630, 100630, 100620, 100620, 
    100620, 100630, 100630, 100630, 100620, 100620, 100640, 100630, 100620, 
    100600, 100590, 100610, 100590, 100600, 100610, 100630, 100650, 100650, 
    100660, 100670, 100680, 100680, 100700, 100710, 100720, 100730, 100770, 
    100770, 100810, 100820, 100820, 100820, 100830, 100820, 100820, 100820, 
    100840, 100840, 100840, 100840, 100860, 100840, 100830, 100830, 100810, 
    100780, 100790, 100780, 100770, 100780, 100780, 100780, 100760, 100750, 
    100720, 100670, 100630, 100630, 100610, 100580, 100590, 100570, 100570, 
    100570, 100560, 100530, 100480, 100440, 100430, 100390, 100360, 100300, 
    100290, 100280, 100240, 100250, 100260, 100230, 100140, 100080, 99980, 
    99900, 99860, 99830, 99770, 99760, 99760, 99780, 99810, 99810, 99820, 
    99820, 99820, 99830, 99810, 99820, 99820, 99810, 99780, 99750, 99760, 
    99760, 99750, 99720, 99710, 99690, 99700, 99700, 99700, 99700, 99690, 
    99710, 99740, 99760, 99780, 99800, 99810, 99820, 99860, 99910, 99960, 
    100000, 100060, 100110, 100160, 100220, 100290, 100330, 100380, 100410, 
    100460, 100510, 100560, 100620, 100690, 100740, 100800, 100860, 100900, 
    100940, 100960, 100990, 101040, 101110, 101160, 101200, 101250, 101300, 
    101350, 101420, 101450, 101470, 101490, 101510, 101520, 101530, 101570, 
    101570, 101580, 101590, 101610, 101620, 101640, 101640, 101620, 101630, 
    101640, 101650, 101660, 101660, 101670, 101710, 101720, 101720, 101700, 
    101710, 101690, 101660, 101660, 101670, 101680, 101680, 101690, 101690, 
    101670, 101680, 101680, 101670, 101650, 101650, 101640, 101630, 101620, 
    101640, 101630, 101640, 101620, 101610, 101620, 101620, 101580, 101560, 
    101520, 101520, 101490, 101470, 101450, 101430, 101420, 101390, 101360, 
    101300, 101260, 101220, 101200, 101190, 101200, 101230, 101270, 101280, 
    101300, 101300, 101340, 101380, 101420, 101450, 101480, 101510, 101540, 
    101580, 101600, 101610, 101660, 101670, 101700, 101720, 101730, 101740, 
    101760, 101800, 101810, 101850, 101880, 101900, 101920, 101940, 101940, 
    101950, 101960, 101960, 101990, 102000, 102030, 102050, 102080, 102090, 
    102100, 102120, 102130, 102130, 102140, 102130, 102130, 102130, 102150, 
    102180, 102200, 102220, 102210, 102220, 102220, 102220, 102220, 102210, 
    102200, 102210, 102200, 102180, 102180, 102150, 102130, 102130, 102110, 
    102100, 102080, 102060, 102050, 102030, 102020, 102010, 102040, 102040, 
    102020, 102010, 102000, 102010, 102000, 101990, 101960, 101940, 101940, 
    101950, 101960, 101950, 101940, 101930, 101900, 101860, 101840, 101830, 
    101790, 101760, 101740, 101730, 101710, 101680, 101630, 101610, 101560, 
    101540, 101510, 101460, 101430, 101390, 101370, 101360, 101350, 101330, 
    101320, 101310, 101290, 101270, 101290, 101290, 101300, 101290, 101290, 
    101290, 101300, 101300, 101300, 101320, 101310, 101310, 101320, 101340, 
    101340, 101340, 101350, 101370, 101390, 101370, 101330, 101290, 101250, 
    101210, 101170, 101140, 101100, 101040, 100950, 100880, 100890, 100890, 
    100900, 100920, 100920, 100920, 100930, 100930, 100930, 100920, 100920, 
    100930, 100960, 100970, 100980, 100960, 100950, 100930, 100930, 100930, 
    100940, 100930, 100930, 100940, 100960, 100960, 100980, 101020, 101020, 
    101030, 101030, 101050, 101030, 101040, 101060, 101070, 101090, 101110, 
    101130, 101160, 101170, 101170, 101160, 101170, 101180, 101200, 101230, 
    101240, 101290, 101320, 101330, 101350, 101380, 101360, 101360, 101380, 
    101370, 101350, 101350, 101360, 101360, 101360, 101360, 101350, 101340, 
    101310, 101280, 101250, 101240, 101220, 101240, 101250, 101280, 101290, 
    101270, 101270, 101250, 101240, 101220, 101190, 101170, 101150, 101120, 
    101110, 101100, 101090, 101060, 101040, 101010, 100990, 100960, 100930, 
    100910, 100890, 100890, 100900, 100910, 100910, 100880, 100850, 100840, 
    100820, 100800, 100770, 100750, 100730, 100700, 100710, 100690, 100680, 
    100680, 100670, 100660, 100660, 100640, 100610, 100600, 100590, 100570, 
    100590, 100570, 100580, 100580, 100580, 100570, 100560, 100540, 100510, 
    100500, 100470, 100460, 100460, 100450, 100450, 100450, 100440, 100440, 
    100420, 100390, 100380, 100330, 100310, 100310, 100290, 100290, 100290, 
    100290, 100280, 100250, 100240, 100240, 100230, 100220, 100230, 100220, 
    100230, 100240, 100240, 100250, 100250, 100240, 100230, 100230, 100210, 
    100200, 100190, 100170, 100170, 100140, 100120, 100110, 100080, 100050, 
    100020, 100000, 99980, 99950, 99930, 99920, 99910, 99900, 99900, 99890, 
    99870, 99850, 99830, 99820, 99820, 99800, 99790, 99780, 99780, 99790, 
    99810, 99810, 99810, 99800, 99790, 99770, 99780, 99760, 99770, 99790, 
    99800, 99830, 99860, 99890, 99920, 99950, 99960, 99970, 99990, 100060, 
    100080, 100100, 100140, 100160, 100180, 100190, 100190, 100200, 100210, 
    100200, 100220, 100220, 100210, 100210, 100210, 100250, 100250, 100230, 
    100190, 100180, 100170, 100180, 100170, 100170, 100170, 100160, 100160, 
    100140, 100120, 100130, 100120, 100100, 100080, 100060, 100030, 100000, 
    99990, 100000, 99990, 99960, 99960, 99950, 99930, 99920, 99950, 99920, 
    99950, 99960, 99990, 100010, 100060, 100070, 100120, 100140, 100170, 
    100200, 100230, 100260, 100290, 100310, 100340, 100360, 100380, 100400, 
    100420, 100420, 100430, 100430, 100430, 100440, 100480, 100480, 100500, 
    100530, 100550, 100580, 100580, 100600, 100610, 100580, 100590, 100590, 
    100580, 100580, 100570, 100550, 100540, 100530, 100540, 100540, 100510, 
    100500, 100480, 100460, 100430, 100410, 100410, 100390, 100390, 100380, 
    100370, 100360, 100370, 100370, 100370, 100370, 100370, 100390, 100430, 
    100460, 100460, 100490, 100510, 100530, 100550, 100560, 100570, 100580, 
    100570, 100580, 100610, 100610, 100600, 100590, 100590, 100590, 100550, 
    100520, 100480, 100420, 100390, 100350, 100310, 100310, 100270, 100250, 
    100250, 100270, 100300, 100360, 100370, 100450, 100500, 100550, 100580, 
    100630, 100660, 100720, 100780, 100840, 100900, 100960, 101010, 101050, 
    101110, 101150, 101170, 101220, 101260, 101310, 101320, 101330, 101330, 
    101320, 101300, 101300, 101300, 101300, 101300, 101300, 101290, 101290, 
    101290, 101300, 101310, 101310, 101310, 101330, 101360, 101400, 101420, 
    101460, 101460, 101470, 101520, 101540, 101540, 101520, 101520, 101510, 
    101480, 101470, 101490, 101470, 101430, 101390, 101370, 101320, 101250, 
    101160, 101100, 101000, 100870, 100780, 100680, 100610, 100550, 100510, 
    100460, 100420, 100400, 100370, 100350, 100370, 100370, 100390, 100430, 
    100470, 100520, 100590, 100670, 100780, 100840, 100880, 100980, 101050, 
    101090, 101150, 101200, 101230, 101230, 101250, 101210, 101200, 101150, 
    101080, 100980, 101020, 101000, 100980, 100960, 100940, 100940, 100950, 
    100940, 100910, 100910, 100920, 100930, 100970, 101000, 101050, 101120, 
    101160, 101210, 101240, 101260, 101260, 101250, 101210, 101180, 101160, 
    101150, 101150, 101130, 101140, 101130, 101110, 101090, 101060, 101040, 
    101010, 100980, 100940, 100900, 100870, 100830, 100790, 100760, 100710, 
    100660, 100610, 100560, 100470, 100390, 100320, 100250, 100220, 100170, 
    100090, 100060, 100030, 99970, 99940, 99960, 99980, 99980, 99960, 100000, 
    100030, 100050, 100070, 100070, 100050, 100100, 100110, 100110, 100150, 
    100180, 100230, 100250, 100280, 100330, 100400, 100420, 100440, 100470, 
    100500, 100550, 100610, 100610, 100600, 100580, 100600, 100590, 100630, 
    100590, 100570, 100550, 100510, 100460, 100450, 100480, 100490, 100510, 
    100550, 100560, 100620, 100660, 100740, 100830, 100910, 100990, 101100, 
    101200, 101300, 101390, 101470, 101550, 101600, 101660, 101730, 101790, 
    101820, 101850, 101860, 101880, 101900, 101920, 101940, 101940, 101930, 
    101940, 101980, 101970, 101920, 101910, 101890, 101860, 101820, 101760, 
    101670, 101610, 101550, 101500, 101440, 101360, 101290, 101240, 101160, 
    101050, 100950, 100890, 100830, 100740, 100660, 100620, 100540, 100460, 
    100380, 100280, 100180, 100090, 100030, 99980, 99960, 99960, 99990, 
    100070, 100120, 100150, 100200, 100210, 100250, 100290, 100330, 100400, 
    100450, 100510, 100550, 100630, 100700, 100730, 100780, 100820, 100840, 
    100860, 100850, 100840, 100830, 100820, 100830, 100840, 100910, 100930, 
    100950, 100970, 100980, 100960, 100980, 100980, 100970, 100950, 100950, 
    100930, 100920, 100900, 100860, 100800, 100760, 100690, 100650, 100600, 
    100560, 100540, 100490, 100460, 100440, 100400, 100380, 100350, 100320, 
    100280, 100220, 100160, 100080, 100020, 99960, 99870, 99760, 99670, 
    99600, 99540, 99540, 99510, 99490, 99450, 99400, 99320, 99200, 99110, 
    99000, 98940, 98880, 98820, 98760, 98720, 98630, 98550, 98490, 98370, 
    98300, 98210, 98180, 98130, 98040, 98010, 97930, 97840, 97810, 97790, 
    97770, 97770, 97820, 97860, 97940, 97980, 98050, 98110, 98170, 98220, 
    98310, 98380, 98450, 98530, 98620, 98720, 98830, 98920, 98980, 99050, 
    99120, 99180, 99220, 99270, 99310, 99330, 99350, 99390, 99420, 99440, 
    99440, 99420, 99420, 99360, 99340, 99290, 99280, 99240, 99230, 99200, 
    99180, 99140, 99110, 99070, 99020, 98980, 98950, 98930, 98930, 98930, 
    98960, 98960, 98980, 99000, 99000, 99000, 99000, 99000, 99000, 99050, 
    99050, 99060, 99070, 99090, 99120, 99130, 99130, 99110, 99110, 99080, 
    99060, 99040, 99050, 99020, 99010, 98990, 98990, 98980, 98960, 98950, 
    98940, 98950, 98960, 98950, 98960, 98970, 98980, 98980, 98980, 98980, 
    98970, 98990, 99010, 99010, 99030, 99060, 99100, 99150, 99200, 99270, 
    99330, 99390, 99440, 99500, 99560, 99650, 99730, 99800, 99860, 99910, 
    99980, 100050, 100110, 100150, 100220, 100290, 100340, 100370, 100410, 
    100450, 100490, 100520, 100560, 100590, 100620, 100630, 100650, 100680, 
    100700, 100700, 100710, 100710, 100720, 100740, 100730, 100720, 100730, 
    100730, 100740, 100750, 100740, 100730, 100740, 100760, 100770, 100770, 
    100770, 100770, 100780, 100800, 100820, 100840, 100850, 100850, 100890, 
    100900, 100920, 100940, 100970, 100990, 101000, 101020, 101070, 101090, 
    101010, 101140, 101160, 101180, 101210, 101240, 101230, 101220, 101230, 
    101240, 101250, 101280, 101250, 101240, 101240, 101230, 101220, 101210, 
    101190, 101160, 101130, 101100, 101090, 101100, 101070, 101030, 101000, 
    100980, 100930, 100910, 100880, 100860, 100840, 100820, 100800, 100770, 
    100750, 100690, 100650, 100620, 100600, 100560, 100540, 100520, 100490, 
    100470, 100430, 100440, 100430, 100440, 100410, 100420, 100410, 100440, 
    100460, 100490, 100530, 100580, 100630, 100660, 100710, 100760, 100790, 
    100830, 100880, 100910, 100940, 100990, 101040, 101080, 101120, 101150, 
    101180, 101210, 101210, 101260, 101290, 101310, 101350, 101400, 101440, 
    101480, 101500, 101520, 101540, 101530, 101560, 101570, 101570, 101590, 
    101620, 101640, 101660, 101680, 101700, 101720, 101730, 101730, 101740, 
    101770, 101760, 101750, 101790, 101820, 101830, 101870, 101860, 101850, 
    101860, 101860, 101850, 101850, 101890, 101900, 101940, 101950, 101950, 
    101940, 101930, 101940, 101940, 101930, 101910, 101890, 101860, 101840, 
    101840, 101840, 101810, 101770, 101750, 101730, 101710, 101660, 101630, 
    101600, 101580, 101570, 101570, 101560, 101550, 101510, 101500, 101480, 
    101430, 101380, 101370, 101360, 101360, 101370, 101370, 101320, 101370, 
    101330, 101310, 101330, 101350, 101350, 101340, 101340, 101330, 101340, 
    101380, 101400, 101360, 101370, 101410, 101400, 101410, 101420, 101410, 
    101430, 101450, 101490, 101500, 101530, 101540, 101540, 101540, 101540, 
    101550, 101570, 101550, 101560, 101560, 101570, 101590, 101600, 101580, 
    101550, 101530, 101550, 101530, 101490, 101460, 101420, 101380, 101350, 
    101340, 101300, 101270, 101240, 101120, 101040, 100980, 100860, 100740, 
    100610, 100480, 100350, 100270, 100190, 100090, 99980, 99860, 99740, 
    99670, 99590, 99500, 99400, 99290, 99180, 99090, 99030, 98980, 98950, 
    98960, 98970, 98980, 99010, 99030, 99060, 99130, 99150, 99210, 99300, 
    99420, 99500, 99580, 99700, 99820, 99960, 100080, 100160, 100250, 100330, 
    100450, 100560, 100670, 100750, 100820, 100860, 100940, 101010, 101100, 
    101150, 101200, 101270, 101350, 101400, 101450, 101500, 101530, 101560, 
    101580, 101620, 101640, 101660, 101690, 101700, 101720, 101720, 101730, 
    101720, 101710, 101670, 101690, 101690, 101690, 101670, 101640, 101610, 
    101580, 101550, 101510, 101470, 101400, 101280, 101260, 101240, 101190, 
    101100, 101000, 100920, 100850, 100760, 100680, 100640, 100590, 100510, 
    100470, 100370, 100370, 100340, 100300, 100290, 100280, 100280, 100300, 
    100330, 100350, 100350, 100350, 100350, 100340, 100320, 100270, 100180, 
    100090, 99990, 99890, 99760, 99590, 99420, 99270, 99060, 98940, 98870, 
    98760, 98700, 98750, 98850, 98900, 98990, 99180, 99280, 99440, 99630, 
    99890, 100030, 100120, 100140, 100260, 100320, 100380, 100440, 100470, 
    100480, 100490, 100500, 100530, 100560, 100580, 100630, 100700, 100760, 
    100840, 100910, 100950, 100970, 101020, 101030, 101070, 101090, 101090, 
    101100, 101110, 101140, 101190, 101180, 101190, 101180, 101200, 101220, 
    101260, 101290, 101340, 101400, 101430, 101430, 101420, 101380, 101340, 
    101240, 101160, 101010, 100840, 100650, 100550, 100510, 100580, 100660, 
    100700, 100730, 100710, 100750, 100780, 100800, 100830, 100880, 100980, 
    101040, 101050, 101080, 101110, 101130, 101120, 101070, 101020, 100970, 
    100920, 100930, 100930, 100960, 101010, 101050, 101080, 101140, 101200, 
    101290, 101360, 101430, 101490, 101550, 101610, 101640, 101710, 101740, 
    101780, 101810, 101780, 101770, 101770, 101720, 101720, 101670, 101630, 
    101610, 101580, 101540, 101520, 101530, 101510, 101510, 101520, 101520, 
    101510, 101510, 101540, 101560, 101570, 101560, 101550, 101540, 101540, 
    101510, 101500, 101510, 101520, 101520, 101540, 101550, 101570, 101570, 
    101580, 101590, 101590, 101570, 101540, 101520, 101500, 101490, 101490, 
    101490, 101490, 101510, 101520, 101520, 101520, 101500, 101510, 101640, 
    101510, 101510, 101510, 101540, 101560, 101580, 101580, 101610, 101610, 
    101610, 101630, 101660, 101690, 101700, 101710, 101720, 101750, 101770, 
    101790, 101800, 101790, 101790, 101810, 101800, 101800, 101790, 101790, 
    101810, 101810, 101800, 101780, 101740, 101700, 101640, 101590, 101560, 
    101510, 101450, 101390, 101310, 101240, 101170, 101090, 100990, 100910, 
    100840, 100730, 100660, 100630, 100590, 100570, 100560, 100580, 100590, 
    100610, 100590, 100580, 100580, 100550, 100530, 100490, 100470, 100430, 
    100440, 100440, 100410, 100370, 100350, 100310, 100280, 100260, 100250, 
    100230, 100200, 100200, 100210, 100220, 100240, 100230, 100230, 100220, 
    100220, 100230, 100220, 100230, 100200, 100180, 100210, 100230, 100210, 
    100180, 100190, 100190, 100160, 100130, 100110, 100030, 100090, 100040, 
    100020, 100010, 99960, 99910, 99880, 99840, 99780, 99700, 99640, 99610, 
    99530, 99470, 99390, 99300, 99260, 99190, 99080, 99020, 99970, 98930, 
    98880, 98810, 98770, 98720, 98720, 98690, 98710, 98710, 98740, 98730, 
    98770, 98760, 98770, 98790, 98800, 98810, 98840, 98850, 98850, 98890, 
    98920, 98860, 98860, 98880, 98870, 98850, 98820, 98830, 98850, 98830, 
    98840, 98820, 98820, 98780, 98810, 98810, 98830, 98880, 98920, 98970, 
    98980, 99000, 98990, 99030, 99050, 99060, 99060, 99090, 99100, 99130, 
    99160, 99210, 99290, 99350, 99400, 99450, 99510, 99560, 99620, 99680, 
    99760, 99810, 99870, 99930, 100010, 100110, 100200, 100290, 100380, 
    100470, 100560, 100670, 100770, 100890, 100990, 101070, 101150, 101240, 
    101280, 101300, 101300, 101260, 101260, 101320, 101320, 101380, 101440, 
    101520, 101580, 101730, 101860, 102010, 102120, 102220, 102270, 102270, 
    102310, 102310, 102270, 102240, 102210, 102180, 102140, 102080, 101990, 
    101880, 101810, 101760, 101730, 101680, 101690, 101630, 101560, 101460, 
    101380, 101330, 101260, 101160, 101050, 100920, 100770, 100610, 100500, 
    100440, 100380, 100360, 100380, 100400, 100450, 100490, 100490, 100500, 
    100560, 100660, 100740, 100860, 100980, 101100, 101230, 101370, 101490, 
    101610, 101760, 101910, 102080, 102150, 102220, 102330, 102410, 102460, 
    102550, 102610, 102610, 102600, 102640, 102610, 102610, 102580, 102550, 
    102500, 102390, 102290, 102180, 102060, 101950, 101820, 101700, 101560, 
    101430, 101350, 101210, 101080, 101000, 100940, 100880, 100850, 100880, 
    101060, 101090, 101130, 101160, 101110, 101100, 101100, 101260, 101320, 
    101500, 101610, 101730, 101830, 101940, 102020, 102120, 102200, 102260, 
    102300, 102330, 102360, 102410, 102460, 102520, 102530, 102540, 102580, 
    102610, 102620, 102650, 102690, 102730, 102750, 102760, 102790, 102810, 
    102820, 102820, 102830, 102820, 102800, 102750, 102760, 102740, 102730, 
    102690, 102650, 102590, 102550, 102490, 102440, 102410, 102350, 102330, 
    102290, 102240, 102190, 102170, 102090, 102040, 102000, 101960, 101880, 
    101820, 101800, 101730, 101720, 101690, 101700, 101700, 101690, 101660, 
    101660, 101670, 101640, 101640, 101650, 101650, 101640, 101630, 101620, 
    101610, 101580, 101550, 101490, 101430, 101370, 101290, 101200, 101110, 
    101070, 101000, 100950, 100850, 100760, 100670, 100620, 100590, 100600, 
    100610, 100630, 100670, 100740, 100800, 100850, 100910, 100960, 101020, 
    101060, 101130, 101150, 101180, 101200, 101250, 101280, 101350, 101400, 
    101440, 101470, 101500, 101520, 101530, 101540, 101550, 101580, 101600, 
    101630, 101660, 101680, 101700, 101710, 101740, 101760, 101790, 101810, 
    101840, 101830, 101870, 101910, 101940, 101960, 101980, 102010, 102020, 
    102040, 102090, 102090, 102090, 102090, 102110, 102110, 102110, 102110, 
    102100, 102110, 102090, 102050, 101990, 101930, 101840, 101760, 101680, 
    101590, 101490, 101380, 101300, 101220, 101150, 101070, 100990, 100950, 
    100880, 100790, 100740, 100700, 100630, 100550, 100530, 100470, 100410, 
    100380, 100300, 100230, 100150, 100050, 99970, 99920, 99900, 99980, 
    100010, 100070, 100050, 100040, 100170, 100300, 100380, 100370, 100410, 
    100490, 100510, 100610, 100700, 100750, 100810, 100830, 100960, 101060, 
    101140, 101230, 101290, 101330, 101370, 101420, 101470, 101510, 101520, 
    101520, 101500, 101520, 101490, 101480, 101460, 101420, 101410, 101400, 
    101400, 101400, 101420, 101440, 101450, 101430, 101440, 101470, 101470, 
    101470, 101480, 101500, 101490, 101500, 101510, 101500, 101500, 101490, 
    101490, 101480, 101470, 101450, 101440, 101470, 101480, 101490, 101490, 
    101470, 101470, 101470, 101470, 101500, 101500, 101500, 101530, 101550, 
    101560, 101560, 101550, 101520, 101530, 101530, 101510, 101500, 101530, 
    101510, 101490, 101490, 101490, 101490, 101500, 101490, 101480, 101450, 
    101450, 101440, 101410, 101410, 101400, 101400, 101410, 101410, 101400, 
    101370, 101360, 101340, 101340, 101330, 101310, 101310, 101330, 101320, 
    101320, 101290, 101320, 101330, 101280, 101270, 101280, 101280, 101260, 
    101260, 101280, 101310, 101350, 101380, 101390, 101360, 101320, 101290, 
    101260, 101240, 101230, 101190, 101150, 101110, 101010, 101000, 100880, 
    100850, 100820, 100710, 100700, 100690, 100660, 100680, 100690, 100790, 
    100820, 100890, 100920, 100970, 101050, 101100, 101210, 101290, 101370, 
    101420, 101520, 101600, 101660, 101690, 101690, 101690, 101730, 101730, 
    101710, 101720, 101720, 101780, 101820, 101910, 101990, 102090, 102170, 
    102240, 102320, 102400, 102470, 102520, 102560, 102580, 102630, 102660, 
    102670, 102660, 102790, 102660, 102660, 102660, 102650, 102660, 102680, 
    102710, 102720, 102720, 102710, 102760, 102780, 102760, 102750, 102770, 
    102760, 102770, 102760, 102790, 102830, 102810, 102840, 102840, 102800, 
    102800, 102760, 102720, 102700, 102670, 102620, 102600, 102590, 102580, 
    102560, 102550, 102490, 102440, 102410, 102350, 102280, 102210, 102160, 
    102100, 102010, 101940, 101880, 101820, 101750, 101690, 101610, 101550, 
    101470, 101400, 101340, 101280, 101230, 101190, 101150, 101110, 101080, 
    101040, 101000, 100960, 100940, 100910, 100900, 100910, 100900, 100910, 
    100900, 100870, 100850, 100830, 100790, 100780, 100770, 100770, 100750, 
    100760, 100760, 100740, 100730, 100710, 100710, 100700, 100670, 100640, 
    100610, 100570, 100530, 100540, 100540, 100560, 100580, 100590, 100610, 
    100610, 100600, 100620, 100630, 100650, 100670, 100690, 100740, 100780, 
    100800, 100810, 100840, 100860, 100840, 100830, 100840, 100820, 100780, 
    100780, 100780, 100800, 100820, 100820, 100820, 100840, 100870, 100890, 
    100900, 100920, 100950, 100970, 101020, 101080, 101120, 101120, 101180, 
    101200, 101210, 101270, 101330, 101410, 101440, 101560, 101600, 101630, 
    101670, 101710, 101730, 101760, 101820, 101850, 101960, 102010, 102070, 
    102130, 102200, 102270, 102310, 102410, 102490, 102540, 102580, 102630, 
    102650, 102680, 102690, 102730, 102760, 102790, 102820, 102860, 102900, 
    102950, 102970, 103000, 103020, 103040, 103060, 103090, 103100, 103130, 
    103140, 103160, 103180, 103180, 103200, 103200, 103210, 103190, 103180, 
    103190, 103210, 103210, 103220, 103200, 103200, 103180, 103160, 103140, 
    103110, 103090, 103080, 103070, 103070, 103070, 103080, 103070, 103060, 
    103060, 103070, 103060, 103040, 103050, 103060, 103080, 103090, 103100, 
    103100, 103100, 103090, 103090, 103060, 103050, 103050, 103050, 103050, 
    103010, 103020, 103020, 103020, 103000, 102970, 102950, 102920, 102880, 
    102850, 102820, 102780, 102760, 102720, 102690, 102680, 102650, 102620, 
    102590, 102560, 102540, 102530, 102510, 102480, 102480, 102470, 102460, 
    102480, 102490, 102490, 102490, 102500, 102520, 102540, 102560, 102540, 
    102560, 102590, 102610, 102610, 102630, 102640, 102660, 102670, 102690, 
    102700, 102700, 102700, 102720, 102730, 102760, 102790, 102800, 102800, 
    102810, 102810, 102810, 102820, 102820, 102830, 102830, 102840, 102820, 
    102820, 102820, 102800, 102770, 102750, 102730, 102700, 102690, 102640, 
    102590, 102550, 102510, 102490, 102450, 102400, 102360, 102300, 102250, 
    102210, 102160, 102120, 102080, 102070, 102050, 102040, 102020, 102030, 
    102020, 102030, 102040, 102050, 102070, 102100, 102120, 102150, 102190, 
    102200, 102190, 102200, 102210, 102200, 102200, 102190, 102200, 102170, 
    102140, 102100, 102070, 102010, 101940, 101870, 101780, 101720, 101650, 
    101590, 101510, 101430, 101380, 101340, 101290, 101220, 101170, 101100, 
    101040, 100950, 100880, 100800, 100750, 100670, 100600, 100530, 100460, 
    100370, 100300, 100220, 100150, 100050, 99990, 99920, 99830, 99740, 
    99660, 99570, 99520, 99450, 99400, 99330, 99260, 99190, 99080, 99000, 
    98910, 98860, 98780, 98750, 98620, 98540, 98480, 98390, 98310, 98260, 
    98250, 98250, 98330, 98460, 98610, 98810, 98990, 99110, 99250, 99450, 
    99600, 99670, 99790, 99920, 99970, 100050, 100110, 100140, 100200, 
    100210, 100240, 100270, 100290, 100330, 100380, 100450, 100490, 100530, 
    100590, 100650, 100740, 100840, 100940, 101050, 101110, 101120, 101220, 
    101290, 101340, 101390, 101430, 101470, 101530, 101580, 101640, 101640, 
    101670, 101700, 101710, 101730, 101770, 101790, 101840, 101890, 101920, 
    101970, 101990, 102020, 102030, 102060, 102070, 102070, 102080, 102070, 
    102060, 102020, 102010, 102000, 102000, 101970, 101920, 101850, 101840, 
    101790, 101760, 101710, 101660, 101660, 101660, 101640, 101600, 101580, 
    101540, 101480, 101480, 101450, 101420, 101360, 101340, 101320, 101280, 
    101250, 101240, 101200, 101130, 101080, 101040, 100980, 100960, 100890, 
    100830, 100820, 100800, 100770, 100740, 100700, 100650, 100630, 100610, 
    100610, 100580, 100570, 100560, 100560, 100510, 100480, 100470, 100440, 
    100420, 100390, 100370, 100330, 100290, 100250, 100220, 100200, 100190, 
    100160, 100130, 100120, 100100, 100050, 100050, 100030, 99990, 99950, 
    99900, 99840, 99780, 99720, 99630, 99510, 99430, 99330, 99270, 99120, 
    99060, 98970, 98850, 98710, 98510, 98240, 98040, 97830, 97620, 97440, 
    97260, 97140, 97060, 97020, 96970, 96820, 96790, 96770, 96790, 96850, 
    96970, 97080, 97170, 97260, 97350, 97360, 97420, 97470, 97530, 97590, 
    97700, 97800, 97900, 97990, 98070, 98150, 98240, 98270, 98320, 98370, 
    98380, 98410, 98390, 98380, 98340, 98300, 98210, 98090, 97950, 97870, 
    97790, 97720, 97670, 97630, 97570, 97500, 97430, 97420, 97320, 97270, 
    97250, 97270, 97300, 97390, 97740, 97740, 98010, 98260, 98510, 98750, 
    98960, 99130, 99250, 99410, 99560, 99630, 99750, 99870, 99970, 100030, 
    100120, 100230, 100340, 100440, 100510, 100610, 100690, 100780, 100860, 
    100970, 101040, 101100, 101160, 101210, 101240, 101270, 101290, 101320, 
    101340, 101370, 101370, 101390, 101400, 101400, 101410, 101370, 101360, 
    101340, 101340, 101340, 101320, 101290, 101250, 101220, 101200, 101210, 
    101190, 101190, 101120, 101080, 101030, 100990, 100950, 100900, 100850, 
    100780, 100770, 100750, 100710, 100690, 100670, 100630, 100570, 100520, 
    100470, 100440, 100400, 100360, 100310, 100280, 100240, 100220, 100200, 
    100200, 100170, 100170, 100170, 100190, 100200, 100220, 100210, 100200, 
    100220, 100200, 100210, 100230, 100250, 100320, 100350, 100390, 100420, 
    100480, 100520, 100530, 100550, 100570, 100610, 100610, 100680, 100710, 
    100740, 100780, 100830, 100880, 100940, 100970, 101000, 101040, 101070, 
    101100, 101150, 101180, 101210, 101240, 101270, 101300, 101300, 101300, 
    101300, 101320, 101330, 101340, 101350, 101360, 101370, 101400, 101450, 
    101460, 101470, 101500, 101510, 101510, 101510, 101510, 101510, 101510, 
    101530, 101560, 101550, 101560, 101530, 101520, 101530, 101520, 101530, 
    101530, 101530, 101540, 101530, 101530, 101550, 101580, 101570, 101580, 
    101580, 101570, 101590, 101580, 101560, 101570, 101590, 101600, 101600, 
    101600, 101610, 101630, 101650, 101630, 101630, 101620, 101610, 101630, 
    101620, 101650, 101680, 101710, 101740, 101770, 101890, 101760, 101770, 
    101760, 101750, 101750, 101740, 101750, 101760, 101770, 101750, 101750, 
    101730, 101690, 101660, 101640, 101610, 101580, 101550, 101530, 101500, 
    101490, 101480, 101460, 101410, 101370, 101330, 101320, 101320, 101300, 
    101280, 101340, 101380, 101410, 101390, 101360, 101350, 101370, 101380, 
    101370, 101400, 101400, 101410, 101410, 101430, 101440, 101460, 101450, 
    101430, 101470, 101460, 101470, 101480, 101510, 101500, 101550, 101550, 
    101550, 101570, 101610, 101630, 101650, 101630, 101720, 101750, 101760, 
    101800, 101820, 101840, 101850, 101880, 101900, 101910, 101900, 101890, 
    101860, 101850, 101840, 101820, 101800, 101790, 101770, 101720, 101660, 
    101590, 101540, 101480, 101430, 101380, 101320, 101240, 101190, 101130, 
    101090, 101030, 100970, 100920, 100850, 100790, 100740, 100650, 100600, 
    100570, 100550, 100530, 100530, 100500, 100480, 100450, 100390, 100360, 
    100330, 100320, 100280, 100260, 100230, 100200, 100220, 100290, 100320, 
    100320, 100360, 100370, 100360, 100410, 100440, 100460, 100480, 100510, 
    100510, 100520, 100540, 100510, 100540, 100600, 100650, 100710, 100730, 
    100740, 100760, 100790, 100850, 100880, 100910, 100970, 100980, 101000, 
    101030, 101070, 101100, 101100, 101120, 101160, 101200, 101250, 101290, 
    101280, 101300, 101350, 101370, 101400, 101420, 101430, 101470, 101510, 
    101540, 101570, 101620, 101670, 101680, 101700, 101710, 101740, 101760, 
    101790, 101830, 101840, 101860, 101860, 101850, 101850, 101850, 101840, 
    101840, 101820, 101780, 101770, 101750, 101730, 101710, 101680, 101660, 
    101620, 101580, 101540, 101490, 101460, 101420, 101370, 101320, 101280, 
    101230, 101190, 101130, 101060, 101010, 100970, 100930, 100890, 100860, 
    100830, 100830, 100830, 100840, 100830, 100800, 100780, 100760, 100720, 
    100690, 100680, 100630, 100580, 100580, 100550, 100500, 100450, 100410, 
    100360, 100290, 100250, 100200, 100160, 100150, 100120, 100080, 100020, 
    99990, 99950, 99910, 99850, 99780, 99720, 99730, 99720, 99760, 99790, 
    99810, 99860, 99930, 100000, 100030, 100090, 100140, 100200, 100230, 
    100290, 100300, 100320, 100350, 100370, 100440, 100490, 100570, 100640, 
    100760, 100870, 100950, 101010, 101080, 101180, 101210, 101230, 101220, 
    101260, 101290, 101300, 101270, 101260, 101220, 101190, 101160, 101150, 
    101130, 101100, 101050, 101040, 101000, 100950, 100910, 100870, 100850, 
    100820, 100800, 100770, 100760, 100750, 100770, 100790, 100780, 100780, 
    100770, 100750, 100750, 100750, 100750, 100740, 100750, 100720, 100740, 
    100730, 100710, 100690, 100640, 100620, 100600, 100550, 100520, 100470, 
    100410, 100360, 100340, 100310, 100250, 100200, 100170, 100120, 100040, 
    99970, 99900, 99850, 99820, 99810, 99780, 99830, 99860, 99900, 99930, 
    99960, 100000, 100070, 100120, 100140, 100190, 100260, 100330, 100370, 
    100410, 100500, 100570, 100610, 100680, 100710, 100730, 100780, 100870, 
    100920, 100990, 101060, 101150, 101210, 101270, 101330, 101380, 101390, 
    101440, 101450, 101490, 101510, 101530, 101580, 101600, 101600, 101640, 
    101640, 101640, 101620, 101630, 101640, 101640, 101650, 101680, 101670, 
    101640, 101640, 101600, 101560, 101530, 101490, 101450, 101410, 101390, 
    101340, 101310, 101260, 101210, 101160, 101110, 101070, 101020, 100960, 
    100900, 100860, 100840, 100810, 100790, 100790, 100760, 100750, 100740, 
    100740, 100700, 100690, 100650, 100640, 100620, 100590, 100580, 100600, 
    100580, 100570, 100590, 100570, 100560, 100540, 100500, 100490, 100520, 
    100520, 100530, 100510, 100540, 100540, 100540, 100510, 100500, 100500, 
    100510, 100530, 100560, 100580, 100610, 100630, 100650, 100660, 100650, 
    100670, 100660, 100660, 100650, 100660, 100690, 100680, 100690, 100680, 
    100690, 100680, 100710, 100720, 100720, 100720, 100710, 100730, 100750, 
    100750, 100750, 100730, 100680, 100640, 100620, 100580, 100570, 100540, 
    100530, 100500, 100480, 100480, 100470, 100450, 100440, 100420, 100390, 
    100370, 100350, 100320, 100280, 100240, 100220, 100200, 100140, 100110, 
    100090, 100050, 100030, 100000, 100000, 99950, 99950, 99940, 99950, 
    99980, 100020, 100020, 100000, 99970, 99950, 99930, 99900, 99820, 99730, 
    99690, 99650, 99620, 99570, 99510, 99450, 99400, 99370, 99350, 99320, 
    99290, 99290, 99310, 99360, 99410, 99490, 99570, 99620, 99710, 99800, 
    99870, 99910, 99940, 99950, 100010, 100070, 100100, 100090, 100040, 
    100060, 99990, 99940, 99900, 99870, 99830, 99760, 99700, 99670, 99610, 
    99580, 99540, 99490, 99480, 99450, 99410, 99370, 99340, 99310, 99280, 
    99250, 99230, 99200, 99170, 99160, 99160, 99160, 99160, 99160, 99150, 
    99160, 99160, 99180, 99180, 99200, 99210, 99220, 99260, 99290, 99310, 
    99320, 99340, 99360, 99420, 99490, 99550, 99630, 99670, 99690, 99720, 
    99770, 99680, 99650, 99580, 99540, 99460, 99330, 99180, 99030, 98760, 
    98560, 98320, 97980, 97750, 97470, 97190, 96930, 96710, 96490, 96410, 
    96500, 96520, 96570, 96620, 96670, 96730, 96780, 96860, 96880, 96970, 
    97130, 97300, 97400, 97480, 97610, 97750, 97860, 97970, 98020, 98010, 
    98020, 98020, 98010, 98000, 97980, 97950, 97930, 97860, 97720, 97530, 
    97330, 97030, 96750, 96510, 96370, 96360, 96390, 96320, 96290, 96330, 
    96370, 96360, 96380, 96370, 96250, 96210, 96200, 96250, 96300, 96340, 
    96410, 96430, 96480, 96530, 96530, 96570, 96550, 96530, 96550, 96570, 
    96550, 96630, 96670, 96700, 96740, 96720, 96710, 96710, 96690, 96650, 
    96700, 96690, 96690, 96730, 96750, 96720, 96720, 96740, 96780, 96790, 
    96810, 96850, 96880, 96950, 97000, 97030, 97100, 97130, 97160, 97190, 
    97250, 97290, 97300, 97340, 97380, 97400, 97420, 97440, 97460, 97450, 
    97450, 97450, 97460, 97470, 97480, 97490, 97500, 97560, 97610, 97630, 
    97650, 97660, 97710, 97760, 97790, 97800, 97820, 97850, 97870, 97900, 
    97940, 97970, 98010, 98020, 98050, 98060, 98070, 98080, 98100, 98120, 
    98120, 98140, 98150, 98190, 98210, 98190, 98170, 98170, 98170, 98150, 
    98100, 98060, 98020, 98000, 98020, 97980, 97940, 97910, 97890, 97860, 
    97820, 97790, 97770, 97760, 97770, 97760, 97790, 97860, 97880, 97880, 
    97860, 97860, 97900, 97910, 98020, 98130, 98260, 98400, 98560, 98720, 
    98840, 98960, 99100, 99240, 99330, 99470, 99610, 99750, 99820, 99950, 
    100110, 100220, 100340, 100410, 100500, 100620, 100700, 100750, 100770, 
    100810, 100860, 100930, 100990, 101050, 101100, 101120, 101130, 101150, 
    101150, 101130, 101120, 101050, 100970, 100830, 100680, 100510, 100320, 
    100160, 99940, 99650, 99440, 99220, 99020, 98780, 98570, 98410, 98260, 
    98190, 98110, 98110, 98020, 98090, 98070, 98180, 98240, 98360, 98470, 
    98600, 98720, 98810, 98890, 98970, 99060, 99090, 99150, 99280, 99330, 
    99460, 99560, 99640, 99750, 99820, 99910, 99940, 99970, 100000, 100030, 
    100040, 100000, 99960, 100000, 100010, 100070, 100130, 100120, 100130, 
    100110, 100150, 100100, 100130, 100190, 100240, 100310, 100380, 100420, 
    100460, 100510, 100510, 100550, 100600, 100650, 100690, 100720, 100790, 
    100860, 100940, 101000, 101110, 101170, 101270, 101340, 101460, 101540, 
    101570, 101630, 101670, 101770, 101840, 101920, 101990, 102000, 102030, 
    102050, 102070, 102080, 102110, 102120, 102120, 102110, 102120, 102160, 
    102160, 102160, 102150, 102120, 102110, 102110, 102110, 102110, 102100, 
    102120, 102110, 102110, 102080, 102050, 102010, 101990, 101960, 101920, 
    101870, 101810, 101790, 101770, 101750, 101750, 101710, 101690, 101630, 
    101600, 101570, 101520, 101500, 101480, 101440, 101440, 101390, 101400, 
    101410, 101400, 101390, 101420, 101440, 101440, 101440, 101450, 101480, 
    101510, 101560, 101580, 101590, 101630, 101660, 101680, 101700, 101660, 
    101710, 101690, 101670, 101680, 101720, 101730, 101720, 101730, 101710, 
    101660, 101620, 101600, 101560, 101520, 101470, 101450, 101380, 101280, 
    101240, 101160, 101080, 100990, 100940, 100910, 100830, 100790, 100760, 
    100750, 100730, 100760, 100730, 100660, 100580, 100490, 100370, 100220, 
    100030, 99820, 99660, 99570, 99440, 99280, 99120, 98980, 98870, 98730, 
    98660, 98610, 98680, 98750, 98720, 98710, 98790, 98850, 98860, 98890, 
    98930, 98940, 98960, 99020, 99030, 99010, 99000, 98990, 98970, 98910, 
    98860, 98750, 98670, 98560, 98480, 98450, 98340, 98350, 98370, 98380, 
    98360, 98450, 98490, 98530, 98570, 98590, 98630, 98660, 98650, 98740, 
    98770, 98820, 98860, 98890, 98940, 98970, 98970, 98980, 99030, 99070, 
    99080, 99110, 99160, 99240, 99260, 99290, 99290, 99290, 99300, 99300, 
    99300, 99280, 99260, 99220, 99210, 99210, 99220, 99220, 99220, 99200, 
    99180, 99180, 99170, 99150, 99150, 99190, 99190, 99190, 99240, 99260, 
    99270, 99300, 99340, 99360, 99320, 99360, 99400, 99420, 99430, 99440, 
    99470, 99510, 99520, 99520, 99560, 99570, 99580, 99570, 99590, 99570, 
    99560, 99550, 99580, 99570, 99550, 99560, 99550, 99550, 99550, 99540, 
    99520, 99480, 99480, 99450, 99440, 99460, 99450, 99410, 99360, 99340, 
    99290, 99240, 99190, 99180, 99120, 99110, 99070, 99030, 99000, 98960, 
    98900, 98850, 98810, 98740, 98690, 98630, 98580, 98530, 98510, 98480, 
    98450, 98410, 98380, 98380, 98400, 98410, 98410, 98430, 98460, 98480, 
    98530, 98580, 98630, 98660, 98730, 98750, 98810, 98840, 98890, 98920, 
    98940, 98980, 99030, 99070, 99130, 99160, 99170, 99190, 99210, 99200, 
    99180, 99210, 99230, 99270, 99310, 99340, 99360, 99400, 99400, 99400, 
    99410, 99410, 99410, 99410, 99400, 99410, 99430, 99450, 99460, 99460, 
    99470, 99490, 99460, 99480, 99480, 99480, 99480, 99480, 99490, 99480, 
    99480, 99490, 99500, 99510, 99470, 99460, 99440, 99410, 99410, 99430, 
    99450, 99480, 99500, 99510, 99510, 99520, 99550, 99580, 99600, 99600, 
    99620, 99660, 99700, 99760, 99760, 99800, 99820, 99850, 99910, 99940, 
    99960, 99990, 100040, 100090, 100120, 100170, 100200, 100250, 100290, 
    100340, 100400, 100420, 100390, 100420, 100440, 100450, 100420, 100470, 
    100490, 100470, 100440, 100360, 100280, 100200, 100090, 99940, 99770, 
    99600, 99400, 99170, 98940, 98670, 98450, 98220, 98010, 97840, 97670, 
    97650, 97640, 97560, 97610, 97570, 97550, 97490, 97410, 97300, 97210, 
    97140, 97040, 96890, 96780, 96760, 96850, 96870, 96850, 96780, 96800, 
    96750, 96880, 96900, 96930, 97020, 97130, 97310, 97490, 97720, 97950, 
    98170, 98300, 98410, 98440, 98470, 98510, 98490, 98450, 98380, 98320, 
    98260, 98240, 98240, 98210, 98210, 98190, 98200, 98240, 98290, 98270, 
    98240, 98260, 98220, 98170, 98130, 98080, 98010, 97920, 97870, 97820, 
    97750, 97700, 97690, 97690, 97730, 97750, 97790, 97840, 97860, 97930, 
    98020, 98030, 98040, 98090, 98130, 98180, 98230, 98300, 98310, 98330, 
    98360, 98390, 98390, 98370, 98360, 98420, 98480, 98530, 98630, 98730, 
    98800, 98850, 98920, 98980, 99020, 99070, 99150, 99220, 99280, 99390, 
    99530, 99660, 99740, 99790, 99820, 99830, 99850, 99790, 99880, 99990, 
    100070, 100140, 100260, 100290, 100350, 100450, 100550, 100650, 100770, 
    100820, 100940, 101000, 101060, 101080, 101130, 101190, 101240, 101270, 
    101270, 101280, 101300, 101300, 101280, 101260, 101280, 101300, 101310, 
    101270, 101280, 101250, 101230, 101210, 101180, 101180, 101150, 101120, 
    101110, 101110, 101090, 101060, 101030, 101010, 100970, 100940, 100930, 
    100890, 100860, 100830, 100820, 100800, 100790, 100750, 100710, 100690, 
    100650, 100590, 100540, 100510, 100440, 100370, 100300, 100250, 100200, 
    100170, 100120, 100050, 99930, 99850, 99770, 99670, 99580, 99470, 99350, 
    99260, 99140, 98990, 98860, 98780, 98620, 98490, 98360, 98260, 98200, 
    98200, 98230, 98250, 98280, 98290, 98300, 98290, 98280, 98250, 98240, 
    98230, 98200, 98170, 98140, 98160, 98220, 98230, 98220, 98240, 98300, 
    98350, 98370, 98430, 98520, 98600, 98720, 98820, 98960, 99130, 99280, 
    99430, 99590, 99730, 99890, 100020, 100200, 100350, 100470, 100620, 
    100740, 100820, 100940, 101020, 101070, 101120, 101120, 101140, 101150, 
    101150, 101180, 101180, 101180, 101200, 101170, 101130, 101110, 101030, 
    101010, 100940, 100900, 100840, 100820, 100770, 100720, 100640, 100540, 
    100460, 100360, 100270, 100230, 100170, 100110, 100100, 100110, 100200, 
    100280, 100330, 100400, 100480, 100540, 100600, 100670, 100680, 100710, 
    100740, 100760, 100770, 100780, 100760, 100770, 100770, 100780, 100780, 
    100780, 100750, 100740, 100740, 100770, 100790, 100810, 100800, 100780, 
    100720, 100680, 100620, 100520, 100510, 100440, 100340, 100300, 100270, 
    100230, 100190, 100150, 100100, 100050, 99960, 99920, 99930, 99950, 
    99940, 99930, 99950, 99980, 99970, 99970, 99960, 99970, 100000, 100020, 
    100040, 100080, 100150, 100190, 100230, 100290, 100320, 100360, 100400, 
    100440, 100480, 100560, 100620, 100650, 100760, 100810, 100790, 100870, 
    100920, 100960, 100960, 100980, 101030, 101080, 101200, 101260, 101280, 
    101330, 101420, 101510, 101600, 101650, 101720, 101760, 101870, 101900, 
    101940, 101950, 102010, 102030, 102090, 102120, 102160, 102160, 102130, 
    102140, 102150, 102150, 102120, 102110, 102070, 102060, 102050, 102020, 
    101990, 101940, 101890, 101820, 101750, 101680, 101600, 101540, 101470, 
    101390, 101310, 101240, 101160, 101100, 101050, 100970, 100940, 100890, 
    100830, 100780, 100710, 100690, 100670, 100680, 100670, 100640, 100600, 
    100590, 100580, 100550, 100510, 100480, 100470, 100450, 100440, 100430, 
    100400, 100360, 100330, 100320, 100310, 100290, 100250, 100200, 100170, 
    100150, 100130, 100110, 100080, 100040, 100040, 100020, 99970, 99940, 
    99900, 99870, 99850, 99850, 99860, 99870, 99890, 99920, 99960, 100010, 
    100060, 100100, 100170, 100210, 100320, 100390, 100480, 100560, 100600, 
    100630, 100630, 100680, 100690, 100650, 100640, 100600, 100550, 100520, 
    100510, 100480, 100490, 100490, 100510, 100510, 100500, 100470, 100440, 
    100460, 100440, 100430, 100460, 100510, 100540, 100540, 100510, 100490, 
    100500, 100530, 100550, 100560, 100600, 100600, 100640, 100650, 100700, 
    100730, 100740, 100790, 100800, 100890, 100950, 100990, 101020, 101070, 
    101130, 101200, 101280, 101300, 101350, 101400, 101450, 101470, 101510, 
    101520, 101530, 101500, 101490, 101470, 101440, 101410, 101350, 101310, 
    101300, 101300, 101290, 101270, 101260, 101320, 101410, 101470, 101530, 
    101600, 101640, 101640, 101700, 101720, 101770, 101830, 101920, 102010, 
    102060, 102080, 102150, 102300, 102360, 102400, 102410, 102460, 102470, 
    102550, 102570, 102670, 102720, 102790, 102820, 102860, 102890, 102870, 
    102820, 102810, 102840, 102870, 102890, 102890, 102930, 102940, 102990, 
    103020, 103010, 103050, 103100, 103090, 103070, 103060, 103050, 103090, 
    103070, 103090, 103060, 103110, 103160, 103150, 103150, 103150, 103190, 
    103180, 103200, 103220, 103200, 103180, 103140, 103100, 103080, 103050, 
    103000, 102950, 102920, 102850, 102780, 102720, 102680, 102610, 102550, 
    102460, 102330, 102220, 102090, 101970, 101850, 101720, 101570, 101450, 
    101330, 101280, 101240, 101180, 101170, 101220, 101230, 101280, 101300, 
    101300, 101310, 101270, 101250, 101240, 101190, 101100, 101020, 100880, 
    100740, 100560, 100430, 100280, 100120, 100080, 99920, 99790, 99630, 
    99440, 99340, 99130, 98880, 98660, 98440, 98170, 97940, 97780, 97720, 
    97700, 97720, 97780, 97860, 98000, 98220, 98460, 98680, 98840, 98990, 
    99170, 99290, 99340, 99350, 99440, 99480, 99570, 99560, 99500, 99480, 
    99500, 99490, 99510, 99570, 99670, 99800, 99920, 100050, 100190, 100370, 
    100530, 100680, 100790, 100960, 101160, 101300, 101480, 101610, 101740, 
    101880, 102010, 102120, 102220, 102300, 102370, 102400, 102470, 102560, 
    102580, 102550, 102550, 102620, 102540, 102440, 102360, 102260, 102160, 
    102090, 101980, 101840, 101750, 101620, 101530, 101420, 101330, 101250, 
    101120, 101010, 100900, 100810, 100740, 100660, 100590, 100550, 100500, 
    100490, 100500, 100540, 100590, 100630, 100680, 100750, 100780, 100800, 
    100900, 100940, 101050, 101100, 101110, 101100, 101130, 101180, 101190, 
    101170, 101150, 101160, 101200, 101190, 101170, 101180, 101160, 101130, 
    101120, 101080, 101070, 101070, 101060, 101070, 101070, 101040, 101030, 
    101000, 100980, 100960, 100940, 100910, 100890, 100870, 100860, 100860, 
    100870, 100880, 100870, 100860, 100870, 100840, 100830, 100820, 100800, 
    100810, 100810, 100810, 100820, 100810, 100800, 100760, 100730, 100700, 
    100690, 100670, 100620, 100580, 100590, 100580, 100580, 100540, 100510, 
    100460, 100420, 100390, 100330, 100270, 100230, 100170, 100100, 100050, 
    99990, 99900, 99830, 99760, 99680, 99590, 99450, 99330, 99220, 99080, 
    98950, 98860, 98770, 98620, 98470, 98280, 98150, 98110, 98100, 98130, 
    98140, 98130, 98140, 98150, 98150, 98190, 98200, 98180, 98170, 98160, 
    98190, 98130, 98090, 98070, 98020, 97950, 97910, 97810, 97720, 97720, 
    97700, 97710, 97740, 97770, 97800, 97860, 97870, 97860, 97850, 97870, 
    97890, 97970, 97990, 98060, 98170, 98280, 98390, 98560, 98690, 98860, 
    99040, 99180, 99410, 99420, 99480, 99620, 99700, 99820, 99800, 99840, 
    99860, 99950, 100020, 100000, 99990, 99930, 99940, 99920, 99860, 99860, 
    99820, 99820, 99820, 99820, 99770, 99760, 99820, 99830, 99770, 99780, 
    99800, 99790, 99730, 99740, 99720, 99730, 99710, 99730, 99730, 99690, 
    99710, 99730, 99700, 99730, 99700, 99700, 99700, 99690, 99670, 99700, 
    99660, 99660, 99600, 99590, 99560, 99530, 99500, 99500, 99480, 99510, 
    99560, 99570, 99610, 99650, 99690, 99750, 99780, 99830, 99850, 99930, 
    99920, 99990, 100030, 100110, 100130, 100190, 100200, 100200, 100260, 
    100280, 100310, 100340, 100370, 100380, 100430, 100460, 100490, 100530, 
    100580, 100610, 100630, 100640, 100690, 100720, 100750, 100820, 100870, 
    100930, 100960, 100990, 101030, 101070, 101080, 101130, 101180, 101220, 
    101260, 101290, 101330, 101370, 101410, 101460, 101480, 101510, 101510, 
    101560, 101580, 101620, 101650, 101700, 101750, 101780, 101790, 101810, 
    101830, 101870, 101910, 101950, 101960, 102010, 102060, 102080, 102100, 
    102110, 102110, 102080, 102040, 102050, 102060, 102060, 102030, 101990, 
    101970, 101960, 101930, 101850, 101820, 101780, 101740, 101670, 101630, 
    101580, 101530, 101510, 101460, 101390, 101320, 101260, 101210, 101130, 
    101110, 101070, 101050, 101010, 100960, 100910, 100910, 100910, 100900, 
    100880, 100840, 100820, 100780, 100760, 100770, 100770, 100760, 100740, 
    100720, 100750, 100740, 100750, 100740, 100720, 100700, 100680, 100660, 
    100670, 100700, 100640, 100620, 100610, 100610, 100620, 100640, 100640, 
    100650, 100620, 100600, 100590, 100580, 100590, 100580, 100570, 100590, 
    100600, 100600, 100570, 100570, 100560, 100550, 100560, 100570, 100580, 
    100570, 100590, 100610, 100640, 100680, 100690, 100690, 100740, 100790, 
    100840, 100880, 100930, 100980, 101040, 101080, 101130, 101160, 101190, 
    101240, 101280, 101290, 101320, 101330, 101330, 101360, 101390, 101410, 
    101450, 101480, 101460, 101470, 101490, 101500, 101490, 101490, 101480, 
    101460, 101430, 101390, 101370, 101360, 101300, 101230, 101150, 101110, 
    101090, 101030, 100990, 100930, 100930, 100910, 100880, 100870, 100850, 
    100830, 100800, 100790, 100760, 100740, 100720, 100680, 100650, 100610, 
    100590, 100530, 100480, 100470, 100410, 100410, 100400, 100420, 100420, 
    100430, 100470, 100500, 100570, 100630, 100690, 100750, 100850, 100960, 
    101040, 101120, 101230, 101290, 101330, 101370, 101420, 101460, 101490, 
    101510, 101530, 101490, 101510, 101460, 101390, 101360, 101360, 101340, 
    101330, 101340, 101320, 101290, 101230, 101260, 101210, 101170, 101130, 
    101110, 101110, 101090, 101100, 101120, 101130, 101110, 101100, 101100, 
    101060, 101020, 100990, 100940, 100890, 100860, 100830, 100820, 100770, 
    100720, 100670, 100630, 100610, 100580, 100570, 100580, 100590, 100590, 
    100570, 100560, 100550, 100560, 100550, 100530, 100520, 100510, 100520, 
    100550, 100560, 100620, 100690, 100740, 100800, 100840, 100870, 100890, 
    100930, 100920, 100950, 100970, 101000, 101040, 101050, 101060, 101100, 
    101100, 101080, 101080, 101080, 101090, 101110, 101130, 101130, 101130, 
    101110, 101110, 101110, 101100, 101080, 101050, 101010, 100950, 100900, 
    100860, 100790, 100710, 100630, 100510, 100400, 100220, 100040, 99840, 
    99610, 99560, 99450, 99430, 99390, 99390, 99360, 99350, 99480, 99610, 
    99690, 99780, 99830, 99890, 99960, 100000, 100060, 100080, 100150, 
    100170, 100180, 100200, 100170, 100130, 100080, 100040, 99980, 99910, 
    99870, 99830, 99800, 99790, 99720, 99730, 99700, 99690, 99680, 99640, 
    99660, 99680, 99720, 99760, 99800, 99860, 99910, 100060, 100080, 100150, 
    100270, 100410, 100460, 100540, 100590, 100700, 100760, 100790, 100820, 
    100830, 100830, 100870, 100890, 100900, 100870, 100850, 100800, 100750, 
    100650, 100560, 100460, 100370, 100270, 100130, 100000, 99890, 99780, 
    99710, 99670, 99650, 99610, 99580, 99530, 99470, 99420, 99380, 99360, 
    99340, 99320, 99300, 99280, 99250, 99200, 99140, 99060, 98970, 98840, 
    98710, 98580, 98480, 98370, 98310, 98210, 98100, 98050, 97950, 97890, 
    97800, 97740, 97670, 97580, 97500, 97430, 97380, 97360, 97330, 97330, 
    97340, 97330, 97320, 97350, 97380, 97430, 97470, 97490, 97520, 97580, 
    97680, 97680, 97700, 97740, 97780, 97820, 97870, 97920, 97970, 98000, 
    98040, 98060, 98120, 98150, 98190, 98190, 98230, 98250, 98290, 98330, 
    98340, 98330, 98370, 98400, 98410, 98330, 98390, 98390, 98350, 98350, 
    98350, 98360, 98370, 98310, 98320, 98310, 98330, 98360, 98310, 98270, 
    98240, 98250, 98240, 98210, 98190, 98160, 98160, 98170, 98210, 98210, 
    98240, 98250, 98220, 98250, 98220, 98230, 98230, 98260, 98270, 98280, 
    98270, 98280, 98290, 98290, 98280, 98280, 98280, 98280, 98250, 98230, 
    98240, 98260, 98240, 98230, 98230, 98220, 98210, 98220, 98200, 98200, 
    98200, 98190, 98220, 98210, 98240, 98220, 98230, 98220, 98240, 98270, 
    98280, 98290, 98320, 98360, 98370, 98390, 98400, 98410, 98430, 98440, 
    98440, 98420, 98410, 98390, 98390, 98400, 98400, 98410, 98430, 98470, 
    98490, 98530, 98580, 98610, 98620, 98660, 98700, 98760, 98820, 98860, 
    98910, 98970, 99020, 99090, 99140, 99170, 99220, 99240, 99310, 99390, 
    99420, 99450, 99520, 99560, 99620, 99650, 99710, 99740, 99780, 99810, 
    99820, 99830, 99860, 99870, 99910, 99940, 99960, 99980, 99970, 99970, 
    99970, 100000, 100020, 100010, 100010, 100000, 100000, 100000, 99990, 
    99980, 99980, 99950, 99910, 99870, 99870, 99850, 99820, 99800, 99770, 
    99750, 99750, 99720, 99690, 99660, 99610, 99560, 99520, 99460, 99410, 
    99350, 99340, 99260, 99210, 99190, 99140, 99060, 99020, 99000, 99000, 
    99000, 99000, 99030, 99050, 99090, 99120, 99150, 99180, 99190, 99250, 
    99320, 99400, 99470, 99590, 99610, 99700, 99760, 99830, 99830, 99870, 
    99890, 99890, 99890, 99890, 99870, 99870, 99870, 99850, 99870, 99870, 
    99860, 99850, 99810, 99800, 99800, 99840, 99860, 99890, 99900, 99930, 
    99960, 100000, 100030, 100040, 100050, 100020, 100010, 99970, 99930, 
    99860, 99790, 99800, 99690, 99600, 99500, 99410, 99260, 99100, 98950, 
    98810, 98640, 98520, 98430, 98340, 98270, 98210, 98180, 98180, 98210, 
    98260, 98320, 98360, 98440, 98560, 98630, 98770, 98960, 99130, 99220, 
    99440, 99590, 99680, 99750, 99830, 99870, 99950, 100000, 100020, 100080, 
    100110, 100060, 100090, 100100, 100100, 100120, 100100, 100110, 100130, 
    100170, 100240, 100330, 100330, 100410, 100480, 100490, 100590, 100680, 
    100720, 100730, 100780, 100840, 100860, 100910, 100970, 101050, 101030, 
    101070, 101070, 101150, 101150, 101220, 101280, 101280, 101290, 101350, 
    101360, 101360, 101380, 101370, 101350, 101300, 101290, 101340, 101350, 
    101380, 101410, 101410, 101390, 101390, 101360, 101340, 101310, 101290, 
    101240, 101210, 101170, 101140, 101120, 101110, 101080, 101060, 101020, 
    100980, 100940, 100920, 100900, 100910, 100930, 100940, 100930, 100940, 
    100910, 100910, 100880, 100850, 100820, 100810, 100800, 100790, 100810, 
    100810, 100800, 100800, 100790, 100830, 100860, 100880, 100890, 100890, 
    100880, 100870, 100850, 100850, 100820, 100820, 100820, 100820, 100820, 
    100810, 100790, 100770, 100770, 100780, 100780, 100780, 100760, 100770, 
    100770, 100750, 100740, 100710, 100700, 100700, 100700, 100680, 100710, 
    100700, 100700, 100720, 100710, 100730, 100770, 100780, 100810, 100830, 
    100850, 100880, 100890, 100900, 100950, 100980, 101000, 101040, 101020, 
    101060, 101090, 101110, 101130, 101150, 101180, 101190, 101220, 101260, 
    101300, 101320, 101360, 101380, 101400, 101380, 101390, 101400, 101390, 
    101390, 101370, 101370, 101340, 101320, 101310, 101290, 101200, 101100, 
    101070, 101030, 100990, 100930, 100840, 100770, 100720, 100670, 100630, 
    100560, 100490, 100400, 100330, 100290, 100230, 100190, 100160, 100120, 
    100080, 100070, 100030, 100000, 100040, 100020, 100020, 100010, 100080, 
    100110, 100200, 100290, 100330, 100390, 100420, 100460, 100500, 100520, 
    100520, 100540, 100560, 100570, 100560, 100590, 100610, 100590, 100580, 
    100590, 100580, 100590, 100600, 100630, 100650, 100650, 100670, 100690, 
    100670, 100660, 100640, 100640, 100630, 100630, 100660, 100650, 100640, 
    100660, 100680, 100740, 100790, 100810, 100840, 100880, 100910, 100930, 
    100910, 100890, 100870, 100880, 100890, 100890, 100890, 100900, 100880, 
    100880, 100880, 100870, 100880, 100890, 100920, 100920, 100990, 101000, 
    101000, 101010, 101040, 101060, 101080, 101120, 101140, 101170, 101220, 
    101190, 101200, 101210, 101210, 101240, 101260, 101270, 101290, 101310, 
    101330, 101370, 101390, 101410, 101430, 101440, 101430, 101440, 101460, 
    101450, 101460, 101480, 101490, 101510, 101500, 101520, 101530, 101520, 
    101510, 101510, 101470, 101440, 101430, 101420, 101390, 101380, 101380, 
    101380, 101370, 101380, 101380, 101360, 101350, 101300, 101270, 101250, 
    101210, 101200, 101170, 101150, 101160, 101140, 101100, 101050, 101010, 
    100980, 100960, 100960, 100980, 100970, 100980, 100990, 100980, 100960, 
    100960, 100920, 100910, 100890, 100850, 100820, 100810, 100760, 100750, 
    100740, 100710, 100700, 100670, 100660, 100670, 100660, 100680, 100700, 
    100720, 100770, 100800, 100800, 100800, 100810, 100860, 100880, 100900, 
    100920, 100950, 100970, 101010, 101030, 101060, 101090, 101130, 101160, 
    101180, 101200, 101250, 101280, 101320, 101320, 101370, 101400, 101440, 
    101470, 101510, 101540, 101580, 101600, 101630, 101660, 101690, 101680, 
    101710, 101730, 101760, 101810, 101840, 101840, 101860, 101890, 101910, 
    101940, 101940, 101950, 101970, 102010, 102060, 102080, 102100, 102120, 
    102140, 102150, 102150, 102170, 102170, 102170, 102180, 102170, 102180, 
    102210, 102220, 102220, 102220, 102220, 102230, 102210, 102190, 102170, 
    102160, 102170, 102160, 102160, 102170, 102160, 102150, 102140, 102120, 
    102110, 102070, 102050, 102020, 101990, 101990, 101970, 101940, 101890, 
    101850, 101800, 101750, 101710, 101680, 101690, 101760, 101830, 101910, 
    101950, 102000, 102030, 102060, 102100, 102180, 102190, 102230, 102220, 
    102230, 102250, 102260, 102270, 102280, 102290, 102310, 102300, 102310, 
    102340, 102350, 102380, 102360, 102350, 102340, 102350, 102340, 102350, 
    102370, 102330, 102310, 102310, 102290, 102280, 102250, 102280, 102280, 
    102290, 102290, 102310, 102300, 102270, 102270, 102270, 102250, 102250, 
    102240, 102220, 102220, 102200, 102180, 102170, 102150, 102160, 102160, 
    102140, 102150, 102130, 102130, 102130, 102120, 102120, 102110, 102110, 
    102090, 102080, 102070, 102070, 102060, 102050, 102020, 101980, 101980, 
    101950, 101940, 101930, 101890, 101880, 101860, 101840, 101840, 101810, 
    101790, 101780, 101770, 101780, 101780, 101770, 101750, 101750, 101760, 
    101790, 101790, 101760, 101760, 101780, 101790, 101800, 101800, 101810, 
    101840, 101830, 101810, 101810, 101810, 101790, 101790, 101780, 101790, 
    101780, 101760, 101780, 101770, 101770, 101760, 101740, 101710, 101670, 
    101640, 101620, 101620, 101620, 101610, 101590, 101580, 101580, 101560, 
    101540, 101510, 101480, 101460, 101440, 101430, 101410, 101390, 101370, 
    101370, 101350, 101310, 101280, 101260, 101220, 101210, 101200, 101190, 
    101210, 101230, 101230, 101220, 101180, 101180, 101160, 101110, 101100, 
    101120, 101130, 101170, 101210, 101240, 101240, 101240, 101240, 101200, 
    101200, 101180, 101130, 101120, 101130, 101090, 101130, 101130, 101110, 
    101100, 101090, 101100, 101110, 101100, 101140, 101220, 101270, 101310, 
    101280, 101380, 101400, 101410, 101450, 101460, 101470, 101520, 101530, 
    101540, 101560, 101580, 101610, 101650, 101660, 101650, 101670, 101670, 
    101660, 101640, 101640, 101650, 101670, 101680, 101690, 101700, 101710, 
    101700, 101680, 101660, 101670, 101650, 101630, 101590, 101600, 101630, 
    101650, 101680, 101660, 101650, 101640, 101620, 101610, 101600, 101650, 
    101640, 101660, 101680, 101700, 101720, 101720, 101730, 101700, 101710, 
    101690, 101670, 101660, 101670, 101660, 101660, 101660, 101660, 101680, 
    101650, 101640, 101630, 101610, 101600, 101600, 101600, 101590, 101600, 
    101610, 101590, 101580, 101560, 101530, 101500, 101490, 101470, 101440, 
    101430, 101420, 101410, 101400, 101380, 101380, 101380, 101360, 101360, 
    101370, 101360, 101350, 101340, 101350, 101360, 101370, 101380, 101380, 
    101400, 101410, 101430, 101430, 101450, 101440, 101440, 101460, 101470, 
    101490, 101500, 101510, 101510, 101500, 101500, 101480, 101470, 101440, 
    101420, 101400, 101380, 101320, 101240, 101160, 101110, 101050, 101000, 
    100970, 100920, 100890, 100870, 100850, 100860, 100880, 100890, 100870, 
    100890, 100910, 100910, 100910, 100910, 100880, 100870, 100850, 100850, 
    100830, 100810, 100780, 100730, 100690, 100640, 100570, 100530, 100460, 
    100420, 100390, 100370, 100360, 100390, 100450, 100550, 100630, 100740, 
    100790, 100860, 100850, 100900, 100910, 100930, 100950, 100950, 100940, 
    100930, 100970, 100970, 101040, 101080, 101120, 101170, 101210, 101240, 
    101280, 101330, 101360, 101450, 101500, 101590, 101690, 101800, 101930, 
    102050, 102160, 102240, 102370, 102460, 102530, 102570, 102630, 102700, 
    102710, 102730, 102740, 102750, 102780, 102790, 102830, 102870, 102870, 
    102890, 102900, 102890, 102860, 102820, 102780, 102770, 102760, 102740, 
    102710, 102690, 102670, 102630, 102560, 102530, 102510, 102490, 102410, 
    102330, 102270, 102230, 102190, 102180, 102130, 102090, 102050, 102030, 
    102000, 101960, 101940, 101900, 101880, 101870, 101870, 101890, 101890, 
    101890, 101880, 101900, 101880, 101910, 101940, 101970, 102020, 102080, 
    102120, 102170, 102230, 102290, 102340, 102390, 102440, 102450, 102470, 
    102510, 102530, 102550, 102560, 102570, 102570, 102560, 102570, 102580, 
    102580, 102550, 102510, 102470, 102420, 102390, 102300, 102250, 102150, 
    102030, 101900, 101770, 101650, 101560, 101460, 101390, 101330, 101240, 
    101200, 101120, 101100, 101040, 101000, 100990, 100950, 100930, 100870, 
    100890, 100880, 100880, 100860, 100860, 100880, 100820, 100860, 100920, 
    100970, 101000, 101040, 101110, 101190, 101210, 101320, 101420, 101480, 
    101540, 101630, 101680, 101760, 101860, 101910, 101980, 102030, 102120, 
    102200, 102300, 102370, 102420, 102480, 102550, 102590, 102630, 102630, 
    102660, 102670, 102680, 102710, 102710, 102730, 102730, 102740, 102730, 
    102710, 102700, 102660, 102640, 102630, 102620, 102620, 102630, 102680, 
    102630, 102720, 102750, 102780, 102770, 102780, 102830, 102830, 102830, 
    102850, 102890, 102880, 102860, 102900, 102880, 102880, 102900, 102910, 
    102920, 102900, 102910, 102930, 102950, 102970, 102980, 102970, 102970, 
    102980, 102970, 102960, 102990, 103000, 103050, 103040, 103060, 103060, 
    103080, 103090, 103070, 103080, 103080, 103090, 103100, 103110, 103090, 
    103130, 103130, 103140, 103140, 103170, 103150, 103130, 103130, 103110, 
    103080, 103070, 103060, 103060, 103040, 103020, 103020, 102990, 102960, 
    102950, 102940, 102920, 102890, 102900, 102920, 102930, 102940, 102960, 
    102980, 103020, 103040, 103070, 103090, 103120, 103160, 103190, 103240, 
    103260, 103290, 103300, 103320, 103320, 103300, 103290, 103280, 103250, 
    103320, 103200, 103190, 103170, 103180, 103150, 103120, 103090, 103080, 
    103050, 103020, 102990, 102960, 102930, 102920, 102930, 102920, 102890, 
    102860, 102850, 102820, 102800, 102780, 102750, 102710, 102710, 102710, 
    102720, 102730, 102720, 102720, 102710, 102700, 102700, 102690, 102680, 
    102700, 102700, 102710, 102720, 102720, 102740, 102750, 102750, 102750, 
    102770, 102760, 102750, 102740, 102760, 102760, 102760, 102780, 102790, 
    102800, 102800, 102790, 102790, 102780, 102770, 102760, 102760, 102770, 
    102780, 102800, 102800, 102800, 102800, 102800, 102820, 102800, 102790, 
    102790, 102800, 102820, 102840, 102840, 102850, 102870, 102890, 102900, 
    102900, 102920, 102920, 102920, 102920, 102930, 102930, 102950, 102960, 
    102950, 102930, 102930, 102940, 102940, 102940, 102930, 102920, 102910, 
    102890, 102870, 102850, 102830, 102770, 102730, 102670, 102600, 102540, 
    102440, 102300, 102230, 102130, 102060, 101980, 101910, 101780, 101680, 
    101560, 101540, 101520, 101510, 101480, 101460, 101450, 101450, 101490, 
    101490, 101530, 101540, 101570, 101600, 101640, 101660, 101690, 101710, 
    101740, 101760, 101780, 101800, 101810, 101820, 101840, 101840, 101820, 
    101810, 101820, 101830, 101840, 101880, 101880, 101880, 101890, 101880, 
    101870, 101890, 101890, 101880, 101890, 101900, 101920, 101950, 101940, 
    101960, 101970, 101980, 101960, 101980, 101970, 101980, 101980, 101990, 
    101990, 102010, 102020, 102030, 102040, 102040, 102030, 102010, 102000, 
    102000, 102000, 101980, 101970, 101970, 101960, 101950, 101940, 101920, 
    101900, 101880, 101860, 101860, 101850, 101840, 101840, 101840, 101850, 
    101860, 101870, 101870, 101870, 101860, 101840, 101820, 101800, 101800, 
    101810, 101810, 101820, 101810, 101790, 101790, 101790, 101800, 101790, 
    101780, 101790, 101810, 101830, 101850, 101860, 101850, 101840, 101860, 
    101860, 101850, 101830, 101820, 101810, 101810, 101810, 101810, 101820, 
    101790, 101780, 101770, 101720, 101710, 101680, 101650, 101630, 101630, 
    101620, 101640, 101630, 101620, 101590, 101580, 101530, 101500, 101490, 
    101470, 101440, 101420, 101400, 101370, 101380, 101350, 101340, 101320, 
    101310, 101270, 101230, 101190, 101160, 101150, 101110, 101070, 101050, 
    101020, 100950, 100910, 100850, 100800, 100760, 100700, 100660, 100640, 
    100640, 100640, 100660, 100670, 100650, 100640, 100660, 100650, 100660, 
    100690, 100680, 100680, 100710, 100750, 100750, 100740, 100760, 100780, 
    100790, 100800, 100800, 100810, 100830, 100880, 100870, 100900, 100900, 
    100910, 100930, 100930, 100930, 100920, 100920, 100920, 100900, 100920, 
    100950, 100960, 100950, 100980, 100960, 100960, 100950, 100950, 100950, 
    100980, 100980, 100970, 100960, 100960, 100990, 101000, 101010, 101020, 
    101020, 101010, 101030, 101030, 101030, 101050, 101060, 101080, 101090, 
    101100, 101120, 101130, 101150, 101160, 101180, 101190, 101210, 101210, 
    101220, 101230, 101240, 101240, 101260, 101270, 101290, 101300, 101310, 
    101330, 101340, 101380, 101410, 101430, 101450, 101470, 101490, 101510, 
    101530, 101530, 101540, 101540, 101550, 101550, 101560, 101570, 101580, 
    101590, 101590, 101610, 101590, 101580, 101570, 101570, 101550, 101550, 
    101540, 101550, 101540, 101520, 101500, 101510, 101520, 101530, 101510, 
    101500, 101510, 101530, 101570, 101570, 101610, 101650, 101690, 101720, 
    101760, 101780, 101780, 101800, 101830, 101870, 101890, 101920, 101930, 
    101980, 102000, 102010, 102010, 102020, 102010, 102010, 102020, 102010, 
    102010, 102010, 102030, 102030, 102030, 102010, 102020, 102000, 101980, 
    101950, 101950, 101950, 101960, 101970, 101980, 101990, 102000, 102010, 
    102000, 102000, 102000, 101990, 101980, 101990, 102010, 102000, 101970, 
    101940, 101890, 101830, 101790, 101760, 101690, 101640, 101600, 101520, 
    101490, 101440, 101370, 101330, 101280, 101180, 101090, 101130, 101050, 
    101000, 100950, 100980, 100970, 100980, 100980, 100980, 101010, 101020, 
    101090, 101100, 101130, 101160, 101210, 101240, 101270, 101300, 101260, 
    101240, 101260, 101250, 101250, 101360, 101380, 101390, 101360, 101470, 
    101530, 101550, 101620, 101630, 101660, 101690, 101750, 101770, 101760, 
    101780, 101810, 101790, 101800, 101790, 101790, 101790, 101780, 101780, 
    101790, 101810, 101820, 101880, 101910, 101910, 101950, 101990, 102020, 
    102110, 102190, 102240, 102250, 102290, 102340, 102360, 102430, 102480, 
    102500, 102550, 102590, 102620, 102650, 102680, 102690, 102740, 102770, 
    102790, 102830, 102860, 102870, 102880, 102890, 102890, 102880, 102880, 
    102900, 102900, 102890, 102890, 102870, 102880, 102870, 102860, 102840, 
    102840, 102830, 102800, 102800, 102770, 102740, 102700, 102670, 102640, 
    102610, 102580, 102560, 102520, 102470, 102440, 102420, 102380, 102340, 
    102310, 102290, 102290, 102280, 102250, 102230, 102220, 102210, 102220, 
    102210, 102200, 102200, 102200, 102190, 102180, 102170, 102190, 102200, 
    102190, 102210, 102210, 102220, 102240, 102250, 102250, 102270, 102260, 
    102270, 102290, 102320, 102310, 102290, 102290, 102310, 102310, 102310, 
    102300, 102280, 102280, 102250, 102260, 102230, 102200, 102190, 102190, 
    102160, 102140, 102130, 102080, 102060, 102030, 102030, 102010, 101970, 
    101920, 101900, 101870, 101850, 101830, 101800, 101780, 101770, 101750, 
    101690, 101680, 101650, 101630, 101620, 101590, 101560, 101550, 101530, 
    101510, 101530, 101500, 101520, 101520, 101500, 101550, 101580, 101580, 
    101600, 101630, 101660, 101670, 101690, 101720, 101760, 101800, 101810, 
    101850, 101880, 101890, 101920, 101940, 101930, 101920, 101930, 101940, 
    101950, 101950, 101920, 101910, 101930, 101950, 101960, 101980, 101990, 
    102030, 102050, 102080, 102100, 102140, 102150, 102170, 102200, 102240, 
    102290, 102290, 102300, 102320, 102370, 102380, 102430, 102460, 102490, 
    102500, 102520, 102550, 102570, 102600, 102610, 102610, 102610, 102610, 
    102640, 102670, 102690, 102710, 102720, 102740, 102750, 102770, 102770, 
    102770, 102790, 102790, 102800, 102820, 102780, 102780, 102790, 102780, 
    102780, 102780, 102760, 102730, 102700, 102690, 102690, 102660, 102640, 
    102600, 102600, 102600, 102590, 102570, 102570, 102550, 102550, 102550, 
    102550, 102550, 102530, 102520, 102520, 102520, 102510, 102500, 102470, 
    102420, 102370, 102330, 102320, 102280, 102250, 102200, 102160, 102110, 
    102090, 102050, 102000, 101950, 101890, 101850, 101810, 101780, 101760, 
    101740, 101700, 101670, 101630, 101600, 101560, 101520, 101490, 101450, 
    101430, 101390, 101370, 101340, 101320, 101300, 101270, 101210, 101170, 
    101130, 101090, 101060, 101040, 101020, 101010, 100990, 100970, 100970, 
    100950, 100930, 100920, 100890, 100870, 100860, 100840, 100820, 100810, 
    100800, 100790, 100750, 100740, 100730, 100730, 100700, 100670, 100650, 
    100660, 100660, 100650, 100620, 100610, 100610, 100590, 100570, 100540, 
    100490, 100470, 100440, 100420, 100400, 100370, 100320, 100300, 100270, 
    100250, 100220, 100180, 100150, 100110, 100090, 100090, 100060, 100050, 
    100060, 100050, 100020, 100020, 100020, 100030, 100040, 100040, 100050, 
    100040, 100050, 100050, 100060, 100050, 100050, 100050, 100050, 100030, 
    100010, 100000, 100000, 99990, 100010, 100020, 100030, 100030, 100010, 
    100010, 100000, 99980, 99980, 99950, 99960, 99960, 99970, 99970, 99980, 
    100000, 100020, 100050, 100080, 100090, 100120, 100140, 100190, 100240, 
    100270, 100310, 100350, 100400, 100430, 100440, 100470, 100500, 100530, 
    100560, 100590, 100620, 100660, 100680, 100700, 100730, 100740, 100760, 
    100770, 100750, 100770, 100770, 100780, 100770, 100770, 100790, 100790, 
    100790, 100790, 100780, 100750, 100730, 100710, 100700, 100680, 100660, 
    100670, 100650, 100660, 100660, 100660, 100630, 100600, 100580, 100560, 
    100560, 100580, 100590, 100600, 100600, 100620, 100610, 100620, 100620, 
    100630, 100610, 100600, 100600, 100600, 100610, 100610, 100620, 100620, 
    100630, 100620, 100610, 100590, 100580, 100560, 100550, 100570, 100560, 
    100560, 100590, 100590, 100570, 100560, 100560, 100540, 100540, 100540, 
    100530, 100520, 100510, 100510, 100500, 100500, 100490, 100520, 100530, 
    100540, 100550, 100550, 100570, 100600, 100660, 100690, 100710, 100710, 
    100730, 100730, 100750, 100770, 100810, 100810, 100830, 100850, 100860, 
    100870, 100890, 100910, 100900, 100920, 100920, 100940, 100940, 100950, 
    100970, 100980, 101000, 101020, 101000, 101010, 101030, 101050, 101040, 
    101040, 101030, 101040, 101050, 101050, 101050, 101050, 101040, 101070, 
    101070, 101070, 101070, 101060, 101060, 101070, 101080, 101090, 101070, 
    101060, 101050, 101050, 101060, 101050, 101030, 101020, 101010, 100990, 
    100980, 100980, 100980, 100980, 100980, 100970, 100980, 101000, 101000, 
    101000, 100990, 101000, 101000, 100990, 101010, 101020, 101030, 101020, 
    101020, 101000, 101010, 101010, 100990, 100970, 100960, 100930, 100900, 
    100890, 100900, 100910, 100900, 100900, 100900, 100870, 100860, 100850, 
    100860, 100860, 100850, 100870, 100870, 100860, 100860, 100860, 100860, 
    100860, 100860, 100840, 100820, 100830, 100840, 100840, 100840, 100860, 
    100860, 100860, 100860, 100830, 100820, 100810, 100810, 100800, 100780, 
    100800, 100800, 100800, 100780, 100770, 100730, 100730, 100730, 100720, 
    100700, 100680, 100680, 100650, 100630, 100620, 100590, 100570, 100550, 
    100510, 100480, 100440, 100410, 100390, 100370, 100360, 100340, 100320, 
    100300, 100260, 100240, 100230, 100200, 100190, 100170, 100170, 100170, 
    100160, 100150, 100140, 100130, 100110, 100110, 100110, 100100, 100110, 
    100100, 100100, 100100, 100120, 100120, 100120, 100130, 100120, 100110, 
    100110, 100130, 100130, 100100, 100090, 100080, 100090, 100070, 100050, 
    100040, 100010, 99990, 99940, 99930, 99900, 99870, 99860, 99860, 99840, 
    99810, 99780, 99780, 99760, 99730, 99700, 99710, 99700, 99720, 99730, 
    99750, 99760, 99810, 99830, 99850, 99890, 99930, 99960, 99990, 100030, 
    100080, 100110, 100160, 100220, 100260, 100300, 100350, 100400, 100470, 
    100530, 100590, 100650, 100720, 100780, 100860, 100930, 100990, 101060, 
    101110, 101170, 101210, 101240, 101260, 101300, 101330, 101350, 101400, 
    101430, 101460, 101480, 101500, 101510, 101530, 101560, 101580, 101570, 
    101590, 101640, 101660, 101680, 101690, 101690, 101710, 101690, 101680, 
    101670, 101640, 101630, 101620, 101590, 101580, 101590, 101570, 101550, 
    101530, 101500, 101480, 101440, 101410, 101380, 101360, 101360, 101340, 
    101350, 101350, 101340, 101330, 101300, 101290, 101270, 101260, 101240, 
    101240, 101230, 101240, 101250, 101220, 101220, 101220, 101220, 101220, 
    101210, 101210, 101190, 101190, 101190, 101180, 101200, 101210, 101210, 
    101210, 101210, 101200, 101160, 101130, 101100, 101070, 101060, 101040, 
    101030, 101050, 101040, 101040, 100990, 100940, 100920, 100850, 100840, 
    100800, 100750, 100720, 100700, 100630, 100570, 100550, 100510, 100480, 
    100450, 100410, 100370, 100330, 100320, 100290, 100260, 100250, 100210, 
    100190, 100160, 100140, 100100, 100060, 100040, 100020, 100010, 100020, 
    100020, 100020, 100020, 100010, 100010, 99990, 100010, 100020, 100020, 
    100030, 100050, 100080, 100110, 100150, 100170, 100200, 100220, 100250, 
    100290, 100300, 100320, 100350, 100370, 100410, 100440, 100500, 100570, 
    100590, 100600, 100630, 100650, 100660, 100660, 100690, 100690, 100730, 
    100770, 100810, 100840, 100860, 100850, 100870, 100860, 100850, 100860, 
    100850, 100840, 100860, 100870, 100880, 100880, 100880, 100860, 100830, 
    100810, 100800, 100780, 100770, 100760, 100730, 100710, 100690, 100670, 
    100630, 100580, 100560, 100530, 100490, 100440, 100410, 100370, 100330, 
    100290, 100280, 100250, 100210, 100170, 100130, 100110, 100090, 100050, 
    100030, 100010, 99990, 100000, 100010, 100020, 100030, 100000, 100010, 
    99990, 100000, 100010, 100020, 100040, 100060, 100090, 100140, 100160, 
    100210, 100240, 100260, 100280, 100300, 100320, 100340, 100350, 100380, 
    100390, 100400, 100410, 100420, 100410, 100420, 100420, 100410, 100440, 
    100450, 100490, 100520, 100540, 100580, 100620, 100630, 100650, 100670, 
    100660, 100680, 100710, 100730, 100750, 100780, 100790, 100800, 100800, 
    100800, 100800, 100810, 100810, 100820, 100810, 100810, 100810, 100810, 
    100820, 100820, 100820, 100810, 100800, 100780, 100770, 100770, 100750, 
    100730, 100720, 100700, 100680, 100670, 100670, 100680, 100670, 100640, 
    100630, 100620, 100610, 100610, 100610, 100610, 100610, 100620, 100610, 
    100600, 100590, 100590, 100570, 100570, 100550, 100560, 100560, 100580, 
    100570, 100570, 100560, 100560, 100570, 100570, 100580, 100590, 100600, 
    100610, 100610, 100630, 100610, 100620, 100600, 100600, 100590, 100560, 
    100530, 100510, 100490, 100470, 100440, 100400, 100380, 100320, 100280, 
    100260, 100230, 100180, 100150, 100120, 100090, 100040, 100030, 100000, 
    99970, 99960, 99960, 99960, 99970, 99970, 99960, 99950, 99910, 99900, 
    99980, 100050, 100120, 100190, 100250, 100290, 100370, 100450, 100490, 
    100590, 100660, 100760, 100860, 100930, 101010, 101060, 101070, 101080, 
    101130, 101140, 101180, 101210, 101240, 101260, 101270, 101280, 101310, 
    101320, 101320, 101300, 101280, 101250, 101260, 101250, 101220, 101170, 
    101140, 101100, 101120, 101060, 101030, 100940, 100880, 100820, 100740, 
    100690, 100620, 100490, 100390, 100330, 100270, 100210, 100150, 100090, 
    100000, 99940, 99920, 99890, 99890, 99900, 99900, 99890, 99930, 99960, 
    99980, 99980, 99990, 99980, 99970, 99930, 99890, 99920, 99900, 99940, 
    99960, 100010, 100030, 100080, 100150, 100160, 100180, 100240, 100310, 
    100380, 100450, 100470, 100520, 100600, 100650, 100680, 100720, 100750, 
    100750, 100810, 100860, 100850, 100880, 100920, 100930, 100950, 100960, 
    100970, 100950, 100970, 100930, 100880, 100860, 100840, 100820, 100800, 
    100810, 100800, 100780, 100730, 100720, 100690, 100670, 100680, 100660, 
    100670, 100650, 100650, 100650, 100650, 100670, 100690, 100720, 100720, 
    100740, 100760, 100800, 100840, 100870, 100910, 100940, 100980, 100990, 
    101000, 101000, 101010, 101030, 101000, 100990, 100960, 100910, 100850, 
    100800, 100730, 100660, 100600, 100550, 100490, 100480, 100500, 100520, 
    100530, 100550, 100560, 100580, 100620, 100640, 100690, 100730, 100780, 
    100790, 100810, 100840, 100880, 100930, 101000, 101050, 101110, 101170, 
    101250, 101320, 101360, 101400, 101420, 101450, 101490, 101540, 101590, 
    101650, 101700, 101720, 101750, 101780, 101800, 101820, 101850, 101860, 
    101860, 101840, 101830, 101850, 101850, 101860, 101880, 101850, 101810, 
    101750, 101700, 101660, 101610, 101570, 101540, 101460, 101440, 101410, 
    101390, 101410, 101460, 101500, 101540, 101560, 101620, 101660, 101680, 
    101710, 101720, 101780, 101850, 101860, 101850, 101820, 101830, 101840, 
    101850, 101850, 101840, 101840, 101830, 101830, 101820, 101830, 101800, 
    101800, 101790, 101760, 101750, 101740, 101720, 101710, 101680, 101650, 
    101630, 101590, 101540, 101470, 101440, 101420, 101360, 101350, 101340, 
    101320, 101290, 101240, 101220, 101210, 101210, 101200, 101180, 101170, 
    101160, 101180, 101200, 101220, 101240, 101270, 101280, 101270, 101270, 
    101270, 101280, 101300, 101310, 101330, 101350, 101360, 101390, 101410, 
    101420, 101420, 101420, 101410, 101400, 101390, 101380, 101360, 101330, 
    101300, 101290, 101280, 101240, 101200, 101180, 101140, 101110, 101060, 
    101030, 101010, 100980, 100970, 100930, 100890, 100870, 100840, 100790, 
    100750, 100740, 100720, 100710, 100680, 100650, 100610, 100590, 100580, 
    100560, 100550, 100550, 100520, 100490, 100480, 100480, 100450, 100450, 
    100440, 100440, 100420, 100410, 100400, 100390, 100380, 100370, 100400, 
    100420, 100450, 100490, 100510, 100550, 100590, 100630, 100680, 100710, 
    100750, 100790, 100800, 100890, 100910, 100930, 100960, 101020, 101050, 
    101060, 101080, 101090, 101120, 101120, 101140, 101160, 101160, 101180, 
    101210, 101220, 101240, 101240, 101260, 101280, 101260, 101270, 101280, 
    101270, 101280, 101310, 101330, 101350, 101350, 101370, 101350, 101330, 
    101310, 101320, 101300, 101300, 101300, 101300, 101340, 101340, 101330, 
    101330, 101310, 101320, 101310, 101290, 101290, 101310, 101320, 101310, 
    101320, 101330, 101300, 101290, 101260, 101220, 101200, 101180, 101150, 
    101140, 101140, 101110, 101100, 101060, 101050, 101030, 101010, 100980, 
    100960, 100930, 100940, 100930, 100950, 100960, 100970, 100970, 100960, 
    100940, 100910, 100880, 100880, 100860, 100830, 100800, 100840, 100840, 
    100810, 100790, 100780, 100780, 100780, 100750, 100720, 100710, 100700, 
    100720, 100700, 100730, 100730, 100760, 100760, 100760, 100770, 100770, 
    100780, 100790, 100790, 100800, 100800, 100840, 100850, 100880, 100880, 
    100870, 100870, 100860, 100870, 100860, 100880, 100880, 100910, 100920, 
    100920, 100950, 101000, 100980, 100960, 100970, 100980, 100970, 100960, 
    100950, 100960, 100970, 100970, 100970, 100980, 100980, 100960, 100950, 
    100920, 100890, 100900, 100900, 100910, 100920, 100930, 100940, 100940, 
    100950, 100960, 100960, 100970, 100970, 100970, 100980, 100980, 100970, 
    100980, 101000, 101010, 101010, 101010, 101000, 101000, 100980, 100980, 
    100980, 101000, 101020, 101030, 101050, 101060, 101070, 101070, 101090, 
    101090, 101090, 101100, 101110, 101130, 101140, 101150, 101190, 101220, 
    101240, 101270, 101280, 101290, 101280, 101280, 101290, 101310, 101320, 
    101320, 101330, 101340, 101350, 101360, 101340, 101340, 101340, 101340, 
    101350, 101380, 101400, 101410, 101430, 101450, 101450, 101460, 101450, 
    101430, 101440, 101430, 101420, 101420, 101430, 101440, 101460, 101450, 
    101450, 101450, 101460, 101450, 101430, 101420, 101420, 101410, 101420, 
    101420, 101430, 101430, 101430, 101430, 101420, 101420, 101410, 101410, 
    101400, 101430, 101430, 101450, 101460, 101480, 101510, 101520, 101530, 
    101530, 101530, 101530, 101550, 101570, 101590, 101600, 101640, 101670, 
    101690, 101710, 101740, 101750, 101760, 101760, 101760, 101780, 101810, 
    101850, 101870, 101890, 101920, 101940, 101940, 101950, 101940, 101940, 
    101940, 101960, 101970, 101970, 101980, 101980, 101980, 101970, 101950, 
    101930, 101900, 101860, 101840, 101820, 101830, 101800, 101780, 101750, 
    101700, 101680, 101650, 101600, 101570, 101540, 101530, 101530, 101520, 
    101520, 101520, 101500, 101510, 101500, 101480, 101470, 101450, 101440, 
    101430, 101400, 101400, 101380, 101370, 101370, 101350, 101340, 101310, 
    101290, 101270, 101240, 101220, 101200, 101200, 101200, 101180, 101170, 
    101140, 101090, 101060, 101040, 101010, 101000, 100990, 101000, 100970, 
    100960, 100930, 100910, 100860, 100800, 100760, 100710, 100660, 100620, 
    100570, 100530, 100490, 100490, 100460, 100430, 100390, 100350, 100360, 
    100360, 100320, 100290, 100260, 100230, 100180, 100180, 100170, 100140, 
    100120, 100100, 100080, 100070, 100060, 100060, 100030, 100030, 100010, 
    99980, 99960, 99940, 99910, 99870, 99850, 99820, 99810, 99780, 99770, 
    99750, 99720, 99700, 99680, 99650, 99630, 99610, 99560, 99520, 99490, 
    99430, 99400, 99370, 99360, 99330, 99310, 99290, 99260, 99250, 99240, 
    99230, 99220, 99200, 99180, 99180, 99180, 99180, 99200, 99200, 99210, 
    99230, 99240, 99250, 99270, 99300, 99320, 99340, 99360, 99380, 99410, 
    99460, 99480, 99490, 99490, 99470, 99460, 99480, 99470, 99470, 99460, 
    99450, 99450, 99450, 99420, 99390, 99390, 99380, 99370, 99340, 99350, 
    99380, 99370, 99380, 99380, 99420, 99500, 99600, 99730, 99850, 100010, 
    100130, 100230, 100350, 100440, 100540, 100650, 100740, 100780, 100820, 
    100820, 100860, 100870, 100880, 100880, 100900, 100900, 100930, 100940, 
    100960, 100970, 101010, 101040, 101060, 101090, 101110, 101130, 101160, 
    101170, 101200, 101230, 101230, 101250, 101270, 101280, 101300, 101300, 
    101290, 101310, 101350, 101360, 101390, 101410, 101410, 101400, 101380, 
    101370, 101370, 101370, 101360, 101370, 101370, 101380, 101390, 101380, 
    101370, 101390, 101370, 101360, 101360, 101340, 101330, 101330, 101330, 
    101330, 101310, 101300, 101280, 101240, 101220, 101160, 101150, 101130, 
    101100, 101100, 101100, 101080, 101080, 101060, 101060, 101050, 101040, 
    101000, 100960, 100920, 100910, 100900, 100900, 100900, 100900, 100870, 
    100870, 100850, 100850, 100810, 100790, 100790, 100760, 100750, 100730, 
    100750, 100750, 100740, 100740, 100740, 100740, 100730, 100710, 100700, 
    100700, 100700, 100700, 100710, 100720, 100740, 100740, 100740, 100750, 
    100730, 100710, 100690, 100680, 100670, 100700, 100720, 100760, 100770, 
    100790, 100820, 100850, 100880, 100910, 100910, 100950, 100980, 101000, 
    101050, 101090, 101140, 101190, 101220, 101240, 101260, 101270, 101290, 
    101310, 101330, 101360, 101390, 101430, 101470, 101480, 101520, 101540, 
    101540, 101530, 101550, 101570, 101590, 101580, 101590, 101620, 101640, 
    101650, 101670, 101680, 101670, 101680, 101680, 101670, 101680, 101670, 
    101680, 101710, 101700, 101710, 101720, 101730, 101720, 101710, 101710, 
    101720, 101720, 101710, 101710, 101700, 101680, 101630, 101610, 101560, 
    101520, 101470, 101450, 101430, 101420, 101370, 101330, 101280, 101250, 
    101220, 101210, 101180, 101140, 101120, 101040, 101010, 100970, 100950, 
    100950, 100940, 100900, 100840, 100840, 100820, 100820, 100770, 100740, 
    100700, 100700, 100690, 100670, 100660, 100630, 100610, 100590, 100540, 
    100490, 100470, 100440, 100420, 100400, 100390, 100380, 100340, 100330, 
    100320, 100330, 100350, 100340, 100370, 100380, 100410, 100450, 100480, 
    100510, 100530, 100570, 100570, 100560, 100550, 100560, 100560, 100550, 
    100520, 100500, 100500, 100520, 100530, 100530, 100510, 100500, 100480, 
    100470, 100430, 100390, 100350, 100320, 100280, 100220, 100160, 100120, 
    100060, 100000, 99950, 99890, 99860, 99810, 99790, 99780, 99740, 99740, 
    99730, 99710, 99680, 99660, 99620, 99620, 99590, 99580, 99560, 99520, 
    99490, 99460, 99450, 99420, 99410, 99410, 99400, 99370, 99350, 99330, 
    99330, 99320, 99310, 99320, 99300, 99290, 99290, 99260, 99230, 99190, 
    99130, 99100, 99060, 99020, 99000, 98970, 98920, 98880, 98830, 98810, 
    98770, 98750, 98720, 98710, 98710, 98730, 98720, 98770, 98810, 98850, 
    98880, 98920, 98960, 99010, 99040, 99030, 99080, 99110, 99140, 99170, 
    99200, 99230, 99280, 99330, 99370, 99390, 99440, 99490, 99550, 99590, 
    99660, 99720, 99800, 99850, 99930, 100010, 100050, 100120, 100160, 
    100200, 100250, 100280, 100330, 100360, 100420, 100460, 100470, 100500, 
    100550, 100560, 100570, 100590, 100590, 100600, 100610, 100650, 100640, 
    100640, 100640, 100620, 100630, 100630, 100620, 100620, 100610, 100620, 
    100620, 100640, 100650, 100640, 100640, 100650, 100650, 100650, 100650, 
    100650, 100660, 100650, 100650, 100640, 100650, 100650, 100650, 100660, 
    100660, 100630, 100610, 100590, 100570, 100550, 100520, 100490, 100440, 
    100410, 100400, 100350, 100260, 100160, 100060, 99990, 99930, 99890, 
    99840, 99810, 99810, 99770, 99710, 99670, 99620, 99580, 99530, 99540, 
    99540, 99600, 99710, 99880, 99970, 100060, 100170, 100260, 100330, 
    100420, 100500, 100580, 100670, 100760, 100840, 100940, 101040, 101140, 
    101220, 101280, 101350, 101400, 101440, 101500, 101550, 101630, 101710, 
    101770, 101830, 101890, 101930, 101960, 101940, 101950, 101980, 102000, 
    102000, 102040, 102050, 102070, 102130, 102140, 102150, 102150, 102150, 
    102120, 102120, 102120, 102100, 102090, 102120, 102120, 102130, 102140, 
    102140, 102130, 102130, 102120, 102100, 102090, 102100, 102060, 102060, 
    102060, 102090, 102090, 102070, 102030, 102010, 102000, 101960, 101920, 
    101860, 101830, 101810, 101780, 101770, 101750, 101720, 101670, 101660, 
    101630, 101590, 101550, 101530, 101530, 101540, 101520, 101520, 101480, 
    101440, 101410, 101390, 101380, 101370, 101370, 101360, 101360, 101360, 
    101380, 101400, 101420, 101410, 101460, 101480, 101500, 101500, 101520, 
    101570, 101610, 101630, 101670, 101690, 101710, 101740, 101760, 101780, 
    101820, 101820, 101810, 101800, 101760, 101760, 101770, 101780, 101780, 
    101780, 101770, 101800, 101820, 101860, 101860, 101880, 101900, 101930, 
    101940, 101910, 101880, 101880, 101900, 101900, 101890, 101870, 101850, 
    101830, 101800, 101790, 101760, 101730, 101700, 101710, 101690, 101670, 
    101660, 101650, 101610, 101590, 101570, 101570, 101570, 101550, 101550, 
    101510, 101500, 101470, 101460, 101460, 101460, 101450, 101440, 101380, 
    101360, 101350, 101360, 101340, 101320, 101270, 101250, 101220, 101190, 
    101190, 101190, 101190, 101170, 101170, 101140, 101130, 101130, 101130, 
    101110, 101100, 101120, 101100, 101100, 101070, 101100, 101070, 101110, 
    101110, 101050, 101060, 101030, 101000, 101010, 101000, 101000, 101020, 
    101040, 101080, 101100, 101130, 101150, 101180, 101180, 101210, 101230, 
    101250, 101270, 101270, 101310, 101340, 101370, 101430, 101430, 101430, 
    101450, 101460, 101500, 101550, 101570, 101560, 101600, 101640, 101680, 
    101710, 101730, 101750, 101780, 101800, 101840, 101900, 101890, 101940, 
    101970, 101980, 102010, 102040, 102070, 102070, 102090, 102110, 102120, 
    102140, 102150, 102170, 102170, 102160, 102160, 102150, 102120, 102130, 
    102110, 102080, 102060, 102060, 102030, 102010, 101970, 101950, 101930, 
    101900, 101870, 101860, 101830, 101830, 101800, 101800, 101780, 101760, 
    101730, 101730, 101740, 101750, 101720, 101710, 101670, 101660, 101650, 
    101650, 101620, 101610, 101600, 101590, 101550, 101530, 101500, 101470, 
    101410, 101380, 101320, 101310, 101270, 101230, 101190, 101160, 101140, 
    101120, 101050, 100990, 100910, 100850, 100810, 100750, 100690, 100650, 
    100620, 100580, 100560, 100540, 100530, 100530, 100540, 100570, 100590, 
    100650, 100690, 100740, 100810, 100830, 100890, 100930, 100980, 101040, 
    101070, 101140, 101170, 101210, 101240, 101260, 101270, 101300, 101320, 
    101350, 101390, 101380, 101350, 101310, 101280, 101240, 101260, 101260, 
    101240, 101200, 101150, 101100, 101080, 101050, 101020, 101020, 101000, 
    100970, 100990, 101020, 101040, 101060, 101070, 101060, 101060, 101030, 
    101040, 101030, 101010, 101030, 101070, 101100, 101180, 101300, 101420, 
    101550, 101680, 101820, 101920, 102040, 102160, 102250, 102340, 102430, 
    102500, 102560, 102630, 102710, 102770, 102810, 102860, 102880, 102890, 
    102920, 102900, 102940, 102950, 102960, 103000, 102990, 102980, 102960, 
    102940, 102900, 102890, 102870, 102860, 102850, 102840, 102840, 102850, 
    102840, 102840, 102820, 102810, 102780, 102790, 102770, 102760, 102760, 
    102740, 102740, 102730, 102740, 102730, 102700, 102670, 102620, 102580, 
    102540, 102500, 102460, 102430, 102380, 102330, 102290, 102220, 102150, 
    102100, 102040, 101990, 101930, 101860, 101820, 101760, 101740, 101720, 
    101700, 101690, 101650, 101640, 101630, 101620, 101590, 101580, 101590, 
    101580, 101570, 101540, 101520, 101490, 101420, 101310, 101220, 101040, 
    100940, 100860, 100880, 100880, 100910, 100930, 100910, 100910, 100840, 
    100780, 100780, 100750, 100750, 100860, 100880, 100970, 101050, 101180, 
    101270, 101340, 101450, 101530, 101610, 101670, 101740, 101810, 101920, 
    102010, 102100, 102210, 102310, 102360, 102440, 102530, 102570, 102600, 
    102660, 102710, 102740, 102750, 102740, 102740, 102690, 102670, 102600, 
    102510, 102440, 102420, 102410, 102380, 102360, 102370, 102350, 102370, 
    102350, 102310, 102230, 102190, 102090, 101980, 101870, 101850, 101770, 
    101720, 101770, 101710, 101730, 101720, 101710, 101760, 101810, 101840, 
    101860, 101900, 101940, 101950, 101990, 102050, 102110, 102130, 102160, 
    102170, 102160, 102170, 102210, 102240, 102240, 102260, 102270, 102260, 
    102270, 102240, 102210, 102180, 102210, 102240, 102270, 102290, 102350, 
    102390, 102410, 102450, 102440, 102430, 102420, 102450, 102450, 102450, 
    102480, 102490, 102510, 102540, 102560, 102580, 102600, 102620, 102630, 
    102640, 102630, 102600, 102630, 102670, 102690, 102760, 102830, 102840, 
    102790, 102770, 102770, 102760, 102760, 102760, 102770, 102790, 102780, 
    102770, 102780, 102790, 102810, 102810, 102820, 102830, 102800, 102820, 
    102750, 102760, 102750, 102720, 102690, 102650, 102600, 102560, 102520, 
    102490, 102470, 102460, 102470, 102470, 102480, 102450, 102420, 102410, 
    102390, 102390, 102380, 102370, 102400, 102410, 102430, 102450, 102500, 
    102530, 102530, 102500, 102530, 102540, 102550, 102550, 102550, 102560, 
    102560, 102550, 102530, 102480, 102470, 102410, 102390, 102370, 102370, 
    102310, 102290, 102270, 102210, 102240, 102240, 102220, 102170, 102120, 
    102080, 102060, 102010, 101970, 101960, 101950, 101980, 101940, 101900, 
    101900, 101880, 101850, 101800, 101760, 101730, 101690, 101650, 101580, 
    101510, 101440, 101400, 101360, 101320, 101270, 101220, 101160, 101070, 
    101000, 100930, 100870, 100830, 100780, 100740, 100680, 100650, 100650, 
    100600, 100510, 100410, 100350, 100360, 100370, 100350, 100300, 100210, 
    100210, 100230, 100170, 100150, 100120, 100100, 100080, 100060, 100050, 
    100020, 100010, 100000, 99980, 99980, 99970, 99970, 99950, 99930, 99890, 
    99870, 99870, 99860, 99860, 99880, 99860, 99850, 99850, 99860, 99870, 
    99880, 99880, 99910, 99940, 99960, 99970, 99980, 100020, 100040, 100060, 
    100070, 100090, 100070, 100070, 100070, 100080, 100090, 100120, 100150, 
    100180, 100190, 100230, 100220, 100230, 100250, 100270, 100290, 100310, 
    100350, 100370, 100400, 100440, 100460, 100510, 100550, 100580, 100620, 
    100650, 100690, 100710, 100730, 100780, 100830, 100880, 100920, 100950, 
    100990, 101030, 101060, 101110, 101140, 101160, 101190, 101220, 101240, 
    101260, 101280, 101280, 101280, 101300, 101300, 101300, 101310, 101320, 
    101330, 101340, 101360, 101370, 101390, 101400, 101410, 101410, 101440, 
    101440, 101450, 101450, 101440, 101460, 101450, 101460, 101470, 101480, 
    101480, 101470, 101460, 101460, 101470, 101460, 101440, 101440, 101460, 
    101480, 101490, 101480, 101490, 101490, 101480, 101460, 101440, 101450, 
    101440, 101430, 101430, 101430, 101450, 101430, 101400, 101390, 101390, 
    101380, 101370, 101380, 101350, 101350, 101340, 101350, 101400, 101450, 
    101470, 101500, 101520, 101550, 101570, 101600, 101600, 101620, 101640, 
    101650, 101650, 101650, 101640, 101640, 101630, 101610, 101610, 101610, 
    101600, 101610, 101590, 101620, 101650, 101680, 101690, 101680, 101680, 
    101680, 101680, 101690, 101680, 101690, 101690, 101700, 101720, 101720, 
    101700, 101690, 101660, 101660, 101660, 101650, 101660, 101670, 101650, 
    101670, 101680, 101660, 101650, 101630, 101630, 101620, 101600, 101590, 
    101600, 101590, 101590, 101580, 101570, 101560, 101560, 101530, 101500, 
    101460, 101450, 101430, 101420, 101420, 101410, 101420, 101450, 101470, 
    101460, 101440, 101430, 101420, 101410, 101390, 101380, 101370, 101360, 
    101340, 101320, 101310, 101290, 101300, 101310, 101310, 101300, 101300, 
    101310, 101320, 101350, 101370, 101400, 101400, 101390, 101340, 101330, 
    101310, 101270, 101250, 101250, 101210, 101210, 101220, 101210, 101200, 
    101170, 101150, 101110, 101100, 101070, 101030, 101070, 101040, 101060, 
    101040, 101020, 101040, 101040, 101030, 101040, 101000, 100960, 100940, 
    100960, 100920, 100930, 100940, 100960, 100970, 100990, 101000, 101030, 
    101040, 101050, 101020, 101050, 101070, 101080, 101110, 101110, 101130, 
    101120, 101100, 101100, 101070, 101050, 101030, 101000, 100970, 100930, 
    100920, 100900, 100880, 100840, 100830, 100790, 100750, 100680, 100680, 
    100660, 100640, 100630, 100620, 100630, 100620, 100620, 100590, 100590, 
    100590, 100600, 100620, 100630, 100660, 100690, 100710, 100730, 100730, 
    100730, 100760, 100760, 100790, 100810, 100850, 100890, 100940, 100980, 
    101030, 101070, 101080, 101110, 101140, 101170, 101200, 101220, 101250, 
    101270, 101320, 101360, 101370, 101390, 101420, 101450, 101480, 101500, 
    101530, 101550, 101590, 101620, 101660, 101680, 101720, 101750, 101780, 
    101810, 101830, 101850, 101860, 101870, 101870, 101880, 101890, 101890, 
    101890, 101910, 101910, 101890, 101890, 101890, 101900, 101880, 101880, 
    101860, 101860, 101860, 101850, 101850, 101860, 101840, 101820, 101810, 
    101780, 101720, 101680, 101630, 101580, 101530, 101500, 101460, 101400, 
    101350, 101310, 101270, 101260, 101220, 101220, 101200, 101210, 101210, 
    101240, 101260, 101290, 101320, 101340, 101370, 101390, 101410, 101430, 
    101470, 101460, 101500, 101500, 101530, 101550, 101550, 101570, 101560, 
    101580, 101580, 101590, 101610, 101600, 101630, 101650, 101650, 101650, 
    101650, 101680, 101680, 101680, 101710, 101710, 101710, 101740, 101760, 
    101770, 101810, 101820, 101840, 101810, 101830, 101840, 101840, 101830, 
    101790, 101770, 101740, 101700, 101690, 101640, 101600, 101570, 101480, 
    101430, 101400, 101330, 101270, 101210, 101170, 101110, 101050, 101050, 
    101010, 100940, 100860, 100860, 100830, 100810, 100800, 100770, 100710, 
    100670, 100640, 100610, 100610, 100560, 100540, 100560, 100590, 100610, 
    100660, 100710, 100740, 100790, 100850, 100900, 100930, 100970, 101020, 
    101050, 101030, 101040, 101030, 101010, 101020, 101020, 100990, 100970, 
    100920, 100860, 100840, 100780, 100730, 100660, 100630, 100590, 100570, 
    100570, 100560, 100520, 100520, 100500, 100510, 100500, 100510, 100470, 
    100490, 100490, 100490, 100490, 100510, 100510, 100530, 100540, 100480, 
    100450, 100460, 100440, 100400, 100390, 100420, 100420, 100410, 100400, 
    100360, 100300, 100290, 100270, 100260, 100180, 100110, 100020, 99990, 
    99930, 99880, 99780, 99670, 99570, 99490, 99410, 99320, 99260, 99170, 
    99080, 98980, 98880, 98770, 98710, 98660, 98590, 98510, 98440, 98370, 
    98360, 98350, 98370, 98380, 98370, 98380, 98400, 98420, 98410, 98420, 
    98420, 98460, 98480, 98510, 98510, 98530, 98550, 98610, 98620, 98610, 
    98610, 98630, 98690, 98730, 98720, 98760, 98800, 98820, 98870, 98900, 
    98950, 99000, 99050, 99060, 99030, 99050, 99040, 99010, 99060, 99080, 
    99150, 99200, 99230, 99230, 99190, 99230, 99390, 99260, 99400, 99400, 
    99500, 99500, 99500, 99520, 99560, 99560, 99460, 99380, 99450, 99400, 
    99400, 99460, 99410, 99460, 99500, 99560, 99540, 99550, 99500, 99480, 
    99470, 99460, 99450, 99420, 99430, 99440, 99450, 99450, 99540, 99550, 
    99570, 99560, 99560, 99560, 99560, 99580, 99570, 99570, 99580, 99550, 
    99520, 99520, 99500, 99490, 99510, 99500, 99500, 99490, 99500, 99530, 
    99540, 99560, 99590, 99620, 99630, 99620, 99620, 99610, 99620, 99640, 
    99640, 99620, 99620, 99610, 99630, 99640, 99630, 99600, 99590, 99580, 
    99570, 99570, 99550, 99550, 99550, 99560, 99550, 99520, 99500, 99460, 
    99420, 99360, 99330, 99290, 99260, 99230, 99180, 99130, 99060, 99040, 
    99010, 98950, 98870, 98840, 98810, 98760, 98730, 98700, 98660, 98640, 
    98600, 98500, 98500, 98470, 98440, 98400, 98360, 98340, 98310, 98290, 
    98260, 98250, 98230, 98230, 98200, 98160, 98150, 98150, 98130, 98130, 
    98140, 98150, 98170, 98190, 98200, 98200, 98210, 98190, 98190, 98190, 
    98140, 98140, 98100, 98130, 98130, 98130, 98130, 98130, 98160, 98170, 
    98210, 98250, 98300, 98360, 98470, 98600, 98770, 98890, 98980, 99050, 
    99160, 99260, 99320, 99380, 99420, 99520, 99570, 99620, 99660, 99740, 
    99790, 99840, 99840, 99920, 99910, 99930, 99970, 100020, 100060, 100100, 
    100180, 100260, 100330, 100360, 100420, 100450, 100510, 100560, 100620, 
    100630, 100680, 100730, 100770, 100820, 100850, 100880, 100900, 100940, 
    100990, 101020, 101050, 101070, 101110, 101150, 101190, 101220, 101250, 
    101300, 101310, 101340, 101370, 101400, 101450, 101470, 101510, 101550, 
    101580, 101620, 101660, 101670, 101690, 101720, 101750, 101800, 101830, 
    101850, 101880, 101910, 101950, 101990, 102040, 102080, 102080, 102120, 
    102130, 102140, 102140, 102130, 102140, 102140, 102100, 102080, 102070, 
    102040, 102050, 101990, 101940, 101910, 101850, 101820, 101760, 101690, 
    101710, 101670, 101590, 101560, 101530, 101490, 101440, 101380, 101280, 
    101220, 101140, 101060, 101040, 101040, 100970, 100900, 100880, 100780, 
    100730, 100670, 100620, 100540, 100470, 100490, 100480, 100430, 100410, 
    100380, 100360, 100320, 100330, 100340, 100360, 100350, 100320, 100290, 
    100290, 100310, 100270, 100280, 100250, 100230, 100300, 100350, 100410, 
    100470, 100480, 100450, 100410, 100390, 100370, 100370, 100400, 100410, 
    100340, 100320, 100330, 100300, 100300, 100260, 100250, 100200, 100170, 
    100170, 100160, 100160, 100110, 100040, 100010, 99990, 99920, 99920, 
    99850, 99870, 99890, 99880, 99890, 99890, 99890, 99880, 99840, 99810, 
    99830, 99840, 99860, 99870, 99860, 99880, 99890, 99890, 99870, 99870, 
    99860, 99850, 99840, 99860, 99900, 99930, 99950, 99980, 99950, 99960, 
    99990, 99990, 100000, 100020, 100030, 100030, 100040, 100040, 100060, 
    100100, 100100, 100120, 100130, 100150, 100150, 100160, 100170, 100180, 
    100200, 100210, 100200, 100200, 100230, 100240, 100250, 100240, 100240, 
    100260, 100280, 100290, 100320, 100330, 100330, 100350, 100370, 100390, 
    100400, 100410, 100440, 100450, 100480, 100490, 100510, 100530, 100560, 
    100560, 100560, 100600, 100610, 100620, 100620, 100610, 100610, 100620, 
    100610, 100610, 100630, 100650, 100690, 100720, 100720, 100750, 100750, 
    100750, 100810, 100840, 100870, 100900, 100940, 100970, 101010, 101050, 
    101070, 101080, 101080, 101070, 101100, 101150, 101180, 101190, 101230, 
    101240, 101270, 101280, 101290, 101290, 101310, 101320, 101320, 101360, 
    101390, 101420, 101420, 101410, 101400, 101400, 101410, 101410, 101420, 
    101410, 101440, 101440, 101460, 101470, 101460, 101450, 101440, 101440, 
    101450, 101460, 101440, 101420, 101410, 101390, 101390, 101380, 101360, 
    101350, 101340, 101330, 101300, 101320, 101340, 101340, 101340, 101370, 
    101380, 101390, 101410, 101410, 101410, 101430, 101410, 101440, 101450, 
    101480, 101520, 101630, 101620, 101690, 101730, 101780, 101840, 101870, 
    101890, 101930, 101940, 101960, 101980, 102020, 102050, 102100, 102110, 
    102150, 102160, 102190, 102180, 102190, 102200, 102230, 102250, 102280, 
    102320, 102360, 102400, 102420, 102460, 102460, 102490, 102480, 102470, 
    102460, 102480, 102500, 102540, 102570, 102600, 102610, 102630, 102640, 
    102680, 102700, 102710, 102700, 102740, 102820, 102860, 102890, 102910, 
    102940, 102970, 103020, 103060, 103110, 103140, 103190, 103210, 103250, 
    103310, 103360, 103390, 103400, 103400, 103410, 103430, 103440, 103480, 
    103510, 103540, 103600, 103630, 103660, 103710, 103690, 103680, 103660, 
    103660, 103610, 103610, 103580, 103570, 103600, 103610, 103620, 103630, 
    103630, 103590, 103580, 103560, 103550, 103550, 103530, 103540, 103550, 
    103570, 103600, 103640, 103640, 103660, 103680, 103680, 103670, 103680, 
    103700, 103720, 103740, 103720, 103720, 103700, 103690, 103670, 103640, 
    103670, 103650, 103590, 103580, 103570, 103590, 103590, 103570, 103550, 
    103510, 103470, 103470, 103480, 103430, 103400, 103380, 103370, 103330, 
    103320, 103270, 103240, 103210, 103170, 103150, 103130, 103110, 103040, 
    103030, 103020, 103000, 102990, 102980, 102930, 102910, 102870, 102840, 
    102810, 102790, 102760, 102750, 102710, 102690, 102640, 102620, 102580, 
    102540, 102500, 102470, 102400, 102370, 102320, 102260, 102210, 102160, 
    102130, 102120, 102090, 102030, 101970, 101880, 101830, 101780, 101730, 
    101700, 101650, 101610, 101570, 101510, 101470, 101440, 101380, 101330, 
    101270, 101220, 101160, 101090, 101050, 101020, 100980, 100950, 100910, 
    100860, 100800, 100740, 100690, 100650, 100600, 100550, 100510, 100480, 
    100470, 100430, 100390, 100360, 100290, 100240, 100210, 100180, 100150, 
    100160, 100180, 100190, 100240, 100280, 100320, 100330, 100370, 100390, 
    100430, 100450, 100480, 100510, 100550, 100590, 100630, 100670, 100690, 
    100700, 100740, 100770, 100820, 100850, 100840, 100860, 100870, 100890, 
    100910, 100930, 100920, 100920, 100930, 100990, 101000, 100990, 101010, 
    101040, 101110, 101170, 101170, 101190, 101200, 101220, 101220, 101210, 
    101200, 101200, 101190, 101190, 101170, 101140, 101140, 101170, 101170, 
    101160, 101140, 101140, 101140, 101150, 101160, 101160, 101160, 101160, 
    101130, 101110, 101110, 101090, 101060, 101010, 100970, 100920, 100890, 
    100870, 100830, 100790, 100730, 100720, 100710, 100650, 100530, 100450, 
    100350, 100260, 100230, 100180, 100090, 99990, 99890, 99760, 99670, 
    99580, 99450, 99330, 99250, 99210, 99150, 99170, 99150, 99140, 99170, 
    99170, 99140, 99110, 99100, 99070, 99030, 99000, 98960, 98940, 98910, 
    98940, 98920, 98920, 98920, 98920, 98900, 98890, 98880, 98870, 98890, 
    98880, 98850, 98840, 98820, 98810, 98800, 98770, 98710, 98720, 98670, 
    98620, 98630, 98580, 98550, 98540, 98520, 98530, 98540, 98530, 98520, 
    98500, 98470, 98460, 98430, 98430, 98410, 98430, 98440, 98460, 98450, 
    98430, 98450, 98440, 98500, 98530, 98580, 98700, 98770, 98880, 98930, 
    99010, 99110, 99180, 99300, 99380, 99440, 99490, 99540, 99610, 99640, 
    99690, 99740, 99780, 99820, 99870, 99900, 99970, 99990, 100070, 100100, 
    100140, 100170, 100210, 100230, 100260, 100290, 100290, 100310, 100300, 
    100320, 100340, 100330, 100350, 100380, 100410, 100410, 100420, 100430, 
    100460, 100450, 100460, 100470, 100460, 100470, 100490, 100520, 100520, 
    100540, 100530, 100530, 100520, 100510, 100500, 100490, 100480, 100480, 
    100490, 100500, 100500, 100540, 100550, 100570, 100600, 100620, 100650, 
    100680, 100710, 100720, 100740, 100740, 100750, 100790, 100810, 100790, 
    100810, 100830, 100850, 100880, 100870, 100870, 100920, 100910, 100940, 
    100950, 100980, 100980, 100990, 100970, 100960, 100950, 100950, 100940, 
    100940, 100950, 100950, 101000, 101060, 101070, 101060, 101120, 101160, 
    101170, 101160, 101210, 101230, 101250, 101290, 101350, 101390, 101400, 
    101430, 101440, 101470, 101490, 101530, 101560, 101620, 101680, 101720, 
    101770, 101800, 101810, 101760, 101760, 101770, 101760, 101760, 101790, 
    101810, 101800, 101810, 101840, 101890, 101910, 101880, 101850, 101820, 
    101760, 101720, 101700, 101680, 101650, 101630, 101630, 101610, 101570, 
    101530, 101490, 101460, 101420, 101370, 101350, 101320, 101300, 101280, 
    101280, 101260, 101240, 101220, 101190, 101150, 101150, 101090, 101080, 
    101070, 101070, 101050, 101050, 101060, 101090, 101090, 101120, 101120, 
    101120, 101120, 101100, 101090, 101060, 101040, 101030, 101060, 101000, 
    100930, 100860, 100810, 100780, 100740, 100720, 100710, 100680, 100650, 
    100610, 100560, 100510, 100490, 100470, 100430, 100410, 100360, 100320, 
    100300, 100210, 100160, 100110, 100060, 100000, 99930, 99890, 99860, 
    99780, 99760, 99700, 99670, 99620, 99580, 99520, 99510, 99490, 99430, 
    99390, 99330, 99300, 99280, 99250, 99220, 99190, 99190, 99170, 99140, 
    99120, 99120, 99110, 99110, 99120, 99150, 99190, 99210, 99220, 99230, 
    99240, 99270, 99250, 99270, 99250, 99280, 99280, 99330, 99330, 99390, 
    99420, 99450, 99460, 99500, 99490, 99550, 99630, 99670, 99690, 99760, 
    99800, 99800, 99930, 99930, 99980, 100000, 100010, 100030, 100030, 
    100030, 100050, 100050, 100040, 100040, 100060, 100070, 100110, 100130, 
    100120, 100130, 100120, 100120, 100120, 100120, 100120, 100110, 100110, 
    100110, 100100, 100120, 100120, 100110, 100100, 100090, 100080, 100070, 
    100050, 100030, 100020, 100020, 100020, 100010, 99990, 99980, 99950, 
    99950, 99940, 99910, 99900, 99890, 99870, 99850, 99830, 99800, 99780, 
    99760, 99740, 99700, 99700, 99670, 99700, 99610, 99560, 99560, 99600, 
    99610, 99610, 99620, 99630, 99630, 99630, 99660, 99700, 99750, 99790, 
    99840, 99860, 99890, 99920, 99950, 99990, 100040, 100080, 100100, 100130, 
    100150, 100170, 100210, 100250, 100270, 100320, 100360, 100400, 100420, 
    100420, 100430, 100460, 100470, 100430, 100410, 100390, 100390, 100400, 
    100410, 100400, 100360, 100290, 100210, 100130, 100020, 99890, 99780, 
    99720, 99550, 99440, 99280, 99010, 98760, 98470, 98130, 97830, 97450, 
    97090, 96800, 96590, 96380, 96170, 95990, 95800, 95680, 95590, 95540, 
    95460, 95420, 95360, 95330, 95360, 95400, 95450, 95520, 95610, 95670, 
    95720, 95730, 95700, 95710, 95800, 95890, 95970, 96040, 96110, 96180, 
    96250, 96260, 96430, 96500, 96550, 96570, 96610, 96670, 96730, 96780, 
    96860, 96920, 96990, 97070, 97160, 97230, 97320, 97410, 97470, 97550, 
    97630, 97700, 97770, 97830, 97880, 97970, 98030, 98120, 98210, 98240, 
    98310, 98390, 98490, 98560, 98630, 98690, 98760, 98800, 98830, 98840, 
    98890, 98880, 98880, 98850, 98840, 98840, 98820, 98800, 98770, 98760, 
    98780, 98800, 98830, 98860, 98900, 98960, 99010, 99050, 99100, 99090, 
    99110, 99150, 99230, 99290, 99360, 99440, 99490, 99530, 99620, 99690, 
    99720, 99760, 99820, 99890, 99910, 99980, 100020, 100040, 100080, 100090, 
    100130, 100180, 100180, 100190, 100220, 100220, 100270, 100270, 100290, 
    100290, 100300, 100290, 100330, 100370, 100390, 100440, 100460, 100520, 
    100560, 100590, 100630, 100680, 100730, 100790, 100860, 100940, 100990, 
    101050, 101100, 101190, 101240, 101260, 101300, 101330, 101350, 101340, 
    101380, 101420, 101470, 101510, 101530, 101550, 101560, 101520, 101560, 
    101550, 101550, 101570, 101560, 101550, 101530, 101470, 101340, 101240, 
    101120, 101010, 100850, 100720, 100610, 100510, 100490, 100470, 100440, 
    100380, 100370, 100350, 100380, 100400, 100370, 100350, 100430, 100480, 
    100480, 100480, 100480, 100470, 100390, 100370, 100370, 100300, 100240, 
    100140, 99990, 99800, 99640, 99450, 99220, 98970, 98720, 98410, 98160, 
    98260, 98460, 98550, 98520, 98540, 98630, 98660, 98640, 98700, 98760, 
    98780, 98810, 98860, 98850, 98910, 98980, 99040, 99110, 99190, 99290, 
    99390, 99470, 99530, 99590, 99660, 99700, 99770, 99830, 99870, 99940, 
    100030, 100100, 100170, 100240, 100280, 100350, 100390, 100450, 100510, 
    100560, 100580, 100620, 100690, 100730, 100770, 100820, 100820, 100820, 
    100830, 100850, 100850, 100850, 100870, 100910, 100930, 100930, 100940, 
    100940, 100920, 100900, 100900, 100880, 100890, 100870, 100850, 100820, 
    100810, 100820, 100800, 100770, 100760, 100720, 100720, 100710, 100720, 
    100720, 100730, 100750, 100760, 100780, 100790, 100780, 100760, 100770, 
    100770, 100770, 100760, 100750, 100750, 100730, 100710, 100720, 100700, 
    100660, 100640, 100640, 100620, 100580, 100560, 100540, 100520, 100540, 
    100530, 100510, 100470, 100440, 100410, 100380, 100350, 100370, 100340, 
    100340, 100350, 100370, 100370, 100380, 100380, 100390, 100390, 100370, 
    100370, 100350, 100330, 100340, 100360, 100370, 100410, 100440, 100440, 
    100460, 100460, 100480, 100480, 100490, 100500, 100510, 100520, 100540, 
    100530, 100540, 100550, 100540, 100520, 100510, 100510, 100510, 100510, 
    100530, 100530, 100570, 100590, 100600, 100610, 100640, 100650, 100650, 
    100670, 100670, 100670, 100680, 100690, 100690, 100700, 100690, 100700, 
    100700, 100690, 100690, 100680, 100660, 100650, 100650, 100640, 100660, 
    100690, 100700, 100680, 100690, 100690, 100640, 100670, 100660, 100660, 
    100690, 100700, 100700, 100700, 100710, 100760, 100760, 100750, 100740, 
    100730, 100710, 100720, 100730, 100760, 100780, 100790, 100750, 100750, 
    100700, 100670, 100610, 100560, 100490, 100450, 100420, 100400, 100370, 
    100340, 100310, 100230, 100200, 100110, 100080, 100050, 100020, 100000, 
    100000, 100020, 100040, 100140, 100150, 100200, 100190, 100180, 100160, 
    100230, 100260, 100310, 100320, 100320, 100330, 100340, 100270, 100220, 
    100210, 100170, 100110, 100050, 99990, 99960, 99930, 99860, 99870, 99860, 
    99820, 99760, 99700, 99690, 99690, 99680, 99680, 99700, 99680, 99700, 
    99720, 99770, 99740, 99740, 99760, 99820, 99860, 99920, 99940, 99970, 
    100050, 100160, 100250, 100360, 100420, 100490, 100570, 100630, 100670, 
    100700, 100760, 100820, 100870, 100900, 100930, 100920, 100940, 100960, 
    101010, 101010, 101020, 101030, 101040, 101070, 101070, 101070, 101080, 
    101110, 101100, 101090, 101110, 101130, 101150, 101130, 101160, 101190, 
    101230, 101230, 101250, 101230, 101260, 101270, 101250, 101270, 101300, 
    101310, 101300, 101270, 101280, 101290, 101300, 101320, 101340, 101350, 
    101330, 101320, 101320, 101330, 101340, 101340, 101360, 101390, 101400, 
    101420, 101410, 101410, 101430, 101410, 101410, 101400, 101390, 101400, 
    101400, 101420, 101470, 101500, 101520, 101510, 101520, 101500, 101460, 
    101440, 101390, 101360, 101300, 101240, 101210, 101180, 101130, 101070, 
    101020, 100950, 100900, 100810, 100760, 100710, 100660, 100600, 100560, 
    100580, 100580, 100590, 100640, 100700, 100730, 100790, 100820, 100860, 
    100890, 100840, 100810, 100760, 100660, 100590, 100470, 100350, 100250, 
    100160, 100070, 99950, 99880, 99790, 99650, 99560, 99410, 99380, 99320, 
    99190, 99110, 99060, 98970, 98880, 98800, 98700, 98620, 98580, 98580, 
    98640, 98730, 98790, 98850, 99010, 99040, 99120, 99190, 99240, 99310, 
    99320, 99360, 99400, 99420, 99420, 99400, 99330, 99290, 99270, 99250, 
    99230, 99240, 99210, 99200, 99140, 99090, 99060, 99050, 99060, 99070, 
    99060, 99070, 99110, 99150, 99190, 99230, 99260, 99260, 99250, 99350, 
    99360, 99380, 99410, 99450, 99480, 99520, 99570, 99610, 99620, 99620, 
    99620, 99590, 99590, 99580, 99610, 99490, 99560, 99580, 99600, _, 99600, 
    99610, 99640, 99650, 99680, 99700, 99720, 99650, 99710, 99760, 99800, 
    99820, 99880, 99930, 99970, 100030, 100080, 100130, 100160, 100250, 
    100320, 100400, 100490, 100590, 100650, 100700, 100740, 100810, 100880, 
    100900, 100930, 100960, 100980, 100990, 101040, 101100, 101140, 101150, 
    101180, 101210, 101170, 101140, 101120, 101120, 101130, 101140, 101140, 
    101140, 101090, 101010, 100980, 100960, 100860, 100840, 100860, 100900, 
    100990, 101060, 101180, 101280, 101340, 101390, 101430, 101470, 101480, 
    101490, 101510, 101600, 101620, 101630, 101640, 101660, 101680, 101670, 
    101660, 101660, 101670, 101660, 101650, 101660, 101640, 101610, 101610, 
    101620, 101560, 101520, 101490, 101460, 101400, 101350, 101320, _, 
    101160, 101120, 101090, 101060, 101050, 100990, 100950, 100930, 100930, 
    100930, 100950, 100940, 100960, 101010, 101070, 101120, 101150, 101180, 
    101220, 101250, 101280, 101310, 101320, _, 101420, 101450, 101490, 
    101510, 101510, 101500, 101500, 101500, 101500, 101500, 101500, 101610, 
    101610, 101600, 101580, 101590, 101590, 101560, 101520, 101500, 101460, 
    101430, 101430, _, 101470, 101470, 101500, 101530, 101540, 101540, 
    101550, 101560, 101530, 101510, 101530, 101590, 101590, 101590, 101590, 
    101600, 101600, 101600, 101620, 101620, 101630, 101620, 101620, 101640, 
    101670, 101700, 101720, 101720, 101740, 101730, 101700, 101660, 101630, 
    101620, 101620, 101600, 101600, 101590, 101570, 101560, 101510, 101480, 
    101460, 101440, 101410, 101370, 101360, 101310, 101300, 101280, 101260, 
    101250, 101240, 101230, 101190, 101180, 101160, 101120, 101110, 101030, 
    101030, 101050, 101040, 101020, 101020, 101000, 100990, 100990, 100970, 
    100940, 100920, 100930, 100920, 100970, 101000, 100980, 100980, 100960, 
    100960, 100940, 100960, 100970, 100950, 100940, 100940, 100940, 100960, 
    100960, 100950, 100950, 100950, 100930, 100900, 100870, 100880, 100770, 
    100790, 100780, 100790, 100770, 100760, 100790, 100840, 100850, 100870, 
    100910, 100960, 100930, 100930, 100920, 100920, 100970, 101010, 101050, 
    101070, 101070, 101070, 101070, 101050, 101120, 101120, 101140, 101140, 
    101160, 101140, 101140, 101090, 101030, 100990, 100930, 100900, 100830, 
    100780, 100730, 100690, 100660, 100640, 100610, 100560, 100520, 100490, 
    100470, 100440, 100490, 100500, 100500, 100530, 100560, 100580, 100620, 
    100640, 100640, 100650, 100670, 100730, 100820, 100880, 100890, 100940, 
    100990, 101040, 101090, 101110, 101130, 101150, 101170, 101210, 101080, 
    101130, 101180, 101220, 101240, 101260, 101290, 101330, 101330, 101330, 
    101340, 101380, 101400, 101450, 101480, 101490, 101510, 101530, 101560, 
    101580, 101600, 101620, 101630, 101610, 101530, 101550, 101570, 101600, 
    101630, 101670, 101680, 101680, 101640, 101610, 101630, 101680, 101630, 
    101630, 101620, 101640, 101650, 101670, 101670, 101690, 101720, 101720, 
    101700, 101690, 101650, 101700, 101750, 101810, 101850, 101840, 101850, 
    101910, 101970, 101990, 101970, 101960, 102030, 102080, 102130, 102200, 
    102250, 102280, 102280, 102310, 102370, 102410, 102420, 102430, 102450, 
    102470, 102510, 102540, 102590, 102590, 102570, 102550, 102540, 102520, 
    102510, 102490, 102440, 102420, 102410, 102410, 102370, 102340, 102300, 
    102250, 102180, 102140, 102120, 102070, 101980, 101970, 101940, 101900, 
    101870, 101830, 101790, 101760, 101720, 101630, 101580, 101520, 101510, 
    101490, 101460, 101440, 101430, 101410, 101390, 101360, 101300, 101280, 
    101280, 101280, 101200, 101220, 101230, 101250, 101250, 101240, 101220, 
    101190, 101150, 101140, 101090, 101040, 100960, 100920, 100890, 100810, 
    100720, 100690, 100620, 100550, 100480, 100410, 100310, 100220, 100050, 
    99910, 99800, 99770, 99740, 99700, 99650, 99590, 99540, 99530, 99520, 
    99480, 99310, 99130, 98980, 98810, 98610, 98240, 97840, 97520, 97230, 
    97130, 97200, 97220, 97180, 97230, 97320, 97410, 97530, 97690, 97860, 
    97990, 98110, 98230, 98300, 98380, 98470, 98560, 98630, 98680, 98740, 
    98820, 98900, 99010, 99170, 99330, 99510, 99660, 99910, 100100, 100280, 
    100430, 100510, 100550, 100570, 100580, 100570, 100550, 100640, 100770, 
    100950, 101010, 101030, 101050, 101080, 101060, 101020, 100930, 100790, 
    100630, 100490, 100380, 100120, 99980, 99800, 99600, 99380, 99210, 99090, 
    98970, 98880, 98790, 98730, 98660, 98700, 98650, 98610, 98570, 98540, 
    98510, 98490, 98430, 98390, 98360, 98370, 98380, 98450, 98460, 98500, 
    98550, 98590, 98660, 98710, 98760, 98830, 98880, 98900, 98930, 99020, 
    99060, 99090, 99120, 99130, 99120, 99130, 99130, 99120, 99070, 99030, 
    99000, 99170, 99200, 99260, 99300, 99350, 99400, 99480, 99540, 99580, 
    99580, 99580, 99630, 99650, 99640, 99620, 99570, 99500, 99400, 99410, 
    99390, 99400, 99390, 99350, 99330, 99330, 99340, 99290, 99230, 99180, 
    99090, 98950, 98760, 98620, 98520, 98410, 98350, 98320, 98380, 98510, 
    98660, 98780, 98930, 99070, 99130, 99130, 99140, 99130, 99180, 99030, 
    98910, 99050, 99310, 99550, 99670, 99800, 99890, 100000, 100110, 100230, 
    100320, 100360, 100420, 100480, 100530, 100560, 100590, 100630, 100660, 
    100690, 100740, 100780, 100810, 100790, 100820, 100860, 100920, 100960, 
    100980, 100990, 101000, 101020, 101040, 101050, 101070, 101150, 101170, 
    101210, 101230, 101240, 101260, 101290, 101300, 101310, 101290, 101280, 
    101280, 101260, 101260, 101290, 101310, 101320, 101330, 101310, 101280, 
    101240, 101210, 101210, 101220, 101210, 101220, 101220, 101210, 101200, 
    101200, 101200, 101210, 101230, 101230, 101220, 101190, 101210, 101230, 
    101270, 101300, 101330, 101350, 101360, 101370, 101370, 101370, 101370, 
    101390, 101440, 101440, 101430, 101410, 101420, 101450, 101460, 101470, 
    101480, 101470, 101460, 101470, 101560, 101580, 101620, 101620, 101640, 
    101660, 101670, 101690, 101700, 101740, 101740, 101750, 101750, 101790, 
    101820, 101840, 101860, 101880, 101910, 101950, 101950, 101930, 101920, 
    101930, 102030, 102060, 102080, 102120, 102160, 102200, 102240, 102250, 
    102240, 102250, 102250, 102290, 102340, 102360, 102380, 102420, 102430, 
    102440, 102460, 102490, 102510, 102520, 102520, 102540, 102510, 102530, 
    102560, 102600, 102640, 102680, 102700, 102740, 102790, 102830, 102870, 
    102890, 102870, 102910, 102950, 102970, 103000, 103020, 103020, 103040, 
    103070, 103070, 103070, 103060, 103030, 103050, 103060, 103090, 103110, 
    103120, 103130, 103140, 103140, 103140, 103130, 103130, 103090, 103080, 
    103070, 103080, 103080, 103070, 103060, 103060, 103070, 103060, 103040, 
    103010, 103070, 103070, 103080, 103100, 103130, 103120, 103110, 103110, 
    103100, 103080, 103050, 103020, 103010, 102970, 102940, 102920, 102900, 
    102870, 102870, 102870, 102870, 102850, 102820, 102800, 102860, 102850, 
    102850, 102850, 102860, 102880, 102890, 102890, 102910, 102920, 102930, 
    102950, 103030, 103080, 103090, 103070, 103060, 103080, 103120, 103150, 
    103120, 103090, 103080, 103090, 103080, 103070, 103070, 103120, 103150, 
    103160, 103160, 103170, 103160, 103160, 103160, 103180, 103150, 103190, 
    103220, 103250, 103270, 103280, 103320, 103330, 103330, 103320, 103310, 
    103290, 103310, 103330, 103360, 103360, 103370, 103370, 103370, 103390, 
    103390, 103410, 103400, 103420, 103530, 103550, 103580, 103580, 103550, 
    103560, 103550, 103520, 103510, 103470, 103420, 103370, 103290, 103260, 
    103240, 103260, 103240, 103230, 103220, 103210, 103180, 103150, 103130, 
    103110, 103130, 103110, 103100, 103120, 103140, 103200, 103260, 103330, 
    103410, 103470, 103570, 103660, _, 103820, 103910, 103980, 104060, 
    104010, 104090, 104150, 104160, 104170, 104170, 104210, 104230, 104260, 
    104310, 104330, 104350, 104350, 104330, 104250, 104240, 104210, 104160, 
    104100, _, 104050, 104000, 103940, 103860, 103790, 103760, 103730, 
    103640, 103590, 103580, 103580, 103630, 103530, 103470, 103450, 103450, 
    103450, 103460, 103510, 103560, 103590, 103580, 103570, _, 103740, 
    103720, 103730, 103720, 103630, 103530, 103440, 103300, 103230, 103130, 
    103090, 103060, 103080, 103020, 102930, 102860, 102830, 102750, 102630, 
    102520, 102420, 102310, 102230, _, 101990, 101910, 101830, 101710, 
    101560, 101420, 101260, 101150, 101090, 101030, 101000, 101310, 101370, 
    101460, 101550, 101630, 101790, 101970, 102120, 102260, 102360, 102460, 
    102610, 102610, 102710, 102820, 102920, 102900, 102990, 103070, 103120, 
    103200, 103230, 103280, 103330, 103370, 103410, 103440, 103470, 103500, 
    103540, 103530, 103500, 103480, 103470, 103480, 103470, 103470, 103480, 
    103470, 103470, 103490, 103490, 103480, 103470, 103440, 103440, 103460, 
    103440, 103430, 103380, 103400, 103390, 103370, 103370, 103340, 103320, 
    103310, 103270, 103210, 103150, 103110, 103080, 103050, 103040, 103040, 
    103030, 103020, 102990, 102950, 102920, 102880, 102880, 102830, 102790, 
    102780, 102760, 102760, 102750, 102740, 102740, 102760, 102750, 102740, 
    102740, 102770, 102740, 102760, 102800, 102810, 102820, 102850, 102850, 
    102860, 102890, 102890, 102880, 102890, 102870, 102900, 102920, 102950, 
    102970, 102970, 102980, 103000, 103000, 103010, 103030, 103030, 103050, 
    103080, 103100, 103140, 103160, 103160, 103160, 103150, 103160, 103150, 
    103150, 103150, 103130, 103150, 103160, 103170, 103150, 103130, 103100, 
    103090, 103070, 103050, 103040, 103040, 103050, 103050, 103050, 103040, 
    103040, 103020, 103020, 103000, 102990, 103000, 103000, 103010, 102970, 
    102960, 102950, 102940, 102920, 102900, 102890, 102880, 102870, 102860, 
    102840, 102810, 102800, 102800, 102820, 102810, 102820, 102810, 102790, 
    102780, 102770, 102760, 102750, 102720, 102730, 102710, 102710, 102700, 
    102690, 102690, 102660, 102650, 102660, 102640, 102630, 102640, 102640, 
    102660, 102690, 102690, 102690, 102690, 102690, 102690, 102700, 102690, 
    102680, 102680, 102690, 102700, 102710, 102720, 102710, 102710, 102690, 
    102700, 102700, 102700, 102700, 102720, 102730, 102740, 102780, 102790, 
    102790, 102790, 102800, 102800, 102820, 102820, 102820, 102820, 102830, 
    102850, 102870, 102890, 102890, 102900, 102900, 102900, 102910, 102910, 
    102900, 102910, 102930, 102960, 102980, 102980, 102980, 103000, 103010, 
    103010, 103010, 103000, 103010, 103020, 103060, 103060, 103050, 103050, 
    103050, 103030, 103020, 103020, 103010, 103000, 103010, 103010, 103020, 
    103010, 103030, 103040, 103030, 103010, 103010, 102990, 102990, 102990, 
    102970, 102950, 102950, 102960, 102950, 102930, 102900, 102880, 102840, 
    102820, 102800, 102770, 102740, 102690, 102670, 102660, 102670, 102630, 
    102600, 102560, 102530, 102500, 102490, 102460, 102440, 102450, 102460, 
    102460, 102470, 102440, 102410, 102390, 102350, 102330, 102310, 102310, 
    102300, 102300, 102290, 102310, 102320, 102320, 102310, 102320, 102320, 
    102310, 102310, 102310, 102320, 102330, 102330, 102330, 102370, 102380, 
    102380, 102380, 102360, 102370, 102370, 102380, 102370, 102380, 102400, 
    102410, 102420, 102430, 102420, 102430, 102440, 102420, 102430, 102440, 
    102440, 102440, 102450, 102440, 102440, 102460, 102440, 102430, 102440, 
    102450, 102420, 102410, 102430, 102430, 102440, 102470, 102510, 102500, 
    102530, 102530, 102540, 102560, 102570, 102570, 102580, 102590, 102580, 
    102600, 102600, 102610, 102600, 102610, 102600, 102580, 102580, 102570, 
    102560, 102580, 102580, 102560, 102530, 102530, 102520, 102480, 102500, 
    102460, 102420, 102380, 102340, 102260, 102230, 102220, 102180, 102150, 
    102110, 102060, 102000, 101940, 101910, 101850, 101810, 101770, 101730, 
    101690, 101660, 101660, 101630, 101540, 101500, 101450, 101380, 101290, 
    101170, 101090, 101000, 100900, 100800, 100660, 100520, 100360, 100170, 
    100000, 99800, 99590, 99400, 99210, 99030, 98860, 98700, 98550, 98370, 
    98270, 98140, 98070, 98030, 98000, 97990, 97950, 98020, 98110, 98210, 
    98330, 98480, 98600, 98740, 98950, 99230, 99430, 99560, 99810, 100040, 
    100180, 100370, 100540, 100690, 100810, 100950, 101080, 101230, 101370, 
    101470, 101530, 101560, 101650, 101730, 101770, 101790, 101840, 101860, 
    101880, 101910, 101940, 101980, 101990, 102040, 102060, 102080, 102100, 
    102080, 102100, 102090, 102090, 102060, 102040, 102000, 101960, 101930, 
    101920, 101890, 101840, 101790, 101740, 101650, 101590, 101560, 101520, 
    101470, 101450, 101410, 101370, 101320, 101280, 101220, 101170, 101160, 
    101120, 101090, 101040, 100990, 100980, 100940, 100920, 100900, 100850, 
    100790, 100760, 100740, 100710, 100670, 100630, 100630, 100630, 100590, 
    100600, 100610, 100630, 100630, 100630, 100660, 100710, 100740, 100780, 
    100780, 100810, 100820, 100850, 100880, 100920, 100920, 100920, 100920, 
    100910, 100880, 100870, 100850, 100830, 100780, 100750, 100700, 100670, 
    100630, 100600, 100590, 100570, 100570, 100520, 100520, 100500, 100520, 
    100520, 100530, 100540, 100560, _, 100560, 100580, 100590, 100600, 
    100630, 100610, 100600, 100580, 100600, 100610, 100610, 100610, 100650, 
    100670, 100700, 100760, 100830, 100900, 100950, 100980, 101020, 101050, 
    101070, 101100, 101090, 101120, 101110, 101160, 101260, 101300, 101320, 
    101360, 101410, 101440, 101450, 101470, 101480, 101460, 101490, 101530, 
    101550, 101620, 101660, 101710, 101740, 101750, 101750, 101760, 101770, 
    101770, 101780, 101770, 101770, 101770, 101770, 101780, 101830, 101850, 
    101870, 101880, 101910, 101910, 101890, 101880, 101850, 101840, 101780, 
    101730, 101700, 101630, 101580, 101550, 101440, 101420, 101420, 101380, 
    101350, 101320, 101300, 101290, 101290, 101320, 101300, 101290, 101270, 
    101260, 101240, 101230, 101210, 101220, 101180, 101180, 101200, 101190, 
    101190, 101170, 101150, 101130, 101110, 101110, 101090, 101060, 101070, 
    101060, 101050, 101040, 101070, 101040, 101070, 101050, 101010, 100960, 
    _, 100860, 100850, 100800, 100730, 100670, 100620, 100550, 100480, 
    100440, 100390, 100370, 100350, 100350, 100340, 100360, 100400, 100440, 
    100480, 100520, 100560, 100600, 100630, 100670, 100700, 100730, 100780, 
    100820, 100860, 100880, 100910, 100940, _, 100980, 101000, 101020, 
    101040, 101050, 101080, 101100, 101130, 101160, 101190, 101200, 101190, 
    101180, 101170, 101190, 101160, 101170, 101160, 101170, 101170, 101180, 
    101170, 101170, 101140, 101140, 101110, 101100, 101080, 101070, 101070, 
    101050, 101050, 101050, 101050, 101040, 101030, 100990, 100980, 100970, 
    100960, 100960, 100960, 100980, 100990, 101000, 101010, 101010, 101020, 
    101020, 101010, 101030, 101040, 101040, 101070, 101090, 101120, 101140, 
    101170, 101190, 101210, _, 101240, 101230, 101260, 101290, 101310, 
    101350, 101380, 101430, 101470, 101510, _, 101550, _, 101620, 101650, 
    101710, 101790, 101880, 101930, 101990, 102050, 102080, 102130, 102180, 
    102210, 102240, 102280, 102310, 102350, 102370, 102410, 102460, 102500, 
    102510, 102530, 102540, 102560, 102600, 102610, 102650, 102700, 102720, 
    102720, 102760, 102770, 102790, 102790, 102780, 102790, 102780, 102790, 
    102810, 102840, 102850, 102860, 102850, 102880, 102860, 102840, 102810, 
    102800, 102810, 102780, 102790, 102780, 102760, 102740, 102750, 102730, 
    102700, 102690, 102670, 102640, _, 102600, 102570, 102570, 102560, 
    102560, 102550, 102540, 102540, 102540, 102510, 102500, 102460, 102470, 
    102450, 102430, 102430, 102400, 102380, 102380, 102350, 102310, 102290, 
    _, _, 102230, 102200, 102180, 102190, 102180, 102150, 102120, 102110, 
    102070, 102030, 102000, 101960, 101940, 101930, 101900, 101870, 101850, 
    101830, 101810, 101790, 101750, 101720, 101690, 101660, 101660, 101660, 
    101660, 101640, 101640, 101620, 101600, 101620, 101630, 101610, 101620, 
    101610, 101620, 101630, 101620, 101650, 101680, 101680, 101690, 101700, 
    101690, 101680, 101690, _, _, 101720, 101740, 101750, 101750, 101760, 
    101780, _, _, 101800, 101800, 101800, 101790, 101810, 101810, 101790, 
    101800, 101790, 101800, 101810, 101810, 101800, 101790, 101790, 101770, 
    101760, 101750, 101750, 101740, 101730, 101710, 101710, 101720, 101700, 
    101690, 101680, 101670, 101670, 101660, 101660, 101620, 101610, 101580, 
    101580, 101560, 101560, 101540, 101520, 101490, 101460, 101440, 101390, 
    101370, 101340, 101310, 101260, 101220, 101170, 101090, 101020, 100940, 
    100860, 100810, 100730, 100610, 100480, 100370, 100260, 100170, 100080, 
    100030, _, 99980, 99980, 100050, 100040, 100100, 100150, 100190, 100230, 
    100310, 100360, 100450, 100510, 100570, 100640, 100730, 100810, 100840, 
    100890, 100950, 100990, 101030, 101060, 101060, 101070, 101060, 101040, 
    101030, 101030, 101040, 100980, 100930, 100950, 100910, 100880, 100800, 
    100770, 100750, 100700, 100690, 100640, 100590, 100510, 100450, 100350, 
    100300, 100300, 100290, 100300, 100320, 100370, 100410, 100530, 100590, 
    100670, 100700, 100750, 100780, 100790, 100850, 100880, 100840, 100870, 
    100860, 100810, 100830, 100780, 100710, 100610, 100470, 100370, 100280, 
    100220, 100150, 100090, 100070, 100060, 100080, 100090, 100130, 100170, 
    100210, 100250, 100290, 100310, 100340, 100400, 100460, 100520, 100600, 
    100690, 100750, 100820, 100900, 100990, 101070, 101140, 101190, 101220, 
    101270, 101330, 101370, 101410, 101480, 101530, 101540, 101580, 101600, 
    101620, 101640, 101670, 101670, 101680, 101720, 101730, 101730, 101710, 
    101690, 101670, 101620, 101560, 101490, 101440, 101420, 101450, 101510, 
    101550, 101580, 101650, 101680, 101720, 101740, 101760, 101760, 101750, 
    101760, 101770, 101780, 101790, 101770, 101730, 101720, 101700, 101650, 
    101600, 101540, 101480, 101430, 101430, 101390, 101340, 101300, 101230, 
    101210, 101170, 101150, 101120, 101110, 101090, 101080, 101100, 101110, 
    101130, 101120, 101110, 101100, 101090, 101080, 101060, 101020, 100990, 
    100980, 100960, 100960, 100930, 100920, 100910, 100890, 100900, 100910, 
    100940, 100940, 101010, 101090, 101170, 101230, 101300, 101360, 101420, 
    101480, 101540, 101600, 101640, 101700, 101730, 101800, 101870, 101930, 
    101990, 102020, 102020, 102020, 102080, 102120, 102150, 102170, 102160, 
    102150, 102200, 102230, 102290, 102300, 102350, 102390, 102400, 102390, 
    102420, 102450, 102460, 102490, 102510, 102550, 102610, 102640, 102670, 
    102670, 102690, 102700, 102720, 102740, 102760, 102740, 102750, 102750, 
    102750, 102750, 102740, 102720, 102700, 102680, 102640, 102580, 102520, 
    102470, 102430, 102370, 102340, 102290, 102240, 102180, 102130, 102050, 
    102010, 101940, 101900, 101840, 101780, 101720, 101680, 101650, 101610, 
    101550, 101510, 101430, 101360, 101290, 101240, 101180, 101140, 101100, 
    101060, 101040, 101000, 100950, 100910, 100870, _, 100770, 100710, 
    100660, 100620, 100580, 100550, 100520, 100470, 100390, 100380, 100370, 
    100390, 100410, 100440, 100470, 100460, 100470, 100500, 100530, 100540, 
    100590, 100620, 100650, 100690, 100740, 100760, 100790, 100810, 100830, 
    100860, 100880, 100900, 100900, 100920, 100900, 100930, 100920, 100950, 
    100960, 100980, 100980, 101000, 100990, 100990, 100990, 100940, 100920, 
    100880, 100850, 100820, 100770, 100730, 100700, 100670, 100630, 100610, 
    100590, 100570, 100520, 100500, 100510, 100520, _, 100570, 100560, 
    100570, 100590, 100610, 100630, 100620, 100630, 100620, 100620, 100620, 
    100610, 100640, 100630, 100640, 100640, 100630, 100610, 100580, 100560, 
    100550, 100550, 100560, _, 100550, 100550, 100550, 100550, 100550, 
    100540, 100530, 100520, 100510, 100500, _, 100520, 100520, 100530, 
    100530, 100550, 100560, 100570, 100580, 100590, 100590, 100600, 100620, 
    100630, 100650, 100660, _, 100710, 100720, 100750, 100760, 100770, 
    100790, 100800, 100830, 100860, 100880, 100910, 100930, 100950, 100980, 
    101010, 101020, 101040, 101060, 101090, 101110, _, 101170, 101200, 
    101220, 101220, 101240, 101270, 101280, 101290, 101290, 101300, 101320, 
    101340, 101360, 101380, 101420, 101420, 101440, 101450, 101450, 101450, 
    101470, 101480, 101490, 101520, 101520, 101510, 101500, 101490, 101480, 
    101460, 101450, 101440, 101420, 101400, 101370, 101360, 101350, 101340, 
    101300, 101250, 101210, 101170, 101160, 101120, 101090, 101070, 101050, 
    101040, 101030, 101020, 100980, 100950, 100930, 100920, 100920, 100910, 
    100890, 100890, 100900, 100920, 100940, 100960, 100970, 100970, 100990, 
    101020, 101040, 101040, 101040, 101060, 101070, _, 101080, 101120, 
    101120, 101130, 101150, 101160, 101160, 101160, 101160, 101180, 101200, 
    101220, 101240, 101250, 101270, 101290, 101320, 101330, 101350, 101330, 
    101350, 101370, 101380, 101380, 101410, 101430, 101450, 101460, 101480, 
    101490, 101510, 101550, 101560, 101560, 101590, 101620, 101620, 101650, 
    101660, 101680, 101720, 101740, 101770, 101780, 101770, 101760, 101770, 
    101800, 101810, 101830, 101850, 101860, 101860, 101880, 101890, 101890, 
    101890, 101900, 101900, 101920, 101940, 101970, 102000, 102020, 102010, 
    102010, 102020, 101970, 101940, 101900, 101870, 101870, 101870, 101860, 
    101830, 101880, 101860, 101860, 101850, 101840, 101820, 101780, 101760, 
    101760, 101740, 101710, 101680, 101640, 101640, 101610, 101570, 101530, 
    101510, 101480, 101460, 101440, 101360, 101300, 101250, 101230, 101200, 
    101160, 101130, 101060, 100990, 100970, 100910, 100880, 100850, 100850, 
    100800, 100780, 100800, 100800, 100840, 100840, 100850, 100850, 100860, 
    100870, 100880, 100880, 100850, 100810, 100780, 100760, 100730, 100650, 
    100590, 100530, 100480, 100380, 100310, 100290, 100210, 100120, 100070, 
    99980, 99870, 99760, 99670, 99590, 99580, 99710, 99780, 99820, 99850, 
    99880, 99900, 99920, 99930, 99910, 99900, 99860, 99820, 99730, 99670, 
    99600, 99540, 99470, 99300, 99150, 99040, 99000, 98980, 97980, 99010, 
    99100, 99180, 99250, 99330, 99410, 99470, 99540, 99610, 99670, 99750, 
    99820, 99880, 99950, 100000, 100090, 100140, 100190, 100220, 100280, 
    100280, 100290, 100300, 100300, 100270, 100240, 100230, 100240, 100260, 
    100290, 100290, 100270, 100290, 100260, 100210, 100160, 100130, 100110, 
    100100, 100090, 100110, 100110, 100120, 100130, 100180, 100190, 100250, 
    100330, 100390, 100460, 100510, 100560, 100610, 100670, 100720, 100770, 
    100780, 100800, 100770, 100760, 100770, 100710, 100650, 100560, 100470, 
    100380, 100290, 100170, 100050, 99900, 99740, 99560, 99410, 99300, 99200, 
    99170, 99160, 99160, 99200, 99280, 99370, 99500, 99610, 99740, 99850, 
    99980, 100100, 100210, 100320, 100420, 100530, 100620, 100720, 100790, 
    100860, 100950, 101030, 101070, 101130, 101170, 101230, 101260, 101290, 
    101280, 101280, 101270, 101290, 101290, 101280, 101260, 101270, 101260, 
    101220, 101200, 101170, 101120, 101040, 100930, 100830, 100690, 100590, 
    100530, 100470, 100420, 100390, 100370, 100380, 100410, 100440, 100470, 
    100490, 100530, 100590, 100650, 100730, 100810, 100900, 100970, 101060, 
    101120, 101190, 101260, 101310, 101380, 101450, 101510, 101580, 101650, 
    101700, 101730, 101770, 101810, 101800, 101780, 101760, 101710, 101660, 
    101590, 101510, 101470, 101410, 101370, 101320, 101290, 101290, 101290, 
    101250, 101360, 101430, 101550, 101660, 101750, 101870, 101900, 102030, 
    102110, 102210, 102280, _, 102360, 102380, 102430, 102480, 102540, 
    102540, 102530, 102550, 102590, 102590, 102580, 102540, _, 102440, 
    102390, 102340, 102290, 102250, 102200, 102150, 102100, 102040, 101980, 
    101910, 101820, 101780, 101740, 101710, 101660, 101630, 101610, 101570, 
    101520, 101500, 101450, 101390, 101360, 101320, 101300, 101300, 101250, 
    101270, 101250, 101220, 101160, 101120, 101120, 101060, 100990, 100950, 
    100970, 100990, 100990, 100990, 100990, 100970, 100980, 100960, 100940, 
    100940, 100900, 100870, 100850, 100820, 100760, 100710, 100630, 100540, 
    100450, 100400, 100310, 100240, 100150, 100010, 99950, 99910, 99930, 
    99960, 99980, 99920, 99910, 99890, 99900, 99950, 99940, 99940, 99950, 
    99960, 99970, 99960, 99960, 99950, 99970, _, 99960, 99960, 99980, 99980, 
    100000, 100020, _, 100020, 100030, 100010, 100010, 100010, 99990, 99950, 
    99930, 99910, 99900, 99880, _, 99850, 99820, 99800, 99770, 99740, 99720, 
    99680, 99670, 99670, 99680, 99680, 99670, 99670, 99660, 99650, 99680, 
    99680, 99700, 99710, 99730, 99720, 99740, 99760, 99780, 99820, 99850, 
    99870, 99920, 99960, 99990, 100000, 100010, 100030, 100060, 100080, 
    100100, 100080, 100090, 100070, 100050, 100040, 99990, 99940, 99880, 
    99790, 99770, 99750, 99710, 99670, 99660, 99660, 99670, 99670, 99700, 
    99720, 99760, 99780, 99840, 99900, 99950, 100000, 100060, 100120, 100160, 
    100210, 100250, 100290, 100330, 100350, _, 100450, _, 100510, 100540, 
    100560, 100580, 100580, 100580, 100600, 100600, 100600, 100600, 100630, 
    100620, 100630, 100650, 100670, 100680, 100690, 100710, 100730, 100750, 
    100780, 100810, 100850, 100900, 100930, 100980, 101020, 101070, 101110, 
    101140, 101180, 101180, 101190, 101230, 101250, 101270, 101350, 101390, 
    101420, 101450, 101450, 101440, 101400, 101360, 101320, 101270, 101240, 
    101200, 101150, 101070, 100980, 100900, 100840, 100760, 100690, 100630, 
    100590, 100550, 100500, 100460, 100430, 100400, 100380, 100380, 100380, 
    100380, 100400, 100430, 100450, 100480, 100520, 100560, 100580, 100640, 
    100680, 100740, 100800, 100870, 100890, 100920, 100930, 100970, 100970, 
    101010, 101000, 100970, 100920, 100890, 100820, 100740, 100650, 100570, 
    100490, 100390, 100300, 100250, 100240, 100230, 100220, 100220, 100230, 
    100270, 100300, 100350, 100410, 100490, 100560, 100650, 100710, 100780, 
    100830, 100900, 100950, 101020, 101090, 101150, 101210, 101270, 101310, 
    101310, 101340, 101370, 101410, 101430, 101410, 101370, 101320, 101290, 
    101290, 101310, 101270, 101250, 101270, _, 101250, 101220, 101150, 
    101080, 101020, 100930, 100860, _, _, 100690, _, 100610, 100590, 100590, 
    100630, 100640, 100680, 100720, 100760, 100800, 100860, 100910, 100970, 
    101040, 101090, 101110, 101140, 101190, 101210, 101230, 101240, 101260, 
    101270, 101310, 101310, 101310, 101310, 101310, 101310, 101310, 101390, 
    101460, 101490, 101530, 101560, 101600, 101640, 101680, 101720, 101750, 
    101730, 101710, 101720, 101730, 101730, 101740, 101750, 101760, 101800, 
    101830, 101860, 101900, 101930, 101960, 102020, 102070, 102120, 102160, 
    102220, 102260, 102260, 102290, 102290, 102290, 102290, 102270, 102230, 
    102210, _, _, 102100, 102050, 102010, 101950, 101900, 101800, 101740, 
    101650, 101550, 101440, 101350, 101230, 101130, 101050, 100950, 100840, 
    100740, 100660, 100530, 100440, 100370, 100290, 100250, 100220, 100190, 
    100170, 100170, 100150, 100140, 100160, 100180, 100180, 100200, 100220, 
    100230, 100240, 100260, 100280, 100290, 100310, 100340, 100280, 100280, 
    100260, 100260, 100250, 100230, 100220, 100200, 100160, 100130, 100100, 
    100060, 100040, 100020, 99980, 99950, 99940, 99920, 99910, 99900, 99890, 
    99880, 99890, 99880, 99870, 99850, 99850, 99850, 99850, 99850, 99850, 
    99850, 99820, 99800, 99780, 99770, 99760, 99750, 99720, 99710, 99700, 
    99680, 99710, 99710, 99710, 99700, 99710, 99740, 99750, 99780, 99790, 
    99820, 99850, 99880, 99930, 99970, 100010, 100050, 100090, 100160, 
    100210, 100270, 100340, 100420, 100480, 100550, 100620, 100710, 100780, 
    100850, 100910, 100980, 101050, 101080, 101120, 101130, 101160, 101210, 
    101230, 101240, 101290, 101320, 101320, 101320, 101350, 101340, 101350, 
    101360, 101360, 101370, 101360, 101360, _, 101350, 101350, 101360, 
    101370, 101340, 101330, 101320, 101300, 101250, 101230, 101230, 101190, 
    101180, 101130, 101120, 101110, 101080, 101030, 101010, 100950, 100920, 
    100930, 100900, 100880, 100840, 100820, 100830, 100790, 100750, 100730, 
    100700, 100670, 100650, 100600, 100580, 100540, 100530, 100490, 100470, 
    100480, 100450, 100390, 100340, 100320, 100270, 100210, 100170, 100100, 
    100070, 100020, 99970, 99890, 99820, 99760, 99720, 99700, 99650, 99630, 
    99630, 99600, 99570, 99570, 99570, 99600, 99630, 99670, 99700, 99730, 
    99790, 99860, 99930, _, 100060, 100140, 100200, 100270, 100330, 100360, 
    100410, 100480, 100530, 100580, 100640, 100710, 100760, 100810, 100860, 
    100910, 100950, 100980, 101040, 101050, 101100, 101130, 101170, 101200, 
    101220, 101230, 101240, 101260, 101270, 101270, 101270, 101250, 101260, 
    101260, 101280, 101280, 101280, 101290, 101290, 101280, 101280, 101280, 
    101280, 101290, 101300, 101300, 101290, 101310, 101310, 101310, 101300, 
    101330, 101340, 101350, 101360, 101380, 101380, 101390, 101390, 101380, 
    101400, 101400, 101400, 101410, 101420, 101400, 101380, 101370, 101370, 
    101370, 101340, 101340, 101340, 101320, 101290, 101270, _, 101190, 
    101170, 101130, 101110, 101090, 101090, 101040, 101000, 100940, 100890, 
    100880, 100860, 100790, 100720, 100660, 100630, 100600, 100580, 100540, 
    100480, 100470, 100440, 100410, 100350, 100330, 100280, 100240, 100190, 
    100140, 100080, 100030, 99960, 99920, 99880, 99840, 99790, 99740, 99700, 
    99660, 99630, 99600, 99590, 99580, 99590, 99580, 99570, 99580, 99590, 
    99600, 99600, 99620, 99630, 99630, 99640, 99680, 99710, 99730, 99760, 
    99780, 99830, 99850, 99880, 99900, 99920, 99940, 99990, 100030, 100070, 
    100110, 100140, 100190, 100220, 100250, 100290, 100310, 100350, 100390, 
    100430, 100480, 100520, 100570, 100590, 100630, 100650, 100690, 100720, 
    100740, 100740, 100720, 100760, 100770, 100770, 100760, 100710, 100640, 
    100600, 100560, 100430, 100340, 100220, 100180, 100160, 100040, 99980, 
    99890, 99860, 99880, 99870, 99890, 99840, 99800, 99810, 99810, 99800, 
    99790, 99750, 99750, 99730, 99730, _, 99680, 99600, 99600, 99590, 99590, 
    99560, 99490, 99440, 99390, 99360, 99340, 99310, 99290, 99280, 99260, 
    99280, 99320, 99410, 99480, 99560, 99650, 99740, 99800, 99890, 99960, 
    100010, 100090, 100110, 100140, 100200, 100250, 100310, 100370, 100430, 
    100510, 100560, 100610, 100680, 100730, 100790, 100820, 100860, 100920, 
    100970, 100990, 101000, 101010, 101020, 101010, 101000, 100950, 100960, 
    100930, 100900, 100870, 100840, 100800, 100740, 100690, 100630, 100560, 
    100460, 100400, 100350, 100310, 100260, 100270, 100190, 100100, 100000, 
    99890, 99810, 99750, 99700, 99600, 99560, 99530, 99500, 99460, 99430, 
    99410, 99390, 99370, 99370, 99380, 99400, 99420, 99460, 99510, 99570, 
    99640, 99700, 99770, 99840, 99920, 100000, 100070, 100120, 100170, 
    100220, 100280, 100310, 100350, 100400, 100440, 100470, 100490, 100530, 
    100560, 100600, 100600, 100610, 100640, 100700, 100720, 100760, 100790, 
    100810, 100840, 100870, 100900, 100910, 100940, 100930, 100960, 100970, 
    100980, 100990, 100990, 101010, 101020, 101020, 101030, 101010, 101040, 
    101040, 101060, 101050, 101050, 101070, 101090, 101100, 101090, 101070, 
    101070, 101070, 101070, 101040, 101030, 101030, 101040, 101040, 101030, 
    101030, 101010, 101010, 101000, 100980, 100970, 100960, 100950, 100940, 
    100980, 100990, 100950, 100940, 100920, 100900, 100870, 100840, 100810, 
    100720, 100690, 100640, 100620, 100570, 100540, 100480, 100440, 100410, 
    100370, 100350, 100290, 100200, 100170, 100130, 100080, 100020, 99990, 
    99960, 99900, 99850, 99800, 99800, 99770, 99720, 99690, 99690, 99690, 
    99700, 99700, 99690, 99690, 99690, 99690, 99700, 99710, 99710, 99720, 
    99730, 99760, 99770, 99780, 99800, 99790, 99770, 99730, 99700, 99670, 
    99640, 99640, 99600, 99570, 99540, 99510, 99450, 99420, 99390, 99350, 
    99310, 99250, 99210, 99170, 99140, 99110, 99060, _, 98990, 98950, 98950, 
    98940, 98910, 98900, 98900, 98920, 98920, 98960, 98990, 99000, 99020, 
    99040, 99070, 99090, 99100, 99140, 99170, 99240, 99320, 99380, 99440, 
    99500, 99510, 99550, 99600, 99630, 99660, 99700, 99740, 99770, 99830, 
    99870, 99910, 99940, 99980, 100010, 100040, 100060, 100090, 100110, 
    100120, 100160, 100180, 100220, 100240, 100260, 100270, 100280, 100290, 
    100290, 100290, 100300, 100320, 100320, 100340, 100370, 100370, _, 
    100420, 100400, 100400, 100410, 100410, 100410, 100420, 100450, 100460, 
    100510, 100500, _, 100560, 100560, 100580, 100590, 100590, 100600, 
    100620, 100630, 100680, 100690, 100730, 100730, 100780, 100780, 100840, 
    100870, 100900, 100930, 100930, 100940, 100950, 100970, 100960, 100950, 
    100950, 100980, 100990, 100970, 100980, 100970, 100990, 101020, 101050, 
    101040, 101060, 101050, 101050, 101040, 101010, 100980, 100960, 100920, 
    100890, 100860, 100830, 100790, 100750, 100680, 100620, 100560, 100490, 
    100430, 100350, 100300, 100260, 100280, 100300, 100350, 100450, 100520, 
    100610, 100670, 100730, 100780, 100830, 100880, 100950, 101000, 101070, 
    101140, 101180, 101240, 101280, 101320, 101350, 101360, 101380, 101380, 
    101400, 101410, 101410, 101440, 101420, 101410, 101410, 101430, 101410, 
    101410, 101390, 101390, 101410, 101410, 101430, 101410, 101400, 101440, 
    101430, 101420, 101410, 101400, 101410, 101410, 101400, 101390, 101360, 
    101370, 101380, 101380, 101380, 101360, 101350, 101360, 101330, 101310, 
    101300, 101300, 101310, 101290, 101300, 101290, 101280, 101250, 101260, 
    101260, 101260, 101250, 101250, 101250, 101250, 101240, 101250, 101250, 
    101240, 101220, 101210, 101200, 101180, 101160, 101180, 101190, 101190, 
    101190, 101200, 101200, 101200, 101210, 101170, 101140, 101140, 101130, 
    101130, 101150, 101160, 101180, 101170, 101180, 101200, 101180, 101180, 
    101200, 101200, 101220, 101220, 101250, 101260, 101260, 101280, 101280, 
    101300, 101300, 101280, 101270, 101240, 101240, 101230, 101220, 101210, 
    101220, 101200, 101190, 101180, 101160, 101130, 101070, 101030, 101020, 
    101020, _, 100970, 100970, 100950, 100950, 100970, 100980, 100980, 
    100960, 100920, 100900, 100870, 100830, 100780, 100750, 100710, 100660, 
    100600, 100540, 100510, 100470, 100410, 100340, 100320, 100290, 100260, 
    100240, 100210, 100240, 100260, 100250, 100270, 100260, 100270, 100270, 
    100300, 100360, 100350, 100320, 100310, 100330, 100360, 100370, 100400, 
    100420, 100460, 100490, 100530, 100570, 100610, 100620, 100660, 100660, 
    100660, 100670, 100640, 100640, 100620, 100590, 100540, 100520, 100500, 
    100480, 100430, 100390, 100340, 100280, 100210, 100170, 100120, 100070, 
    100090, 100090, 100130, 100150, 100090, 100050, 100020, 99970, 99910, 
    99870, 99810, 99810, 99780, 99780, 99830, 99810, 99870, 99900, 99990, 
    100030, 100120, 100200, 100260, 100310, 100370, 100430, 100510, 100560, 
    100570, 100570, 100550, 100560, 100570, 100580, 100600, 100630, 100660, 
    100690, 100730, 100760, 100790, 100820, 100810, 100840, 100820, 100820, 
    100790, 100730, 100680, 100620, 100530, 100420, 100360, 100280, 100210, 
    100160, 100120, 100120, 100100, 100110, 100140, 100170, 100180, 100210, 
    100250, 100280, 100300, 100330, 100340, 100370, 100370, 100410, 100450, 
    100510, 100550, 100620, 100670, 100710, 100760, 100800, 100810, 100820, 
    100830, 100820, 100810, 100810, 100810, 100780, 100740, 100720, 100690, 
    100620, 100560, 100470, 100400, 100330, 100260, 100240, 100200, 100150, 
    100130, 100110, 100090, 100100, 100110, 100130, 100170, 100210, 100250, 
    100300, 100360, 100380, 100470, 100490, 100530, 100580, 100600, 100610, 
    100630, 100640, 100650, 100650, 100650, 100650, 100630, 100640, 100630, 
    100610, 100600, 100560, 100530, 100510, 100480, 100450, 100470, 100470, 
    100470, 100430, 100390, 100400, 100360, 100330, 100290, 100240, 100240, 
    100280, 100290, 100330, 100370, 100410, 100470, 100520, 100540, 100570, 
    100640, 100710, 100750, 100800, 100820, 100880, 100900, 100940, 101010, 
    101040, 101060, 101060, 101080, 101100, 101130, 101150, 101180, 101180, 
    101210, 101220, 101230, 101240, 101260, 101290, 101310, 101340, 101360, 
    101400, 101450, 101490, 101540, 101580, 101620, 101660, 101680, 101700, 
    101730, 101710, 101720, 101710, 101720, 101720, 101680, 101680, 101670, 
    101640, 101610, 101590, 101560, 101550, 101550, 101560, 101600, 101610, 
    101600, 101610, 101630, 101650, 101610, 101610, 101590, 101560, 101550, 
    101490, 101450, 101380, 101300, 101220, 101180, 101100, 101000, 100920, 
    100850, 100720, 100650, 100570, 100500, 100450, 100370, 100370, 100380, 
    100370, 100360, 100320, 100260, 100240, 100190, 100150, 100120, 100070, 
    100050, 100030, 100040, 100050, 100070, 100070, 100070, 100060, 100050, 
    100070, 100090, 100120, 100160, 100190, 100230, 100280, 100320, 100350, 
    100380, 100410, 100450, 100490, _, 100570, _, 100670, 100730, 100790, 
    100830, 100860, 100880, 100920, 100950, 100980, 101000, 101020, 101030, 
    101040, 101020, 101010, 100960, 100940, 100900, 100870, 100860, 100820, 
    100780, 100750, 100730, 100710, 100670, 100610, 100570, 100500, 100470, 
    100440, 100410, 100400, 100400, 100380, 100350, 100360, 100340, 100330, 
    100290, 100280, 100250, 100220, 100210, 100190, 100170, 100160, 100190, 
    100160, 100150, _, _, 100060, 100050, 100040, 99990, 100000, 99970, 
    99970, 99940, 99910, 99880, 99850, 99820, 99790, 99810, 99820, 99840, 
    99850, 99870, 99910, 99950, 100010, 100100, 100160, 100180, 100220, 
    100250, 100290, 100380, 100430, 100460, 100520, 100550, 100610, 100650, 
    100670, 100680, 100690, 100720, 100720, 100730, 100710, 100690, 100660, 
    100650, 100630, 100580, 100550, 100520, 100460, 100440, 100420, 100410, 
    100380, 100370, 100400, 100420, 100430, 100440, 100420, 100410, 100390, 
    100390, 100430, 100490, 100530, 100630, 100740, 100810, 100860, 100860, 
    100910, 100940, 100960, 100950, 100980, 100980, 101020, 101030, 101060, 
    101080, 101110, 101140, 101140, 101150, 101150, 101180, 101160, 101210, 
    101290, 101360, 101470, _, 101550, 101610, 101630, 101620, 101660, 
    101650, 101640, 101600, 101550, 101480, 101410, 101350, 101290, 101240, 
    101220, 101230, 101210, 101210, 101240, 101260, 101270, 101320, 101320, 
    101350, 101410, 101420, 101450, 101470, 101500, 101500, 101530, 101530, 
    101530, 101550, 101560, 101540, 101520, 101520, 101510, 101520, 101520, 
    101530, 101510, 101520, 101550, 101610, 101650, 101660, 101690, 101720, 
    101740, 101730, 101740, 101780, 101790, 101840, 101890, 101930, 101940, 
    101980, 102010, 102040, 102060, 102070, 102070, 102090, 102080, 102070, 
    102070, 102080, 102090, 102090, 102090, 102110, 102100, 102100, 102090, 
    102050, 102030, 102030, 102030, 102030, 102030, 102010, 102000, 101980, 
    101980, 101970, 101940, 101900, 101870, 101850, 101850, 101870, 101860, 
    101840, 101830, 101790, 101760, 101750, 101710, 101650, 101670, 101680, 
    101730, 101740, 101740, 101750, 101730, 101730, 101730, 101730, 101730, 
    101740, 101740, 101700, 101690, 101700, 101730, 101750, 101720, 101710, 
    101720, 101700, 101670, 101620, 101630, 101640, 101630, 101640, 101620, 
    101590, 101580, 101590, 101580, 101570, 101590, 101590, _, 101620, 
    101620, 101630, 101630, _, 101650, 101700, 101730, 101760, 101800, 
    101830, 101830, 101860, 101860, 101870, 101860, 101870, 101870, 101860, 
    101860, 101870, 101850, 101840, 101820, 101800, 101800, 101790, _, 
    101790, 101760, 101750, 101730, 101700, 101680, 101650, 101630, 101590, 
    101560, 101540, 101510, 101510, 101480, 101460, 101430, 101410, 101380, 
    101350, 101320, 101280, 101270, 101260, 101250, 101230, 101210, 101200, 
    101180, 101140, 101130, 101100, 101090, 101070, 101070, 101070, 101060, 
    101070, 101040, 101070, 101060, 101070, 101080, 101070, _, 101100, 
    101130, 101160, 101190, _, 101220, _, 101240, 101240, 101250, 101220, 
    101190, 101210, 101190, 101190, 101190, 101190, 101160, 101140, 101120, 
    101080, 101050, 100990, 100910, 100890, 100850, 100840, 100810, 100780, 
    100750, 100720, 100700, 100670, 100620, 100590, 100570, 100500, 100480, 
    100430, 100380, 100360, 100280, 100230, 100200, 100080, 100110, 100080, 
    100040, 100020, 99980, 99910, 99870, 99810, 99780, 99730, 99730, 99710, 
    _, 99640, 99610, 99600, 99630, 99600, 99660, 99720, 99680, 99710, 99770, 
    99770, 99780, 99820, 99810, 99820, 99850, 99880, 99910, 99940, 99970, 
    99990, 100010, 100020, 100030, 100050, 100070, 100100, 100130, 100150, 
    100180, 100200, 100210, 100220, 100220, 100240, 100240, 100230, 100240, 
    100260, 100280, 100290, _, 100300, 100310, 100340, 100350, 100360, 
    100360, 100390, 100400, 100410, 100440, 100460, 100510, 100540, 100560, 
    100580, 100600, 100640, 100640, 100650, 100670, 100700, 100730, 100770, 
    100790, 100820, 100850, 100860, 100880, 100890, 100910, 100930, 100940, 
    100940, 100960, 100990, 101020, 101030, 101050, 101050, 101060, 101070, 
    101060, 101060, 101030, 101040, 101050, 101040, 101060, 101040, 101030, 
    101020, 101010, 100990, 100960, 100950, 100930, 100930, 100920, 100910, 
    100910, 100900, 100870, 100880, 100880, 100860, 100830, 100820, 100810, 
    100800, 100790, 100780, 100800, 100800, 100800, 100800, 100800, 100780, 
    100770, 100750, 100760, 100780, 100780, 100790, 100800, 100780, 100780, 
    100780, 100780, 100770, 100780, 100770, 100750, 100740, 100720, 100730, 
    100720, 100730, 100720, 100710, 100710, 100700, 100700, 100690, _, 
    100680, 100670, 100640, 100640, 100630, 100660, 100650, 100670, 100670, 
    100670, 100660, 100650, 100640, 100640, 100640, 100660, 100660, 100680, 
    100680, 100690, 100680, 100680, 100680, 100670, 100660, 100650, 100650, 
    100660, 100680, 100690, 100710, 100700, 100720, 100720, 100720, 100720, 
    100720, 100730, 100740, _, 100760, 100780, 100780, 100790, 100800, 
    100810, 100810, 100820, 100840, 100850, 100850, 100870, 100900, 100910, 
    100930, 100950, 100980, 100970, 100980, 100990, 101010, 101020, 101030, 
    101040, 101050, 101060, 101040, 101030, 101020, 101010, 101020, 100980, 
    100960, 100940, 100960, 100940, 100920, 100900, 100890, 100860, 100830, 
    100790, 100740, 100690, 100650, 100590, 100550, 100520, 100490, 100410, 
    _, 100310, 100250, 100180, 100130, 100050, 99970, 99870, 99790, 99710, 
    99580, 99470, 99410, 99290, 99150, 99020, 98860, 98690, 98550, 98470, 
    98450, 98390, 98370, 98340, 98360, 98340, 98330, 98330, 98300, 98310, 
    98310, 98300, 98330, 98340, 98340, 98360, 98360, 98360, 98350, 98360, 
    98360, 98350, 98360, 98370, 98380, 98380, 98400, 98400, 98430, 98430, 
    98450, 98460, 98470, 98470, 98470, 98480, 98480, 98490, 98510, 98530, 
    98540, 98540, 98540, 98550, 98550, 98540, 98550, 98550, 98580, 98600, 
    98610, 98630, 98640, 98650, 98680, 98720, _, 98800, 98830, 98860, 98920, 
    98970, 99020, 99040, 99080, 99130, 99140, 99160, 99170, 99190, 99260, 
    99300, 99360, 99380, 99440, 99470, 99510, 99550, 99580, 99630, 99670, 
    99690, 99730, 99750, 99810, 99840, 99860, 99900, 99930, 99930, 99930, 
    99960, 99990, 100010, 100010, 100020, 100040, 100060, 100100, 100120, 
    100150, 100190, 100190, 100220, 100270, 100350, 100360, 100380, 100420, 
    100450, 100480, 100510, 100550, 100560, 100580, 100600, 100610, 100650, 
    100670, 100710, 100720, 100760, 100790, 100820, 100830, 100870, 100890, 
    100870, 100880, 100910, 100920, 100920, 100920, 100930, 100940, 100960, 
    100970, 100960, 100960, 100960, 100960, 100960, 100970, 100980, 100980, 
    101000, 101000, 101000, 101020, 101030, 101030, 101020, 101030, 101040, 
    101030, 101040, 101050, 101060, 101070, 101070, 101060, 101060, 101030, 
    100990, 100960, 100960, 100940, 100910, 100860, 100810, 100740, 100720, 
    100680, 100630, 100630, 100530, 100500, 100420, 100350, 100300, 100230, 
    100180, 100140, 100090, 100040, 99990, 99930, 99910, 99880, 99850, 99830, 
    99820, 99810, 99820, 99830, 99840, 99870, 99900, 99920, 99960, 100010, 
    100050, 100090, 100130, 100180, 100240, 100270, 100330, 100360, 100390, 
    100400, 100430, 100430, 100450, 100480, 100500, 100510, 100510, 100520, 
    100530, 100540, 100550, 100560, 100570, 100570, 100580, 100600, 100600, 
    100600, 100610, 100620, 100640, 100660, 100690, 100700, 100720, 100750, 
    100780, 100820, 100860, 100900, 100930, 100990, 101030, 101060, 101090, 
    101120, 101150, 101180, 101220, 101250, 101270, 101270, 101280, 101280, 
    _, 101260, 101240, 101200, 101170, 101130, 101110, 101070, 101050, 
    101040, 101090, 101090, 101090, 101090, 101070, 101050, 101030, 101000, 
    100930, 100870, 100810, 100710, 100680, 100640, 100590, 100520, 100440, 
    100360, 100260, 100150, 100060, 99950, 99850, 99740, 99590, 99480, 99310, 
    99120, 98950, 98790, 98620, 98600, 98790, 98940, 98970, 99050, 99030, 
    98970, 98960, 98960, 99050, 99060, 99020, 99060, 99100, _, 99270, 99400, 
    99500, 99620, 99700, 99770, 99920, 100070, 100200, 100320, 100390, 
    100420, 100540, 100590, 100700, 100770, 100850, 100870, 100880, 100890, 
    100900, 100880, 100860, 100860, 100840, 100810, 100820, 100840, 100870, 
    100890, 100880, 100860, 100830, 100820, 100820, 100780, 100770, 100720, 
    100710, 100680, 100640, 100560, 100500, 100420, 100390, 100330, 100280, 
    100260, 100250, 100270, 100260, 100270, _, 100230, 100220, 100190, 
    100150, 100130, 100090, 100070, 100050, 100020, 100010, 100010, 100010, 
    100000, 99970, 99900, 99850, 99820, 99790, 99710, 99660, 99530, 99410, 
    99290, 99170, 99070, 99000, 98960, 98950, 98980, 99050, 99110, 99190, 
    99280, 99360, 99470, 99560, 99660, 99760, 99850, 99950, 100060, 100170, 
    100270, 100370, 100480, 100570, 100670, 100770, 100870, 100950, 101000, 
    101080, 101130, 101210, 101290, 101370, 101450, 101520, 101570, 101600, 
    101640, 101690, 101710, 101720, 101750, 101770, 101790, 101780, 101770, 
    101730, _, _, 101580, 101510, 101430, 101350, 101290, 101240, 101190, 
    101120, 101060, 100980, 100940, 100920, 100850, 100860, 100920, 100950, 
    100990, 101020, 101050, 101070, 101130, 101180, 101230, 101270, 101320, 
    101370, 101410, 101460, 101520, 101580, 101640, 101690, 101740, 101780, 
    101810, 101850, 101870, 101900, 101900, 101910, 101910, 101860, 101860, 
    101840, 101810, 101760, 101710, 101650, 101630, 101580, 101550, 101490, 
    101450, 101440, 101430, 101440, 101430, 101440, 101470, 101460, 101460, 
    101450, 101450, 101440, 101440, 101470, 101440, 101440, 101420, 101390, 
    101380, 101360, 101330, 101300, 101270, 101260, 101220, 101200, 101200, 
    101190, 101180, 101180, 101200, 101200, 101190, 101210, 101210, 101210, 
    101240, 101250, 101280, 101310, 101340, 101380, 101420, 101450, 101480, 
    101500, 101520, 101540, 101550, 101550, 101560, 101570, 101560, 101550, 
    101540, 101570, 101600, 101600, 101580, 101560, 101530, 101540, 101530, 
    101540, 101540, 101520, 101500, 101480, 101480, 101490, 101480, 101450, 
    101430, 101440, 101460, 101460, 101480, 101480, 101470, 101440, 101440, 
    101430, 101420, 101420, 101380, 101350, 101350, 101330, 101290, 101290, 
    101250, 101230, 101190, 101170, 101150, 101120, 101080, 101040, 101010, 
    100970, 100960, 100920, 100880, 100860, 100850, 100820, 100790, 100760, 
    100750, 100720, 100680, 100670, 100670, 100710, 100700, 100650, 100650, 
    100680, 100670, 100690, 100680, 100710, 100720, 100710, 100720, 100730, 
    100730, 100720, 100720, 100700, 100670, 100640, 100600, 100580, 100570, 
    100560, 100550, 100540, 100530, 100520, 100510, 100490, 100470, 100430, 
    100400, 100370, 100340, 100320, 100310, 100300, 100270, 100270, 100250, 
    100240, 100240, 100250, 100230, 100250, 100300, 100330, 100360, 100400, 
    100410, 100440, 100470, 100480, 100490, 100490, 100500, 100500, 100520, 
    100540, 100570, 100570, 100590, 100580, 100560, 100560, 100580, 100590, 
    100590, 100590, 100610, 100650, 100700, 100750, 100790, 100790, 100810, 
    100840, 100860, 100890, 100920, 100960, 101000, 101030, 101070, 101110, 
    101130, 101150, 101170, 101200, 101210, 101230, 101270, 101280, 101310, 
    101330, 101360, 101370, 101380, 101410, 101420, 101420, 101430, 101430, 
    101460, 101460, 101480, 101490, 101490, 101510, 101500, 101480, 101460, 
    101470, 101450, 101450, 101450, 101460, 101420, 101410, 101390, 101370, 
    101340, 101300, 101240, 101230, 101210, 101180, 101180, 101160, 101150, 
    101150, 101140, 101130, 101100, 101080, 101090, 101090, 101090, 101090, 
    101090, 101110, 101110, 101110, 101110, 101140, 101130, 101130, 101140, 
    101150, 101160, 101180, 101210, 101230, 101260, 101270, 101280, 101290, 
    101290, 101300, 101330, 101330, 101350, 101370, 101380, 101370, 101370, 
    101360, 101350, 101360, 101340, 101330, 101320, 101330, 101330, 101330, 
    101320, 101310, 101280, 101280, 101220, 101190, 101180, 101140, 101140, 
    101100, 101080, 101060, 101040, 100990, 100970, 100970, 100930, 100910, 
    100910, 100880, 100860, 100830, 100800, 100810, 100790, 100760, 100690, 
    100680, 100700, 100680, 100650, 100640, 100600, 100560, 100530, 100500, 
    100490, 100520, 100510, 100500, 100510, 100510, 100460, 100430, 100430, 
    100430, 100440, 100430, 100420, 100400, 100400, 100390, 100390, 100400, 
    100420, 100440, 100440, 100440, 100450, 100430, 100380, 100380, 100350, 
    100320, 100340, 100360, 100340, 100300, 100280, 100270, 100270, 100260, 
    100280, 100220, 100200, 100150, 100150, 100100, 100040, 99970, 99920, 
    99850, 99750, 99690, 99620, 99500, 99370, 99230, 99130, 99000, 98980, 
    98900, 98780, 98660, 98620, 98520, 98430, 98270, 98130, 98000, 97960, 
    97890, 97800, 97770, 97770, 97740, 97700, 97700, 97670, 97640, 97600, 
    97610, 97610, 97620, 97610, 97590, 97590, 97590, 97580, 97560, 97560, 
    97540, 97550, 97570, 97590, 97600, 97600, 97620, 97650, 97660, 97660, 
    97680, 97700, 97740, 97760, 97790, 97830, 97860, 97910, 97960, 97990, 
    98040, 98070, 98110, 98130, 98150, 98150, 98170, 98200, 98240, 98270, 
    98280, 98270, 98290, 98290, 98300, 98300, 98300, 98330, 98350, 98380, 
    98410, 98460, 98510, 98540, 98560, 98590, 98630, 98660, 98690, 98730, 
    98750, 98790, 98830, 98840, 98870, 98890, 98900, 98910, 98920, 98920, 
    98930, 98950, 98970, 98990, 99030, 99070, 99090, 99110, 99120, 99140, 
    99150, 99200, 99220, 99250, 99260, 99300, 99320, 99320, 99330, 99340, 
    99350, 99360, 99380, 99360, 99390, 99380, 99370, 99390, 99390, 99400, 
    99400, 99420, 99410, 99420, 99420, 99420, 99420, 99420, 99400, 99410, 
    99440, 99440, 99450, 99450, 99440, 99480, 99510, 99550, 99590, 99630, 
    99660, 99700, 99720, 99780, 99800, 99820, 99840, 99880, 99890, 99910, 
    99910, 99960, 99980, 100020, 100060, 100110, 100110, 100120, 100140, 
    100170, 100190, 100190, 100230, 100280, 100320, 100350, 100380, 100440, 
    100500, 100540, 100580, 100630, 100670, 100700, 100750, 100780, 100810, 
    100840, 100850, 100870, 100900, 100880, 100870, 100840, 100830, 100810, 
    100770, 100740, 100730, 100710, 100700, 100680, 100650, 100630, 100600, 
    100550, 100510, 100450, 100410, 100390, 100380, 100350, 100350, 100320, 
    100330, 100310, 100300, 100290, 100290, 100290, 100290, 100290, 100300, 
    100290, 100280, 100280, 100280, 100290, 100280, 100300, 100310, 100320, 
    100330, 100350, 100350, 100350, 100410, 100440, 100470, 100450, 100470, 
    100520, 100520, 100520, 100520, 100550, 100550, 100540, 100570, 100600, 
    100630, 100630, 100630, 100630, 100620, 100620, 100600, 100600, 100570, 
    100560, 100540, 100530, 100480, 100460, 100430, 100400, 100380, 100360, 
    100330, 100300, 100280, 100280, 100290, 100280, 100280, 100280, 100270, 
    100260, 100250, 100230, 100190, 100160, 100130, 100090, 100030, 100010, 
    99960, 99900, 99870, 99780, 99700, 99590, 99510, 99440, 99380, 99330, 
    99260, 99190, 99130, 99040, 98960, 98890, 98810, 98750, 98670, 98610, 
    98560, 98500, 98450, 98420, 98370, 98370, 98370, 98350, 98350, 98350, 
    98340, 98360, 98410, 98460, 98520, 98560, 98620, 98680, 98720, 98760, 
    98760, 98790, 98820, 98830, 98870, 98900, 98940, 98970, 98970, 98990, 
    99010, 99030, 99060, 99080, 99100, 99110, 99120, 99180, 99220, 99240, 
    99270, 99300, 99330, 99300, 99280, 99270, 99280, 99270, 99260, 99240, 
    99220, 99210, 99170, 99140, 99100, 99050, 99010, 98970, 98950, 98910, 
    98880, 98870, 98860, 98860, 98850, 98840, 98820, 98800, 98770, 98770, 
    98750, 98740, 98750, 98750, 98740, 98740, 98740, 98720, 98710, 98700, 
    98690, 98670, 98640, 98640, 98640, 98660, 98680, 98690, 98700, 98710, 
    98720, 98730, 98740, 98760, 98790, 98820, 98850, 98890, 98930, 98970, 
    99010, 99040, 99100, 99150, 99200, 99250, 99310, 99380, 99420, 99510, 
    99590, 99660, 99740, 99810, 99870, 99950, 100010, 100050, 100140, 100210, 
    100280, 100360, 100430, 100500, 100550, 100570, 100620, 100660, 100660, 
    100690, 100740, 100780, 100850, 100920, 100990, 101060, 101110, 101150, 
    101210, 101270, 101320, 101360, 101390, 101430, 101470, 101500, 101530, 
    101560, 101570, 101570, 101540, 101500, 101490, 101500, 101520, 101520, 
    101530, 101560, 101590, 101620, 101630, 101650, 101630, 101640, 101640, 
    101630, 101630, 101610, 101570, 101540, 101500, 101440, 101400, 101350, 
    101290, 101290, 101210, 101180, 101100, 101030, 100990, 100930, 100830, 
    100720, 100660, 100600, 100490, 100380, 100270, 100140, 99990, 99900, 
    99770, 99670, 99570, 99360, 99270, 99080, 99020, 98950, 98930, 98840, 
    98780, 98690, 98640, 98570, 98510, 98440, 98410, 98420, 98480, 98540, 
    98610, 98750, 98810, 98870, 98880, 98920, 98980, 98970, 98980, 98960, 
    98970, 98960, 98930, 98890, 98880, 98880, 98890, 98890, 98890, 98920, 
    98940, 98960, 98980, 98980, 98990, 99000, 99020, 99010, 99020, 99030, 
    99030, 99030, 99030, 99020, 99040, 99020, 99050, 99070, 99080, 99100, 
    99140, 99190, 99270, 99320, 99380, 99420, 99460, 99530, 99590, 99650, 
    99720, 99770, 99830, 99890, 99930, 99980, 100020, 100060, 100090, 100120, 
    100130, 100150, 100170, 100170, 100190, 100200, 100220, 100220, 100210, 
    100200, 100200, 100170, 100130, 100110, 100080, 100030, 100010, 99980, 
    99950, 99910, 99900, 99870, 99840, 99790, 99760, 99730, 99690, 99670, 
    99670, 99690, 99700, 99690, 99700, 99700, 99710, 99730, 99740, 99760, 
    99800, 99830, 99850, 99890, 99930, 100000, 100050, 100100, 100150, 
    100200, 100260, 100320, 100360, 100420, 100480, 100550, 100620, 100690, 
    100740, 100810, 100880, 100910, 100940, 100950, 100980, 101010, 101010, 
    101020, 101060, 101050, 101030, 101010, 100980, 100950, 100910, 100860, 
    100810, 100790, 100780, 100700, 100670, 100640, 100590, 100520, 100430, 
    100320, 100220, 100120, 100040, 99930, 99840, 99720, 99620, 99540, 99460, 
    99350, 99280, 99180, 99050, 98960, 98950, 98870, 98810, 98760, 98710, 
    98650, 98590, 98530, 98520, 98470, 98390, 98350, 98270, 98220, 98170, 
    98140, 98080, 98040, 98010, 98000, 97960, 97950, 97940, 97930, 97930, 
    97930, 97980, 97990, 98030, 98060, 98120, 98160, 98180, 98190, 98220, 
    98270, 98310, 98360, 98390, 98450, 98540, 98580, 98630, 98720, 98820, 
    98920, 98980, 99100, 99210, 99300, 99400, 99510, 99670, 99800, 99940, 
    99990, 100070, 100120, 100250, 100300, 100380, 100420, 100510, 100540, 
    100620, 100670, 100740, 100740, 100810, 100840, 100890, 100930, 100960, 
    101000, 101060, 101090, 101110, 101130, 101170, 101200, 101230, 101250, 
    101290, 101320, 101310, 101330, 101400, 101400, 101450, 101460, 101480, 
    101490, 101510, 101540, 101570, 101580, 101630, 101660, 101710, 101710, 
    101750, 101810, 101870, 101920, 101960, 101980, 102010, 102030, 102050, 
    102090, 102120, 102150, 102190, 102220, 102260, 102280, 102310, 102360, 
    102400, 102450, 102500, 102550, 102620, 102690, 102750, 102780, 102810, 
    102850, 102870, 102930, 102960, 102960, 102990, 103010, 103040, 103020, 
    103000, 102990, 102970, 102950, 102900, 102890, 102870, 102810, 102780, 
    102690, 102710, 102690, 102670, 102610, 102560, 102530, 102470, 102440, 
    102420, 102360, 102300, 102240, 102200, 102150, 102070, 102040, 101980, 
    101910, 101830, 101760, 101710, 101660, 101580, 101510, 101470, 101410, 
    101350, 101290, 101170, 101110, 101020, 100930, 100860, 100780, 100650, 
    100560, 100490, 100420, 100360, 100290, 100170, 100090, 100010, 99940, 
    99890, 99860, 99820, 99820, 99850, 99920, 100000, 100080, 100130, 100190, 
    100230, 100250, 100240, 100240, 100270, 100370, 100480, 100610, 100740, 
    100830, 100890, 101030, 101170, 101220, 101340, 101430, 101560, 101700, 
    101790, 101890, 101980, 101980, 101970, 102010, 102000, 101950, 101910, 
    101870, 101820, 101780, 101740, 101700, 101650, 101640, 101620, 101550, 
    101510, 101450, 101370, 101300, 101240, 101180, 101140, 101110, 101090, 
    101070, 101030, 100990, 100980, 100950, 100920, 100930, 100930, 100940, 
    100940, 100940, 100940, 100940, 100960, 100960, 100950, 100980, 100980, 
    100990, 101010, 101020, 101070, 101130, 101160, 101220, 101260, 101300, 
    101330, 101370, 101400, 101420, 101450, 101470, 101510, 101520, 101540, 
    101590, 101630, 101620, 101650, 101680, 101700, 101730, 101770, 101790, 
    101820, 101860, 101920, 101920, 101940, 101960, 101980, 101980, 101990, 
    101980, 101980, 102010, 101990, 101980, 101960, 101930, 101910, 101840, 
    101810, 101780, 101700, 101650, 101620, 101580, 101540, 101510, 101500, 
    101480, 101460, 101470, 101410, 101390, 101320, 101290, 101290, 101290, 
    101250, 101250, 101210, 101170, 101130, 101080, 101010, 100940, 100870, 
    100790, 100700, 100600, 100550, 100540, 100500, 100440, 100440, 100410, 
    100380, 100310, 100240, 100210, 100150, 100070, 100010, 99980, 99950, 
    99890, 99870, 99810, 99770, 99720, 99690, 99690, 99690, 99740, 99780, 
    99820, 99830, 99890, 99920, 99960, 100010, 100100, 100100, 100130, 
    100210, 100260, 100340, 100360, 100420, 100470, 100530, 100530, 100550, 
    100600, 100610, 100640, 100670, 100680, 100730, 100830, 100890, 100950, 
    100980, 101030, 101090, 101120, 101190, 101250, 101310, 101410, 101470, 
    101550, 101610, 101680, 101730, 101810, 101850, 101900, 101940, 101930, 
    101950, 101970, 101990, 102020, 102070, 102150, 102220, 102280, 102330, 
    102370, 102390, 102400, 102420, 102450, 102510, 102510, 102530, 102540, 
    102570, 102590, 102610, 102620, 102630, 102660, 102660, 102670, 102720, 
    102760, 102780, 102790, 102810, 102820, 102810, 102820, 102840, 102780, 
    102750, 102750, 102730, 102720, 102720, 102710, 102660, 102670, 102640, 
    102620, 102600, 102550, 102490, 102430, 102400, 102400, 102350, 102300, 
    102260, 102230, 102180, 102110, 102060, 102020, 101950, 101900, 101840, 
    101790, 101750, 101670, 101590, 101520, 101450, 101380, 101270, 101180, 
    101140, 101090, 101050, 100990, 100960, 100890, 100840, 100770, 100700, 
    100650, 100620, 100540, 100460, 100390, 100370, 100370, 100350, 100320, 
    100300, 100320, 100320, 100320, 100360, 100380, 100400, 100370, 100420, 
    100400, 100410, 100410, 100450, 100470, 100490, 100480, 100500, 100510, 
    100550, 100560, 100570, 100570, 100610, 100610, 100600, 100620, 100620, 
    100640, 100640, 100620, 100600, 100600, 100610, 100590, 100570, 100560, 
    100580, 100560, 100580, 100570, 100620, 100640, 100650, 100680, 100720, 
    100750, 100770, 100850, 100870, 100890, 100900, 100920, 100940, 100960, 
    100990, 101000, 101030, 101060, 101090, 101120, 101130, 101130, 101170, 
    101180, 101210, 101220, 101230, 101240, 101240, 101250, 101270, 101280, 
    101280, 101290, 101300, 101300, 101280, 101270, 101240, 101200, 101180, 
    101170, 101150, 101090, 101040, 101010, 100960, 100920, 100880, 100830, 
    100800, 100730, 100700, 100660, 100610, 100560, 100490, 100430, 100390, 
    100330, 100290, 100280, 100270, 100260, 100290, 100290, 100340, 100370, 
    100400, 100430, 100490, 100520, 100560, 100590, 100620, 100670, 100730, 
    100780, 100850, 100890, 100990, 101070, 101100, 101150, 101200, 101250, 
    101300, 101360, 101380, 101390, 101430, 101420, 101420, 101420, 101430, 
    101430, 101420, 101410, 101440, 101470, 101520, 101580, 101640, 101730, 
    101810, 101920, 102040, 102130, 102210, 102320, 102350, 102410, 102470, 
    102580, 102680, 102770, 102800, 102880, 103020, 103000, 103030, 102990, 
    102950, 102860, 102770, 102670, 102480, 102340, 102210, 102070, 101950, 
    101840, 101680, 101520, 101360, 101180, 101080, 101040, 101020, 101040, 
    101020, 100970, 100970, 100930, 100850, 100770, 100710, 100590, 100490, 
    100320, 100170, 99990, 99820, 99770, 99660, 99570, 99450, 99370, 99380, 
    99360, 99500, 99570, 99650, 99660, 99680, 99700, 99740, 99760, 99910, 
    100070, 100250, 100430, 100670, 100980, 101250, 101550, 101650, 101940, 
    102070, 102200, 102280, 102390, 102440, 102550, 102600, 102660, 102740, 
    102810, 102830, 102850, 102830, 102780, 102710, 102600, 102570, 102470, 
    102360, 102250, 102110, 101980, 101850, 101690, 101670, 101640, 101620, 
    101620, 101600, 101600, 101690, 101720, 101780, 101850, 101880, 101910, 
    101950, 101970, 101980, 102030, 102050, 102050, 102040, 102070, 102060, 
    102020, 101990, 101950, 101890, 101840, 101800, 101740, 101630, 101520, 
    101440, 101320, 101200, 101130, 101000, 100870, 100750, 100640, 100480, 
    100330, 100200, 100060, 99950, 99850, 99720, 99600, 99500, 99400, 99330, 
    99290, 99260, 99290, 99330, 99420, 99530, 99640, 99730, 99860, 99940, 
    100030, 100100, 100200, 100320, 100390, 100470, 100500, 100570, 100640, 
    100710, 100780, 100800, 100850, 100900, 100920, 100930, 100970, 100950, 
    100970, 100980, 100990, 101020, 101050, 101100, 101120, 101160, 101180, 
    101170, 101170, 101190, 101220, 101270, 101280, 101320, 101330, 101330, 
    101340, 101350, 101370, 101380, 101390, 101400, 101420, 101450, 101490, 
    101500, 101530, 101540, 101540, 101550, 101560, 101560, 101570, 101550, 
    101570, 101580, 101600, 101610, 101630, 101610, 101620, 101630, 101650, 
    101660, 101630, 101630, 101640, 101630, 101660, 101670, 101670, 101670, 
    101660, 101640, 101610, 101570, 101520, 101480, 101430, 101390, 101330, 
    101280, 101200, 101120, 101000, 100910, 100840, 100740, 100610, 100480, 
    100350, 100260, 100130, 100050, 99930, 99870, 99890, 99860, 99830, 99840, 
    99800, 99710, 99690, 99670, 99650, 99620, 99580, 99550, 99520, 99480, 
    99450, 99440, 99450, 99480, 99520, 99520, 99560, 99580, 99600, 99610, 
    99560, 99520, 99480, 99320, 99130, 99270, 99510, 99610, 99610, 99680, 
    99810, 99860, 99850, 99800, 99770, 99760, 99830, 99850, 99890, 99960, 
    100060, 100110, 100130, 100110, 100070, 100140, 100080, 100090, 100130, 
    100120, 100160, 100080, 100110, 100110, 100120, 100110, 100110, 100120, 
    100110, 100120, 100160, 100170, 100210, 100210, 100220, 100260, 100230, 
    100260, 100260, 100240, 100200, 100200, 100230, 100280, 100280, 100280, 
    100310, 100300, 100300, 100310, 100320, 100320, 100350, 100340, 100330, 
    100260, 100280, 100270, 100270, 100260, 100260, 100250, 100220, 100180, 
    100180, 100140, 100160, 100120, 100090, 100060, 100060, 100010, 99990, 
    99950, 99880, 99830, 99770, 99730, 99660, 99620, 99560, 99540, 99530, 
    99560, 99560, 99570, 99560, 99540, 99540, 99530, 99530, 99490, 99480, 
    99490, 99510, 99500, 99490, 99520, 99500, 99470, 99420, 99420, 99420, 
    99380, 99350, 99330, 99340, 99340, 99350, 99310, 99280, 99260, 99220, 
    99200, 99160, 99150, 99150, 99160, 99120, 99100, 99110, 99090, 99090, 
    99070, 99060, 99050, 99020, 99040, 99040, 99050, 99060, 99070, 99080, 
    99090, 99080, 99120, 99140, 99160, 99160, 99160, 99130, 99180, 99180, 
    99170, 99150, 99130, 99100, 99080, 99090, 99070, 99040, 99010, 99000, 
    98980, 98980, 98990, 98990, 98980, 98940, 98930, 98940, 98930, 98960, 
    98970, 98970, 98970, 99000, 99040, 99080, 99100, 99120, 99140, 99170, 
    99200, 99210, 99230, 99250, 99280, 99290, 99340, 99360, 99380, 99380, 
    99390, 99400, 99400, 99400, 99390, 99360, 99340, 99360, 99360, 99310, 
    99240, 99210, 99170, 99150, 99160, 99100, 99080, 99050, 99040, 99020, 
    99010, 98990, 98950, 98960, 98970, 98970, 98970, 98950, 98970, 98970, 
    98980, 98980, 99010, 99030, 99020, 99030, 99060, 99060, 99090, 99100, 
    99120, 99140, 99170, 99210, 99220, 99250, 99270, 99280, 99270, 99280, 
    99290, 99310, 99330, 99320, 99320, 99370, 99440, 99430, 99480, 99510, 
    99530, 99580, 99590, 99650, 99690, 99740, 99790, 99860, 99930, 100000, 
    100040, 100050, 100080, 100150, 100200, 100240, 100260, 100290, 100290, 
    100350, 100380, 100430, 100460, 100490, 100550, 100580, 100620, 100670, 
    100690, 100730, 100770, 100830, 100870, 100850, 100810, 100770, 100710, 
    100690, 100670, 100700, 100750, 100750, 100750, 100780, 100780, 100790, 
    100790, 100740, 100660, 100590, 100500, 100430, 100340, 100280, 100170, 
    100090, 99990, 99880, 99780, 99760, 99770, 99800, 99910, 100030, 100120, 
    100170, 100230, 100320, 100410, 100470, 100480, 100540, 100580, 100560, 
    100600, 100570, 100550, 100540, 100540, 100540, 100500, 100470, 100420, 
    100380, 100330, 100250, 100190, 100090, 100040, 99910, 99820, 99680, 
    99520, 99310, 99030, 98790, 98620, 98550, 98550, 98530, 98520, 98560, 
    98650, 98760, 98830, 98910, 98950, 98950, 98970, 98960, 98930, 98880, 
    98820, 98870, 98940, 99010, 99120, 99180, 99250, 99350, 99470, 99610, 
    99780, 99880, 99940, 100030, 100130, 100170, 100250, 100270, 100300, 
    100290, 100280, 100260, 100220, 100170, 100090, 100010, 99940, 99820, 
    99710, 99610, 99510, 99450, 99360, 99310, 99270, 99250, 99240, 99250, 
    99280, 99270, 99290, 99310, 99300, 99320, 99310, 99310, 99310, 99300, 
    99290, 99250, 99210, 99230, 99310, 99420, 99580, 99760, 99810, 99890, 
    100010, 100100, 100210, 100280, 100400, 100490, 100550, 100630, 100660, 
    100710, 100720, 100730, 100740, 100740, 100730, 100740, 100780, 100860, 
    100890, 100900, 100950, 101010, 101050, 101070, 101130, 101200, 101290, 
    101340, 101430, 101490, 101590, 101670, 101760, 101820, 101900, 101950, 
    101970, 102020, 102140, 102200, 102240, 102300, 102330, 102370, 102400, 
    102410, 102440, 102440, 102440, 102420, 102400, 102390, 102360, 102320, 
    102310, 102270, 102190, 102080, 101950, 101880, 101860, 101800, 101740, 
    101700, 101690, 101690, 101640, 101570, 101530, 101480, 101380, 101330, 
    101300, 101290, 101260, 101280, 101270, 101250, 101240, 101230, 101200, 
    101200, 101180, 101210, 101260, 101290, 101320, 101330, 101320, 101360, 
    101390, 101420, 101430, 101450, 101450, 101420, 101400, 101380, 101360, 
    101360, 101370, 101340, 101310, 101280, 101240, 101220, 101180, 101160, 
    101120, 101120, 101110, 101070, 101070, 101060, 101030, 101020, 100980, 
    100920, 100890, 100870, 100850, 100820, 100760, 100730, 100710, 100690, 
    100660, 100650, 100600, 100570, 100540, 100490, 100440, 100380, 100320, 
    100240, 100180, 100120, 100050, 99970, 99890, 99800, 99720, 99620, 99490, 
    99300, 99150, 99020, 98880, 98770, 98700, 98580, 98470, 98390, 98340, 
    98260, 98210, 98220, 98180, 98230, 98320, 98420, 98570, 98680, 98790, 
    98890, 99010, 99120, 99200, 99280, 99370, 99470, 99530, 99610, 99740, 
    99800, 99860, 99880, 99900, 99940, 100010, 100060, 100130, 100200, 
    100220, 100280, 100300, 100360, 100380, 100410, 100400, 100380, 100380, 
    100340, 100270, 100190, 100150, 100120, 100070, 99990, 99900, 99860, 
    99800, 99740, 99710, 99680, 99660, 99630, 99630, 99610, 99620, 99610, 
    99610, 99630, 99650, 99670, 99700, 99730, 99750, 99750, 99800, 99840, 
    99870, 99900, 99910, 99930, 99960, 99930, 99920, 99910, 99930, 99920, 
    99900, 99880, 99880, 99880, 99880, 99860, 99860, 99880, 99890, 99880, 
    99890, 99910, 99960, 99990, 100000, 100010, 100000, 100060, 100080, 
    100100, 100100, 100110, 100120, 100120, 100130, 100170, 100220, 100240, 
    100240, 100270, 100270, 100320, 100320, 100340, 100350, 100360, 100390, 
    100400, 100440, 100440, 100470, 100470, 100500, 100490, 100510, 100520, 
    100530, 100520, 100520, 100490, 100450, 100400, 100390, 100290, 100260, 
    100220, 100190, 100180, 100170, 100170, 100190, 100200, 100270, 100290, 
    100290, 100260, 100190, 100120, 100030, 99960, 99860, 99760, 99680, 
    99640, 99550, 99450, 99360, 99280, 99210, 99200, 99210, 99210, 99250, 
    99300, 99380, 99460, 99520, 99600, 99660, 99700, 99730, 99780, 99820, 
    99840, 99850, 99850, 99900, 99980, 100050, 100120, 100190, 100260, 
    100340, 100410, 100460, 100520, 100520, 100540, 100550, 100570, 100590, 
    100600, 100610, 100600, 100590, 100580, 100570, 100570, 100560, 100550, 
    100550, 100580, 100620, 100650, 100660, 100700, 100720, 100730, 100730, 
    100700, 100680, 100670, 100690, 100700, 100670, 100670, 100630, 100620, 
    100590, 100550, 100510, 100420, 100360, 100310, 100270, 100230, 100220, 
    100240, 100260, 100300, 100330, 100380, 100410, 100450, 100490, 100550, 
    100590, 100670, 100740, 100800, 100850, 100890, 100940, 100970, 101030, 
    101070, 101130, 101170, 101210, 101250, 101310, 101370, 101420, 101460, 
    101520, 101560, 101580, 101580, 101640, 101630, 101650, 101690, 101680, 
    101680, 101680, 101650, 101630, 101620, 101560, 101490, 101440, 101370, 
    101260, 101140, 101020, 100890, 100780, 100690, 100600, 100530, 100450, 
    100390, 100330, 100280, 100230, 100230, 100210, 100230, 100250, 100270, 
    100290, 100350, 100390, 100430, 100500, 100530, 100560, 100600, 100610, 
    100620, 100660, 100720, 100730, 100740, 100760, 100740, 100750, 100770, 
    100790, 100830, 100860, 100840, 100850, 100830, 100840, 100820, 100790, 
    100740, 100690, 100660, 100640, 100620, 100590, 100560, 100550, 100570, 
    100570, 100550, 100540, 100550, 100560, 100520, 100480, 100460, 100400, 
    100390, 100390, 100350, 100250, 100150, 100160, 100130, 100050, 99970, 
    99900, 99870, 99850, 99870, 99800, 99790, 99720, 99720, 99700, 99720, 
    99680, 99660, 99660, 99630, 99630, 99630, 99580, 99550, 99560, 99620, 
    99570, 99580, 99590, 99610, 99610, 99600, 99600, 99620, 99670, 99700, 
    99710, 99700, 99690, 99750, 99760, 99830, 99910, 99940, 99960, 99960, 
    99950, 99950, 99970, 100040, 100010, 100020, 100110, 100190, 100270, 
    100370, 100460, 100530, 100620, 100710, 100780, 100830, 100900, 100920, 
    100940, 100980, 101040, 101100, 101140, 101160, 101170, 101180, 101180, 
    101190, 101170, 101130, 101110, 101070, 100990, 100950, 100890, 100820, 
    100750, 100670, 100620, 100540, 100440, 100370, 100270, 100170, 100100, 
    100060, 100040, 100040, 100000, 99960, 99960, 99970, 99950, 99910, 99830, 
    99770, 99730, 99640, 99610, 99480, 99340, 99210, 99100, 98920, 98750, 
    98590, 98400, 98360, 98240, 98180, 98100, 98080, 98030, 97940, 97940, 
    98010, 98150, 98250, 98370, 98510, 98620, 98770, 98890, 98930, 99140, 
    99210, 99400, 99540, 99680, 99640, 99750, 99840, 99900, 99920, 99910, 
    99980, 99990, 100000, 100000, 100020, 100070, 100080, 100060, 100090, 
    100110, 100120, 100160, 100160, 100150, 100140, 100140, 100130, 100070, 
    100040, 100040, 100040, 100040, 100010, 99980, 99960, 99930, 99910, 
    99880, 99860, 99820, 99790, 99740, 99710, 99660, 99630, 99580, 99560, 
    99510, 99460, 99430, 99410, 99360, 99350, 99320, 99280, 99240, 99190, 
    99160, 99160, 99140, 99130, 99160, 99190, 99230, 99260, 99290, 99280, 
    99290, 99340, 99380, 99430, 99470, 99470, 99510, 99550, 99590, 99610, 
    99640, 99650, 99690, 99750, 99780, 99820, 99850, 99870, 99910, 99950, 
    99970, 100000, 100020, 100030, 100050, 100080, 100110, 100160, 100150, 
    100140, 100120, 100110, 100110, 100140, 100130, 100120, 100130, 100140, 
    100140, 100150, 100160, 100160, 100160, 100160, 100180, 100180, 100170, 
    100170, 100150, 100150, 100150, 100160, 100160, 100160, 100150, 100130, 
    100140, 100150, 100120, 100120, 100130, 100120, 100120, 100140, 100130, 
    100100, 100100, 100080, 100060, 100050, 100050, 100040, 100050, 100050, 
    100050, 100060, 100060, 100040, 100030, 100040, 100040, 100040, 100060, 
    100060, 100050, 100070, 100090, 100110, 100090, 100060, 100050, 100040, 
    100040, 100050, 100070, 100060, 100040, 100030, 100030, 100030, 100010, 
    99990, 99950, 99930, 99920, 99900, 99880, 99860, 99840, 99840, 99850, 
    99860, 99860, 99860, 99850, 99850, 99830, 99830, 99820, 99830, 99820, 
    99820, 99820, 99860, 99890, 99900, 99920, 99900, 99910, 99910, 99940, 
    99980, 100020, 100050, 100090, 100100, 100130, 100190, 100220, 100260, 
    100300, 100330, 100380, 100410, 100450, 100490, 100550, 100590, 100650, 
    100690, 100730, 100750, 100810, 100840, 100880, 100910, 100950, 101010, 
    101050, 101120, 101150, 101170, 101180, 101220, 101250, 101280, 101300, 
    101320, 101340, 101360, 101400, 101430, 101450, 101480, 101510, 101510, 
    101540, 101550, 101550, 101570, 101610, 101640, 101680, 101710, 101730, 
    101770, 101760, 101770, 101790, 101810, 101830, 101850, 101870, 101860, 
    101860, 101910, 101920, 101920, 101930, 101950, 101970, 101990, 102000, 
    102020, 102060, 102100, 102120, 102170, 102180, 102210, 102220, 102250, 
    102270, 102290, 102310, 102340, 102370, 102400, 102430, 102480, 102500, 
    102510, 102510, 102540, 102560, 102570, 102580, 102600, 102630, 102650, 
    102670, 102680, 102700, 102710, 102710, 102710, 102750, 102750, 102740, 
    102760, 102760, 102780, 102790, 102800, 102800, 102800, 102800, 102780, 
    102770, 102770, 102750, 102720, 102740, 102740, 102720, 102680, 102670, 
    102630, 102620, 102620, 102580, 102600, 102570, 102570, 102530, 102510, 
    102490, 102480, 102450, 102410, 102400, 102390, 102380, 102350, 102320, 
    102300, 102320, 102320, 102320, 102320, 102310, 102300, 102280, 102290, 
    102290, 102280, 102270, 102270, 102260, 102260, 102250, 102240, 102230, 
    102190, 102160, 102150, 102110, 102060, 102040, 102010, 101990, 101950, 
    101910, 101850, 101820, 101760, 101710, 101680, 101630, 101610, 101540, 
    101510, 101460, 101420, 101390, 101360, 101320, 101290, 101230, 101190, 
    101150, 101110, 101060, 101030, 101000, 101000, 101000, 101030, 101020, 
    101020, 101050, 101050, 101070, 101070, 101060, 101050, 101060, 101070, 
    101100, 101110, 101130, 101150, 101170, 101220, 101220, 101240, 101280, 
    101290, 101300, 101320, 101340, 101370, 101370, 101330, 101360, 101370, 
    101370, 101360, 101360, 101380, 101390, 101400, 101400, 101400, 101390, 
    101390, 101370, 101370, 101370, 101350, 101370, 101310, 101310, 101290, 
    101300, 101290, 101270, 101270, 101230, 101180, 101200, 101170, 101160, 
    101140, 101120, 101100, 101110, 101100, 101110, 101100, 101070, 101050, 
    101020, 100990, 100960, 100940, 100920, 100890, 100870, 100860, 100820, 
    100780, 100740, 100690, 100660, 100640, 100560, 100530, 100520, 100540, 
    100590, 100660, 100720, 100770, 100810, 100860, 100920, 100960, 101030, 
    101070, 101130, 101180, 101250, 101320, 101410, 101460, 101520, 101590, 
    101640, 101690, 101760, 101820, 101890, 101970, 102050, 102110, 102180, 
    102210, 102240, 102270, 102290, 102330, 102370, 102420, 102460, 102500, 
    102550, 102580, 102620, 102650, 102650, 102660, 102670, 102700, 102710, 
    102730, 102760, 102770, 102800, 102830, 102830, 102830, 102820, 102800, 
    102790, 102790, 102770, 102760, 102760, 102750, 102740, 102730, 102720, 
    102700, 102640, 102590, 102540, 102520, 102490, 102450, 102400, 102370, 
    102320, 102300, 102280, 102260, 102260, 102250, 102230, 102200, 102190, 
    102180, 102190, 102220, 102230, 102250, 102270, 102270, 102250, 102230, 
    102200, 102190, 102200, 102200, 102200, 102190, 102200, 102190, 102180, 
    102170, 102150, 102130, 102100, 102080, 102080, 102070, 102070, 102080, 
    102070, 102070, 102080, 102060, 102030, 102020, 101990, 101980, 101960, 
    101960, 101970, 101980, 102000, 101990, 101990, 102000, 101990, 102010, 
    102000, 101990, 102000, 101990, 102010, 102010, 102030, 102040, 102050, 
    102070, 102070, 102050, 102050, 102050, 102050, 102050, 102060, 102080, 
    102080, 102080, 102090, 102080, 102050, 102020, 102000, 101950, 101910, 
    101880, 101860, 101880, 101850, 101830, 101780, 101760, 101700, 101650, 
    101590, 101530, 101480, 101420, 101360, 101330, 101280, 101230, 101180, 
    101120, 101050, 101030, 101000, 100970, 100920, 100890, 100880, 100870, 
    100850, 100830, 100820, 100820, 100820, 100790, 100740, 100730, 100710, 
    100680, 100670, 100670, 100680, 100680, 100680, 100700, 100700, 100710, 
    100680, 100670, 100700, 100700, 100730, 100740, 100730, 100740, 100730, 
    100710, 100700, 100710, 100710, 100700, 100670, 100650, 100660, 100650, 
    100630, 100610, 100580, 100560, 100510, 100480, 100480, 100430, 100430, 
    100430, 100410, 100410, 100420, 100410, 100390, 100370, 100360, 100340, 
    100310, 100300, 100280, 100280, 100260, 100240, 100220, 100200, 100180, 
    100160, 100140, 100110, 100080, 100050, 100050, 100060, 100060, 100070, 
    100080, 100060, 100070, 100080, 100060, 100050, 100030, 100020, 100020, 
    100010, 100010, 100000, 100000, 100020, 100010, 100000, 100030, 100040, 
    100040, 100050, 100080, 100090, 100110, 100150, 100180, 100190, 100200, 
    100240, 100280, 100310, 100320, 100330, 100360, 100370, 100370, 100420, 
    100420, 100460, 100480, 100460, 100480, 100500, 100510, 100530, 100550, 
    100560, 100560, 100600, 100600, 100630, 100640, 100650, 100660, 100640, 
    100630, 100600, 100570, 100560, 100550, 100520, 100490, 100470, 100440, 
    100420, 100390, 100370, 100350, 100320, 100310, 100310, 100300, 100330, 
    100340, 100340, 100360, 100360, 100360, 100330, 100350, 100350, 100320, 
    100290, 100280, 100250, 100240, 100220, 100180, 100140, 100100, 100070, 
    100020, 99950, 99860, 99780, 99710, 99670, 99610, 99570, 99500, 99440, 
    99390, 99350, 99320, 99300, 99300, 99280, 99290, 99300, 99330, 99380, 
    99420, 99470, 99510, 99540, 99630, 99680, 99740, 99780, 99830, 99910, 
    99960, 100000, 100060, 100100, 100130, 100170, 100210, 100210, 100240, 
    100270, 100280, 100300, 100320, 100360, 100360, 100350, 100310, 100300, 
    100280, 100260, 100260, 100250, 100260, 100270, 100300, 100330, 100350, 
    100380, 100400, 100440, 100490, 100560, 100630, 100690, 100770, 100840, 
    100900, 100950, 101000, 101030, 101080, 101130, 101190, 101250, 101270, 
    101320, 101350, 101440, 101480, 101540, 101580, 101630, 101660, 101680, 
    101690, 101710, 101710, 101690, 101680, 101680, 101670, 101690, 101690, 
    101650, 101630, 101600, 101550, 101530, 101500, 101510, 101480, 101440, 
    101430, 101400, 101370, 101340, 101290, 101250, 101210, 101150, 101130, 
    101110, 101080, 101080, 101030, 101000, 100970, 100930, 100910, 100850, 
    100810, 100750, 100700, 100660, 100620, 100600, 100590, 100580, 100540, 
    100530, 100500, 100490, 100480, 100460, 100450, 100480, 100490, 100490, 
    100510, 100540, 100540, 100520, 100520, 100530, 100540, 100550, 100560, 
    100570, 100590, 100600, 100620, 100650, 100620, 100600, 100590, 100510, 
    100470, 100400, 100340, 100290, 100250, 100200, 100200, 100210, 100230, 
    100240, 100260, 100300, 100350, 100380, 100430, 100490, 100510, 100540, 
    100570, 100560, 100550, 100590, 100570, 100510, 100430, 100330, 100220, 
    100040, 99890, 99790, 99710, 99640, 99610, 99520, 99470, 99440, 99370, 
    99330, 99210, 99080, 98960, 98810, 98640, 98480, 98330, 98180, 98090, 
    98010, 97980, 97970, 97950, 97950, 97950, 97980, 98000, 98040, 98100, 
    98150, 98210, 98280, 98380, 98470, 98540, 98660, 98790, 98880, 98990, 
    99100, 99180, 99270, 99340, 99390, 99450, 99520, 99520, 99550, 99590, 
    99580, 99610, 99590, 99580, 99500, 99430, 99390, 99340, 99260, 99170, 
    99170, 99130, 99130, 99140, 99180, 99250, 99320, 99420, 99510, 99610, 
    99790, 99910, 100030, 100190, 100390, 100570, 100680, 100790, 100910, 
    101010, 101110, 101180, 101260, 101280, 101310, 101370, 101410, 101440, 
    101490, 101480, 101490, 101490, 101490, 101430, 101410, 101390, 101370, 
    101390, 101390, 101430, 101420, 101410, 101420, 101420, 101380, 101350, 
    101280, 101230, 101230, 101210, 101220, 101240, 101220, 101180, 101040, 
    100970, 100920, 100850, 100770, 100640, 100540, 100490, 100490, 100480, 
    100470, 100440, 100430, 100450, 100450, 100450, 100480, 100510, 100520, 
    100610, 100660, 100690, 100750, 100800, 100830, 100860, 100900, 100920, 
    100920, 100880, 100860, 100860, 100850, 100820, 100830, 100800, 100800, 
    100780, 100770, 100770, 100710, 100690, 100730, 100720, 100740, 100760, 
    100810, 100810, 100880, 100930, 100930, 100980, 100960, 100960, 101000, 
    101030, 101010, 101050, 101010, 101060, 101100, 101090, 101110, 101120, 
    101120, 101090, 101130, 101130, 101100, 101080, 101120, 101100, 101060, 
    101030, 100980, 100930, 100870, 100850, 100780, 100730, 100640, 100580, 
    100520, 100440, 100330, 100210, 100110, 100060, 100050, 100030, 99980, 
    99960, 99960, 99940, 99970, 99950, 99970, 99980, 99910, 99900, 99890, 
    99890, 99850, 99820, 99800, 99780, 99760, 99760, 99740, 99740, 99740, 
    99730, 99730, 99720, 99800, 99820, 99850, 99920, 99900, 99960, 99950, 
    99960, 99900, 99980, 99980, 99990, 100030, 100040, 100040, 100060, 
    100100, 100110, 100100, 100020, 100030, 99970, 99950, 99890, 99790, 
    99760, 99710, 99640, 99630, 99560, 99560, 99520, 99490, 99480, 99450, 
    99420, 99400, 99360, 99340, 99290, 99250, 99210, 99180, 99150, 99100, 
    99060, 99070, 99060, 99080, 99100, 99120, 99120, 99160, 99210, 99230, 
    99220, 99180, 99230, 99200, 99210, 99200, 99170, 99210, 99250, 99320, 
    99370, 99380, 99390, 99420, 99420, 99430, 99430, 99480, 99490, 99560, 
    99680, 99740, 99870, 99990, 100050, 100100, 100180, 100290, 100330, 
    100330, 100380, 100420, 100440, 100430, 100440, 100490, 100530, 100500, 
    100570, 100600, 100600, 100560, 100610, 100620, 100640, 100650, 100650, 
    100670, 100670, 100680, 100700, 100720, 100730, 100730, 100730, 100740, 
    100730, 100740, 100750, 100740, 100760, 100750, 100740, 100720, 100720, 
    100720, 100740, 100740, 100780, 100790, 100800, 100800, 100800, 100800, 
    100750, 100740, 100720, 100710, 100670, 100660, 100630, 100590, 100570, 
    100550, 100510, 100490, 100460, 100390, 100350, 100330, 100310, 100270, 
    100270, 100210, 100210, 100160, 100130, 100070, 100010, 99980, 99930, 
    99890, 99890, 99890, 99860, 99840, 99850, 99830, 99820, 99830, 99810, 
    99800, 99810, 99830, 99830, 99850, 99860, 99880, 99890, 99900, 99920, 
    99930, 99940, 99960, 99980, 99980, 100010, 100050, 100080, 100120, 
    100140, 100160, 100190, 100220, 100260, 100280, 100310, 100310, 100350, 
    100380, 100410, 100430, 100460, 100460, 100450, 100450, 100450, 100460, 
    100470, 100450, 100450, 100450, 100440, 100430, 100440, 100430, 100420, 
    100380, 100370, 100340, 100330, 100320, 100300, 100290, 100270, 100290, 
    100260, 100220, 100230, 100220, 100190, 100180, 100190, 100190, 100190, 
    100230, 100220, 100220, 100200, 100210, 100190, 100180, 100190, 100180, 
    100170, 100160, 100170, 100190, 100210, 100210, 100210, 100180, 100170, 
    100150, 100140, 100100, 100080, 100050, 100050, 100010, 100000, 99990, 
    99980, 99950, 99920, 99920, 99890, 99870, 99870, 99850, 99850, 99850, 
    99870, 99870, 99850, 99840, 99810, 99800, 99780, 99780, 99770, 99740, 
    99750, 99730, 99750, 99770, 99760, 99760, 99770, 99790, 99780, 99740, 
    99760, 99800, 99820, 99850, 99860, 99890, 99910, 99910, 99940, 99950, 
    99980, 100000, 100030, 100060, 100090, 100140, 100160, 100190, 100210, 
    100230, 100250, 100300, 100300, 100300, 100300, 100320, 100340, 100350, 
    100360, 100370, 100390, 100400, 100400, 100410, 100410, 100430, 100440, 
    100450, 100470, 100490, 100450, 100440, 100440, 100440, 100450, 100420, 
    100420, 100390, 100380, 100350, 100360, 100360, 100330, 100360, 100360, 
    100290, 100320, 100330, 100350, 100330, 100330, 100300, 100290, 100300, 
    100320, 100310, 100310, 100320, 100290, 100230, 100190, 100130, 100060, 
    99890, 99770, 99660, 99540, 99450, 99280, 99100, 99020, 98850, 98900, 
    98990, 99080, 99140, 99330, 99540, 99730, 99870, 99930, 99980, 100120, 
    100170, 100230, 100260, 100290, 100360, 100440, 100490, 100520, 100590, 
    100590, 100570, 100510, 100470, 100410, 100310, 100240, 100170, 100140, 
    100010, 99920, 99750, 99560, 99430, 99300, 99170, 99040, 98890, 98770, 
    98630, 98550, 98460, 98450, 98420, 98440, 98460, 98510, 98580, 98660, 
    98740, 98820, 98870, 98920, 98960, 99030, 99080, 99100, 99080, 99090, 
    99060, 99040, 99030, 98970, 98940, 98900, 98900, 98880, 98830, 98790, 
    98740, 98720, 98710, 98680, 98630, 98580, 98530, 98510, 98460, 98410, 
    98330, 98270, 98240, 98150, 98080, 97970, 97860, 97840, 97790, 97770, 
    97750, 97740, 97750, 97770, 97770, 97800, 97850, 97900, 97970, 98030, 
    98030, 98080, 98100, 98140, 98130, 98110, 98080, 98040, 97970, 97960, 
    97920, 97880, 97860, 97800, 97790, 97800, 97800, 97770, 97770, 97780, 
    97800, 97850, 97880, 97950, 97970, 98000, 98040, 98110, 98170, 98230, 
    98300, 98360, 98430, 98510, 98570, 98630, 98700, 98770, 98860, 98900, 
    98990, 99040, 99060, 99110, 99120, 99140, 99200, 99220, 99250, 99220, 
    99200, 99240, 99260, 99250, 99210, 99170, 99160, 99140, 99190, 99320, 
    99390, 99460, 99500, 99650, 99730, 99780, 99890, 99980, 100010, 100070, 
    100140, 100210, 100270, 100340, 100460, 100490, 100560, 100590, 100630, 
    100620, 100670, 100700, 100670, 100660, 100640, 100650, 100650, 100650, 
    100650, 100620, 100590, 100510, 100440, 100390, 100330, 100260, 100200, 
    100140, 100070, 100040, 99990, 99950, 99890, 99820, 99780, 99720, 99680, 
    99630, 99580, 99540, 99520, 99490, 99450, 99410, 99350, 99300, 99310, 
    99290, 99260, 99180, 99140, 99080, 99060, 99030, 98950, 98890, 98850, 
    98760, 98690, 98620, 98540, 98510, 98460, 98390, 98340, 98340, 98320, 
    98260, 98210, 98150, 98090, 98040, 97980, 97920, 97830, 97760, 97680, 
    97600, 97550, 97460, 97430, 97510, 97520, 97510, 97480, 97500, 97510, 
    97570, 97650, 97730, 97750, 97740, 97800, 97820, 97770, 97910, 97960, 
    98030, 98100, 98200, 98280, 98330, 98430, 98530, 98610, 98650, 98740, 
    98780, 98870, 98940, 98980, 99000, 99050, 99080, 99110, 99110, 99120, 
    99110, 99140, 99140, 99200, 99240, 99280, 99300, 99330, 99320, 99320, 
    99330, 99310, 99310, 99300, 99270, 99310, 99360, 99330, 99310, 99290, 
    99320, 99350, 99340, 99330, 99360, 99400, 99380, 99390, 99370, 99390, 
    99430, 99430, 99430, 99470, 99470, 99480, 99480, 99500, 99490, 99520, 
    99530, 99530, 99550, 99560, 99600, 99620, 99640, 99670, 99680, 99690, 
    99670, 99660, 99650, 99680, 99670, 99700, 99730, 99770, 99780, 99810, 
    99810, 99810, 99850, 99860, 99840, 99870, 99900, 99960, 100000, 100020, 
    100030, 100070, 100100, 100130, 100170, 100190, 100220, 100260, 100280, 
    100330, 100370, 100410, 100430, 100450, 100460, 100500, 100500, 100510, 
    100520, 100550, 100590, 100650, 100660, 100690, 100730, 100750, 100780, 
    100800, 100810, 100860, 100880, 100910, 100950, 100980, 101060, 101090, 
    101100, 101110, 101170, 101200, 101190, 101220, 101240, 101270, 101290, 
    101320, 101370, 101380, 101380, 101370, 101350, 101280, 101220, 101090, 
    100950, 100840, 100700, 100510, 100380, 100230, 100050, 99890, 99860, 
    99770, 99800, 99830, 99900, 99930, 99960, 100010, 100070, 100130, 100240, 
    100330, 100450, 100510, 100590, 100640, 100660, 100660, 100680, 100690, 
    100680, 100670, 100540, 100520, 100470, 100450, 100420, 100400, 100400, 
    100420, 100470, 100510, 100590, 100660, 100740, 100800, 100910, 101080, 
    101170, 101300, 101450, 101570, 101690, 101810, 101880, 101970, 102040, 
    102100, 102150, 102230, 102300, 102390, 102430, 102490, 102540, 102580, 
    102620, 102640, 102650, 102660, 102670, 102650, 102660, 102660, 102680, 
    102690, 102730, 102790, 102850, 102860, 102870, 102900, 102930, 102970, 
    103040, 103080, 103090, 103120, 103150, 103160, 103190, 103220, 103240, 
    103260, 103270, 103270, 103280, 103260, 103260, 103250, 103250, 103240, 
    103170, 103100, 103060, 103020, 102990, 102890, 102820, 102770, 102670, 
    102570, 102460, 102380, 102320, 102290, 102250, 102210, 102180, 102150, 
    102110, 102080, 102030, 102000, 101970, 101930, 101890, 101840, 101780, 
    101720, 101680, 101640, 101600, 101550, 101480, 101450, 101390, 101360, 
    101330, 101300, 101280, 101260, 101270, 101270, 101250, 101260, 101270, 
    101290, 101310, 101320, 101340, 101370, 101420, 101440, 101470, 101470, 
    101490, 101520, 101540, 101580, 101640, 101690, 101760, 101830, 101870, 
    101920, 101960, 101990, 102020, 102040, 102060, 102070, 102100, 102110, 
    102150, 102130, 102120, 102130, 102130, 102110, 102090, 102050, 102030, 
    102010, 101980, 101950, 101900, 101870, 101840, 101820, 101780, 101720, 
    101670, 101620, 101600, 101540, 101510, 101500, 101470, 101410, 101430, 
    101380, 101360, 101320, 101290, 101260, 101260, 101220, 101220, 101260, 
    101280, 101260, 101260, 101280, 101250, 101240, 101190, 101180, 101120, 
    101110, 101140, 101150, 101160, 101130, 101140, 101160, 101180, 101110, 
    101010, 100960, 100870, 100810, 100730, 100630, 100640, 100600, 100610, 
    100640, 100700, 100700, 100710, 100740, 100770, 100800, 100850, 100900, 
    100960, 101020, 101070, 101150, 101270, 101370, 101460, 101560, 101660, 
    101750, 101810, 101900, 101990, 102010, 102030, 102040, 102020, 101980, 
    101920, 101860, 101830, 101800, 101750, 101690, 101640, 101570, 101500, 
    101500, 101450, 101400, 101420, 101380, 101360, 101390, 101410, 101460, 
    101480, 101490, 101500, 101480, 101430, 101370, 101330, 101320, 101270, 
    101190, 101140, 101120, 101110, 101120, 101110, 101160, 101210, 101280, 
    101320, 101380, 101430, 101510, 101590, 101650, 101710, 101760, 101780, 
    101800, 101790, 101800, 101780, 101740, 101700, 101670, 101610, 101550, 
    101540, 101510, 101500, 101440, 101410, 101390, 101390, 101350, 101310, 
    101310, 101310, 101320, 101320, 101310, 101310, 101320, 101310, 101310, 
    101300, 101260, 101220, 101160, 101120, 101100, 101100, 101130, 101100, 
    101050, 101030, 101050, 101030, 101000, 100980, 100980, 100990, 100980, 
    100950, 100920, 100890, 100800, 100700, 100600, 100490, 100400, 100310, 
    100200, 100080, 100040, 100020, 100020, 100010, 100030, 100170, 100320, 
    100440, 100530, 100610, 100660, 100710, 100660, 100700, 100720, 100700, 
    100680, 100620, 100520, 100440, 100390, 100280, 100160, 100080, 100050, 
    100000, 99980, 99940, 99870, 99830, 99810, 99800, 99810, 99800, 99800, 
    99810, 99840, 99900, 99940, 99970, 100010, 100040, 100110, 100230, 
    100310, 100400, 100480, 100550, 100630, 100720, 100800, 100870, 100950, 
    101020, 101050, 101090, 101130, 101170, 101210, 101260, 101290, 101310, 
    101300, 101310, 101300, 101290, 101250, 101200, 101190, 101160, 101120, 
    101060, 101040, 101030, 101010, 100990, 100940, 100910, 100910, 100890, 
    100880, 100900, 100910, 100930, 100960, 100990, 101020, 101040, 101080, 
    101120, 101150, 101190, 101230, 101260, 101310, 101340, 101390, 101450, 
    101500, 101560, 101630, 101690, 101760, 101820, 101900, 101960, 102020, 
    102080, 102120, 102190, 102250, 102260, 102300, 102320, 102300, 102320, 
    102290, 102280, 102260, 102260, 102300, 102310, 102320, 102330, 102330, 
    102340, 102350, 102360, 102360, 102330, 102340, 102350, 102350, 102360, 
    102360, 102360, 102330, 102330, 102290, 102270, 102220, 102170, 102150, 
    102110, 102110, 102100, 102120, 102100, 102100, 102100, 102110, 102130, 
    102130, 102160, 102180, 102190, 102210, 102260, 102320, 102350, 102390, 
    102430, 102470, 102510, 102530, 102540, 102570, 102590, 102610, 102630, 
    102670, 102660, 102670, 102670, 102650, 102630, 102620, 102590, 102580, 
    102570, 102570, 102570, 102570, 102560, 102530, 102500, 102480, 102460, 
    102430, 102400, 102370, 102340, 102320, 102300, 102280, 102250, 102230, 
    102220, 102220, 102220, 102230, 102230, 102250, 102270, 102300, 102320, 
    102350, 102380, 102400, 102410, 102450, 102480, 102470, 102470, 102490, 
    102510, 102540, 102550, 102570, 102570, 102560, 102550, 102550, 102500, 
    102460, 102410, 102360, 102300, 102270, 102220, 102140, 102090, 101980, 
    101870, 101780, 101690, 101590, 101550, 101570, 101600, 101690, 101770, 
    101780, 101790, 101870, 101910, 101960, 101980, 101970, 101960, 101960, 
    101990, 101980, 102000, 101960, 101940, 101910, 101910, 101840, 101870, 
    101830, 101810, 101780, 101710, 101710, 101700, 101710, 101710, 101660, 
    101640, 101590, 101550, 101520, 101490, 101480, 101480, 101520, 101560, 
    101600, 101620, 101660, 101720, 101660, 101720, 101800, 101880, 101970, 
    101990, 102140, 102220, 102350, 102390, 102450, 102420, 102420, 102470, 
    102510, 102590, 102570, 102600, 102610, 102590, 102570, 102580, 102550, 
    102450, 102300, 102250, 102140, 101990, 101830, 101680, 101600, 101460, 
    101320, 101220, 101150, 101080, 101020, 100950, 100990, 100930, 100900, 
    100880, 100860, 100860, 100870, 100910, 100960, 101010, 100990, 101010, 
    101070, 101040, 101120, 101140, 101140, 101180, 101210, 101240, 101250, 
    101310, 101340, 101390, 101420, 101500, 101560, 101630, 101680, 101770, 
    101810, 101860, 101910, 101940, 101990, 102000, 102030, 102040, 102060, 
    102110, 102140, 102110, 102150, 102180, 102210, 102200, 102200, 102190, 
    102200, 102190, 102200, 102160, 102170, 102160, 102150, 102150, 102150, 
    102170, 102150, 102120, 102100, 102080, 102070, 102030, 102030, 101990, 
    101950, 101930, 101920, 101900, 101880, 101900, 101930, 101940, 101930, 
    101930, 101960, 101970, 101990, 102000, 102010, 102030, 102040, 102020, 
    102010, 102020, 102060, 102100, 102140, 102150, 102190, 102230, 102250, 
    102260, 102300, 102320, 102320, 102340, 102380, 102380, 102390, 102400, 
    102400, 102410, 102420, 102450, 102380, 102380, 102400, 102390, 102420, 
    102450, 102480, 102500, 102540, 102520, 102570, 102600, 102590, 102600, 
    102600, 102630, 102650, 102670, 102690, 102670, 102660, 102650, 102640, 
    102610, 102590, 102570, 102540, 102490, 102460, 102430, 102360, 102340, 
    102300, 102260, 102220, 102170, 102110, 102030, 101940, 101910, 101880, 
    101830, 101850, 101840, 101840, 101810, 101810, 101810, 101820, 101840, 
    101850, 101860, 101880, 101900, 101950, 101980, 102060, 102140, 102200, 
    102250, 102300, 102340, 102390, 102410, 102450, 102470, 102520, 102580, 
    102620, 102640, 102670, 102680, 102700, 102730, 102760, 102780, 102820, 
    102850, 102890, 102920, 102950, 102960, 102970, 102980, 102970, 102970, 
    102970, 102960, 102960, 102980, 102980, 102980, 102980, 102960, 102950, 
    102950, 102930, 102920, 102910, 102920, 102930, 102940, 102960, 102950, 
    102950, 102970, 103000, 102990, 102960, 102940, 102950, 102970, 102950, 
    102970, 103010, 103030, 103010, 103030, 103020, 102960, 102920, 102910, 
    102880, 102860, 102850, 102840, 102830, 102810, 102790, 102720, 102660, 
    102630, 102610, 102510, 102460, 102420, 102370, 102320, 102320, 102290, 
    102220, 102220, 102070, 101930, 101870, 101840, 101750, 101660, 101720, 
    101580, 101570, 101530, 101480, 101410, 101360, 101310, 101270, 101220, 
    101180, 101130, 101100, 101070, 101070, 101010, 100960, 100950, 100870, 
    100830, 100800, 100760, 100700, 100650, 100620, 100610, 100600, 100600, 
    100570, 100570, 100580, 100580, 100600, 100610, 100610, 100620, 100640, 
    100670, 100690, 100720, 100740, 100760, 100790, 100830, 100890, 100920, 
    100940, 100960, 100980, 101000, 101040, 101060, 101100, 101120, 101140, 
    101200, 101210, 101240, 101270, 101260, 101280, 101350, 101410, 101470, 
    101510, 101560, 101630, 101700, 101750, 101800, 101830, 101860, 101900, 
    101940, 102000, 102040, 102070, 102090, 102100, 102130, 102150, 102170, 
    102180, 102210, 102220, 102250, 102260, 102270, 102290, 102300, 102330, 
    102340, 102360, 102390, 102380, 102380, 102430, 102420, 102440, 102450, 
    102470, 102490, 102500, 102540, 102550, 102590, 102580, 102600, 102610, 
    102630, 102650, 102680, 102730, 102740, 102750, 102770, 102770, 102790, 
    102760, 102790, 102780, 102780, 102800, 102820, 102830, 102840, 102820, 
    102810, 102810, 102800, 102810, 102820, 102820, 102820, 102840, 102850, 
    102880, 102900, 102910, 102910, 102930, 102940, 102930, 102910, 102900, 
    102890, 102890, 102910, 102890, 102900, 102880, 102880, 102850, 102840, 
    102830, 102830, 102830, 102840, 102850, 102860, 102870, 102900, 102890, 
    102890, 102900, 102900, 102900, 102900, 102890, 102880, 102890, 102890, 
    102880, 102870, 102880, 102880, 102870, 102860, 102840, 102830, 102820, 
    102820, 102820, 102830, 102830, 102830, 102830, 102810, 102810, 102810, 
    102800, 102820, 102840, 102860, 102880, 102920, 102960, 102970, 103010, 
    103020, 103020, 103010, 103010, 103010, 103000, 103000, 102980, 102950, 
    102930, 102910, 102890, 102860, 102840, 102790, 102750, 102730, 102680, 
    102650, 102630, 102580, 102610, 102580, 102550, 102550, 102490, 102450, 
    102410, 102390, 102350, 102310, 102300, 102240, 102230, 102200, 102150, 
    102090, 102040, 101980, 101930, 101880, 101830, 101820, 101770, 101730, 
    101690, 101660, 101580, 101600, 101590, 101570, 101560, 101540, 101530, 
    101510, 101490, 101500, 101520, 101510, 101510, 101500, 101510, 101510, 
    101480, 101490, 101490, 101500, 101530, 101560, 101570, 101600, 101620, 
    101650, 101630, 101620, 101620, 101590, 101560, 101540, 101530, 101480, 
    101460, 101420, 101400, 101370, 101340, 101330, 101310, 101270, 101240, 
    101210, 101200, 101170, 101170, 101190, 101230, 101220, 101220, 101220, 
    101250, 101250, 101280, 101320, 101360, 101410, 101420, 101490, 101550, 
    101560, 101570, 101580, 101580, 101580, 101600, 101630, 101650, 101650, 
    101670, 101680, 101710, 101730, 101740, 101740, 101750, 101770, 101770, 
    101770, 101780, 101800, 101770, 101770, 101760, 101760, 101730, 101710, 
    101680, 101650, 101650, 101640, 101620, 101620, 101600, 101580, 101520, 
    101510, 101470, 101430, 101370, 101370, 101330, 101290, 101270, 101260, 
    101250, 101240, 101240, 101260, 101260, 101270, 101270, 101280, 101270, 
    101280, 101290, 101300, 101320, 101340, 101360, 101370, 101410, 101440, 
    101470, 101510, 101570, 101630, 101700, 101750, 101780, 101830, 101880, 
    101910, 101940, 101970, 102010, 102040, 102070, 102110, 102130, 102130, 
    102120, 102150, 102180, 102190, 102210, 102220, 102160, 102150, 102120, 
    102110, 102170, 102110, 102070, 102020, 101990, 101980, 101970, 101950, 
    101910, 101870, 101820, 101780, 101740, 101710, 101670, 101690, 101620, 
    101520, 101490, 101500, 101580, 101800, 101550, 101530, 101480, 101550, 
    101530, 101510, 101530, 101600, 101620, 101620, 101630, 101610, 101630, 
    101660, 101660, 101660, 101640, 101630, 101630, 101670, 101670, 101680, 
    101670, 101660, 101660, 101640, 101640, 101640, 101690, 101700, 101710, 
    101720, 101650, 101640, 101600, 101570, 101550, 101510, 101520, 101500, 
    101470, 101440, 101400, 101390, 101350, 101300, 101270, 101230, 101170, 
    101140, 101120, 101140, 101120, 101110, 101110, 101100, 101060, 101030, 
    101010, 101010, 101000, 100990, 101000, 100990, 100980, 100980, 100970, 
    100960, 100970, 100950, 100930, 100930, 100900, 100910, 100900, 100900, 
    100920, 100910, 100910, 100900, 100900, 100880, 100860, 100830, 100790, 
    100760, 100740, 100740, 100720, 100710, 100700, 100700, 100710, 100690, 
    100700, 100700, 100700, 100720, 100720, 100740, 100750, 100750, 100770, 
    100790, 100780, 100790, 100800, 100790, 100790, 100800, 100810, 100810, 
    100840, 100840, 100860, 100870, 100860, 100860, 100850, 100860, 100860, 
    100870, 100900, 100900, 100920, 100940, 100930, 100950, 100930, 100910, 
    100910, 100910, 100920, 100940, 100950, 100960, 100970, 100980, 100970, 
    100950, 100980, 100990, 100980, 100980, 100990, 101000, 101020, 101030, 
    101050, 101050, 101060, 101080, 101100, 101110, 101120, 101150, 101170, 
    101180, 101200, 101230, 101250, 101280, 101310, 101330, 101360, 101350, 
    101360, 101370, 101380, 101430, 101430, 101470, 101500, 101500, 101540, 
    101550, 101550, 101550, 101530, 101520, 101520, 101530, 101560, 101590, 
    101620, 101630, 101620, 101620, 101640, 101640, 101680, 101680, 101710, 
    101710, 101740, 101780, 101790, 101830, 101840, 101860, 101870, 101900, 
    101920, 101940, 101960, 102000, 102040, 102080, 102100, 102110, 102140, 
    102130, 102160, 102170, 102170, 102180, 102210, 102220, 102220, 102220, 
    102250, 102240, 102240, 102240, 102230, 102230, 102230, 102210, 102220, 
    102210, 102230, 102230, 102240, 102230, 102220, 102210, 102190, 102160, 
    102120, 102120, 102120, 102120, 102140, 102140, 102180, 102160, 102150, 
    102170, 102190, 102210, 102220, 102230, 102260, 102260, 102290, 102330, 
    102350, 102360, 102370, 102370, 102360, 102370, 102350, 102350, 102350, 
    102360, 102360, 102390, 102390, 102390, 102400, 102390, 102400, 102400, 
    102400, 102390, 102390, 102390, 102390, 102410, 102420, 102440, 102430, 
    102450, 102470, 102470, 102470, 102490, 102500, 102550, 102560, 102620, 
    102640, 102650, 102670, 102670, 102680, 102670, 102630, 102670, 102630, 
    102650, 102630, 102620, 102630, 102600, 102570, 102560, 102490, 102460, 
    102430, 102370, 102340, 102260, 102220, 102180, 102120, 102090, 102040, 
    101970, 101960, 101940, 101940, 101920, 101880, 101890, 101850, 101860, 
    101840, 101800, 101770, 101760, 101720, 101670, 101710, 101710, 101720, 
    101750, 101780, 101810, 101830, 101800, 101780, 101730, 101680, 101670, 
    101620, 101590, 101510, 101430, 101390, 101320, 101280, 101210, 101160, 
    101100, 101030, 100990, 100970, 100950, 100910, 100890, 100890, 100890, 
    100910, 100930, 100950, 100950, 100930, 100950, 100950, 100980, 100990, 
    101010, 101010, 101000, 101030, 101020, 100990, 100930, 100890, 100870, 
    100870, 100860, 100930, 100860, 100860, 100880, 100850, 100820, 100810, 
    100780, 100770, 100780, 100790, 100800, 100770, 100770, 100740, 100740, 
    100760, 100750, 100760, 100770, 100760, 100740, 100750, 100750, 100750, 
    100760, 100760, 100780, 100810, 100840, 100850, 100860, 100850, 100840, 
    100850, 100840, 100840, 100830, 100820, 100810, 100800, 100780, 100760, 
    100750, 100740, 100720, 100710, 100700, 100680, 100650, 100680, 100680, 
    100680, 100670, 100700, 100730, 100750, 100760, 100750, 100760, 100790, 
    100780, 100780, 100770, 100750, 100740, 100740, 100730, 100710, 100700, 
    100680, 100650, 100630, 100640, 100650, 100690, 100710, 100740, 100760, 
    100770, 100770, 100780, 100790, 100780, 100790, 100800, 100830, 100870, 
    100890, 100900, 100950, 100970, 101000, 101010, 101020, 101040, 101060, 
    101090, 101130, 101160, 101200, 101230, 101260, 101280, 101310, 101320, 
    101340, 101340, 101340, 101360, 101390, 101400, 101430, 101440, 101440, 
    101440, 101440, 101430, 101420, 101400, 101380, 101360, 101350, 101350, 
    101360, 101330, 101310, 101310, 101290, 101290, 101270, 101260, 101250, 
    101240, 101240, 101240, 101250, 101260, 101240, 101260, 101270, 101250, 
    101240, 101230, 101200, 101200, 101220, 101230, 101230, 101220, 101240, 
    101250, 101260, 101270, 101270, 101270, 101270, 101270, 101280, 101280, 
    101310, 101330, 101350, 101360, 101370, 101380, 101380, 101400, 101400, 
    101410, 101440, 101460, 101490, 101510, 101530, 101550, 101550, 101570, 
    101580, 101560, 101570, 101570, 101580, 101570, 101600, 101600, 101580, 
    101580, 101560, 101550, 101520, 101490, 101460, 101430, 101390, 101380, 
    101350, 101320, 101300, 101250, 101240, 101210, 101170, 101120, 101080, 
    101060, 101030, 101010, 100980, 100960, 100940, 100890, 100870, 100830, 
    100800, 100760, 100720, 100690, 100690, 100680, 100640, 100640, 100630, 
    100610, 100590, 100570, 100550, 100510, 100500, 100500, 100490, 100480, 
    100480, 100480, 100470, 100480, 100440, 100430, 100390, 100360, 100340, 
    100340, 100310, 100270, 100240, 100220, 100170, 100140, 100080, 100020, 
    99970, 99900, 99830, 99760, 99700, 99650, 99590, 99520, 99470, 99430, 
    99370, 99340, 99300, 99270, 99260, 99290, 99320, 99340, 99390, 99430, 
    99440, 99470, 99510, 99540, 99540, 99560, 99550, 99550, 99570, 99580, 
    99590, 99660, 99690, 99720, 99750, 99810, 99870, 99940, 99970, 100030, 
    100060, 100110, 100160, 100180, 100210, 100240, 100260, 100250, 100290, 
    100310, 100310, 100300, 100320, 100310, 100300, 100300, 100240, 100230, 
    100250, 100220, 100200, 100250, 100310, 100290, 100290, 100320, 100340, 
    100370, 100390, 100420, 100430, 100470, 100510, 100520, 100520, 100580, 
    100670, 100730, 100800, 100850, 100870, 100940, 100960, 100960, 101030, 
    101060, 101120, 101140, 101160, 101180, 101160, 101140, 101120, 101080, 
    101080, 101080, 101000, 100900, 100840, 100770, 100740, 100690, 100590, 
    100560, 100510, 100460, 100440, 100450, 100410, 100370, 100320, 100280, 
    100320, 100290, 100270, 100300, 100330, 100350, 100380, 100440, 100470, 
    100470, 100450, 100450, 100460, 100430, 100400, 100360, 100280, 100330, 
    100370, 100370, 100350, 100370, 100340, 100370, 100390, 100380, 100360, 
    100390, 100400, 100450, 100540, 100610, 100620, 100640, 100660, 100680, 
    100700, 100750, 100780, 100810, 100830, 100840, 100900, 100960, 100990, 
    101060, 101100, 101160, 101210, 101240, 101280, 101320, 101340, 101380, 
    101430, 101470, 101490, 101530, 101550, 101580, 101610, 101620, 101650, 
    101680, 101710, 101720, 101730, 101760, 101760, 101790, 101790, 101810, 
    101830, 101860, 101870, 101860, 101890, 101870, 101860, 101860, 101860, 
    101860, 101820, 101870, 101870, 101850, 101830, 101760, 101710, 101670, 
    101670, 101670, 101630, 101590, 101540, 101520, 101500, 101480, 101530, 
    101510, 101510, 101460, 101450, 101500, 101450, 101500, 101520, 101560, 
    101590, 101640, 101680, 101700, 101690, 101680, 101690, 101730, 101740, 
    101740, 101760, 101780, 101820, 101850, 101860, 101880, 101920, 101940, 
    101930, 101950, 101990, 102020, 102000, 101990, 102020, 102050, 102090, 
    102130, 102160, 102180, 102200, 102210, 102240, 102240, 102240, 102240, 
    102230, 102240, 102260, 102280, 102300, 102300, 102320, 102320, 102320, 
    102310, 102300, 102310, 102320, 102310, 102320, 102310, 102290, 102280, 
    102240, 102230, 102210, 102190, 102180, 102170, 102170, 102180, 102170, 
    102160, 102150, 102150, 102110, 102100, 102110, 102110, 102110, 102110, 
    102090, 102100, 102110, 102110, 102100, 102080, 102060, 102040, 102040, 
    102010, 102270, 102010, 102020, 101990, 101970, 101930, 101900, 101880, 
    101850, 101820, 101800, 101740, 101710, 101680, 101660, 101630, 101590, 
    101570, 101520, 101480, 101460, 101410, 101380, 101350, 101330, 101330, 
    101330, 101320, 101300, 101290, 101270, 101250, 101230, 101240, 101220, 
    101230, 101220, 101210, 101220, 101210, 101190, 101190, 101190, 101180, 
    101180, 101180, 101170, 101160, 101180, 101200, 101200, 101210, 101200, 
    101220, 101220, 101220, 101200, 101210, 101200, 101180, 101180, 101190, 
    101200, 101200, 101200, 101200, 101200, 101200, 101210, 101190, 101190, 
    101180, 101180, 101150, 101170, 101200, 101210, 101210, 101230, 101240, 
    101250, 101260, 101280, 101280, 101290, 101310, 101320, 101340, 101350, 
    101340, 101340, 101330, 101320, 101340, 101330, 101320, 101340, 101370, 
    101420, 101420, 101420, 101420, 101430, 101400, 101380, 101380, 101390, 
    101380, 101360, 101370, 101360, 101370, 101380, 101380, 101400, 101400, 
    101390, 101400, 101400, 101400, 101390, 101400, 101440, 101450, 101450, 
    101430, 101420, 101420, 101440, 101460, 101460, 101470, 101470, 101490, 
    101510, 101520, 101520, 101520, 101530, 101530, 101530, 101530, 101540, 
    101540, 101540, 101560, 101570, 101580, 101580, 101580, 101580, 101600, 
    101590, 101590, 101600, 101600, 101600, 101620, 101630, 101650, 101680, 
    101690, 101690, 101710, 101720, 101730, 101740, 101760, 101760, 101780, 
    101820, 101860, 101870, 101310, 101860, 101880, 101900, 101920, 101950, 
    101990, 102000, 102020, 102040, 102080, 102110, 102110, 102120, 102120, 
    102110, 102110, 102090, 102080, 102060, 102040, 102010, 101990, 101990, 
    101930, 101900, 101860, 101820, 101740, 101690, 101630, 101530, 101450, 
    101380, 101280, 101230, 101170, 101080, 100990, 100880, 100810, 100700, 
    100620, 100570, 100510, 100470, 100450, 100460, 100450, 100450, 100450, 
    100470, 100520, 100590, 100670, 100720, 100770, 100830, 100890, 101000, 
    101060, 101110, 101160, 101210, 101230, 101240, 101260, 101290, 101320, 
    101340, 101350, 101350, 101380, 101380, 101370, 101350, 101340, 101350, 
    101340, 101320, 101320, 101320, 101280, 101280, 101280, 101270, 101230, 
    101190, 101160, 101160, 101150, 101130, 101140, 101140, 101130, 101120, 
    101140, 101120, 101100, 101080, 101080, 101070, 101040, 101020, 101020, 
    101010, 101030, 101050, 101080, 101080, 101100, 101090, 101120, 101130, 
    101120, 101100, 101110, 101120, 101120, 101120, 101140, 101120, 101120, 
    101090, 101070, 101070, 101040, 101040, 101030, 101040, 101040, 101030, 
    101060, 101030, 101010, 101010, 101010, 100990, 100970, 100960, 100960, 
    100970, 100970, 100990, 101000, 100970, 100960, 100950, 100900, 100900, 
    100910, 100910, 100910, 100910, 100940, 100980, 101000, 101000, 101030, 
    101050, 101050, 101070, 101110, 101130, 101160, 101210, 101270, 101290, 
    101320, 101330, 101370, 101390, 101390, 101410, 101430, 101430, 101480, 
    101500, 101530, 101530, 101540, 101550, 101530, 101530, 101540, 101530, 
    101520, 101530, 101510, 101520, 101540, 101550, 101540, 101510, 101480, 
    101470, 101490, 101510, 101530, 101560, 101600, 101610, 101640, 101660, 
    101710, 101780, 101850, 101870, 101870, 101870, 101890, 101900, 101930, 
    101950, 101990, 102000, 102020, 102030, 102030, 102020, 102030, 102050, 
    102080, 102090, 102110, 102150, 102140, 102160, 102170, 102180, 102180, 
    102180, 102170, 102170, 102180, 102200, 102210, 102230, 102250, 102260, 
    102270, 102280, 102260, 102280, 102280, 102290, 102310, 102330, 102370, 
    102420, 102460, 102520, 102560, 102590, 102640, 102670, 102690, 102710, 
    102760, 102810, 102830, 102880, 102940, 102970, 102980, 103000, 103050, 
    103050, 103080, 103090, 103100, 103140, 103150, 103180, 103200, 103220, 
    103240, 103240, 103230, 103240, 103230, 103220, 103210, 103190, 103180, 
    103190, 103210, 103200, 103190, 103190, 103190, 103170, 103160, 103170, 
    103170, 103170, 103170, 103180, 103200, 103220, 103230, 103270, 103280, 
    103270, 103270, 103270, 103270, 103280, 103280, 103270, 103270, 103270, 
    103250, 103240, 103230, 103220, 103180, 103190, 103180, 103140, 103120, 
    103100, 103090, 103070, 103050, 103010, 102950, 102900, 102870, 102810, 
    102770, 102740, 102710, 102680, 102630, 102620, 102590, 102550, 102510, 
    102480, 102470, 102430, 102430, 102410, 102390, 102370, 102320, 102310, 
    102280, 102260, 102220, 102190, 102150, 102120, 102080, 102060, 102060, 
    102040, 102020, 102020, 102010, 102000, 101970, 101950, 101950, 101940, 
    101990, 102020, 102050, 102080, 102130, 102170, 102190, 102210, 102240, 
    102250, 102270, 102270, 102280, 102310, 102310, 102310, 102320, 102330, 
    102310, 102330, 102320, 102310, 102290, 102260, 102240, 102230, 102180, 
    102170, 102180, 102180, 102160, 102150, 102150, 102130, 102110, 102100, 
    102090, 102070, 102080, 102080, 102060, 102060, 102050, 102040, 102030, 
    102020, 102000, 102010, 102000, 101990, 101990, 101990, 102010, 102010, 
    102020, 102020, 102020, 102010, 102010, 102010, 102000, 102000, 102000, 
    101990, 101980, 101980, 101970, 101950, 101950, 101940, 101940, 101910, 
    101940, 101930, 101940, 101940, 101960, 101960, 101940, 101950, 101940, 
    101920, 101900, 101890, 101890, 101890, 101870, 101850, 101850, 101850, 
    101830, 101810, 101780, 101760, 101750, 101720, 101710, 101710, 101700, 
    101700, 101710, 101740, 101750, 101760, 101760, 101770, 101790, 101790, 
    101790, 101790, 101800, 101800, 101800, 101810, 101810, 101790, 101810, 
    101800, 101810, 101790, 101800, 101800, 101800, 101790, 101800, 101810, 
    101810, 101800, 101780, 101770, 101750, 101720, 101700, 101680, 101660, 
    101640, 101620, 101610, 101590, 101570, 101550, 101530, 101510, 101530, 
    101530, 101530, 101540, 101580, 101610, 101610, 101630, 101640, 101650, 
    101640, 101650, 101630, 101640, 101650, 101660, 101670, 101690, 101700, 
    101710, 101700, 101680, 101660, 101660, 101650, 101630, 101610, 101610, 
    101610, 101610, 101610, 101610, 101610, 101610, 101590, 101590, 101590, 
    101600, 101590, 101610, 101600, 101600, 101620, 101620, 101620, 101630, 
    101620, 101620, 101630, 101630, 101630, 101630, 101650, 101640, 101660, 
    101670, 101680, 101690, 101690, 101680, 101670, 101660, 101650, 101650, 
    101660, 101660, 101680, 101700, 101700, 101710, 101720, 101740, 101740, 
    101730, 101710, 101710, 101730, 101740, 101770, 101770, 101770, 101770, 
    101770, 101770, 101750, 101740, 101740, 101750, 101750, 101750, 101730, 
    101750, 101740, 101750, 101740, 101720, 101710, 101690, 101720, 101720, 
    101760, 101750, 101770, 101730, 101740, 101740, 101740, 101730, 101720, 
    101710, 101680, 101650, 101640, 101630, 101630, 101610, 101580, 101550, 
    101520, 101500, 101490, 101490, 101480, 101470, 101480, 101490, 101470, 
    101480, 101480, 101490, 101470, 101460, 101430, 101420, 101400, 101390, 
    101370, 101370, 101370, 101350, 101340, 101330, 101290, 101280, 101270, 
    101250, 101250, 101230, 101210, 101230, 101180, 101190, 101190, 101170, 
    101120, 101110, 101060, 101040, 101010, 100980, 100950, 100930, 100900, 
    100880, 100850, 100800, 100760, 100730, 100660, 100610, 100550, 100480, 
    100470, 100470, 100390, 100370, 100280, 100190, 100160, 100120, 100080, 
    100080, 100070, 100070, 100050, 100040, 100030, 100010, 99980, 99950, 
    99920, 99910, 99890, 99840, 99820, 99790, 99760, 99740, 99740, 99720, 
    99700, 99700, 99690, 99680, 99660, 99650, 99650, 99640, 99620, 99630, 
    99610, 99580, 99570, 99560, 99570, 99560, 99570, 99580, 99590, 99610, 
    99630, 99660, 99680, 99720, 99730, 99750, 99750, 99760, 99760, 99750, 
    99770, 99780, 99790, 99800, 99810, 99810, 99810, 99790, 99750, 99720, 
    99690, 99680, 99680, 99680, 99690, 99700, 99740, 99750, 99760, 99790, 
    99810, 99820, 99870, 99890, 99930, 99930, 99970, 100010, 100040, 100070, 
    100100, 100130, 100150, 100150, 100180, 100210, 100250, 100270, 100280, 
    100310, 100360, 100390, 100420, 100440, 100460, 100470, 100490, 100510, 
    100530, 100560, 100570, 100590, 100610, 100630, 100650, 100660, 100680, 
    100690, 100720, 100720, 100730, 100750, 100770, 100780, 100800, 100810, 
    100820, 100820, 100820, 100840, 100840, 100830, 100850, 100870, 100870, 
    100850, 100850, 100850, 100830, 100850, 100860, 100840, 100830, 100830, 
    100810, 100780, 100780, 100770, 100750, 100720, 100690, 100660, 100620, 
    100600, 100560, 100520, 100480, 100410, 100360, 100290, 100230, 100200, 
    100140, 100100, 100070, 100050, 100010, 100000, 100010, 99990, 99990, 
    100030, 100020, 100040, 100090, 100130, 100160, 100210, 100280, 100350, 
    100390, 100450, 100510, 100570, 100640, 100710, 100750, 100840, 100880, 
    100910, 100980, 101030, 101050, 101110, 101160, 101210, 101250, 101290, 
    101330, 101370, 101390, 101400, 101410, 101420, 101440, 101450, 101460, 
    101480, 101490, 101490, 101490, 101500, 101510, 101500, 101490, 101500, 
    101500, 101520, 101520, 101540, 101550, 101570, 101580, 101570, 101570, 
    101590, 101520, 101580, 101620, 101640, 101650, 101670, 101720, 101710, 
    101720, 101720, 101720, 101730, 101750, 101760, 101790, 101800, 101820, 
    101810, 101820, 101830, 101820, 101840, 101590, 101700, 101740, 101780, 
    101800, 101850, 101870, 101870, 101860, 101850, 101850, 101840, 101820, 
    101800, 101770, 101730, 101710, 101700, 101690, 101680, 101660, 101660, 
    101660, 101630, 101610, 101600, 101590, 101570, 101750, 101570, 101570, 
    101550, 101560, 101550, 101550, 101550, 101540, 101530, 101530, 101550, 
    101560, 101570, 101640, 101670, 101690, 101710, 101730, 101740, 101770, 
    101790, 101830, 101550, 101600, 101860, 101900, 101950, 101980, 102020, 
    102040, 102040, 102050, 102030, 102030, 102040, 102050, 102060, 102040, 
    102030, 102040, 101920, 101880, 101930, 101990, 102030, 102060, 102040, 
    101800, 101720, 101710, 101640, 101620, 101540, 101440, 101400, 101350, 
    101300, 101190, 101130, 101060, 100980, 100970, 100930, 100870, 100830, 
    100800, 100750, 100720, 100690, 100680, 101740, 101240, 100640, 100630, 
    100630, 100630, 100670, 100710, 100730, 100740, 100730, 100710, 100680, 
    100660, 100670, 100700, 100740, 100760, 100790, 100830, 100860, 100860, 
    100880, 100880, 100920, 100930, 100930, 100940, 100950, 100930, 100920, 
    100920, 100870, 100870, 100830, 100770, 100740, 100690, 100620, 100590, 
    100530, 100510, 100470, 100450, 100410, 100390, 100370, 100330, 100320, 
    100310, 100290, 100330, 100320, 100290, 100310, 100310, 100270, 100230, 
    100230, 100220, 100200, 100200, 100210, 100210, 100190, 100160, 100150, 
    100220, 100230, 100260, 100250, 100260, 100220, 100290, 100300, 100350, 
    100380, 100410, 100450, 100490, 100490, 100530, 100550, 100560, 100570, 
    100580, 100630, 100660, 100660, 100670, 100680, 100670, 100670, 100660, 
    100670, 100660, 100640, 100590, 100610, 100650, 100630, 100620, 100610, 
    100610, 100600, 100590, 100580, 100580, 100580, 100580, 100610, 100610, 
    100600, 100600, 100660, 100650, 100610, 100610, 100610, 100600, 100580, 
    100590, 100570, 100610, 100600, 100600, 100530, 100540, 100520, 100510, 
    100500, 100530, 100500, 100480, 100480, 100510, 100580, 100510, 100540, 
    100490, 100500, 100470, 100440, 100410, 100380, 100360, 100340, 100320, 
    100310, 100220 ;

 wind_from_direction_10m = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, 327, 310, _, _, 332, 316, 299, 14, 328, 339, 344, 324, 
    311, 322, 332, 308, 311, 326, 343, 343, 302, 312, 346, 300, 327, 0, 340, 
    334, 73, _, 78, 68, 32, 31, 31, 34, 31, 32, 43, 43, 29, 28, 358, 353, 1, 
    299, 262, 280, 20, 268, 30, 356, 45, 34, 41, 38, 34, 26, 30, 37, 180, 
    220, 109, 329, 131, 191, 271, 355, 16, 150, 215, 131, 2, 278, _, _, 353, 
    318, 308, 304, 303, 304, 314, 308, 313, 305, _, _, _, _, _, _, _, _, _, 
    318, 317, 325, 314, 350, 308, _, 309, 323, 312, 324, 316, 315, 315, 310, 
    309, 282, 289, 298, 321, 325, 320, 322, 302, 326, 319, 329, _, 319, 311, 
    313, 307, 325, 303, 264, _, _, 91, 86, 82, 86, 93, 67, 93, 89, 95, 97, 
    102, 90, 100, 100, _, _, 88, 82, 79, 84, 91, 92, 86, 86, 94, 78, 92, 93, 
    98, 95, 92, 93, 97, 95, 94, 93, 91, 84, 82, 85, 83, _, 83, 98, 86, 93, 
    117, 121, 123, 96, 107, 95, 90, 90, 96, 94, 98, 98, 98, 94, 99, 92, _, 
    89, 88, 262, 316, 90, 85, 82, 86, 81, 61, 9, 5, 63, 59, 311, 9, 78, 86, 
    64, 81, 70, 64, 44, 49, _, 52, 52, 50, 285, 59, 51, 63, 66, 87, 69, 71, 
    97, 102, 98, 75, 63, 72, 69, 64, 68, 64, 69, 49, 328, 330, 301, 324, 294, 
    346, 66, 295, 306, 303, 291, 297, 308, 295, 262, 344, _, 80, 70, 67, 68, 
    92, 84, _, 63, 55, 65, 70, 75, 74, 69, 76, 74, 68, 78, 68, 58, 129, 317, 
    191, 262, 313, 304, 332, 20, 315, 292, 329, _, 7, 313, 357, 333, 3, 331, 
    0, 334, 344, 303, 45, 300, 302, 35, 323, 331, 328, 342, 318, 321, _, 0, 
    327, 333, 42, 312, 359, 32, 321, 78, 344, 306, 323, 336, 338, 303, 25, 
    331, 359, _, 329, 344, 326, 306, 49, 8, _, 360, 36, 69, 51, 292, 353, 
    311, 330, 344, 308, 66, 59, 346, 4, 39, 356, 331, 54, 332, 22, 24, 314, 
    288, 312, 322, 311, 304, 341, 328, 305, 60, 293, 321, 331, 330, 292, 19, 
    308, 10, 344, 359, 318, 335, 306, 337, _, 353, 344, 352, 305, 329, 336, 
    333, 313, 352, 307, 271, 33, 300, 299, 313, 66, 358, _, _, 72, 0, 335, 
    83, 358, 19, 308, 360, 343, 337, 325, 331, 288, 313, 292, 16, 301, 299, 
    294, 305, 299, 308, 301, 297, 303, 301, 295, 341, 298, 341, 319, 322, 
    341, 327, 34, 351, 341, 85, 305, 1, 308, 358, 4, 318, 328, 100, 60, 355, 
    351, 314, 342, 85, _, 357, 40, 346, 325, 350, 333, 18, 330, 321, 20, 82, 
    90, 95, 100, 98, 97, 95, 71, 72, 93, 84, 72, 68, 84, 164, _, 307, 35, 
    336, _, _, 311, 3, 95, 310, _, 86, 319, 296, 296, 73, 344, 359, 312, 323, 
    352, 354, 360, 345, 290, 332, 305, 267, 97, 155, 155, 47, 68, 42, 308, 
    314, 295, 25, 323, 14, 64, 331, 48, 70, 318, 311, 301, 307, 334, 327, 42, 
    331, 91, 2, 1, 315, 300, 328, 349, 344, 1, 304, 354, 323, 57, 34, 17, 
    325, 324, 296, 3, 342, 311, 356, 314, 344, _, 318, _, 40, 303, 36, 311, 
    317, 323, 6, 310, 348, 31, 334, 348, 8, 341, 314, 308, 326, _, 300, 348, 
    0, 333, 343, 35, 324, 334, 327, 324, 0, 330, 339, 32, 286, 358, 348, 315, 
    11, 26, 0, _, 324, 355, 29, 43, 44, 332, 353, 333, 316, 96, 54, 328, 291, 
    320, 360, 344, 302, 5, 314, 37, 305, 301, 318, 348, 325, 357, 343, 327, 
    19, _, 342, 328, 320, 0, 314, 311, 306, 10, 351, 337, 4, 297, 290, 290, 
    49, 47, 35, 42, 35, 33, _, 34, 37, 39, 35, 52, 56, 49, 48, 56, 42, 51, 
    27, 320, 280, 4, 170, 354, 291, 314, 359, _, 18, 54, 25, 348, 342, 326, 
    307, 302, 315, 320, 306, 308, 317, 309, 332, 310, 348, 335, 323, 273, 
    302, 295, _, 276, 311, 325, 331, 1, 0, 0, 70, 270, 283, 292, 297, 290, 
    297, 312, 331, 311, 36, 323, 346, 306, 49, 315, 306, _, 305, 305, _, 291, 
    340, 349, 19, 311, _, 311, 76, 319, 307, 352, 316, 326, 310, 309, 100, 
    313, 351, 313, 2, _, 22, 37, 298, 302, 309, 248, 303, 239, 255, 275, 290, 
    346, 132, 4, 56, 295, 284, 290, 290, 284, 283, 300, _, 287, 293, 285, 
    272, 273, 281, _, 273, 280, 287, 288, 280, 255, 278, 300, 287, 296, 299, 
    307, 324, 311, 298, 279, 320, _, 204, _, _, 315, _, 291, 352, 303, 316, 
    284, 342, 322, 316, 303, 324, 275, 314, 316, 290, 305, 312, _, 319, 348, 
    13, 353, 21, 353, 348, 98, 211, 44, 303, 327, 359, 355, 36, 29, 49, 45, 
    38, 29, 40, 10, 299, 298, _, 281, 303, 312, 320, 317, 327, 321, 306, 303, 
    316, 312, 296, 260, 318, 3, 317, 305, 334, 266, 290, 327, 359, 5, 356, 
    279, 320, 325, _, 279, 327, 316, 306, 288, 336, 300, 352, 334, 347, 357, 
    352, 359, 21, 10, 1, 6, 22, 11, 14, 6, 317, 316, 305, 300, 316, 319, 304, 
    316, 348, 323, 322, 337, 270, 284, 319, 304, 317, 308, 331, 323, 314, 
    315, 337, 323, 345, 5, 47, 317, 299, 303, 315, 325, 320, 293, 320, 26, 
    320, 39, 355, 334, 346, 328, 315, _, 342, 43, 359, 30, 19, 57, 60, 152, 
    214, 191, 238, 184, 337, 149, 305, 300, 310, 310, 295, 314, 319, 320, 
    283, 307, 323, 307, 297, 301, 321, 283, 245, 247, 235, 285, 204, 286, 
    299, 289, 279, 46, 342, _, 314, 308, 301, 290, 303, 48, 313, 294, 48, 
    359, 94, 84, 96, 94, 93, 85, 87, 82, 105, 106, 98, 97, 96, 85, 92, 96, 
    98, 100, 97, _, _, 96, 98, 97, 98, 98, 98, 97, 94, 96, 96, 100, 99, 93, 
    97, 96, 94, 94, 94, 92, 83, 78, 83, 79, 80, 88, 90, 88, 89, 85, 88, 78, 
    87, 88, 92, 90, 95, 77, 84, 79, 85, 90, 86, 75, 86, 111, 84, _, _, 50, 
    114, 294, 113, 84, 87, 75, 74, 77, 74, 79, 80, 78, 89, 64, 73, 104, 82, 
    64, 77, 84, 72, 70, _, 100, 89, 324, 16, 330, 341, 351, 325, 101, 356, 
    331, 341, 314, 122, 75, 89, 94, 114, 116, 112, 109, 112, 98, 96, 91, 93, 
    _, 348, 321, 324, 1, 281, 325, 327, 317, 325, 329, 325, 5, 332, 324, 323, 
    37, 359, 0, 308, 82, 21, 30, 2, 333, 284, 77, 295, 96, 22, 17, 303, 360, 
    349, 90, 337, 101, 144, 143, 94, 124, 114, 73, 76, _, _, 283, 12, 17, 
    291, 318, 291, 354, 346, 347, 314, 48, 87, 16, 0, 0, 92, 73, 298, 48, 
    291, 307, 329, 296, 275, 281, 296, 292, _, 266, 290, 300, 293, 300, 280, 
    295, 309, 305, 300, 300, 308, 313, 305, 330, 286, 320, 307, 318, 352, 
    349, 298, 308, 335, 314, 33, 313, 306, 46, 289, 317, 335, 324, 4, 310, 
    311, 295, 287, 301, 307, 315, 304, 307, _, _, 332, 300, 293, 107, 330, 
    316, 297, 304, 332, 311, 346, 34, 346, 326, 72, 27, 335, 321, 318, 3, 
    318, 298, 300, 294, 326, 340, _, 36, 359, 56, 286, 295, 282, 287, 295, 
    251, 262, 285, 286, 299, 287, 296, _, 287, 283, 291, 286, 253, 286, 313, 
    294, 289, 314, 291, 292, 309, 293, 278, 271, 273, 285, 295, 307, 305, 
    294, 10, 348, 312, 323, 13, _, _, 314, 322, 28, 320, 58, 295, 357, 12, 
    347, 356, 321, 306, 301, 327, 311, 300, 318, 286, 304, 296, 300, 305, 68, 
    291, 307, _, 2, 132, 245, 29, 317, 154, 75, 350, 334, 331, 298, 301, 272, 
    299, 333, 343, 317, 346, 318, 350, 321, 296, 6, 308, 332, 1, 315, 306, 
    352, 317, 301, 359, 313, 17, 323, 349, 344, 351, 319, 18, 355, 311, 350, 
    8, _, 336, 26, 339, 315, 322, 98, 17, 329, 346, 334, 69, 313, 309, 312, 
    335, 342, 308, 306, 329, 299, 324, 84, 83, 84, 87, 88, _, 88, _, 319, 
    300, 319, 280, 293, 292, 310, 304, 290, 299, 286, 332, 327, 60, _, 352, 
    77, 333, _, 276, 337, 340, 1, 61, 295, 329, 294, 74, 42, 39, 332, 276, 
    28, 209, 23, 17, 28, 34, 50, 43, 27, 57, _, 71, 307, 290, 268, 321, 302, 
    308, 290, 341, 352, 355, _, 47, 353, 19, 1, 304, 359, 29, 337, 320, 317, 
    320, 324, 356, 284, 325, _, _, 39, 337, 16, 304, 318, 346, 311, 335, 320, 
    22, 308, 322, 345, 0, 358, 268, 319, 349, _, 109, 317, 315, 346, 296, 
    274, 3, 250, 104, 58, _, 325, 302, 304, 306, 316, 328, 2, 74, 19, 106, 
    106, 103, 104, _, 111, 109, 115, 58, 68, 1, 55, 46, 56, 354, 281, 320, 
    304, 300, 311, 332, 332, 322, 71, 284, 118, 97, 160, 36, 359, 27, 6, 33, 
    320, 269, 84, 63, 253, 64, 46, 36, 49, _, 359, _, 353, 27, 338, 343, 118, 
    241, _, 28, 42, 45, 46, 73, 1, 57, 47, 43, 41, 47, 52, 61, 45, 55, 74, 
    67, 25, 310, 318, 290, 331, 304, 183, _, 284, 324, 318, 325, 331, 345, 
    321, 358, 347, 10, 333, 347, 318, 299, 312, 348, 315, 5, 346, 291, _, 
    342, 305, 81, 57, 289, 311, 313, 309, 314, 310, 342, 342, 319, 299, 343, 
    315, 318, 310, _, 312, 311, 321, 285, 298, 286, _, 320, 310, 318, 324, 
    297, 313, 289, 325, 306, 334, 314, 313, 310, 317, 340, 330, 301, 320, 
    336, 320, 306, 310, 334, _, _, 321, 321, 311, 322, 333, 330, 329, 331, 
    314, 330, 314, 310, 298, 11, 317, 331, 359, 339, 331, 310, 328, 313, 312, 
    314, 306, 12, 359, 355, 312, 356, 0, 310, 299, _, 323, 334, 310, 313, 
    320, _, 354, 287, _, 304, 354, 313, _, 324, 346, 359, 318, 338, 300, 62, 
    342, 6, 332, 303, 28, 358, 360, 305, 353, 8, 305, 342, 342, 359, _, _, 
    301, _, _, 356, _, 327, 54, 340, _, _, 346, 349, _, _, 324, 323, 324, 
    319, _, 334, 325, 315, 329, 287, 4, 303, 302, 328, 359, 337, 78, 304, 
    308, 349, 327, 302, 40, 305, 59, 52, 80, _, 66, 91, 62, 62, 69, 50, 56, 
    34, 97, 108, 69, 92, 71, 66, 56, 68, 48, 303, 265, 2, 337, 303, 306, 308, 
    323, 320, 325, 324, 38, 10, _, 302, 323, 350, 359, 288, 334, 17, 341, 
    355, 320, 21, 358, 333, 35, 1, 311, 328, 3, 0, 310, 343, 310, 27, 29, 
    344, 346, 2, 70, 322, 3, 3, 345, 343, 326, 20, 344, 310, 53, 5, 327, 342, 
    49, 338, 353, 64, 355, 58, 342, 46, 333, 89, 0, 60, 50, 5, 19, 21, 333, 
    72, 305, 299, 356, 338, 301, 324, 20, 316, 17, 87, 86, _, 294, 274, _, 
    333, 12, 337, 309, 283, 318, 340, 307, 282, 316, 44, 48, 339, 325, 4, 10, 
    353, 329, 331, 305, 333, 77, 316, 88, 59, 323, 20, 62, 13, 37, 323, 298, 
    14, 321, 359, 55, 356, 97, 347, 25, 320, 22, 357, 349, 352, 360, 42, 315, 
    2, _, 340, 84, 324, 304, 301, 292, 300, 89, 325, 320, 68, 21, 331, 340, 
    324, 26, 316, 337, 103, 0, 77, 67, 0, 18, 292, 34, 303, 301, 314, 332, 
    314, 339, 84, 24, 0, 297, 324, 335, 314, 356, 333, 48, 333, 307, 85, 356, 
    310, 353, 332, 5, 355, 325, 28, 76, 86, 358, 7, 340, 3, 322, 334, 322, 
    304, 311, 327, 323, 320, 313, 316, 0, 346, _, 294, 311, 307, 300, 181, 
    356, 99, 114, 300, 297, 288, 319, 327, 241, 353, 5, 322, _, 332, 0, 317, 
    321, 318, 326, 304, 85, 348, 286, 343, 319, 313, 0, 313, 73, 356, 354, 6, 
    298, 296, 301, 313, 311, 305, 328, 313, 346, 305, 301, 328, 275, 255, 
    350, 19, 355, 70, 315, 106, 86, 327, 283, 341, 339, 291, 250, 273, 286, 
    299, 293, 301, 297, 296, _, 298, 294, 303, 303, 324, 309, 329, 303, 346, 
    307, 317, 357, 338, 66, 314, 0, 339, _, 66, 45, 356, 303, 341, 347, 312, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 307, 333, 339, 34, 74, 
    97, 58, 50, 211, 261, 40, 29, 359, 200, 276, 217, 180, 321, 327, 331, 
    329, 315, _, 310, 304, 344, 341, 322, 303, 348, 43, 319, 315, 343, 315, 
    315, 295, 360, 10, 321, 310, 88, 0, 0, 342, 102, 337, 71, 54, 350, 115, 
    330, 19, 329, 13, 322, 291, 44, 359, 332, 348, 330, 13, 5, 311, 310, 316, 
    293, 155, 344, _, 34, 35, 44, 38, 41, 53, _, 39, 57, 49, 27, 20, 353, 21, 
    26, 18, 15, 354, 359, 306, 354, 305, 329, 1, 54, 15, 359, 311, 280, 313, 
    318, 327, 308, 301, _, 354, 307, 286, 344, 338, 0, 351, 343, 348, 350, _, 
    30, 74, 86, 80, 73, 66, 61, 57, 67, 48, 58, 61, 53, 18, 12, 10, 32, 67, 
    28, 21, 4, 283, _, 275, 356, _, 328, 330, 343, 349, 307, 308, 320, 304, 
    313, 325, 315, 330, 352, 325, 329, 339, 18, 306, 313, 286, 347, 305, 276, 
    348, 275, 329, 44, 82, 85, 87, 93, 104, 96, 83, 80, 92, 82, 80, 58, 65, 
    82, 64, 47, 47, _, 25, _, 305, 303, 349, 323, 307, 312, 18, 49, 346, 334, 
    344, 323, 327, 311, 53, 299, 323, 0, 11, 319, 46, 341, 352, _, 306, 302, 
    10, 318, 312, 332, 11, 342, 36, 340, 315, 357, 360, 36, _, 309, 109, 330, 
    10, 311, 346, 323, 0, 62, 359, 326, 356, 325, 71, 90, 80, 98, 104, 98, 
    91, 65, 85, 99, 91, 97, 322, 315, 280, 297, 292, 321, 318, _, 313, 317, 
    314, 314, _, 338, 314, 334, 330, 359, 307, 16, 339, 329, 59, 338, 356, 1, 
    70, 326, 75, 330, 320, 42, 327, 53, 342, _, 311, 92, 93, 96, 93, 87, 85, 
    89, 90, 89, 89, 86, 88, 50, 70, 76, 79, 86, 73, 90, 75, 295, 293, 299, 
    318, 334, 285, 325, 77, 315, 9, 326, 359, 0, 0, 306, 4, 16, 46, 310, 319, 
    77, 46, 339, 320, 28, 94, 333, 2, 344, 322, 77, 350, 332, 343, 346, 236, 
    2, 0, 320, 0, 65, 326, 80, 313, 359, 47, 323, 332, 316, _, 0, 306, 336, 
    326, 43, 317, 22, 4, 2, 109, 95, 280, 323, 319, 319, 42, 30, 52, 21, 64, 
    69, 48, 66, 330, 56, 22, 335, 30, 320, 295, 330, 324, 308, 9, 83, 77, 90, 
    42, 39, 39, 59, 88, 66, 323, _, 319, 3, 311, 321, 357, 324, 310, 308, 
    311, 345, 99, 205, 28, 305, 148, 328, 303, 317, 321, 131, 10, 67, 326, 
    353, 65, 348, 88, 83, 111, 44, 48, 55, 88, 60, 45, 122, 137, 137, 110, 
    95, 301, 109, 117, 59, 87, 57, 61, 95, 61, 67, 43, 22, 50, 353, 10, 11, 
    5, 335, 279, 318, 356, 314, 316, 310, 306, 293, 311, 312, 59, 353, 300, 
    273, _, 349, 318, 8, 349, 335, 0, 347, 358, 1, 29, 352, 349, 75, 343, 18, 
    25, 343, 338, 355, 51, 345, 301, 7, 324, 10, _, 349, 6, 17, 345, 324, 12, 
    66, 297, 341, 15, 326, 0, 312, 357, 315, _, 321, 277, 305, 68, 305, 351, 
    315, 333, 342, 291, 230, 181, 318, 279, 213, 312, 335, 51, 33, 45, 44, 
    24, 57, 8, 70, 41, 14, 211, _, _, 47, 26, 276, 30, 146, 351, 293, 305, _, 
    80, 73, 97, 27, 355, 343, 295, 354, 32, 97, 10, 8, 313, _, _, 273, _, 
    341, _, _, _, _, _, 299, 28, 305, 320, 327, _, 307, 47, 49, 333, 337, 
    323, 31, 219, _, 24, 32, 19, 346, 20, 274, 188, 152, 336, 304, 285, 190, 
    340, 77, 42, 355, 13, 297, 328, 19, 22, 345, 296, 316, 315, 3, 5, 21, 
    354, 55, 310, 359, 0, 320, 4, 322, 103, 67, 334, 296, 260, 6, 19, 33, 
    143, 79, 182, 68, 15, 349, _, 339, 336, 332, 334, 10, _, 291, 292, 348, 
    318, 352, 15, 0, 328, 41, 345, 342, 2, 3, 343, _, 24, 348, 0, 16, 34, 26, 
    303, 330, 290, 297, 297, 319, 290, 327, 61, 352, 308, 311, 324, 24, 37, 
    24, 35, _, 317, 343, 53, 347, 63, 310, 304, 37, 17, 30, 71, 29, 8, 346, 
    41, 59, 357, 49, 336, 62, 326, 346, 42, 85, 348, 329, _, 21, 79, 78, 30, 
    22, 344, 323, 77, 61, 338, 331, 300, 329, 350, 28, 87, 69, 313, 323, 87, 
    _, 75, 75, 81, 81, 79, 80, 80, 77, 87, 84, 94, 67, 77, 95, 95, 57, 86, 
    71, 67, 58, 101, 99, 99, _, 89, 99, 104, 122, 71, 68, 318, 338, 40, 118, 
    272, 14, 206, 151, 68, 341, 337, 337, 329, 348, 332, 348, 357, 57, 353, 
    326, 357, 323, 16, 2, 325, 356, 314, 295, 12, 65, 101, 65, 12, 353, 60, 
    325, 341, 339, 28, 334, 349, _, 28, 107, 316, 0, 30, 344, 357, 313, 354, 
    356, 45, 356, 89, 0, 94, 326, 22, 0, 321, 43, 56, 325, 94, _, _, 16, 352, 
    30, 314, 27, 130, 317, 102, 1, 330, 90, 320, 137, 359, 35, 298, 350, 104, 
    20, 324, 3, 136, 300, 261, 60, 65, 17, 31, 73, 209, 197, 38, 42, 45, 27, 
    29, 46, 50, 16, _, 33, 22, 162, 296, 292, 27, _, 226, 43, 47, 53, 204, 
    43, 13, 21, 352, 47, 148, 210, 35, 18, 271, 16, 324, 12, 343, 324, 303, 
    341, _, _, _, 327, 307, 308, 313, 356, 343, 330, 302, 356, 356, 359, 347, 
    0, 0, 341, 348, 93, 357, 20, 63, 23, 74, 286, 351, 286, 40, _, _, 350, 
    295, 277, 281, 242, 306, 99, 243, 226, 284, 189, 238, 228, 357, 51, 89, 
    106, 175, _, 20, 41, 58, 66, 87, 57, 56, 68, 64, 111, 84, 64, 76, 90, 70, 
    102, 37, 79, 72, 66, 70, 76, 89, _, 74, 86, 89, 73, 74, 60, 73, 94, 15, 
    83, 79, 74, 69, 68, 69, 77, 75, 73, 17, 343, 302, 325, 310, 313, 329, 
    279, 324, 307, 346, 303, 279, 313, 326, 325, 92, 325, 117, 333, 11, 352, 
    337, 349, 345, 0, 324, 5, 337, _, 294, 297, 331, 310, 307, 2, 1, 36, 301, 
    343, 50, 36, 51, 56, 263, 247, 248, 308, 351, 321, 2, 307, 322, _, 52, 
    350, 172, 259, 307, 304, _, 331, 294, 300, 287, _, 5, _, 46, 350, 333, 
    37, 349, 9, _, _, 28, 0, 0, 0, 0, 14, 0, 339, 85, 1, 312, 126, 0, 356, 
    88, 334, 22, _, _, 321, 43, 344, 66, 359, 101, _, 336, 76, 339, 312, 329, 
    108, 0, 89, 359, 100, 81, 360, 315, 12, 36, 302, 329, 349, _, 87, 321, _, 
    _, _, 313, 354, 0, 25, 74, 307, 8, 323, 280, 305, 71, 101, 2, 336, 90, 5, 
    352, 288, 325, 331, 87, 355, 104, 341, 305, 261, 302, 264, 328, 140, 263, 
    319, 255, 53, 357, 357, 6, 21, 21, 13, 36, 28, 110, 21, 19, 17, 13, _, 
    42, 60, 65, _, 67, 171, 39, 36, 41, 80, 38, 35, _, 44, 29, 43, 35, 94, 
    343, 342, 359, _, 267, _, 341, 357, 51, 61, 360, 360, 268, 348, 49, 302, 
    317, 207, 296, 340, _, 46, 43, 40, 42, 43, 12, _, 43, 27, 31, 27, 33, 38, 
    30, 22, 32, 16, 15, 168, 199, 120, 222, 272, 107, 28, 66, 37, 317, 278, 
    191, 302, 2, _, 23, 23, 356, _, 345, 283, 275, 280, 101, 321, 196, 49, 
    62, 39, 49, 69, 35, 35, 37, 63, 156, _, 283, 26, 25, 304, 334, 345, 337, 
    328, 317, 323, 283, 281, 266, 260, 272, 282, 283, 281, 328, 329, 304, 
    347, 319, 357, 7, 33, 14, 2, 349, 342, 357, 79, 138, 343, 1, 295, 294, 4, 
    256, 335, 220, 223, 266, 338, 276, 101, 238, 123, 216, 211, 147, 98, 220, 
    224, 21, 323, 146, 171, 131, 153, 288, 98, 158, 62, 235, 128, 12, 348, 
    306, 330, 316, 74, 325, 17, 359, 0, 62, 20, 0, 46, 337, 0, 0, 312, 111, 
    12, 130, 349, 356, 1, 315, 0, 335, _, 23, _, 356, 299, 2, 310, 106, 306, 
    317, 115, 0, 39, 349, 358, 9, 165, 0, 343, 297, 297, 107, 313, 0, 352, 
    51, 354, 0, 94, 314, 63, 0, 0, 348, 7, 359, 88, 0, 358, 268, 305, 341, 
    346, 359, 346, 32, 14, 333, 322, 292, 286, 329, _, 25, 16, 74, 310, 329, 
    48, _, _, 119, 354, 277, 286, 279, 307, 295, 41, 346, _, 0, _, 358, 344, 
    344, 345, 350, 331, 2, 348, 325, 15, 68, 111, 82, 355, 358, 336, 262, 
    305, 351, 317, 314, 299, 297, 336, 320, 309, 4, 285, 346, 2, 37, 105, 34, 
    327, 355, 239, 231, 288, 185, 157, 32, 210, 189, 190, 200, 207, 348, 320, 
    333, 354, 349, 345, 354, 336, 355, 2, 91, 126, 133, 131, 190, 178, 157, 
    161, 173, 196, 89, _, 89, 43, 354, _, 323, 289, 327, 1, 324, 7, 10, 359, 
    329, 325, 0, 322, 0, 215, 193, 268, 281, 261, 275, 305, _, _, _, 14, 355, 
    358, 22, 345, 332, 68, 26, 0, 63, 359, 100, 5, 14, 273, 0, 277, 311, 322, 
    348, 311, 297, 41, _, 44, 316, 336, 358, 36, 0, 356, 84, 348, 37, 60, 3, 
    331, 355, 305, 13, 0, 293, 0, 6, 344, 131, 69, 70, 88, 82, _, _, 88, 79, 
    75, 76, 99, 67, 98, 69, 110, 56, _, 359, 293, 311, 303, 308, 294, 77, 
    250, 277, 315, 314, 307, 79, 289, 300, 286, 324, 314, _, _, _, 67, 299, 
    _, _, 356, 170, 0, 348, 330, 321, 36, _, 45, 357, 323, 334, 15, 338, 38, 
    234, 178, 204, 187, 350, 225, 116, 8, 216, 248, 258, 22, 319, 315, 49, 
    66, 93, 14, 0, _, 328, 89, 41, 356, 96, 310, 9, 25, 18, 355, 0, 302, 345, 
    63, 123, 1, 301, 297, 304, 260, 231, 354, 238, 358, 124, 303, 352, 104, 
    0, 3, 216, 0, 357, 226, 329, 26, 324, 335, 323, 323, 354, 347, 356, 326, 
    0, 358, 323, 0, 32, 1, 135, 53, _, 311, 44, 81, 98, 87, 70, 105, 121, 2, 
    156, 318, 255, 125, 91, 359, 16, 313, 348, _, 266, 336, 320, 114, 161, 
    219, 212, 212, 55, 299, 7, 38, 66, 51, 42, 305, 140, 313, 270, 209, 333, 
    33, 266, 123, 15, 187, 56, 217, 325, 292, 1, _, 99, 322, 261, 173, 262, 
    244, 278, 271, 267, 92, 13, 345, 292, 341, 323, 55, 327, 317, 335, 74, 
    220, 282, 333, 114, 4, 322, 122, 0, 159, 343, 5, 279, 88, 4, 323, _, 324, 
    97, 82, _, 90, 105, 99, 91, 103, 107, 104, 110, 107, 101, 100, 81, 114, 
    122, 111, 101, _, 114, 95, 320, 308, 325, 303, 83, 324, 347, 301, 284, 
    72, 7, 331, 341, 340, 303, 353, 266, 295, 354, 10, 161, 289, 329, 358, 
    353, 297, 303, 0, 351, 357, 356, 9, 310, 93, 80, 0, 358, 131, 358, 236, 
    271, 270, 271, 268, 264, 287, 114, 246, 56, 294, 300, 276, _, 300, _, 
    270, 270, 276, 263, 270, 308, 288, 249, 330, 238, 137, 240, 239, 295, 
    339, 233, 6, 355, 325, 346, 311, 335, 0, 6, _, 326, 3, 90, 62, 118, 163, 
    75, 297, 99, 51, 54, 63, 61, 26, 50, 49, 21, 280, 251, 336, 43, 47, 48, 
    352, 359, 298, 355, 59, 249, 244, 264, 292, 271, 271, 272, 281, 268, 286, 
    255, 286, 266, 352, 5, 332, 321, 285, 333, 299, 301, 280, 290, 287, 272, 
    273, 245, 281, 110, 112, 122, 131, 100, 105, 114, 120, 100, _, 91, 96, 
    336, 320, 343, 316, 293, 306, 294, 274, 278, 10, 281, 176, 149, 114, 98, 
    114, 357, 162, 304, 320, 325, 323, 297, 305, 328, 329, 329, 312, 8, 306, 
    267, 360, 0, _, 279, 270, 277, 284, 270, 287, 286, 45, 359, 71, 325, 352, 
    0, 326, 281, 79, 84, 304, 304, 207, 291, 313, 275, 285, 290, 280, 281, 
    273, 121, 94, 16, 134, 137, 360, 319, _, 318, 14, 5, 338, 1, 267, 300, 
    248, _, _, _, 251, 2, 176, 145, 98, 66, 65, 72, 68, 66, 78, 69, _, 66, 
    29, 26, 339, 30, 312, 33, 0, 348, 35, 332, 268, 262, 263, 262, 210, 349, 
    256, 270, 263, 269, 253, 56, 353, 358, 89, 329, 303, 86, 99, 0, 313, 281, 
    108, 348, 268, 250, 296, 136, 131, 164, 123, 149, 152, 77, 141, 107, _, 
    93, 83, 87, 144, 129, 118, 100, 119, 128, 107, 138, 132, 101, 121, 151, 
    171, 30, 137, 128, 124, 169, 128, 75, _, 168, 132, 113, 139, 277, 136, 
    137, 105, 101, 117, 113, 92, 130, 121, 152, 164, 126, 131, 133, 122, 131, 
    125, 98, 94, 84, 26, 19, 98, 23, 2, 299, 305, 299, 316, 115, 129, 117, 
    124, 38, 139, 186, 219, 201, 208, 79, 327, 88, _, 84, 130, 122, 70, 116, 
    0, 89, 261, 270, 22, 275, 292, 54, 347, 41, 208, 88, 98, 98, 92, 87, 84, 
    90, _, 85, 81, 60, 71, 61, 67, 304, 293, 124, 106, 117, 130, 298, 310, 
    351, 265, 267, 173, 81, 189, 279, 241, 323, 18, 67, 83, 49, 53, 7, 353, 
    15, 102, 305, 245, 257, 173, 125, 284, 287, 269, 260, 274, 137, 276, 214, 
    269, 278, _, 295, 313, 304, 299, 307, 120, 184, 70, 86, 298, 300, 294, 
    56, 114, 293, 273, 320, 128, 124, 131, 125, _, 120, _, 273, 324, 330, 
    303, 351, 343, 356, 85, 135, 128, 139, 67, 325, 348, 313, 269, 277, 267, 
    272, 165, 19, 169, 209, 218, 187, 238, 202, 206, 250, 236, 259, 163, 349, 
    223, 229, 247, 290, 40, 46, 44, 46, 42, 50, 49, 66, 43, 113, _, 83, 82, 
    95, 90, 84, 103, 109, 142, 0, 243, 76, 28, 334, 73, 20, 141, 251, 272, 
    264, 265, 292, _, 359, _, _, 136, 101, 1, 112, 87, 327, 120, 108, 0, 273, 
    137, 177, 320, 0, 356, 358, 167, 360, 331, 3, 32, 39, 23, 31, 24, 40, 48, 
    47, 39, 46, 47, 48, 51, 54, 53, 52, 50, 60, 63, 55, 57, 59, 61, 49, 53, 
    47, _, 304, 303, 295, 296, 74, 327, 339, 245, 356, 0, 358, 152, 183, 230, 
    249, _, 233, 287, 164, 147, _, _, 265, _, 308, 19, 22, 60, 0, 1, 61, 108, 
    14, 92, 151, 260, 155, 164, 147, 159, 254, 257, 270, 269, 269, 344, 150, 
    116, 175, 349, 227, 345, 90, 148, 280, 276, 300, 254, 258, 272, 267, 263, 
    179, 164, 139, 243, 255, 239, 151, 340, 321, _, 14, 60, 99, 211, 299, 
    269, 243, 269, 273, 271, 280, 285, _, 256, 270, 269, 208, 166, 164, 311, 
    167, _, 175, 168, 127, 28, 53, 355, 291, 294, 27, 0, 242, 278, 280, 301, 
    303, _, _, 346, 52, 0, 128, 38, 112, 0, 0, 294, 74, 19, 93, 67, 303, 342, 
    0, 310, 135, 339, 278, 336, 114, 298, 267, 333, 149, 345, 163, 128, 126, 
    303, 358, _, 358, 360, 0, _, 131, 111, 130, 124, 162, 134, 141, _, 254, 
    232, 252, 201, 158, 270, 269, 268, 285, _, 272, 273, 7, 0, 321, 93, 0, 
    90, 355, 267, 135, 149, 235, 137, 128, 265, 168, 164, 234, 149, 139, _, 
    161, 293, 247, 114, 276, 335, 333, 128, 354, 299, 10, 9, 292, 284, 290, 
    294, 211, 260, 119, 147, 30, 280, 8, 112, 70, 198, 300, _, 124, 143, 320, 
    305, 302, 314, 317, 306, 303, 272, 265, 285, 287, 272, 275, 279, 282, 
    274, 290, 288, 281, _, _, _, 310, 26, 8, 1, 306, 294, 230, 124, 302, 306, 
    314, 320, 310, 304, 294, 295, 290, 306, _, _, 272, _, 262, 302, 295, 296, 
    308, 296, 293, 282, 273, 271, 292, 304, 121, 166, 173, 197, 284, 286, 
    296, 295, 174, 162, 171, 158, 151, 92, 84, 88, 115, 93, 111, 1, 288, 277, 
    274, 275, 272, 269, 291, 51, 49, 72, 51, 93, 76, 271, 109, _, 283, 62, 
    357, 305, 274, 297, 285, 287, 268, 272, 264, 260, 264, 269, 267, 263, 
    248, 244, 250, _, 263, _, 261, _, 256, 254, 274, 274, 279, 253, 270, 276, 
    290, 268, 275, 300, 295, 273, 290, 286, 102, 295, _, 198, 43, 42, 15, 20, 
    129, 79, 57, 38, 46, _, 47, 67, 33, 88, 158, 137, 124, 156, 167, 153, 
    109, 112, 97, 68, 68, 58, 58, 46, 63, 53, 62, 257, 54, 3, 240, 49, 72, 
    331, 229, 69, 65, 158, 159, 127, 149, 163, 152, 184, 182, _, 257, _, 269, 
    266, 276, 279, 284, 284, 273, 277, 269, 278, 267, 275, 301, 131, 114, _, 
    98, 66, 119, 96, 59, 63, 38, 41, 10, 60, 45, 247, 54, 54, 178, 65, 340, 
    296, 304, 312, 288, 293, 274, 280, 295, 270, 270, 268, 270, 268, 266, 
    270, 288, 286, 284, 275, 271, 277, 275, 272, 273, 266, 271, 286, 290, 
    288, 298, 306, 312, 304, 296, 294, 291, 285, 267, _, 281, 277, 280, 286, 
    290, 301, 312, 200, 157, 339, 334, 51, 52, 29, 48, _, 57, 42, 57, 40, 44, 
    26, 29, 61, 53, 18, _, 86, 69, 197, 270, 292, 254, 313, 303, 295, 303, 
    296, 268, 282, 288, 275, 270, 281, 301, 301, 294, 276, 287, 293, 296, 
    301, 295, 290, 289, 286, 285, 295, 297, 294, 288, 273, 278, 273, 267, 
    269, 259, 260, 266, 265, 280, _, 272, 284, 293, 295, 295, 291, 286, 292, 
    302, 267, 287, 301, 91, 96, 78, 101, 262, 295, 93, 110, 127, 293, 315, 
    303, 310, 292, 295, 288, 297, 302, 286, 176, 20, 184, 59, 124, 6, 48, 94, 
    77, 270, 314, 300, 317, 309, 107, 90, 116, 288, 279, _, 269, 243, 76, 
    250, 249, 107, 64, 14, 353, 293, 121, 124, 144, 128, 132, 122, 118, 123, 
    133, 134, _, 287, 300, 288, 277, 60, 290, 88, 40, 105, 147, 96, 109, 90, 
    127, 128, 122, 130, 130, 142, 126, 146, 111, 125, 115, 119, 136, 4, 125, 
    349, 291, 249, 298, 289, 255, 36, 285, 154, 114, 126, 135, 132, 105, 110, 
    94, 109, 96, 113, 167, 102, 85, 98, 60, 327, 276, 31, 137, 142, 229, 203, 
    166, 297, 147, 167, 173, 173, 187, 231, 274, 269, 265, 272, _, 277, 282, 
    281, 284, 294, 277, 279, 272, 271, 271, 274, 293, 288, 287, 299, 279, 
    269, 268, 174, 176, 169, 158, _, _, _, _, _, 124, 116, 138, 137, _, 85, 
    168, 11, 294, 292, 285, 258, 180, 175, 168, 159, 160, 162, 161, 178, 181, 
    172, 182, _, 295, 292, 294, 228, 171, 291, 291, 280, 289, 290, 291, 181, 
    172, 118, 126, 105, 0, 125, 144, _, 289, _, 320, 331, 337, 358, 180, 220, 
    293, 291, 287, 280, 293, 292, 275, 281, 267, 287, 290, 285, 296, 295, 
    295, 302, 290, 309, 318, 326, 304, 296, 302, 195, 301, 281, 301, 250, 
    312, 297, 297, 290, 271, 190, _, 152, 160, 115, 152, 131, 164, 75, 335, 
    116, 294, 86, 349, 74, 5, 106, 113, 5, 28, 137, 169, 120, 126, 136, 134, 
    133, 123, 120, 95, 295, 305, 122, 121, 2, 122, 183, 55, 155, 286, 296, 
    153, 141, 290, 13, 136, 113, 168, 155, 58, 82, 107, _, 123, 269, 285, 
    291, 291, 305, 278, _, 277, 309, 0, 120, 354, 290, 113, 265, 293, 352, 5, 
    20, 43, 20, 131, 122, 122, 354, 295, 272, 258, 108, 76, 313, 294, 315, 
    310, 9, 0, 120, 287, 261, 122, 303, 272, 294, 125, 111, 351, 115, 121, 
    130, 116, 319, 123, 146, 0, 24, 7, 78, 81, 328, 134, 9, 74, 32, 139, 175, 
    163, 148, 107, 78, 94, _, 85, 95, 107, 118, 106, 124, 301, 309, 349, 108, 
    95, 104, 317, 308, 249, 134, 332, 262, 109, 128, 117, _, 108, _, 109, 71, 
    110, 89, 93, 116, 122, 127, 105, 127, 115, 103, 122, 117, 125, 125, 109, 
    107, 100, 101, 150, 180, 162, 99, 129, 110, 100, 302, 275, 340, 288, 10, 
    59, 10, 134, 309, 66, 322, 127, 0, 30, 95, 115, 109, 187, 298, 139, _, 
    14, 39, 331, 300, 330, 167, 322, 118, 0, 346, 0, 15, 61, 122, 154, 83, 
    186, 290, 82, 105, 153, 205, 99, _, 341, 61, 17, 318, 238, 282, 317, 269, 
    63, 136, 105, 246, 244, 343, 196, 185, 274, 137, 127, 121, 131, 125, 140, 
    124, 123, 142, 102, 136, 133, 141, 144, 113, 132, 145, 181, 225, 332, 40, 
    9, 173, _, 318, 144, 151, 120, 161, 266, _, 265, 263, 271, 277, 267, 262, 
    271, 278, 279, 289, 290, 285, 293, 291, 190, 53, 47, 213, 250, 54, 78, 
    64, 84, 73, 291, 21, 42, 33, 41, 15, 194, 15, 14, 2, 15, 21, 53, 257, 71, 
    78, 326, 219, 341, 56, 88, 55, 33, 234, 60, 66, 199, 56, 183, 329, 309, 
    302, 32, 0, 344, 0, 286, 182, 263, 293, 85, 63, 71, 62, 80, 71, 76, _, 
    159, 180, 71, 207, 279, 0, 335, 332, 330, 8, 15, 351, 346, 219, 5, 117, 
    124, 121, 81, 64, _, 76, 105, _, 70, 73, 130, 295, 134, 201, 293, 326, 
    326, 256, 297, 359, 30, 335, 75, 65, 66, 57, 91, 59, 60, 42, 70, _, 91, 
    88, 138, 123, 78, 118, 94, 94, 54, 63, 69, 347, 3, 43, 88, 243, 0, 89, 
    335, 151, 57, 34, 170, _, 75, 110, 69, 84, 66, 259, 25, 43, 40, 35, 19, 
    53, 105, 113, 103, 111, 57, 68, 40, 79, _, _, 146, _, 61, 93, 55, 41, 60, 
    191, 65, 76, _, 295, 252, 120, 129, 115, 95, 93, 96, 165, 159, 155, 129, 
    130, 129, 146, 135, 146, 149, 134, 129, 89, 0, 24, 0, 316, 10, 0, 107, 
    82, 110, _, 104, 133, 132, 138, 143, 133, 145, _, 145, 124, 97, 119, 122, 
    96, 111, 64, 87, 125, 105, 78, 206, 141, 125, 133, 164, 184, 142, 107, _, 
    _, 109, _, 100, 93, 99, 124, 117, 128, 113, 85, 117, 131, 113, 71, 71, 
    112, 104, 48, 114, 123, 102, 105, 123, 85, 102, 118, 116, 114, 100, 123, 
    112, 137, _, 109, 109, 115, 102, 123, 199, 7, 177, 212, 269, 293, 307, 
    267, 246, 263, 273, _, 286, 274, 295, 289, 293, 290, 288, 294, 313, 296, 
    297, 308, 295, 295, 292, 262, 271, 267, 271, 272, 276, _, 294, _, 274, 
    279, 294, 299, 272, _, 289, 300, 300, 318, 278, 306, 338, _, _, 302, 195, 
    175, 199, 173, 167, _, 169, 164, 126, 146, 161, 155, 80, 90, 247, 81, 89, 
    122, 92, 80, 126, 131, 128, 134, 159, 148, 159, 177, 144, 357, 172, _, 
    105, 104, 130, 132, 134, 113, 122, 36, 0, 315, 359, _, 354, 70, 181, 238, 
    273, 264, 265, 266, 285, _, 279, _, 246, 177, 175, 153, 172, 172, 175, 
    180, 182, 70, 325, 318, 300, 297, 297, 130, 147, 112, 175, 155, 135, 136, 
    147, 171, 336, 166, 181, 132, 99, 54, 202, 301, 284, 295, 254, 256, 303, 
    302, 247, 276, 262, 189, 169, 145, 110, 112, 130, 145, 175, 166, 293, 
    280, 262, 264, 265, 269, 288, 258, 273, 273, 298, 271, 283, 278, 183, 
    180, 117, 128, 169, 160, 150, 140, 133, 132, 0, 359, 144, 0, 123, 115, 5, 
    56, 123, 155, 315, 98, 283, 277, 282, 175, 168, 170, 172, 165, 102, 89, 
    119, 306, 62, 74, 93, 108, 96, 53, 107, 102, 27, 0, 280, 112, 119, 317, 
    280, 15, 166, 260, 132, 126, 122, 110, 132, 169, 157, 342, 10, 306, 307, 
    302, 110, 195, 155, 74, 223, 34, 358, 137, 88, 115, 2, 124, 347, _, _, 
    111, 126, 162, 142, 131, 314, 104, 142, 120, 123, 85, 170, 164, 165, 78, 
    3, 14, 2, 129, 110, _, 213, 271, 229, 355, 108, 293, 264, 320, 350, 327, 
    320, 312, 277, 5, 100, 130, 128, 340, 138, 359, 4, 0, 109, 135, 0, 114, 
    120, 169, 167, 156, 26, 0, 138, 152, 88, 88, 111, 121, 315, 295, 215, 
    237, 222, 251, 195, 226, 102, 130, 153, 123, 108, 128, 102, 106, 111, 
    112, 109, 129, 102, 117, 143, 279, 114, 296, 134, 111, 96, 130, 140, 87, 
    120, 133, 123, 121, 108, 124, 128, 114, 102, 123, 332, 237, 170, 70, 61, 
    40, 51, 193, 185, 46, 66, 197, 220, 230, 111, 82, 71, 66, 83, 99, 116, 
    130, 104, 353, 94, 97, 262, 305, 306, 285, 288, 292, 276, 128, 126, 76, 
    356, 159, 139, 159, 157, 149, 125, 130, 132, 160, 136, 145, 144, 6, 358, 
    335, 355, 83, 27, 49, 335, 280, 0, 274, 351, 0, 299, 287, 329, _, 99, 
    105, 113, 3, 0, 88, 102, 106, 95, 314, 317, 14, 9, 355, 285, _, 279, 158, 
    111, 51, 170, 191, 186, 206, 315, 174, 47, 98, 304, 254, 328, 340, 353, 
    354, 0, 232, 232, 334, 146, 303, 280, 118, 67, 102, 75, 59, 71, 55, 220, 
    _, 157, 72, 157, 122, 98, 87, 303, 283, 283, 274, _, 271, 271, 268, 279, 
    286, 279, 275, 306, 303, 269, _, 268, 105, 51, 22, 171, 72, 240, 28, 68, 
    3, 61, 2, 80, 335, 0, 289, 314, 271, 269, 265, 242, 265, 272, 270, 267, 
    288, 265, 264, 255, 264, 276, 298, 276, 328, 318, 315, 330, 315, 324, 
    319, 314, 305, 105, 144, 91, 164, 144, 143, 70, _, 349, 129, 144, 118, 
    108, 358, 303, 310, 315, 314, 334, _, 275, 265, 284, 278, 260, 332, 1, 6, 
    _, _, 154, 248, 141, 74, 53, 48, 43, 86, 288, 60, 276, 261, 295, 281, 
    259, 257, 249, 311, 75, 119, 99, 211, 278, 355, 299, 293, 302, 302, 310, 
    213, 202, 297, 303, 288, 291, 296, 301, 311, 304, 302, 312, 334, 109, 88, 
    120, 338, 296, 334, 0, 105, 276, 277, 275, 329, 3, 313, 50, 8, 357, 0, 
    86, 312, 347, 95, 116, 331, 136, 5, 342, 356, 5, _, 33, 89, 1, 113, 100, 
    123, 0, 77, 107, 286, 25, 0, 86, 48, 300, 122, 354, 118, 120, 357, 278, 
    18, 40, 134, 138, 312, 80, 156, 80, 123, 109, 126, 118, 123, 5, 80, 69, 
    80, 93, 73, 69, 93, 84, 83, 94, 90, 87, 98, 83, 96, _, 81, 81, 302, 312, 
    357, 340, 61, 84, 68, 7, 329, 105, 351, 320, 46, 122, 263, 122, 100, 263, 
    _, 61, 129, 238, 231, 268, 353, 117, 159, 41, 9, _, 358, 34, 314, 130, _, 
    _, 315, 129, 123, 121, 73, 128, 101, 77, 78, 322, 265, 293, 285, 303, 
    301, 317, 305, 330, 332, 302, 93, 0, 310, 315, 59, 9, _, 98, 212, 125, 
    124, 72, 82, _, 145, 303, 130, 324, 357, 357, 337, 317, 349, 329, 22, 
    317, 21, 143, 103, 99, 119, 137, 110, 111, _, 113, 124, 97, 124, 112, 
    114, 129, 119, 104, 103, 326, 241, 94, 83, 357, 292, 301, 295, 209, 154, 
    _, 128, 74, 96, 92, 80, 55, 34, 289, 267, _, _, 290, 15, 109, 352, 22, 
    337, 36, 73, 139, 358, 133, 104, 108, 137, 145, 137, 115, 132, 109, 126, 
    112, 359, 85, 114, 134, 139, 121, 139, 107, 84, 94, 85, 102, 95, 92, 113, 
    122, 135, 161, 170, 162, 127, 113, 128, 304, 280, 7, 103, 341, 15, 97, 
    83, 83, 343, 113, 101, 312, 43, 339, 293, _, 314, 300, 109, 45, 83, 94, 
    94, 93, 92, 89, 70, 88, 84, 87, 88, 100, 108, 116, 110, 92, 94, _, 100, 
    105, 101, 106, 105, 97, 94, 98, 97, 94, 95, 71, 86, 69, 80, 74, 77, 74, 
    84, 76, 101, 353, 316, 109, 73, 78, 74, 76, 91, 80, 93, 92, 76, 90, 93, 
    74, 89, 91, 105, 44, 49, 37, 31, 355, 52, 84, 82, 61, 247, _, 304, 112, 
    16, _, 8, 23, 12, 80, 90, 48, 75, 333, 339, 15, 330, 345, 192, 154, 236, 
    126, 79, 55, 189, 67, 142, 56, 102, 87, 59, 64, 81, 287, 329, 26, 50, 56, 
    61, 60, 76, 49, 44, 36, 61, 71, 58, 81, 39, 57, 60, 96, 349, 76, _, 54, 
    46, 56, 37, 87, 0, 82, 353, 2, _, 71, _, _, _, 288, 359, 0, _, _, 169, 
    156, 167, 168, 185, 179, 181, 173, 140, 160, 127, 114, 108, 106, 343, 
    319, 319, 315, 304, 350, 290, 321, 156, 144, 140, 171, 169, 153, 91, 144, 
    153, 178, 79, 201, 328, 6, 38, 48, 318, 314, 284, 340, 2, 5, 264, 274, 
    266, 259, 113, 169, 176, 159, 296, 302, 287, 322, 323, 26, 356, 352, 82, 
    50, 60, 62, 317, 308, 306, 330, 346, 355, 275, _, 159, 126, 111, 105, 91, 
    87, 88, 91, 208, 234, 67, 290, 221, 337, _, 175, 321, 230, 225, 274, 306, 
    315, 313, 314, _, 233, 259, 288, 300, 312, 314, 297, 315, 316, 331, 318, 
    322, 299, 310, 296, 298, 307, 303, 276, 251, 252, 252, 262, 255, 274, 
    270, _, 256, 265, 298, 295, 296, 286, 288, 268, 259, 280, 280, 288, 276, 
    295, 294, 288, 278, 267, 275, _, 276, 278, 270, 276, 291, 282, 317, 308, 
    10, 59, 108, 326, 325, 285, 306, 296, 295, 354, 6, 98, 303, _, 101, _, 
    111, 31, 274, 295, 314, 303, 313, 317, 311, 315, 315, 295, 322, 324, 312, 
    322, 334, 335, 0, 356, 1, _, 13, 7, 127, 197, 130, 84, 47, 40, 46, 32, 2, 
    15, 33, 24, 354, 17, 10, _, 219, 353, 348, 13, 139, 305, 70, _, 77, 63, 
    87, 93, 99, 98, 109, 112, 119, 79, 87, 325, 264, 306, 290, 283, 313, 293, 
    285, 329, 309, _, 76, _, 278, 297, 283, 271, 272, 282, 287, 284, 268, 
    349, 301, 295, 82, 21, 237, 283, 18, _, 356, 282, 258, 288, 77, 96, 10, 
    198, 237, 267, 278, 268, 298, _, 287, 313, 335, 333, 32, 360, 336, 191, 
    332, 86, 89, 74, 78, 99, 116, _, 114, 82, 86, 101, 90, 78, 79, 89, 82, 
    76, 62, 307, 303, 336, 301, 29, 312, 304, 302, 319, 306, _, 316, _, 297, 
    306, 319, 303, 290, 314, 161, 317, 19, 340, 329, 320, 325, 325, _, 346, 
    316, 328, 348, 41, 41, 356, 345, 158, 99, 227, 318, 138, 360, 352, 322, 
    359, 19, 360, 326, 0, 0, 49, 326, 331, 1, 30, 0, 357, 346, 109, 356, _, 
    88, 1, 353, _, 82, 326, 300, 7, 52, 349, 9, 4, 48, 45, 24, _, 316, 81, 
    296, 338, 59, _, 334, _, 121, 0, 357, 0, 303, 120, _, 348, 105, 80, 125, 
    330, 297, 33, _, 1, 315, 68, 287, _, 29, _, 0, 0, 43, 355, 347, 360, 338, 
    320, 10, 314, 321, 7, 95, 92, 354, 92, 328, 335, 106, 358, 355, 349, 353, 
    32, 326, _, 133, 261, 271, 107, 287, 355, 352, 1, 53, 48, 33, 109, 353, 
    65, 109, 347, 8, 342, 358, 312, 314, _, _, 340, 343, 51, 29, 338, 83, 
    113, 73, 70, 66, 72, 77, 74, 71, 311, 294, 299, 311, 312, 96, 15, 331, 
    341, 94, _, 80, 87, 64, 57, 83, 81, 101, 112, 115, 94, 104, 110, 100, 91, 
    79, _, 109, 97, 105, 104, 116, 86, 107, 99, 105, 96, 35, 44, 106, 116, 
    106, 96, 310, 317, 102, 135, 0, 309, 350, 329, 106, 92, 59, 47, 332, _, 
    _, 276, 299, 275, 10, 305, 300, 313, 314, 11, 75, 56, 353, 313, 25, 0, 9, 
    0, 335, 356, 323, _, 353, 358, 340, 0, 313, 205, 4, 359, 113, 101, 96, 
    98, 104, 336, 309, 354, 301, 0, 349, _, 335, 339, 0, 358, 330, 341, 322, 
    338, 283, 195, 250, 181, 266, 337, _, 288, 342, 290, 278, 341, 357, 341, 
    7, 313, 0, 0, 0, 0, 0, 0, 331, 272, 354, 291, 351, 327, 308, 296, 332, 
    307, 311, 342, 357, 0, 333, 25, 0, 45, 316, 308, 22, 45, 311, _, 317, 
    355, 306, 301, 1, 323, 313, 313, 324, 78, 3, 49, 86, 339, 307, 100, 332, 
    _, 357, 357, 77, 9, 310, 301, 356, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 315, 322, 122, 315, 341, 64, 30, 
    96, 87, 47, 51, _, 30, 314, 305, 349, 0, 89, 7, 340, _, 15, 318, 4, 54, 
    _, 47, 57, 284, 284, 71, 288, 312, 23, 332, 57, 76, 8, 312, 302, 309, 
    314, 318, 310, 254, 99, 99, 89, 301, 307, 300, _, 320, _, 322, 304, 294, 
    293, 299, 311, 319, 313, 317, 316, 310, 323, 193, 197, 175, 181, _, 83, 
    129, 143, 0, 287, 302, 296, 296, 278, 291, 279, 310, 294, 295, 297, 302, 
    309, 312, 307, 305, 291, _, 292, 288, 302, 296, 312, 297, 290, 318, 307, 
    308, 305, 337, 338, 294, 320, 344, 31, 304, 329, 42, 325, 298, 313, 323, 
    317, 309, 301, 296, 294, 13, 318, 305, 320, 339, 358, 67, 336, 135, 307, 
    158, 45, 19, 21, 46, 20, 10, 26, 27, 263, 221, 221, 212, 323, 260, 318, 
    277, 318, 314, 320, 36, 15, 60, 77, 71, 63, 51, 54, 78, 70, 72, 94, _, 
    97, 95, 98, 93, 90, 91, 105, 100, 95, 87, _, 101, 102, 105, 102, 82, 89, 
    101, 104, 95, 93, 98, 94, 94, 85, 94, 99, 97, 105, _, 103, 102, 89, 100, 
    84, 88, 86, 70, 71, 112, 80, 104, 67, 18, 35, 84, 114, 99, 207, 11, 28, 
    350, 76, 78, 76, 67, 75, 85, 73, 59, 58, 52, 50, 60, 72, 67, 60, 70, 60, 
    69, 39, 337, 316, 286, 322, 295, 293, 328, 253, 347, 77, 87, 73, 70, 64, 
    71, 108, 88, 79, 89, _, 323, 324, 309, 296, 8, 342, 331, 30, _, _, 346, 
    9, 340, _, 206, 53, 317, 328, 292, 324, 79, 30, 109, 235, 34, 50, 74, 11, 
    36, 48, 46, _, 315, 326, 304, 303, 312, 305, 332, 324, 328, 332, 315, 
    299, 313, 328, 305, 308, 317, 313, 322, 310, _, 308, 317, 259, 335, 340, 
    344, 325, 316, 310, 33, 269, 320, 328, 281, 64, 301, 281, 327, 319, 307, 
    307, 62, 318, 312, 305, 333, 333, 316, 295, 61, 310, 48, 338, 338, 317, 
    351, 310, 338, 326, 312, 30, 313, 311, 302, 316, 59, 326, 107, 98, 102, 
    _, 94, 98, 102, 98, 103, 106, 90, 93, 83, 100, 66, 64, 66, 58, 33, 60, 
    62, 34, 49, 7, _, 39, 323, 49, 339, 335, 321, 306, 297, 324, 324, 329, 
    327, 315, 351, 1, 342, 315, 352, 299, 324, 337, 316, 357, 304, 289, 298, 
    307, 342, 332, 329, 316, 327, 328, 322, 338, 309, 312, 315, 316, 316, 
    331, 333, 33, 27, 24, 22, 43, 46, 66, 58, _, 30, 136, 45, 55, 62, 16, 3, 
    6, 360, 352, 350, 348, 9, 1, 359, 358, 4, 352, 4, 17, 28, 16, 11, 17, 
    114, 19, 206, 10, 10, 18, 269, 257, 293, 105, 339, 5, 24, 354, 339, 9, 
    357, _, 303, 313, 312, 352, 326, 339, 315, 300, 312, 314, 296, 315, 321, 
    19, 352, 70, 48, 60, 93, 54, 77, 107, 202, 294, 275, 296, 285, 346, 353, 
    _, 323, 307, 317, 331, 285, 323, 296, 340, 332, 308, 302, 304, 328, 294, 
    324, 310, 313, 312, 352, 353, 306, 317, 53, 316, 326, 306, 315, 324, 306, 
    341, 349, 57, 343, 26, 330, 1, 297, 329, 317, 308, 321, _, 346, 344, 359, 
    322, 314, 1, 315, 313, 324, 333, 332, 9, 294, 304, 323, 326, 311, 349, 
    340, 355, 344, 305, 334, 53, 53, 45, 31, 17, 293, 1, 33, 79, 246, 340, 
    327, 329, 311, 285, 15, 295, 317, 315, 6, 318, 324, 6, 310, 307, 55, 24, 
    306, 310, 304, 318, 311, 344, 339, 323, 281, 308, 317, 321, 307, 309, 
    285, 294, 304, 336, 308, 309, 342, _, 336, 336, 322, 326, 318, 327, 327, 
    2, _, _, _, 323, 294, 310, 302, 316, 318, 170, 314, 324, 301, 344, 317, 
    312, 328, 337, 300, 308, 336, 285, 302, 319, 341, 304, 315, 313, 325, 
    296, 311, 320, 294, 301, 358, 321, 303, 322, 336, 318, 319, 325, 321, 
    346, _, 358, 319, 292, 315, 303, 280, 353, 296, 304, 314, 339, 320, 349, 
    322, 0, 333, 327, 58, _, 15, 330, 0, 2, 329, 346, 350, 354, 56, 33, 51, 
    18, 334, 18, 7, 14, 1, 23, 12, 27, 41, 50, 43, 59, 48, 52, 97, 104, 80, 
    110, 97, 92, 88, 87, 94, 99, 102, _, _, 96, 65, 57, 221, 334, 308, 329, 
    266, 276, 317, 301, 303, 321, 318, 336, 322, 67, 315, 345, 307, 312, 311, 
    316, 314, 310, 299, 306, 343, 333, 298, 331, 339, 337, 335, 341, 353, 
    320, 342, 354, 48, 291, 350, 3, 314, 359, 313, 312, 359, 320, 320, 308, 
    357, 313, 337, 338, 338, 310, 301, 315, 315, 315, 297, 299, 325, 296, 
    296, 315, 286, 304, 77, 98, 86, 91, 96, 93, 68, 75, 295, 290, 284, 277, 
    288, 298, 304, 125, 77, 40, 60, 73, 51, 320, 212, 57, 300, 213, 228, 360, 
    3, 6, 253, 250, 242, 271, 318, 310, 308, 304, 303, 314, 323, 317, 321, 
    315, 321, 323, 313, 323, 306, 292, 306, 90, 301, 330, 335, 2, 8, 360, 
    259, 320, 301, 314, 320, 317, 326, 37, 55, 84, 83, 98, 104, 96, 110, 118, 
    110, 110, 103, 89, 95, 95, 92, 97, 99, 92, 96, 96, 67, 176, 312, 324, 
    304, 312, 313, 296, 305, 318, 304, 231, 298, 295, 270, 261, 308, 271, 
    271, 293, 281, 291, 274, 283, 243, 280, 282, 274, 292, 282, 281, 282, 
    315, 294, 318, 323, 283, 305, 298, 291, 292, 285, 298, 295, 292, 296, 
    295, 269, 301, 317, 288, 319, 97, 36, 352, 320, 291, 303, 320, 296, 262, 
    269, 77, 279, 20, 332, 305, 306, 307, 276, 296, 327, 309, 305, 313, 314, 
    305, 62, 311, 328, 11, 330, 318, 324, 326, 325, 325, _, _, _, _, _, 294, 
    295, 296, 305, 310, 286, 313, 298, 306, 311, 318, 2, 292, 304, 306, 311, 
    310, 317, 306, 354, 328, 327, 308, 300, 283, 331, 322, 332, 289, 14, 0, 
    301, 338, 317, 298, 312, 309, 305, 4, 343, 305, 329, 108, 340, 131, 360, 
    345, 360, 13, 34, 44, 45, 359, 113, 44, 215, 38, 43, 201, 42, 294, 309, 
    281, 293, 278, 316, 271, 291, 319, 300, 303, 315, 317, 314, 313, 299, 1, 
    350, 327, 324, 298, 353, 353, 332, 338, 324, 332, 309, 359, 8, 309, 312, 
    293, 287, 314, 267, 45, 4, 29, 318, 19, 203, 4, 3, 15, 32, 272, 63, 280, 
    315, 318, 313, 307, 317, 335, 1, 350, 41, 322, 290, 329, 314, 316, 309, 
    310, 305, 332, 296, 279, 293, 299, 283, 299, 325, 354, 325, 30, 0, 307, 
    310, 326, 317, 319, 320, 323, 68, 59, 73, 83, 60, 49, 60, 77, 85, 16, 0, 
    341, 337, 356, 359, 26, 35, 32, 31, 30, 29, 25, 29, 31, 35, 34, 32, 34, 
    32, 32, 34, 38, 31, 26, 27, 27, 33, 39, 46, 35, 44, 29, 27, 26, 312, 292, 
    247, 304, 312, 335, 297, 338, 303, 301, 289, 309, 316, 310, 297, 351, 
    342, 325, 287, 310, 307, 305, 316, 291, 295, 299, 300, 313, 309, 334, 
    253, 320, 337, 319, 301, 323, 343, 4, 342, 336, 346, 305, 306, 307, 321, 
    313, 326, 299, 302, 275, 297, 310, 314, 345, 319, 320, 271, 22, 354, 10, 
    6, 360, 3, 26, 357, 3, 35, 30, 33, 22, 28, 36, 17, 36, 17, 32, 2, 4, 77, 
    328, 2, 1, 274, 322, 311, 310, 310, 323, 315, 315, 303, 313, 306, 333, 
    313, 317, 330, 350, 314, 308, 300, 25, 359, 334, 327, 330, 16, 327, 297, 
    304, 313, 24, 311, 320, 309, 305, 314, 321, 306, 331, 313, 307, 326, 300, 
    65, 178, 40, 110, 119, 94, 94, 89, 89, 88, 81, 74, 72, 73, 73, 88, 91, 
    93, 91, 90, 92, 90, 76, 56, 66, 70, 52, 257, 70, 310, 216, 172, 78, 86, 
    81, 70, 65, 39, 85, 329, 322, 310, 305, 289, 15, 353, 359, 172, 291, 251, 
    102, 215, 73, 70, 22, 323, 330, 340, 350, 352, 150, 182, 112, 293, 35, 4, 
    42, 40, 42, 42, 40, 40, 38, 42, 40, 41, 41, 37, 23, 34, 35, 37, 27, 1, 
    308, 317, 336, 292, 289, 269, 9, 310, 329, 280, 321, 311, 307, 313, 318, 
    313, 312, 344, 298, 295, 283, 299, 296, 273, 295, 331, 263, 294, 316, 
    314, 309, 311, 326, 275, 312, 340, 285, 320, 22, 327, 272, 352, 26, 332, 
    19, 1, 88, 337, 324, 6, 312, 232, 263, 282, 292, 261, 345, 187, 336, 328, 
    295, 341, 334, 330, 313, 315, 300, 337, 334, 55, 325, 320, 296, 321, 317, 
    257, 307, 316, 302, 326, 290, 352, 337, 317, 292, 316, 311, 316, 328, 
    337, 318, 305, 315, 303, 317, 343, 352, 333, 18, 15, 320, 331, 14, 310, 
    13, 355, 320, 331, 328, 330, 317, 290, 300, 318, 314, 291, 273, 277, 321, 
    52, 22, 5, 14, 10, 7, 15, 12, 279, 9, 1, 26, 346, 266, 287, 288, 305, 
    283, 314, 297, 320, 313, 307, 276, 228, 331, 18, 338, 296, 286, 322, 307, 
    288, 293, 307, 304, 338, 251, 333, 78, 18, 333, 315, 309, 319, 284, 329, 
    324, 320, 331, 37, 321, 326, 324, 346, 355, 345, 338, 1, 339, 329, 335, 
    317, 343, 321, 301, 313, 282, 339, 351, 308, 298, 319, 335, 317, 311, 
    339, 353, 288, 250, 349, 26, 37, 30, 49, 38, 40, 39, 32, 35, 39, 47, 2, 
    190, 333, 358, 39, 5, 65, 31, 30, 30, 41, 58, 195, 127, 59, 19, 340, 269, 
    295, 288, 173, 58, 27, 31, 20, 235, 339, 4, 5, 154, 258, 7, 6, 341, 10, 
    29, 177, 300, 173, 38, 17, 130, 136, 103, 297, 320, 358, 320, 27, 9, 43, 
    24, 54, 53, 50, 45, 40, 30, 188, 266, 208, 286, 290, 317, 343, 279, 290, 
    310, 214, 315, 312, 262, 294, 309, 323, 296, 299, 271, 303, 334, 339, 
    357, 325, 8, 12, 288, 165, 332, 173, 266, 287, 105, 10, 334, 326, 317, 
    339, 322, 326, 323, 297, 302, 315, 318, 326, 302, 350, 319, 320, 322, 
    335, 334, 252, 30, 316, 322, 77, 303, 315, 317, 357, 346, 337, 340, 326, 
    19, 359, 2, 8, 336, 327, 28, 325, 319, 348, 7, 342, 2, 341, 12, 10, 54, 
    333, 18, 46, 298, 23, 338, 297, 295, 334, 353, 73, 79, 94, 82, 90, 100, 
    80, 79, 60, 73, 60, 23, 31, 29, 33, 56, 15, 27, 156, 48, 53, 71, 9, 13, 
    7, 30, 5, 341, 345, 347, 6, 11, 13, 19, 18, 17, 23, 19, 18, 25, 360, 360, 
    3, 6, 26, 12, 14, 12, 5, 25, 24, 21, 37, 341, 134, 100, 39, 340, 360, 20, 
    346, 360, 17, 0, 356, 306, 280, 316, 307, 308, 329, 304, 276, 301, 302, 
    307, 3, 310, 83, 86, 329, 60, 26, 300, 294, 294, 301, 304, 309, 296, 298, 
    299, 328, 320, 295, 294, 300, 292, 301, 311, 315, 89, 38, 353, 304, 329, 
    10, 327, 314, 313, 324, 312, 310, 311, 336, 335, 327, 299, 6, 343, 84, 
    88, 82, 93, 91, 39, 107, 90, 59, 49, 30, 18, 42, 10, 83, 96, 135, 100, 
    123, 63, 69, 63, 74, 74, 74, 66, 67, 79, 69, 66, 113, 85, 47, 357, 75, 
    73, 51, 86, 92, 93, 88, 16, 329, 297, 302, 290, 280, 265, 250, 233, 262, 
    270, 269, 273, 275, 298, 313, 314, 299, 303, 285, 300, 342, 317, 316, 
    353, 349, 2, 334, 297, 18, 336, 75, 1, 29, 346, 352, 297, 294, 308, 327, 
    317, 310, 305, 304, 335, 307, 321, 357, 101, 358, 345, 340, 288, 65, 316, 
    356, 342, 329, 60, 46, 316, 52, 3, 72, 360, 303, 13, 91, 22, 255, 1, 28, 
    313, 359, 339, 328, 292, 314, 318, 328, 325, 303, 313, 341, 310, 318, 
    301, 303, 309, 286, 304, 299, 304, 36, 319, 81, 289, 297, 304, 345, 311, 
    304, 319, 318, 303, 120, 304, 77, 316, 301, 305, 307, 316, 310, 307, 78, 
    75, 74, 67, 92, 72, 85, 86, 95, 122, 117, 84, 88, 68, 78, 76, 105, 77, 
    74, 94, 85, 96, 85, 85, 94, 87, 93, 98, 109, 95, 90, 89, 91, 84, 78, 81, 
    92, 78, 87, 81, 81, 59, 51, 58, 57, 75, 76, 54, 95, 83, 81, 87, 55, 107, 
    94, 71, 81, 89, 91, 71, 89, 102, 94, 92, 94, 85, 105, 95, 101, 86, 67, 
    94, 96, 78, 92, 90, 95, 88, 79, 83, 82, 80, 87, 85, 82, 92, 86, 88, 86, 
    91, 90, 91, 94, 95, 92, 72, 91, 80, 65, 73, 57, 55, 61, 57, 58, 58, 58, 
    51, 45, 47, 63, 44, 85, 83, 74, 94, 120, 97, 79, 74, 73, 51, 310, 77, 67, 
    58, 76, 77, 80, 86, 80, 79, 78, 89, 81, 84, 76, 303, 313, 296, 198, 69, 
    90, 91, 95, 93, 98, 79, 73, 75, 75, 85, 86, 74, 85, 96, 97, 97, 109, 108, 
    84, 70, 76, 67, 84, 292, 304, 299, 315, 325, 347, 299, 292, 335, 306, 
    312, 314, 309, 313, 333, 300, 347, 336, 336, 338, 359, 0, 301, 317, 41, 
    300, 299, 316, 359, 353, 328, 48, 338, 5, 345, 356, 7, 292, 342, 332, 
    302, 359, 18, 338, 0, 12, 11, 349, 324, 48, 301, 302, 303, 16, 321, 8, 
    342, 48, 354, 347, 335, 316, 0, 339, 351, 308, 311, 290, 353, 47, 312, 
    117, 9, 319, 132, 96, 310, 315, 319, 2, 346, 19, 206, 345, 311, 301, 291, 
    307, 301, 304, 304, 296, 260, 299, 307, 331, 296, 301, 315, 0, 314, 330, 
    310, 308, 321, 331, 343, 110, 68, 328, 37, 320, 313, 310, 325, 71, 324, 
    315, 328, 345, 327, 50, 42, 331, 359, 312, 357, 70, 332, 50, 360, 9, 259, 
    321, 339, 309, 5, 95, 67, 68, 70, 72, 72, 67, 82, 69, 70, 85, 101, 100, 
    98, 96, 97, 93, 91, 100, 115, 125, 91, 91, 79, 72, 73, 285, 292, 108, 
    295, 316, 354, 314, 339, 309, 325, 33, 305, 64, 311, 218, 73, 89, 40, 
    285, 293, 320, 286, 306, 312, 323, 310, 308, 312, 304, 290, 308, 321, 
    299, 352, 316, 316, 306, 29, 7, 337, 356, 36, 354, 2, 350, 328, 0, 338, 
    348, 327, 313, 354, 357, 45, 348, 23, 58, 317, 317, 65, 356, 3, 357, 83, 
    331, 314, 3, 334, 352, 360, 360, 328, 6, 358, 0, 27, 359, 347, 343, 27, 
    298, 8, 331, 77, 88, 1, 332, 335, 74, 316, 328, 351, 353, 85, 1, 68, 355, 
    346, 287, 350, 300, 97, 305, 334, 329, 120, 0, 351, 313, 357, 355, 23, 
    339, 1, 106, 92, 307, 248, 222, 218, 247, 305, 247, 214, 273, 298, 286, 
    308, 91, 70, 3, 306, 359, 294, 304, 309, 320, 331, 349, 357, 0, 337, 310, 
    296, 309, 320, 360, 22, 313, 314, 288, 350, 100, 360, 352, 360, 2, 10, 
    30, 38, 360, 360, 0, 304, 297, 311, 305, 360, 90, 306, 337, 355, 17, 115, 
    297, 9, 12, 356, 360, 347, 330, 313, 329, 43, 358, 356, 352, 30, 333, 64, 
    30, 13, 350, 34, 96, 350, 324, 37, 29, 39, 357, 348, 358, 15, 344, 35, 
    321, 107, 311, 4, 308, 311, 312, 309, 360, 50, 4, 52, 306, 357, 339, 353, 
    348, 99, 325, 341, 348, 35, 74, 342, 313, 65, 350, 1, 327, 304, 72, 92, 
    348, 336, 289, 313, 0, 359, 354, 360, 73, 23, 316, 331, 88, 327, 301, 
    319, 26, 0, 360, 18, 26, 330, 66, 305, 350, 232, 6, 360, 237, 234, 221, 
    244, 309, 290, 287, 289, 262, 243, 267, 235, 258, 221, 232, 207, 193, 
    169, 198, 191, 220, 273, 277, 268, 273, 262, 291, 290, 287, 278, 322, 
    302, 306, 315, 328, 284, 301, 312, 310, 312, 286, 311, 313, 304, 244, 
    269, 259, 282, 272, 263, 279, 254, 258, 248, 262, 259, 264, 292, 294, 
    309, 296, 301, 312, 311, 7, 13, 322, 325, 335, 346, 316, 321, 341, 309, 
    26, 335, 5, 334, 63, 316, 32, 22, 24, 25, 88, 33, 182, 318, 51, 297, 331, 
    317, 351, 295, 112, 351, 5, 301, 0, 315, 48, 0, 316, 340, 21, 328, 3, 84, 
    38, 0, 0, 0, 0, 0, 360, 37, 305, 298, 303, 304, 263, 290, 311, 326, 336, 
    324, 308, 304, 319, 345, 340, 304, 325, 330, 326, 14, 71, 17, 325, 99, 
    319, 309, 5, 310, 32, 353, 284, 360, 75, 306, 313, 339, 357, 68, 352, 59, 
    99, 344, 344, 0, 0, 0, 0, 0, 290, 299, 298, 321, 324, 292, 299, 187, 99, 
    288, 88, 124, 300, 327, 47, 334, 86, 94, 335, 314, 92, 313, 326, 320, 
    318, 6, 329, 300, 324, 106, 302, 1, 359, 65, 350, 1, 315, 307, 317, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 341, 0, 0, 325, 91, 83, 86, 89, 86, 74, 328, 80, 80, 87, 89, 54, 
    308, 6, 331, 60, 309, 69, 17, 68, 323, 351, 299, 304, 71, 89, 118, 101, 
    300, 316, 335, 321, 12, 328, 296, 19, 17, 327, 15, 20, 19, 327, 349, 319, 
    72, 9, 315, 62, 297, 332, 298, 314, 293, 318, 311, 314, 309, 350, 65, 
    329, 325, 1, 296, 301, 296, 347, 67, 349, 318, 313, 12, 285, 299, 301, 
    345, 327, 303, 329, 294, 300, 310, 320, 335, 277, 303, 17, 28, 360, 305, 
    312, 2, 56, 73, 316, 70, 351, 82, 29, 56, 336, 306, 309, 315, 315, 106, 
    23, 7, 1, 113, 76, 327, 313, 319, 320, 326, 1, 325, 83, 68, 349, 321, 19, 
    353, 321, 343, 64, 2, 27, 97, 58, 309, 97, 113, 97, 69, 297, 314, 319, 
    315, 320, 100, 32, 336, 348, 5, 66, 24, 5, 38, 358, 0, 0, 360, 66, 359, 
    8, 27, 48, 319, 360, 15, 35, 64, 9, 313, 15, 326, 318, 50, 106, 16, 74, 
    360, 304, 71, 325, 87, 66, 76, 82, 77, 83, 68, 68, 274, 295, 78, 82, 90, 
    95, 94, 84, 93, 80, 99, 88, 80, 98, 97, 94, 86, 92, 92, 93, 93, 86, 79, 
    85, 77, 309, 63, 315, 11, 35, 5, 359, 111, 350, 2, 287, 74, 5, 324, 316, 
    113, 307, 59, 9, 354, 57, 299, 322, 342, 301, 25, 293, 100, 73, 85, 35, 
    16, 28, 318, 341, 360, 81, 89, 354, 351, 331, 357, 322, 350, 331, 52, 59, 
    351, 77, 22, 323, 99, 350, 350, 351, 352, 331, 334, 52, 84, 84, 80, 64, 
    77, 72, 79, 78, 73, 73, 75, 79, 75, 92, 94, 95, 77, 71, 119, 72, 100, 
    234, 70, 74, 92, 87, 100, 97, 81, 93, 101, 86, 83, 90, 93, 86, 93, 86, 
    72, 74, 321, 248, 89, 96, 88, 80, 77, 75, 70, 66, 94, 78, 314, 87, 64, 
    87, 74, 75, 65, 78, 88, 114, 89, 95, 94, 94, 84, 105, 98, 87, 73, 92, 
    103, 107, 103, 66, 92, 62, 100, 292, 340, 329, 356, 130, 68, 83, 87, 96, 
    101, 116, 96, 95, 82, 85, 75, 54, 86, 106, 96, 94, 88, 116, 80, 144, 93, 
    303, 76, 108, 90, 341, 319, 97, 100, 288, 22, 318, 9, 315, 308, 315, 360, 
    18, 52, 98, 348, 348, 353, 312, 322, 42, 38, 324, 298, 308, 18, 326, 325, 
    56, 128, 75, 40, 95, 65, 57, 78, 166, 107, 143, 90, 105, 43, 38, 81, 67, 
    100, 177, 150, 124, 154, 93, 98, 96, 92, 99, 97, 84, 78, 130, 99, 84, 80, 
    84, 91, 91, 76, 80, 86, 81, 75, 91, 83, 81, 87, 77, 78, 97, 95, 98, 93, 
    90, 86, 82, 80, 76, 78, 99, 97, 111, 76, 81, 93, 94, 95, 81, 82, 88, 87, 
    91, 91, 80, 95, 64, 58, 74, 82, 81, 93, 80, 86, 85, 105, 88, 83, 58, 89, 
    100, _, 102, 80, 59, 314, 308, 87, 71, 77, 68, 65, 83, 67, 46, 49, 301, 
    334, 338, 330, 343, 355, 107, 121, 12, 27, 2, 315, 284, 296, 260, 88, 4, 
    47, 14, 45, 360, 20, 45, 44, 53, 70, 50, 338, 11, 317, 353, 60, 71, 75, 
    65, 83, 85, 81, 98, 103, 85, 79, 79, 86, 78, 85, 83, 80, 90, 87, 83, 88, 
    88, 88, 77, 78, 85, 87, 76, 80, 87, 84, 69, 65, 94, 64, 48, 39, 27, 73, 
    274, 58, 354, 90, 329, 320, 27, 356, 350, 342, 354, 81, 360, 304, 52, 
    360, 304, 310, 329, 328, 36, 360, 320, 296, 298, 310, 320, 339, 111, 180, 
    306, 312, 299, 297, 290, 292, 289, 275, 270, 289, 291, 284, 270, 292, 
    300, 300, 303, 295, 294, 312, 300, 325, 313, 298, 296, 281, 305, 290, 
    297, 307, 318, 307, 300, 307, 314, 306, 310, 318, 328, 312, 315, 2, 342, 
    70, 3, 350, 4, 15, 325, 296, 355, 311, 65, 314, 330, 316, 273, 69, 324, 
    321, 49, 316, 320, 302, 6, 299, 50, 315, 351, 305, 323, 321, 327, 317, 
    299, 323, 162, 316, 63, 39, 67, 50, 39, 330, 32, 42, 25, 27, 42, 38, 48, 
    60, 39, 50, 69, 44, 64, 58, 71, 50, 52, 55, 57, 58, 59, 80, 48, 50, 65, 
    44, 65, 65, 64, 61, 60, 77, 85, 62, 41, 41, 42, 48, 37, 49, 57, 75, 75, 
    69, 67, 35, 251, 354, 328, 26, 359, 342, 344, 0, 326, 37, 353, 354, 23, 
    32, 29, 337, 334, 18, 295, 307, 297, 288, 285, 290, 296, 291, 311, 37, 
    64, 269, 20, 38, 57, 294, 334, 323, 23, 287, 289, 270, 289, 296, 312, 
    289, 278, 335, 5, 354, 6, 358, 321, 322, 341, 0, 303, 76, 359, 308, 343, 
    54, 162, 289, 131, 336, 306, 299, 296, 360, 97, 194, 85, 317, 336, 1, 
    359, 12, 272, 227, 193, 284, 298, 322, 312, 293, 330, 36, 249, 300, 315, 
    315, 336, 347, 330, 341, 332, 330, 328, 290, 328, 331, 322, 261, 120, 
    312, 316, 356, 8, 48, 0, 328, 340, 331, 6, 0, 17, 360, 288, 322, 316, 
    331, 323, 314, 316, 4, 331, 313, 326, 263, 352, 78, 71, 51, 67, 356, 43, 
    244, 297, 281, 325, 307, 330, 321, _, _, _, _, _, _, 36, 32, 35, 32, 19, 
    304, 5, 328, 350, 83, 12, 16, 338, 328, 293, 341, 327, 310, 312, 28, 15, 
    89, 333, 354, 72, 299, 314, 308, 307, 293, 296, 20, 33, 32, 19, 313, 309, 
    307, 308, 320, 332, 13, 13, 303, 89, 329, 300, 317, 79, 17, 307, 317, 11, 
    7, 318, 107, 72, 263, 83, 104, 93, 92, 92, 73, 72, 82, 70, 77, 76, 68, 
    87, 99, 98, 101, 97, 91, 105, 293, 6, 330, 30, 63, 18, 123, 77, 99, 88, 
    86, 78, 73, 92, 92, 91, 80, 78, 92, 105, 103, 79, 88, 100, 113, 79, 78, 
    81, 77, 136, 128, 65, 114, 47, 60, 323, 319, 316, 112, 22, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 70, 83, 68, 78, 106, 82, 90, 92, 101, 68, 
    84, 75, 93, 95, 76, 80, 79, 79, 271, 287, 111, 91, 65, 72, 77, 318, 290, 
    302, 300, 11, 10, 358, 343, 356, 356, 322, 336, 35, 325, 15, 337, 305, 
    252, 0, 359, 300, 305, 313, 347, 1, 0, 348, 360, 22, 8, 25, 328, 5, 33, 
    356, 63, 95, 71, 28, 30, 42, 346, 188, 42, 7, 12, 26, 32, 40, 164, 129, 
    306, 277, 336, 319, 305, 343, 19, 330, 6, 340, 326, 319, 0, 321, 57, 313, 
    334, 37, 7, 3, 79, 309, 317, 23, 322, 44, 59, 305, 11, 335, 323, 60, 318, 
    36, 301, 352, 39, 355, 3, 9, 9, 24, 360, 339, 340, 356, 8, 59, 3, 309, 
    32, 61, 64, 349, 2, 334, 360, 56, 12, 197, 100, 73, 3, 329, 344, 317, 
    319, 269, 308, 326, 307, 270, 314, 314, 55, 360, 348, 352, 345, 326, 26, 
    34, 336, 358, 343, 333, 352, 357, 10, 1, 348, 59, 313, 337, 10, 356, 84, 
    3, 74, 302, 284, 291, 299, 20, 323, 320, 24, 229, 187, 311, 234, 74, 164, 
    49, 155, 302, 223, 358, 253, 267, 228, 253, 279, 258, 346, 271, 316, 312, 
    35, 94, 117, 95, 161, 264, 260, 115, 265, 328, 325, 164, 135, 338, 310, 
    305, 301, 283, 289, 285, 233, 35, 351, 335, 50, 201, 96, 9, 277, 13, 283, 
    334, 302, 305, 343, 316, 305, 296, 317, 300, 320, 334, 4, 34, 346, 314, 
    41, 1, 8, 351, 70, 352, 321, 343, 101, 322, 333, 89, 309, 98, 293, 328, 
    25, 311, 64, 337, 323, 318, 0, 356, 58, 349, 304, 338, 340, 26, 327, 343, 
    5, 353, 321, 289, 58, 343, 357, 84, 1, 340, 43, 357, 356, 322, 12, 326, 
    317, 346, 308, 308, 305, 322, 9, 317, 355, 313, 54, 44, 4, 1, 310, 312, 
    73, 43, 335, 87, 77, 356, 319, 359, 359, 319, 345, 27, 331, 51, 18, 349, 
    328, 2, 96, 1, 26, 320, 322, 315, 312, 319, 320, 307, 320, 3, 330, 19, 
    346, 52, 2, 352, 33, 50, 60, 18, 328, 341, 12, 38, 297, 360, 11, 346, 26, 
    352, 347, 312, 0, 1, 10, 343, 321, 2, 99, 360, 4, 324, 348, 100, 309, 99, 
    83, 301, 290, 299, 352, 338, 310, 315, 316, 316, 205, 13, 30, 22, 16, 
    119, 64, 343, 55, 319, 312, 300, 269, 90, 309, 110, 10, 330, 333, 318, 
    330, 325, 318, 12, 6, 338, 342, 29, 12, 323, 354, 58, 321, 57, 308, 34, 
    319, 72, 317, 57, 309, 320, 355, 320, 308, 110, 20, 287, 125, 348, 99, 
    354, 18, 4, 360, 109, 61, 0, 358, 99, 322, 355, 300, 270, 276, 279, 278, 
    277, 277, 284, 283, 283, 268, 300, 297, 295, 47, 40, 42, 135, 51, 223, 
    20, 38, 98, 281, 88, 172, 139, 80, 58, 88, 50, 212, 176, 89, 56, 55, 57, 
    12, 254, 49, 341, 303, 339, 13, 312, 329, 15, 250, 348, 287, 269, 210, 
    32, 117, 312, 288, 293, 285, 336, 311, 321, 331, 291, 283, 348, 318, 310, 
    278, 282, 317, 321, 314, 56, 312, 136, 20, 100, 169, 107, 117, 35, 247, 
    338, 336, 325, 53, 36, 39, 56, 5, 341, 297, 285, 348, 335, 311, 296, 316, 
    339, 326, 343, 308, 16, 12, 220, 265, 326, 12, 228, 230, 230, 185, 104, 
    58, 10, 199, 320, 120, 181, 151, 73, 132, 51, 169, 16, 103, 260, 294, 
    291, 295, 324, 210, 209, 289, 324, 347, 340, 334, 285, 331, 329, 87, 20, 
    30, 34, 96, 8, 10, 6, 41, 19, 337, 294, 304, 0, 360, 11, 53, 345, 350, 
    325, 330, 351, 321, 84, 339, 27, 348, 0, 68, 297, 311, 65, 0, 317, 90, 0, 
    47, 259, 53, 217, 19, 46, 275, 347, 69, 340, 58, 290, 270, 7, 350, 331, 
    323, 32, 5, 0, 6, 336, 305, 284, 97, 8, 295, 339, 233, 28, 22, 360, 350, 
    278, 280, 19, 288, 357, 147, 160, 338, 262, 109, 177, 123, 28, 236, 285, 
    296, 319, 291, 192, 211, 339, 318, 277, 33, 301, 335, 313, 16, 340, 270, 
    261, 337, 320, 321, 303, 72, 360, 325, 95, 288, 77, 353, 39, 344, 312, 
    17, 315, 19, 19, 355, 336, 52, 18, 324, 91, 4, 325, 297, 0, 287, 114, 
    335, 0, 114, 0, 336, 290, 305, 16, 0, 34, 69, 25, 359, 271, 79, 327, 0, 
    307, 274, 13, 310, 13, 0, 46, 110, 2, 348, 349, 294, 308, 65, 45, 314, 
    310, 293, 340, 314, 335, 329, 44, 62, 31, 72, 66, 72, 70, 73, 52, 52, 48, 
    34, 16, 45, 35, 17, 33, 47, 349, 164, 217, 80, 21, 40, 1, 359, 307, 283, 
    302, 297, 300, 289, 6, 352, 353, 40, 46, 26, 40, 33, 38, 38, 39, 46, 44, 
    28, 356, 40, 346, 359, 342, 9, 341, 326, 230, 359, 25, 19, 70, 349, 26, 
    35, 173, 353, 354, 337, 9, 330, 19, 66, 322, 52, 318, 21, 11, 312, 63, 
    310, 352, 324, 330, 288, 95, 0, 304, 354, 87, 347, 319, 90, 0, 356, 344, 
    341, 327, 317, 350, 338, 314, 359, 27, 329, 73, 66, 346, 106, 0, 351, 0, 
    0, 132, 357, 65, 334, 84, 39, 339, 304, 325, 323, 303, 49, 333, 336, 320, 
    280, 312, 288, 310, 62, 306, 287, 118, 299, 286, 325, 95, 36, 3, 36, 4, 
    307, 309, 316, 40, 306, 359, 309, 284, 87, 90, 100, 83, 84, 81, 73, 53, 
    46, 38, 55, 86, 207, 156, 22, 34, 33, 13, 17, 34, 28, 36, 25, 354, 340, 
    43, 32, 88, 74, 51, 40, 3, 37, 72, 56, 37, 89, 57, 64, 35, 50, 83, 339, 
    359, 12, 295, 314, 0, 338, 300, 290, 285, 278, 297, 281, 306, 279, 345, 
    275, 270, 54, 338, 318, 12, 71, 307, 327, 0, 315, 339, 343, 355, 243, 
    260, 267, 292, 249, 293, 291, 283, 334, 80, 89, 320, 340, 334, 332, 332, 
    338, 355, 307, 3, 77, 324, 354, 47, 2, 359, 351, 301, 331, 293, 214, 343, 
    332, 291, 284, 19, 14, 55, 301, 76, 293, 117, 84, 332, 313, 314, 360, 14, 
    325, 33, 282, 150, 139, 10, 255, 194, 271, 340, 350, 4, 59, 359, 47, 31, 
    35, 49, 35, 7, 70, 61, 197, 45, 53, 26, 282, 232, 172, 202, 292, 56, 245, 
    270, 268, 309, 326, 41, 348, 338, 56, 46, 317, 73, 12, 321, 303, 307, 58, 
    137, 358, 313, 282, 290, 284, 15, 328, 277, 292, 102, 348, 74, 50, 314, 
    32, 326, 326, 306, 305, 296, 1, 328, 243, 308, 348, 360, 89, 168, 84, 92, 
    97, 295, 312, 74, 183, 319, 85, 315, 324, 328, 351, 347, 28, 329, 332, 
    75, 0, 0, 0, 268, 263, 183, 258, 51, 350, 8, 299, 341, 329, 172, 90, 120, 
    49, 83, 315, 100, 97, 4, 335, 351, 319, 291, 290, 286, 283, 330, 10, 100, 
    120, 130, 360, 5, 210, 350, 43, 355, 30, 356, 340, 346, 28, 317, 318, 
    330, 58, 71, 78, 48, 51, 63, 43, 45, 282, 257, 290, 358, 288, 71, 73, 
    338, 11, 332, 352, 334, 298, 299, 91, 109, 100, 91, 71, 106, 80, 135, 
    100, 151, 146, 285, 284, 32, 53, 315, 16, 81, 319, 8, 305, 316, 345, 300, 
    276, 293, 112, 90, 43, 52, 139, 328, 339, 186, 101, 127, 52, 344, 1, 316, 
    257, 317, 357, 93, 296, 73, 182, 6, 350, 225, 359, 51, 84, 1, 351, 51, 
    168, 79, 175, 225, 349, 351, 71, 56, 9, 324, 289, 280, 319, 39, 56, 36, 
    78, 107, 86, 94, 88, 98, 111, 108, 124, 126, 119, 123, 93, 51, 40, 42, 
    38, 34, 23, 113, 68, 60, 52, 248, 7, 338, 305, 310, 261, 273, 280, 275, 
    280, 270, 259, 265, 292, 251, 319, 353, 346, 293, 8, 318, 356, 5, 338, 
    329, 350, 318, 355, 320, 305, 263, 222, 183, 147, 250, 258, 267, 267, 15, 
    30, 34, 0, 0, 319, 79, 328, 0, 341, 10, 0, 0, 0, 342, 134, 0, 157, 360, 
    7, 255, 248, 264, 266, 44, 325, 74, 19, 325, 294, 76, 93, 303, 102, 326, 
    304, 143, 329, 359, 136, 303, 312, 261, 143, 281, 139, 107, 100, 343, 2, 
    105, 96, 278, 294, 315, 323, 294, 316, 324, 302, 69, 101, 102, 106, 95, 
    93, 84, 305, 316, 324, 318, 322, 311, 293, 304, 321, 319, 314, 327, 320, 
    302, 310, 299, 301, 296, 311, 296, 300, 297, 266, 296, 289, 293, 276, 
    287, 289, 283, 277, 277, 270, 275, 284, 282, 277, 276, 275, 288, 286, 
    276, 280, 287, 86, 142, 182, 193, 213, 284, 0, 266, 253, 310, 248, 77, 
    70, 267, 325, 265, 0, 289, 305, 25, 13, 126, 0, 272, 282, 275, 344, 1, 
    239, 0, 0, 70, 242, 189, 257, 41, 329, 5, 359, 337, 331, 329, 318, 3, 12, 
    39, 18, 36, 30, 338, 29, 23, 44, 64, 61, 61, 8, 25, 33, 27, 37, 39, 37, 
    39, 18, 28, 26, 38, 45, 54, 53, 64, 61, 59, 55, 45, 242, 55, 54, 60, 54, 
    41, 39, 37, 300, 312, 319, 352, 293, 82, 0, 306, 288, 277, 273, 271, 272, 
    266, 274, 258, 246, 70, 206, 185, 95, 54, 29, 11, 37, 40, 356, 256, 12, 
    6, 10, 291, 260, 164, 276, 217, 219, 226, 57, 57, 63, 51, 45, 45, 359, 3, 
    24, 32, 37, 50, 60, 55, 47, 42, 38, 37, 38, 40, 47, 52, 46, 47, 40, 39, 
    59, 69, 59, 38, 35, 30, 37, 50, 41, 1, 2, 332, 354, 339, 357, 302, 295, 
    300, 262, 155, 157, 246, 268, 271, 276, 271, 264, 287, 271, 261, 279, 
    279, 310, 346, 322, 128, 50, 274, 296, 300, 350, 221, 270, 281, 258, 275, 
    272, 277, 274, 285, 278, 281, 299, 298, 3, 104, 154, 91, 274, 283, 290, 
    270, 256, 225, 280, 273, 283, 282, 271, 285, 292, 290, 297, 292, 337, 
    289, 226, 77, 213, 62, 194, 324, 36, 43, 50, 27, 21, 41, 39, 35, 278, 
    255, 265, 221, 257, 263, 261, 276, 232, 250, 268, 97, 289, 344, 105, 328, 
    21, 107, 359, 274, 88, 250, 277, 277, 172, 272, 274, 266, 162, 271, 269, 
    268, 282, 270, 125, 100, 33, 40, 51, 0, 305, 18, 0, 342, 7, 31, 1, 199, 
    223, 198, 274, 173, 180, 184, 223, 252, 117, 136, 164, 241, 288, 346, 
    352, 312, 315, 119, 287, 301, 57, 304, 310, 324, 289, 296, 291, 288, 301, 
    303, 292, 286, 292, 288, 294, 265, 201, 289, 167, 3, 267, 319, 357, 70, 
    0, 321, 267, 235, 287, 268, 265, 228, 258, 227, 179, 195, 301, 230, 254, 
    117, 133, 313, 89, 349, 325, 356, 0, 297, 336, 88, 355, 298, 285, 288, 
    278, 10, 123, 143, 0, 0, 259, 273, 251, 262, 3, 0, 350, 0, 348, 4, 308, 
    293, 325, 0, 358, 312, 290, 264, 265, 265, 265, 273, 53, 60, 41, 58, 54, 
    62, 239, 50, 346, 173, 358, 335, 18, 28, 14, 13, 270, 2, 354, 269, 267, 
    154, 175, 156, 223, 238, 184, 182, 0, 280, 282, 89, 70, 318, 350, 108, 
    296, 0, 0, 346, 349, 143, 314, 274, 270, 267, 179, 269, 260, 267, 277, 
    222, 0, 153, 304, 288, 345, 324, 329, 289, 311, 298, 308, 299, 257, 286, 
    269, 254, 263, 266, 260, 256, 251, 260, 265, 260, 263, 269, 272, 278, 
    274, 282, 289, 299, 298, 299, 291, 279, 285, 290, 296, 301, 281, 300, 
    277, 286, 284, 304, 297, 296, 316, 326, 44, 96, 114, 298, 0, 0, 287, 0, 
    46, 96, 61, 47, 273, 301, 309, 281, 299, 314, 293, 291, 296, 298, 320, 
    286, 295, 322, 311, 273, 301, 316, 322, 319, 312, 309, 304, 297, 298, 
    307, 332, 269, 61, 26, 3, 134, 335, 357, 0, 342, 0, 35, 333, 311, 325, 0, 
    308, 352, 58, 140, 3, 9, 256, 184, 149, 100, 69, 111, 303, 147, 120, 194, 
    154, 204, 195, 187, 198, 243, 348, 287, 169, 129, 201, 51, 92, 109, 107, 
    106, 108, 39, 99, 130, 174, 203, 170, 170, 183, 147, 145, 140, 122, 129, 
    112, 299, 251, 304, 262, 212, 168, 18, 260, 268, 294, 273, 5, 302, 271, 
    275, 282, 268, 268, 282, 293, 292, 302, 300, 319, 323, 298, 299, 310, 
    286, 309, 201, 102, 100, 89, 64, 70, 92, 95, 82, 111, 218, 55, 58, 246, 
    66, 59, 264, 263, 112, 342, 20, 241, 171, 20, 17, 172, 133, 124, 122, 
    132, 132, 128, 122, 137, 140, 271, 270, 271, 277, 275, 66, 80, 7, 27, 
    109, 133, 0, 53, 43, 137, 167, 286, 148, 136, 137, 121, 159, 263, 130, 
    133, 168, 268, 305, 159, 0, 323, 89, 348, 0, 12, 0, 186, 249, 265, 137, 
    120, 137, 166, 259, 163, 157, 172, 95, 145, 117, 123, 279, 159, 342, 299, 
    297, 301, 335, 314, 315, 296, 304, 302, 298, 281, 141, 164, 119, 149, 
    201, 283, 211, 140, 132, 277, 291, 303, 279, 263, 356, 322, 310, 318, 
    294, 304, 306, 302, 313, 299, 298, 290, 296, 316, 285, 282, 288, 287, 
    266, 278, 283, 296, 322, 318, 324, 302, 308, 297, 144, 137, 111, 128, 
    152, 173, 232, 196, 179, 175, 221, 197, 206, 176, 191, 138, 275, 133, 
    308, 349, 0, 10, 261, 110, 160, 173, 157, 161, 137, 143, 157, 281, 292, 
    167, 118, 137, 127, 110, 72, 87, 120, 64, 276, 0, 0, 163, 135, 79, 300, 
    275, 316, 288, 297, 285, 187, 175, 181, 179, 195, 311, 173, 182, 163, 15, 
    300, 314, 308, 124, 331, 136, 66, 141, 116, 163, 87, 60, 59, 53, 81, 122, 
    111, 102, 94, 89, 92, 74, 96, 67, 76, 178, 49, 324, 128, 0, 310, 14, 123, 
    127, 127, 119, 137, 268, 257, 270, 268, 273, 272, 273, 281, 277, 283, 
    276, 283, 281, 292, 291, 288, 279, 272, 289, 238, 360, 6, 33, 311, 286, 
    264, 296, 307, 47, 40, 339, 237, 280, 297, 293, 290, 318, 42, 49, 39, 54, 
    55, 56, 66, 85, 84, 55, 315, 26, 119, 76, 116, 284, 13, 360, 304, 328, 
    152, 35, 12, 151, 355, 77, 245, 44, 338, 37, 65, 140, 147, 136, 137, 132, 
    130, 126, 128, 150, 274, 282, 292, 292, 309, 280, 302, 286, 179, 76, 118, 
    132, 102, 87, 93, 250, 273, 274, 218, 133, 178, 87, 65, 125, 111, 108, 
    99, 115, 99, 95, 100, 107, 113, 118, 112, 116, 110, 108, 117, 106, 114, 
    124, 131, 132, 103, 52, 54, 62, 32, 175, 9, 46, 24, 28, 48, 95, 323, 345, 
    48, 38, 33, 59, 96, 76, 329, 61, 50, 55, 60, 84, 352, 38, 41, 54, 71, 79, 
    78, 94, 45, 28, 52, 67, 51, 41, 54, 37, 65, 125, 122, 111, 106, 280, 118, 
    52, 69, 42, 201, 106, 58, 58, 54, 52, 65, 53, 54, 59, 51, 54, 53, 327, 
    71, 52, 51, 252, 227, 128, 110, 128, 160, 148, 167, 165, 167, 160, 158, 
    159, 160, 134, 113, 106, 91, 78, 152, 152, 147, 127, 129, 156, 164, 152, 
    157, 161, 165, 165, 165, 163, 165, 160, 170, 121, 112, 111, 129, 143, 
    120, 121, 110, 147, 102, 98, 92, 105, 124, 118, 112, 78, 81, 77, 140, 
    133, 135, 137, 267, 259, 334, 332, 236, 288, 292, 290, 278, 275, 264, 
    267, 245, 294, 270, 160, 155, 165, 326, 68, 264, 175, 356, 270, 286, 285, 
    289, 304, 279, 287, 297, 273, 175, 10, 129, 115, 114, 155, 168, 171, 150, 
    204, 288, 282, 286, 296, 273, 291, 313, 296, 0, 336, 307, 298, 274, 286, 
    293, 304, 324, 300, 271, 142, 168, 137, 204, 177, 279, 252, 293, 268, 
    280, 305, 296, 301, 339, 293, 209, 200, 152, 314, 233, 339, 159, 127, 
    130, 126, 134, 159, 131, 114, 127, 128, 126, 126, 107, 134, 167, 138, 
    108, 105, 114, 93, 297, 291, 274, 239, 120, 122, 147, 99, 126, 117, 102, 
    111, 113, 132, 127, 182, 190, 158, 139, 135, 150, 2, 0, 287, 70, 146, 
    316, 15, 28, 120, 135, 26, 157, 135, 149, 120, 79, 108, 109, 110, 105, 
    100, 111, 106, 108, 111, 100, 77, 87, 69, 59, 236, 95, 89, 83, 90, 114, 
    139, 108, 128, 126, 58, 53, 282, 112, 109, 98, 157, 150, 179, 163, 86, 
    179, 118, 123, 92, 103, 120, 117, 104, 114, 127, 259, 325, 177, 170, 183, 
    238, 241, 265, 272, 269, 270, 271, 258, 280, 205, 15, 164, 138, 126, 92, 
    119, 173, 119, 126, 123, 132, 134, 123, 128, 127, 132, 127, 128, 131, 
    119, 117, 107, 95, 97, 109, 284, 290, 266, 290, 292, 263, 103, 124, 127, 
    122, 155, 150, 127, 339, 176, 24, 167, 171, 17, 89, 86, 127, 20, 0, 314, 
    306, 299, 290, 268, 149, 119, 227, 166, 112, 108, 167, 179, 169, 186, 
    198, 178, 137, 169, 142, 156, 183, 252, 240, 235, 176, 190, 171, 170, 
    179, 234, 128, 133, 133, 131, 117, 125, 114, 131, 132, 142, 147, 141, 
    128, 305, 292, 295, 286, 292, 292, 281, 288, 294, 169, 160, 175, 174, 
    177, 175, 175, 175, 178, 174, 293, 207, 178, 162, 181, 124, 88, 104, 117, 
    124, 125, 151, 120, 127, 119, 112, 131, 131, 131, 135, 136, 142, 130, 
    120, 113, 65, 176, 103, 107, 336, 323, 62, 352, 326, 10, 0, 208, 93, 117, 
    100, 145, 132, 144, 135, 114, 131, 120, 98, 118, 270, 280, 165, 141, 109, 
    156, 165, 161, 159, 161, 117, 141, 141, 136, 141, 150, 164, 145, 161, 
    121, 154, 105, 153, 124, 92, 85, 88, 134, 97, 123, 0, 0, 0, 156, 134, 
    117, 133, 120, 343, 123, 349, 15, 115, 104, 122, 119, 226, 241, 301, 101, 
    58, 349, 245, 176, 36, 95, 88, 100, 179, 281, 277, 253, 272, 279, 283, 
    272, 292, 293, 295, 257, 290, 299, 310, 305, 317, 309, 284, 305, 272, 
    254, 289, 282, 133, 95, 71, 79, 93, 126, 153, 291, 267, 285, 282, 287, 
    269, 268, 267, 278, 259, 274, 287, 281, 285, 290, 299, 272, 278, 283, 
    276, 282, 266, 287, 285, 271, 273, 302, 264, 270, 292, 312, 287, 280, 
    294, 287, 307, 303, 317, 321, 302, 310, 311, 171, 176, 176, 163, 165, 
    162, 165, 171, 164, 167, 175, 155, 144, 133, 130, 129, 90, 59, 25, 343, 
    0, 349, 337, 97, 101, 147, 129, 131, 118, 114, 90, 121, 140, 153, 164, 
    97, 104, 83, 86, 92, 95, 90, 87, 110, 114, 75, 158, 131, 120, 142, 123, 
    131, 143, 140, 160, 135, 133, 116, 147, 126, 121, 90, 314, 298, 308, 300, 
    297, 294, 291, 303, 92, 83, 76, 81, 170, 110, 115, 121, 116, 123, 96, 
    138, 91, 68, 99, 100, 100, 115, 105, 22, 0, 0, 360, 307, 315, 296, 172, 
    150, 156, 70, 112, 121, 99, 115, 120, 130, 335, 260, 185, 10, 286, 299, 
    319, 315, 300, 291, 303, 301, 332, 284, 295, 291, 294, 297, 285, 293, 
    288, 219, 316, 239, 85, 113, 333, 291, 284, 267, 290, 270, 263, 279, 309, 
    338, 318, 303, 308, 314, 272, 325, 181, 297, 260, 343, 211, 225, 194, 
    256, 267, 273, 284, 296, 311, 305, 287, 297, 289, 291, 293, 294, 291, 
    289, 289, 280, 270, 273, 272, 242, 275, 209, 278, 266, 175, 176, 165, 
    304, 191, 307, 172, 312, 319, 64, 89, 100, 92, 95, 103, 113, 110, 108, 
    97, 104, 115, 114, 122, 102, 128, 116, 136, 130, 125, 100, 360, 2, 0, 71, 
    105, 9, 360, 360, 121, 101, 142, 189, 138, 160, 136, 0, 296, 305, 178, 
    325, 296, 313, 329, 343, 332, 331, 183, 1, 52, 162, 126, 124, 132, 150, 
    179, 173, 227, 277, 242, 272, 264, 290, 311, 297, 293, 298, 289, 290, 
    289, 300, 188, 318, 74, 224, 156, 140, 123, 125, 145, 138, 141, 140, 116, 
    89, 104, 46, 129, 103, 163, 286, 255, 6, 170, 106, 356, 279, 343, 20, 
    343, 317, 84, 257, 126, 96, 161, 157, 116, 112, 115, 95, 37, 112, 289, 
    291, 75, 356, 360, 90, 107, 98, 329, 332, 298, 292, 94, _, 293, 294, 299, 
    182, 162, 164, 165, 170, 226, 79, 82, 97, 348, 326, 0, 0, 295, 130, 128, 
    116, 113, 98, 102, 166, 209, 108, 135, 138, 236, 263, 182, 145, 123, 163, 
    0, 359, 174, 342, 0, 305, 228, 270, 95, 129, 158, 147, 115, 153, 295, 
    211, 126, 141, 108, 54, 90, 67, 113, 60, 78, 306, 287, 197, 341, 248, 94, 
    249, 198, 31, 287, 20, 64, 65, 55, 49, 23, 85, 90, 99, 128, 161, 113, 
    182, 270, 287, 290, 285, 285, 293, 288, 281, 298, 307, 283, 275, 296, 
    315, 266, 272, 269, 267, 296, 270, 269, 266, 282, 290, 290, 280, 291, 
    280, 305, 79, 284, 250, 314, 223, 174, 335, 308, 64, 59, 76, 56, 80, 76, 
    190, 59, 60, 263, 72, 174, 271, 234, 80, 338, 313, 250, 0, 309, 282, 217, 
    0, 15, _, _, _, 127, 50, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, 129, 136, _, 114, 117, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 162, 163, 173, 169, 167, 167, _, _, 129, 152, 148, 134, 
    116, 155, 167, 179, 166, 170, 180, 185, 302, 175, 151, 93, 116, 109, 139, 
    118, 107, 128, 159, 156, 152, 200, 200, 240, 240, 281, 309, 291, 300, 
    315, 327, 283, 276, 96, 92, 88, 84, 98, 91, 100, 123, 124, 123, 120, 100, 
    73, 170, 147, 146, 161, 155, 148, 140, 133, 125, 118, 155, 284, 305, 282, 
    57, 311, 304, 314, 14, 326, 354, 253, 200, 157, 171, _, _, _, _, _, 54, 
    62, 0, _, _, _, 293, 184, _, _, _, _, _, _, _, _, _, _, _, _, _, 359, 
    163, 93, 34, 0, 0, 47, 251, _, _, _, _, 112, 119, 107, 108, _, 123, 119, 
    118, 121, 124, 119, _, _, _, _, _, _, _, 97, 113, 151, _, 114, 112, 158, 
    137, 113, 119, 103, _, 118, _, 113, _, 96, 102, 102, 102, 105, 77, 270, 
    288, 8, _, _, _, 307, 128, 116, 155, 132, 129, 143, 132, 132, 129, 127, 
    126, 126, 0, 353, 51, 0, 100, 95, 105, 110, 90, 115, 80, 110, 149, 130, 
    146, 117, 104, 133, 123, 122, 120, 119, 126, 100, 54, 31, 351, 309, 356, 
    339, 322, 319, 280, 288, 282, 238, 332, 274, 185, 160, 111, 280, 251, 
    214, 176, 142, 109, 75, 44, 13, 89, 359, 322, 312, 178, 284, 4, 57, _, 
    244, 207, 182, 179, 127, _, _, _, 241, 114, _, _, 140, 285, 299, 194, 
    336, 314, 89, 152, 12, _, _, _, 290, 100, 129, 115, 241, 190, 100, 106, 
    107, 262, 127, 79, 225, 227, 230, 313, 112, 97, 343, 353, 35, 337, 124, 
    130, 138, 127, 158, 99, 194, 136, 90, 21, _, _, 60, _, 0, _, 315, 63, 
    355, 83, 97, 77, 163, _, _, _, 204, 120, 162, 101, 111, _, 198, 121, 116, 
    _, _, _, _, _, _, _, _, _, _, 315, 5, 341, 122, 69, 142, 130, 253, 147, 
    144, 88, 62, 146, 53, 129, _, 77, _, _, _, _, _, _, _, 157, 339, _, _, 
    146, _, _, 274, _, 94, 70, 80, 137, _, 87, 53, 239, 340, _, _, 304, 316, 
    355, 319, 305, 14, _, _, _, 350, 139, _, 125, 129, 139, 148, 128, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 89, 15, 275, _, 249, 256, 73, 62, 
    148, _, _, _, _, _, _, _, _, 63, 68, 74, 106, 47, 87, _, _, 68, 67, _, _, 
    68, 93, 77, _, 77, _, _, _, _, _, _, _, 325, 315, _, 327, 329, 37, 279, 
    358, _, 291, _, _, 89, 77, 69, 63, 75, 216, 248, 274, 318, _, _, 315, _, 
    0, 33, 5, 324, _, 0, 0, _, 143, 136, 131, 129, 139, 140, 126, 131, 123, 
    130, _, 138, 310, 9, 29, 0, 358, 58, 74, _, _, 0, 295, 292, 284, 298, 
    293, 277, 262, 158, 133, 140, 121, 130, 130, 123, 339, 337, 317, _, _, _, 
    _, 356, 339, 306, 0, 275, 256, 132, 136, 139, 132, 92, 150, _, 99, 128, 
    0, 308, 116, 302, 323, 299, 321, _, 29, 341, 277, 294, 322, 322, 109, 
    341, 99, 358, 112, 107, 71, 231, 296, 270, 278, 257, 241, 253, 265, 270, 
    269, 260, 269, 278, 288, 283, 282, 268, 268, 266, 265, 266, 266, 288, 
    292, 288, 289, 288, 268, 281, 279, 277, 282, 275, 298, 307, 310, 309, 
    298, 304, 295, 286, 278, 291, 263, 263, 294, 284, 197, 292, 274, 289, 
    290, 291, 329, 342, 359, 351, 346, 326, 322, 336, 322, 320, 319, 308, 
    269, 262, 266, 290, 271, 268, 266, 268, 272, 274, 288, 274, 271, 280, 
    288, 309, 301, 283, 324, 325, 328, 263, 35, 323, 84, 85, 78, 72, 63, 67, 
    67, 64, 59, 50, 285, 209, 263, 340, 302, 10, 0, 325, 0, 358, 353, 357, 
    339, 347, 342, 219, 96, 96, 133, 95, 92, 88, 92, 89, 88, 108, 103, 99, 
    94, 99, 110, 109, 118, 121, 118, 120, 119, 120, 119, 118, 113, 113, 106, 
    115, 110, 111, 113, 115, 114, 113, 112, 111, 110, 110, 109, 108, 107, 
    106, 105, 116, 96, 101, 108, 102, 100, 113, 110, 110, 105, 115, 120, 120, 
    150, 150, 140, 28, 310, 298, 302, 303, 312, 315, 321, 313, 310, 307, 348, 
    123, 358, 59, 181, 177, 164, _, _, _, _, _, _, 321, 58, 339, 320, 275, 
    299, 301, 349, 308, _, _, _, _, 284, 270, 106, 155, 300, 285, 295, 290, 
    293, _, _, _, 216, 185, 11, 38, 43, 51, 54, 51, _, _, _, _, _, _, 90, 56, 
    23, 58, 44, 36, 332, 62, 64, _, _, _, 318, 301, 328, 351, 0, 308, 71, 
    300, 251, 0, 47, 250, 83, 73, 96, 0, 67, 0, _, _, 278, 319, 275, 298, 26, 
    320, 310, 292, _, 87, 25, 215, 242, 32, 139, 145, 173, _, 99, 357, 328, 
    316, 355, 338, 345, _, _, _, _, _, _, _, 266, 299, 314, 295, 13, _, 311, 
    284, 218, 261, 311, 293, 330, 300, 1, 303, 13, _, _, _, _, _, _, _, _, 
    338, 301, 281, 297, 313, 277, 290, 102, 47, 128, 300, 323, 89, 360, 342, 
    303, 324, 322, _, _, _, 293, 317, 304, 320, 9, 53, 50, 8, 83, 17, 304, 
    250, 351, 301, 239, 7, 282, _, _, _, 25, 37, 246, 311, 250, 336, 97, 319, 
    _, _, _, 306, 299, 314, 319, 309, 306, 314, 303, 296, _, _, 313, 304, 
    294, 290, _, 293, 285, 293, 291, _, 284, 284, 286, 280, 293, 282, 281, 
    283, 273, 270, 286, 281, _, 287, 286, 285, _, _, 311, 310, 325, 309, 41, 
    357, 301, 351, 348, 257, 233, 266, 233, 294, 348, 0, 292, 236, 66, _, _, 
    _, _, 336, 301, 157, 326, 290, 149, 97, 322, 118, _, _, 97, 353, 27, 58, 
    0, 82, 58, 285, 301, _, _, 301, 270, 281, _, 276, 269, 263, 281, 296, 
    287, _, _, 274, 273, 281, 278, 271, 271, 281, 290, 295, _, _, 290, 292, 
    286, 291, 288, 290, 284, 290, 294, _, _, 289, 288, 282, 294, 289, 287, 
    284, 297, _, _, _, _, _, _, _, _, 286, _, 274, 281, 282, 289, 282, 280, 
    275, _, 277, 287, 293, 289, 295, 319, 292, 317, 316, _, _, _, _, _, 0, _, 
    306, _, 355, _, _, _, 310, _, 290, 355, 306, 316, 327, 265, _, 353, 259, 
    _, 114, 234, _, 6, 3, 0, 15, _, 158, 264, 320, 207, 310, 30, _, _, _, _, 
    _, _, _, 244, 22, 10, 350, 309, 320, _, 334, _, _, _, _, _, 327, 317, 
    271, 294, 0, 0, 359, _, _, _, _, 300, 63, 60, 32, _, 267, 311, 291, _, _, 
    322, 309, 340, 325, 33, _, _, 297, _, _, 290, 299, 295, 273, 288, 298, _, 
    283, 268, 254, _, 278, 302, _, 281, _, _, _, 302, 304, 306, 313, 298, _, 
    _, 321, 283, 312, 299, 302, 296, 279, 306, _, _, _, _, _, 316, 209, _, 4, 
    317, 329, _, 90, 22, _, 126, 90, 111, 88, 101, _, 123, 130, 79, 80, 319, 
    290, 356, _, _, _, 178, 279, _, 48, 57, 29, 41, 57, 54, 71, 74, 44, 47, 
    34, 26, _, 290, _, 73, _, 241, _, 89, _, 205, 272, 151, 201, 41, _, 18, 
    _, 65, 21, 72, _, _, _, 192, _, 324, 224, _, _, 252, 226, 341, 54, 355, 
    4, 347, 246, 4, 328, _, _, _, 63, 39, 156, 75, 56, 65, 56, 63, _, _, _, 
    14, 300, 5, _, _, 40, 3, 0, _, 157, 359, 294, 320, 284, _, 302, 304, 306, 
    _, 354, 4, 333, 286, 329, 282, 271, 332, 337, _, _, _, 317, 311, 337, 
    340, _, 301, 135, 267, _, _, _, 294, _, 313, 0, _, 334, _, 346, _, _, _, 
    _, _, _, _, 290, 306, 293, _, 304, 1, 293, 286, 301, 313, 279, 332, _, 
    105, _, _, 74, _, _, 70, 312, _, 285, 310, 62, 23, 318, 22, 119, 322, 0, 
    _, _, _, 352, _, _, _, 348, 293, 327, _, _, _, 308, 9, 338, 358, 312, 
    299, _, _, 68, _, 302, 349, 337, 327, _, 89, _, _, 90, _, 91, _, 77, _, 
    75, 81, 87, _, 94, 60, 92, 65, 71, 65, 326, 324, 42, _, _, 75, _, _, 318, 
    318, _, 83, 297, _, _, _, _, _, _, _, _, _, _, 79, 337, 312, 46, _, 286, 
    20, 311, 322, _, 340, 334, _, 309, _, 312, _, _, _, _, _, 318, _, 297, _, 
    300, 305, _, 309, _, 311, _, 286, _, _, 294, 327, 343, _, 312, 322, _, _, 
    312, 312, 249, _, 329, 184, 198, 190, 233, 3, 115, 215, _, _, _, _, _, 
    296, 301, 131, 343, 315, 284, 306, 325, 314, 318, 294, 293, 311, 252, 
    312, 294, _, 282, 301, 327, 327, 288, 277, 0, 308, 296, 282, _, _, _, 
    323, 268, 281, 287, 331, 0, 300, 321, 313, 339, 333, _, _, _, _, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, _, 0, 0, 0, 19, 312, 273, 323, 331, 15, _, 310, 335, 
    331, 318, _, 322, 349, 310, 310, _, 294, 319, 312, 278, 0, 221, 32, 344, 
    358, _, 319, 336, 308, _, 307, _, 331, 315, 329, _, 320, 1, 332, 325, 4, 
    52, 340, 314, 357, _, _, 327, _, 310, 353, 318, 332, 348, _, _, 10, 45, 
    21, _, 53, 1, 303, 334, 339, _, 297, 289, 298, 295, 313, 273, 308, 290, 
    7, _, _, 287, 278, 287, 268, 350, 300, 314, 295, 310, _, _, _, 280, 302, 
    306, 295, 283, 322, 313, 301, 301, _, _, 279, _, 49, 35, 38, 56, 47, 57, 
    50, _, _, 188, 303, 264, 259, 297, 322, 332, 312, _, 9, 320, 338, 311, 
    333, 340, 325, 299, 340, _, _, _, _, 12, 18, 32, 49, 25, 107, _, 28, 11, 
    _, 351, 312, 353, 36, 47, 44, 39, 37, _, _, _, 42, 28, 43, 40, 35, 44, 
    26, 34, 33, _, 35, 274, 232, 329, 353, 1, 256, 277, _, _, _, 299, 319, 
    310, 311, 321, 318, 318, 322, 326, _, _, _, 321, 287, 308, 293, 260, 281, 
    288, 320, _, _, _, _, _, _, _, _, _, 296, 316, 352, 340, 293, 297, 294, 
    277, 291, 303, 294, _, 287, 293, 300, 305, _, _, _, _, _, _, 324, 329, 
    298, 293, 310, 322, 352, 24, _, _, 312, 352, 353, 318, 316, 351, 340, 
    351, 315, _, 308, 347, 301, 316, 308, 11, 349, 332, 83, 351, 320, 8, 316, 
    61, 331, _, 322, 337, 334, 336, _, _, _, 322, _, _, _, _, 322, 1, 326, 
    350, 358, 297, 305, 293, 308, _, _, _, _, 45, 10, 109, 13, 78, 31, 51, 
    324, _, _, _, _, _, _, _, _, _, 288, 340, 310, 329, 34, 330, 44, 303, 
    318, _, _, 350, 308, 265, 311, 28, 318, 347, 304, _, _, _, _, 96, 80, 81, 
    89, 97, 112, 83, 55, 306, _, 321, _, _, _, 89, 78, 86, 70, 88, _, _, 96, 
    85, 86, 94, 92, 89, 85, 90, 87, _, _, 308, 316, 67, 359, 22, 52, 323, 7, 
    346, _, _, 78, 96, 77, 87, 79, 90, 92, 86, 84, _, 89, 81, 77, 90, 95, 85, 
    99, 101, 104, _, _, _, 91, 120, 109, 103, 69, 59, 46, 43, _, _, _, 41, 
    44, 50, 63, 48, 53, 79, 82, _, _, _, _, _, 97, 76, 96, 98, 102, 95, 95, 
    111, 95, 110, 98, 91, 96, 94, 88, 97, 97, 94, 99, 100, 98, 98, _, 97, 98, 
    97, _, _, _, _, _, 100, 94, 88, 92, 83, 100, 96, 86, 82, 84, 94, 105, 91, 
    79, 73, 116, 103, 90, 94, 81, 93, 94, 89, 69, 58, 70, 75, 72, 275, 304, 
    315, 295, 320, 292, 293, 314, 303, 0, 0, 301, 303, 297, 322, 324, 316, 
    302, 315, 4, 305, 40, 350, 355, 319, 339, 318, 283, 310, 290, 300, 286, 
    292, 358, 323, 317, 341, 328, 324, 343, 336, 0, 319, 7, 0, 346, 316, 352, 
    320, 296, 318, 309, 314, 337, 344, 296, 326, 303, 318, 1, 347, 336, 333, 
    347, 2, 298, 276, 326, 337, 327, 335, 312, 354, 342, 59, 60, 79, 77, 50, 
    55, 46, 46, 50, 39, 37, 57, 53, 12, 12, 348, 39, 81, 69, 44, 140, 275, 
    281, 287, 306, 302, 287, 285, 328, 261, 289, 281, 324, 338, 59, 270, 45, 
    314, 235, 294, 266, 303, 302, 318, 303, 301, 297, 310, 295, 278, 292, 
    291, 286, 307, 304, 287, 278, 278, 287, 296, 295, 280, 284, 296, 307, 
    305, 327, 323, 0, 325, _, 296, 323, 329, 329, 48, 8, 26, 184, 9, 269, 
    102, 334, 310, 348, 331, 328, 309, 326, 320, 311, 313, 319, 317, 313, 
    304, 320, 313, 310, 316, 310, 313, 307, 301, 309, 323, 9, 302, 313, 347, 
    344, 299, 285, 69, 82, 87, 89, 87, 74, 76, 57, 74, 304, 304, 317, 59, 
    320, 329, 23, 37, 328, 2, 58, 37, 44, 49, 57, 42, 39, 50, 48, 9, 18, 33, 
    64, 145, 13, 79, 48, _, 16, 48, 32, 37, 38, 37, 34, 37, 29, 25, 22, 7, _, 
    3, 16, 10, 7, 13, 359, 17, 22, 39, 35, 36, 38, 39, 45, 45, 44, 39, 38, 
    25, 13, 15, 327, 240, 299, 302, 307, 306, 329, 313, 317, 330, 339, 298, 
    267, 311, 320, 300, 338, 312, 285, 314, 314, 296, 324, 335, 340, 14, 340, 
    342, 358, 194, 46, 47, 204, 201, 345, 300, 318, 293, 288, 315, 289, 290, 
    301, 331, 323, 294, 312, 311, 307, 303, 325, 315, 303, 324, 300, 261, 
    310, 295, 300, 307, 271, 300, 287, 295, 311, 280, 299, 290, 351, 299, 
    276, 339, 166, 225, 296, 90, 296, 226, 203, 138, 345, 262, 28, 312, 157, 
    18, 311, 360, 6, 311, 306, 302, 312, 298, 320, 320, 295, 292, 342, 290, 
    295, 324, 300, 310, 336, 313, 289, 354, 316, 257, 284, 322, 319, 326, 
    315, 297, 303, 315, 334, 36, 314, 57, 263, 257, 274, 301, 295, 292, 280, 
    289, 270, 281, 275, 286, 281, 269, 297, 301, 317, 310, 344, 4, 271, 10, 
    334, 316, 246, 326, 66, 323, 43, 319, 323, 328, 321, 319, 347, 328, 325, 
    310, 304, 316, 314, 301, 310, 318, 315, 281, 321, 330, 359, 299, 21, 57, 
    26, 319, 0, 324, 336, 314, 10, 339, 320, 9, 307, 318, 327, 287, 296, 316, 
    50, 100, 311, 283, 345, 358, 299, 302, 19, 317, 338, 325, 303, 275, 11, 
    324, 335, 40, 320, 349, 48, 47, 352, 325, 314, 54, 337, 323, 359, 62, 
    354, 15, 341, 13, 321, 43, 45, 38, 40, 51, 131, 29, 19, 46, 47, 330, 310, 
    298, 320, 5, 309, 341, 311, 324, 298, 342, 315, 318, 244, 305, 330, 315, 
    48, 329, 288, 277, 290, 108, 97, 92, 85, 81, 323, 284, 300, 289, 285, 
    333, 304, 298, 321, 0, 312, 354, 31, 75, 297, 317, 5, 347, 305, 350, 17, 
    307, 15, 359, 0, 37, 328, 293, 12, 23, 337, 27, 283, 299, 23, 294, 306, 
    295, 294, 278, 301, 289, 296, 302, 269, 309, 288, 309, 306, 316, 305, 
    313, 330, 306, 289, 288, 299, 288, 279, 280, 289, 296, 272, 286, 268, 
    289, 270, 262, 273, 274, 275, 270, 263, 339, 296, 20, 47, 48, 11, 360, 
    248, 347, 330, 316, 329, 329, 312, 303, 356, 352, 347, 320, 287, 276, 
    292, 322, 301, 313, 359, 7, 6, 1, 63, 40, 27, 0, 318, 4, 135, 32, 294, 
    94, 34, 23, 336, 45, 81, 356, 18, 8, 303, 12, 311, 345, 313, 354, 335, 
    119, 24, 76, 58, 83, 109, 293, 307, 277, 290, 297, 318, 312, 330, 99, 13, 
    12, 14, 337, 8, 346, 307, 131, 298, 75, 360, 352, 273, 290, 10, 326, 333, 
    299, 200, 168, 276, 314, 320, 282, 316, 311, 330, 313, 316, 315, 310, 
    300, 296, 279, 288, 35, 197, 296, 324, 330, 355, 331, 318, 27, 1, 24, 29, 
    350, 10, 291, 339, 331, 277, 310, 320, 338, 293, 286, 336, 306, 302, 274, 
    310, 288, 293, 321, 320, 314, 299, 300, 318, 348, 315, 10, 70, 13, 4, 
    290, 0, 31, 331, 15, 322, 304, 272, 305, 309, 69, 9, 73, 0, 14, 80, 92, 
    306, 19, 31, 322, 41, 355, 317, 351, 0, 321, 95, 281, 349, 307, 316, 320, 
    312, 300, 298, 101, 88, 98, 97, 102, 95, 109, 96, 117, 92, 94, 100, 118, 
    96, 100, 95, 96, 93, 95, 95, 95, 94, 95, 98, 96, 95, 98, 97, 95, 95, 94, 
    90, 94, 95, 91, 97, 95, 107, 109, 115, 120, 112, 97, 107, 110, 88, 79, 
    111, 84, 95, 99, 89, 95, 111, 101, 104, 98, 98, 47, 47, 89, 96, 46, 67, 
    76, 62, 68, 118, 80, 63, 56, 284, 283, 323, 340, 342, 351, 335, 332, 293, 
    320, 306, 334, 304, 332, 313, 293, 285, 300, 308, 313, 285, 58, 98, 97, 
    103, 98, 98, 80, 76, 90, 109, 104, 107, 116, 110, 103, 102, 90, 95, 103, 
    108, 117, 120, 123, 137, 115, 65, 48, 78, 348, 30, 228, 316, 76, 37, 91, 
    336, 281, 9, 352, 357, 3, 34, 35, 30, 26, 32, 1, 358, 333, 84, 42, 70, 
    89, 73, 61, 50, 62, 50, 42, 75, 64, 82, 99, 67, 51, 37, 36, 83, 38, 37, 
    2, 33, 14, 16, 360, 44, 22, 39, 38, 38, 36, 34, 36, 34, 42, 46, 45, 19, 
    16, 310, 328, 331, 316, 328, 315, 322, 308, 301, 305, 337, 340, 349, 334, 
    292, 23, 323, 310, 311, 305, 297, 284, 306, 304, 305, 299, 313, 360, 16, 
    5, 342, 328, 328, 327, 282, 316, 311, 322, 25, 305, 315, 321, 333, 322, 
    19, 95, 177, 165, 23, 202, 11, 19, 20, 13, 30, 338, 340, 350, 356, 357, 
    82, 200, 280, 300, 355, 319, 354, 3, 4, 25, 32, 27, 2, 356, 345, 59, 28, 
    345, 292, 281, 243, 326, 338, 360, 20, 24, 324, 306, 303, 54, 323, 4, 44, 
    147, 162, 124, 97, 187, 182, 306, 205, 250, 241, 300, 314, 317, 293, 303, 
    297, 302, 300, 299, 291, 301, 300, 275, 271, 310, 286, 316, 345, 350, 
    323, 229, 316, 2, 360, 333, 322, 295, 348, 325, 33, 353, 309, 67, 4, 334, 
    350, 357, 352, 43, 319, 65, 143, 2, 130, 288, 322, 275, 323, 293, 300, 
    302, 293, 300, 317, 307, 305, 289, 285, 282, 273, 273, 278, 287, 274, 
    291, 287, 289, 305, 309, 324, 318, 319, 320, 324, 327, 307, 299, 358, 
    351, 92, 12, 64, 96, 14, 315, 316, 317, 300, 296, 284, 275, 290, 275, 
    290, 294, 284, 280, 299, 312, 297, 311, 285, 297, 321, 304, 303, 318, 
    348, 5, 354, 332, 346, 327, 335, 39, 40, 306, 320, 354, 330, 322, 314, 
    324, 340, 43, 15, 327, 13, 318, 303, 339, 333, 320, 337, 37, 221, 317, 
    247, 345, 129, 246, 321, 299, 28, 354, 21, 52, 37, 19, 318, 286, 252, 17, 
    26, 6, 220, 215, 251, 21, 217, 301, 17, 12, 11, 12, 35, 35, 12, 360, 282, 
    357, 49, 331, 263, 6, 28, 355, 21, 3, 213, 75, 332, 353, 32, 54, 202, 43, 
    45, 314, 336, 321, 305, 61, 332, 35, 353, 344, 314, 355, 347, 345, 335, 
    357, 6, 22, 26, 336, 347, 37, 307, 9, 319, 11, 6, 338, 345, 335, 309, 
    355, 323, 313, 312, 317, 346, 343, 336, 346, 342, 327, 330, 335, 314, 
    293, 270, 272, 61, 40, 185, 25, 162, 337, 174, 340, 281, 346, 161, 355, 
    276, 284, 68, 338, 292, 240, 334, 35, 229, 202, 254, 305, 301, 200, 131, 
    312, 6, 267, 129, 14, 138, 174, 313, 310, 30, 18, 21, 213, 11, 199, 335, 
    330, 360, 328, 300, 204, 295, 3, 4, 5, 7, 360, 32, 314, 12, 272, 21, 29, 
    23, 13, 68, 308, 117, 328, 17, 5, 360, 321, 273, 347, 303, 160, 123, 332, 
    40, 360, 342, 310, 30, 190, 180, 239, 178, 296, 295, 346, 35, 121, 306, 
    187, 299, 321, 341, 331, 311, 339, 313, 327, 338, 293, 305, 298, 318, 
    323, 333, 329, 325, 320, 324, 317, 307, 312, 324, 59, 354, 58, 330, 321, 
    2, 92, 337, 109, 332, 360, 358, 19, 319, 81, 101, 333, 325, 316, 283, 
    341, 76, 83, 87, 83, 70, 82, 90, 90, 83, 95, 93, 98, 100, 108, 107, 92, 
    100, 106, 111, 121, 75, 50, 352, 285, 290, 299, 126, 319, 80, 303, 10, 
    324, 321, 324, 343, 103, 94, 107, 98, 87, 79, 79, 73, 96, 97, 90, 105, 
    67, 91, 88, 95, 80, 75, 24, 34, 29, 32, 36, 9, 33, 40, 48, 11, 42, 34, 
    55, 44, 44, 44, 58, 48, 355, 133, 108, 333, 352, 13, 19, 303, 66, 1, 330, 
    340, 359, 340, 325, 43, 355, 23, 321, 17, 320, 33, 20, 347, 329, 306, 
    360, 1, 72, 351, 354, 315, 69, 309, 328, 335, 333, 326, 8, 318, 0, 357, 
    7, 356, 324, 307, 78, 67, 344, 136, 0, 341, 59, 2, 50, 0, 0, 0, 0, 0, 0, 
    0, 0, 72, 110, 92, 105, 101, 94, 57, 85, 87, 63, 76, 89, 81, 82, 89, 87, 
    81, 78, 109, 53, 319, 320, 340, 353, 331, 344, 322, 315, 311, 311, 345, 
    333, 350, 349, 25, 358, 323, 15, 329, 352, 55, 29, 327, 333, 314, 20, 
    314, 345, 324, 359, 35, 327, 330, 341, 336, 309, 42, 62, 307, 276, 293, 
    258, 303, 337, 311, 313, 334, 42, 86, 323, 326, 321, 340, 353, 331, 322, 
    356, 320, 305, 286, 1, 356, 62, 70, 61, 3, 84, 104, 41, 21, 171, 94, 109, 
    71, 90, 112, 84, 83, 87, 70, 86, 87, 79, 63, 314, 309, 303, 0, 308, 81, 
    284, 332, 339, 86, 288, 284, 355, 310, 325, 37, 315, 15, 354, 354, 74, 
    98, 84, 87, 93, 74, 87, 91, 89, 82, 95, 107, 91, 84, 84, 141, 66, 66, 78, 
    75, 70, 64, 66, 58, 89, 64, 68, 63, 60, 337, 53, 50, 45, 1, 330, 314, 
    307, 292, 56, 360, 354, 1, 282, 46, 360, 317, 309, 18, 80, 325, 326, 35, 
    356, 317, 64, 41, 62, 81, 115, 110, 99, 99, 94, 69, 108, 98, 95, 87, 69, 
    62, 64, 63, 72, 87, 346, 284, 304, 302, 302, 320, 303, 325, 359, 339, 0, 
    317, 354, 22, 359, 296, 320, 3, 1, 353, 39, 334, 352, 360, 4, 67, 20, 
    311, 21, 333, 324, 321, 356, 350, 343, 321, 11, 14, 8, 100, 66, 119, 115, 
    113, 114, 57, 60, 78, 80, 66, 327, 318, 320, 69, 75, 80, 76, 79, 60, 66, 
    70, 94, 106, 77, 99, 285, 330, 335, 311, 287, 331, 33, 315, 326, 294, 
    330, 321, 322, 325, 322, 296, 326, 10, 327, 298, 325, 311, 319, 316, 321, 
    8, 320, 346, 319, 333, 300, 296, 314, 310, 312, 322, 320, 325, 311, 85, 
    93, 91, 84, 110, 33, 82, 73, 103, 81, 310, 281, 323, 301, 282, 341, 292, 
    307, 316, 318, 345, 287, 356, 332, 292, 306, 294, 327, 318, 317, 320, 
    321, 314, 330, 340, 352, 18, 307, 333, 342, 322, 351, 325, 25, 343, 0, 7, 
    6, 301, 308, 345, 304, 319, 47, 319, 72, 294, 349, 85, 46, 329, 0, 351, 
    126, 34, 294, 318, 302, 305, 311, 313, 306, 355, 60, 354, 305, 296, 321, 
    295, 287, 309, 100, 101, 0, 360, 14, 296, 285, 291, 290, 298, 280, 290, 
    301, 315, 306, 313, 300, 284, 306, 286, 291, 299, 307, 315, 300, 297, 
    324, 325, 319, 112, 18, 304, 334, 349, 324, 0, 335, 57, 315, 6, 16, 310, 
    322, 327, 325, 322, 70, 311, 318, 93, 340, 307, 86, 110, 304, 353, 59, 
    324, 352, 288, 290, 300, 298, 78, 326, 0, 0, 277, 268, 271, 274, 268, 
    268, 268, 281, _, 277, 276, 262, 262, 265, _, 260, 269, 259, 262, 269, 
    260, 280, 256, 267, 263, 265, 262, 267, 270, _, 243, 288, 300, 284, 307, 
    276, 307, 52, 335, 340, 62, 323, 26, 54, 352, 32, 332, 60, 39, 294, 360, 
    55, 336, 11, 13, 292, 309, 317, 77, 11, 323, 343, 234, 39, 85, 80, 86, 
    107, 86, 77, 76, 93, 318, 92, 62, 66, 133, 324, 45, 208, 45, 347, 0, 351, 
    15, 58, 316, 61, 23, 1, 110, 90, 86, 81, 80, 99, 98, 100, 107, 97, 112, 
    107, 97, 99, 105, 111, 110, 111, 112, 104, 112, 111, _, 104, 84, 123, 96, 
    _, 87, _, _, 99, _, 96, 78, 86, 102, 98, 88, _, _, 70, 353, 103, 118, 57, 
    9, 13, 334, _, 317, _, 321, 16, 325, _, 26, _, 347, 328, _, 313, 314, 
    295, 69, 307, 356, 48, 345, 0, 340, 360, 358, 331, 340, 347, 76, 73, 80, 
    60, 39, 66, 320, 5, 317, 358, 328, 69, 347, 311, 82, 359, 344, 27, 333, 
    349, 337, 305, 26, 333, 297, 24, 337, 347, 47, 305, 65, 340, 58, 312, 
    357, 82, 320, 313, 31, 336, 67, 70, 80, 88, 35, 356, 360, 335, 93, 9, 
    354, 90, 312, 355, 356, 90, 70, 63, 70, 88, 359, 331, 18, 172, 316, 87, 
    357, 13, 355, 300, 342, 310, 312, 312, 350, 315, 22, 333, 360, 0, 333, 
    65, 72, 305, 342, 324, 328, 279, 338, 303, 331, 326, 319, 14, 30, 65, 
    360, 0, 329, 54, 73, 79, 320, 310, 296, 323, 348, 348, 91, 86, 333, 31, 
    354, 284, 89, 360, 342, 43, 24, 314, 360, 39, 90, 338, 12, 99, _, 300, _, 
    87, _, 315, 84, 107, 332, 114, 345, 280, 245, 248, 216, 212, 211, 205, 
    223, 203, 209, 209, 207, 205, 205, 207, 180, 48, 178, 106, 115, 110, 88, 
    13, 131, 145, 155, 87, 90, 103, 157, 138, 169, 142, 149, 300, 305, 13, 
    188, 257, 293, 238, 230, 162, 257, 23, 210, 196, 187, 28, 33, 55, 257, 
    108, 98, 354, 31, _, 329, 293, _, 308, 315, _, _, _, _, 295, 299, 306, 
    274, 187, 13, 293, 196, 286, 45, 247, 215, 270, _, 260, 225, _, 263, 307, 
    _, 297, 256, _, 41, 309, _, 313, 289, _, 19, 292, 11, 7, 9, 10, _, _, 
    356, _, 26, _, 24, 213, 12, _, 198, _, 142, 313, 319, 293, 302, 327, 342, 
    _, 12, 43, _, 324, 358, 4, 356, _, _, _, 308, 337, 311, 61, 334, 91, _, 
    7, 69, 68, 327, 306, 5, 13, 329, 312, 345, 314, 305, 23, 355, _, 356, 
    334, 318, 9, 0, 308, 34, 348, 352, 307, 294, 70, 327, 329, 340, 7, 5, 
    338, 6, 341, 5, 73, 57, 99, 62, _, 88, 80, 25, 39, 74, 260, 144, 233, _, 
    297, 248, 240, 11, 133, 82, 31, 315, 11, 59, 261, 80, _, 76, 162, 49, 70, 
    306, 128, 11, 59, 100, 126, 163, 336, 314, 302, 315, 341, 270, 100, 344, 
    359, 309, 301, 343, 325, 358, 325, 327, 323, 7, 328, 306, 317, 333, 325, 
    309, 341, 323, 71, 339, 29, 45, 360, 46, 21, 303, 309, 343, 357, 52, 55, 
    15, 329, 12, 344, 355, 331, 5, 319, 17, 60, 104, 350, 81, 293, 316, 31, 
    62, 64, 308, 311, 46, 88, 98, 5, 47, 90, 341, 319, 72, 89, 97, 90, 87, 
    88, 90, 93, 75, 76, 307, 298, 317, 187, 115, 326, 31, 234, 342, 53, 45, 
    106, 92, 31, 285, 300, 282, 278, 276, 195, 273, 253, 309, 278, 274, 280, 
    277, 277, 277, 287, 292, 310, 303, 304, 79, 48, 15, 359, 21, 322, 335, 
    307, 336, 327, 309, 322, 68, 89, 325, 96, 338, 342, 18, 332, 30, _, _, 5, 
    31, 36, 35, 37, 38, 36, 35, 31, 27, 40, 38, 39, 352, 27, 42, 31, 35, 40, 
    40, 42, 43, 36, 40, 45, 69, 41, 40, 42, 27, 15, 95, 66, 346, 280, 353, 
    328, 316, 354, 330, 261, 309, 309, 324, 163, 277, 229, 303, 353, 276, 
    315, 312, 329, 321, 317, 68, 336, 76, 25, 316, 335, 57, 302, 327, 349, 6, 
    38, 349, 330, 317, 324, 360, 56, 348, 26, 304, 70, 64, 353, 109, 6, 331, 
    42, 9, 307, 31, 335, 325, 88, 241, 17, 346, 308, 3, 349, 89, 316, 334, 3, 
    5, 309, 78, 92, 336, 325, 82, 61, 324, 332, 15, 118, 320, 329, 72, 66, 0, 
    6, 51, 320, 112, 313, 84, 4, 59, 303, 37, 76, 323, 324, 344, 1, 96, 353, 
    329, 333, 59, 3, 68, 324, 86, 313, 336, 337, 339, 111, 63, 289, 348, 4, 
    57, 281, 67, 85, 94, 93, 98, 112, 101, 99, 105, 92, 72, 78, 94, 111, 124, 
    124, 117, 104, 104, 74, 76, 58, 75, 87, 82, 76, 81, 88, 63, 89, 310, 14, 
    334, 333, 350, 13, 134, 77, 322, 349, 0, 317, 332, 332, 329, 329, 322, 
    305, 311, 316, 360, 66, 73, 347, 356, 340, 312, 39, 79, 325, 2, 81, 319, 
    _, 73, 318, 335, 325, 344, 86, 309, 45, 95, 309, 304, 62, 308, 69, 306, 
    336, 91, 11, 15, 327, 350, 121, 338, 83, 95, 294, 318, 352, 319, 98, 75, 
    346, 344, 66, 326, 72, 23, 328, 102, 82, 92, 92, 78, 80, 86, 100, _, 95, 
    100, _, 102, 92, 89, 98, 91, 105, 99, 99, 96, 101, 110, 97, 98, 98, 95, 
    93, 93, 94, 88, 98, 101, _, 101, _, 87, _, 92, 101, 67, 94, 99, 98, 103, 
    127, 118, 100, 91, 90, 87, 101, 90, 75, 87, _, 83, 84, 296, 5, 313, 309, 
    309, 313, 101, 340, 112, 0, 310, 7, 0, 66, 61, 315, 322, 333, 4, 336, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 66, 326, 107, 324, 283, 282, 
    286, 85, 8, 84, 238, 271, 266, 265, 257, 259, 254, 251, 252, 258, 255, 
    245, 219, 224, 272, 262, 276, 281, 273, 276, 289, 274, 287, 300, 295, _, 
    _, 283, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, 314, 115, 318, 281, 7, 61, 329, 349, 318, 357, 
    _, 316, 329, 25, 0, 92, 76, 356, 331, 302, 350, 354, 75, 36, 38, 39, 26, 
    339, 42, 43, 26, 42, 46, 39, 91, 12, 25, 39, _, _, 22, 346, 52, 38, 23, 
    48, 59, 354, 18, 275, 288, 352, 53, 47, 355, 316, 352, 26, 15, _, 259, 
    26, 176, 49, 81, 278, 95, 72, 217, 338, 293, 327, 340, 352, 346, 329, 
    322, 337, 11, 335, 358, _, _, 343, 359, 309, 327, 110, 282, 57, 30, 81, 
    7, 359, 76, 318, 72, 296, 20, 333, 63, 14, 71, _, 294, _, 349, 297, 95, 
    311, _, _, 322, 97, _, _, _, 322, 81, 314, 81, 1, 301, 348, _, 82, 357, 
    _, 78, 103, 81, _, 312, 322, _, 298, 350, _, 321, _, 294, 275, 333, 304, 
    316, 49, 108, 74, 76, _, 65, 315, 305, _, 342, 18, 308, 354, 343, 49, 
    327, 321, 322, 328, 349, 15, 43, 301, 10, 357, 312, 21, 329, 357, 351, 
    102, 330, 81, 54, 339, 97, 345, 83, 22, 340, 93, 131, 17, 346, 340, 310, 
    5, 265, 321, 37, 174, 328, 293, 44, _, 335, 319, 305, 311, 294, 285, 297, 
    343, 302, 32, 266, 268, 260, 259, 252, 264, 263, 264, 272, 262, 262, _, 
    308, _, 314, 321, 223, 266, 308, 100, 331, 295, 328, 326, _, 314, _, 65, 
    15, 310, 296, 89, 106, 90, 327, 3, 0, 0, 107, 123, 276, _, 8, 0, 0, 0, 
    32, 93, 186, 314, 325, 325, 327, 321, 329, 115, 44, 32, 349, 319, 310, _, 
    50, 59, 12, 42, 44, 355, 15, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, 105, 61, 91, 92, 105, 75, 111, 101, 290, 
    112, 65, 105, _, _, _, 50, 36, _, _, _, 41, _, 39, _, 31, 38, 48, _, _, 
    37, 41, 33, 42, 37, 58, 58, 73, 15, _, 14, 2, 22, 14, 0, 8, 8, 7, 9, 12, 
    23, 18, 19, 18, 27, 31, 34, 37, 34, 32, 24, _, 14, 27, 38, 29, 13, 35, 
    35, 28, 34, 38, 29, 32, 32, 30, 30, 36, 38, 41, 31, 45, 53, 25, 44, _, 
    32, 25, 38, 59, 31, _, _, 69, 318, 318, 306, 343, 324, 326, 288, 81, 52, 
    357, 310, 294, 354, 56, 10, 358, 325, _, 328, 79, 331, 356, 95, 306, 88, 
    296, 138, 116, 322, 127, 64, 33, 324, 95, 91, 334, 107, 323, _, 43, 4, _, 
    21, 332, 75, 319, 94, 318, 226, 71, 119, 65, 47, 112, 111, 80, 68, 80, 
    100, 90, 83, 105, 97, _, 86, 92, 59, 77, 122, 92, _, 106, 93, 101, 109, 
    122, 121, 75, 90, 63, 102, 34, 340, 11, 20, 40, 359, 330, 14, _, 323, 63, 
    _, 306, 65, 299, 294, 313, 269, 303, 303, 65, 104, 0, 262, 28, 323, 65, 
    303, 27, _, 314, 328, _, 358, 84, 348, 116, 2, 103, 354, 45, 351, 77, 
    331, 106, 332, 141, 354, 322, 12, 341, 338, 328, 328, _, _, 340, 351, 
    320, 352, 353, _, 104, 124, 98, 118, 357, 322, 198, 28, 277, 34, 351, 1, 
    30, 27, 354, 321, 333, 31, 236, 263, 232, _, 235, 189, 270, 272, 194, 
    218, 58, 56, 148, 22, 44, 30, 50, 49, 50, 42, 350, 350, 2, 17, 17, 34, 
    356, 74, 308, 61, 353, 291, 25, 0, 156, 0, 325, 76, 20, 347, 89, 324, 
    291, 325, 307, 294, 92, 0, 354, 86, 288, 14, 349, 307, 1, 305, 313, 354, 
    69, 65, 52, 288, 277, 67, 57, 73, 71, 316, 70, 83, 95, 92, 90, 91, 78, 
    74, 48, 87, 102, 93, 87, 77, 79, 84, 17, 319, 11, 47, 299, 286, 283, 297, 
    290, 256, 274, 262, 271, 309, 316, 324, 51, 351, 314, 14, 304, 72, 74, 
    71, 311, 322, 81, 338, 36, 319, 70, 101, 84, 93, 95, 74, 82, 72, 117, 
    126, 150, 197, 340, 99, 127, 272, 312, 298, 252, 298, 297, 301, 287, 284, 
    269, 287, 283, 284, 269, 280, 266, 292, 305, 319, 313, 332, 303, 304, 
    101, 326, 271, 258, 304, 313, 71, 105, 96, 266, 304, 19, 308, 0, 0, 93, 
    0, 0, 317, 135, 338, 327, 261, 23, 24, 13, 257, 237, 49, 330, 274, 305, 
    121, 229, 54, 46, 222, 185, 339, 309, 220, 17, 2, 298, 320, 302, 100, 
    311, 330, 76, 2, 28, 69, 281, 5, 256, 62, 292, 98, 156, 122, 356, 272, 
    298, 347, 56, 303, 350, 334, 270, 79, 358, 295, 332, 40, 21, 331, 349, 
    268, 300, 286, 277, 279, 271, 39, 323, 69, 304, 335, 297, 286, 321, 110, 
    42, 43, 42, 42, 39, 21, 8, 21, 18, 18, 17, 25, 26, 34, 33, 27, 32, 30, 
    32, 27, 33, 23, 17, 23, 343, 351, 288, 244, 352, 336, 289, 68, 317, 286, 
    296, 294, 284, 68, 133, 329, 355, 98, 45, 72, 128, 85, 274, 273, 131, 49, 
    77, 132, 109, 281, 202, 255, 244, 238, 36, 65, 39, 21, 285, 9, 209, 11, 
    347, 17, 36, 125, 253, 286, 239, 306, 46, 64, 44, 6, 44, 12, 326, 212, 
    109, 14, 17, 54, 43, 14, 17, 24, 31, 307, 95, 82, 22, 25, 339, 344, 244, 
    90, 359, 3, 348, 49, 13, 8, 22, 226, 237, 49, 46, 326, 331, 116, 114, 
    102, 247, 35, 189, 206, 191, 221, 162, 39, 139, 213, 162, 33, 129, 307, 
    55, 330, 327, 307, 259, 276, 257, 298, 270, 276, 337, 345, 18, 338, 333, 
    100, 0, 2, 345, 247, 271, 128, 236, 268, 275, 278, 301, 276, 4, 341, 320, 
    120, 2, 0, 261, 232, 292, 231, 271, 267, 5, 297, 47, 313, 321, 309, 338, 
    358, 93, 317, 3, 324, 101, 41, 110, 105, 151, 22, 1, 233, 201, 117, 116, 
    333, 356, 236, 236, 220, 169, 157, 160, 167, 181, 53, 31, 359, 290, 134, 
    358, 312, 347, 291, 113, 16, 91, 17, 0, 250, 0, 359, 250, 248, 298, 258, 
    263, 345, 277, 275, 11, 302, 354, 93, 359, 117, 2, 128, 26, 137, 317, 
    346, 6, 180, 15, 273, 93, 1, 54, 306, 65, 128, 93, 73, 100, 105, 75, 107, 
    118, 89, 78, 119, 132, 98, 102, 78, 106, 124, 183, 218, 72, 72, 123, 108, 
    97, 332, 59, 296, 248, 308, 213, 254, 115, 56, 55, 240, 44, 57, 49, 20, 
    42, 13, 9, 58, 16, 18, 187, 165, 224, 221, 217, 265, 73, 358, 46, 318, 
    329, 42, 64, 88, 75, 97, 93, 28, 300, 339, 334, 310, 292, 18, 321, 311, 
    297, 300, 304, 303, 300, 315, 316, 298, 295, 294, 293, 288, 287, 289, 
    298, 267, 285, 289, 288, 294, 309, 303, 88, 310, 301, 134, 300, 228, 17, 
    155, 134, 264, 128, 177, 173, 139, 337, 5, 126, 66, 18, 40, 48, 50, 45, 
    40, 38, 90, 93, 103, 98, 94, 102, 284, 305, 95, 314, 294, 301, 304, 282, 
    285, 122, 116, 279, 311, 305, 303, 307, 304, 50, 91, 22, 356, 3, 100, 42, 
    269, 268, 270, 266, 239, 254, 242, 264, 268, 269, 271, 306, 280, 290, 
    289, 265, 282, 281, 285, 323, 296, 258, 233, 158, 140, 131, 171, 350, 
    298, 11, 283, 265, 359, 294, 283, 317, 123, 291, 275, 294, 293, 114, 120, 
    145, 17, 0, 150, 284, 3, 329, 317, 317, 316, 316, 343, 0, 89, 94, 37, 
    294, 304, 314, 316, 316, 260, 180, 358, 100, 104, 121, 106, 97, 82, 305, 
    289, 279, 295, 304, 304, 279, 271, 270, 277, 292, 278, 254, 259, 261, 
    179, 163, 116, 329, 114, 132, 153, 130, 127, 0, 358, 300, 301, 306, 316, 
    240, 58, 54, 46, 112, 344, 300, 285, 260, 272, 262, 256, 294, 283, 299, 
    270, 275, 2, 32, 119, 109, 113, 301, 296, 0, 0, 0, 350, 271, 274, 289, 
    287, 27, 18, 114, 264, 300, 276, 105, 331, 64, 6, 5, 59, 310, 99, 289, 
    202, 22, 77, 360, 283, 343, 214, 255, 2, 36, 212, 203, 181, 67, 121, 172, 
    21, 21, 328, 89, 25, 354, 2, 344, 6, 334, 353, 228, 328, 202, 221, 240, 
    263, 341, 258, 298, 282, 167, 215, 231, 326, 246, 339, 93, 36, 95, 31, 
    60, 67, 69, 51, 88, 43, 38, 24, 37, 43, 42, 60, 38, 59, 34, 244, 121, 39, 
    62, 31, 278, 254, 221, 213, 287, 129, 99, 124, 33, 53, 24, 17, 332, 308, 
    75, 3, 267, 217, 252, 126, 266, 261, 250, 260, 293, 47, 46, 42, 0, 0, 10, 
    203, 215, 209, 115, 185, 181, 162, 237, 210, 207, 338, 248, 306, 311, 
    347, 219, 30, 96, 80, 82, 99, 182, 133, 156, 262, 273, 216, 253, 240, 0, 
    271, 0, 64, 358, 49, 15, 337, 21, 264, 304, 341, 358, 278, 108, 106, 287, 
    331, 216, 239, 218, 131, 163, 205, _, _, _, _, _, _, 334, 288, 298, 302, 
    248, 296, 326, 272, 271, 280, 242, 272, 210, 251, 8, 23, 148, _, 131, 
    347, 5, 337, 96, 11, 340, 3, 357, 287, 332, 80, 116, _, 123, _, 112, 127, 
    84, 117, 111, 98, 96, _, 78, 87, 80, 59, 293, _, _, 15, 330, 65, _, 129, 
    122, 137, 128, 142, 244, 334, 153, _, 265, 204, 260, _, _, _, 358, 305, 
    286, 151, 249, 11, 300, 294, 340, 300, 252, 303, 268, 67, 84, 79, 73, 
    279, 285, 300, 310, 322, _, _, _, _, 307, 345, _, 349, _, _, 68, 55, _, 
    _, 124, 229, 102, 72, 73, 336, 192, 97, 187, _, _, 172, 346, 50, 82, 29, 
    _, 201, 261, 63, 56, 62, 5, 78, 89, 33, 3, 96, 7, _, _, 36, 53, 53, 57, 
    55, 159, 60, _, 190, 23, 45, 28, 287, 260, 59, 24, 57, 79, 64, 77, 46, 
    43, 23, 28, 15, 15, 356, 23, 26, 70, 45, 13, 115, 2, 12, 126, 94, 36, 81, 
    89, 111, 22, 54, 57, 71, 60, 88, 76, 76, 120, _, _, 336, 291, 18, 6, 297, 
    _, 312, 360, 87, 117, 5, 9, 19, 10, 91, 53, 72, 77, 75, 68, 48, 280, 26, 
    55, 51, 81, 175, 46, 24, 22, 39, 66, 6, 107, 96, 119, 184, 309, 157, 100, 
    70, _, 123, 198, 149, 256, 260, 262, 360, 82, 130, 356, 73, 98, 355, 351, 
    316, 283, 268, 85, 89, 132, 179, 207, 177, 171, 182, 154, 200, 272, 262, 
    252, 287, 314, 309, 309, 282, 283, 285, 299, 312, 299, 190, 164, 207, 
    153, 99, 103, 157, 168, 298, 280, 269, 294, 265, 150, 108, 128, 258, 139, 
    260, 190, 163, 144, 94, 98, 95, 93, 115, 105, 92, 90, 84, 95, 98, 116, 
    100, 86, _, 42, _, 70, 13, 6, 45, 17, 5, 346, 4, 7, 11, 29, 27, 14, 50, 
    12, 196, 79, 56, 67, _, 182, _, 51, 54, 208, 44, 11, 36, 360, 314, 174, 
    21, 360, 13, 152, 31, 30, 355, 64, 40, _, 134, _, 115, 83, 108, 87, 125, 
    359, 360, 355, 17, 351, 360, 43, 12, 194, 105, 7, 26, 23, 26, 14, 1, 16, 
    23, 354, 104, 118, 90, _, _, 64, 57, 191, 57, 65, 246, 211, 112, 60, 85, 
    104, 103, 212, 215, 177, 55, 26, 48, 49, 36, 111, _, 80, 64, 55, 59, 36, 
    97, _, 69, 82, 57, 69, 48, 64, 117, 108, 115, _, 96, 85, 85, _, 88, 94, 
    94, 114, 89, 98, 113, 68, 96, 107, 76, 93, 102, 91, 97, 99, 97, 92, 34, 
    129, 127, 188, 127, 173, 121, 109, 114, _, _, 333, 120, 120, 125, 99, 
    319, 273, 339, 163, 90, 355, 118, 205, 169, 232, 287, 202, 163, 119, 111, 
    102, 121, 136, 315, 312, 345, 307, 187, 127, 163, 335, 32, 252, 175, 132, 
    125, 131, 145, 158, 145, 90, 147, 134, 125, 132, 84, 50, 30, 53, 54, 248, 
    335, 6, 0, 26, 328, 333, 213, 99, 80, 86, 69, 91, 68, 213, 145, 152, 167, 
    180, 190, 210, 97, 73, 173, 317, 25, 147, 137, 179, 209, 161, 234, 190, 
    174, 161, 162, 151, 123, 165, 163, 159, 171, 168, 130, 134, _, 117, 104, 
    60, 110, 114, 109, 133, 124, 129, 136, 149, 143, 129, 158, 157, 156, 142, 
    162, 151, 153, 162, 113, _, _, 127, 128, 88, 151, 304, 66, 88, 79, 115, 
    145, 118, 114, 134, 136, 139, 129, 128, 129, 131, 174, 168, 137, 121, 66, 
    45, 58, 306, 311, 31, 40, 48, 55, 65, 69, 66, 118, 118, 104, 142, 156, 
    155, 147, 171, 173, 152, 172, 64, 72, 80, 166, 216, 183, 90, 102, 268, 
    182, 63, 73, 95, 155, 155, 159, 167, 69, 48, 181, 249, 272, 273, 287, _, 
    287, 295, 317, 295, 285, 333, 315, 305, 317, 300, 257, 332, 300, 282, 
    275, 188, 214, 233, 277, 273, 171, _, 172, 302, 298, 143, 126, 97, 89, 
    106, 125, _, 135, 152, 131, 166, 168, 169, 156, 167, 165, 161, 174, 170, 
    166, 158, 171, 138, 88, 115, 238, 314, 343, 120, 93, 46, 40, 146, 182, 
    175, 175, 258, 190, 181, 266, 272, 271, 196, 292, 279, 304, 307, 283, 
    266, 269, 296, 282, 282, 284, 271, 265, 341, 267, 295, 341, 159, 174, _, 
    197, 175, 170, 169, 157, 110, 121, 135, 99, 66, 65, 62, 57, 66, 50, 38, 
    67, 94, 120, 101, 124, 125, 123, 124, 123, 129, 103, 109, 111, 95, 95, 
    102, 135, 118, 115, 120, 126, 135, 315, 295, 296, 272, 276, 293, 239, 
    241, 15, 16, 53, 358, 10, 345, 66, 6, 93, 69, 164, 128, 92, 197, 31, 76, 
    222, 119, 51, 176, 159, 67, 260, 70, 66, 153, 246, 184, 87, 137, 143, 
    134, 171, 95, 21, 297, 308, 319, 323, 331, 328, 270, 293, 260, 291, 277, 
    263, 282, 268, 282, 271, 268, 269, 256, 280, 269, 261, 291, 290, 294, 
    275, 267, 249, 283, 288, 285, 285, 273, 263, 268, 265, 251, 248, 282, 
    272, 280, 288, 292, 281, 276, 339, 75, _, 325, 317, 350, 217, 104, 82, 5, 
    56, 2, 31, 57, 50, 81, 60, 54, 37, 36, 297, 63, 87, 81, 212, 80, 27, 266, 
    146, 358, 0, 334, 352, _, 84, 67, 81, 71, 69, 82, 73, 61, 60, 126, 78, 
    84, 84, 209, 115, 153, 182, 174, 160, 313, 290, 264, 283, 127, 99, 125, 
    120, 113, 126, 152, 144, 137, 136, 162, 170, 159, 126, 180, 163, 122, _, 
    107, 85, 108, 101, 79, 63, 109, 124, 138, 152, 170, 157, 168, 125, 137, 
    124, 67, 76, 52, 64, 54, 67, 212, 217, 247, 77, 6, 87, 85, 8, 212, 30, 
    346, 35, 77, 46, 65, 68, 61, 19, 360, _, 12, 341, 240, 23, 36, 48, 75, 
    64, 202, 75, 62, 47, 77, 132, 103, 54, 47, 52, 92, 132, 108, 100, 103, 
    96, 80, 57, 93, 107, _, _, 70, 329, 95, 342, 243, 174, 263, 171, 285, 
    233, 228, 127, 233, 161, 127, 184, 230, 162, 115, 185, 189, 186, 184, 
    337, 170, 159, 136, 31, 162, 360, 329, 159, 352, 292, 267, 316, 243, 176, 
    163, 152, 180, 170, 172, 268, 242, 255, 127, 353, 37, 53, 0, 0, 349, 68, 
    _, 120, 89, 117, 120, 129, 125, 139, 138, 130, _, 132, 121, 128, 109, 
    119, 128, _, _, 171, 33, 142, 71, 69, 151, 160, 327, 135, 130, 155, 135, 
    119, 121, 140, 136, 133, 134, 120, 127, 139, _, 159, 158, 89, 151, 133, 
    140, 126, 138, 172, 190, 165, 152, 99, 138, 126, 135, 122, 111, 124, 133, 
    137, 121, 123, 124, 128, 272, 296, 0, 13, 343, 251, 258, 249, 73, 61, 88, 
    96, 116, 274, 118, 35, _, 82, 114, 205, 163, 190, 233, _, 262, 286, 239, 
    154, 59, 73, 332, 308, 135, 130, 179, 75, 78, _, 157, 80, 86, 359, 72, 
    92, 66, _, 41, 63, 53, 43, 58, 159, 126, 74, 134, 104, 228, 69, 358, 343, 
    337, 96, 280, 9, 310, 55, 16, 157, 44, 54, 355, 287, 210, 223, 287, 168, 
    160, 194, 223, 250, 298, 5, 240, 150, 193, 65, 35, 220, _, 179, 171, 297, 
    243, 205, 277, _, 178, 260, 267, 195, 242, 324, 75, 93, 269, 120, 124, 
    101, 108, _, 81, 102, 97, 87, _, 62, 50, 96, 217, 57, 76, 62, 81, 75, 70, 
    100, 104, 126, 119, 94, 91, 141, 119, 105, 112, 108, 98, 89, 72, 63, 70, 
    67, 75, 90, 75, 115, 22, 83, 100, 64, 34, 349, 110, 124, 137, 107, 158, 
    130, 134, 137, _, 128, 128, 133, 122, 113, 129, _, 0, 351, 83, 0, 93, 
    112, 131, 108, 107, 123, 296, 198, 80, _, 151, 122, 80, 103, 96, 137, 
    318, _, 186, 228, 177, 323, 312, 194, 4, 338, 8, 13, 294, 128, 106, 141, 
    81, 66, 91, 79, 64, 69, _, 147, 27, 348, 61, 53, 329, 41, 348, 34, 36, 
    46, 46, 57, 28, 18, 67, 35, 73, 63, 53, 331, 320, 313, 38, 79, 91, 184, 
    125, 67, 360, _, 20, 180, 81, 76, 75, 64, 10, 181, 194, 119, 12, _, 112, 
    84, 69, 73, 69, 33, 16, _, 355, 277, 0, 288, 104, 167, 127, 32, 0, 98, 
    111, 78, 156, 172, 173, 167, 184, _, 165, 199, 285, 186, 282, 290, 273, 
    276, 279, 282, 293, 291, 20, 310, 169, 272, 170, 175, 251, 301, 305, 180, 
    173, 166, _, 173, 172, 127, _, 127, 137, 174, 117, 122, 106, 212, 53, 
    140, 133, 23, 79, 94, 39, 68, 82, _, 113, 109, 151, 138, 154, 141, 158, 
    _, 120, 140, 162, 271, 356, 145, 254, 130, 104, 108, 101, 95, 103, 99, 
    115, 112, 108, 109, 117, _, 115, 92, 183, 98, 116, 88, 89, 92, 103, 96, 
    90, 58, 359, 108, 29, 14, 307, 156, 164, 157, 73, 142, _, 139, 87, 129, 
    _, 143, 13, 356, 6, 128, 342, 352, 36, 310, 360, 108, 287, 5, 260, 52, 
    137, _, 134, 140, 171, 149, 129, 105, 81, _, _, 79, 109, 349, 85, 324, 
    273, 335, 320, 12, 110, 136, 97, 112, 85, 132, 123, 87, 85, 84, _, _, 
    102, 97, 74, 66, 78, 97, 333, 308, 325, 1, 325, 324, 325, 125, 109, 117, 
    75, 102, 87, 92, _, _, 88, 98, 101, 127, 106, 269, 126, _, 82, 105, 89, 
    295, 305, 314, 145, 26, 102, 129, 231, 127, 130, 90, 83, 101, 162, 169, 
    100, 106, 133, 20, 4, 299, 333, 327, 338, 96, 336, 130, 136, 269, 143, 
    147, 124, 140, 148, 145, 162, 111, _, _, 76, 114, 136, 109, 116, 128, 
    106, 116, 52, 119, 123, 116, 129, 117, 132, 120, 126, 134, 128, 130, _, 
    126, 130, 283, _, 148, 117, 300, 300, 276, 102, 0, 0, 0, 0, 110, 282, 
    315, 112, 338, 326, 159, 65, 113, 121, 148, 94, 113, 78, 90, _, 300, 306, 
    305, 298, 296, 321, 98, 115, 84, 118, 134, 130, 145, 115, 126, 155, 146, 
    144, 156, _, _, 109, 93, 112, 127, 254, 131, 87, 105, 107, 104, 172, 171, 
    163, 92, 179, 171, 166, 170, 176, 178, _, 90, 85, 88, 93, 106, 131, 113, 
    123, 110, 124, 114, 193, 159, 119, 106, 138, 125, 139, 127, 131, 138, 
    143, _, 151, 130, 136, 145, 103, 131, _, 203, 96, 84, 69, 93, 109, 88, 
    89, 115, 95, 93, 96, 94, 108, 137, 120, 110, 99, 104, _, _, 127, 120, 16, 
    48, 120, 102, 142, 335, 297, 289, 120, 119, 139, 158, 269, 135, 122, 126, 
    101, 113, 127, 119, 111, 112, 117, 77, 77, 317, 28, 93, 72, 203, 73, 17, 
    95, 263, 132, 150, 105, 165, 138, 0, 264, 247, 246, 285, 85, 94, 110, 99, 
    106, 112, 70, 125, 56, 0, 31, 81, 110, 353, 342, 124, 89, 132, 126, 131, 
    111, 102, 128, 125, 87, 49, 11, 2, 180, 206, 213, 172, 340, 321, 10, 340, 
    286, 284, 34, 149, 137, 267, 194, 244, 193, 219, 227, 217, 206, 196, 198, 
    307, 283, 300, 321, 331, 327, 315, 355, 321, 78, 353, 350, 278, 323, 104, 
    150, 163, 160, 169, 144, 131, 152, 140, 151, 171, 166, 94, 85, 98, 84, 
    95, 135, 164, 157, 173, 163, 24, 159, 110, 166, 168, 167, 157, 114, 125, 
    121, 117, 108, 100, 121, 114, 0, 266, 111, 185, 241, 0, 4, 145, 127, 129, 
    124, 132, 124, 147, 156, 2, 202, 275, 347, 349, 294, 317, 0, 355, 0, 110, 
    70, 96, 341, 9, 357, 0, 291, 359, 334, 68, 36, 97, 104, 121, 138, 121, 
    359, 50, 114, 126, 122, 22, 354, 314, 274, 268, 252, 280, 300, 324, 197, 
    282, 294, 308, 269, 269, 265, 278, 267, 282, 277, 283, 297, 295, 276, 
    281, 281, 245, 298, 283, 294, 241, 304, 226, 271, 268, 271, 279, 274, 
    272, 280, 282, 272, 261, 251, 268, 275, 293, 286, 295, 280, 315, 292, 
    312, 313, 310, 309, 322, 204, 265, 302, 285, 285, 288, 287, 282, 287, 
    105, 121, 134, 95, 81, 105, 326, 336, 323, 309, 318, 333, 10, 305, 353, 
    8, 250, 73, 104, 120, 114, 108, 130, 110, 88, 147, 122, 90, 72, 51, 62, 
    266, 195, 0, 335, 319, 41, 34, 27, 20, 54, 13, 214, 198, 142, 104, 120, 
    116, 111, 107, 100, 101, 106, 98, 85, 89, 67, 77, 92, 177, 72, 61, 73, 
    76, 84, 93, 62, 60, 82, 229, 303, 291, 149, 111, 99, 138, 133, 124, 117, 
    58, 111, 93, 89, 0, 321, 0, 114, 108, 113, 360, 136, 119, 0, 134, 125, 
    124, 126, 38, 359, 73, 183, 186, 337, 334, 315, 47, 175, 358, 292, 355, 
    95, 107, 4, 102, 102, 121, 130, 122, 114, 150, 143, 138, 132, 127, 288, 
    314, 322, 153, 308, 234, 11, 307, 0, 3, 331, 339, 334, 227, 2, 128, 130, 
    133, 105, 111, 102, 115, 107, 126, 122, 123, 117, 316, 352, 27, 352, 72, 
    119, 116, 113, 112, 97, 121, 126, 77, 27, 108, 126, 115, 173, 155, 151, 
    289, 312, 303, 326, 317, 0, 320, 307, 309, 347, 346, 0, 343, 330, 85, 
    134, 98, 111, 121, 116, 107, 105, 101, 106, 105, 105, 93, 100, 96, 3, 37, 
    341, 328, 298, 288, 300, 294, 296, 0, 0, 0, 0, 316, 358, 6, 315, 358, 30, 
    25, 40, 47, 58, 23, 19, 200, 51, 38, 31, 44, 37, 37, 54, 47, 61, 100, 
    112, 91, 106, 119, 100, 109, 107, 96, 121, 130, 126, 128, 125, 88, 71, 
    76, 74, 51, 29, 82, 33, 34, 37, 43, 70, 97, 118, 84, _, _, 11, 355, 13, 
    14, 12, 39, 29, 19, 280, 30, 36, 44, 35, 28, 26, 23, _, 38, 55, 39, 51, 
    61, 62, 51, 28, 39, 60, 50, 26, 89, 110, 57, 25, 168, 302, 302, 283, 292, 
    250, 186, 294, 280, 349, 345, 83, 268, 70, 33, 313, 310, 296, 325, 317, 
    347, 155, 125, 308, 275, 350, 52, 334, 196, 202, 272, _, 2, 346, 15, 19, 
    15, _, _, 27, 35, 16, 215, 339, 61, 347, 29, 46, 211, 161, 211, 283, 333, 
    352, 329, 356, 311, 0, 63, 58, 60, 89, 225, 149, 128, 14, 62, 46, 351, 
    52, 39, 42, 21, 350, 29, 314, 317, 295, 307, 299, 353, 171, 347, 260, 
    118, 111, 105, 0, 1, 34, 0, 0, 318, 0, 0, 314, 312, 341, 0, 0, 318, 353, 
    274, _, 283, 130, 132, 156, 27, 0, 118, 103, 193, 108, 3, 321, 321, 246, 
    303, 0, 309, 0, 22, 330, 7, 344, 338, 10, 75, _, 63, 62, 69, 62, 320, 
    298, 283, 270, 277, 273, 289, 267, 271, 286, 285, 289, 303, 299, 312, 
    286, 280, 274, 269, 269, 272, 274, 270, 288, 275, 276, 290, 287, 301, 
    308, 309, 297, 272, 323, 328, 316, 292, 307, 300, 309, 303, _, 279, 264, 
    260, 228, 219, 283, 294, 302, 302, 355, 310, _, 297, 219, 305, 360, 323, 
    312, 279, 289, _, 310, 91, 55, 79, _, 28, _, _, 89, 10, 62, 298, 296, 
    301, 284, 281, 308, 342, 345, 1, 0, 0, 0, 0, 0, 0, 0, 327, 332, 0, 354, 
    80, 26, 313, 321, 317, 285, 307, 290, 292, 294, 276, 294, 287, 303, 283, 
    299, 292, 287, 302, _, 268, 269, 279, 263, 284, 287, _, 301, 125, 0, 0, 
    333, 334, 341, 21, 18, 297, 314, 308, 278, _, 304, 305, 290, 317, _, 304, 
    310, 275, 332, 340, 306, 313, 305, 71, 138, 324, 274, 296, 34, 291, 49, 
    336, 334, 61, 0, 291, 34, 299, 335, 356, 0, 112, 13, 358, 356, 354, 309, 
    100, 0, 284, 75, 82, 118, 360, 291, 359, 36, 330, 56, 45, _, 149, 97, 
    247, 326, 355, 58, _, 313, 310, 299, 0, 331, 96, 87, 55, 303, 333, 3, 0, 
    341, _, 307, 358, 340, 0, 352, 320, 295, _, 282, 295, 311, 311, 339, 0, 
    9, 355, 326, 343, 101, 124, 306, 333, 329, 325, 91, _, 352, 242, _, 145, 
    95, 45, 222, 357, 39, 67, 74, 100, 358, 329, 321, 293, 353, 324, 27, 301, 
    306, 6, 339, 45, _, 264, 66, 232, 154, 335, 278, _, 350, 347, 0, 0, 347, 
    54, 351, 38, 328, 35, 1, 9, 8, _, 300, 294, 176, 88, 97, 321, 294, _, _, 
    315, 303, 322, 313, 319, 340, 310, 355, 37, 320, 0, 0, 340, 0, 310, 29, 
    337, 285, 290, 266, 309, 14, 68, 75, 64, 352, 296, 325, 306, 313, 287, 
    305, 309, 319, 52, 338, 356, 346, 0, 337, 360, _, 8, 335, 299, 288, 303, 
    282, 285, 293, 14, 66, 14, 112, 0, 304, 39, 355, 328, 304, 284, 306, 61, 
    344, 351, 101, 349, 300, 307, 348, _, 347, 290, 296, 107, 251, 119, 358, 
    331, 337, 95, 355, 341, 309, 89, 60, 0, 334, 110, 0, 310, 103, _, 113, 
    318, 358, 10, 360, 353, 334, 40, 339, 345, 323, 358, 344, 356, 353, 325, 
    332, 359, 32, 2, _, 0, 103, 255, _, 53, 323, 33, 77, _, 309, 345, 13, 0, 
    0, 337, 325, 359, 0, 16, 1, _, 313, 337, 334, 325, 324, 0, 0, _, _, 344, 
    337, 8, 359, 45, 52, 9, 7, 0, 40, 9, 57, 5, 332, 356, 105, 43, 278, 17, 
    _, _, 339, 202, 322, 20, 44, 6, 353, 354, 331, 317, 9, 2, 322, 0, 0, 351, 
    53, 0, 0, 0, _, 0, 0, 0, 353, 329, 323, 331, 0, _, 24, 10, 6, _, 343, 
    335, 310, 303, 292, 323, 83, _, 136, 90, 341, 331, 341, 137, 337, 355, 
    346, 0, 322, 322, 276, 217, 94, 351, 322, 350, 81, 334, 323, 74, 318, 
    298, 357, 331, 320, 342, _, 316, 23, 72, 71, 59, 50, 51, 32, 38, _, 8, 
    17, 20, 10, 6, 273, 282, 289, 303, 321, 322, _, _, 333, 324, 299, 289, 
    295, 312, 289, _, 287, 278, 291, 316, 306, 293, 338, 326, 314, 306, 301, 
    _, 325, 325, 312, 310, 306, 286, 280, 278, _, 279, 284, 271, 303, 332, 0, 
    19, 220, 347, 1, 25, 357, 23, 351, 98, 119, 69, 81, 257, _, 260, 2, 105, 
    83, 312, 310, 313, 343, 320, 0, 331, 0, 337, 347, 355, 0, 330, 319, 323, 
    344, 294, _, _, 287, 70, 344, 309, 306, 290, 3, 351, 353, 332, 325, 339, 
    312, 353, 42, 313, 1, 301, 298, 334, 331, 93, 333, 315, 155, 98, 290, 
    289, _, 309, 18, 325, 328, 322, 328, 360, 303, 308, 336, 334, 322, 345, 
    312, 314, 329, 342, 313, 343, _, 345, 357, 344, 359, 320, 0, 352, 303, 
    302, 300, 307, 336, 273, 294, 320, 334, 287, 292, 328, 338, 348, _, _, 
    334, 19, 0, 291, 0, 0, 311, 317, 310, 352, 20, 38, 332, 320, 0, 314, 75, 
    331, 358, 32, 347, 309, 310, 327, 41, 34, 335, 25, _, 325, 310, 302, 82, 
    325, 337, 334, 0, 309, 0, 44, 6, 10, 359, 327, 59, 0, 0, 34, _, 339, 54, 
    336, 350, 337, 295, 66, 7, 26, 0, 0, 17, 0, 338, 15, 0, 0, 340, 344, 81, 
    352, _, _, 352, 11, 356, 358, 336, 318, 2, 312, 315, 305, 35, 37, 329, 
    27, 35, 304, 13, 324, 357, 309, 76, 311, 334, 48, 14, 71, 17, 348, _, 
    305, 66, 75, 334, 336, 70, 307, 354, 315, 326, 333, 70, 339, 314, 84, 9, 
    337, 352, 44, _, 360, 355, 13, 357, 14, 8, 24, 79, 335, 327, 334, 282, 
    343, 97, 312, 345, 299, 1, 80, 338, 290, _, _, 0, 32, 0, 317, 27, 6, 337, 
    311, 326, 0, 321, 0, 284, 6, 0, 318, 323, 309, 2, 357, 60, 79, 342, 346, 
    0, 324, 0, 0, 327, 305, 331, 313, 324, 53, 316, 325, 0, 305, 347, 64, 
    304, 333, _, 24, 339, 304, 302, 325, 92, 62, 93, 91, 84, 99, 142, 94, 78, 
    78, 85, 61, 316, 316, 305, 353, 334, 304, 64, 54, 329, 359, _, _, 0, 342, 
    9, 339, 328, 331, 0, 344, 54, 19, 5, 0, 0, 334, 293, 291, 295, 297, 293, 
    302, 302, 294, 294, 304, 300, 304, 300, 288, 287, 301, 314, 304, 322, 
    343, 354, 354, 18, 51, 21, 353, 349, 36, 16, 342, 313, 341, 56, 336, 320, 
    323, 308, 312, 305, 340, 333, 2, 344, 360, 6, 314, 359, 299, 35, 319, 
    322, 338, 283, 91, 321, 319, _, _, 310, 300, 309, 301, 312, 9, 311, 287, 
    286, 298, 85, 0, 325, 314, 301, 88, 0, 0, 0, 0, 283, 299, 78, 77, _, 253, 
    261, 271, 264, 255, 292, 307, 312, 77, 58, 38, 33, 33, 34, 35, 34, 36, _, 
    39, 33, 32, 38, 42, 50, 43, 17, 38, 44, 42, 48, 49, 50, 46, 69, _, 65, 
    60, 66, 78, 67, 62, 63, 60, 103, 82, 56, _, 73, 62, 75, 81, 81, 91, 100, 
    74, 84, 87, 89, 79, 84, 73, 76, 90, 92, 95, 98, 93, _, 83, 101, 98, 96, 
    93, 90, 95, 90, 95, 97, 99, 86, 109, 96, 91, 89, 101, 99, 95, 93, 103, _, 
    95, 94, 106, 103, 92, 99, 81, 93, 100, 97, 88, 78, 84, 80, 83, 84, 86, 
    100, 100, 80, 92, 74, 51, 343, 74, 33, 338, 331, _, _, 301, 6, 315, 335, 
    36, 41, 39, 36, 34, 31, 50, 45, 18, 21, 25, 350, 16, 77, 354, 4, 1, 50, 
    26, 196, 346, 59, 66, 70, 80, 80, 62, 68, 65, 64, 4, 6, 8, 11, 7, 356, 
    308, 1, 9, 5, 2, 202, 267, 208, 5, 34, 31, 29, 23, 15, 20, 331, 24, 333, 
    185, 352, 335, 346, 335, 313, 300, 313, 317, 294, 354, 349, _, 305, 327, 
    316, 322, 329, 330, 330, 342, 21, 27, 347, 344, 325, 352, 337, 322, 317, 
    293, 306, 280, 309, 347, 329, 311, 300, 304, 309, 299, 290, 297, 307, 
    314, 297, 296, 322, 349, 315, 354, 300, 304, 314, 306, 288, 311, 293, 
    312, 315, 314, 331, 356, 313, 0, 299, 359, 355, 304, 326, 0, 310, 291, 
    297, 292, 305, 69, 93, 94, 88, 58, 354, 0, 0, _, _, 302, 320, 318, 312, 
    310, 314, 311, 312, 312, 316, 304, 311, 302, 307, 324, 315, 304, 313, _, 
    317, 317, 300, 298, 301, 311, 302, 304, 264, 77, 55, 315, 252, 313, 167, 
    333, 31, 159, 3, 246, 294, 312, 111, 16, 274, 353, 32, 4, 49, 326, 65, 
    22, 7, 335, 327, 61, 8, 31, 0, 0, 355, 341, 0, 15, 23, 335, 10, 0, 357, 
    10, 12, 351, 0, 349, 345, 353, 315, 180, 20, 19, 27, 36, 38, 33, 37, 34, 
    44, 41, 38, 45, 42, _, 31, 35, 49, 62, 355, 110, 78, 8, 24, 351, 26, 33, 
    358, 24, 356, 303, 310, 4, 338, 344, 325, 2, 50, _, 271, _, 353, 330, 
    348, 336, 328, 326, 303, 248, 42, 46, 38, 33, 41, _, 176, 43, 216, 265, 
    303, _, 273, 288, 307, 315, 310, 295, _, 286, 321, 308, 309, 314, 308, 
    307, 308, 309, 320, 314, 309, 354, 327, 313, 344, 308, 314, _, 310, 329, 
    329, 301, 284, 338, 288, 23, 319, 319, 309, 304, 299, 320, 353, 319, 313, 
    354, 306, 336, 290, 266, 307, _, 333, 292, 339, 328, 302, 324, 328, 316, 
    336, 1, 6, 341, 286, 24, 312, 337, 315, 14, 332, 313, 346, _, 95, 311, 
    294, 329, 313, 342, _, 303, 325, 356, 84, 301, 305, 314, 307, 214, 95, 
    32, 350, 354, _, 1, 281, 353, 302, 322, 317, 319, 312, 317, 14, 305, 1, 
    323, 46, 80, 323, 310, 2, 329, 326, 295, 357, 322, 325, 338, 89, 75, 88, 
    81, 103, 86, 93, 91, 91, 103, 85, 91, 100, 95, 75, 79, 85, 94, 92, 85, 
    80, 87, 83, 88, 80, _, 68, 57, 102, 103, 352, 73, _, 89, 59, 121, 102, 
    91, 99, 95, 119, 78, 104, 133, 121, 112, 184, 45, 110, 131, 117, 111, 
    116, 95, _, 131, 137, 106, 148, 90, 95, 115, 133, 117, 131, 119, 105, 78, 
    96, 67, 64, 61, 109, 117, 117, 91, 84, 79, 70, 63, 79, 63, 64, 82, 78, 
    81, 85, 76, 84, 102, 107, 97, 96, 87, 93, 88, 80, _, _, 77, 93, 83, 104, 
    103, _, 95, 77, 72, 73, 71, 80, 73, 90, 68, 85, 74, 93, 67, 54, 52, 58, 
    44, 38, 50, 47, 43, _, _, 56, 22, 36, 35, 41, 21, 35, 82, 69, 74, 69, _, 
    74, 64, 88, 82, 84, 73, 72, 63, _, 75, 57, 57, 59, 79, 80, 3, 193, 334, 
    39, 349, 27, 1, 335, 0, 315, 339, 313, 319, 301, _, _, 293, 326, 323, 
    328, 296, _, 314, 335, 360, 323, 57, 356, 350, 0, 356, 35, 48, 41, 42, _, 
    41, 50, 35, 24, 37, 30, 30, _, 23, 325, 292, 356, 25, 35, 35, 33, 52, 
    340, 28, 99, 62, 118, 52, 95, 105, 119, 83, 104, _, 90, 54, 41, 42, 59, 
    318, 296, 188, 293, 36, 128, 254, 285, 206, 312, 168, 320, 310, 320, 293, 
    277, _, 222, 290, 250, 311, 335, 328, 340, 315, _, 299, 340, 315, 313, 
    305, 308, 355, 339, 304, 319, 326, 307, 317, 311, 293, 297, 301, 304, 
    306, _, 346, 327, 314, 357, 337, 319, 310, 287, 313, 314, 315, 301, 351, 
    355, 0, 293, 289, 272, 311, 294, _, 350, 18, 13, 24, 312, 38, 297, 321, 
    295, 318, 294, 296, 291, 310, 316, 318, 296, 299, 291, 286, 296, _, _, 
    305, 302, 292, 317, 354, 1, 357, 128, 339, 53, 27, _, 302, 277, 267, 229, 
    271, 279, 309, _, 188, 282, 282, 290, 252, 325, 301, _, 244, 257, 92, 
    291, 3, 60, 246, 228, 263, 107, 196, 262, 54, 86, 201, 76, 158, 178, 304, 
    354, 344, 282, 357, 349, 59, 314, 277, 274, 66, 66, 65, 60, 66, 66, 67, 
    74, 75, 64, 79, 82, 79, 321, _, 353, _, 29, 57, 69, 66, 76, 70, _, 81, 
    86, 76, 85, 78, 97, 92, 96, 95, 93, 80, _, 61, 69, 65, 56, 76, 87, 83, 
    26, _, 48, 47, 77, 81, 83, 102, 118, 90, 84, 81, 73, 77, 77, 50, 82, 79, 
    80, 86, 98, 88, _, 86, 78, 63, 74, 72, 64, 59, 64, 79, 69, 72, 85, 79, 
    87, 68, 60, 70, 73, 75, 77, _, _, _, 116, 88, 85, 105, 90, 95, _, 60, 32, 
    37, 18, 28, 48, 39, 32, 33, 18, 40, _, 118, 48, 31, 52, 51, 45, 47, 53, 
    _, 46, 58, _, 39, 77, _, 92, 95, 91, 104, 93, 91, 93, 89, 97, 98, 95, 98, 
    96, 100, 89, 93, 96, 71, 74, 72, 59, 141, 83, 345, 84, 60, 71, 82, 292, 
    293, 315, 306, 312, 317, 310, _, _, 346, 333, 92, 311, 345, 328, 46, 292, 
    306, 34, 301, 315, 12, 336, 299, 316, 323, 329, 13, _, 71, 80, 76, 281, 
    35, 40, 41, 304, _, 332, 355, 352, 99, 4, 319, 15, 339, 215, 281, 328, 6, 
    29, 72, 200, 222, 298, 33, 43, 121, 285, _, 30, 32, 34, 33, 37, 17, 11, 
    10, 220, 289, _, 188, 356, 5, 266, 16, 329, 267, 9, _, _, 296, 1, 278, 
    311, 166, 126, 204, 36, 70, 141, 114, 95, 100, 93, 97, 89, 89, 95, 76, _, 
    64, 84, 80, 72, 62, 60, 63, 65, _, 47, 68, 34, 15, 44, 48, 55, 42, 52, 
    47, 61, 57, 45, 60, 63, 51, 55, 302, 350, 338, 352, 31, 326, 307, 303, 
    23, 327, 350, 330, 324, 336, 356, 13, 317, 310, 278, 252, 291, 329, 283, 
    326, _, _, 309, 316, 315, 328, 324, 328, 324, 303, 349, 302, 339, 331, 
    308, 328, 335, 320, 309, 318, 330, 278, 315, 317, 320, 313, 339, 22, 34, 
    21, 45, 55, 341, 360, 26, 302, 304, 322, 335, 317, 289, 323, 332, 300, 
    312, 327, 312, 327, 304, 301, 310, 310, 313, 322, 323, 341, 347, 6, 323, 
    60, 308, 282, 287, 296, 306, 284, 297, 298, 284, 290, 300, 295, _, _, 
    303, 22, 355, 310, 302, 314, 1, 40, 34, 44, 47, 41, 43, 39, 41, 39, 43, 
    41, 45, 51, 54, 242, 226, 349, 216, 142, 352, 236, 343, 289, 318, 253, 
    173, 258, 142, 153, 43, 272, 332, 93, 281, 320, 298, 310, 297, 275, 301, 
    292, 324, 310, 322, 308, 292, _, 306, 297, 335, 254, 358, 298, 319, 313, 
    320, 321, 326, 314, 312, 314, 330, 324, _, _, 323, _, 29, 14, 321, 323, 
    358, 52, 3, 65, 97, 54, 66, 5, 16, 42, 350, 11, 8, 58, 22, 358, 325, 337, 
    319, 5, 334, 3, 337, 4, 338, 343, 37, 360, 6, 0, 324, 320, 202, 295, 146, 
    32, _, 45, 39, 21, 356, 6, 47, 338, 335, 37, 308, 12, 342, 311, 357, 322, 
    315, 318, 311, 316, 292, 326, 318, 302, 326, 323, 335, 306, 288, _, 107, 
    57, 90, 67, 353, 305, 282, 273, 327, 113, 88, 99, 93, 110, 97, 95, 102, 
    93, 97, 95, 100, 92, 95, 95, 93, 91, 91, 96, 94, 93, 95, 95, 96, 98, 95, 
    92, 91, 90, 92, 89, 92, 92, 93, 97, 96, 95, 94, 94, 93, 89, 87, _, 88, 
    98, 97, 134, 118, 88, 87, 94, 94, 88, 88, 93, 85, 96, 101, 93, 84, 93, 
    97, _, 89, 69, 88, 90, 83, 75, 88, 73, 86, 73, 70, 89, 79, 73, 68, 76, 
    47, 32, 80, 78, 40, 41, 57, 50, 327, 320, 314, 47, 352, 335, 321, 295, 
    13, 328, 335, 317, 326, 8, 326, 54, 296, 355, 233, 319, 331, 279, 297, 1, 
    53, 37, 64, 49, 302, 306, 337, 61, 322, 304, 329, 316, 307, 314, 321, 
    312, 332, 20, 331, 303, 298, 100, 67, _, 40, 69, 74, 83, 74, 66, 64, 65, 
    310, 311, 294, 296, 284, 305, 295, 306, 300, 297, 309, _, 278, 76, 316, 
    337, 350, 315, 0, 0, 17, 328, 354, 358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 38, 
    17, 39, 41, 34, 28, 32, 15, 20, 11, 8, 12, 14, 14, 14, 29, 25, 28, 27, 
    33, 19, 15, 13, 18, 24, 25, 13, 12, 4, _, 319, 294, 296, 291, 304, 288, 
    304, 299, 289, 294, 298, 294, 297, 305, 304, 296, 298, 304, 311, _, 333, 
    333, 296, 311, 315, 312, 304, 305, 329, 308, 290, 304, 325, 322, 307, 
    305, 331, 309, 295, 305, 284, 288, 290, _, 305, 297, 306, 317, 329, 324, 
    339, 320, 326, 12, 253, 292, 304, 294, 288, 313, 94, 292, 312, 49, 95, 
    341, 301, 299, 281, 292, 316, 96, _, 333, 1, 358, 9, 5, 313, 312, 346, 
    343, 333, 302, 220, 52, 285, 290, 269, 291, 143, _, 351, 276, 20, 314, 
    323, 321, 267, 317, 322, 303, 302, 118, 73, 309, 358, 317, 313, 39, 5, 
    304, 296, 345, 315, 336, 11, 319, 1, 304, 359, 36, 72, 182, 21, 296, 281, 
    298, 314, 311, 107, 300, 289, 277, 272, 296, 297, _, 270, 284, 258, 296, 
    83, 359, _, 12, 340, 358, 15, 347, 331, 2, 85, 75, 313, 308, 308, 321, 
    39, 30, 217, 284, 317, _, 224, 329, 77, 314, 358, 332, 351, 318, 284, 
    311, 316, 317, 305, 76, 312, 312, 323, 318, 264, 266, _, 269, _, _, 30, 
    86, 220, 333, 287, 301, 237, 238, 211, 199, 226, 261, 324, 232, 249, 270, 
    267, 240, 237, 267, 281, _, 296, 313, 314, 298, 287, 279, _, 297, 299, 
    297, 299, 322, 311, 310, 315, 352, 297, 314, 313, 267, 295, 303, 309, 
    287, 274, 303, 343, 316, _, 314, 322, 306, 323, 327, 301, 310, 288, 302, 
    293, 314, 305, 297, 299, 294, 315, 339, 314, 294, _, _, 282, 297, 301, 
    294, 276, 301, 330, 293, 279, 310, 306, 300, 300, 316, 358, 320, 326, 
    333, 314, 290, 294, _, 293, 38, 327, 71, 86, 355, _, 34, 84, 92, 77, 53, 
    45, 48, 44, 43, 34, 12, 38, 48, 38, 19, 40, 49, 29, 34, 299, 321, 328, 
    333, 302, 79, 94, 87, 74, 72, 74, 81, 83, 95, 96, 104, 103, 111, 106, 73, 
    84, 84, 70, 73, 75, 78, 80, 83, 64, 62, 293, 309, 315, 302, 287, 76, 90, 
    75, 68, 71, 221, 68, 80, 68, 70, 73, 75, 275, 307, 319, 324, 290, 302, 
    305, 327, 307, 327, 75, 63, 61, 16, 138, 66, 61, 305, 2, 103, 102, 70, 
    94, 69, 75, 83, 105, 103, 101, 91, 82, 96, 94, 89, 88, 90, 87, 89, 93, 
    75, 81, 80, 56, 296, 299, 310, 321, 334, 324, 316, 324, 24, 330, 346, 1, 
    35, 0, 45, 331, 319, 7, 312, 357, 341, 344, 299, 356, 353, 306, 358, 360, 
    312, 345, 8, 301, 353, 288, 309, 0, 296, 333, 330, 332, 0, 313, 318, 316, 
    359, 333, 321, 0, 351, 341, 343, 316, 5, 318, 349, 324, 356, 2, 20, 80, 
    301, 300, 306, 316, 292, 291, 277, 291, 288, 305, 298, 298, 291, 298, 
    317, 3, 313, 291, 313, 305, 94, 0, 0, 334, 82, 34, 358, 329, 321, 329, 
    337, 326, 308, 333, 275, 326, 314, 287, 335, 83, 294, 310, 324, 322, 329, 
    299, 332, 260, _, 124, 138, 8, 36, 200, 15, 54, 34, 115, 83, 83, 86, 102, 
    64, 132, 63, 12, 44, 302, 77, 309, 284, 298, 95, 70, 326, 320, 312, 288, 
    299, 320, 333, _, 72, 308, 305, 313, 289, 314, 318, 302, 344, 83, 77, 90, 
    83, 72, 91, 76, 88, 78, 61, 174, 58, 116, 72, 51, 325, 302, 307, 327, 73, 
    274, 299, _, 105, 348, 28, 336, 352, 350, _, 23, 13, 62, 59, 78, 25, 319, 
    306, 353, 307, 309, _, 335, 355, 3, 341, 359, 51, 313, 336, 58, 0, 0, 
    328, 323, 331, 25, 322, 319, 327, 0, 0, 24, 66, 330, 321, 304, 316, 323, 
    325, 320, 316, 14, 331, 312, 54, 339, 324, 18, 357, 333, 302, 301, 269, 
    343, 312, 2, 12, 71, 355, 64, 32, 58, _, 71, 312, 346, 58, 8, 360, 359, 
    26, 0, 78, 316, 289, 283, 350, 322, 355, 315, 360, 292, 0, 0, 313, 286, 
    2, 296, 301, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, 301, 324, 316, 87, 60, 4, 328, 351, 321, 346, 71, 
    97, 321, 146, 39, 34, 4, _, 45, 30, 59, 47, 334, 351, 134, 189, 152, 82, 
    357, 58, 96, 44, 6, 179, 103, 8, 140, _, 131, 115, 121, 109, 99, 134, 90, 
    88, _, 94, 96, 94, 84, 92, 94, 95, 86, 92, 93, 97, _, 94, 96, 103, 93, 
    85, 90, 100, 83, 91, 96, 73, 88, 89, 87, 64, 79, 84, 81, 62, 37, 58, 60, 
    51, 62, 57, 55, 54, 61, 65, 74, _, 64, 69, 73, 75, 69, 85, 64, 67, 91, 
    59, 35, 33, 41, 39, 33, 54, 45, 60, 60, _, 67, 53, 80, 68, 51, 49, 20, 
    26, _, 34, 37, 27, 33, 126, 37, 316, 349, 343, 317, 335, 326, 349, 329, 
    315, 326, 289, 339, 301, 296, 294, 299, 68, 67, 94, 69, 77, 81, 78, 83, 
    81, 89, 92, 83, 80, 82, 56, 40, 45, 64, 67, 73, _, 68, 79, 82, 59, 56, 
    61, 36, 243, 91, 60, 42, 3, 254, 173, 331, 60, 110, 84, 59, 48, 81, 277, 
    30, 57, 28, 75, 47, 48, 81, 58, 60, 49, 66, 58, 54, 61, 69, 69, 76, 70, 
    60, 59, 65, 76, 86, 69, 75, 47, 58, 90, 99, 91, 98, 99, 129, 272, 130, 
    86, 79, 105, 71, 92, 95, 70, 93, 6, 99, 82, 73, 56, 81, _, _, 83, 103, 
    93, 90, 52, 66, 66, 120, 113, 90, 79, 75, 64, 54, 58, 17, 360, 349, 63, 
    63, 272, 48, 12, 209, 68, 27, 69, 60, 53, 69, 97, 62, 112, 92, 106, 92, 
    74, 89, 21, 277, 308, 346, 319, 313, 306, 360, 311, 317, _, 305, 317, 
    306, 301, 317, 321, 304, 358, 307, 306, 325, 315, 338, 316, 329, 348, 
    322, 308, 330, 299, 314, _, _, 3, 337, 6, 331, 348, 350, 321, 328, 306, 
    314, 308, 302, 280, 289, 332, 336, 335, 340, 310, 41, 357, 334, 359, 290, 
    296, 35, 352, 335, 308, 310, 349, 34, 335, 19, 311, 319, 210, 286, 327, 
    13, 344, _, 296, 339, 343, _, 309, 90, 76, _, 314, 304, 88, 72, 66, 65, 
    77, 78, 70, 60, 249, 54, 347, 10, 36, 29, 214, 14, 355, _, _, _, 5, 18, 
    23, 38, 31, 21, 25, 6, 360, 9, 176, 90, 191, 205, 16, 104, 126, 206, _, 
    250, 220, 124, 219, 235, 259, 61, 26, 42, 36, 358, 59, 218, 76, 359, 234, 
    360, 360, 328, 308, 322, 309, _, 310, 308, 311, 313, 310, 311, 320, _, 
    307, 312, 357, 323, 358, 317, 351, 358, 311, 355, 324, 349, 3, 0, 355, 
    356, 0, 335, 307, _, _, _, 41, 332, 327, 314, 296, 318, 292, 302, 313, 
    325, 330, 337, 303, 49, 344, 15, 329, 320, _, 324, 317, 323, 341, 14, 
    319, 332, 306, 346, 323, 328, 343, 333, 300, 308, 3, 331, 322, 333, 357, 
    337, 349, _, 295, 339, 329, 317, 354, 0, 10, 343, 115, 322, 8, 336, 354, 
    305, 326, 42, 79, 95, 80, 89, 60, 59, 81, 96, 87, 78, 82, 85, 72, _, 97, 
    99, 106, 94, 95, 88, 93, 80, 79, 69, 40, 318, 18, 318, 41, 31, 78, 88, _, 
    2, 314, 295, 287, 294, 272, 293, 358, 309, 1, 0, 0, 353, 285, 308, 339, 
    309, 7, 326, 306, 44, 323, _, 186, 346, 58, 47, 313, 86, 43, 130, 349, 
    353, 323, 347, 2, 274, 69, 74, 76, 62, 79, 81, 99, 87, 72, 107, 98, 97, 
    92, 88, 87, _, 64, 327, 305, 308, 292, 323, 325, 318, 12, 97, 93, 333, 
    321, 55, 64, 41, 318, 316, _, 79, 319, 316, 6, 320, 304, 313, 352, 301, 
    84, 74, 345, 334, 359, 339, 327, 337, 38, 26, 353, 334, 351, _, 357, 344, 
    10, 71, 31, 11, 10, 301, 342, 8, 58, 24, 20, 306, 317, 78, 36, 310, 344, 
    6, 333, 109, 95, 324, 316, 332, 91, 344, _, _, 48, 338, 90, 6, 33, 313, 
    323, 9, 351, 55, 113, 350, 3, 29, 39, 27, 43, 45, _, 48, 30, 3, 17, 20, 
    5, 17, 16, 2, 40, 32, 42, 32, 32, 29, 31, _, 34, 37, 31, 26, 305, 306, 
    319, 26, 317, 318, 306, 299, 357, 342, 337, 14, 73, 186, 250, 148, 343, 
    34, 14, 2, 218, 9, 72, 41, 93, 53, 59, 66, 64, 73, _, _, 66, 72, 65, 69, 
    74, 66, 71, 104, 74, 97, 78, 96, 62, 107, 104, 289, 324, 338, _, 300, 
    310, 356, 321, 346, 335, 308, 323, 344, 350, 354, 21, 341, 157, 337, 6, 
    354, 1, 329, 305, _, 304, _, 312, 279, 341, 347, 307, 349, 278, 329, 335, 
    309, 238, 350, 57, 325, 69, 121, 55, 218, 88, 63, 234, 117, 195, 72, 343, 
    353, 26, 352, 2, _, 336, 316, 324, 352, 0, 332, 330, 50, 55, 312, 343, 
    307, 346, 328, 329, 311, 315, 319, 320, 357, 335, 320, 0, 357, 353, 330, 
    345, 297, 349, 317, 353, 345, 345, 3, 336, 360, 355, 3, 322, 10, 315, 74, 
    74, 74, 353, 334, 9, 359, 340, 347, 1, 318, 291, 1, 301, 20, 360, 16, 19, 
    26, 304, 100, 341, 0, 331, 333, 335, 64, 356, 335, 84, 16, 307, 42, 323, 
    304, 332, 332, 9, 303, 355, 309, 289, 75, 332, _, 330, 68, 321, 303, 354, 
    12, 29, 13, 324, 81, 75, 91, 95, 55, 46, 59, 307, 319, 307, 102, 65, 348, 
    84, 22, 46, 318, 322, _, 63, 65, 69, 106, 110, 97, 65, 53, 60, 47, 60, 
    62, 87, 77, 91, _, 54, 316, 302, 355, 334, 345, 307, 51, 95, 325, 104, 
    74, 307, _, 317, 305, 345, 326, 318, 62, 302, 315, 84, 72, 89, 301, 299, 
    _, 314, 278, 119, 340, 10, 77, 11, 0, 299, 349, 0, 359, 0, 51, 0, 312, 
    86, 347, 64, 16, 40, 341, 93, 85, 354, 31, 322, _, 301, 302, 301, 308, 
    314, 322, 315, 306, 284, 319, 348, 319, 301, 307, 328, 302, 324, 0, 16, 
    0, 13, 35, 347, 345, 355, 323, 309, 315, 300, _, 330, 321, 3, 57, 301, 
    323, 23, 325, 0, 333, 321, 291, 310, _, 350, 3, 14, 352, 324, 358, 97, 
    14, 352, 355, 37, 352, 358, 356, 339, 319, 36, 13, 343, 60, 344, 356, 38, 
    338, 347, 348, 50, _, 40, 305, 99, 347, 45, 49, 28, 12, 355, 0, 312, 63, 
    72, 77, 267, 301, 44, 65, 113, 45, 34, 0, 344, 16, 349, 76, 79, 312, 82, 
    349, 331, _, 13, 5, 81, 12, 310, 0, 332, 357, 355, 343, 4, 330, 71, 340, 
    332, 37, 316, 339, 86, 14, 296, 106, 342, 318, 67, 23, 17, 86, 347, 333, 
    316, 307, 75, 110, 2, 305, 305, 289, 130, _, 304, 324, 308, 315, 305, 
    255, 315, 315, 323, 315, 303, 322, 357, 311, 202, 199, 239, 245, 243, 
    237, 234, 243, 239, 254, _, 261, 293, 274, 271, 254, 234, 211, 252, 95, 
    340, 314, 307, 301, 288, 264, 300, 281, 262, _, 264, 268, 256, 270, 259, 
    269, 273, 281, _, 291, 313, 305, 344, 279, 307, 311, 303, 326, 323, 315, 
    _, 302, 323, 302, 17, 111, 294, 326, 275, 290, 281, 298, 88, 299, 72, 74, 
    5, 356, 29, 45, _, 24, 40, 32, 20, 50, 38, 49, 53, 44, 40, _, 349, 344, 
    38, 249, 360, 354, 319, 311, 295, 349, 34, 37, 29, 45, 25, 359, 23, 295, 
    254, _, 280, 287, 286, 20, 278, 317, 330, 139, _, 300, 324, 307, 310, 
    322, 206, 182, 244, 285, 288, 6, 62, 49, 276, 305, 291, 292, 358, 16, 8, 
    152, 353, 354, 297, 278, 353, 339, 6, 28, 37, 60, 345, 175, 27, 37, 217, 
    25, 271, 290, 249, 22, 249, _, 303, 6, 250, 354, 16, 257, 226, 274, 336, 
    269, 162, 86, 236, 181, 198, 238, 172, 39, 202, 315, 235, 47, 347, 329, 
    183, 292, 303, 48, _, 34, 103, 303, 205, 172, 324, 298, 355, 311, 298, 
    292, 336, 318, 320, 288, 302, 298, 308, 275, 355, 280, 300, 306, 282, 
    301, 296, 257, 300, 303, 306, 331, 285, 309, 280, 311, 305, 282, 266, 
    296, 303, 296, 324, _, 303, 1, 298, 9, 6, 35, 23, 20, 325, 336, 304, 316, 
    325, 295, 307, 348, 330, 304, 327, 3, 320, 293, 340, 289, 351, 322, 316, 
    328, 314, 352, 272, 352, 326, 275, 302, 290, 27, 153, 237, 321, 27, 267, 
    269, 301, 325, 279, 338, 308, 326, 0, 328, 281, 316, 0, 309, 320, 325, 
    347, 326, 354, 12, 327, 328, 328, 283, 329, 306, 339, 317, 0, 338, _, 
    353, 347, 354, 317, 332, 355, 1, 345, 45, 320, 357, 329, 299, 354, 335, 
    311, 356, 307, 9, 102, 76, 107, 300, 340, 81, 345, 8, 39, 342, 360, 30, 
    78, 94, 352, 357, 35, 64, 77, 53, 81, 124, 241, 105, 180, 197, 51, 21, 
    79, 281, 11, 76, 5, 349, 32, 73, 73, 307, 246, 64, 65, 74, 77, 84, 88, 
    85, 58, 59, 52, 54, 73, 96, _, _, 86, 93, 65, 283, 281, 80, 311, 73, 84, 
    77, 105, 89, 87, 82, 97, 101, 108, 119, 95, 324, 260, 326, 81, 76, 316, 
    303, 301, 300, 301, 309, 309, 295, 308, 296, 303, 321, 312, 303, 277, 
    297, 5, 1, 0, 347, 287, 350, 73, 8, 356, 295, 347, 16, 46, 64, 357, 339, 
    344, 51, 337, 23, 334, 312, 312, 329, 8, 197, 333, 20, 44, 43, _, _, 45, 
    38, 23, 7, 4, 3, 2, 8, 3, 9, 3, 3, 2, 3, 11, 13, 18, 42, 37, 36, 32, 43, 
    29, 41, 25, 26, 343, _, 190, 282, 173, 202, 272, 358, 27, 349, 346, 284, 
    298, 314, _, 338, 320, 294, 332, _, 45, 315, 357, _, 339, 4, 352, 316, 
    316, 355, 21, 9, 196, 336, 295, 24, 300, 167, 327, 137, 10, 355, 6, _, _, 
    _, 357, 40, 328, 0, 360, 342, 354, 287, 342, 331, 10, 345, 0, 360, 330, 
    304, 303, 305, _, 314, 329, 315, 343, 322, 334, 327, 319, 75, 353, 26, 
    319, 306, 314, 311, 293, 313, 304, 305, 296, 330, _, _, 311, 300, 306, 
    284, 298, 308, 309, _, 320, 299, 330, 11, 0, 78, 358, 81, 87, 77, 105, 
    82, 34, 78, 289, 305, 318, 263, 267, 105, _, _, 15, 43, 64, 84, 8, 10, 
    346, 337, 341, 37, 1, 32, 344, 70, 274, 317, 53, 33, _, 101, 305, 322, 
    101, 334, 0, 81, 304, 303, 9, 10, 354, 320, 0, 0, 0, 351, 0, 124, 0, 0, 
    21, _, 287, 0, 0, 0, 343, 18, 3, _, 0, 0, 325, 8, 339, 0, 10, 358, 329, 
    360, 10, 0, 0, 324, 294, 58, 45, 0, 66, 309, _, _, 330, 45, 23, 11, 352, 
    353, 28, _, 328, 349, 353, 346, 0, 351, 284, 275, 287, 76, _, 355, 20, 
    30, 20, 22, 28, 353, 38, 26, 34, 14, 15, 55, 30, 32, 36, 44, 52, 58, 54, 
    43, 49, _, 38, 46, 53, 43, 211, 285, 236, 321, 52, 227, 27, 282, 306, 
    115, 35, 14, 2, 333, 56, 29, 208, 73, 87, 13, 240, 245, 309, 6, _, _, 20, 
    32, 280, 254, 269, 335, 314, 270, 293, 288, 303, 286, 21, 327, 305, 53, 
    313, 349, _, 285, _, 54, 76, 218, 302, 27, 199, 71, 211, 117, 57, 339, 
    339, 106, 327, 327, 300, 268, 320, 284, 234, _, 173, 74, 50, 322, 270, 
    324, 317, 253, 315, 356, 34, 290, 10, 149, 274, 13, 68, 112, 8, 10, 61, 
    42, 5, 334, 41, 14, 1, 26, _, _, 37, 52, 37, 344, 348, 239, 262, 353, 
    310, 25, 25, 43, 32, 356, 40, 31, 34, 11, _, 9, _, 33, 9, 47, 39, 67, 
    237, 55, 151, 177, 143, 350, 170, 35, 199, 289, 269, 78, 205, _, 236, _, 
    223, 169, 263, 291, 305, 334, 345, 304, 314, 134, 355, 254, 296, 36, 289, 
    111, 95, 323, 335, 23, 43, 169, 142, 37, 25, 31, 26, 41, _, _, 34, 38, 
    29, 34, 27, 28, 32, 358, 278, 70, 54, 221, 282, 179, 313, 282, 257, 236, 
    _, 224, 212, 222, 116, 146, 68, 54, 302, 32, 319, 309, 326, 349, 276, 
    265, 271, 349, 356, 350, 276, 271, 257, _, 272, 269, 280, 274, 322, 335, 
    321, 354, 315, 306, 325, 343, 36, 329, 313, 0, 294, 340, _, 322, 331, 
    268, 274, 258, 273, 280, 257, 350, 301, _, 86, 356, 324, 99, 8, 351, 310, 
    335, 344, 338, 22, 323, 355, 270, 273, 277, 275, 245, _, 94, 179, 262, 
    30, 1, 292, 181, 239, 209, 167, 192, 51, 8, 83, 286, 55, 347, 77, 47, 24, 
    352, 149, 329, 306, 282, 318, 10, 0, 117, 104, 107, 30, 50, 7, 0, 68, 40, 
    4, 58, 66, 1, 334, 0, 0, 121, 103, 270, 250, 321, 69, 143, 263, _, 96, 
    57, 52, 43, 317, 27, 38, 36, 25, 17, 322, 67, 141, 124, 105, 117, 152, 
    157, 309, 190, 203, 181, 173, 45, 219, 25, 205, 163, 356, 359, 315, 33, 
    5, 197, 2, 327, 224, 181, 199, 203, 254, 193, 287, 88, 278, 0, 0, 44, 30, 
    122, 0, 0, 0, 321, 347, 342, 64, 350, 329, 0, 283, 269, 321, 279, 264, 
    279, 278, 261, 302, 203, 56, _, 314, 74, 81, 110, 76, 79, 93, 287, 309, 
    280, 303, 291, 338, 279, 291, 280, 277, 259, 90, 113, 105, 82, 298, 335, 
    303, 332, 298, 29, 309, 337, 55, 305, 2, 309, 355, 0, 0, 13, 244, 160, 
    225, _, 241, 259, 269, 2, 0, 346, 66, 322, 67, 328, 319, 305, 20, 52, 
    302, 90, 0, 302, 288, 65, 154, 116, 270, 5, 325, 292, 294, 6, 360, _, 30, 
    14, 70, 299, 114, 0, 93, 288, 99, 344, 20, 45, 41, _, 332, 274, 343, 154, 
    0, 0, 267, 353, 100, 0, 292, 0, 343, 319, 360, 0, 1, 344, 307, 292, 87, 
    335, 41, 329, 127, 77, 344, 33, 85, 105, 111, 344, 1, 344, 344, 309, 84, 
    42, 314, 322, 318, 97, 350, 304, 0, 351, 124, 308, 154, 144, 188, 242, 
    355, 100, 285, 98, 148, _, 0, 32, 0, 0, 0, 114, 133, 316, 338, 330, 146, 
    117, 156, _, 170, 150, 146, 179, 131, 119, 100, 97, 109, 104, 107, 124, 
    315, 305, 129, 74, 348, 124, 310, 279, 194, 162, 155, 149, 156, 122, 168, 
    _, 145, 145, 122, 104, 124, 152, 127, 103, 86, 72, 91, 82, 86, 72, 75, 
    62, 72, 92, 107, 93, 112, 96, 96, 93, 99, 108, 110, 113, 110, 113, 102, 
    105, 107, 100, 77, 68, 59, 277, 303, 269, 267, 282, 265, _, 273, 118, 
    123, 100, 100, 97, 95, 96, _, 93, 95, 97, 99, 96, 101, 91, 88, 90, 101, 
    106, 100, 114, 92, 104, 107, 122, 117, 118, 115, 114, 112, 112, 112, 113, 
    107, 103, 94, 84, 76, 88, 88, 308, 276, 293, 263, 278, 201, 133, 100, 
    100, 106, 135, 104, 91, 107, 112, 85, 22, 303, 301, 311, 5, 0, 343, 26, 
    344, 8, 224, 290, 337, 267, _, 125, 35, 158, 0, 166, 11, 149, 10, 154, 
    354, 1, 317, 318, 316, 315, 296, 117, 72, 128, 298, 318, 266, 271, 274, 
    275, 274, 294, 269, 164, 124, 224, 278, 291, 52, 46, 279, 293, 297, 342, 
    285, 304, 95, 79, 91, 84, 87, 90, 93, 96, 97, 97, 86, 87, 95, 100, 101, 
    97, 97, 84, 87, 89, 90, 104, 100, 99, 102, 94, 102, 105, 108, 104, 104, 
    106, 100, 85, 78, 84, 94, 94, 84, 85, 79, 90, 92, 90, 80, 80, 89, 89, 83, 
    85, 87, 88, 89, 95, 97, 95, 93, 96, 100, 97, 97, 95, 95, 82, 80, 87, 83, 
    101, 104, 102, 88, 92, 83, 104, 37, 82, 41, 47, 40, 29, 8, 8, 19, 46, 
    258, 16, 66, 46, 70, 9, 53, 18, 43, 42, 46, 43, 44, 61, 43, 77, 129, 278, 
    282, 168, 171, 165, 229, 279, 224, 261, 256, 269, 285, 282, 90, 78, 79, 
    76, 91, 50, 62, 85, 77, 85, 79, 120, 63, 70, 104, 117, 108, 114, 121, 
    121, 121, 107, 79, 115, 338, 353, 346, 2, 331, 74, 0, 91, 118, 45, 115, 
    100, 99, 104, 109, 107, 105, 103, 114, 54, 15, 60, 39, 39, 81, 122, 70, 
    90, 69, 145, 72, 74, 35, 37, 68, 41, 44, 58, 58, 56, 44, 45, 65, 8, 10, 
    11, 34, 49, 39, 34, 39, 35, 40, 26, 35, 45, 41, 34, 50, 156, 159, 141, 
    251, 163, 170, 173, 173, 153, 188, 108, 175, 224, 254, 217, 17, 0, 360, 
    244, 357, 177, 246, 223, 264, 334, 328, 254, 231, 283, 208, 210, 177, 
    166, 144, 122, 64, 274, 298, 308, 297, 350, 230, 20, 121, 268, 253, 244, 
    128, 159, 135, 273, 274, 287, 253, 267, 257, 269, 271, 271, 286, 284, 
    311, 314, 325, 308, 315, 324, 313, 303, 296, 300, 262, 192, 108, 158, 
    136, 150, 173, 206, 256, 270, 283, 261, 257, 293, 334, 3, 0, 302, 101, 
    56, 98, 93, 173, 103, 106, 263, 123, 121, 164, 160, 146, 134, 122, 358, 
    160, 138, 129, 0, 258, 0, 16, 2, 106, 0, 70, 93, 350, 163, 165, 229, 180, 
    171, 193, 189, 184, 208, 112, 77, 201, 62, 202, 150, 60, 114, 64, 55, 
    172, 93, 79, 53, 62, 64, 76, 68, 84, 48, 87, 128, 168, 154, 139, 67, 143, 
    92, 183, 164, 292, 328, 167, 334, 212, 294, 126, 153, 75, 270, 283, 290, 
    280, 296, 286, 274, 263, 251, 109, 55, 83, 330, 309, 1, 8, 65, 358, 225, 
    245, 333, 146, 132, 71, 128, 117, 136, 74, 94, 199, _, 294, 309, 298, 
    293, 305, 302, 286, 260, 252, 242, 267, 292, 298, 285, 267, 256, 266, 
    259, _, 267, 266, 268, 267, 255, 270, 266, 272, 273, 285, 280, 307, 324, 
    322, 113, 95, 317, 320, 329, 136, 124, 40, 129, 130, 120, 130, 122, 147, 
    _, _, _, 262, 261, 249, 274, 317, 113, 117, 113, 6, 253, 258, 266, 287, 
    262, 123, 123, 268, 104, _, 156, 166, _, 168, 171, 149, 159, 134, 112, 
    114, 119, 135, 124, 5, 118, 120, 139, 118, 137, 131, 140, _, 146, 139, 
    143, 146, 179, 291, 159, 133, 142, 142, 153, 90, 143, 171, 69, 108, 140, 
    178, 153, 148, 122, 52, 93, 333, 228, 231, 254, 313, _, 157, 80, 76, 74, 
    61, 260, 176, 211, 300, _, 130, 109, 85, 11, 183, 169, 179, 163, 170, 
    197, _, 131, 135, _, 207, 51, 28, 23, 56, 30, 30, 357, 25, 94, 25, 55, 
    27, 61, 39, 85, 347, 74, 128, _, 32, 52, 354, 18, 36, 98, 63, _, 56, 61, 
    70, 48, 55, 73, 93, 61, 71, 68, 15, 139, 42, 31, 116, 66, 100, 54, 310, 
    18, _, 49, 48, 49, 48, 47, 51, 44, 39, 56, 108, 336, 132, 68, 64, 46, 67, 
    60, 70, 69, _, 67, 82, _, 78, 73, 67, 66, 63, 73, 72, 57, 65, 54, 58, 
    260, 74, 56, 80, 83, 85, _, 60, _, 54, _, 66, 68, _, 57, 50, 65, 70, _, 
    95, 27, 46, 224, _, 172, 81, 5, 221, _, 120, 135, 163, 157, _, 167, 153, 
    _, _, _, 165, 160, 82, 241, _, 121, 90, 79, 306, 240, 242, 289, 334, 76, 
    265, 29, _, 32, _, 26, _, _, 31, 89, 89, 68, 95, 112, 90, 325, 45, _, 
    161, 169, 23, 98, _, 131, 356, _, 98, _, 128, 241, 250, 284, _, 276, 278, 
    _, 288, _, 291, 282, 69, 167, _, 144, 82, 187, 85, _, 127, 106, 163, 168, 
    _, 39, 278, 271, _, _, 287, 285, 116, 259, _, 271, 278, 285, 189, 71, 
    160, 71, 67, 45, 55, 51, _, 72, _, 79, 83, 77, 54, 69, 60, 60, 37, 47, 
    56, 41, 61, 81, 149, 52, 88, 92, 72, 77, 86, 109, _, _, 75, 62, 101, 133, 
    _, 170, 128, 142, 172, _, 171, 226, 172, 138, _, 74, 97, 103, 108, _, 
    176, 179, 173, 157, _, 141, 153, 147, 157, _, 164, 141, 132, 74, _, 169, 
    130, 17, _, 82, 132, 131, 120, 117, 145, 161, 150, 152, _, 144, 142, 130, 
    144, 137, 131, 118, 103, 82, 114, 51, 137, _, 44, 128, 115, 261, 57, 44, 
    60, 216, _, 53, 81, 122, 259, 64, _, 360, 359, 32, 69, _, 209, 224, 272, 
    263, _, 216, 298, 144, 129, _, 99, 100, 98, 128, 140, 249, 269, 99, 126, 
    _, 118, 36, 140, 40, _, 144, 202, 192, 336, 129, 13, 308, 294, 292, 306, 
    252, 315, 291, _, 149, 163, 129, 115, 119, 273, 285, 272, 278, 205, 336, 
    151, _, 138, 116, 283, 267, _, 304, 116, 268, 251, 111, 95, 135, 119, 
    123, 136, 127, 160, 170, 169, _, 287, 59, 167, 0, 249, 261, 296, 343, 
    163, _, 131, 141, 120, 246, _, 255, 268, 264, 269, _, 258, 289, 241, 273, 
    279, 297, 275, 286, 271, 288, 285, _, 249, 275, 288, 258, _, 254, 256, 
    256, 266, 266, 230, 246, 270, 265, _, 292, 277, 257, 271, _, 294, 296, 
    314, 312, _, 293, 260, 306, 292, 291, 282, 297, 270, 269, _, 259, 285, 
    287, 288, _, 276, 162, 49, 105, _, 138, 123, 118, 120, _, _, _, 106, 171, 
    _, 167, 179, 270, 272, _, 285, 288, 284, 312, 295, 312, _, 314, 277, 274, 
    264, 304, 268, 311, 312, 287, 308, 296, 291, 292, 286, 273, 285, 298, 
    280, 284, _, 301, 290, 290, 287, 293, 285, 296, 306, 300, 311, 315, 299, 
    259, 270, 269, 255, 248, 257, 272, 287, 273, 266, 291, 285, 305, 305, 
    320, 322, 314, 170, 162, 76, 81, 300, 143, 152, _, 106, 122, 123, 91, 68, 
    140, 135, 132, 136, 136, 127, 126, 145, 121, 104, 320, 332, 121, 133, 
    346, 283, _, 281, 302, 109, 132, 125, 135, 126, 253, 289, 300, 301, 299, 
    262, 293, 300, 296, 297, 90, 78, 284, 299, 301, 300, 295, 276, 293, 105, 
    103, 292, 147, 180, 299, 182, 175, 170, 119, 120, 136, 97, 146, 155, 0, 
    111, 0, 125, 0, 131, 108, 145, _, 123, 134, 127, 125, 128, 123, 116, 166, 
    168, 159, 146, 146, 164, 124, 302, 195, 304, _, 59, 130, 122, _, 146, 
    118, 123, 122, 134, 143, 64, 126, 284, 236, 124, 103, 118, 107, 318, 92, 
    81, 219, 269, 255, 230, 228, 175, 168, 137, 127, 106, 119, 147, 140, 140, 
    125, 126, 132, 131, 143, 147, 134, 160, 139, 131, 116, 169, 133, 156, 
    128, 134, 126, _, _, 143, 132, 152, 138, 132, 146, 135, _, 127, 118, 116, 
    126, 127, 131, 131, 0, 358, 6, 0, 0, 62, _, 183, 173, 151, 168, 122, 101, 
    134, _, 97, 104, 115, 102, 116, 97, 94, 108, 39, 110, 328, 29, 59, 0, 89, 
    8, 126, 172, 176, 249, 147, 124, 271, 86, 261, 71, 82, 42, 65, 51, 75, 
    45, 288, 240, 233, 298, 33, 50, 334, 221, 220, 286, 28, 231, 241, 282, 
    302, 49, 86, 105, 89, 6, 161, 285, 198, 201, 109, 237, 170, 12, 103, 62, 
    170, _, 52, 80, 78, 71, 2, 64, 77, 165, 163, 164, 150, 123, 125, 81, 98, 
    118, 78, 127, 51, 100, 302, 333, 20, 144, 172, 122, 125, 133, 143, 146, 
    151, 164, 136, 142, 156, 129, 166, 159, 110, _, 109, 118, _, 118, 95, 
    130, 137, 127, 123, 116, 126, 123, 123, 112, 114, 102, 109, 116, 109, 
    111, 69, 97, 117, 100, 89, 86, 74, 67, 79, 70, 68, 117, 152, 150, 127, 
    97, 112, 109, 111, 112, 124, 113, 113, 117, 100, 97, 108, 108, 98, 74, 
    182, 86, 77, 76, 94, 99, 97, 128, 117, 148, 114, 103, 132, 112, 138, 133, 
    139, 114, 104, 82, 85, 94, 105, 93, 113, 242, 292, 47, 133, 138, 115, 
    145, 145, 119, 146, 146, 132, 134, 141, 112, 117, 115, 108, 122, 76, 142, 
    135, 91, 96, 111, 143, 155, 143, 131, 116, 160, 132, 124, 167, 61, 158, 
    _, 144, 63, 85, 180, 119, 122, 107, 142, 117, 88, 89, 111, 100, 73, 88, 
    99, 90, 100, 85, 112, 91, 131, 127, 98, 110, 104, 105, 99, 115, 108, 111, 
    122, 35, 324, 313, 347, 314, 307, 360, 46, 19, 147, 119, 304, 114, 137, 
    313, 56, 277, 317, 237, 130, 11, 98, 133, 31, 12, 67, 276, 2, 321, 331, 
    69, 90, 143, 136, 12, 223, 123, 217, 252, _, 254, 332, 152, 57, 154, 161, 
    297, 249, 358, 332, 1, 283, 194, 294, 24, 172, 234, 4, 235, 183, 253, 
    300, 269, 145, 141, 143, 112, 117, 126, 126, 125, 166, 60, 313, 343, 233, 
    200, 319, 13, 220, 233, 179, 232, 195, 128, 137, 124, 156, 136, 146, 116, 
    115, 108, 111, 122, 104, 123, 125, 113, _, 136, 309, 341, 132, 116, 109, 
    115, 125, 133, 142, 118, 121, 111, 53, 110, 125, 67, 161, 118, 326, 319, 
    236, 171, 165, 1, 116, 74, 114, 125, 109, 100, 102, _, 281, 83, 77, 13, 
    117, 114, 90, 89, 111, 100, 97, 86, 60, 49, 61, 56, 146, 103, 43, 74, 52, 
    _, 24, _, 73, 125, 131, 111, 145, 106, 103, 98, 85, 114, 88, 131, 0, 55, 
    109, 119, 101, 89, 95, 94, 108, _, 109, 111, 131, 102, 112, 116, 107, 84, 
    296, 118, 260, 97, 111, 104, 109, _, 100, 308, _, 316, 278, 273, 279, 
    271, 236, 255, 237, _, 225, 275, 269, 267, 264, 265, 273, 275, 291, 292, 
    _, 316, 320, 309, 309, 314, 152, 111, 189, 156, 161, 165, 149, 360, 256, 
    251, 272, 267, 233, 267, 288, 181, 173, 182, 236, 301, 355, 177, 112, 88, 
    110, 128, 147, 144, 122, 123, 127, 131, 116, 127, 117, 105, 100, 120, 
    125, 123, 122, 112, 358, 133, 120, 119, _, 101, 106, 106, 114, 359, 139, 
    168, 175, 185, 169, 168, 174, 167, 57, 175, 148, 129, 98, 94, _, 126, 97, 
    60, 76, 330, 304, 247, 30, _, 67, 147, 71, 74, 238, 98, 63, 86, 65, 64, 
    8, 4, 69, 27, 273, 303, 303, 345, 91, 272, _, 94, 20, 224, 170, 160, 117, 
    134, 137, 145, 123, 127, 127, 129, 135, 128, 0, 91, 319, 0, 315, 353, _, 
    126, 100, 139, 131, 121, 151, 147, 125, 160, 119, 132, 123, 126, 119, 
    112, 109, 75, 339, 321, _, 322, 346, 352, 48, 344, 328, 195, 288, 259, 
    261, _, 225, 219, 217, 241, 265, 234, 240, 249, 268, 266, 286, 299, 308, 
    324, 296, 294, 297, 292, _, 347, _, 280, 213, 42, 70, 68, 64, 55, 75, 61, 
    62, 70, 55, 300, 99, 282, 330, 73, 175, 90, _, 3, 49, 71, 71, 69, 70, 96, 
    124, 122, 168, 141, 116, 97, 122, 136, 188, 276, 273, 291, _, 51, 49, 47, 
    66, 65, 50, 77, 54, _, 72, 69, 96, 51, 33, 224, 65, 72, 88, 69, 252, 65, 
    67, 310, 72, 48, 65, 48, 317, 27, _, _, _, 61, 18, 199, 95, 60, 63, 80, 
    65, 306, 55, 339, 83, 52, 343, 54, 316, 324, 326, 335, 1, _, 262, 33, 75, 
    159, 133, 120, 100, 119, 115, 116, 106, 172, 39, 267, 269, 280, 117, 174, 
    _, 70, 346, 159, 166, 176, 333, 191, 288, 284, 258, 251, 270, 237, 178, 
    176, 192, 266, 274, 269, 278, 268, 272, 249, 254, 251, 258, 243, 261, 
    266, _, 235, 225, 236, 246, 177, 318, 304, 182, 235, 199, 298, 237, 292, 
    283, 294, 294, 293, 283, 285, 265, 276, 334, 269, 204, 258, 192, 244, 
    235, 148, 126, 134, 124, 135, 142, 119, 103, 111, 118, 88, 116, 102, 83, 
    89, 114, 129, 75, 38, 113, 130, 140, 133, 145, 136, 127, 163, 131, 110, 
    104, 167, 171, 186, 346, 177, 105, 96, 145, 341, 306, 280, 280, 281, 274, 
    266, 258, 266, 213, 83, 126, 125, 126, 157, 146, 157, 133, 141, 142, 138, 
    202, 317, 16, 316, 355, 304, 300, 295, 291, 301, 346, 250, 272, 175, 218, 
    210, 195, 176, 139, 78, 53, 23, 39, 21, 17, 8, 33, 13, 38, 42, 48, 44, 
    16, 4, 189, 159, 69, 89, 120, 105, 140, 113, 72, 27, 52, 38, 45, 49, 33, 
    106, 4, 7, 43, 278, 350, 350, 81, 337, 352, 341, 75, 219, 69, 69, 75, 68, 
    66, 69, 80, 75, 58, 43, 129, 44, 41, 41, 27, 34, 42, 49, 106, 103, 82, 
    351, 79, 62, 58, 71, 77, 133, 121, 103, 87, 142, 185, 195, 70, 341, 358, 
    359, 19, 155, 264, 88, 126, 131, 135, 119, 147, 174, 173, 177, 65, 104, 
    124, 105, 62, 125, 300, 276, 339, 166, 0, 43, 0, 0, 0, 0, 13, 157, 101, 
    116, 109, 113, 115, 127, 115, 127, 118, 100, 213, 242, 286, 211, 32, 296, 
    255, 250, 231, 293, 355, 71, 258, 233, 243, 256, 262, 274, 280, 283, 271, 
    274, 272, 273, 291, 305, 311, 299, 288, 295, 302, 303, 304, 320, 328, 
    330, 287, 236, 233, 261, 223, 235, 272, 235, 264, 276, 281, 282, 269, 
    275, 298, 307, 317, 0, 0, 113, 286, 0, 0, 355, 254, 295, 121, 159, 148, 
    178, 135, 118, 101, 100, 101, 121, 124, 96, 116, 90, 77, 102, 128, 127, 
    181, 309, 0, 192, 0, 351, 330, 291, 58, 351, 0, 283, 106, 109, 109, 143, 
    329, 298, 298, 298, 292, 288, 294, 292, 296, 303, 298, 291, 303, 288, 
    305, 298, 281, 225, 136, 102, 250, 311, 284, 114, 243, 315, 307, 299, 
    291, 283, 308, 292, 297, 291, 283, 272, 314, 306, 307, 312, 315, 315, 
    290, 307, 58, 305, 301, 304, 288, 294, 303, 324, 300, 315, 310, 339, 320, 
    311, 288, 201, 34, 106, 86, 101, 126, 114, 117, 117, 0, 151, 122, 326, 
    312, 319, 288, 305, 101, 293, 289, 295, 286, 276, 256, 288, 277, 272, 
    297, 302, 299, 288, 275, 263, 272, 269, 269, 268, 286, 282, 304, 289, 
    309, 317, 312, 307, 321, 316, 322, 325, 294, 295, 290, 290, 293, 279, 
    276, 284, 285, 296, 276, 287, 269, 289, 307, 297, 288, 289, 356, 25, 352, 
    39, 47, 54, 90, 297, 77, 61, 75, 55, 32, 25, 70, 344, 317, 287, 297, 295, 
    304, 308, 321, 309, 326, 349, 330, 311, 301, 354, 85, 85, 29, 283, 295, 
    285, 178, 173, 162, 183, 176, 193, 270, 292, 309, 0, 63, 108, 110, 341, 
    9, 267, 303, 283, 16, 40, 11, 27, 39, 57, 290, 311, 76, 58, 61, 49, 48, 
    11, 353, 77, 242, 54, 98, 167, 350, 293, 317, 259, 83, 77, 249, 157, 47, 
    71, 318, 266, 239, 78, 87, 102, 247, 11, 345, 28, 350, 0, 0, 340, _, 357, 
    111, 52, 72, 26, 352, 355, _, 35, 157, 172, 135, 310, 320, 331, 32, 350, 
    342, 327, 323, 308, _, 289, 66, 341, 223, 60, 46, 17, 333, 293, 281, 290, 
    290, 301, 292, 288, 301, 279, 293, 278, 281, 284, 273, 266, 292, 292, 
    279, 293, 285, 282, 301, 290, 286, 286, 288, 284, 302, 311, 294, 319, 
    302, 304, 272, 308, 12, 35, 105, 183, 245, 115, 23, 46, 37, 1, 20, 54, 
    59, 85, 96, 66, 86, 118, 61, 74, 84, 95, 63, 121, 283, 298, 296, 281, _, 
    344, 334, 356, _, 187, 358, 294, 257, 246, 333, 271, 278, 325, 186, 221, 
    150, 129, 250, 124, 85, _, 95, 349, 70, 341, _, 353, 343, 331, 355, 222, 
    298, 277, 179, _, 179, _, 125, 197, 314, 128, 85, 65, 92, 57, 0, 2, 297, 
    353, 0, 121, 0, 356, 38, 266, 81, 142, 183, 297, 299, 269, 271, 269, 275, 
    272, 267, 274, 253, 277, 272, 280, 267, 289, 302, 309, 314, 309, 297, 
    325, _, 281, 57, 110, 169, 127, 126, 119, 110, 84, 71, 76, 72, _, 74, 
    278, 306, 291, 301, 321, 344, 355, 25, 178, 355, 218, 148, 150, 129, 105, 
    98, 108, 128, 109, 130, 38, 337, 317, 316, 325, 327, 340, 296, _, 357, _, 
    324, 0, 266, 158, 125, 132, 140, 132, 126, 97, 121, 136, 166, 311, 298, 
    290, 322, 297, 238, 10, 306, 25, 79, 293, 322, 0, 306, 268, 259, 264, 
    119, 129, 0, 267, 139, 39, 6, 14, 316, 294, 330, 315, 297, 333, 357, 338, 
    348, 355, 303, 292, 266, 183, 5, 168, 97, 105, 110, 69, 141, 144, 161, 
    300, 305, 299, 284, 342, 39, _, 319, _, 8, 79, 0, 74, 79, 122, 4, 146, 
    127, 93, 110, 126, 136, 90, 360, 111, 29, 0, 359, 343, _, 22, 352, _, 26, 
    348, 299, 354, _, 153, 119, 155, 153, 155, 139, 25, 217, 78, 132, 312, 
    125, 305, 0, 358, 44, 357, 359, 0, 3, _, 19, 0, 0, 269, 132, 151, 138, 
    127, 143, 134, 95, 142, _, 309, 79, 316, 46, 337, 347, 28, 59, _, 5, 360, 
    65, 331, 17, 276, 50, 101, 315, 293, 109, 103, 0, 353, 14, 349, 41, 315, 
    347, 334, _, 310, 326, 82, 315, 7, 25, 8, 0, 292, 115, 168, 228, 165, 
    345, 129, 130, 354, 305, 354, 10, 0, 325, 43, 313, 343, 85, 50, 12, 12, 
    32, 336, 108, 4, 345, 0, 126, 250, 293, 130, 255, 306, 312, 318, 352, 6, 
    50, 331, 329, 314, 298, 300, 75, 65, 347, 29, 318, 290, 318, 318, 110, 
    337, 73, 296, 287, 275, 317, 313, 301, 299, 317, 293, 298, 302, 293, 294, 
    324, 308, 324, 332, 332, 313, 329, 334, 102, 100, 137, 102, 60, 87, 56, 
    40, 321, 311, 310, 88, 320, 302, 123, 0, 319, 307, 311, 206, 4, 119, 101, 
    118, 125, 123, 87, 126, 109, 76, _, 305, 308, 296, 288, 326, 350, 336, 
    33, 280, 92, 315, 355, 49, 320, 324, 352, 290, 98, 319, 303, 61, 334, 
    293, 328, 308, 307, 296, 331, 314, _, 321, _, 281, 102, 290, 35, 265, 
    331, 108, 283, 289, 280, 74, 48, 358, 53, 64, 76, 55, 327, 264, _, 258, 
    270, 270, 266, 267, _, 278, 272, 297, 302, 288, 277, 291, 292, 292, 295, 
    292, 301, 307, _, 298, 294, 339, 334, 306, 306, 11, 7, 344, 322, 354, 23, 
    348, 13, 124, 0, 309, 349, 288, 300, 291, 284, 290, 285, 298, 101, 301, 
    7, 348, _, 293, _, 88, 81, 39, 78, 290, 297, 262, 273, 278, 273, 267, 
    271, 285, 273, 269, 274, 281, 323, 325, 316, 297, 315, 305, 238, 43, _, 
    304, 23, 283, 285, 78, 58, 271, 267, 263, 255, 253, 286, 287, _, 298, 
    292, 293, 286, 251, 281, 333, 323, 317, 310, 301, 331, 310, 301, 37, 13, 
    310, 303, 92, 43, 69, 328, 310, 352, 0, 36, 115, 350, 0, _, 1, _, 2, 0, 
    0, 116, 28, 324, 107, 0, 0, 30, 0, 0, 310, 5, 21, 290, 142, 93, _, 329, 
    0, 303, 327, 332, 314, _, 0, 358, 321, 0, 0, 0, 25, 104, 61, 349, 329, 
    100, 1, _, 337, 9, 293, 305, 333, 356, 22, 59, 48, 27, _, 338, 100, 81, 
    336, 88, 128, 300, 286, 127, 96, 324, 106, 338, 95, 95, 51, 346, 50, _, 
    289, 310, 344, 322, 316, 83, 325, 354, 358, 357, 2, 351, 280, 74, 199, 
    291, 305, 320, 316, 78, 103, 104, _, 285, 4, 31, 343, 313, 310, 23, 8, 
    11, 32, 325, 102, 259, 330, 43, 64, 316, 341, _, 323, 346, 342, 343, 0, 
    87, 352, 63, _, 288, _, 11, 5, 23, 44, 353, 27, 48, 23, 39, 55, 58, 54, 
    63, 37, 57, 129, 143, 64, _, 45, _, 81, 76, 92, 214, 228, 340, 360, 358, 
    3, 8, 5, 12, 19, 22, 19, 22, 32, 39, 44, _, _, 25, 20, 24, 19, 16, 16, 
    21, 14, 7, 20, 10, 10, 34, 43, 53, 9, 19, 36, 40, 230, 257, 228, 229, 
    212, 201, 271, 191, 243, 22, 19, 125, 8, 16, 76, 107, 360, 248, 82, 347, 
    32, 0, 16, 307, 297, 323, 341, 354, 35, 40, 305, 300, 44, 319, 315, 319, 
    288, 290, 293, 300, 333, 311, 323, 289, 290, 298, 309, 291, 282, 288, 
    316, _, _, 338, 323, 312, 333, 315, 0, 305, 314, 290, _, 295, 286, 293, 
    310, 75, 0, 318, 345, 71, 298, 8, 310, 320, 308, 33, 78, 290, 101, 316, 
    _, 309, 311, 44, 80, 68, 319, 306, 295, 301, 299, 314, 326, 327, 313, 53, 
    334, 351, 40, 360, 326, 330, 346, 86, 54, 148, 20, 359, 277, 287, 296, 
    300, 333, 317, 12, 57, 74, 321, 281, 294, 334, 325, 317, 308, 111, 91, 
    103, 303, 290, 290, 281, 277, 267, 266, 273, 288, 272, 271, 285, 272, 
    313, _, 289, 236, 296, 284, 268, _, 298, 289, 273, 290, 303, 304, 342, 
    323, 215, 297, 37, 348, 334, 304, 0, 357, 27, 4, 0, 329, 91, 67, 330, 
    343, 345, 351, 321, 279, 321, 353, 319, 24, 89, 315, 253, 289, 308, 311, 
    258, 355, 309, 317, 311, 299, 319, _, _, 310, 310, 300, 274, 255, 291, 
    279, 284, 254, 301, 294, 313, 319, 310, 306, 313, 316, 274, 304, 310, 
    312, 305, 299, 319, _, 317, 322, 313, 307, 299, 313, 323, 319, 66, 88, 
    317, 309, 320, 325, 70, 46, 0, 14, 0, 341, 327, 0, 2, 56, 76, 322, 347, 
    342, 0, 350, 276, 299, 317, 310, 307, 303, 300, 329, 305, 350, 112, 88, 
    0, 122, 116, 68, 107, 332, 330, 332, 354, 351, 102, 85, 309, 0, 304, 294, 
    294, 299, 303, 0, 26, 324, 313, 294, 299, 340, 54, 88, 281, 307, 311, 
    287, 290, 292, 308, 291, 286, 72, 18, 0, 308, 1, 63, 300, 292, 294, 287, 
    278, _, 263, 297, 284, 269, 276, 299, 300, 305, 286, 280, 297, 285, 283, 
    294, 273, 271, 269, 279, 295, 290, 278, 280, 286, 294, 293, 287, 284, 
    269, 278, 290, 286, 293, 296, 302, 291, 294, 292, 299, 310, 301, 308, 
    336, 337, 44, 75, 90, 78, 40, _, 266, 300, 311, _, 286, 349, 18, 317, 99, 
    315, 357, 337, 315, 301, 287, 336, 10, 63, 290, 333, 334, 0, _, 286, 303, 
    298, 332, 301, 328, 322, 336, 346, 353, 338, 288, 327, 332, 334, 355, 
    339, 334, 8, 327, 1, 1, 0, 300, 0, 17, _, 300, 304, 308, 320, 8, 313, 
    337, 61, 3, 43, 360, 0, 15, 309, 322, 0, 326, 31, 341, 331, 357, 33, _, 
    319, 305, _, 68, 299, 295, 301, 304, 306, 310, 309, 306, 302, 297, 305, 
    316, 316, 304, 303, 282, 288, _, 279, 300, 281, 276, _, _, _, _, 258, 
    243, 251, 262, 259, 252, 277, 280, 271, 274, 268, 284, 281, 271, 276, 
    258, 262, 251, 284, 289, 287, 296, 288, 294, 293, 298, 288, 323, 316, 
    315, 22, 120, 355, 147, 42, 55, 225, 357, 304, 0, 357, 288, 0, 358, _, 
    307, 304, 56, 52, 0, 3, 320, 315, 313, 303, 283, 287, 299, 300, 304, 307, 
    295, 302, _, 305, 308, 300, 303, 336, 302, 318, _, 321, 96, 8, 334, 0, 
    315, 0, 359, 359, 322, 323, 317, 313, 50, 6, 355, 103, 22, 93, 38, 349, 
    38, 333, 333, 311, 77, 70, 84, 85, 81, 84, 83, 319, 338, 355, 320, 4, 49, 
    343, 58, 353, 322, 291, 304, 360, 8, 358, 358, 355, 86, 54, 331, 306, 
    296, 327, 348, 341, 17, 59, 335, 357, 305, 53, 30, 6, 30, 289, 309, 295, 
    165, 66, 76, 86, 86, 92, 73, 81, 104, 70, 90, 92, 70, 87, 73, 80, 92, 86, 
    80, 84, 88, 85, _, 103, 79, 94, 92, 80, 81, 88, 92, 96, 99, 88, 89, 87, 
    68, 88, 96, 90, 68, 71, 56, 65, 60, 84, 70, _, 94, 81, 94, 116, 127, 83, 
    47, 66, 75, 67, 104, 73, 68, 21, 47, 46, 37, 330, _, 284, 311, _, 103, 
    95, 100, 100, 89, 98, 86, 92, 92, 71, 97, 102, 99, 107, 106, 96, 103, 
    294, 330, 321, _, 321, 306, 287, _, 303, 307, 309, 323, 285, 325, 328, 
    15, 313, 331, 298, 307, 25, 0, 352, 294, 320, 10, 319, 304, 260, 42, 1, 
    322, 314, 350, 5, 319, 315, 342, 331, 332, 348, 350, 330, 326, 356, 336, 
    334, 10, 21, 18, 358, 72, 49, 321, 300, 277, 277, 263, 280, 296, 334, 
    292, 309, 291, 348, 348, 296, 354, 58, 0, 339, 325, 0, 360, 3, 317, 328, 
    0, 324, 13, 10, 9, 339, 339, 346, 0, 344, 352, 0, 351, 333, 285, 298, 
    300, 303, 307, 0, 92, 0, 356, 348, 4, 360, 360, 322, 316, 315, 315, 283, 
    64, 0, 349, 327, 76, 77, 312, 325, 335, 344, 287, 33, 311, 358, 360, 347, 
    62, 0, 297, 289, 306, 316, 305, 300, 0, 9, 18, 360, 339, 298, 323, 302, 
    305, 329, 290, 296, 307, 319, 330, 342, 306, 297, 312, 303, 292, 302, 
    320, 318, 2, 63, 336, 43, 271, 250, 259, 273, 250, 240, 255, 266, 271, 
    263, 265, 237, 286, 283, 270, 233, 232, 229, 238, 256, 278, 212, 216, 
    255, 232, 240, 232, 270, 274, 285, 289, 289, 294, 288, 270, 268, 234, 
    243, 242, 247, 251, 262, 269, 285, 277, 266, 276, 270, 283, 277, 265, 
    269, 277, 297, 281, 282, _, 295, 289, 293, 285, 212, 318, 350, 259, 286, 
    355, 306, 332, 0, 347, 314, 328, 359, 7, 311, 310, 308, 312, 302, 313, 
    314, 301, 306, 310, 310, 308, _, 289, 309, 285, 281, 298, 315, 312, 311, 
    330, 317, 318, 315, 322, 309, 43, 317, 359, 337, _, 35, _, _, 322, 357, 
    4, 10, 48, 351, 294, 319, 50, 322, 301, 21, 309, 312, 287, 349, 307, 319, 
    _, 37, 70, 290, 49, 311, 328, _, 340, 83, _, 25, 358, 314, 296, 25, 0, 0, 
    0, 0, _, 2, 319, 133, 107, 15, 120, 91, 198, 62, 309, _, 62, 70, 51, 40, 
    77, 309, 13, 328, 344, 319, 296, 3, 3, 333, 312, 51, 354, 95, _, 328, _, 
    _, 333, 1, 319, 286, 293, 317, 316, 308, 323, 358, 37, 78, 74, 135, 126, 
    112, 74, 70, _, 258, 336, 58, 77, 215, 210, 207, 237, 266, 267, 268, 262, 
    280, 242, 244, 269, 247, 256, 257, 270, 282, 286, 290, 291, 307, 294, 4, 
    90, 324, 291, 322, 307, 351, 305, 64, 57, 61, 78, 82, 89, 82, 88, 92, 98, 
    123, 93, 79, 81, 71, _, 69, _, _, 276, 283, 276, 291, 292, 311, 307, 329, 
    338, 300, 0, 308, 307, 321, 6, 355, 302, _, _, 297, 290, 83, 307, 274, 
    310, 329, 316, 324, 93, 64, 3, 1, 40, 319, 319, 52, 74, 68, _, 81, 95, 
    72, 95, 88, 56, 80, 64, 73, 81, 73, 91, 95, 103, 106, 100, 90, 79, 85, 
    69, 81, 84, 88, 91, 125, 122, 89, 64, 53, _, 68, 62, 74, 58, 55, 49, 54, 
    46, 61, 58, 61, 60, 49, 59, 56, 110, 54, 63, 45, 57, 67, 43, _, 119, 103, 
    104, 80, 80, 48, 65, 112, 123, 122, 61, 73, 87, 122, 112, 104, 106, 95, 
    _, 114, 87, 77, 81, 295, 327, 328, 324, 316, 337, 7, 104, 0, 310, 9, 61, 
    87, 86, 86, 74, 38, 52, 358, 20, 267, 272, 314, 322, 7, _, 152, _, 70, 
    74, 65, 49, 60, 69, 105, 156, 106, 73, 55, 45, 64, 32, 87, 60, 52, 70, 
    83, 323, 300, 286, 301, 322, 324, 290, 24, 104, 65, 64, 69, 84, 82, 57, 
    96, 92, 57, 0, 318, 310, 305, 328, 326, 321, 354, 313, 322, 292, 335, 
    348, 305, 315, 346, 316, 323, 0, 307, 322, 272, 302, 256, 280, 21, 39, 
    15, 39, 35, 59, 15, 30, 45, 40, 23, 359, 196, 10, 15, 13, 10, 56, 47, 77, 
    95, 121, 198, 179, 63, 65, 45, 19, 320, 236, 235, 233, 306, 267, 198, 10, 
    18, 2, 3, 4, 15, 291, 344, 341, 313, 342, 252, 316, 334, 312, 13, 343, 
    322, 289, 348, 330, 304, 315, 321, 322, 308, 12, 333, 346, 327, 303, 313, 
    303, 319, 285, 304, 308, 297, 281, 291, 358, 43, 105, 136, 136, 135, 137, 
    121, 101, 89, 79, 97, 103, 110, 99, 99, 91, 83, 92, 96, 94, 99, 101, 98, 
    100, 97, 90, 80, 70, 83, 93, 95, 88, 95, 110, 99, 87, 89, 71, 64, 60, 29, 
    46, 44, 33, 50, 60, 67, 63, 25, 39, 62, 42, 60, 44, 56, 64, 65, 47, 60, 
    50, 42, 238, 357, 46, 44, 42, 54, 220, 53, 331, 332, 327, 301, 315, 314, 
    315, 314, 52, 332, 296, 302, 275, 290, 310, 317, 288, 322, 313, 307, 295, 
    352, 294, 315, 298, 298, 315, 291, 305, 297, 316, 349, 294, 337, 329, 
    355, 273, 299, 298, 326, 322, 313, 305, 321, 293, 317, 326, 275, 306, 96, 
    308, 297, 70, 341, 307, 322, 339, 356, 0, 337, 328, 27, 360, 21, 36, 17, 
    45, 36, 35, 42, 32, 40, 27, 12, 11, 16, 29, 37, 30, 28, 42, 29, 31, 45, 
    37, 16, 345, 332, 316, 345, 329, 37, 90, 42, 33, 25, 33, 39, 46, 48, 38, 
    40, 51, 28, 118, 303, 220, 202, 278, 327, 0, 341, 6, 304, 342, 281, 281, 
    313, 348, 349, 321, 51, 40, 38, 41, 353, 34, 36, 33, 36, 33, 34, 358, 16, 
    37, 32, 38, 29, 41, 27, 32, 41, 197, 324, 331, 300, 278, 236, 265, 304, 
    300, 283, 299, 307, 315, 297, 287, 278, 314, 311, 294, 288, 322, 311, 
    310, 302, 289, 282, 317, 305, 19, 310, 0, 316, 306, 306, 323, 342, 291, 
    31, 349, 2, 335, 304, 289, 302, 253, 10, 325, 322, 328, 313, 320, 286, 
    304, 298, 24, 29, 360, 310, 321, 4, 357, 333, 296, 312, 267, 295, 320, 
    338, 2, 347, 321, 309, 344, 323, 336, 314, 301, 329, 309, 318, 297, 333, 
    295, 349, 327, 312, 314, 313, 345, 322, 305, 311, 347, 335, 315, 309, 
    298, 314, 304, 318, 324, 320, 315, 326, 0, 321, 306, 13, 328, 341, 314, 
    325, 351, 328, 301, 315, 299, 301, 273, 312, 310, 323, 327, 318, 289, 
    312, 316, 297, 300, 317, 315, 316, 326, 324, 324, 305, 323, 313, 331, 
    305, 312, 328, 330, 316, 301, 325, 313, 300, 296, 315, 317, 330, 316, 
    318, 327, 338, 358, 352, 346, 324, 335, 318, 321, 313, 319, 312, 321, 
    332, 39, 335, 344, 348, 345, 344, 23, 0, 315, 294, 68, 323, 332, 328, 
    355, 322, 90, 46, 352, 52, 29, 359, 347, 301, 321, 330, 57, 3, 271, 327, 
    151, 314, 360, 29, 320, 304, 301, 293, 311, 307, 318, 338, 300, 350, 29, 
    45, 0, 325, 2, 326, 314, 315, 317, 292, 307, 299, 317, 312, 30, 317, 314, 
    95, 119, 310, 59, 342, 321, 359, 15, 68, 311, 342, 334, 31, 60, 31, 314, 
    340, 348, 337, 59, 333, 16, 334, 286, 286, 298, 304, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 295, 320, 300, 303, 329, 301, 316, 300, 293, 304, 295, 289, 300, 
    313, 291, 329, 292, 341, 313, 344, 333, 282, 324, 307, 2, 36, 90, 104, 
    93, 87, 76, 70, 55, 285, 280, 295, 285, 294, 286, 306, 305, 325, 284, 
    278, 273, 314, 302, 308, 286, 302, 304, 300, 360, 16, 5, 319, 297, 280, 
    326, 61, 74, 354, 312, 81, 72, 79, 92, 85, 83, 59, 0, 335, 303, 307, 230, 
    289, 315, 218, 41, 40, 39, 293, 306, 329, 342, 88, 314, 3, 113, 343, 350, 
    326, 341, 299, 85, 3, 330, 83, 60, 50, 347, 358, 107, 77, 175, 70, 59, 
    82, 82, 70, 101, 86, 76, 72, 65, 74, 76, 6, 352, 324, 313, 350, 341, 30, 
    344, _, _, 356, 300, 326, 317, 359, 315, 318, 350, 308, 326, 30, 309, 
    349, 232, _, 183, 291, 194, 235, 127, 9, 49, 328, 306, 56, 353, 328, 355, 
    324, 321, 337, 358, 341, 4, 334, 320, 15, 3, 320, _, 306, 288, 306, _, 
    354, 310, 310, 309, 350, 359, 341, 322, 298, 316, 311, 308, 304, 306, 
    315, 295, 350, 319, 128, 153, 210, 117, 33, 25, 335, 332, _, _, _, 46, 
    68, 72, 64, 62, 66, 52, 38, 37, 70, 32, 68, 96, 28, 183, 73, 109, 284, 
    296, 306, 303, 347, 329, 314, 294, 305, 296, 328, 16, 332, 297, 329, 332, 
    344, 315, 332, 307, 331, 84, 85, 97, 88, _, 87, 95, 91, 94, 94, 96, 96, 
    94, 94, 92, 96, 96, 87, 91, 94, 93, 94, 93, 94, 96, 94, 93, 89, _, 84, 
    81, 85, _, 80, 81, 82, 90, 78, 84, 96, 96, 95, 96, 85, 100, 100, 100, 98, 
    104, 114, 86, 96, 97, 102, 97, 90, 118, 83, 91, 71, 62, 65, 72, 64, 51, 
    62, 65, 65, 69, 68, 53, 47, 35, 26, 10, 51, _, 22, _, 63, 77, 66, 74, 61, 
    34, 68, 286, 73, 352, 43, 57, 41, 59, 33, 45, 40, 38, 344, 48, 35, 50, 
    42, 40, 54, _, 27, 343, 323, 291, 348, 37, 334, 55, 313, 70, 78, 86, 307, 
    47, 70, 82, 55, _, 335, 324, 321, 351, 286, 293, 77, 70, 85, 72, 79, 101, 
    86, 96, 135, 121, 105, 328, 3, 333, 27, 297, 324, 341, 298, _, 300, _, 
    326, 324, 319, 337, 326, 342, 13, 312, 34, 332, 343, 15, 334, 333, 317, 
    303, 313, 1, 319, 2, 348, 336, 323, 22, 343, _, _, 309, 324, 317, 334, 
    308, 348, 313, 333, 283, 301, 326, 308, 329, 202, 277, 204, 212, 221, 
    222, 205, 281, 291, 299, _, 285, 292, 305, 307, 309, 342, 339, 47, 3, 
    344, 351, 312, 323, 320, 73, 335, 327, 174, _, 35, _, _, 52, 53, 69, 87, 
    65, 78, 97, 57, 137, 123, 352, 44, 34, 39, 41, 38, 41, _, _, 42, 28, 32, 
    46, 33, 33, 15, _, 22, 284, 337, 277, 313, 322, 328, 151, 346, 351, 343, 
    _, 32, 25, 36, 41, 38, 40, 37, 33, 43, 26, 7, 359, 57, 353, 350, 352, 6, 
    32, 53, 38, 12, 10, 11, 23, 13, 6, 11, 11, 9, _, 356, 286, _, 349, 294, 
    287, 302, 310, 344, 293, 320, 258, 292, 320, 316, 276, 294, 292, 298, 
    309, _, _, 310, 306, 298, 304, 304, _, 304, 309, 311, 308, 18, 358, 28, 
    65, 0, 79, 22, 349, 342, _, 311, 338, 297, 313, 326, 350, _, 337, 313, 
    340, 314, 295, 302, 318, 352, 357, 312, 264, 317, 3, 109, 0, 250, 4, 302, 
    18, 307, 326, 333, _, 300, 333, _, 311, 312, 310, 311, 305, 35, 302, 312, 
    303, 324, 335, 336, 308, 348, 303, 340, 334, _, _, 240, 8, 340, 352, 336, 
    _, 350, 29, 323, 219, 315, 51, 180, 191, 186, 296, 305, _, 339, _, 338, 
    _, 304, 300, 287, 296, 8, 56, 21, 319, 317, 334, 317, 316, 6, 355, 15, 
    317, 334, 313, 356, 346, 20, 346, 306, 333, 7, 325, 325, _, 349, 291, _, 
    291, 5, 299, 316, 317, 344, 34, 312, 268, 304, 310, 322, 338, 325, 312, 
    293, 311, 6, _, 183, 183, 181, 356, 36, 287, 202, 259, 301, 274, 235, 
    216, 265, 213, 215, 249, 237, _, 251, _, 269, 285, 280, 279, 269, 268, 
    303, 273, 278, 284, 299, 291, 300, 296, 312, 317, 325, 321, 294, 345, 34, 
    341, 333, 333, 353, 310, 309, 318, 2, _, 309, 69, 46, 296, 259, 28, 341, 
    341, 335, 319, 315, 315, 295, 301, 326, 305, 315, 324, 308, 320, 322, 
    303, 22, 21, 15, 322, 308, 309, 292, 294, 330, 331, 315, 300, 317, 304, 
    312, 323, 293, 21, 301, _, 301, 331, 344, 326, 318, 338, 332, 323, 319, 
    328, 324, 319, 307, 304, 342, 329, 312, 315, 327, 309, 301, 320, 307, 
    312, 285, 96, 247, 268, 320, _, 277, 94, 90, 349, 9, 31, 41, 31, 34, 47, 
    275, 349, 320, 79, 53, 358, 348, 339, 359, 7, 303, 316, _, 347, 1, 358, 
    29, 6, 346, 343, 353, 324, 332, 309, 292, 308, 12, 307, 337, 13, 329, _, 
    349, 314, 345, 335, 47, 326, 2, 347, 33, 37, 341, 78, 29, 342, 4, 13, 0, 
    327, 320, 46, 6, 335, 35, 21, 359, 328, 5, 103, 68, _, 345, 68, 83, 307, 
    115, 16, 60, 59, 39, 34, 43, 35, 20, 35, 36, 39, 25, 31, 19, 13, _, 29, 
    16, 11, 12, 22, 16, 12, 15, 16, 16, 25, 17, 10, 10, 15, 16, 25, 38, 3, 
    359, _, 33, 27, 34, 223, 29, _, 310, 329, 320, 307, 315, 252, 318, 309, 
    300, 14, 260, 272, 309, 337, 283, 302, 305, 321, 298, 298, 359, 303, 322, 
    _, 337, 6, 24, 19, 10, 36, 10, 177, 110, 317, 310, 311, 308, 345, 273, 
    331, 296, 312, 304, 317, _, _, 306, 356, 328, 356, 353, 325, 345, 336, 0, 
    303, 318, 320, 321, 319, 305, 348, 337, 43, 105, 12, 302, _, 295, 355, 6, 
    _, 38, 15, 24, 356, 14, 345, 169, 353, 287, 249, 63, 309, 302, 297, 324, 
    56, 49, 49, 299, 322, 327, 28, 338, _, 139, 338, 30, 45, 41, 20, 197, 
    306, 323, 350, 360, 1, 3, 12, 15, 18, 9, 288, 300, 298, 315, 347, _, 54, 
    304, 270, 20, 61, 37, 298, 319, 350, 330, 325, 324, 324, 311, 286, 311, 
    324, 318, 317, 3, 300, 302, 313, 349, 327, 305, 2, 312, 47, 344, 315, 55, 
    77, 1, 50, 54, 331, 351, 60, 302, 41, 345, 334, 305, 299, 35, 308, 305, 
    313, 321, 335, 353, 70, 33, 24, 318, 332, 11, 333, 356, 313, 341, 20, 
    307, 298, 315, 314, 306, 322, _, _, _, 308, 292, 316, 319, 278, 302, 290, 
    307, 304, 307, 113, 82, 40, 94, 24, 327, 334, 196, 72, 288, 357, 3, 333, 
    352, _, _, 306, 304, 360, 20, 82, 79, 344, 145, 30, 0, 0, 308, 345, 89, 
    81, 95, 304, 293, 299, 258, _, 270, 299, 299, 304, 277, 305, 275, 301, 
    300, 304, 303, 310, 285, 300, 299, 302, 301, 323, 56, 239, 286, 285, 294, 
    _, _, 292, 300, 301, 240, 296, 298, 301, 282, 287, 298, 272, 269, 271, 
    268, 274, 283, 275, 268, 292, 286, 289, 289, 282, 300, _, 270, 263, 261, 
    262, 245, 275, 248, 273, 288, 281, 300, 303, 299, 306, 305, 311, 289, 
    305, _, 303, 305, 302, 286, 295, 305, 321, 298, 307, 303, 315, 317, 287, 
    305, 299, 282, 297, 288, 300, 317, 297, 294, 291, 300, 298, 276, _, 314, 
    304, 308, 288, 279, 281, 283, 305, 284, 284, 283, 302, 302, 301, 310, 
    313, 315, 261, 291, 291, 286, 261, 265, 294, 273, 292, 275, 254, 261, 
    256, 298, 253, 228, 257, 263, 251, 265, 271, 270, 286, 246, 264, 268, 
    272, _, 267, 267, _, 263, 267, 283, 290, 286, 286, 297, 295, 300, 292, 
    303, 290, 259, 222, 83, 90, 79, 294, 336, 75, 51, 18, _, _, 355, 356, 
    121, 102, 61, 8, 129, 48, 59, 15, 132, 39, 41, 326, 64, 1, 76, 53, 35, 
    34, 37, 35, 35, 42, 43, 45, 43, 45, 26, 19, 9, 7, 360, 315, 297, 270, 52, 
    32, 324, 24, 18, 292, 301, 275, 300, 307, 279, 305, 314, 52, 271, 278, 
    308, 299, 296, 296, 284, 355, 300, 334, 313, 69, 317, 321, 315, 304, 8, 
    331, 73, 47, 45, 40, 37, 33, 37, 32, 39, 37, 32, 39, 46, 38, 44, 22, 29, 
    30, 359, 36, 166, 289, 238, 288, 149, 359, 262, 275, 65, 357, 280, 279, 
    298, 317, 342, 54, 272, 297, 207, 292, 341, 352, 308, 282, 300, 306, 296, 
    295, 300, 311, 11, 179, 41, 346, 318, 327, 324, 339, 290, 354, 284, 308, 
    345, 314, 301, 300, 313, 331, 309, 307, 325, 270, 299, 315, 314, 320, 
    330, 335, 310, 303, 276, 297, 289, 283, 55, 333, 309, 0, 325, 33, 298, 
    347, 296, 332, 70, 65, 64, 60, 39, 36, 32, 35, 33, 35, 47, 45, 55, 36, 
    40, 49, 39, 30, 38, 35, 1, 60, 240, 4, 206, 230, 200, 167, 41, 49, 62, 
    78, 71, 73, 76, 78, 94, 83, 80, 91, 93, 90, 92, 99, 98, 103, 95, 93, 88, 
    85, 82, 73, 83, 80, 75, 74, 62, 69, 55, 73, 88, 61, 84, 62, 73, 69, 71, 
    48, 48, 57, 269, 35, 104, 101, 83, 52, 249, 329, 37, 20, 7, 1, 353, 352, 
    350, 55, 31, 283, 340, 288, 317, 340, 345, 304, 219, 314, 300, 291, 295, 
    298, 348, 9, 295, 291, 304, 20, 36, 189, 181, 165, 129, 80, 87, 74, 323, 
    23, 23, 336, 2, 9, 5, 48, 41, 35, 27, 33, 33, 32, 32, 17, 79, 132, 240, 
    255, 328, 322, 261, 204, 200, 360, 185, 234, 303, 202, 254, 346, 77, 178, 
    85, 275, 176, 328, 307, 219, 133, 258, 204, 329, 358, 329, 342, 317, 297, 
    41, 331, 307, 298, 313, 319, 13, 360, 357, 319, 320, 319, 306, 327, 321, 
    320, 316, 321, 316, 295, 338, 312, 358, 350, 332, 353, 340, 320, 311, 
    315, 318, 312, 316, 260, 316, 320, 350, 10, 345, 9, 309, 23, 310, 35, 
    347, 298, 358, 336, 353, 330, 322, 20, 18, 354, 341, 339, 344, 53, 13, 
    299, 0, 12, 318, 358, 354, 25, 285, 352, 3, 1, 298, 35, 298, 85, 324, 
    317, 328, 282, 353, 360, 4, 360, 360, 0, 338, 37, 323, 325, 353, 351, 1, 
    349, 321, 357, 339, 319, 35, 340, 36, 66, 360, 305, 354, 68, 336, 317, 0, 
    0, 0, 332, 317, 338, 356, 339, 311, 328, 354, 2, 336, 8, 318, 320, 344, 
    317, 315, 314, 39, 0, 76, 89, 320, 318, 85, 327, 335, 28, 347, 0, 26, 
    360, 326, 273, 123, 316, 310, 306, 96, 322, 68, 343, 0, 360, 316, 360, 
    46, 0, 316, 53, 333, 104, 345, 340, 24, 332, 327, 315, 322, 341, 49, 315, 
    0, 360, 360, 350, 346, 5, 323, 318, 325, 300, 214, 236, 53, 100, 178, 19, 
    254, 161, 72, 8, 334, 4, 309, 360, 28, 78, 36, 0, 16, 326, 326, 326, 307, 
    317, 332, 289, 299, 354, 326, 82, 327, 329, 3, 112, 350, 306, 287, 92, 0, 
    352, 313, 3, 339, 360, 65, _, 1, 0, 355, 0, 310, 26, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 302, 307, 305, 296, 328, 360, 39, 38, 41, 12, 19, 
    24, 306, 309, 320, 30, 25, 46, 56, 60, 71, 69, 63, 65, 70, 71, 70, 66, 
    72, 64, 330, 301, 288, 297, 337, 279, 306, 298, 320, 296, 327, 304, 301, 
    284, 0, 255, 0, 65, 3, 40, 77, 46, 32, 44, 27, 15, 58, 326, 360, 19, 23, 
    143, 47, 42, 26, 51, 39, 2, 58, 59, 356, 300, 285, 291, 313, 45, 46, 50, 
    52, 59, 68, 58, 292, 299, 303, 181, 342, 33, 327, 185, 58, 360, 338, 138, 
    350, 177, 325, 328, 330, 351, 172, 31, 314, 315, 298, 18, 309, 337, 315, 
    306, 293, 298, 304, 318, 60, 351, 66, 357, 312, 77, 316, 320, 328, 26, 
    316, 303, 47, 72, 47, 0, 41, 357, 356, 356, 0, 67, 353, 71, 14, 307, 2, 
    70, 40, 360, 323, 106, 319, 128, 79, 290, 309, 290, 80, 323, 329, 300, 
    296, 260, 325, 33, 62, 355, 47, 360, 357, 355, 344, 313, 340, 201, 110, 
    109, 43, 103, 106, 340, 37, 27, 11, 33, 16, 13, 15, 15, 20, 34, 27, 29, 
    28, 27, 32, 30, 30, 28, 26, 33, 27, 36, 33, 34, 34, 33, 34, 34, 32, 33, 
    35, 38, 28, 42, 40, 37, 39, 38, 36, 35, 33, 32, 36, 37, 44, 41, 41, 44, 
    24, 32, 36, 51, 26, 44, 5, 40, 11, 47, 24, 360, 349, 55, 14, 351, 16, 
    334, 325, 325, 160, 245, 106, 70, 0, 311, 330, 342, 313, 310, 0, 359, 0, 
    0, 340, 2, 328, 328, 41, 315, 342, 330, 324, 0, 313, 331, 300, 312, 316, 
    274, 349, 0, 28, 301, 342, 329, 335, 328, 316, 317, 333, 344, 360, 81, 
    360, 357, 342, 320, 341, 320, 348, 360, 5, 49, 0, 1, 52, 49, 4, 22, 26, 
    315, 15, 10, 5, 319, 360, 50, 329, 320, 320, 0, 20, 348, 0, 5, 81, 343, 
    347, 7, 15, 54, 38, 7, 351, 321, 336, 337, 353, 351, 358, 300, 328, 330, 
    332, 12, 345, 352, 349, 13, 1, 307, 80, 76, 127, 130, 86, 107, 324, 282, 
    17, 8, 315, 59, 360, 300, 310, 357, 114, 326, 317, 298, 328, 56, 303, 
    306, 304, 268, 289, 283, 310, 302, 313, 311, 302, 205, 203, 210, 360, 
    347, 320, 32, 41, 3, 331, 284, 345, 0, 326, 88, 184, 300, 324, 234, 45, 
    351, 70, 57, 178, 80, 36, 24, 329, 82, 24, 30, 32, 358, 94, 26, 319, 332, 
    108, 75, 81, 83, 78, 80, 51, 69, 54, 64, 37, 42, 43, 45, 40, 39, 40, 44, 
    42, 46, 211, 260, 220, 192, 55, 280, 235, 100, 103, 227, 101, 55, 73, 
    121, 188, 229, 300, 341, 182, 64, 117, 80, 78, 79, 80, 80, 143, 161, 268, 
    256, 283, 145, 224, 194, 78, 23, 176, 191, 198, 35, 174, 221, 190, 342, 
    10, 8, 7, 45, 285, 82, 81, 338, 8, 25, 198, 347, 40, 78, 59, 262, 252, 
    88, 353, 20, 360, 311, 309, 320, 300, 293, 278, 311, 275, 296, 307, 315, 
    13, 343, 188, 14, 339, 33, 330, 308, 318, 336, 0, 357, 349, 344, 329, 
    335, 336, 309, 340, 342, 360, 94, 359, 353, 330, 290, 292, 351, 301, 311, 
    311, 334, 321, 355, 0, 340, 360, 352, 37, 7, 322, 100, 0, 347, 338, 292, 
    255, 311, 95, 310, 291, 294, 76, 302, 198, 312, 145, 335, 339, 143, 130, 
    329, 26, 325, 300, 288, 317, 342, 294, 318, 277, 265, 303, 40, 327, 322, 
    322, 292, 343, 337, 289, 343, 360, 8, 328, 3, 56, 308, 329, 98, 0, 116, 
    291, 331, 77, 307, 268, 324, 110, 13, 334, 327, 342, 71, 354, 326, 0, 
    113, 38, 48, 1, 50, 82, 331, 140, 10, 304, 300, 164, 270, 207, 18, 24, 
    26, 144, 332, 240, 224, 267, 246, 355, 344, 346, 330, 17, 20, 90, 92, 
    116, 87, 333, 151, 164, 212, 237, 223, 190, 277, 326, 319, 288, 8, 356, 
    112, 131, 176, 84, 100, 175, 282, 22, 65, 56, 69, 69, 48, 42, 61, 95, 89, 
    78, 85, 75, 76, 339, 350, 347, 309, 38, 234, 300, 324, 325, 330, 314, 
    322, 316, 325, 118, 133, 14, 107, 126, 115, 91, 296, 311, 283, 334, 311, 
    307, 337, 308, 283, 290, 308, 305, 300, 298, 322, 291, 338, 288, 17, 250, 
    347, 109, 66, 312, 74, 334, 46, 0, 88, 356, 6, 324, 17, 327, 360, 61, 0, 
    21, 35, 135, 350, 0, 340, 356, 343, 74, 328, 343, 0, 91, 282, 359, 352, 
    284, 308, 123, 67, 360, 334, 345, 340, 332, 348, 311, 326, 329, 81, 71, 
    75, 74, 77, 80, 83, 75, 78, 77, 81, 74, 86, 103, 76, 91, 100, 5, 3, 40, 
    72, 61, 73, 125, 68, 96, 287, 311, 312, 291, 310, 321, 329, 313, 90, 355, 
    13, 348, 305, 99, 200, 292, 322, 106, 104, 343, 321, 108, 79, 0, 114, 90, 
    72, 309, 114, 344, 358, 19, 346, 5, 342, 15, 13, 360, 315, 347, 335, 331, 
    340, 313, 62, 73, 27, 332, 4, 103, 291, 34, 351, 18, 37, 311, 1, 0, 0, 0, 
    334, 353, 334, 343, 90, 360, 350, 0, 98, 92, 308, 0, 0, 93, 317, 322, 
    356, 295, 315, 359, 294, 299, 328, 89, 358, 319, 320, 344, 357, 108, 356, 
    300, 257, 283, 220, 210, 50, 220, 233, 317, 276, 328, 337, 312, 324, 314, 
    35, 38, 355, 350, 340, 101, 248, 197, 24, 122, 123, 126, 162, 5, 247, 
    110, 204, 83, 77, 96, 317, 11, 293, 123, 25, 274, 39, 13, 322, 103, 351, 
    20, 32, 300, 350, 28, 74, 85, 81, 216, 337, 346, 67, 344, 355, 105, 4, 4, 
    357, 0, 8, 339, 100, 82, 100, 322, 38, 0, 358, 287, 295, 306, 301, 320, 
    333, 297, 323, 306, 285, 312, 84, 73, 113, 193, 310, 311, 320, 317, 306, 
    345, 91, 115, 200, 262, 282, 270, 296, 277, 264, 16, 47, 31, 64, 51, 51, 
    8, 1, 44, 14, 311, 308, 293, 60, 360, 2, 311, 271, 270, 276, 274, 272, 
    270, 272, 304, 65, 300, 66, 19, 318, 304, 80, 315, 339, 340, 320, 319, 
    108, 85, 63, 302, 284, 276, 276, 305, 326, 335, 82, 46, 66, 53, 45, 52, 
    58, 53, 70, 80, 87, 50, 45, 56, 45, 47, 37, 68, 50, 13, 52, 14, 12, 32, 
    42, 57, 38, 48, 61, 50, 337, 31, 39, 102, 331, 335, 68, 330, 301, 360, 
    88, 111, 275, 282, 275, 278, 265, 228, 170, 144, 328, 228, 347, 346, 47, 
    65, 53, 235, 360, 3, 40, 43, 56, 48, 86, 59, 48, 249, 158, 43, 204, 27, 
    27, 223, 143, 256, 82, 18, 348, 289, 147, 120, 112, 60, 31, 345, 336, 
    320, 157, 159, 346, 174, 153, 82, 103, 105, 179, 81, 107, 265, 1, 0, 3, 
    0, 341, 327, 351, 0, 0, 0, 348, 360, 18, 300, 298, 247, 309, 225, 228, 
    230, 270, 274, 277, 291, 0, 360, 353, 0, 0, 57, 360, 318, 342, 41, 130, 
    275, 274, 273, 270, 272, 267, 277, 237, 321, 133, 295, 272, 265, 280, 
    260, 272, 17, 325, 299, 304, 300, 300, 301, 306, 115, 117, 130, 20, 290, 
    286, 257, 7, 115, 336, 355, 95, 360, 336, 12, 317, 346, 80, 77, 241, 261, 
    232, 245, 18, 20, 100, 280, 268, 277, 271, 286, 320, 306, 316, 88, 343, 
    104, 315, 305, 291, 297, 298, 300, 301, 301, 308, 289, 288, 292, 285, 
    290, 281, 266, 292, 267, 114, 113, 120, 131, 277, 290, 316, 308, 317, 0, 
    113, 336, 132, 150, 251, 300, 291, 302, 286, 311, 322, 241, 124, 166, 
    242, 283, 263, 76, 152, 292, 275, 310, 272, 131, 100, 87, 73, 105, 292, 
    300, 322, 300, 275, 345, 344, 229, 124, 120, 130, 155, 276, 16, 0, 34, 0, 
    317, 210, 259, 326, 295, 290, 282, 322, 225, 185, 152, 235, 295, 250, 
    254, 259, 237, 222, 235, 223, 229, 212, 281, 185, 251, 161, 307, 285, 63, 
    114, 300, 326, 303, 322, 124, 117, 278, 282, 286, 279, 280, 342, 105, 
    104, 75, 308, 314, 272, 49, 297, 212, 300, 334, 320, 319, 1, 287, 349, 
    137, 164, 148, 186, 215, 291, 90, 63, 59, 13, 239, 31, 15, 25, 6, 360, 
    221, 8, 8, 340, 31, 35, 40, 58, 36, 184, 52, 99, 273, 262, 118, 29, 58, 
    26, 87, 111, 102, 45, 358, 3, 55, 341, 18, 302, 360, 70, 277, 65, 98, 
    121, 75, 60, 37, 56, 45, 77, 269, 197, 16, 259, 26, 30, 26, 249, 89, 50, 
    32, 52, 40, 294, 356, 24, 91, 258, 253, 73, 63, 94, 127, 100, 299, 268, 
    333, 241, 270, 57, 267, 335, 335, 33, 358, 65, 54, 54, 53, 53, 187, 107, 
    102, 90, 174, 106, 88, 65, 110, 78, 79, 37, 76, 88, 3, 65, 341, 90, 2, 
    323, 360, 26, 133, 148, 147, 241, 164, 174, 122, 142, 144, 212, 171, 179, 
    153, 187, 168, 294, 183, 268, 120, 250, 258, 258, 186, 224, 230, 252, 
    180, 237, 200, 179, 201, 84, 213, 183, 225, 189, 210, 262, 189, 156, 318, 
    113, 309, 21, 358, 298, 100, 60, 360, 324, 181, 166, 131, 222, 176, 259, 
    235, 256, 293, 290, 290, 297, 291, 291, 292, 289, 138, 340, 340, 302, 
    280, 263, 278, 273, 259, 248, 229, 162, 180, 160, 146, 109, 147, 153, 
    139, 239, 233, 286, 280, 286, 286, 300, 308, 29, 0, 271, 106, 267, 155, 
    15, 260, 257, 179, 155, 147, 175, 152, 122, 110, 115, 280, 288, 98, 359, 
    280, 128, 31, 1, 27, 146, 200, 262, 270, 268, 276, 265, 183, 140, 279, 
    126, 99, 188, 171, 184, 330, 309, 289, 290, 118, 92, 87, 291, 290, 288, 
    278, 287, 271, 277, 270, 277, 272, 268, 295, 269, 90, 263, 177, 298, 269, 
    294, 312, 310, 321, 330, 357, 3, 327, 315, 133, 331, 252, 265, 270, 278, 
    205, 202, 148, 129, 85, 224, 290, 91, 315, 255, 242, 118, 253, 278, 353, 
    300, 286, 258, 322, 235, 30, 50, 66, 259, 257, 226, 289, 220, 237, 303, 
    142, 150, 223, 241, 130, 123, 171, 150, 157, 165, 200, 287, 284, 284, 
    284, 264, 262, 200, 181, 151, 134, 125, 132, 165, 116, 126, 102, 123, 
    120, 132, 187, 100, 80, 78, 11, 279, 252, 270, 262, 137, 141, 126, 150, 
    164, 157, 192, 138, 139, 175, 354, 149, 139, 263, 273, 254, 106, 0, 320, 
    310, 269, 133, 154, 268, 277, 162, 161, 162, 147, 138, 155, 271, 292, 
    293, 275, 283, 287, 104, 91, 197, 0, 9, 317, 360, 57, 280, 18, 292, 333, 
    154, 354, 139, 128, 0, 296, 307, 300, 257, 6, 200, 47, 256, 250, 244, 
    131, 279, 255, 32, 43, 28, 67, 74, 61, 10, 9, 44, 55, 51, 20, 75, 81, 
    105, 55, 76, 88, 48, 309, 267, 272, 337, 360, 32, 90, 112, 67, 80, 60, 
    62, 65, 39, 67, 42, 40, 34, 49, 48, 325, 10, 29, 119, 273, 296, 225, 343, 
    278, 250, 232, 237, 36, 153, 180, 199, 177, 209, 146, 155, 195, 154, 114, 
    76, 126, 57, 70, 314, 19, 312, 53, 116, 123, 129, 97, 129, 93, 95, 86, 
    255, 116, 89, 158, 187, 120, 218, 155, 209, 198, 288, 243, 178, 300, 289, 
    277, 290, 282, 280, 278, 276, 247, 233, 134, 177, 158, 134, 294, 280, 
    321, 272, 269, 295, 49, 65, 100, 273, 200, 179, 300, 149, 11, 260, 265, 
    272, 248, 277, 260, 264, 194, 232, 135, 174, 148, 175, 151, 126, 69, 36, 
    233, 296, 257, 195, 220, 254, 268, 245, 220, 96, 103, 146, 139, 126, 112, 
    107, 108, 47, 88, 91, 66, 61, 66, 15, 44, 33, 304, 347, 52, 273, 328, 
    310, 306, 239, 34, 81, 198, 185, 191, 353, 314, 351, 21, 18, 325, 360, 7, 
    21, 141, 48, 20, 9, 38, 360, 351, 300, 265, 110, 351, 13, 333, 355, 79, 
    16, 45, 95, 39, 33, 106, 51, 88, 290, 121, 41, 28, 23, 40, 63, 50, 51, 
    12, 199, 252, 82, 241, 187, 29, 286, 195, 197, 226, 170, 245, 262, 225, 
    48, 148, 2, 119, 136, 332, 110, 69, 200, 283, 295, 168, 130, 172, 173, 
    139, 166, 150, 162, 166, 166, 163, 159, 136, 127, 135, 0, 0, 83, 316, 
    360, 8, 306, 33, 138, 113, 153, 171, 172, 163, 164, 167, 139, 149, 167, 
    150, 180, 145, 159, 175, 167, 253, 221, 208, 208, 120, 118, 141, 164, 
    176, 170, 152, 167, 144, 156, 174, 163, 176, 170, 176, 171, 156, 177, 
    144, 158, 157, 89, 141, 80, 99, 100, 306, 304, 356, 139, 162, 154, 176, 
    169, 141, 126, 106, 146, 175, 209, 278, 12, 247, 68, 40, 26, 16, 20, 112, 
    308, 259, 130, 253, 258, 187, 269, 147, 216, 156, 201, 246, 174, 177, 
    174, 144, 115, 346, 77, 1, 355, 341, 45, 46, 46, 73, 127, 140, 110, 155, 
    105, 112, 92, 99, 113, 89, 98, 71, 148, 95, 305, 303, 311, 183, 349, 316, 
    80, 124, 20, 17, 99, 306, 160, 243, 131, 130, 160, 162, 101, 112, 62, 
    121, 98, 124, 116, 120, 140, 135, 133, 321, 265, 0, 134, 11, 348, 191, 
    158, 275, 270, 275, 262, 231, 166, 159, 155, 129, 155, 157, 249, 83, 89, 
    52, 308, 52, 333, 360, 7, 31, 133, 113, 123, 139, 131, 131, 150, 147, 
    125, 158, 132, 124, 137, 147, 114, 132, 161, 89, 327, 128, 341, 97, 358, 
    355, 119, 9, 63, 70, 142, 149, 175, 119, 127, 51, 0, 348, 260, 124, 54, 
    60, 110, 120, 355, 350, 340, 90, 119, 162, 140, 139, 137, 135, 132, 124, 
    133, 153, 127, 153, 162, 124, 139, 166, 120, 124, 22, 129, 87, 89, 0, 
    351, 127, 127, 130, 131, 119, 129, 166, 151, 152, 145, 141, 152, 149, 
    173, 204, 245, 187, 292, 291, 57, 81, 349, 291, 155, 195, 286, 291, 92, 
    185, 127, 147, 137, 156, 179, 173, 147, 165, 169, 174, 178, 127, 360, 
    347, 119, 125, 360, 314, 292, 181, 169, 170, 177, 152, 180, 138, 82, 98, 
    120, 130, 172, 166, 202, 197, 231, 177, 208, 195, 231, 1, 139, 0, 222, 
    350, 360, 146, 343, 237, 186, 184, 143, 120, 140, 140, 109, 54, 111, 86, 
    97, 95, 83, 102, 151, 181, 288, 290, 291, 144, 111, 111, 316, 94, 163, 0, 
    321, 130, 278, 204, 86, 302, 116, 111, 172, 326, 267, 164, 235, 305, 137, 
    38, 167, 184, 340, 119, 274, 91, 81, 106, 135, 148, 164, 173, 148, 83, 
    275, 284, 219, 244, 184, 173, 173, 156, 131, 176, 172, 156, 153, 149, 
    144, 134, 133, 132, 127, 134, 123, 136, 154, 133, 135, 138, 135, 130, 
    112, 127, 355, 357, 331, 330, 63, 132, 170, 177, 228, 136, 152, 89, 138, 
    265, 294, 283, 118, 94, 131, 102, 165, 154, 172, 162, 100, 84, 288, 286, 
    278, 113, 110, 100, 34, 83, 106, 156, 170, 92, 90, 143, 154, 51, 115, 
    134, 46, 85, 115, 111, 130, 78, 112, 151, 96, 88, 100, 157, 80, 129, 158, 
    155, 169, 149, 144, 159, 168, 160, 114, 159, 180, 121, 136, 98, 278, 287, 
    299, 296, 290, 283, 267, 266, 289, 255, 264, 166, 174, 168, 31, 118, 133, 
    183, 177, 179, 176, 175, 169, 102, 104, 84, 233, 150, 190, 75, 54, 80, 
    67, 71, 120, 130, 80, 72, 139, 102, 140, 162, 156, 48, 130, 100, 74, 59, 
    39, 277, 190, 125, 219, 227, 294, 284, 254, 264, 292, 330, 103, 268, 112, 
    80, 72, 32, 208, 169, 170, 170, 147, 100, 77, 146, 124, 126, 82, 163, 
    108, 134, 146, 161, 166, 172, 201, 235, 178, 179, 173, 324, 186, 126, 
    173, 171, 176, 181, 198, 268, 296, 295, 291, 294, 313, 265, 266, 283, 
    270, 180, 172, 291, 287, 290, 272, 274, 275, 286, 286, 290, 299, 309, 
    311, 288, 296, 295, 298, 299, 292, 289, 296, 299, 299, 279, 257, 278, 
    286, 274, 269, 280, 284, 304, 307, 163, 191, 306, 287, 286, 87, 294, 298, 
    272, 254, 102, 119, 109, 157, 106, 167, 170, 139, 167, 141, 135, 110, 
    112, 352, 321, 297, 287, 290, 291, 302, 275, 305, 298, 297, 311, 294, 
    296, 298, 175, 231, 243, 288, 245, 112, 88, 70, 94, 83, 100, 122, 101, 
    126, 90, 164, 137, 155, 130, 124, 127, 145, 130, 94, 62, 138, 156, 172, 
    163, 89, 112, 60, 71, 55, 60, 100, 126, 62, 100, 167, 185, 19, 31, 12, 
    28, 355, 92, 88, 79, 80, 210, 70, 74, 86, 80, 76, 94, 106, 101, 80, 152, 
    153, 154, 190, 160, 139, 143, 159, 138, 140, 141, 143, 170, 282, 151, 
    160, 127, 115, 117, 111, 115, 99, 97, 97, 97, 96, 94, 94, 98, 94, 112, 
    117, 119, 120, 108, 108, 109, 103, 109, 113, 114, 114, 109, 104, 107, 96, 
    118, 117, 125, 127, 127, 127, 116, 111, 118, 114, 88, 171, 156, 151, 129, 
    155, 150, 139, 157, 138, 134, 174, 175, 177, 177, 64, 0, 100, 117, 103, 
    69, 35, 357, 269, 102, 71, 216, 267, 257, 254, 269, 263, 269, 275, 264, 
    265, 276, 266, 266, 269, 271, 265, 263, 277, 275, 278, 282, 279, 274, 
    264, 254, 259, 247, 235, 238, 235, 235, 246, 281, 257, 249, 254, 257, 
    255, 274, 292, 292, 295, 295, 294, 282, 289, 291, 284, 294, 281, 288, 
    172, 166, 174, 168, 170, 164, 140, 151, 140, 120, 143, 148, 135, 130, 
    127, 92, 117, 57, 124, 124, 21, 94, 288, 288, 287, 260, 288, 265, 271, 
    268, 286, 271, 285, 285, 286, 277, 115, 96, 131, 119, 156, 73, 118, 72, 
    76, 111, 157, 146, 131, 136, 137, 145, 137, 137, 154, 159, 156, 159, 144, 
    113, 139, 100, 88, 129, 160, 100, 158, 135, 141, 129, 136, 143, 142, 157, 
    154, 152, 144, 155, 146, 142, 160, 148, 132, 131, 110, 101, 75, 89, 114, 
    166, 166, 154, 158, 155, 160, 164, 164, 166, 168, 167, 163, 155, 164, 
    163, 139, 140, 162, 144, 160, 162, 113, 89, 124, 150, 160, 171, 150, 130, 
    133, 129, 134, 119, 163, 133, 161, 147, 137, 150, 169, 162, 137, 102, 
    114, 114, 114, 95, 140, 176, 177, 179, 154, 128, 175, 19, 354, 140, 106, 
    160, 132, 130, 117, 38, 111, 141, 126, 276, 270, 268, 271, 283, 279, 285, 
    286, 266, 271, 272, 262, 272, 264, 274, 269, 269, 279, 272, 260, 262, 
    268, 260, 251, 286, 291, 286, 305, 300, 313, 320, 315, 299, 296, 173, 
    127, 109, 123, 140, 118, 128, 130, 99, 133, 128, 338, 125, 1, 125, 342, 
    300, 102, 346, 347, 334, 101, 263, 78, 115, 91, 97, 92, 90, 92, 203, 103, 
    164, 140, 45, 273, 292, 300, 293, 300, 332, 278, 87, 333, 117, 83, 91, 
    75, 86, 86, 40, 107, 110, 142, 133, 134, 173, 168, 168, 208, 339, 297, 
    312, 314, 308, 57, 79, 346, 344, 61, 96, 107, 125, 132, 131, 125, 144, 
    279, 298, 52, 322, 316, 113, 316, 0, 340, 339, 105, 332, 99, 100, 116, 
    125, 124, 134, 120, 105, 128, 106, 140, 142, 159, 105, 131, 142, 120, 80, 
    319, 298, 303, 304, 310, 316, 308, 200, 188, 177, 134, 162, 100, 91, 135, 
    144, 265, 25, 56, 161, 157, 0, 1, 303, 107, 110, 294, 308, 286, 286, 270, 
    299, 278, 300, 315, 304, 303, 273, 253, 294, 289, 295, 280, 258, 250, 
    125, 285, 177, 300, 190, 193, 261, 328, 319, 322, 311, 299, 317, 1, 107, 
    122, 92, 137, 140, 112, 116, 175, 173, 166, 161, 166, 170, 281, 286, 291, 
    303, 291, 279, 267, 270, 265, 273, 246, 248, 265, 245, 260, 265, 267, 
    229, 176, 176, 195, 183, 248, 220, 172, 164, 156, 158, 175, 175, 132, 63, 
    142, 131, 132, 142, 153, 55, 165, 152, 148, 141, 132, 121, 127, 141, 169, 
    153, 162, 171, 133, 130, 97, 117, 99, 93, 20, 67, 101, 89, 76, 80, 61, 
    160, 135, 147, 132, 165, 142, 142, 129, 147, 164, 120, 117, 114, 71, 105, 
    100, 109, 119, 121, 116, 87, 82, 142, 119, 106, 99, 211, 186, 186, 186, 
    179, 210, 200, 279, 285, 290, 283, 247, 274, 292, 250, 302, 22, 343, 268, 
    274, 284, 277, 212, 177, 294, 299, 175, 151, 160, 154, 156, 159, 148, 
    158, 169, 179, 316, 306, 295, 300, 289, 281, 294, 295, 153, 144, 67, 114, 
    56, 132, 56, 59, 70, 62, 82, 81, 60, 47, 43, 180, 239, 172, 109, 59, 246, 
    77, 224, 79, 62, 70, 56, 61, 56, 58, 51, 56, 60, 97, 188, 133, 70, 66, 
    310, 313, 30, 315, 299, 0, 136, 133, 139, 113, 141, 143, 140, 144, 134, 
    127, 131, 131, 132, 128, 131, 135, 136, 141, 266, 327, 350, 166, 146, 
    109, 294, 89, 90, 110, 115, 111, 119, 129, 123, 105, 156, 163, 120, 118, 
    147, 137, 124, 123, 106, 103, 141, 99, 95, 101, 180, 167, 168, 141, 163, 
    166, 163, 151, 112, 156, 160, 142, 121, 122, 122, 116, 100, 98, 90, 73, 
    55, 112, 19, 92, 130, 100, 94, 130, 120, 116, 125, 138, 135, 140, 136, 
    151, 150, 57, 71, 80, 203, 328, 313, 120, 30, 6, 99, 140, 166, 121, 100, 
    115, 133, 124, 115, 134, 177, 167, 156, 152, 143, 114, 89, 101, 86, 113, 
    80, 98, 89, 87, 159, 131, 150, 157, 97, 111, 134, 154, 153, 128, 147, 
    139, 126, 133, 141, 140, 155, 173, 160, 158, 200, 293, 301, 296, 305, 
    293, 297, 301, 290, 206, 245, 296, 174, 162, 153, 112, 108, 112, 104, 
    130, 136, 170, 173, 288, 273, 358, 0, 23, 6, 32, 100, 162, 133, 49, 172, 
    132, 123, 126, 148, 134, 181, 260, 299, 144, 132, 134, 114, 113, 90, 143, 
    117, 90, 89, 89, 358, 92, 92, 140, 318, 176, 81, 120, 121, 98, 106, 90, 
    174, 247, 195, 156, 233, 315, 286, 296, 295, 317, 312, 294, 303, 285, 
    290, 299, 290, 291, 270, 266, 238, 227, 234, 232, 171, 187, 235, 260, 
    295, 260, 258, 283, 270, 269, 296, 302, 280, 268, 283, 283, 296, 276, 
    324, 124, 133, 115, 111, 107, 120, 133, 123, 123, 128, 143, 263, 345, 
    259, 299, 300, 107, 31, 107, 108, 56, 124, 117, 119, 144, 147, 150, 98, 
    134, 121, 107, 118, 82, 359, 0, 297, 58, 342, 73, 94, 72, 94, 88, 91, 
    120, 97, 105, 84, 113, 100, 95, 119, 114, 111, 117, 115, 100, 96, 68, 87, 
    94, 97, 98, 99, 98, 107, 73, 105, 110, 109, 108, 113, 109, 118, 117, 110, 
    106, 111, 106, 105, 101, 101, 96, 99, 105, 115, 100, 97, 89, 94, 96, 100, 
    104, 113, 96, 96, 103, 117, 124, 106, 115, 116, 116, 116, 129, 121, 110, 
    17, 53, 123, 340, 340, 0, 12, 112, 322, 318, 343, 105, 261, 127, 70, 101, 
    57, 85, 76, 61, 47, 50, 59, 270, 346, 55, 296, 318, 232, 49, 307, 19, 
    270, 0, 0, 345, 308, 1, 360, 92, 95, 155, 92, 99, 357, 11, 150, 150, 187, 
    166, 6, 321, 72, 114, 359, 313, 214, 253, 228, 173, 233, 291, 280, 279, 
    268, 285, 270, 290, 281, 290, 290, 280, 292, 284, 285, 291, 296, 295, 
    294, 285, 296, 293, 290, 266, 287, 281, 287, 292, 278, 292, 283, 287, 
    288, 290, 294, 291, 287, 293, 281, 280, 293, 295, 297, 276, 237, 88, 83, 
    127, 122, 152, 137, 140, 133, 133, 144, 72, 76, 129, 90, 63, 307, 316, 
    298, 306, 318, 315, 4, 287, 350, 0, 128, 85, 168, 176, 173, 180, 185, 
    200, 290, 284, 276, 280, 290, 295, 317, 308, 301, 313, 316, 322, 325, 
    319, 322, 334, 92, 109, 108, 93, 50, 65, 92, 80, 69, 165, 88, 62, 255, 
    95, 110, 301, 357, 46, 0, 38, 324, 355, 307, 316, 0, 132, 127, 128, 145, 
    131, 134, 137, 156, 147, 125, 266, 289, 314, 318, 322, 335, 331, 322, 
    300, 281, 128, 81, 48, 54, 60, 194, 59, 94, 219, 247, 70, 74, 71, 81, 
    321, 326, 307, 339, 343, 333, 354, 313, 341, 304, 305, 353, 97, 98, 44, 
    176, 178, 176, 190, 177, 180, 280, 242, 312, 227, 280, 299, 312, 296, 
    269, 257, 282, 294, 202, 294, 344, 160, 165, 182, 149, 167, 126, 131, 
    178, 309, 293, 287, 215, 94, 102, 17, 275, 277, 303, 313, 283, 320, 350, 
    97, 115, 31, 297, 281, 311, 165, 49, 123, 358, 310, 295, 303, 305, 300, 
    294, 294, 295, 295, 300, 312, 323, 313, 295, 300, 277, 264, 275, 273, 
    271, 267, 262, 266, 267, 266, 264, 268, 266, 266, 276, 270, 269, 317, 
    324, 307, 332, 319, 318, 295, 330, 300, 269, 209, 271, 110, 14, 276, 284, 
    297, 178, 182, 100, 89, 113, 328, 0, 318, 315, 349, 323, 354, 17, 9, 350, 
    30, 344, 0, 143, 15, 276, 280, 264, 150, 124, 313, 37, 299, 58, 280, 56, 
    356, 40, 81, 3, 321, 21, 7, 313, 3, 288, 284, 263, 289, 285, 126, 278, 
    268, 17, 39, 324, 85, 84, 85, 84, 311, 341, 67, 313, 148, 306, 268, 322, 
    301, 357, 213, 300, 233, 34, 22, 267, 263, 22, 10, 20, 34, 26, 19, 357, 
    19, 19, 17, 47, 24, 12, 53, 277, 265, 268, 262, 293, 94, 69, 72, 75, 78, 
    80, 114, 172, 76, 276, 7, 341, 349, 360, 5, 319, 312, 350, 311, 334, 291, 
    208, 282, 279, 277, 271, 261, 351, 283, 0, 0, 267, 270, 310, 360, 72, 23, 
    342, 303, 312, 350, 0, 57, 314, 50, 355, 288, 26, 0, 285, 212, 129, 297, 
    308, 20, 295, 247, 292, 352, 336, 30, 176, 78, 65, 70, 64, 101, 325, 311, 
    310, 284, 285, 275, 271, 265, 264, 270, 294, 296, 297, 287, 264, 274, 
    241, 276, 287, 282, 275, 274, 279, 284, 290, 276, 272, 279, 280, 267, 
    263, 272, 269, 275, 268, 271, 286, 300, 335, 300, 8, 2, 350, 322, 307, 
    342, 320, 302, 298, 0, 354, 1, 147, 201, 0, 0, 342, 117, 325, 125, 334, 
    90, 99, 327, 8, 0, 360, 38, 290, 33, 332, 6, 49, 334, 278, 80, 160, 285, 
    151, 239, 127, 100, 80, 90, 102, 97, 98, 70, 71, 80, 85, 87, 54, 315, 
    301, 57, 190, 61, 60, 76, 79, 103, 120, 98, 98, 101, 111, 112, 4, 360, 
    305, 311, 343, 52, 103, 326, 346, 10, 306, 0, 111, 15, 0, 22, 249, 312, 
    156, 355, 28, 347, 0, 8, 78, 349, 0, 360, 11, 322, 0, 3, 95, 317, 318, 
    68, 323, 102, 11, 283, 6, 125, 140, 40, 103, 100, 90, 100, 120, 321, 307, 
    286, 72, 17, 5, 72, 318, 350, 320, 14, 360, 0, 60, 343, 132, 156, 272, 
    145, 87, 125, 97, 103, 83, 80, 81, 84, 98, 65, 87, 91, 82, 79, 62, 77, 
    87, 75, 73, 90, 80, 95, 91, 90, 91, 94, 92, 91, 80, 70, 107, 112, 100, 
    90, 83, 90, 94, 95, 93, 96, 98, 100, 98, 98, 99, 97, 99, 95, 91, 90, 86, 
    98, 93, 97, 100, 107, 96, 102, 93, 97, 95, 93, 95, 96, 97, 97, 109, 110, 
    98, 97, 93, 105, 104, 98, 96, 92, 89, 118, 113, 100, 75, 82, 77, 89, 80, 
    75, 86, 86, 67, 88, 91, 108, 120, 122, 106, 110, 143, 91, 126, 75, 360, 
    312, 321, 315, 329, 356, 360, 321, 25, 310, 319, 17, 340, 349, 297, 335, 
    294, 283, 135, 132, 105, 50, 43, 287, 311, 297, 307, 353, 27, 332, 314, 
    341, 344, 66, 288, 300, 98, 91, 103, 82, 111, 117, 144, 132, 110, 94, 
    340, 289, 292, 301, 329, 330, 0, 350, 25, 0, 325, 32, 328, 306, 179, 0, 
    0, 327, 67, 49, 35, 30, 25, 354, 279, 355, 350, 331, 339, 78, 322, 0, 32, 
    0, 309, 311, 351, 282, 89, 88, 6, 61, 319, 304, 279, 82, 280, 100, 93, 
    200, 282, 273, 282, 275, 292, 308, 316, 315, 317, 313, 318, 310, 295, 
    299, 295, 295, 118, 202, 273, 330, 70, 94, 61, 55, 51, 25, 244, 40, 42, 
    44, 40, 35, 33, 35, 179, 299, 232, 330, 315, 282, 342, 268, 359, 350, 
    300, 294, 300, 350, 360, 0, 358, 0, 0, 0, 309, 292, 341, 0, 0, 315, 315, 
    357, 359, 97, 308, 105, 102, 0, 273, 260, 252, 250, 0, 0, 346, 0, 0, 0, 
    4, 85, 88, 0, 0, 8, 59, 280, 289, 298, 294, 20, 130, 4, 10, 147, 341, 
    360, 0, 17, 14, 0, 344, 346, 298, 331, 340, 296, 19, 336, 337, 306, 291, 
    307, 0, 55, 280, 276, 272, 270, 271, 274, 270, 266, 276, 296, 287, 287, 
    289, 294, 310, 310, 329, 12, 15, 306, 302, 313, 3, 100, 112, 134, 126, 
    100, 49, 360, 354, 220, 349, 332, 303, 330, 92, 330, 340, 311, 330, 298, 
    111, 4, 117, 0, 327, 341, 87, 288, 300, 314, 84, 10, 8, 353, 309, 300, 
    293, 269, 264, 266, 293, 283, 254, 273, 287, 283, 280, 283, 275, 280, 
    282, 291, 307, 296, 296, 298, 293, 282, 294, 311, 297, 306, 296, 298, 
    294, 301, 310, 296, 301, 297, 317, 319, 325, 285, 342, 306, 300, 110, 
    120, 300, 320, 344, 304, 92, 83, 303, 283, 317, 282, 268, 281, 298, 296, 
    301, 288, 171, 44, 291, 316, 104, 45, 41, 301, 301, 303, 318, 122, 24, 
    23, 296, 98, 163, 99, 307, 301, 296, 103, 273, 311, 347, 0, 270, 310, 98, 
    136, 318, 360, 8, 98, 108, 349, 345, 29, 5, 344, 360, 88, 3, 113, 331, 
    320, 103, 0, 0, 20, 344, 309, 80, 54, 100, 143, 150, 302, 0, 333, 53, 1, 
    356, 86, 331, 101, 312, 61, 353, 312, 59, 316, 30, 109, 357, 43, 341, 
    360, 83, 8, 83, 302, 349, 352, 63, 316, 320, 328, 90, 353, 0, 33, 0, 56, 
    11, 0, 29, 0, 40, 355, 35, 319, 24, 360, 354, 79, 0, 344, 356, 312, 313, 
    299, 348, 315, 325, 95, 301, 353, 319, 353, 301, 350, 306, 5, 102, 350, 
    360, 84, 319, 351, 333, 353, 341, 340, 69, 346, 323, 317, 345, _, 130, 
    169, 314, 306, 323, 315, 327, 302, 331, 340, 360, 31, 314, 69, 105, 111, 
    80, 66, 60, 70, 59, 71, 1, 23, 317, 306, 119, 80, 88, 89, 100, 107, 95, 
    95, 109, 125, 124, 122, 118, 119, 119, 116, 115, 97, 81, 74, 80, 314, 
    338, 303, 316, 6, 337, 131, 85, 77, 325, 8, 20, 25, 262, 43, 6, 342, 328, 
    1, 324, 303, 323, 319, 316, 300, 303, 342, 322, 289, 294, 312, 283, 292, 
    297, 300, 326, 331, 349, 307, 344, 297, 357, 328, 351, 313, 305, 302, 
    287, 357, 307, 0, 339, 314, 301, 289, 305, 280, 339, 0, 0, 0, 85, 27, 60, 
    44, 68, 89, 0, 316, 317, 82, 0, 0, 0, 0, 0, 0, 304, 113, 66, 55, 300, 
    322, 322, 315, 257, 353, 18, 10, 355, 349, 298, 320, 304, 327, 340, 323, 
    25, 337, 360, 324, 313, 172, 49, 308, 311, 312, 0, 327, 0, 71, 0, 318, 0, 
    354, 103, 4, 97, 12, 343, 356, 293, 352, 13, 348, 317, 320, 97, 319, 315, 
    79, 309, 0, 0, 9, 0, 42, 357, 344, 58, 353, 40, 301, 359, 324, 271, 301, 
    296, 318, 288, 7, 305, 285, 50, 306, 316, _, 308, 308, 297, 326, 317, 
    308, 310, 80, 73, 252, 335, 8, 84, 72, 64, 81, 74, 84, 78, 71, 76, 73, 
    69, 71, 76, 67, 67, 48, 54, 70, 87, 61, 73, 75, 61, 68, 76, 81, 70, 76, 
    93, 94, 92, 82, 85, 83, 82, 83, 89, 86, 81, 78, 74, 73, 72, 76, 77, 74, 
    76, 83, 86, 93, 97, 84, 90, 87, 83, 89, 96, 100, 80, 95, 85, 70, 86, 102, 
    95, 80, 93, 91, 75, 75, 93, 97, 103, 83, 95, 91, 75, 82, 93, 79, 83, 80, 
    87, 90, 89, 86, 77, 77, 79, 112, 69, 53, 61, 104, 121, 123, 94, 77, 79, 
    80, 317, 283, 312, 311, 273, 288, 323, 336, 335, 70, 74, 64, 12, 334, 
    288, 191, 183, 120, 93, 95, 95, 112, 106, 111, 106, 98, 90, 92, 120, 189, 
    214, 327, 306, 293, 297, 306, 301, 299, 269, 323, 337, 296, 307, 310, 
    331, 296, 307, 312, 337, 281, 355, 336, 302, 329, 315, 311, 319, 354, 
    334, 351, 313, 329, 345, 327, 304, 283, 294, 349, 346, 0, 359, 311, 63, 
    344, 359, 13, 20, 321, 4, 325, 19, 347, 97, 307, 286, 343, 339, 324, 0, 
    0, 324, 276, 283, 275, 356, 11, 79, 79, 79, 341, 55, 7, 346, 316, 0, 338, 
    297, 63, 2, 99, 334, 25, 320, 319, 306, 289, 313, 318, 320, 292, 335, 
    346, 316, 90, 342, 345, 357, 84, 71, 350, 284, 305, 313, 296, 236, 240, 
    80, 318, 303, 316, 314, 317, 322, 308, 300, 278, 272, 283, 291, 307, 306, 
    98, 31, 329, 308, 91, 86, 50, 15, 239, 73, 89, 102, 87, 103, 115, 90, 
    201, 108, 110, 139, 344, 353, 111, 263, 25, 251, 19, 40, 42, 41, 41, 55, 
    43, 35, 47, 47, 19, 41, 118, 97, 68, 32, 290, 320, 346, 308, 300, 288, 
    298, 292, 293, 312, 331, 307, 320, 338, 298, 322, 275, 287, 300, 348, 
    277, 291, 294, 312, 296, 79, 359, 308, 285, 338, 303, 319, 288, 291, 71, 
    89, 90, 97, 108, 94, 88, 93, 85, 94, 104, 93, 90, 72, 80, 85, 91, 109, 
    45, 114, 98, 54, 163, 126, 66, 92, 110, 44, 326, 233, 188, 251, 234, 246, 
    222, 210, 206, 346, 339, 124, 140, 29, _, 274, 340, 237, 155, 126, 125, 
    33, 23, 32, 176, 97, 206, 353, 193, 201, 167, 224, 252, 96, 171, 164, 
    162, 141, 255, 21, 8, 12, 9, 21, 15, 10, 357, 7, 360, 5, 10, 14, 2, 349, 
    2, 6, 359, 348, 345, 342, 8, 1, 91, 265, 270, 294, 74, 11, 87, 312, 92, 
    272, 318, 295, 327, 325, 311, 281, 179, 268, 351, 298, 324, 307, 336, 
    340, 360, 33, 35, 178, 307, 338, 360, 332, 12, 20, 315, 358, 352, 327, 
    337, 319, 0, 318, 320, 341, 359, 40, 340, 299, 330, 304, 306, 314, 309, 
    357, 317, 310, 0, 37, 319, 323, 70, 64, 60, 49, 75, 46, 41, 45, 44, 44, 
    46, 200, 43, 50, 307, 262, 200, 18, 241, 46, 38, 31, 43, 4, 87, 239, 30, 
    42, 16, 44, 10, 18, 7, 6, 304, 302, 231, 153, 355, 353, 341, 321, 335, 
    184, 211, 332, 346, 347, 5, 11, 9, 14, 19, 54, 88, 96, 94, 95, 94, 97, 
    86, 85, 84, 89, 76, 82, 74, 87, 95, 70, 66, 149, 27, 35, 280, 248, 359, 
    11, 18, 16, 20, 24, 47, 33, 49, 57, 45, 357, 338, 83, 73, 359, 318, 343, 
    298, 0, 325, 310, 314, 348, 321, 301, 347, 338, 313, 294, 328, 331, 339, 
    301, 303, 303, 109, 62, 52, 338, 2, 344, 348, 296, 308, 318, 350, 329, 
    351, 307, 321, 320, 316, 320, 321, 322, 327, 332, 2, 319, 305, 341, 34, 
    84, 69, 109, 100, 92, 87, 94, 95, 96, 95, 93, 94, 92, 95, 98, 104, 93, 
    108, 109, 102, 103, 104, 100, 95, 88, 78, 86, 85, 93, 90, 95, 82, 86, 83, 
    92, 91, 86, 88, 88, 88, 89, 79, 80, 90, 92, 90, 82, 96, 91, 90, 73, 81, 
    69, 83, 97, 102, 83, 83, 78, 50, 49, 51, 60, 85, 96, 84, 95, 87, 80, 86, 
    86, 86, 82, 92, 70, 69, 85, 82, 85, 80, 76, 53, 66, 66, 68, 68, 67, 63, 
    67, 67, 65, 69, 69, 55, 60, 60, 68, 65, 58, 53, 43, 60, 70, 70, 56, 40, 
    212, 43, 44, 36, 53, 9, 40, 35, 360, 337, 78, 303, 296, 9, 40, 51, 327, 
    335, 234, 0, 335, 356, 295, 288, 317, 317, 319, 351, 355, 358, 298, 311, 
    17, 357, 318, 352, 331, 0, 0, 355, 360, 42, 91, 314, 54, 43, 43, 30, 49, 
    0, 9, 5, 4, 5, 33, 14, 0, 46, 8, 6, 10, 23, 40, 314, 344, 87, 92, 81, 84, 
    91, 97, 98, 78, 83, 93, 82, 73, 82, 92, 89, 80, 78, 71, 80, 102, 95, 103, 
    91, 105, 100, 70, 107, 113, 103, 106, 360, 359, 360, 100, 102, 80, 77, 
    77, 70, 75, 101, 100, 93, 100, 91, _, _, _, 101, 96, 82, 95, 92, 74, 84, 
    91, 69, 64, 50, 40, 77, 76, 66, 49, 68, 55, 49, 50, 59, 52, 65, 64, 91, 
    113, 93, 105, 81, 111, 125, 105, 104, 105, 116, 108, 115, 114, 100, 90, 
    89, 96, 75, 72, 62, 54, 68, 65, 87, 79, 82, 97, 39, 157, 48, 60, 62, 63, 
    45, 45, 46, 62, 63, 47, 44, 39, 45, 31, 41, 32, 36, 40, 78, 39, 43, 40, 
    38, 94, 95, 98, 86, 78, 80, 100, 98, 99, 103, 100, 96, 98, 95, 98, 100, 
    100, 120, 64, 50, 74, 81, 64, 76, 106, 86, 85, 81, 81, 81, 66, 48, 36, 
    62, 60, 58, 50, 62, 41, 66, 67, 67, 44, 73, 98, 85, 75, 83, 106, 83, 83, 
    85, 107, 88, 92, 87, 87, 70, 74, 77, 81, 92, 85, 80, 57, 81, 78, 100, 89, 
    99, 80, 105, 64, 81, 75, 78, 66, 76, 85, 103, 88, 102, 81, 94, 79, 76, 
    89, 87, 86, 88, 78, 68, 96, 65, 29, 71, 82, 54, 50, 39, 40, 88, 96, 90, 
    88, 89, 89, 85, 83, 95, 285, 305, 315, 295, 297, 318, 312, 326, 310, 324, 
    318, 317, 313, 334, 313, 308, 296, 286, 316, 325, 312, 328, 318, 346, 
    324, 342, 337, 336, 329, 298, 308, 308, 323, 309, 315, 300, 349, 343, 
    304, 305, 333, 330, 306, 305, 305, 319, 340, 317, 307, 317, 317, 309, 
    319, 313, 325, 348, 345, 311, 13, 33, 30, 28, 25, 21, 16, 14, 3, 5, 354, 
    36, 57, 58, 58, 15, 120, 85, 236, 72, 26, 15, 2, 120, _, 297, 307, 307, 
    317, 287, 308, 300, 316, 312, 318, 312, 268, 65, 111, 62, 23, 96, 326, 
    333, 311, 41, 60, 52, 11, 312, 347, 346, 303, 302, 332, 325, 310, 302, 
    304, 314, 312, 301, 338, 309, 321, 330, 298, 351, 315, 308, 325, 325, 
    328, 313, 300, 288, 30, 27, 113, 80, 88, 69, 96, 85, 125, 84, 79, 90, 92, 
    75, 85, 69, 44, 59, 60, 69, 65, 128, 166, 120, 299, 313, 8, 308, 310, 
    319, 299, 328, 315, 325, 308, 321, 4, 149, 260, 222, 323, 22, 25, 17, 26, 
    3, 9, 7, 17, 26, 32, 32, 32, 32, 32, 37, 28, 38, 38, 32, 13, 161, 230, 
    309, 338, 229, 249, 265, 301, 295, 100, 77, 60, 57, 40, 47, 49, 54, 54, 
    70, 43, 61, 55, 70, 59, 63, 67, 68, 56, 68, 52, 63, 67, 48, 71, 70, 74, 
    69, 62, 77, 65, 31, 60, 65, 46, 70, 48, 53, 63, 61, 79, 73, 360, 326, 
    296, 275, 356, 8, 9, 354, 248, 250, 315, 300, 292, 303, 323, 273, 247, 
    30, 78, 65, 52, 81, 322, 209, 270, 140, 43, 27, 44, 46, 46, 46, 50, 52, 
    74, 53, 77, 91, 79, 102, 89, 84, 113, 100, 76, 58, 67, 108, 92, 103, 90, 
    84, 88, 78, 70, 77, 71, 88, 62, 67, 66, 96, 113, 59, 55, 54, 84, 72, 94, 
    87, 87, 84, 88, 86, 96, 110, 94, 77, 49, 69, 69, 69, 97, 86, 61, 70, 74, 
    97, 97, 96, 95, 99, 96, 98, 48, 56, 49, 70, 81, 57, 79, 78, 80, 101, 81, 
    92, 88, 91, 74, 81, 88, 73, 84, 312, 313, 325, 305, 315, 302, 297, 293, 
    324, 340, 278, 291, 311, 311, 307, 352, 305, 0, 313, 237, 66, 70, 73, 62, 
    65, 61, 75, 68, 79, 88, 89, 91, 94, 93, 94, 105, 80, 73, 65, 106, 114, 
    70, 87, 85, 95, 82, 108, 72, 48, 43, 90, 95, 66, 81, 96, 90, 84, 87, 83, 
    74, 85, 44, 65, 65, 71, 65, 87, 98, 84, 109, 108, 107, 77, 56, 92, 46, 
    69, 40, 66, 65, 261, 324, 301, 307, 318, 329, 310, 300, 308, 35, 336, 
    298, 84, 335, 327, 314, 311, 222, 56, 43, 59, 17, 234, 52, 63, 74, 68, 
    64, 70, 50, 85, 171, 97, 115, 100, 73, 351, 76, 85, 88, 169, 95, 321, 1, 
    345, 354, 326, 323, 308, 330, 309, 293, 299, 278, 271, 315, 314, 299, 
    288, 263, 291, 302, 328, 309, 311, 309, 310, 329, 302, 300, 279, 2, 233, 
    257, 275, 240, 178, 344, 346, 321, 304, 302, 308, 257, 301, 334, 309, 
    334, 336, 300, 293, 293, 286, 82, 319, 317, 284, 319, 312, 320, 169, 167, 
    20, 54, 2, 255, 300, 352, 157, 245, 221, 293, 300, 316, 312, 311, 323, 
    315, 304, 7, 360, 294, 317, 315, 327, 318, 358, 359, 338, 306, 18, 325, 
    301, 305, 319, 325, 323, 317, 316, 301, 290, 83, 306, 298, 1, 343, 328, 
    301, 326, 315, 283, 200, 55, 100, 87, 106, 78, 82, 85, 83, 87, 87, 82, 
    88, 88, 89, 78, 66, 302, 360, 68, 360, 314, 74, 78, 326, 311, 345, 306, 
    271, 322, 36, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 291, 298, 
    350, 148, 281, 335, 9, 330, 2, 160, 328, 285, 259, 253, 213, 224, 119, 
    303, 43, 82, 64, 360, 353, 2, 354, 63, 37, 37, 52, 48, 76, 67, 358, 317, 
    329, 336, 277, 35, 2, 4, 6, 3, 260, 40, 34, 40, 48, 55, 41, 45, 48, 62, 
    47, 44, 45, 84, 69, 72, 61, 75, 57, 46, 61, 74, 67, 111, 80, 79, 99, 50, 
    296, 284, 336, 348, 330, 252, 208, 23, 294, 355, 285, 275, 40, 317, 115, 
    30, 353, 250, 60, 240, 53, 360, 331, 3, 15, 7, 11, 9, 29, 30, 33, 44, 18, 
    54, 34, 202, 166, 246, 199, 281, 359, 73, 35, 91, 42, 163, 88, 10, 7, 
    304, 350, 7, 2, 10, 276, 236, 262, 307, 297, 242, 268, 240, 162, 167, 43, 
    76, 238, 328, 360, 30, 324, 66, 11, 9, 10, 8, 9, _, 238, 313, 297, 313, 
    288, 326, 309, 321, 309, 314, 273, 302, 282, 22, 321, 295, 2, 36, 50, 
    268, 280, 283, 283, 285, 289, 312, 316, 290, 339, 4, 350, 12, 58, 17, 98, 
    17, 22, 333, 314, 320, 347, 330, 321, 308, 317, 312, 312, 309, 317, 291, 
    288, 301, 264, 280, 311, 300, 298, 307, 302, 297, 298, 336, 340, 356, 
    301, 323, 306, 312, 302, 271, 303, 314, 327, 305, 290, 325, 301, 322, 
    302, 306, 316, 323, 324, 320, 296, 330, 336, 318, 326, 320, 310, 304, 
    315, 317, 311, 304, 320, 331, 299, 325, 28, 292, 308, 302, 295, 336, 320, 
    331, 318, 340, 296, 300, 309, 320, 337, 309, 325, 316, 8, 342, 311, 302, 
    329, 333, 324, 315, 360, 314, 301, 351, 326, 303, 308, 313, 310, 301, 
    295, 306, 307, 334, 333, 298, 320, 3, 308, 346, 24, 45, 39, 133, 326, 
    245, 105, 12, 340, 283, 319, 12, 172, 175, 15, 12, 360, 324, 53, 333, 
    311, 310, 356, 338, 358, 307, 286, 293, 321, 323, 290, 309, 319, 306, 
    314, 310, 306, 311, 321, 285, 0, 324, 307, 13, 328, 329, 355, 336, 334, 
    318, 337, 359, 316, 324, 326, 330, 349, 359, 41, 306, 300, 280, 289, 310, 
    342, 328, 336, 353, 273, 7, 346, 345, 19, 50, 58, 51, 40, 49, 49, 47, 72, 
    50, 61, 62, 69, 67, 58, 51, 55, 61, 92, 120, 96, 147, 89, 79, 335, 346, 
    347, 302, 309, 309, 288, 332, 351, 313, 314, 312, 336, 337, 85, 360, 342, 
    42, 47, 44, 44, 43, 41, 42, 43, 28, 38, 43, 41, 40, 47, 357, 3, 57, 39, 
    44, 210, 221, 170, 206, 154, 71, 16, 10, 9, 324, 89, 0, 318, 278, 111, 
    351, 58, 62, 329, 347, 349, 0, 62, 335, 69, 360, 354, 324, 330, 355, 301, 
    339, 347, 25, 10, 62, 108, 88, 51, 50, 67, 292, 303, 310, 304, 355, 351, 
    284, 1, 58, 318, 360, 3, 353, 313, 66, 307, 18, 41, 0, 330, 26, 20, 298, 
    61, 69, 347, 322, 0, 0, 0, 0, 0, 0, 0, 49, 0, 309, 339, 324, 320, 321, 
    324, 324, 357, 320, 292, 15, 309, 355, 303, 92, 0, 289, 297, 107, 327, 
    332, 349, 250, 200, 135, 290, 311, 353, 73, 0, 27, 55, 304, 312, 298, 
    311, 313, 302, 347, 87, 208, 282, 318, 312, 300, 294, 0, 0, 0, 17, 293, 
    276, 266, 277, 289, 287, 277, 274, 283, 272, 278, 273, 270, 269, 269, 
    272, 270, 288, 271, 272, 273, 280, 280, 280, 277, 294, 288, 290, 343, 
    294, 338, 281, 302, 309, 302, 306, 79, 10, 22, 345, 335, 106, 0, 77, 88, 
    15, 4, 358, 103, 76, 319, 0, 8, 72, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, 313, 60, 343, 347, 43, 307, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, 281, 74, 333, 40, 59, 297, 77, 73, 
    335, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 40, 41, 31, 48, 339, 303, 
    306, 298, 288, 308, 299, 300, 304, 305, 310, 311, 282, 306, 345, 350, 19, 
    336, 343, 352, 331, 311, 320, 39, 351, 341, 312, 328, 311, 231, 66, 50, 
    78, 80, 275, 273, 67, 307, 22, 237, 346, 249, 158, 30, 148, 116, 76, 332, 
    332, 148, 305, 355, 327, 291, 243, 351, 89, 91, 1, 347, 352, 342, 303, 
    18, 222, 284, 325, 72, 339, 323, 329, 333, 8, 334, 329, 277, 327, 334, 
    336, 350, 260, 308, 360, 49, 339, 112, 88, 63, 302, 246, 279, 329, 328, 
    333, 301, 322, 318, 39, 333, 324, 49, 359, 294, 304, 315, 345, 345, 349, 
    331, 360, 1, 347, 301, 335, 298, 305, 322, 312, 51, 348, 349, 11, 28, 11, 
    25, 316, 0, 321, 86, 345, 2, 3, 360, 37, 346, 47, 38, 32, 0, 4, 318, 121, 
    308, 3, 74, 336, 326, 110, 80, 310, 335, 356, 335, 0, _, 305, 356, 321, 
    345, 71, 328, 317, 100, 304, 360, 3, 0, 81, 350, 88, 349, 35, 15, 86, 2, 
    104, 0, 50, 51, 0, 330, 345, 14, 54, 314, 328, 20, 334, 0, 41, 74, 320, 
    0, 0, 56, 0, 46, 316, 358, 100, 316, 0, 350, 340, 83, 0, 69, 357, 15, 0, 
    0, 45, 7, 0, 0, 359, 332, 81, 5, 44, 0, 25, 9, 339, 11, 0, 345, 346, 350, 
    353, 360, 2, 88, 6, 68, 317, 14, 96, 312, 356, 0, 345, 356, 353, 61, 7, 
    61, 0, 85, 86, 88, 311, 7, 86, 350, 356, 354, 56, 20, 309, 89, 328, 51, 
    10, 1, 25, 3, 83, 16, 323, 41, 345, 357, 5, 8, 325, 50, 0, 23, 10, 0, 
    321, 7, 53, 100, 9, 78, 308, 111, 348, 0, 359, 0, 21, 0, 0, 63, 14, 5, 0, 
    334, 77, 0, 343, 38, 100, 76, 351, 0, 100, 311, 50, 331, 4, 0, 330, 347, 
    0, 5, 5, 3, 360, 353, 334, 344, 75, 70, 77, 73, 337, 347, 91, 321, 48, 
    316, 0, 343, 44, 70, 347, 324, 109, 348, 330, 316, 313, 22, 335, 28, 61, 
    26, 323, 77, 360, 349, 320, 315, 89, 310, 0, 327, 121, 326, 85, 32, 50, 
    72, 0, 141, 340, 300, 21, 355, 345, 70, 332, 49, 351, 77, 299, 138, 7, 
    336, 78, 0, 17, 79, 22, 35, 324, 0, 0, 359, 360, 0, 0, 0, 0, 75, 90, 56, 
    70, 63, 91, 96, 95, 93, 90, 81, 86, 82, 92, 99, 93, 93, 90, 86, 91, 88, 
    88, 89, 83, 78, 79, 85, 82, 75, 73, 59, 67, 73, 69, 65, 59, 54, 46, 71, 
    75, 93, 61, 59, 80, 45, 328, 317, 322, 327, 325, 306, 292, 326, 62, 272, 
    278, 308, 104, 17, 351, 321, 9, 55, 357, 24, 355, 331, 352, 85, 323, 51, 
    76, 78, 359, 36, 342, 13, 40, 86, 308, 186, 200, 313, 313, 292, 316, 257, 
    296, 295, 309, 310, 316, 312, 296, 314, 327, 319, 304, 321, 322, 296, 
    286, 294, 170, 340, 230, 266, 312, 308, 322, 336, 325, 319, 112, 4, 35, 
    360, 341, 317, 62, 345, 326, 102, 359, 72, 76, 35, 304, 290, 269, 279, 
    148, 79, 66, 74, 165, 195, 52, 28, 251, 15, 14, 10, 313, 235, 360, 10, 
    52, 44, 64, 76, 142, 138, 221, 123, 70, 107, 82, 50, 51, 77, 13, 295, 
    306, 347, 7, 132, 99, 85, 63, 87, 39, 298, 291, 294, 294, 317, 49, 184, 
    176, 255, 29, 63, 76, 89, 115, 6, 349, 317, 317, 321, 0, 321, 325, 340, 
    352, 341, 285, 309, 348, 77, 345, 300, 355, 100, 66, 350, 98, 76, 310, 
    57, 322, 318, 293, 95, 75, 231, 241, 154, 336, 59, 85, 53, 42, 153, 150, 
    335, 5, 14, 73, 334, 327, 30, 10, 352, 354, 336, 309, 317, 313, 10, 20, 
    7, 297, 319, 277, 285, 66, 87, 292, 287, 338, 330, 340, 344, 0, 360, 336, 
    0, 343, 67, 330, 321, 305, 0, 18, 13, 348, 310, 139, 356, 26, 55, 71, 80, 
    129, 71, 75, 336, 347, 350, 360, 343, 356, 354, 340, 337, 326, 327, 0, 
    322, 355, 132, 297, 90, 92, 0, 118, 110, 0, 336, 320, 347, 354, 343, 29, 
    18, 53, 330, 0, 325, 85, 7, 337, 73, 346, 30, 325, 353, 108, 316, 327, 
    272, 269, 280, 297, 59, 11, 333, 358, 77, 352, 32, 346, 358, 9, 338, 353, 
    319, 348, 0, 293, 278, 273, 284, 276, _, 124, 266, 337, 249, 328, 349, 
    333, 317, 312, 307, 310, 313, 315, 100, 116, 68, 65, 65, 313, 293, 275, 
    275, 231, 354, 290, 105, 342, 117, 325, 316, 94, 32, 332, 360, 0, 0, 356, 
    17, 318, 315, 342, 87, 75, 309, 50, 135, 299, 17, 279, 356, 83, 10, 324, 
    344, 101, 307, 102, 338, 98, 356, 310, 45, 74, 60, 334, 293, 90, 354, 
    287, 263, 0, 123, 84, 360, 348, 313, 306, 312, 295, 309, 312, 310, 309, 
    307, 308, 308, 6, 44, 334, 317, 304, 301, 108, 94, 299, 32, 50, 100, 108, 
    55, 358, 92, 296, 353, 10, 337, 0, 355, 0, 312, 46, 329, 77, 117, 337, 
    283, 358, 242, 245, 0, 301, 355, 109, 300, 349, 9, 0, 8, 323, 31, 5, 318, 
    5, 347, 329, 99, 82, 351, 351, 16, 117, 259, 139, 52, 352, 360, 90, 104, 
    90, 53, 17, 326, 85, 50, 360, 329, 348, 16, 1, 337, 11, 284, 354, 318, 
    143, 24, 290, 169, 338, 123, 0, 72, 4, 0, 70, 327, 1, 123, 353, 96, 311, 
    72, 69, 9, 316, 346, 64, 339, 114, 2, 339, 357, 113, 0, 340, 302, 6, 343, 
    86, 324, 0, 62, 85, 66, 76, 52, 34, 60, 89, 352, 343, 280, 319, 140, 93, 
    342, 333, 360, 10, 284, 281, 296, 299, 309, 303, 318, 319, 67, 84, 58, 
    345, 328, 355, 107, 342, 319, 18, 67, 117, 353, 321, 330, 98, 0, 77, 94, 
    356, 319, 60, 358, 321, 315, 360, 304, 85, 332, 22, 304, 328, 288, 215, 
    284, 295, 290, 94, 314, 320, 351, 333, 33, 336, 315, 308, 339, 0, 356, 
    337, 6, 108, 110, 292, 138, 359, 357, 279, 256, 307, 300, 284, 100, 111, 
    102, 298, 298, 293, 295, 296, 307, 305, 280, 266, 306, 295, 298, 280, 
    280, 339, 307, 37, 305, 39, 319, 276, 29, 81, 111, 329, 35, 354, 345, 87, 
    330, 354, 327, 14, 8, 0, 90, 333, 306, 335, 131, 278, 16, 15, 319, 298, 
    289, 0, 331, 17, 344, 315, 315, 329, 103, 329, 359, 86, 314, 91, 331, 54, 
    347, 343, 102, 126, 316, 107, 110, 131, 360, 136, 0, 307, 305, 316, 93, 
    297, 298, 353, 344, 110, 329, 114, 308, 0, 353, 129, 74, 291, 13, 328, 
    317, 137, 355, 21, 95, 0, 0, 39, 297, 0, 6, 335, 330, 356, 314, 70, 38, 
    18, 54, 42, 136, 129, 45, 27, 75, 54, 58, 306, 52, 50, 50, 91, 119, 323, 
    38, 12, 14, 207, 237, 316, 290, 158, 338, 169, 291, 310, 288, 350, 186, 
    172, 226, 137, 177, 294, 17, 155, 5, 305, 318, 34, 28, 88, 0, 85, 311, 
    24, 108, 0, 311, 107, 0, 330, 353, 100, 339, 319, 5, 53, 0, 53, 60, 100, 
    98, 1, 322, 295, 108, 305, 63, 318, 329, 120, 344, 0, 269, 270, 171, 284, 
    325, 96, _, _, _, 129, 3, 0, 0, 346, 356, 25, 20, 8, 360, 292, 338, 339, 
    7, 350, 89, 247, 289, 274, 267, 296, 320, 320, 321, 310, 316, 317, 317, 
    93, 306, 305, 347, 70, 326, 322, 328, 8, 343, 0, 0, 59, 96, 302, 330, 
    347, 308, 351, 340, 336, 15, 0, 49, 303, 1, 305, 16, 3, 333, 0, 0, 354, 
    109, 115, 37, 59, 41, 38, 41, 43, 38, 38, 38, 47, 52, 60, 99, 292, 311, 
    350, 333, 278, 325, 290, 336, 273, 278, 274, 280, 278, 275, 275, 82, 0, 
    81, 295, 298, 300, 332, 1, 313, 335, 30, 0, 312, 336, 340, 350, 46, 105, 
    96, 259, 308, 86, 317, 347, 284, 63, 0, 336, 0, 339, 310, 307, 64, 0, 14, 
    330, 116, 315, 20, 111, 98, 351, 0, 358, 342, 0, 277, 283, 274, 11, 36, 
    20, 0, 1, 351, 330, 102, 0, 353, 6, 96, 301, 94, 319, 356, 75, 342, 0, 
    333, 256, 349, 278, 50, 42, 20, 0, 18, 306, 313, 8, 10, 46, 36, 333, 35, 
    0, 59, 309, 89, 56, 292, 285, 278, 289, 99, 114, 307, 0, 311, 14, 92, 
    329, 352, 334, 356, 331, 150, 27, 9, 315, 316, 79, 326, 319, 113, 353, 
    261, 352, 196, 107, 14, 351, 4, 360, 325, 318, 318, 341, 0, 3, 351, 301, 
    94, 131, 3, 91, 0, 237, 264, 124, 0, 282, 88, 357, 0, 137, 0, 332, 96, 
    261, 1, 0, 9, 0, 67, 0, 58, 342, 274, 120, 277, 0, 353, 64, 109, 0, 105, 
    128, 0, 288, 282, 2, 312, 107, 359, 50, 360, 17, 7, 62, 87, 65, 303, 139, 
    93, 353, 273, 49, 261, 98, 336, 293, 302, 33, 80, 118, 89, 47, 54, 47, 
    42, 346, 335, 327, 25, 103, 301, 282, 327, 276, 293, 276, 48, 97, 10, 
    325, 42, 50, 60, 77, 72, 87, 138, 113, 145, 92, 103, 121, 84, 116, 79, 
    118, 127, 60, 71, 30, 312, 310, 275, 313, 305, 300, 76, 289, 54, 68, 35, 
    25, 347, 120, 309, 348, 292, 37, 319, 64, 2, 82, 45, 99, 109, 156, 72, 
    51, 109, 151, 185, 299, 277, 301, 312, 358, 268, 310, 47, 62, 360, 0, 52, 
    307, 310, 333, 94, 94, 30, 44, 47, 286, 47, 360, 339, 168, 163, 75, 74, 
    290, 292, 286, 300, 311, 309, 283, 310, 296, 302, 290, 292, 287, 311, 
    315, 75, 116, 350, 270, 304, 273, 322, 311, 298, 47, 200, 265, 19, 273, 
    320, 298, 16, 55, 159, 65, 156, 197, 181, 281, 313, 303, 299, 306, 295, 
    306, 321, 300, 314, 334, 307, 325, 329, 95, 278, 309, 240, 314, 255, 253, 
    162, 94, 95, 98, 108, 77, 75, 70, 91, 93, 90, 60, 81, 39, 250, 73, 100, 
    88, 145, 87, 296, 180, 91, 163, 340, 91, 278, 279, 295, 289, 119, 125, 
    123, 16, 315, 0, 291, 289, 282, 3, 40, 80, 354, 0, 96, 120, 160, 89, 0, 
    90, 90, 123, 90, 162, 113, 115, 296, 133, 108, 3, 0, 0, 0, 0, 90, 94, 25, 
    351, 344, 296, 297, 305, 302, 114, 17, 327, 0, 308, 29, 325, 360, 28, 
    105, 86, 346, 311, 299, 303, 314, 128, 6, 82, 128, 306, 273, 295, 67, 4, 
    95, 286, 273, 264, 271, 258, 273, 285, 291, 289, 305, 310, 330, 42, 221, 
    20, 260, 283, 304, 272, 270, 165, 140, 156, 170, 211, 288, 181, 280, 270, 
    267, 290, 16, 303, 21, 339, 51, 353, 50, 306, 358, 142, 166, 131, 343, 
    186, 165, 157, 129, 152, 164, 198, 155, 272, 294, 200, 189, 303, 276, 
    142, 353, 297, 276, 123, 115, 261, 277, 86, 133, 121, 139, 2, 349, 86, 
    141, 254, 90, 293, 130, 0, 317, 120, 62, 83, 82, 97, 97, 103, 93, 79, 90, 
    105, 106, 108, 87, 92, 92, 95, 90, 92, 105, 85, 97, 118, 145, 93, 116, 
    135, 99, 101, 50, 30, 155, 79, 99, 111, 106, 110, 123, 135, 59, 173, 278, 
    117, 160, 152, 197, 59, 47, 50, 74, 71, 84, 70, 69, 70, 74, 83, 92, 85, 
    92, 90, 104, 88, 81, 110, 132, 95, 123, 261, 276, 299, 309, 276, 174, 
    155, 300, 337, 276, 305, 103, 140, 125, 130, 168, 148, 138, 163, 164, 
    150, 136, 119, 108, 70, 107, 60, 106, 110, 112, 108, 72, 136, 90, 93, 95, 
    97, 116, 119, 108, 110, 117, 118, 116, 119, 107, 109, 105, 94, 104, 102, 
    102, 103, 103, 110, 112, 131, 117, 121, 128, 156, 165, 151, 165, 164, 
    179, 169, 172, 172, 170, 166, 169, 174, 124, 154, 161, 130, 124, 94, 128, 
    126, 129, 125, 140, 335, 145, 164, 289, 306, 290, 268, 262, 262, 281, 
    306, 303, 292, 310, 174, 86, 88, 356, 107, 127, 353, 276, 298, 287, 290, 
    290, 286, 288, 270, 265, 159, 176, 121, 121, 66, 311, 121, 332, 116, 110, 
    109, 105, 100, 96, 113, 319, 354, 302, 213, 87, 266, 199, 126, 78, 117, 
    98, 139, 100, 82, 93, 95, 96, 50, 49, 54, 51, 48, 45, 46, 59, 53, 46, 56, 
    48, 49, 28, 27, 19, 321, 302, 329, 265, 300, 305, 285, 289, 291, 296, 
    275, 286, 269, 276, 287, 306, 247, 278, 295, 310, 264, 274, 260, 261, 
    270, 274, 300, 262, 273, 161, 111, 137, 140, 160, 163, 250, 286, 282, 
    286, 254, 129, 338, 194, 180, 47, 139, 152, 131, 109, 154, 142, 131, 152, 
    148, 130, 128, 80, 105, 113, 100, 93, 106, 107, 98, 107, 110, 88, 99, 99, 
    101, 106, 103, 106, 108, 130, 189, 136, 5, 160, 126, 12, 347, 234, 289, 
    271, 299, 130, 133, 156, 108, 111, 126, 131, 129, 155, 173, 168, 169, 
    180, 263, 258, 208, 309, 300, 200, 116, 48, 52, 114, 4, 107, 88, 355, 80, 
    134, 213, 245, 182, 142, 87, 191, 112, 107, 101, 109, 94, 79, 61, 75, 82, 
    271, 273, 293, 292, 277, 237, 98, 116, 122, 140, 131, 253, 169, 166, 166, 
    117, 146, 168, 135, 296, 295, 296, 302, 297, 261, 171, 321, 296, 298, 
    299, 271, 126, 140, 164, 122, 127, 152, 164, 130, 129, 270, 172, 300, 
    330, 301, 200, 201, 322, 323, 334, 310, 299, 299, 292, 315, 331, 185, 
    170, 117, 132, 140, 129, 129, 131, 136, 144, 134, 129, 137, 99, 130, 15, 
    132, 130, 18, 162, 137, 153, 144, 102, 179, 109, 118, 104, 104, 125, 126, 
    117, 121, 116, 102, 109, 77, 96, 9, 296, 302, 300, 292, 295, 298, 159, 
    79, 74, 84, 162, 106, 290, 45, 42, 46, 32, 39, 40, 16, 358, 356, 50, 31, 
    17, 39, 31, 35, 39, 17, 20, 56, 25, 35, 52, 47, 55, 50, 250, 39, 36, 8, 
    67, 212, 36, 20, 6, 25, 17, 103, 182, 287, 17, 6, 1, 33, 47, 70, 59, 91, 
    26, 65, 54, 45, 48, 50, 48, 51, 47, 305, 293, 293, 288, 305, 295, 283, 
    318, 79, 52, 48, 100, 286, 316, 313, 283, 300, 331, 54, 155, 130, 132, 
    277, 268, 275, 284, 289, 295, 295, 294, 291, 190, 177, 172, 166, 77, 63, 
    56, 47, 57, 60, 43, 82, 84, 114, 114, 115, 113, 109, 99, 102, 103, 98, 
    108, 100, 106, 95, 92, 102, 94, 93, 93, 89, 107, 114, 115, 113, 89, 92, 
    92, 94, 96, 97, 94, 109, 97, 95, 84, 96, 113, 96, 111, 76, 90, 75, 115, 
    102, 134, 54, 48, 16, 50, 14, 20, 39, 60, 52, 33, 34, 40, 243, 88, 68, 
    44, 112, 238, 7, 315, 68, 64, 63, 69, 163, 6, 53, 114, 138, 30, 22, 18, 
    27, 3, 22, 59, 55, 23, 79, 196, 231, 135, 149, 133, 91, 164, 154, 212, 
    182, 183, 173, 176, 180, 175, 171, 174, 172, 175, 171, 167, 290, 253, 
    293, 298, 295, 337, 188, 184, 298, 298, 277, 278, 266, 244, 287, 263, 
    271, 289, 266, 240, 263, 181, 278, 164, 216, 150, 179, 116, 193, 188, 21, 
    343, 228, 150, 121, 98, 95, 97, 97, 94, 107, 115, 126, 136, 112, 85, 108, 
    96, 94, 94, 95, 96, 109, 108, 109, 109, 315, 309, 289, 231, 124, 139, 
    131, 138, 150, 148, 146, 82, 94, 96, 70, 116, 85, 85, 82, 73, 80, 91, 
    100, 110, 82, 295, 296, 310, 288, 194, 167, 313, 309, 292, 278, 267, 264, 
    280, 283, 294, 302, 300, 290, 285, 282, 267, 269, 274, 276, 266, 260, 
    262, 260, 244, 266, 261, 236, 236, 178, 181, 163, 156, 163, 169, 0, 0, 1, 
    298, 334, 359, 270, 108, 103, 112, 114, 125, 98, 105, 84, 89, 99, 97, 96, 
    115, 126, 119, 127, 132, 129, 128, 60, 99, 141, 103, 129, 80, 108, 132, 
    124, 131, 132, 117, 130, 141, 143, 141, 130, 138, 125, 119, 50, 133, 247, 
    250, 151, 140, 128, 34, 17, 310, 254, 270, 255, 228, 157, 124, 125, 86, 
    118, 117, 132, 161, 254, 285, 300, 298, 180, 302, 123, 109, 105, 130, 
    131, 138, 145, 134, 155, 162, 146, 163, 145, 158, 138, 135, 132, 131, 
    127, 129, 131, 113, 0, 92, 37, 0, 113, 90, 91, 61, 139, 133, 133, 127, 
    125, 134, 138, 126, 117, 130, 20, 297, 132, 147, 114, 89, 116, 0, 120, 
    53, 66, 78, 81, 93, 131, 154, 82, 132, 130, 120, 130, 122, 149, 140, 136, 
    107, 139, 8, 168, 138, 87, 142, 140, 104, 0, 336, 172, 173, 162, 112, 
    156, 159, 192, 170, 174, 135, 163, 154, 176, 170, 168, 194, 161, 170, 
    115, 106, 173, 174, 101, 89, 149, 126, 125, 142, 145, 137, 128, 136, 136, 
    136, 135, 140, 158, 135, 348, 255, 186, 237, 95, 25, 350, 177, 140, 153, 
    169, 161, 283, 266, 261, 159, 116, 37, 149, 150, 150, 72, 85, 79, 124, 
    106, 84, 34, 70, 109, 92, 104, 204, 42, 146, 115, 230, 345, 52, 137, 142, 
    111, 161, 65, 105, 173, 70, 71, 328, 84, 50, 202, 30, 70, 360, 342, 331, 
    38, 335, 13, 209, 129, 40, 49, 62, 178, 170, 164, 73, 358, 50, 66, 74, 
    79, 88, 203, 73, 54, 180, 44, 91, 76, 68, 149, 50, 148, 89, 124, 131, 
    166, 156, 164, 167, 172, 138, 167, 164, 154, 154, 174, 158, 119, 148, 
    179, 164, 179, 153, 169, 166, 173, 179, 181, 168, 164, 158, 172, 159, 
    112, 125, 93, 357, 133, 357, 139, 145, 147, 140, 0, 96, 130, 121, 126, 
    125, 120, 359, 360, 88, 119, 143, 173, 150, 129, 138, 127, 121, 124, 93, 
    134, 129, 142, 162, 118, 323, 329, 354, 69, 57, 79, 83, 67, 92, 117, 115, 
    130, 134, 147, 172, 159, 141, 328, 360, 78, 307, 266, 40, 315, 219, 101, 
    136, 134, 174, 141, 165, 158, 164, 158, 159, 148, 165, 158, 171, 200, 
    317, 273, 193, 183, 166, 307, 159, 305, 107, 167, 176, 147, 67, 121, 112, 
    66, 118, 135, 61, 117, 111, 163, 174, 144, 164, 290, 274, 266, 264, 276, 
    285, 296, 153, 180, 178, 172, 170, 166, 173, 161, 157, 148, 150, 136, 
    133, 134, 140, 133, 136, 125, 167, 50, 80, 69, 81, 89, 63, 106, 279, 300, 
    142, 144, 100, 90, 107, 124, 121, 300, 299, 179, 178, 150, 117, 94, 0, 
    257, 48, 129, 359, 48, 100, 160, 92, 124, 142, 126, 173, 123, 169, 215, 
    256, 259, 253, 297, 279, 298, 292, 298, 255, 303, 315, 307, 297, 300, 
    284, 270, 289, 285, 271, 264, 253, 281, 284, 288, 296, 286, 294, 293, 
    286, 294, 296, 298, 305, 300, 302, 300, 315, 176, 131, 93, 105, 147, 333, 
    221, 250, 282, 256, 270, 295, 291, 283, 242, 285, 280, 278, 282, 286, 
    269, 280, 292, 280, 278, 282, 288, 290, 293, 289, 297, 272, 251, 243, 
    276, 296, 289, 293, 290, 290, 289, 268, 275, 255, 270, 293, 301, 281, 
    300, 299, 290, 278, 322, 282, 174, 14, 127, 172, 285, 285, 120, 300, 296, 
    281, 265, 287, 286, 271, 263, 265, 268, 269, 270, 287, 293, 293, 293, 
    279, 274, 245, 288, 267, 285, 278, 238, 240, 187, 200, 197, 183, 282, 
    163, 208, 216, 167, 157, 175, 179, 116, 125, 144, 5, 122, 156, 124, 124, 
    115, 154, 172, 172, 163, 178, 291, 175, 290, 274, 289, 294, 188, 167, 
    139, 147, 120, 154, 155, 120, 81, 104, 120, 135, 116, 111, 114, 120, 120, 
    124, 119, 114, 109, 107, 151, 316, 90, 134, 7, 160, 335, 318, 238, 166, 
    7, 150, 135, 123, 91, 112, 46, 353, 53, 55, 81, 109, 228, 258, 269, 261, 
    249, 172, 107, 62, 92, 110, 124, 105, 161, 153, 143, 167, 144, 169, 167, 
    166, 149, 132, 115, 148, 160, 162, 139, 158, 115, 129, 125, 96, 113, 131, 
    180, 27, 135, 147, 139, 130, 160, 139, 160, 154, 137, 130, 123, 126, 105, 
    126, 147, 109, 120, 83, 113, 61, 98, 59, 217, 223, 288, 107, 174, 169, 
    125, 124, 167, 120, 299, 169, 129, 128, 320, 85, 311, 301, 298, 302, 306, 
    305, 305, 307, 310, 269, 306, 95, 200, 1, 155, 0, 354, 300, 295, 171, 
    251, 168, 148, 106, 138, 60, 122, 297, 290, 287, 291, 312, 300, 299, 298, 
    302, 305, 308, 300, 289, 282, 267, 264, 287, 289, 293, 323, 321, 289, 
    289, 260, 99, 92, 137, 8, 302, 307, 164, 130, 150, 337, 127, 135, 113, 
    99, 127, 141, 131, 91, 162, 98, 93, 100, 111, 292, 261, 81, 131, 127, 
    113, 118, 123, 197, 161, 153, 151, 151, 150, 217, 90, 130, 142, 135, 137, 
    126, 92, 94, 68, 85, 75, 83, 103, 56, 92, 56, 71, 326, 289, 290, 291, 
    280, 277, 290, 286, 281, 286, 293, 293, 292, 293, 290, 295, 293, 298, 
    299, 281, 299, 298, 300, 299, 170, 175, 320, 115, 121, 35, 122, 0, 223, 
    249, 115, 309, 289, 308, 310, 322, 291, 92, 0, 340, 15, 310, 125, 357, 
    300, 287, 276, 253, 282, 264, 282, 282, 282, 255, 278, 268, 254, 271, 
    283, 294, 287, 279, 282, 267, 273, 258, 289, 270, 286, 273, 270, 267, 
    260, 259, 252, 253, 258, 268, 286, 288, 307, 336, 163, 125, 69, 289, 301, 
    294, 122, 102, 126, 54, 104, 284, 291, 297, 291, 315, 309, 293, 321, 270, 
    301, 296, 300, 316, 360, 13, 319, 326, 105, 72, 105, 136, 119, 129, 115, 
    126, 301, 132, 107, 106, 151, 160, 147, 140, 136, 110, 126, 124, 135, 
    344, 301, 292, 93, 268, 274, 7, 134, 307, 193, 132, 128, 134, 133, 133, 
    123, 106, 131, 130, 137, 130, 128, 120, 53, 0, 0, 318, 26, 132, 78, 297, 
    50, 86, 195, 153, 12, 74, 148, 136, 119, 122, 150, 129, 137, 153, 113, 
    148, 200, 299, 130, 0, 0, 117, 108, 26, 121, 33, 100, 133, 132, 148, 127, 
    123, 129, 108, 110, 131, 127, 159, 110, 348, 19, 278, 301, 33, 357, 321, 
    335, 307, 104, 104, 102, 108, 83, 148, 130, 126, 75, 89, 108, 108, 82, 
    109, 115, 255, 352, 245, 286, 358, 276, 314, 326, 47, 114, 284, 40, 355, 
    30, 20, 17, 355, 168, 130, 163, 12, 123, 135, 136, 165, 128, 318, 6, 0, 
    10, 355, 0, 92, 296, 0, 4, 93, 97, 73, 137, 120, 103, 113, 35, 110, 149, 
    114, 110, 97, 116, 270, 0, 112, 113, 267, 124, 98, 119, 120, 124, 123, 
    128, 122, 130, 134, 120, 107, 137, 135, 129, 127, 129, 130, 119, 346, 95, 
    143, 320, 306, 355, 11, 280, 233, 279, 230, 220, 200, 199, 341, 88, 121, 
    230, 169, 244, 80, 207, 53, 94, 95, 66, 199, 44, 11, 59, 13, 58, 76, 205, 
    137, 164, 76, 43, 28, 55, 74, 62, 70, 77, 100, 44, 64, 86, 100, 58, 136, 
    203, 289, 90, 80, 34, 249, 143, 189, 88, 360, 53, 82, 99, 10, 220, 298, 
    49, 236, 106, 81, 119, 122, 95, 92, 97, 82, 58, 122, 99, 94, 90, 99, 97, 
    95, 95, 67, 86, 86, 17, 105, 102, 72, 288, 295, 296, 279, 292, 264, 255, 
    94, 162, 342, 295, 111, 131, 100, 81, 91, 150, 76, 172, 165, 147, 101, 
    107, 80, 78, 103, 25, 89, 128, 114, 251, 298, 330, 307, 112, 129, 151, 
    129, 114, 106, 117, 118, 138, 142, 132, 133, 164, 121, 140, 34, 6, 56, 
    51, 56, 360, 49, 68, 62, 79, 77, 77, 261, 313, 360, 74, 62, 104, 209, 
    134, 110, 79, 92, 62, 66, 73, 77, 87, 354, 286, 270, 318, 317, 319, 355, 
    350, 41, 108, 141, 173, 69, 114, 113, 175, 214, 237, 300, 353, 236, 320, 
    337, 300, 121, 111, 0, 0, 335, 300, 315, 55, 117, 133, 127, 125, 106, 
    102, 101, 160, 155, 125, 165, 174, 169, 170, 176, 179, 171, 174, 178, 
    169, 166, 138, 51, 116, 153, 122, 122, 124, 99, 172, 128, 186, 179, 174, 
    305, 308, 322, 340, 352, 317, 344, 315, 325, 335, 310, 345, 173, 95, 128, 
    120, 126, 129, 132, 132, 105, 103, 119, 115, 104, 120, 137, 271, 177, 0, 
    0, 94, 67, 89, 81, 87, 102, 118, 128, 128, 181, 187, 155, 140, 135, 147, 
    135, 169, 135, 0, 1, 228, 326, 283, 130, 71, 55, 51, 75, 76, 214, 201, 
    143, 173, 131, 66, 161, 85, 68, 65, 2, 95, 133, 358, 142, 360, 124, 109, 
    112, 114, 112, 117, 139, 0, 150, 44, 129, 145, _, 307, 336, 0, 91, 119, 
    98, 8, 3, 0, 360, 0, 0, 14, 17, 58, 0, 0, 360, 340, 353, 0, 91, 85, 99, 
    358, 87, 64, 81, 74, 43, 50, 55, 342, 10, 110, 347, 0, 6, 321, 7, 342, 
    67, 165, 37, 33, 35, 359, 82, 23, 25, 91, 22, 78, 75, 26, 62, 45, 323, 
    13, 62, 98, 134, 24, 353, 3, 37, 359, 319, 0, 0, 140, 123, 140, 128, 101, 
    86, 72, 69, 77, 24, 306, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 120, 144, 360, 0, 10, 17, 38, 322, 0, 360, 48, 6, 4, 39, 302, 340, 
    220, 359, 0, 36, 36, 35, 45, 70, 66, 64, 58, 53, 55, 49, 48, 47, 39, 48, 
    41, 36, 46, 57, 33, 0, 0, 0, 69, 85, 122, 108, 123, 119, 120, 114, 119, 
    125, 125, 118, 110, 94, 76, 71, 46, 19, 342, 18, 109, 273, 66, 67, 231, 
    355, 360, 9, 11, 330, 4, 0, 8, 359, 27, 34, 69, 14, 316, 317, 304, 314, 
    278, 285, 358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 112, 98, 100, 86, 100, 7, 48, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 14, 15, 101, 63, 97, 143, 284, 269, 
    269, 277, 302, 273, 302, 309, 339, 332, 335, 0, 0, 0, 356, 346, 293, 278, 
    273, 284, 352, 287, 270, 282, 257, 122, 6, 0, 348, 349, 0, 352, 0, 83, 
    61, 48, 311, 320, 359, 320, 0, 344, 356, 113, 349, 360, 20, 40, 99, 62, 
    178, 193, 279, 264, 264, 256, 276, 281, 272, 285, 287, 272, 271, 283, 
    277, 278, 280, 290, 299, 291, 299, 309, 295, 271, 269, 285, 275, 294, 
    289, 301, 284, 307, 322, 335, 324, 347, 342, 358, 359, 292, 359, 354, 
    302, 0, 322, 360, 0, 0, 322, 360, 10, 0, 345, 0, 0, 39, 0, 0, 0, 0, 360, 
    0, 360, 0, 291, 320, 360, 53, 10, 4, 305, 85, 0, 0, 0, 360, 11, 0, 0, 0, 
    349, 0, 346, 0, 0, 352, 0, 60, 345, 358, 0, 29, 102, 72, 44, 30, 63, 113, 
    3, 10, 95, 360, 0, 355, 351, 0, 0, 0, 0, 360, 349, 0, 0, 0, 0, 0, 360, 
    65, 352, 179, 351, 300, 273, 311, 303, 304, 309, 312, 320, 309, 309, 320, 
    335, 300, 302, 291, 0, 0, 175, 180, 250, 281, 314, 212, 232, 286, 323, 
    304, 315, 334, 322, 318, 4, 274, 273, 277, 314, 323, 318, 341, 303, 301, 
    330, 56, 34, 63, 57, 360, 38, 81, 44, 6, 58, 359, 0, 0, 0, 348, 314, 316, 
    320, 321, 360, 0, 347, 6, 359, 295, 287, 298, 280, 277, 296, 306, 306, 
    306, 319, 328, 314, 331, 330, 337, 337, 337, 0, 0, 356, 9, 0, 0, 0, 0, 
    84, 49, 0, 0, 11, 346, 293, 302, 335, 0, 318, 314, 309, 281, 0, 0, 0, 
    304, 312, 314, 178, 277, 286, 284, 281, 283, 275, 290, 305, 272, 309, 
    301, 358, 0, 1, 0, 0, 0, 0, 0, 321, 40, 0, 322, 158, 174, 170, 73, 109, 
    99, 159, 139, 360, 176, 360, 0, 0, 0, 351, 312, 312, 0, 0, 359, 0, 354, 
    47, 90, 99, 98, 103, 106, 119, 119, 106, 111, 122, 111, 126, 115, 119, 
    123, 104, 119, 126, 114, 131, 106, 0, 90, 55, 97, 108, 106, 107, 120, 
    130, 121, 112, 123, 122, 123, 126, 135, 130, 131, 126, 118, 102, 65, 16, 
    329, 327, 0, 0, 0, 0, 350, 8, 1, 360, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 48, 43, 36, 40, 49, 42, 17, 359, 358, 66, 62, 54, 66, 74, 77, 
    67, 64, 0, 37, 0, 360, 0, 0, 328, 0, 355, 335, 352, 300, 0, 0, 326, 306, 
    301, 327, 292, 285, 0, 0, 358, 0, 359, 0, 0, 359, 0, 0, 0, 359, 360, 0, 
    4, 54, 9, 335, 344, 271, 348, 359, 26, 0, 0, 0, 342, 343, 0, 360, 360, 0, 
    309, 342, 0, 355, 68, 354, 0, 92, 103, 123, 133, 118, 126, 118, 120, 120, 
    118, 128, 118, 116, 65, 344, 359, 0, 0, 316, 0, 305, 0, 0, 345, 277, 353, 
    284, 277, 0, 299, 276, 278, 355, 0, 0, 360, 0, 357, 0, 310, 331, 339, 
    333, 0, 359, 360, 0, 356, 281, 312, 311, 355, 121, 359, 102, 101, 84, 94, 
    36, 301, 321, 316, 0, 81, 110, 100, 114, 127, 125, _, 128, 79, 102, 82, 
    110, 126, 125, _, 126, _, 121, 86, 113, 113, 80, 93, 98, 88, 66, 76, 49, 
    35, 62, 43, 45, 70, 70, 74, 63, 43, 62, 52, 60, 49, 84, 79, 84, 300, 314, 
    6, 306, 305, 350, 352, 0, 346, 241, 50, 38, 45, 60, 68, 79, 95, 354, 339, 
    8, 79, 70, 121, 86, 61, 68, 65, 46, 54, 71, 62, 62, 75, 81, 72, 74, 40, 
    87, 60, 93, 94, 118, 100, 72, 60, 56, 73, 79, 55, 61, 14, 54, 55, 33, 42, 
    355, 42, 359, 10, 2, 356, 53, 358, 6, 7, 10, 12, 2, 343, 46, 39, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 5, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, 0, 3, 22, 352, 55, 14, 52, 36, 351, 1, 0, 
    282, 318, 309, 313, 294, 308, 0, 347, 0, 318, 321, 318, 311, 321, 357, 
    327, 308, 316, 300, 319, 316, 306, 293, 310, 331, 331, 325, 321, 322, 
    302, 314, 298, 301, 315, 308, 310, 322, 313, 301, 303, 314, 297, 314, 
    311, 312, 309, 319, 318, 321, 328, 316, 342, 340, 334, 327, 342, 333, 
    324, 335, 329, 0, 0, 0, 0, 0, 0, 0, 360, 0, 0, 300, 358, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 359, 339, 0, 0, 0, 324, 326, 0, 0, 0, 0, 0, 0, 360, 0, 
    0, 0, 0, 0, 350, 0, 0, 357, 0, 0, 0, 0, 0, 0, 0, 310, 276, 166, 341, 357, 
    345, 254, 59, 24, 2, 358, 11, 9, 12, 19, 343, 319, 310, 299, 354, 277, 0, 
    0, 293, 334, 0, 18, 15, 7, 13, 360, 46, 40, 37, 37, 35, 9, 197, 349, 178, 
    266, 357, 359, 357, 356, 0, 13, 342, 0, 360, 346, 0, 357, 0, 335, 0, 64, 
    4, 0, 359, 330, 321, 0, 66, 9, 0, 0, 111, 64, 221, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 356, 0, 296, 294, 333, 343, 324, 330, 346, 0, 317, 360, 0, 
    348, 0, 0, 360, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 355, 323, 317, 0, 0, 0, 0, 0, 0, 0, 356, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 360, 0, 345, 0, 0, 0, 359, 357, 360, 0, 357, 0, 0, 354, 345, 
    360, 0, 344, 314, 332, 357, 341, 320, 325, 330, 321, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 359, 0, 0, 354, 358, 
    0, 0, 0, 0, 0, 0, 0, 0, 360, 359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 355, 0, 0, 2, 0, 0, 0, 0, 325, 339, 0, 355, 296, 332, 0, 0, 328, 0, 0, 
    345, 0, 0, 0, 0, 0, 0, 0, 360, 0, 0, 355, 0, 0, 351, 281, 280, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 342, 304, 346, 0, 0, 356, 0, 33, 0, 0, 0, 
    358, 360, 360, 347, 354, 351, 0, 347, 99, 86, 92, 98, 97, 100, 107, 109, 
    102, 101, 98, 111, 79, 98, 112, 105, 109, 113, 91, 95, 98, 88, 104, 104, 
    98, 64, 317, 279, 323, 17, 0, 353, 288, 1, 357, 342, 348, 350, 359, 359, 
    359, 315, 359, 349, 321, 348, 318, 310, 0, 0, 329, 0, 0, 0, 0, 359, 360, 
    0, 0, 359, 0, 327, 5, 0, 359, 0, 0, 25, 360, 355, 0, 0, 0, 10, 0, 360, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 321, 0, 0, 0, 309, 
    358, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 357, 0, 357, 357, 358, 
    0, 352, 0, 325, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 360, 0, 0, 0, 0, 5, 0, 
    346, 0, 0, 0, 0, 115, 78, 89, 95, 77, 82, 82, 80, 66, 98, 95, 91, 103, 
    90, 92, 94, 88, 93, 89, 96, 95, 97, 109, 102, 94, 70, 83, 80, 87, 84, 59, 
    62, 62, 83, 91, 93, 95, 98, 104, 110, 100, 101, 98, 90, 93, 92, 86, 84, 
    85, 95, 98, 90, 88, 87, 90, 81, 83, 85, 82, 86, 90, 91, 93, 96, 99, 89, 
    77, 119, 103, 82, 104, 105, 100, 86, 117, 90, 95, 79, 76, 65, 66, 69, 64, 
    69, 61, 34, 73, 72, 43, 45, 48, 54, 54, 351, 19, 82, 84, 27, 81, 76, 87, 
    11, 29, 15, 17, 94, 67, 86, 35, 91, 27, 74, 68, 79, 80, 64, 114, 28, 357, 
    1, 354, 38, 81, 33, 40, 59, 85, 87, 87, 57, 7, 83, 97, 45, 71, 35, 58, 
    46, 51, 75, 32, 43, 51, 360, 0, 360, 359, 0, 0, 8, 40, 11, 8, 0, 53, 360, 
    310, 240, 24, 167, 348, 312, 328, 360, 319, 338, 0, 336, 357, 333, 360, 
    0, 0, 0, 359, 0, 0, 353, 0, 0, 0, 342, 0, 358, 346, 0, 335, 332, 327, 0, 
    360, 0, 344, 0, 0, 342, 0, 0, 354, 329, 0, 306, 325, 330, 342, 303, 0, 
    359, 0, 0, 0, 0, 0, 0, 0, 0, 294, 289, 290, 293, 294, 301, 294, 305, 310, 
    316, 321, 323, 326, 0, 326, 0, 0, 358, 342, 357, 0, 358, 0, 0, 0, 0, 353, 
    336, 358, 288, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 360, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 360, 2, 5, 0, 0, 357, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 14, 0, 21, 38, 36, 35, 34, 29, 32, 37, 42, 48, 54, 39, 42, 
    35, 46, 43, 46, 47, 57, 72, 60, 70, 96, 80, 71, 91, 75, 78, 77, 87, 88, 
    100, 95, 89, 92, 104, _, 337, 359, 0, 1, 111, 117, 14, 354, 0, 90, 100, 
    0, 0, 98, 82, 89, 96, 91, 83, 90, 99, 110, 99, 99, 108, 105, 94, 101, 79, 
    34, 61, 114, 121, 109, 75, 103, 87, 70, 93, 51, 106, 103, 96, 93, 101, 
    103, 103, 97, 103, 113, 100, 107, 107, 99, 95, 101, 122, 123, 119, 109, 
    120, 117, 108, 106, 100, 93, 104, 97, 108, 115, 96, 93, 94, 98, 113, 96, 
    101, 104, 98, 100, 110, 120, 107, 108, 116, 111, 113, 80, 109, 105, 77, 
    80, 83, 105, 58, 211, 62, 62, 349, 288, 352, 342, 357, 355, 350, 355, 0, 
    0, 0, 0, 0, 357, 0, 348, 357, 354, 0, 0, 360, 0, 0, 355, 357, 0, 0, 0, 
    358, 0, 334, 353, 0, 360, 0, 0, 0, 0, 0, 351, 0, 314, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 360, 0, 10, 360, 0, 359, 338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 304, 
    359, 0, 0, 358, 344, 12, 359, 0, 0, 345, 360, 0, 1, 51, 311, 324, 315, 
    312, 353, 333, 0, 0, 0, 0, 303, 303, 316, 294, 273, 271, 270, 282, 313, 
    312, 289, 310, 299, 292, 292, 292, 309, 345, 352, 291, 0, 0, 333, 305, 
    317, 355, 340, 315, 307, 322, 323, 330, 334, 356, 316, 311, 306, 0, 350, 
    312, 353, 37, 345, 351, 0, 0, 360, 359, 0, 0, 346, 345, 340, 0, 0, 0, 0, 
    0, 0, 0, 293, 300, 0, 327, 356, 348, 332, 330, 345, 357, 336, 320, 296, 
    291, 351, 357, 0, 0, 359, 0, 49, 344, 0, 0, 0, 328, 330, 359, 360, 360, 
    359, 8, 44, 57, 44, 33, 43, 42, 39, 37, 34, 43, 40, 41, 41, 36, 35, 23, 
    35, 15, 42, 0, 0, 0, 353, 0, 359, 0, 0, 356, 350, 332, 341, 0, 0, 0, 0, 
    0, 359, 0, 357, 0, 358, 335, 354, 343, 0, 0, 359, 360, 297, 325, 354, 0, 
    0, 0, 326, 17, 288, 0, 0, 263, 278, 304, 307, 314, 309, 272, 275, 284, 
    273, 310, 315, 309, 284, 194, 286, 312, 312, 321, 311, 312, 305, 312, 
    299, 308, 284, 319, 260, 304, 280, 300, 300, 309, 295, 261, 307, 284, 
    286, 274, 273, 283, 290, 292, 290, 299, 309, 332, 57, 316, 117, 85, 306, 
    67, 49, 20, 8, 47, 334, 285, 289, 321, 286, 360, 2, 26, 21, 257, 289, 0, 
    301, 308, 358, 0, 45, 22, 334, 318, 298, 298, 300, 298, 0, 360, 0, 0, 0, 
    3, 352, 23, 4, 360, 199, 357, 5, 2, 72, 331, 1, 0, 0, 0, 360, 358, 356, 
    357, 345, 357, 0, 356, 339, 0, 0, 0, 0, 8, 352, 0, 0, 344, 316, 314, 327, 
    67, 79, 78, 61, 70, 95, 103, 104, 107, 102, 103, 107, 114, 121, 123, 87, 
    73, 125, 110, 114, 103, 103, 70, 104, 30, 0, 359, 355, 23, 92, 56, 0, 76, 
    358, 22, 356, 15, 43, 46, 42, 55, 43, 5, 346, 32, 53, 17, 36, 173, 30, 
    37, 46, 360, 90, 0, 0, 0, 358, 0, 353, 348, 355, 354, 7, 347, 350, 0, 0, 
    2, 0, 304, 0, 0, 359, 0, 0, 0, 0, 0, 0, 0, 0, 0, 325, 340, 360, 357, 359, 
    0, 0, 0, 0, 0, 0, 360, 0, 0, 360, 0, 0, 0, 339, 356, 360, 0, 346, 26, 86, 
    102, 95, 84, 78, 124, 129, 310, 313, 311, 300, 292, 298, 321, 330, 316, 
    338, 0, 15, 353, 291, 356, 0, 360, 0, 0, 356, 0, 345, 40, 31, 30, 13, 
    331, 29, 90, 84, 64, 117, 341, 357, 14, 1, 300, 89, 81, 61, 88, 67, 61, 
    50, 52, 50, 39, 10, 39, 41, 64, 63, 81, 41, 36, 57, 25, 42, 63, 57, 70, 
    310, 313, 43, 55, 47, 39, 43, 27, 65, 53, 48, 55, 76, 90, 99, 89, 96, 93, 
    88, 88, 105, 91, 83, 89, 91, 96, 68, 93, 101, 75, 63, 82, 83, 59, 60, 83, 
    96, 98, 92, 94, 97, 105, 48, 75, 44, 41, 26, 73, 35, 45, 41, 35, 34, 52, 
    43, 39, 38, 54, 54, 52, 86, 52, 46, 47, 34, 51, 41, 63, 116, 122, 112, 
    73, 100, 123, 84, 100, 79, 90, 100, 72, 92, 90, 99, 79, 80, 91, 83, 72, 
    96, 65, 56, 58, 102, 80, 65, 70, 72, 68, 76, 93, 68, 69, 67, 108, 114, 
    89, 89, 304, 0, 336, 314, 359, 39, 29, 325, 329, 355, 360, 75, 81, 94, 0, 
    0, 359, 0, 360, 0, 0, 0, 360, 360, 43, 0, 0, 0, 0, 0, 353, 0, 0, 0, 0, 0, 
    0, _, 0, 0, 0, 0, 0, 344, 20, 19, 35, 37, 40, 36, 39, 40, 32, 40, 44, 38, 
    25, 5, 355, 9, 2, 4, 10, 1, 7, 3, 5, 4, 15, 343, 358, 8, 11, 14, 6, 8, 
    24, 18, 10, 25, 14, 345, 352, 8, 359, 15, 10, 39, 26, 40, 30, 14, 29, 44, 
    49, 351, 344, 75, 343, 0, 1, 1, 31, 302, 8, 8, 22, 360, 23, 30, 34, 28, 
    25, 14, 314, 0, 0, 359, 353, 321, 321, 0, 8, 0, 342, 348, 15, 1, 351, 
    360, 44, 45, 42, 47, 40, 39, 41, 325, 310, 312, 310, 324, 332, 297, 278, 
    0, 0, 0, 344, 329, 292, 296, 310, 324, 0, 357, 0, 275, 299, 326, 291, 
    299, 313, 294, 288, 284, 294, 282, 286, 316, 308, 311, 312, 334, 300, 
    299, 291, 319, 358, 357, 323, 313, 334, 326, 356, 359, 0, 360, 354, 342, 
    0, 0, 350, 360, 0, 360, 0, 0, 352, 352, 299, 291, 0, 355, 302, 288, 10, 
    311, 308, 278, 276, 285, 285, 296, 301, 297, 305, 303, 285, 288, 263, 
    295, 289, 296, 312, 322, 321, 329, 2, 358, 317, 0, 0, 319, 329, 349, 294, 
    0, 0, 0, 0, 356, 357, 348, 333, 0, 55, 359, 297, 300, 310, 302, 13, 0, 0, 
    0, 0, 0, 0, 28, 0, 0, 0, 304, 318, 325, 300, 300, 287, 283, 277, 282, 
    292, 275, 279, 300, 302, 304, 311, 295, 323, 318, 0, 333, 349, 346, 0, 
    344, 314, 323, 320, 312, 280, 311, 0, 0, 339, 15, 332, 0, 2, 2, 358, 359, 
    354, 328, 0, 347, 0, 339, 343, 336, 340, 355, 12, 341, 334, 321, 341, 
    319, 339, 342, 354, 0, 350, 334, 338, 327, 354, 0, 289, 314, 292, 0, 0, 
    360, 335, 298, 8, 0, 0, 0, 0, 85, 0, 33, 360, 300, 275, 264, 262, 263, 
    259, 317, 308, 288, 273, 284, 277, 298, 308, 293, 285, 266, 278, 300, 
    289, 270, 259, 265, 287, 290, 300, 305, 291, 312, 337, 317, 0, 0, 0, 0, 
    23, 0, 327, 268, 327, 316, 319, 338, 357, 0, 0, 0, 0, 0, 322, 312, 317, 
    328, 320, 315, 314, 321, 320, 315, 322, 305, 324, 322, 318, 324, 323, 
    268, 0, 1, 349, 2, 2, 0, 0, 357, 0, 0, 72, 57, 76, 71, 50, 43, 42, 40, 8, 
    354, 37, 26, 37, 33, 37, 40, 43, 23, 18, 21, 30, 20, 28, 31, 10, 9, 10, 
    15, 5, 14, 19, 5, 46, 35, 47, 31, 213, 0, 355, 314, 352, 319, 356, 320, 
    333, 313, 313, 319, 313, 313, 313, 302, 357, 340, 340, 352, 355, 346, 
    312, 359, 320, 325, 314, 0, 0, 0, 6, 10, 17, 33, 36, 45, 46, 40, 38, 38, 
    46, 41, 36, 42, 35, 45, 40, 40, 43, 40, 29, 32, 36, 36, 35, 35, 35, 25, 
    25, 22, 21, 19, 23, 25, 36, 39, 34, 34, 34, 37, 35, 35, 40, 39, 40, 37, 
    27, 46, 46, 43, 43, 22, 339, 0, 332, 330, 327, 296, 301, 303, 307, 352, 
    0, 339, 355, 352, 0, 0, 317, 297, 341, 323, 325, 324, 323, 0, 0, 0, 25, 
    357, 19, 354, 334, 302, 305, 341, 318, 344, 342, 316, 271, 321, 315, 318, 
    0, 0, 0, 0, 18, 0, 351, 314, 87, 239, 351, 27, 146, 360, 284, 301, 298, 
    302, 311, 316, 349, 106, 318, 275, 0, 338, 320, 20, 29, 27, 338, 323, 
    302, 307, 303, 303, 325, 324, 321, 305, 0, 0, 0, 0, 342, 0, 10, 345, 331, 
    5, 24, 0, 344, 357, 293, 304, 344, 314, 6, 355, 308, 316, 356, 339, 327, 
    308, 0, 303, 339, 349, 0, 358, 0, 347, 35, 314, 323, 0, 324, 13, 12, 32, 
    346, 0, 12, 6, 290, 316, 297, 289, 299, 12, 320, 311, 300, 279, 302, 298, 
    329, 335, 307, 309, 302, 316, 334, 358, 327, 300, 305, 13, 341, 352, 0, 
    0, 350, 314, 316, 322, 325, 3, 337, 0, 0, 0, 0, 0, 0, 336, 353, 331, 0, 
    349, 344, 337, 359, 0, 0, 0, 3, 0, 0, 7, 0, 0, 0, 0, 360, 0, 0, 354, 0, 
    0, 0, 0, 357, 0, 0, 0, 0, 0, 0, 345, 0, 0, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, 99, 102, 109, 110, 103, 99, 92, 
    96, 95, 95, 90, 90, 100, 106, 111, 105, 99, 96, 98, 101, 105, 96, 97, 
    104, 103, 103, 97, 103, 100, 106, 103, 113, 119, 115, 106, 105, 104, 107, 
    82, 41, 87, 70, 73, 70, 74, 78, 73, 93, 98, 91, 100, 106, 111, 101, 109, 
    110, 107, 105, 98, 97, 108, 108, 105, 108, 100, 105, 115, 77, 86, 90, 
    142, 85, 64, 351, 0, 354, 353, 310, 330, 306, 290, 343, 314, 312, 310, 
    305, 313, 312, 57, 3, 0, 341, 322, 306, 311, 310, 318, 321, 0, 325, 0, 0, 
    0, 313, 0, 358, 0, 117, 119, 113, 96, 83, 97, 110, 92, 68, 83, 77, 57, 
    56, 65, 58, 55, 55, 55, 41, 57, 81, 76, 64, 83, 77, 254, 110, 96, 359, 
    157, 83, 65, 55, 50, 88, 71, 51, 37, 61, 41, 37, 73, 36, 64, 273, 50, 77, 
    20, 6, 360, 357, 37, 31, 43, 32, 324, 278, 330, 325, 3, 359, 356, 342, 
    333, 360, 299, 338, 45, 68, 95, 321, 304, 340, 251, 34, 33, 190, 45, 59, 
    39, 38, 38, 60, 43, 50, 51, 50, 49, 97, 354, 73, 59, 72, 0, 355, 346, 
    335, 329, 325, 339, 314, 353, 317, 322, 0, 358, 2, 328, 345, 10, 4, 359, 
    356, 0, 0, 350, 355, 356, 351, 0, 0, 1, 330, 0, 0, 0, 0, 0, 0, 348, 347, 
    341, 0, 325, 359, 359, 0, 0, 0, 0, 330, 345, 0, 333, 0, 0, 0, 347, 329, 
    352, 348, 0, 0, 0, 350, 329, 346, 0, 356, 0, 360, 0, 0, 305, 0, 358, 354, 
    90, 349, 28, 3, 8, 347, 0, 352, 334, 326, 359, 0, 30, 65, 90, 85, 347, 
    357, 348, 0, 358, 360, 349, 39, 40, 47, 335, 352, 357, 334, 8, 349, 32, 
    14, 15, 15, 14, 23, 37, 40, 37, 37, 38, 41, 38, 37, 38, 38, 29, 37, 40, 
    25, 36, 39, 357, 25, 219, 332, 336, 341, 279, 358, 0, 30, 0, 6, 0, 347, 
    0, 360, 0, 360, 0, 319, 329, 351, 356, 324, 347, 356, 351, 353, 317, 0, 
    322, 341, 0, 0, 356, 9, 352, 0, 0, 12, 359, 0, 0, 0, 0, 0, 0, 0, 356, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 340, 0, 0, 0, 345, 343, 351, 30, 0, 4, 0, 
    0, 346, 359, 0, 336, 351, 341, 4, 345, 350, 0, 305, 78, 340, 31, 0, 332, 
    0, 343, 338, 0, 0, 0, 347, 0, 0, 0, 0, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 360, 0, 0, 351, 343, 0, 354, 61, 359, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 357, 360, 0, 0, 0, 0, 0, 0, 0, 5, 359, 0, 355, 0, 352, 
    358, 360, 355, 350, 349, 0, 0, 335, 346, 0, 359, 343, 344, 319, 327, 315, 
    65, 320, 335, 355, 355, 0, 349, 0, 342, 351, 343, 344, 349, 359, 79, 71, 
    358, 0, 309, 50, 0, 358, 334, 355, 324, 360, 360, 0, 330, 4, 349, 303, 9, 
    346, 352, 78, 82, 80, 77, 76, 84, 84, 87, 96, 93, 91, 94, 108, 100, 100, 
    96, 97, 91, 88, 93, 86, 80, 76, 76, 77, 76, 52, 13, 15, 347, 81, 71, 75, 
    71, 74, 79, 79, 78, 79, 83, 77, 77, 77, 90, 81, 99, 91, 76, 71, 80, 60, 
    0, 36, 60, 4, 13, 343, 295, 302, 343, 305, 310, 341, 0, 52, 360, 360, 4, 
    0, 67, 7, 50, 57, 75, 80, 81, 72, 74, 75, 68, 84, 91, 81, 21, 322, 327, 
    0, 359, 323, 349, 328, 2, 338, 360, 1, 0, 6, 14, 333, 3, 351, 324, 0, 0, 
    5, 350, 360, 11, 17, 18, 11, 37, 0, 4, 34, 79, 104, 16, 66, 72, 80, 92, 
    121, 99, 69, 59, 0, 0, 34, 61, 106, 16, 51, 359, 5, 1, 344, 350, 359, 1, 
    5, 328, 334, 0, 0, 316, 360, 1, 3, 12, 335, 0, 0, 0, 351, 7, 355, 356, 
    43, 3, 317, 33, 353, 305, 327, 340, 0, 359, 315, 350, 345, 0, 353, 0, 0, 
    80, 359, 360, 0, 352, 0, 0, 0, 48, 0, 0, 0, 360, 0, 0, 0, 0, 0, 0, 0, 0, 
    355, 356, 360, 357, 0, 0, 358, 1, 3, 0, 314, 334, 324, 357, 299, 319, 
    292, 314, 317, 296, 354, 72, 69, 71, 67, 78, 64, 80, 83, 70, 68, 60, 58, 
    57, 52, 63, 67, 69, 74, 90, 77, 91, 85, 72, 60, 46, 29, 42, 43, 52, 43, 
    72, 36, 46, 16, 45, 314, 44, 68, 295, 46, 40, 28, 24, 20, 2, 263, 346, 
    336, 357, 353, 303, 359, 345, 47, 37, 36, 70, 94, 319, 0, 337, 340, 351, 
    0, 349, 11, 345, 1, 0, 7, 347, 358, 340, 32, 2, 352, 360, 354, 22, 318, 
    162, 153, 32, 13, 122, 38, 206, 340, 3, 347, 295, 352, 344, 0, 0, 336, 0, 
    9, 0, 0, 0, 30, 13, 13, 16, 339, 350, 358, 359, 359, 10, 12, 16, 347, 5, 
    360, 338, 352, 1, 35, 348, 22, 22, 22, 26, 37, 356, 51, 47, 42, 360, 39, 
    40, 47, 62, 62, 44, 61, 11, 16, 334, 332, 356, 345, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 353, 0, 0, 0, 0, 0, 0, 105, 344, 0, 360, 0, 0, 
    355, 0, 0, 359, 354, 358, 0, 19, 350, 0, 0, 355, 0, 0, 340, 0, 0, 0, 0, 
    0, 38, 0, 0, 356, 0, 3, 175, 0, 0, 0, 4, 41, 0, 0, 348, 340, 324, 0, 0, 
    357, 0, 14, 354, 46, 54, 43, 31, 360, 353, 343, 19, 40, 33, 36, 43, 37, 
    40, 44, 51, 49, 43, 36, 31, 23, 88, 37, 12, 5, 354, 312, 313, 289, 309, 
    314, 310, 304, 291, 300, 309, 309, 292, 297, 305, 318, 326, 272, 275, 
    285, 289, 342, 335, 349, 340, 304, 332, 3, 304, 330, 346, 4, 287, 199, 
    334, 0, 347, 0, 291, 351, 0, 5, 282, 354, 336, 353, 339, 308, 340, 326, 
    0, 318, 357, 330, 325, 343, 350, 0, 0, 319, 352, 341, 350, 357, 0, 0, 0, 
    5, 330, 354, 327, 347, 340, 349, 320, 0, 0, 0, 344, 9, 0, 349, 8, 0, 0, 
    335, 356, 63, 334, 352, 64, 360, 320, 304, 0, 9, 65, 0, 350, 360, 0, 4, 
    12, 349, 0, 0, 67, 0, 319, 0, 347, 349, 15, 0, 321, 0, 0, 0, 0, 288, 279, 
    285, 289, 275, 286, 273, 276, 282, 281, 295, 283, 260, 274, 301, 308, 
    319, 22, 360, 0, 320, 27, 12, 8, 0, 0, 0, 0, 288, 285, 306, 35, 7, 302, 
    329, 316, 329, 340, 338, 8, 0, 0, 360, 18, 30, 63, 359, 330, 328, 4, 330, 
    337, 358, 82, 358, 0, 6, 2, 57, 51, 41, 43, 42, 40, 28, 41, 54, 52, 50, 
    48, 47, 45, 40, 39, 34, 46, 46, 29, 52, 49, 33, 27, 47, 51, 52, 219, 357, 
    345, 47, 347, 345, 344, 0, 356, 345, 336, 330, 329, 0, 0, 0, 6, 0, 358, 
    0, 0, 0, 336, 81, 317, 308, 0, 349, 90, 56, 0, 3, 0, 16, 327, 0, 330, 
    343, 0, 360, 0, 0, 0, 0, 0, 337, 305, 348, 348, 330, 315, 186, 210, 347, 
    360, 19, 346, 4, 86, 15, 61, 327, 51, 13, 38, 21, 27, 47, 33, 340, 26, 
    55, 47, 32, 41, 67, 18, 30, 45, 35, 36, 36, 271, 337, 55, 22, 25, 27, 
    357, 356, 13, 263, 3, 264, 10, 31, 3, 231, 357, 71, 2, 352, 2, 196, 82, 
    52, 341, 349, 341, 354, 338, 0, 0, 353, 10, 25, 48, 48, 67, 71, 10, 80, 
    355, 341, 13, 321, 360, 120, 359, 345, 332, 286, 298, 319, 335, 346, 8, 
    35, 264, 341, 36, 26, 46, 42, 29, 33, 232, 29, 64, 40, 16, 313, 336, 99, 
    211, 359, 360, 226, 225, 225, 26, 151, 353, 183, 145, 358, 50, 29, 103, 
    73, 17, 206, 184, 249, 40, 354, 348, 28, 348, 0, 356, 0, 325, 340, 327, 
    349, 0, 44, 358, 8, 26, 2, 330, 107, 1, 295, 36, 356, 316, 36, 13, 219, 
    333, 288, 83, 189, 176, 44, 56, 115, 360, 305, 185, 210, 224, 156, 14, 
    251, 62, 23, 356, 360, 52, 93, 72, 96, 42, 352, 351, 1, 347, 277, 177, 
    355, 100, 51, 359, 0, 345, 335, 0, 12, 0, 341, 0, 312, 343, 343, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 350, 0, 0, 320, 46, 333, 335, 0, 10, 343, 
    0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 350, 10, 352, 2, 0, 314, 84, 306, 77, 
    311, 0, 313, 360, 39, 329, 358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 322, 0, 348, 62, 78, 
    16, 10, 5, 3, 0, 3, 2, 0, 355, 0, 0, 0, 0, 0, 345, 325, 3, 0, 356, 0, 0, 
    0, 0, 0, 354, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 358, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 360, 2, 0, 0, 0, 0, 336, 20, 13, 
    5, 22, 66, 19, 6, 345, 356, 0, 0, 0, 0, 358, 0, 360, 0, 352, 0, 0, 0, 
    342, 0, 33, 0, 358, 0, 0, 0, 341, 0, 0, 0, 0, 330, 83, 0, 353, 129, 0, 0, 
    350, 355, 352, 352, 0, 41, 0, 0, 0, 0, 307, 13, 354, 346, 347, 333, 360, 
    64, 45, 158, 146, 300, 282, 268, 258, 254, 267, 255, 270, 285, 246, 288, 
    306, 264, 294, 300, 279, 282, 279, 261, 268, 356, 51, 56, 54, 305, 285, 
    0, 312, 0, 16, 40, 59, 307, 86, 79, 89, 89, 86, 76, 89, 86, 88, 87, 130, 
    136, 185, 173, 197, 215, 300, 317, 310, 308, 306, 299, 306, 314, 349, 
    330, 339, 0, 0, 0, 1, 352, 0, 39, 355, 0, 344, 340, 330, 320, 0, 0, 0, 0, 
    331, 360, 7, 0, 0, 0, 81, 13, 334, 340, 351, 336, 57, 360, 82, 355, 352, 
    6, 0, 0, 349, 336, 358, 0, 2, 0, 321, 332, 326, 8, 3, 325, 48, 336, 349, 
    335, 291, 280, 270, 322, 314, 32, 41, 41, 41, 40, 40, 30, 310, 129, 326, 
    0, 332, 358, 352, 336, 24, 353, 33, 49, 67, 273, 323, 239, 101, 60, 52, 
    360, 350, 59, 57, 333, 360, 358, 11, 5, 284, 347, 341, 110, 99, 27, 106, 
    232, 51, 24, 44, 11, 40, 199, 78, 51, 52, 223, 118, 18, 331, 249, 222, 
    260, 295, 327, 226, 352, 354, 0, 0, 347, 339, 360, 58, 0, 0, 318, 322, 
    296, 301, 360, 360, 1, 360, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 360, 2, 354, 
    346, 333, 325, 360, 43, 98, 92, 93, 64, 79, 335, 54, 71, 52, 346, 329, 
    355, 88, 94, 94, 93, 97, 113, 122, 105, 111, 116, 117, 104, 104, 112, 
    105, 112, 124, 126, 134, 78, 30, 3, 6, 4, 107, 60, 49, 16, 6, 3, 10, 42, 
    45, 47, 6, 9, 33, 30, 30, 29, 42, 62, 44, 251, 231, 17, 39, 35, 38, 37, 
    18, 14, 49, 51, 72, 76, 45, 59, 200, 257, 79, 34, 308, 48, 356, 46, 88, 
    322, 26, 8, 337, 333, 12, 33, 44, 241, 296, 72, 182, 209, 36, 7, 189, 
    268, 200, 113, 355, 306, 285, 344, 239, 2, 44, 13, 244, 336, 123, 322, 
    185, 189, 35, 227, 333, 357, 358, 358, 270, 321, 334, 49, 47, 304, 13, 
    14, 69, 17, 55, 9, 14, 32, 339, 45, 0, 318, 72, 54, 54, 41, 31, 74, _, 
    188, 80, 95, 56, 357, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 358, 
    328, 55, 0, 335, 0, 310, 350, 0, 347, 0, 0, 0, 0, 0, 0, 359, 11, 360, 0, 
    0, 0, 0, 358, 0, 330, 328, 58, 0, 0, 350, 295, 294, 292, 292, 5, 321, 
    344, 0, 295, 0, 132, 277, 294, 290, 293, 292, 291, 299, 291, 290, 288, 
    293, 295, 292, 298, 293, 298, 305, 325, 331, 9, 0, 0, 305, 307, 352, 0, 
    0, 330, 0, 2, 30, 329, 340, 355, 118, 352, 87, 187, 300, 3, 34, 332, 71, 
    50, 225, 40, 280, 25, 144, 231, 351, 223, 172, 313, 35, 307, 310, 327, 
    286, 355, 312, 10, 0, 351, 341, 0, 0, 354, 0, 0, 359, 0, 0, 0, 13, 0, 0, 
    352, 0, 56, 309, 339, 0, 0, 0, 6, 360, 0, 0, 0, 0, 0, 0, 16, 359, 0, 0, 
    0, 0, 0, 355, 305, 33, 0, 348, 348, 0, 0, 0, 0, 352, 348, 0, 0, 6, 0, 0, 
    0, 1, 0, 25, 0, 0, 3, 0, 0, 341, 0, 28, 0, 279, 0, 0, 0, 0, 0, 41, 1, 
    360, 347, 332, 352, 1, 348, 346, 348, 0, 334, 78, 336, 357, 321, 78, 346, 
    354, 0, 8, 356, 356, 0, 0, 0, 19, 0, 0, 6, 0, 0, 360, 5, 324, 4, 0, 348, 
    348, 322, 330, 338, 360, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 344, 0, 0, 342, 
    352, 360, 0, 0, 0, 0, 0, 360, 351, 0, 24, 0, 2, 346, 355, 360, 0, 20, 73, 
    0, 0, 332, 65, 2, 360, 360, 357, 0, 0, 0, 311, 286, 287, 0, 360, 0, 39, 
    294, 295, 285, 284, 275, 294, 319, 339, 320, 314, 323, 322, 2, 348, 0, 
    325, 296, 299, 284, 268, 327, 336, 321, 356, 301, 338, 0, 0, 0, 0, 284, 
    275, 278, 295, 283, 308, 302, 299, 290, 288, 298, 300, 310, 299, 309, 
    292, 309, 301, 292, 284, 290, 303, 303, 304, 59, 312, 96, 93, 97, 332, 
    306, 311, 309, 305, 306, 355, 287, 296, 302, 11, 107, 307, 50, 360, 290, 
    326, 358, 330, 322, 315, 328, 307, 316, 302, 292, 300, 279, 294, 301, 
    307, 308, 310, 297, 300, 311, 319, 339, 49, 308, 292, 288, 293, 297, 309, 
    283, 275, 297, 304, 305, 304, 296, 303, 321, 310, 305, 123, 1, 0, 0, 0, 
    0, 8, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 330, 0, 328, 
    349, 312, 357, 321, 324, 310, 200, 208, 225, 31, 45, 41, 46, 42, 49, 51, 
    45, 46, 54, 50, 55, 31, 35, 49, 55, 13, 144, 34, 4, 215, 360, 32, 354, 
    325, 44, 1, 7, 344, 172, 10, 335, 300, 307, 357, 274, 273, 308, 11, 0, 
    272, 354, 92, 310, 10, 0, 320, 312, 0, 0, 0, 360, 0, 0, 0, 0, 338, 282, 
    280, 355, 0, 0, 310, 352, 255, 351, 330, 321, 355, 360, 360, 0, 0, 0, 0, 
    80, 87, 31, 0, 356, 344, 296, 326, 341, 294, 301, 325, 0, 291, 300, 313, 
    111, 339, 338, 0, 359, 0, 84, 0, 0, 359, 324, 324, 360, 67, 344, 355, 0, 
    0, 0, 0, 0, 0, 358, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 
    0, 0, 0, 0, 25, 0, 298, 295, 97, 127, 0, 0, 0, 0, 0, 284, 296, 3, 0, 0, 
    0, 0, 5, 360, 0, 0, 20, 0, 0, 0, 0, 0, 0, 348, 288, 341, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 360, 0, 0, 357, 2, 12, 3, 0, 98, 40, 8, 350, 335, 344, 
    0, 345, 0, 0, 18, 341, 0, 0, 0, 347, 269, 279, 328, 276, 322, 9, 20, 166, 
    141, 38, 38, 28, 36, 258, 214, 329, 19, 356, 86, 232, 294, 242, 340, 360, 
    24, 42, 299, 300, 58, 40, 19, 88, 72, 256, 7, 11, 6, 75, 59, 62, 259, 
    329, 343, 26, 162, 150, 133, 198, 193, 272, 36, 40, 37, 31, 92, 33, 9, 
    120, 66, 62, 69, 90, 10, 3, 4, 173, 3, 56, 55, 70, 360, 359, 168, 180, 
    124, 101, 105, 287, 242, 63, 55, 59, 67, 71, 77, 86, 88, 77, 41, 79, 52, 
    25, 14, 50, 72, 226, 34, 41, 42, 43, 24, 30, 52, 38, 2, 351, 6, 17, 22, 
    33, 59, 47, 45, 66, 57, 46, 46, 47, 47, 34, 56, 41, 44, 53, 81, 67, 15, 
    71, 53, 94, 28, 108, 4, 185, 1, 7, 315, 17, 129, 0, 340, 220, 200, 179, 
    209, 98, 161, 223, 157, 175, 355, 49, 148, 108, 89, 40, 99, 52, 6, 352, 
    84, 79, 73, 82, 99, 206, 323, 272, 277, 288, 347, 177, 174, 153, 301, 
    199, 93, 337, 326, 11, 40, 38, 42, 357, 20, 295, 170, 159, 115, 69, 88, 
    106, 88, 173, 284, 360, 65, 28, 46, 52, 39, 322, 353, 350, 360, 52, 273, 
    358, 358, 29, 38, 354, 79, 82, 77, 72, 66, 61, 56, 53, 78, 49, 42, 62, 
    73, 119, 61, 71, 77, 48, 48, 61, 55, 53, 51, 54, 59, 12, 23, 17, 9, 2, 
    10, 77, 60, 34, 42, 15, 63, 17, 335, 101, 209, 21, 327, 342, 32, 12, 323, 
    0, 212, 268, 200, 189, 267, 283, 200, 161, 175, 240, 239, 261, 281, 271, 
    310, 0, 4, 0, 0, 0, 7, 0, 0, 258, 302, 275, 272, 271, 270, 260, 123, 276, 
    0, 2, 0, 360, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 306, 301, 302, 108, 112, 
    104, 113, 121, 93, 109, 113, 107, 105, 107, 125, 113, 120, 98, 97, 100, 
    97, 100, 110, 109, 0, 339, 112, 96, 101, 82, 360, 353, 115, 110, 119, 
    114, 129, 120, 111, 90, 168, 62, 317, 337, 279, 358, 296, 300, 55, 9, 
    111, 100, 0, 4, _, 0, 116, 65, 0, 360, 107, 46, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 30, 7, 348, 250, 290, 295, _, 280, 292, 301, 303, 297, 
    297, 300, 289, 288, 294, 290, 282, 294, 314, 296, 335, 113, 349, 56, 251, 
    118, 291, 352, 119, 57, 245, 44, 0, 22, 59, 294, 296, 358, 0, 16, 322, 
    42, 309, 353, 355, 360, _, 95, 336, 308, 337, 131, 253, 333, 353, _, 0, 
    0, 0, _, 0, 359, 0, 0, 0, _, 0, 0, 0, 360, 9, 360, 0, 0, 360, 360, 4, 
    360, _, 104, 0, 0, 0, 360, 0, 1, 15, 0, 11, 279, 137, 198, 3, 262, 289, 
    236, 295, 236, 5, 30, 63, 167, 59, 36, 355, 0, 0, 0, 11, 0, 0, 0, 356, 0, 
    26, 353, 360, 36, 353, 43, 79, 75, 64, 53, 57, 57, 56, 57, 60, 66, 57, 
    54, 67, 47, 71, 75, 57, 67, 38, 85, 70, 62, 64, 77, 83, 93, 85, 82, 90, 
    106, 80, 22, 102, 33, 63, 38, 40, 26, 265, 329, 239, 262, 241, 271, 0, 
    270, 261, 268, 323, 11, 112, 111, 102, 12, 70, 40, 36, 56, 38, 179, 233, 
    283, 347, 342, 87, 91, 109, 252, 300, 79, 70, 65, 50, 45, 201, 315, 335, 
    121, 68, 74, 134, 8, 331, 27, 30, 40, 141, 248, 176, 64, 152, 250, 33, 
    47, 12, 41, 33, 41, 45, 42, 43, 38, 38, 36, 314, 63, 211, 280, 246, 351, 
    84, 360, 352, 33, 28, 18, 30, 37, 50, 28, 7, 61, 68, 47, 52, 17, 57, 83, 
    23, 357, 331, 51, 50, 11, 6, 15, 5, 30, 40, 48, 50, 54, 55, 57, 55, 49, 
    50, 43, 65, 112, 57, 99, 68, 122, 34, 84, 198, 306, 236, 354, 347, 330, 
    304, 140, 130, 102, 113, 140, 265, 242, 255, 223, 208, 151, 190, 196, 28, 
    106, 40, 36, 107, 173, 182, 240, 326, 147, 360, 340, 350, 358, 318, 88, 
    40, 250, 73, 100, 147, 51, 246, 76, 308, 245, 348, 0, 300, 355, 356, 315, 
    274, 284, 0, 2, 50, 86, 80, 0, 2, 5, 0, 3, 92, 1, 136, 112, 131, 111, 97, 
    105, 111, 110, 115, 112, 98, 102, 99, 116, 127, 103, 101, 120, 145, 90, 
    115, 101, 102, 105, 90, 121, 114, 118, 107, 88, 84, 100, 53, 64, 54, 61, 
    124, 116, 124, 123, 113, 139, 81, 120, 104, 60, 47, 100, 129, 145, 113, 
    70, 97, 351, 85, 64, 80, 90, 91, 344, 63, 65, 100, 113, 115, 118, 150, 
    164, 155, 121, 116, 130, 121, 133, 360, 110, 111, 88, 100, 332, 0, 0, 27, 
    22, 323, 200, 121, 87, 136, 173, 103, 124, 172, 151, 123, 156, 217, 80, 
    90, 181, 343, 6, 65, 56, 72, 68, 80, 101, 100, 97, 233, 200, 296, 77, 75, 
    247, 217, 283, 165, 174, 150, 143, 1, 134, 137, 328, 299, 283, 354, 360, 
    72, 53, 80, 90, 200, 297, 300, 70, 80, 108, 127, 157, 45, 156, 41, 54, 
    64, 31, 8, 76, 105, 69, 100, 42, 100, 136, 221, 360, 88, 295, 47, 51, 61, 
    68, 119, 153, 164, 137, 203, 85, 293, 283, 224, 350, 289, 304, 309, 140, 
    285, 287, 280, 278, 280, 288, 279, 278, 272, 275, 277, 270, 263, 289, 
    286, 267, 284, 283, 283, 286, 296, 293, 278, 275, 318, 289, 275, 273, 
    275, 278, 270, 269, 266, 265, 268, 264, 266, 270, 276, 273, 269, 278, 
    291, 293, 274, 274, 273, 277, 297, 287, 286, 280, 278, 300, 300, 269, 
    289, 268, 271, 272, 181, 166, 154, 76, 126, 242, 23, 132, 112, 49, 260, 
    76, 33, 36, 40, 83, 70, 66, 74, 88, 84, 88, 69, 100, 165, 120, 102, 79, 
    83, 88, 85, 254, 306, 338, 326, 335, 192, 1, 18, 20, 50, 75, 100, 161, 
    112, 155, 355, 92, 103, 58, 169, 120, 114, 110, 252, 359, 2, 53, 357, 0, 
    0, 0, 286, 300, 355, 268, 158, 160, 153, 168, 166, 169, 164, 167, 173, 
    157, 156, 151, 137, 81, 93, 132, 310, 297, 280, 297, 330, 350, 112, 158, 
    168, 162, 168, 169, 171, 161, 154, 169, 165, 162, 169, 116, 158, 164, 
    173, 60, 321, 169, 342, 115, 8, 170, 200, 294, 280, 269, 270, 270, 274, 
    252, 280, 284, 128, 119, 137, 86, 102, 88, 68, 137, 60, 59, 143, 112, 
    156, 130, 110, 172, 159, 160, 142, 158, 136, 129, 129, 127, 134, 171, 
    161, 141, 6, 1, 21, 129, 329, 354, 66, 104, 200, 115, 126, 116, 146, 165, 
    141, 356, 54, 156, 64, 18, 232, 48, 45, 314, 21, 320, 263, 19, 64, 310, 
    296, 61, 55, 52, 120, 70, 60, 313, 40, 165, 100, 80, 102, 94, 74, 177, 
    67, 66, 71, 62, 79, 45, 98, 167, 69, 184, 100, 72, 193, 123, 162, 152, 
    162, 80, 91, 156, 126, 97, 107, 111, 174, 175, 185, 47, 94, 113, 120, 
    152, 165, 114, 0, 189, 188, 187, 64, 255, 68, 90, 96, 82, 63, 75, 90, 61, 
    68, 43, 226, 357, 0, 0, 1, 92, 90, 80, 74, 100, 160, 162, 147, 148, 285, 
    234, 38, 316, 172, 73, 170, 226, 68, 71, 64, 338, 339, 309, 48, 8, 0, 21, 
    0, 34, 65, 150, 167, 167, 103, 115, 121, 119, 124, 124, 114, 120, 115, 
    122, 135, 119, 6, 348, 0, 6, 2, 133, 137, 138, 131, 134, 134, 151, 157, 
    141, 156, 176, 171, 167, 180, 170, 168, 180, 168, 146, 61, 345, 176, 155, 
    92, 100, 121, 125, 133, 136, 137, 138, 133, 134, 140, 135, 140, 122, 105, 
    130, 116, 85, 117, 175, 108, 112, 118, 93, 110, 117, 120, 149, 136, 138, 
    130, 122, 142, 159, 150, 148, 170, 164, 166, 158, 108, 129, 133, 133, 
    328, 13, 83, 17, 20, 141, 148, 134, 130, 120, 100, 97, 138, 266, 255, 
    190, 287, 275, 272, 280, 284, 310, 266, 280, 302, 308, 358, 296, 302, 
    320, 323, 299, 294, 281, 252, 289, 290, 296, 322, 329, 270, 247, 145, 
    180, 173, 179, 177, 178, 176, 176, 178, 144, 98, 294, 23, 50, 93, 90, 81, 
    19, 191, 276, 75, 88, 248, 45, 84, 319, 32, 40, 59, 76, 189, 52, 14, 62, 
    82, 104, 131, 96, 89, 90, 100, 121, 171, 72, 35, 47, 50, 46, 39, 73, 44, 
    54, 61, 50, 58, 60, 27, 59, 44, 50, 68, 52, 91, 101, 70, 55, 136, 167, 
    81, 76, 109, 61, 56, 61, 56, 153, 336, 7, _, 33, 27, 6, _, 64, 48, 81, 
    25, _, 57, 50, 53, 54, 48, 41, 65, 29, 30, _, 54, 96, 84, 107, 150, 67, 
    113, 65, 98, _, 70, 119, 71, 56, 93, 115, 98, 95, 116, 95, 115, 104, 107, 
    91, 151, 78, 74, 70, 80, 58, 47, 61, 53, 77, 51, 24, 31, 39, 31, 47, 48, 
    44, 43, 42, 32, 78, 83, 85, 61, 50, 55, 174, 60, 58, 70, 211, 80, 101, 
    61, 52, 62, 67, 71, 78, 68, 67, 269, 70, 58, 61, 256, 40, 11, 266, 254, 
    241, 211, 188, 272, 316, 275, 233, 231, 191, 230, 314, 243, 36, 7, 11, 0, 
    0, 346, 330, 328, 174, 205, 5, 0, 2, 5, 0, 0, 358, 0, 0, 0, 19, 85, 130, 
    134, 136, 124, 131, 139, 167, 139, 146, 123, 122, 126, 107, 104, 120, 
    138, 112, 102, 92, 95, 97, 97, 90, 93, 121, 111, 126, 131, 128, 35, 105, 
    114, 95, 148, 91, 96, 125, 106, 359, 115, 66, 90, 111, 325, 21, 302, 303, 
    305, 310, 0, 340, 353, 109, 337, 195, 154, 130, 127, 144, 352, 62, 88, 
    102, 345, 338, 96, 296, 0, 0, 0, 128, 129, 132, 132, 128, 119, 112, 121, 
    123, 112, 120, 134, 133, 144, 347, 0, 11, 103, 0, 156, 116, 116, 156, 7, 
    111, 125, 112, 10, 173, 349, 325, 254, 152, 32, 127, 343, 155, 10, 71, 
    83, 124, 301, 0, 59, 80, 0, 112, 115, 106, 116, 132, 135, 140, 138, 142, 
    136, 138, 138, 152, 154, 137, 337, 329, 0, 128, 322, 327, 118, 120, 120, 
    125, 130, 143, 148, 143, 126, 134, 144, 133, 138, 156, 147, 138, 139, 
    142, 140, 137, 140, 138, 142, 121, 119, 137, 130, 122, 141, 157, 157, 
    168, 160, 141, 146, 147, 132, 132, 149, 145, 159, 158, 157, 164, 359, 3, 
    300, 304, 307, 290, 252, 273, 294, 308, 296, 276, 284, 289, 291, 280, 
    264, 256, 268, 279, 276, 277, 260, 256, 254, 251, 276, 274, 280, 293, 
    316, 298, 269, 297, 299, 295, 294, 281, 279, 292, 249, 299, 332, 270, 
    243, 201, 321, 270, 293, 312, 335, 309, 340, 347, 288, 282, 187, 345, 
    180, 176, 176, 172, 165, 164, 139, 161, 177, 142, 159, 152, 176, 168, 
    154, 158, 157, 166, 174, 172, 178, 169, 175, 172, 169, 144, 149, 146, 
    157, 155, 159, 157, 148, 157, 163, 155, 161, 169, 167, 167, 164, 168, 
    168, 170, 170, 173, 150, 167, 163, 174, 190, 186, 168, 141, 176, 169, 
    186, 180, 180, 166, 166, 177, 170, 160, 164, 167, 172, 170, 174, 156, 
    122, 147, 161, 170, 166, 165, 162, 165, 169, 165, 180, 159, 129, 146, 
    128, 149, 129, 122, 147, 124, 93, 0, 0, 49, 70, 67, 60, 54, 56, 76, 74, 
    66, 124, 133, 266, 261, 265, 272, 253, 268, 279, 269, 287, 292, 271, 275, 
    286, 280, 278, 277, 291, 265, 291, 289, 313, 286, 178, 302, 177, 185, 
    318, 320, 129, 108, 38, 147, 150, 330, 330, 38, 0, 0, 133, 65, 121, 0, 
    113, 159, 146, 161, 162, 167, 172, 155, 172, 151, 153, 13, 86, 283, 299, 
    306, 294, 285, 282, 300, 272, 206, 350, 288, 247, 241, 213, 297, 323, 
    167, 266, 269, 254, 264, 275, 278, 273, 269, 256, 271, 270, 300, 316, 
    316, 319, 290, 290, 270, 288, 271, 180, 309, 166, 153, 178, 174, 169, 
    141, 110, 116, 112, 0, 356, 340, 345, 354, 0, 320, 324, 316, 325, 97, 
    172, 88, 152, 141, 142, 124, 139, 120, 124, 139, 143, 136, 105, 86, 122, 
    105, 104, 200, 226, 343, 344, 62, 57, 60, 61, 64, 115, 247, 98, 125, 360, 
    306, 124, 114, 128, 139, 124, 157, 283, 355, 360, 90, 98, 144, 122, 0, 
    138, 164, 170, 155, 132, 148, 170, 163, 162, 166, 149, 127, 129, 131, 
    131, 121, 75, 105, 0, 0, 0, 112, 3, 111, 360, 113, 125, 140, 145, 139, 
    146, 139, 139, 140, 119, 117, 167, 174, 108, 97, 173, 96, 308, 360, 2, 
    29, 101, 92, 132, 99, 80, 74, 85, 67, 81, 84, 70, 67, 237, 20, 32, 346, 
    81, 16, 335, 12, 10, 5, 356, 300, 272, 111, 111, 170, 228, 141, 210, 189, 
    150, 240, 206, 169, 69, 298, 328, 288, 290, 337, 336, 0, 5, 95, 9, 136, 
    137, 106, 118, 118, 132, 134, 114, 126, 127, 111, 121, 128, 128, 129, 
    124, 128, 130, 136, 100, 80, 115, 100, 0, 119, 115, 135, 118, 120, 125, 
    128, 114, 134, 132, 136, 90, 138, 111, 92, 111, 117, 111, 123, 81, 7, 58, 
    80, 100, 128, 134, 126, 143, 53, 132, 126, 167, 136, 182, 178, 344, 253, 
    332, 130, 84, 109, 328, 307, 301, 310, _, _, 345, 0, 99, 133, 129, 142, 
    138, 130, 148, 83, 126, 97, 99, 93, 79, 128, 176, 175, 195, 175, 322, 
    304, 322, 325, 138, 84, 117, 125, 108, 133, 129, 125, 137, 149, 143, 128, 
    132, 131, 123, 127, 140, 137, 91, 110, 115, 121, 117, 113, 110, 106, 102, 
    131, 137, 132, 133, 132, 133, 134, 125, 116, 144, 137, 88, 150, 174, 174, 
    175, 175, 179, 177, 175, 181, 183, 175, 178, 143, 182, 180, 122, 125, 
    109, 132, 139, 161, 156, 152, 153, 145, 142, 143, 33, 100, 126, _, _, _, 
    1, 0, 145, 140, 128, 139, 140, 149, 151, 142, 133, 140, 134, 118, 143, 
    173, 171, 95, 112, 131, 318, 349, 20, 85, 0, 0, 0, 1, 346, 162, 146, 150, 
    140, 130, 146, 166, 239, 261, 128, 184, 82, 84, 58, 47, 17, 13, 31, 49, 
    54, 29, 64, 92, 250, 70, 82, 97, 120, 144, 138, 123, 148, 126, 144, 173, 
    172, 147, 122, 97, 72, 80, 68, 298, 3, 47, 99, 68, 105, 150, 92, 98, 134, 
    87, 121, 81, 135, 75, 121, 133, 122, 110, 112, 6, 275, 315, 310, 304, 
    306, 343, 7, 240, 240, 48, 250, 292, 196, 56, 293, 330, 350, 16, 33, 74, 
    81, 198, 72, 65, 253, 340, 355, 359, 352, 358, 59, 72, 69, 84, 70, 82, 
    70, 51, 67, 61, 70, 73, 67, 54, 56, 45, 84, 75, 50, 56, 30, 20, 10, 35, 
    51, 68, 96, 70, 78, 56, 63, 78, 87, 70, 71, 81, 83, 57, 63, 88, 39, 203, 
    61, 51, 66, 91, 35, 341, 55, 60, 68, 8, 148, 101, 110, 124, 89, 117, 68, 
    67, 66, 47, 149, 67, 72, 126, 63, 60, 31, 40, 66, 73, 89, 326, 231, 102, 
    41, 50, 105, 66, 61, 80, 132, 152, 122, 131, 17, 284, 289, 282, 281, 293, 
    273, 289, 295, 286, 285, 285, 303, 316, 298, 313, 295, 289, 293, 277, 
    277, 264, 274, 270, 269, 290, 284, 289, 320, 15, 98, 1, 310, 347, 262, 
    351, 137, 106, 178, 180, 162, 152, 320, 181, 137, 176, 357, 69, 79, 325, 
    339, 65, 138, 10, 2, 0, 327, 355, 38, 38, 205, 73, 63, 94, 130, 149, 123, 
    136, 240, 236, 269, 296, 270, 273, 302, 288, 279, 290, 287, 293, 289, 
    297, 292, 291, 284, 276, 266, 275, 271, 293, 289, 270, 283, 291, 295, 
    298, 306, 281, 253, 301, 301, 301, 306, 315, 316, 332, 304, 300, 297, 
    272, 289, 263, 275, 272, 193, 184, 181, 15, 62, 65, 97, 95, 89, 80, 345, 
    325, 351, 0, 0, 0, 0, 112, 97, 38, 160, 127, 137, 141, 123, 119, 124, 
    113, 126, 122, 120, 81, 90, 120, 159, 212, 277, 339, 360, 316, 15, 285, 
    292, 276, 209, 173, 135, 5, 21, 13, 27, 16, 34, 35, 35, 24, 1, 33, 33, 
    33, 36, 40, 32, 360, 257, 83, 126, 164, 110, 103, 253, 192, 90, 75, 42, 
    210, 209, 360, 90, 66, 105, 3, 5, 16, 15, 13, 5, 360, 13, 346, 340, 217, 
    334, 357, 348, 228, 12, 127, 116, 143, 144, 131, 69, 62, 0, 358, 324, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 352, 78, 65, 85, 68, 330, 346, 284, 
    187, 0, 0, 0, 0, 352, 0, 0, 50, 360, 250, 200, 0, 18, 138, 134, 136, 166, 
    137, 56, 178, 257, 184, 294, 269, 274, 350, 0, 14, 358, 283, 250, 270, 
    271, 0, 200, 131, 146, 101, 121, 118, 143, 147, 353, 82, 159, 153, 0, 
    351, 298, 343, 0, 0, 309, 0, 1, 351, 97, 110, 300, 141, 115, 131, 157, 
    126, 112, 128, 121, 131, 87, 84, 359, 349, 12, 103, 91, 100, 98, 120, 
    130, 100, 350, 360, 101, 92, 102, 102, 118, 101, 101, 94, 97, 90, 86, 97, 
    94, 98, 90, 100, 118, 75, 90, 102, 100, 96, 82, 95, 88, 60, 264, 289, 
    285, 272, 237, 156, 125, 348, 302, 292, 95, 350, 358, 29, 322, 0, 0, 0, 
    0, 313, 284, 83, 11, 27, 311, 52, 9, 0, 0, 0, 0, 25, 23, 354, 324, 350, 
    360, 114, 324, 0, 328, 52, 68, 20, 70, 72, 64, 324, 84, 214, 44, 110, 
    354, 242, 63, 12, 357, 348, 109, 5, 346, 330, 332, 0, 118, 129, 100, 91, 
    300, 327, 94, 22, 105, 10, 137, 354, 154, 111, 56, 173, 115, 140, 131, 
    113, 116, 141, 109, 110, 128, 100, 86, 0, 167, 333, 285, 98, 0, 0, 143, 
    22, 0, 314, 0, 355, 0, 302, 299, 311, 320, 0, 360, 343, 285, 305, 230, 
    36, 59, 208, 126, 176, 97, 14, _, 154, 104, 131, 116, 120, 120, 123, 111, 
    121, 113, _, 123, 128, 127, 69, 70, 77, 103, 117, 112, 122, 138, 132, 131 ;
}
