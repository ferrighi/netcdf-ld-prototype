netcdf SN99880-LD {
dimensions:
	time = UNLIMITED ; // (59360 currently)
variables:
	double time(time) ;
		time:cf__standard_name = "cfsn__time" ;
		time:cf__long_name = "Time of measurement" ;
		time:cf__calendar = "standard" ;
		time:cf__units = "seconds since 1970-01-01 00:00:00 UTC" ;
		time:cf__axis = "T" ;
	double latitude ;
		latitude:cf__standard_name = "cfsn__latitude" ;
		latitude:cf__long_name = "latitude" ;
		latitude:cf__units = "degree_north" ;
	double longitude ;
		longitude:cf__standard_name = "cfsn__longitude" ;
		longitude:cf__long_name = "longitude" ;
		longitude:cf__units = "degree_east" ;
	float air_temperature_2m(time) ;
		air_temperature_2m:cf__long_name = "Air temperature" ;
		air_temperature_2m:acdd__coverage_content_type = "coordinate" ;
		air_temperature_2m:cf__standard_name = "cfsn__air_temperature" ;
		air_temperature_2m:cf__units = "K" ;
	float air_pressure_at_sea_level(time) ;
		air_pressure_at_sea_level:cf__long_name = "Air pressure at sea level" ;
		air_pressure_at_sea_level:acdd__coverage_content_type = "coordinate" ;
		air_pressure_at_sea_level:cf__standard_name = "cfsn__air_pressure_at_sea_level" ;
		air_pressure_at_sea_level:cf__units = "Pa" ;
	float air_pressure_at_sea_level_qnh(time) ;
		air_pressure_at_sea_level_qnh:cf__long_name = "Air pressure (QNH)" ;
		air_pressure_at_sea_level_qnh:acdd__coverage_content_type = "coordinate" ;
		air_pressure_at_sea_level_qnh:cf__standard_name = "cfsn__air_pressure_at_sea_level_qnh" ;
		air_pressure_at_sea_level_qnh:cf__units = "hPa" ;
	float wind_speed_10m(time) ;
		wind_speed_10m:cf__long_name = "Mean wind speed" ;
		wind_speed_10m:acdd__coverage_content_type = "coordinate" ;
		wind_speed_10m:cf__standard_name = "cfsn__wind_speed" ;
		wind_speed_10m:cf__units = "m s-1" ;
	float relative_humidity(time) ;
		relative_humidity:cf__long_name = "Relative air humidity" ;
		relative_humidity:acdd__coverage_content_type = "coordinate" ;
		relative_humidity:cf__standard_name = "cfsn__relative_humidity" ;
		relative_humidity:cf__units = "1" ;
	float surface_air_pressure_2m(time) ;
		surface_air_pressure_2m:cf__long_name = "Air pressure at station level" ;
		surface_air_pressure_2m:acdd__coverage_content_type = "coordinate" ;
		surface_air_pressure_2m:cf__standard_name = "cfsn__surface_air_pressure" ;
		surface_air_pressure_2m:cf__units = "Pa" ;
	float wind_from_direction_10m(time) ;
		wind_from_direction_10m:cf__long_name = "Wind direction" ;
		wind_from_direction_10m:acdd__coverage_content_type = "coordinate" ;
		wind_from_direction_10m:cf__standard_name = "cfsn__wind_from_direction" ;
		wind_from_direction_10m:cf__units = "degree" ;
	int prefix_list ;
		prefix_list:bald__ = "https://www.opengis.net/def/binary-array-ld/" ;
		prefix_list:rdf__ = "http://www.w3.org/1999/02/22-rdf-syntax-ns#" ;
		prefix_list:cf__ = "http://def.scitools.org.uk/CFTerms/" ;
		prefix_list:acdd__ = "http://def.scitools.org.uk/ACDD/" ;
		prefix_list:nc__ = "http://def.scitools.org.uk/NetCDF/" ;
		prefix_list:cfsn__ = "http://mmisw.org/ont/cf/parameter/" ;

// global attributes:
		:station_name = "PYRAMIDEN" ;
		:wigos_identifier = "0-20000-0-01024" ;
		:wmo_identifier = "01024" ;
		:acdd__date_created = "2019-09-03T09:58:12.415858+00:00" ;
		:acdd__Conventions = "ACDD-1.3,CF-1.6" ;
		:acdd__title = "Observations from station PYRAMIDEN SN99880" ;
		:acdd__institution = "Norwegian Meteorological Institute" ;
		:acdd__source = "Meterological surface observation via frost.met.no" ;
		:acdd__history = "https://github.com/ferrighi/netcdf-ld-prototype/blob/master/files/data-provenance-sios.ttl" ;
		:acdd__references = "" ;
		:acdd__acknowledgement = "frost.met.no" ;
		:acdd__comment = "Observations based on data from frost.met.no" ;
		:acdd__creator_email = "observasjon@met.no" ;
		:acdd__creator_name = "Norwegian Meteorological Institute" ;
		:acdd__creator_url = "https://met.no" ;
		:acdd__geospatial_bounds = "POINT(16.360300 78.655700)" ;
		:acdd__geospatial_bounds_crs = "latlon" ;
		:acdd__geospatial_lat_max = "78.655700" ;
		:acdd__geospatial_lat_min = "78.655700" ;
		:acdd__geospatial_lon_max = "16.360300" ;
		:acdd__geospatial_lon_min = "16.360300" ;
		:acdd__id = "metno_obs_SN99880" ;
		:acdd__keywords = "observations" ;
		:acdd__metadata_link = "https://oaipmh.met.no/oai/?verb=GetRecord&metadataPrefix=iso&identifier=SN99880" ;
		:acdd__summary = "Surface meteorological observations from the observation network operated by the Norwegian Meteorological Institute. Data are received and quality controlled using the local KVALOBS system. Observation stations are normally operated according to WMO requirements, although specifications are not followed on some remote stations for practical matters. Stations may have more parameters than reported in this dataset." ;
		:acdd__time_coverage_start = "2012-11-16T10:00:00" ;
		:acdd__time_coverage_end = "2019-09-03T10:00:00" ;
		:cf__featureType = "timeSeries" ;
		:bald__isPrefixedBy = "prefix_list" ;
}
